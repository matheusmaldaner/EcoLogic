library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(5119 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);
    signal layer1_outputs : std_logic_vector(5119 downto 0);
    signal layer2_outputs : std_logic_vector(5119 downto 0);
    signal layer3_outputs : std_logic_vector(5119 downto 0);
    signal layer4_outputs : std_logic_vector(5119 downto 0);
    signal layer5_outputs : std_logic_vector(5119 downto 0);
    signal layer6_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= not(inputs(255)) or (inputs(41));
    layer0_outputs(1) <= (inputs(223)) or (inputs(45));
    layer0_outputs(2) <= '1';
    layer0_outputs(3) <= '1';
    layer0_outputs(4) <= (inputs(22)) and not (inputs(237));
    layer0_outputs(5) <= not((inputs(90)) xor (inputs(1)));
    layer0_outputs(6) <= not((inputs(159)) and (inputs(82)));
    layer0_outputs(7) <= (inputs(18)) and (inputs(55));
    layer0_outputs(8) <= not(inputs(152));
    layer0_outputs(9) <= (inputs(163)) and not (inputs(142));
    layer0_outputs(10) <= not(inputs(245));
    layer0_outputs(11) <= not(inputs(40)) or (inputs(148));
    layer0_outputs(12) <= (inputs(233)) or (inputs(229));
    layer0_outputs(13) <= not((inputs(161)) or (inputs(162)));
    layer0_outputs(14) <= '1';
    layer0_outputs(15) <= '1';
    layer0_outputs(16) <= (inputs(225)) and (inputs(64));
    layer0_outputs(17) <= not((inputs(212)) or (inputs(160)));
    layer0_outputs(18) <= (inputs(99)) and not (inputs(49));
    layer0_outputs(19) <= '0';
    layer0_outputs(20) <= not((inputs(149)) xor (inputs(143)));
    layer0_outputs(21) <= not((inputs(168)) or (inputs(53)));
    layer0_outputs(22) <= not(inputs(43)) or (inputs(228));
    layer0_outputs(23) <= '1';
    layer0_outputs(24) <= (inputs(90)) and not (inputs(40));
    layer0_outputs(25) <= not(inputs(3)) or (inputs(157));
    layer0_outputs(26) <= '1';
    layer0_outputs(27) <= inputs(219);
    layer0_outputs(28) <= inputs(145);
    layer0_outputs(29) <= not((inputs(203)) or (inputs(21)));
    layer0_outputs(30) <= '1';
    layer0_outputs(31) <= '0';
    layer0_outputs(32) <= not((inputs(34)) or (inputs(60)));
    layer0_outputs(33) <= not((inputs(165)) xor (inputs(91)));
    layer0_outputs(34) <= (inputs(145)) and not (inputs(32));
    layer0_outputs(35) <= inputs(80);
    layer0_outputs(36) <= not(inputs(218)) or (inputs(58));
    layer0_outputs(37) <= '0';
    layer0_outputs(38) <= '1';
    layer0_outputs(39) <= (inputs(45)) and (inputs(246));
    layer0_outputs(40) <= not(inputs(120)) or (inputs(32));
    layer0_outputs(41) <= inputs(154);
    layer0_outputs(42) <= '0';
    layer0_outputs(43) <= (inputs(130)) and not (inputs(135));
    layer0_outputs(44) <= (inputs(230)) and not (inputs(8));
    layer0_outputs(45) <= not((inputs(47)) and (inputs(180)));
    layer0_outputs(46) <= not(inputs(172));
    layer0_outputs(47) <= (inputs(7)) and not (inputs(157));
    layer0_outputs(48) <= inputs(19);
    layer0_outputs(49) <= (inputs(143)) and not (inputs(92));
    layer0_outputs(50) <= '0';
    layer0_outputs(51) <= not(inputs(60));
    layer0_outputs(52) <= not(inputs(20)) or (inputs(117));
    layer0_outputs(53) <= not(inputs(108)) or (inputs(134));
    layer0_outputs(54) <= (inputs(149)) and (inputs(237));
    layer0_outputs(55) <= not(inputs(72));
    layer0_outputs(56) <= not(inputs(179));
    layer0_outputs(57) <= not((inputs(3)) and (inputs(146)));
    layer0_outputs(58) <= '0';
    layer0_outputs(59) <= not(inputs(69)) or (inputs(145));
    layer0_outputs(60) <= (inputs(133)) and not (inputs(208));
    layer0_outputs(61) <= (inputs(176)) and not (inputs(251));
    layer0_outputs(62) <= '0';
    layer0_outputs(63) <= not((inputs(238)) xor (inputs(194)));
    layer0_outputs(64) <= (inputs(187)) or (inputs(221));
    layer0_outputs(65) <= '1';
    layer0_outputs(66) <= (inputs(187)) or (inputs(158));
    layer0_outputs(67) <= not(inputs(26));
    layer0_outputs(68) <= not(inputs(25));
    layer0_outputs(69) <= not(inputs(212));
    layer0_outputs(70) <= (inputs(161)) or (inputs(246));
    layer0_outputs(71) <= not((inputs(185)) and (inputs(34)));
    layer0_outputs(72) <= inputs(180);
    layer0_outputs(73) <= not(inputs(251)) or (inputs(174));
    layer0_outputs(74) <= not(inputs(33)) or (inputs(12));
    layer0_outputs(75) <= not((inputs(125)) or (inputs(164)));
    layer0_outputs(76) <= (inputs(85)) xor (inputs(78));
    layer0_outputs(77) <= (inputs(113)) or (inputs(168));
    layer0_outputs(78) <= (inputs(141)) and not (inputs(236));
    layer0_outputs(79) <= '1';
    layer0_outputs(80) <= (inputs(23)) or (inputs(199));
    layer0_outputs(81) <= (inputs(193)) and not (inputs(156));
    layer0_outputs(82) <= inputs(112);
    layer0_outputs(83) <= not(inputs(26));
    layer0_outputs(84) <= '1';
    layer0_outputs(85) <= not(inputs(43));
    layer0_outputs(86) <= not(inputs(136)) or (inputs(18));
    layer0_outputs(87) <= inputs(183);
    layer0_outputs(88) <= (inputs(228)) and (inputs(133));
    layer0_outputs(89) <= not(inputs(196)) or (inputs(34));
    layer0_outputs(90) <= (inputs(223)) and not (inputs(83));
    layer0_outputs(91) <= not(inputs(75));
    layer0_outputs(92) <= not(inputs(8));
    layer0_outputs(93) <= (inputs(46)) and (inputs(159));
    layer0_outputs(94) <= (inputs(29)) or (inputs(5));
    layer0_outputs(95) <= '0';
    layer0_outputs(96) <= not(inputs(161)) or (inputs(39));
    layer0_outputs(97) <= (inputs(27)) and (inputs(119));
    layer0_outputs(98) <= not(inputs(174));
    layer0_outputs(99) <= not((inputs(53)) xor (inputs(46)));
    layer0_outputs(100) <= not(inputs(158)) or (inputs(31));
    layer0_outputs(101) <= not((inputs(108)) and (inputs(181)));
    layer0_outputs(102) <= not(inputs(153));
    layer0_outputs(103) <= (inputs(71)) xor (inputs(32));
    layer0_outputs(104) <= not(inputs(234));
    layer0_outputs(105) <= (inputs(233)) and not (inputs(202));
    layer0_outputs(106) <= not(inputs(37));
    layer0_outputs(107) <= not(inputs(149));
    layer0_outputs(108) <= inputs(227);
    layer0_outputs(109) <= not(inputs(254)) or (inputs(133));
    layer0_outputs(110) <= (inputs(39)) or (inputs(221));
    layer0_outputs(111) <= (inputs(163)) or (inputs(238));
    layer0_outputs(112) <= not(inputs(121));
    layer0_outputs(113) <= '1';
    layer0_outputs(114) <= not(inputs(211));
    layer0_outputs(115) <= not((inputs(31)) xor (inputs(73)));
    layer0_outputs(116) <= (inputs(170)) or (inputs(235));
    layer0_outputs(117) <= inputs(137);
    layer0_outputs(118) <= not(inputs(140)) or (inputs(43));
    layer0_outputs(119) <= not(inputs(26)) or (inputs(229));
    layer0_outputs(120) <= not((inputs(157)) or (inputs(117)));
    layer0_outputs(121) <= (inputs(147)) and not (inputs(12));
    layer0_outputs(122) <= not((inputs(248)) or (inputs(89)));
    layer0_outputs(123) <= (inputs(41)) and (inputs(9));
    layer0_outputs(124) <= not(inputs(135));
    layer0_outputs(125) <= not((inputs(193)) or (inputs(33)));
    layer0_outputs(126) <= '1';
    layer0_outputs(127) <= not((inputs(212)) and (inputs(186)));
    layer0_outputs(128) <= (inputs(24)) and not (inputs(114));
    layer0_outputs(129) <= '1';
    layer0_outputs(130) <= '0';
    layer0_outputs(131) <= not(inputs(18)) or (inputs(248));
    layer0_outputs(132) <= '0';
    layer0_outputs(133) <= not(inputs(70));
    layer0_outputs(134) <= not(inputs(216));
    layer0_outputs(135) <= '1';
    layer0_outputs(136) <= '0';
    layer0_outputs(137) <= not((inputs(16)) and (inputs(172)));
    layer0_outputs(138) <= (inputs(213)) and (inputs(141));
    layer0_outputs(139) <= (inputs(58)) and (inputs(54));
    layer0_outputs(140) <= '0';
    layer0_outputs(141) <= not(inputs(63)) or (inputs(26));
    layer0_outputs(142) <= (inputs(165)) and not (inputs(51));
    layer0_outputs(143) <= (inputs(148)) or (inputs(101));
    layer0_outputs(144) <= not(inputs(88));
    layer0_outputs(145) <= not((inputs(164)) or (inputs(141)));
    layer0_outputs(146) <= '1';
    layer0_outputs(147) <= (inputs(108)) and not (inputs(106));
    layer0_outputs(148) <= inputs(177);
    layer0_outputs(149) <= inputs(45);
    layer0_outputs(150) <= (inputs(24)) and not (inputs(114));
    layer0_outputs(151) <= (inputs(83)) and not (inputs(16));
    layer0_outputs(152) <= inputs(202);
    layer0_outputs(153) <= not((inputs(157)) or (inputs(181)));
    layer0_outputs(154) <= inputs(103);
    layer0_outputs(155) <= not(inputs(166));
    layer0_outputs(156) <= not(inputs(238));
    layer0_outputs(157) <= (inputs(186)) and not (inputs(27));
    layer0_outputs(158) <= inputs(25);
    layer0_outputs(159) <= inputs(39);
    layer0_outputs(160) <= '0';
    layer0_outputs(161) <= '1';
    layer0_outputs(162) <= not((inputs(90)) or (inputs(59)));
    layer0_outputs(163) <= not((inputs(24)) and (inputs(232)));
    layer0_outputs(164) <= inputs(231);
    layer0_outputs(165) <= '0';
    layer0_outputs(166) <= '0';
    layer0_outputs(167) <= (inputs(139)) xor (inputs(194));
    layer0_outputs(168) <= (inputs(217)) and (inputs(223));
    layer0_outputs(169) <= '1';
    layer0_outputs(170) <= (inputs(234)) and (inputs(74));
    layer0_outputs(171) <= inputs(187);
    layer0_outputs(172) <= not(inputs(211));
    layer0_outputs(173) <= '0';
    layer0_outputs(174) <= not(inputs(119));
    layer0_outputs(175) <= not((inputs(85)) or (inputs(27)));
    layer0_outputs(176) <= not(inputs(172)) or (inputs(198));
    layer0_outputs(177) <= inputs(186);
    layer0_outputs(178) <= inputs(161);
    layer0_outputs(179) <= not(inputs(149));
    layer0_outputs(180) <= not(inputs(13));
    layer0_outputs(181) <= not(inputs(251)) or (inputs(96));
    layer0_outputs(182) <= not(inputs(183)) or (inputs(46));
    layer0_outputs(183) <= not(inputs(142));
    layer0_outputs(184) <= (inputs(58)) and (inputs(47));
    layer0_outputs(185) <= '1';
    layer0_outputs(186) <= not((inputs(235)) or (inputs(213)));
    layer0_outputs(187) <= '1';
    layer0_outputs(188) <= inputs(77);
    layer0_outputs(189) <= not(inputs(16));
    layer0_outputs(190) <= inputs(30);
    layer0_outputs(191) <= not(inputs(184));
    layer0_outputs(192) <= (inputs(99)) and not (inputs(247));
    layer0_outputs(193) <= inputs(164);
    layer0_outputs(194) <= not((inputs(229)) and (inputs(44)));
    layer0_outputs(195) <= not(inputs(118)) or (inputs(108));
    layer0_outputs(196) <= not((inputs(210)) and (inputs(188)));
    layer0_outputs(197) <= not(inputs(191)) or (inputs(190));
    layer0_outputs(198) <= '0';
    layer0_outputs(199) <= (inputs(163)) or (inputs(33));
    layer0_outputs(200) <= '0';
    layer0_outputs(201) <= not(inputs(59)) or (inputs(173));
    layer0_outputs(202) <= not((inputs(64)) or (inputs(88)));
    layer0_outputs(203) <= (inputs(84)) or (inputs(229));
    layer0_outputs(204) <= (inputs(132)) and not (inputs(64));
    layer0_outputs(205) <= (inputs(163)) and (inputs(108));
    layer0_outputs(206) <= inputs(217);
    layer0_outputs(207) <= inputs(230);
    layer0_outputs(208) <= (inputs(42)) and not (inputs(93));
    layer0_outputs(209) <= not(inputs(113)) or (inputs(14));
    layer0_outputs(210) <= '0';
    layer0_outputs(211) <= not(inputs(151));
    layer0_outputs(212) <= (inputs(194)) and (inputs(146));
    layer0_outputs(213) <= not(inputs(131)) or (inputs(199));
    layer0_outputs(214) <= not((inputs(48)) or (inputs(148)));
    layer0_outputs(215) <= not(inputs(1)) or (inputs(112));
    layer0_outputs(216) <= inputs(144);
    layer0_outputs(217) <= inputs(106);
    layer0_outputs(218) <= '1';
    layer0_outputs(219) <= (inputs(28)) or (inputs(113));
    layer0_outputs(220) <= not(inputs(187));
    layer0_outputs(221) <= (inputs(57)) and not (inputs(132));
    layer0_outputs(222) <= not((inputs(203)) or (inputs(234)));
    layer0_outputs(223) <= not((inputs(160)) xor (inputs(6)));
    layer0_outputs(224) <= (inputs(136)) and not (inputs(53));
    layer0_outputs(225) <= '0';
    layer0_outputs(226) <= not(inputs(185)) or (inputs(152));
    layer0_outputs(227) <= (inputs(150)) xor (inputs(227));
    layer0_outputs(228) <= '1';
    layer0_outputs(229) <= '1';
    layer0_outputs(230) <= not(inputs(84));
    layer0_outputs(231) <= not(inputs(166)) or (inputs(144));
    layer0_outputs(232) <= (inputs(38)) and not (inputs(204));
    layer0_outputs(233) <= (inputs(94)) and not (inputs(139));
    layer0_outputs(234) <= (inputs(191)) or (inputs(16));
    layer0_outputs(235) <= (inputs(6)) or (inputs(22));
    layer0_outputs(236) <= inputs(207);
    layer0_outputs(237) <= '0';
    layer0_outputs(238) <= not(inputs(184));
    layer0_outputs(239) <= not(inputs(6));
    layer0_outputs(240) <= inputs(74);
    layer0_outputs(241) <= not(inputs(3));
    layer0_outputs(242) <= inputs(1);
    layer0_outputs(243) <= inputs(228);
    layer0_outputs(244) <= not(inputs(19)) or (inputs(24));
    layer0_outputs(245) <= '1';
    layer0_outputs(246) <= '1';
    layer0_outputs(247) <= not(inputs(189));
    layer0_outputs(248) <= '1';
    layer0_outputs(249) <= not(inputs(243)) or (inputs(215));
    layer0_outputs(250) <= (inputs(132)) and (inputs(228));
    layer0_outputs(251) <= (inputs(140)) or (inputs(89));
    layer0_outputs(252) <= not(inputs(26)) or (inputs(230));
    layer0_outputs(253) <= '1';
    layer0_outputs(254) <= (inputs(105)) or (inputs(38));
    layer0_outputs(255) <= '0';
    layer0_outputs(256) <= not((inputs(164)) xor (inputs(114)));
    layer0_outputs(257) <= '1';
    layer0_outputs(258) <= '1';
    layer0_outputs(259) <= not((inputs(15)) or (inputs(132)));
    layer0_outputs(260) <= inputs(1);
    layer0_outputs(261) <= (inputs(254)) and (inputs(253));
    layer0_outputs(262) <= inputs(206);
    layer0_outputs(263) <= inputs(110);
    layer0_outputs(264) <= not(inputs(50)) or (inputs(184));
    layer0_outputs(265) <= '1';
    layer0_outputs(266) <= inputs(27);
    layer0_outputs(267) <= inputs(106);
    layer0_outputs(268) <= inputs(131);
    layer0_outputs(269) <= (inputs(23)) or (inputs(244));
    layer0_outputs(270) <= not(inputs(2)) or (inputs(12));
    layer0_outputs(271) <= (inputs(247)) or (inputs(149));
    layer0_outputs(272) <= '1';
    layer0_outputs(273) <= '0';
    layer0_outputs(274) <= not(inputs(244));
    layer0_outputs(275) <= not(inputs(235));
    layer0_outputs(276) <= '1';
    layer0_outputs(277) <= not(inputs(103)) or (inputs(164));
    layer0_outputs(278) <= (inputs(217)) and (inputs(145));
    layer0_outputs(279) <= not((inputs(183)) or (inputs(99)));
    layer0_outputs(280) <= not((inputs(250)) and (inputs(225)));
    layer0_outputs(281) <= (inputs(45)) and not (inputs(150));
    layer0_outputs(282) <= '0';
    layer0_outputs(283) <= not((inputs(205)) and (inputs(200)));
    layer0_outputs(284) <= '0';
    layer0_outputs(285) <= (inputs(119)) and (inputs(202));
    layer0_outputs(286) <= '0';
    layer0_outputs(287) <= not(inputs(159)) or (inputs(39));
    layer0_outputs(288) <= '1';
    layer0_outputs(289) <= not(inputs(236)) or (inputs(149));
    layer0_outputs(290) <= (inputs(122)) and not (inputs(86));
    layer0_outputs(291) <= not(inputs(194));
    layer0_outputs(292) <= not(inputs(106)) or (inputs(246));
    layer0_outputs(293) <= not(inputs(220)) or (inputs(34));
    layer0_outputs(294) <= inputs(68);
    layer0_outputs(295) <= not((inputs(103)) or (inputs(193)));
    layer0_outputs(296) <= '0';
    layer0_outputs(297) <= not(inputs(27)) or (inputs(157));
    layer0_outputs(298) <= inputs(48);
    layer0_outputs(299) <= not(inputs(170)) or (inputs(151));
    layer0_outputs(300) <= (inputs(204)) and not (inputs(135));
    layer0_outputs(301) <= inputs(0);
    layer0_outputs(302) <= not(inputs(69));
    layer0_outputs(303) <= (inputs(175)) and not (inputs(129));
    layer0_outputs(304) <= not(inputs(100));
    layer0_outputs(305) <= inputs(232);
    layer0_outputs(306) <= not(inputs(136));
    layer0_outputs(307) <= (inputs(79)) and (inputs(254));
    layer0_outputs(308) <= inputs(217);
    layer0_outputs(309) <= not(inputs(86));
    layer0_outputs(310) <= '0';
    layer0_outputs(311) <= not(inputs(193)) or (inputs(249));
    layer0_outputs(312) <= (inputs(84)) and (inputs(40));
    layer0_outputs(313) <= inputs(110);
    layer0_outputs(314) <= '0';
    layer0_outputs(315) <= (inputs(190)) xor (inputs(254));
    layer0_outputs(316) <= (inputs(5)) or (inputs(6));
    layer0_outputs(317) <= (inputs(193)) or (inputs(205));
    layer0_outputs(318) <= (inputs(53)) and not (inputs(191));
    layer0_outputs(319) <= (inputs(39)) and not (inputs(7));
    layer0_outputs(320) <= (inputs(117)) and not (inputs(140));
    layer0_outputs(321) <= inputs(220);
    layer0_outputs(322) <= not(inputs(145)) or (inputs(130));
    layer0_outputs(323) <= '1';
    layer0_outputs(324) <= '0';
    layer0_outputs(325) <= inputs(20);
    layer0_outputs(326) <= not(inputs(18));
    layer0_outputs(327) <= (inputs(14)) or (inputs(17));
    layer0_outputs(328) <= not((inputs(222)) xor (inputs(254)));
    layer0_outputs(329) <= (inputs(219)) and not (inputs(90));
    layer0_outputs(330) <= not((inputs(187)) and (inputs(51)));
    layer0_outputs(331) <= (inputs(70)) and not (inputs(151));
    layer0_outputs(332) <= not(inputs(37));
    layer0_outputs(333) <= '1';
    layer0_outputs(334) <= not((inputs(73)) and (inputs(251)));
    layer0_outputs(335) <= inputs(144);
    layer0_outputs(336) <= not((inputs(119)) or (inputs(97)));
    layer0_outputs(337) <= '1';
    layer0_outputs(338) <= '1';
    layer0_outputs(339) <= not(inputs(53));
    layer0_outputs(340) <= '1';
    layer0_outputs(341) <= inputs(13);
    layer0_outputs(342) <= (inputs(0)) and not (inputs(94));
    layer0_outputs(343) <= inputs(191);
    layer0_outputs(344) <= '1';
    layer0_outputs(345) <= (inputs(163)) and not (inputs(57));
    layer0_outputs(346) <= (inputs(254)) and not (inputs(239));
    layer0_outputs(347) <= not(inputs(122));
    layer0_outputs(348) <= (inputs(126)) xor (inputs(98));
    layer0_outputs(349) <= not(inputs(235)) or (inputs(152));
    layer0_outputs(350) <= not(inputs(208));
    layer0_outputs(351) <= not((inputs(83)) or (inputs(75)));
    layer0_outputs(352) <= (inputs(171)) and (inputs(44));
    layer0_outputs(353) <= not(inputs(9)) or (inputs(198));
    layer0_outputs(354) <= (inputs(192)) or (inputs(251));
    layer0_outputs(355) <= not((inputs(30)) xor (inputs(113)));
    layer0_outputs(356) <= not((inputs(62)) and (inputs(156)));
    layer0_outputs(357) <= '0';
    layer0_outputs(358) <= '1';
    layer0_outputs(359) <= not(inputs(113)) or (inputs(155));
    layer0_outputs(360) <= '0';
    layer0_outputs(361) <= inputs(237);
    layer0_outputs(362) <= not(inputs(32));
    layer0_outputs(363) <= inputs(147);
    layer0_outputs(364) <= inputs(202);
    layer0_outputs(365) <= inputs(118);
    layer0_outputs(366) <= (inputs(80)) or (inputs(179));
    layer0_outputs(367) <= (inputs(172)) and not (inputs(125));
    layer0_outputs(368) <= not((inputs(60)) or (inputs(29)));
    layer0_outputs(369) <= not(inputs(210));
    layer0_outputs(370) <= not(inputs(61));
    layer0_outputs(371) <= (inputs(201)) and not (inputs(144));
    layer0_outputs(372) <= '1';
    layer0_outputs(373) <= not((inputs(93)) or (inputs(175)));
    layer0_outputs(374) <= '1';
    layer0_outputs(375) <= not((inputs(192)) xor (inputs(5)));
    layer0_outputs(376) <= '1';
    layer0_outputs(377) <= (inputs(187)) and not (inputs(238));
    layer0_outputs(378) <= not(inputs(180));
    layer0_outputs(379) <= not((inputs(51)) and (inputs(160)));
    layer0_outputs(380) <= not((inputs(202)) xor (inputs(246)));
    layer0_outputs(381) <= inputs(150);
    layer0_outputs(382) <= (inputs(192)) and (inputs(206));
    layer0_outputs(383) <= (inputs(233)) and not (inputs(34));
    layer0_outputs(384) <= inputs(173);
    layer0_outputs(385) <= inputs(155);
    layer0_outputs(386) <= not((inputs(254)) or (inputs(168)));
    layer0_outputs(387) <= not(inputs(233));
    layer0_outputs(388) <= inputs(198);
    layer0_outputs(389) <= inputs(198);
    layer0_outputs(390) <= (inputs(220)) or (inputs(240));
    layer0_outputs(391) <= (inputs(128)) and not (inputs(203));
    layer0_outputs(392) <= not(inputs(85));
    layer0_outputs(393) <= not(inputs(52)) or (inputs(124));
    layer0_outputs(394) <= not(inputs(37)) or (inputs(96));
    layer0_outputs(395) <= (inputs(247)) and not (inputs(29));
    layer0_outputs(396) <= not((inputs(215)) and (inputs(107)));
    layer0_outputs(397) <= not((inputs(102)) or (inputs(136)));
    layer0_outputs(398) <= (inputs(177)) and not (inputs(84));
    layer0_outputs(399) <= not(inputs(246));
    layer0_outputs(400) <= inputs(180);
    layer0_outputs(401) <= (inputs(163)) and not (inputs(18));
    layer0_outputs(402) <= '1';
    layer0_outputs(403) <= not((inputs(38)) xor (inputs(142)));
    layer0_outputs(404) <= inputs(81);
    layer0_outputs(405) <= not(inputs(159));
    layer0_outputs(406) <= '0';
    layer0_outputs(407) <= not(inputs(188));
    layer0_outputs(408) <= not((inputs(28)) and (inputs(230)));
    layer0_outputs(409) <= not((inputs(230)) or (inputs(83)));
    layer0_outputs(410) <= inputs(120);
    layer0_outputs(411) <= (inputs(95)) and (inputs(128));
    layer0_outputs(412) <= not(inputs(11));
    layer0_outputs(413) <= '1';
    layer0_outputs(414) <= (inputs(84)) or (inputs(76));
    layer0_outputs(415) <= (inputs(55)) and (inputs(161));
    layer0_outputs(416) <= not(inputs(107)) or (inputs(235));
    layer0_outputs(417) <= (inputs(225)) and (inputs(35));
    layer0_outputs(418) <= not(inputs(166)) or (inputs(179));
    layer0_outputs(419) <= inputs(78);
    layer0_outputs(420) <= (inputs(179)) or (inputs(229));
    layer0_outputs(421) <= (inputs(129)) xor (inputs(148));
    layer0_outputs(422) <= not(inputs(187)) or (inputs(236));
    layer0_outputs(423) <= inputs(179);
    layer0_outputs(424) <= not(inputs(149));
    layer0_outputs(425) <= (inputs(104)) and (inputs(201));
    layer0_outputs(426) <= not(inputs(56)) or (inputs(228));
    layer0_outputs(427) <= '1';
    layer0_outputs(428) <= inputs(37);
    layer0_outputs(429) <= not((inputs(77)) or (inputs(157)));
    layer0_outputs(430) <= inputs(120);
    layer0_outputs(431) <= inputs(77);
    layer0_outputs(432) <= '1';
    layer0_outputs(433) <= (inputs(119)) and (inputs(115));
    layer0_outputs(434) <= (inputs(82)) and (inputs(33));
    layer0_outputs(435) <= '0';
    layer0_outputs(436) <= not(inputs(62));
    layer0_outputs(437) <= (inputs(208)) or (inputs(234));
    layer0_outputs(438) <= (inputs(249)) or (inputs(245));
    layer0_outputs(439) <= '0';
    layer0_outputs(440) <= not((inputs(61)) or (inputs(175)));
    layer0_outputs(441) <= (inputs(19)) and (inputs(235));
    layer0_outputs(442) <= not(inputs(212));
    layer0_outputs(443) <= not((inputs(43)) or (inputs(144)));
    layer0_outputs(444) <= '1';
    layer0_outputs(445) <= (inputs(17)) and not (inputs(122));
    layer0_outputs(446) <= (inputs(15)) or (inputs(34));
    layer0_outputs(447) <= '1';
    layer0_outputs(448) <= '0';
    layer0_outputs(449) <= (inputs(88)) or (inputs(243));
    layer0_outputs(450) <= '1';
    layer0_outputs(451) <= not(inputs(23));
    layer0_outputs(452) <= '1';
    layer0_outputs(453) <= inputs(219);
    layer0_outputs(454) <= not(inputs(123)) or (inputs(9));
    layer0_outputs(455) <= not((inputs(45)) or (inputs(134)));
    layer0_outputs(456) <= not(inputs(31));
    layer0_outputs(457) <= (inputs(181)) and not (inputs(73));
    layer0_outputs(458) <= (inputs(82)) or (inputs(29));
    layer0_outputs(459) <= not((inputs(33)) xor (inputs(250)));
    layer0_outputs(460) <= inputs(181);
    layer0_outputs(461) <= not(inputs(253)) or (inputs(74));
    layer0_outputs(462) <= (inputs(203)) and not (inputs(35));
    layer0_outputs(463) <= not(inputs(100));
    layer0_outputs(464) <= inputs(211);
    layer0_outputs(465) <= '0';
    layer0_outputs(466) <= not(inputs(210));
    layer0_outputs(467) <= (inputs(144)) or (inputs(230));
    layer0_outputs(468) <= not(inputs(185)) or (inputs(27));
    layer0_outputs(469) <= (inputs(233)) and (inputs(10));
    layer0_outputs(470) <= (inputs(199)) and (inputs(60));
    layer0_outputs(471) <= not(inputs(193)) or (inputs(164));
    layer0_outputs(472) <= not(inputs(205)) or (inputs(147));
    layer0_outputs(473) <= (inputs(198)) xor (inputs(2));
    layer0_outputs(474) <= (inputs(64)) and not (inputs(35));
    layer0_outputs(475) <= not(inputs(175)) or (inputs(74));
    layer0_outputs(476) <= '1';
    layer0_outputs(477) <= not(inputs(31)) or (inputs(44));
    layer0_outputs(478) <= not((inputs(136)) or (inputs(235)));
    layer0_outputs(479) <= inputs(130);
    layer0_outputs(480) <= not(inputs(88)) or (inputs(179));
    layer0_outputs(481) <= not((inputs(218)) or (inputs(175)));
    layer0_outputs(482) <= '0';
    layer0_outputs(483) <= (inputs(208)) or (inputs(4));
    layer0_outputs(484) <= inputs(166);
    layer0_outputs(485) <= inputs(166);
    layer0_outputs(486) <= not(inputs(229));
    layer0_outputs(487) <= inputs(62);
    layer0_outputs(488) <= (inputs(130)) or (inputs(125));
    layer0_outputs(489) <= (inputs(144)) or (inputs(237));
    layer0_outputs(490) <= inputs(116);
    layer0_outputs(491) <= '1';
    layer0_outputs(492) <= inputs(36);
    layer0_outputs(493) <= not(inputs(222)) or (inputs(157));
    layer0_outputs(494) <= not(inputs(168));
    layer0_outputs(495) <= inputs(255);
    layer0_outputs(496) <= (inputs(72)) xor (inputs(22));
    layer0_outputs(497) <= not((inputs(92)) and (inputs(244)));
    layer0_outputs(498) <= inputs(23);
    layer0_outputs(499) <= inputs(26);
    layer0_outputs(500) <= '0';
    layer0_outputs(501) <= not(inputs(166)) or (inputs(186));
    layer0_outputs(502) <= (inputs(67)) and (inputs(179));
    layer0_outputs(503) <= not(inputs(23)) or (inputs(129));
    layer0_outputs(504) <= not(inputs(42)) or (inputs(234));
    layer0_outputs(505) <= '0';
    layer0_outputs(506) <= not((inputs(70)) or (inputs(86)));
    layer0_outputs(507) <= not(inputs(215));
    layer0_outputs(508) <= inputs(84);
    layer0_outputs(509) <= (inputs(46)) or (inputs(56));
    layer0_outputs(510) <= inputs(67);
    layer0_outputs(511) <= not(inputs(156)) or (inputs(28));
    layer0_outputs(512) <= not(inputs(104));
    layer0_outputs(513) <= (inputs(215)) and not (inputs(169));
    layer0_outputs(514) <= not(inputs(210));
    layer0_outputs(515) <= (inputs(77)) and (inputs(228));
    layer0_outputs(516) <= (inputs(167)) and not (inputs(130));
    layer0_outputs(517) <= not(inputs(53)) or (inputs(34));
    layer0_outputs(518) <= inputs(166);
    layer0_outputs(519) <= not(inputs(227)) or (inputs(89));
    layer0_outputs(520) <= '1';
    layer0_outputs(521) <= inputs(24);
    layer0_outputs(522) <= inputs(149);
    layer0_outputs(523) <= inputs(106);
    layer0_outputs(524) <= '1';
    layer0_outputs(525) <= inputs(24);
    layer0_outputs(526) <= '1';
    layer0_outputs(527) <= not((inputs(251)) and (inputs(82)));
    layer0_outputs(528) <= not((inputs(50)) xor (inputs(10)));
    layer0_outputs(529) <= (inputs(241)) and (inputs(193));
    layer0_outputs(530) <= inputs(118);
    layer0_outputs(531) <= '0';
    layer0_outputs(532) <= not(inputs(94));
    layer0_outputs(533) <= (inputs(138)) and not (inputs(214));
    layer0_outputs(534) <= not(inputs(230));
    layer0_outputs(535) <= not(inputs(127)) or (inputs(12));
    layer0_outputs(536) <= not((inputs(88)) and (inputs(153)));
    layer0_outputs(537) <= inputs(148);
    layer0_outputs(538) <= (inputs(25)) and not (inputs(204));
    layer0_outputs(539) <= not((inputs(104)) or (inputs(103)));
    layer0_outputs(540) <= not(inputs(192));
    layer0_outputs(541) <= not(inputs(151)) or (inputs(44));
    layer0_outputs(542) <= not(inputs(36));
    layer0_outputs(543) <= not((inputs(53)) or (inputs(232)));
    layer0_outputs(544) <= '1';
    layer0_outputs(545) <= not(inputs(16));
    layer0_outputs(546) <= (inputs(123)) and not (inputs(115));
    layer0_outputs(547) <= (inputs(127)) and not (inputs(3));
    layer0_outputs(548) <= inputs(64);
    layer0_outputs(549) <= (inputs(25)) and not (inputs(18));
    layer0_outputs(550) <= '1';
    layer0_outputs(551) <= not((inputs(204)) or (inputs(236)));
    layer0_outputs(552) <= not((inputs(87)) or (inputs(140)));
    layer0_outputs(553) <= (inputs(107)) and not (inputs(36));
    layer0_outputs(554) <= (inputs(32)) or (inputs(171));
    layer0_outputs(555) <= '0';
    layer0_outputs(556) <= not((inputs(146)) or (inputs(188)));
    layer0_outputs(557) <= (inputs(0)) or (inputs(60));
    layer0_outputs(558) <= '0';
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= not((inputs(121)) and (inputs(4)));
    layer0_outputs(561) <= not(inputs(34));
    layer0_outputs(562) <= inputs(209);
    layer0_outputs(563) <= not(inputs(111));
    layer0_outputs(564) <= not(inputs(222)) or (inputs(65));
    layer0_outputs(565) <= inputs(120);
    layer0_outputs(566) <= inputs(239);
    layer0_outputs(567) <= not(inputs(99));
    layer0_outputs(568) <= (inputs(48)) and not (inputs(120));
    layer0_outputs(569) <= not(inputs(238));
    layer0_outputs(570) <= (inputs(76)) and not (inputs(22));
    layer0_outputs(571) <= (inputs(124)) and not (inputs(222));
    layer0_outputs(572) <= (inputs(141)) and not (inputs(150));
    layer0_outputs(573) <= '0';
    layer0_outputs(574) <= '0';
    layer0_outputs(575) <= '1';
    layer0_outputs(576) <= not(inputs(119));
    layer0_outputs(577) <= (inputs(55)) xor (inputs(40));
    layer0_outputs(578) <= inputs(150);
    layer0_outputs(579) <= (inputs(1)) or (inputs(208));
    layer0_outputs(580) <= inputs(37);
    layer0_outputs(581) <= not((inputs(243)) or (inputs(13)));
    layer0_outputs(582) <= (inputs(255)) and (inputs(191));
    layer0_outputs(583) <= '1';
    layer0_outputs(584) <= '1';
    layer0_outputs(585) <= inputs(210);
    layer0_outputs(586) <= (inputs(156)) or (inputs(162));
    layer0_outputs(587) <= not(inputs(191)) or (inputs(174));
    layer0_outputs(588) <= inputs(165);
    layer0_outputs(589) <= (inputs(5)) or (inputs(90));
    layer0_outputs(590) <= inputs(105);
    layer0_outputs(591) <= not((inputs(38)) or (inputs(149)));
    layer0_outputs(592) <= inputs(51);
    layer0_outputs(593) <= (inputs(114)) and not (inputs(96));
    layer0_outputs(594) <= not((inputs(235)) and (inputs(54)));
    layer0_outputs(595) <= (inputs(174)) or (inputs(171));
    layer0_outputs(596) <= (inputs(153)) and not (inputs(87));
    layer0_outputs(597) <= not(inputs(16));
    layer0_outputs(598) <= not((inputs(141)) xor (inputs(143)));
    layer0_outputs(599) <= not((inputs(220)) and (inputs(42)));
    layer0_outputs(600) <= (inputs(81)) and not (inputs(107));
    layer0_outputs(601) <= not((inputs(176)) and (inputs(202)));
    layer0_outputs(602) <= (inputs(74)) and not (inputs(17));
    layer0_outputs(603) <= inputs(36);
    layer0_outputs(604) <= inputs(182);
    layer0_outputs(605) <= not((inputs(40)) or (inputs(128)));
    layer0_outputs(606) <= (inputs(233)) and not (inputs(157));
    layer0_outputs(607) <= (inputs(147)) or (inputs(158));
    layer0_outputs(608) <= '0';
    layer0_outputs(609) <= '1';
    layer0_outputs(610) <= (inputs(206)) and (inputs(248));
    layer0_outputs(611) <= inputs(52);
    layer0_outputs(612) <= (inputs(40)) and (inputs(82));
    layer0_outputs(613) <= inputs(109);
    layer0_outputs(614) <= inputs(74);
    layer0_outputs(615) <= not((inputs(94)) and (inputs(11)));
    layer0_outputs(616) <= inputs(2);
    layer0_outputs(617) <= not(inputs(106));
    layer0_outputs(618) <= (inputs(45)) and (inputs(58));
    layer0_outputs(619) <= not((inputs(35)) or (inputs(194)));
    layer0_outputs(620) <= not(inputs(111)) or (inputs(21));
    layer0_outputs(621) <= inputs(106);
    layer0_outputs(622) <= (inputs(65)) or (inputs(99));
    layer0_outputs(623) <= (inputs(29)) and not (inputs(251));
    layer0_outputs(624) <= not((inputs(53)) or (inputs(171)));
    layer0_outputs(625) <= '1';
    layer0_outputs(626) <= inputs(168);
    layer0_outputs(627) <= inputs(120);
    layer0_outputs(628) <= inputs(223);
    layer0_outputs(629) <= '1';
    layer0_outputs(630) <= not((inputs(161)) or (inputs(147)));
    layer0_outputs(631) <= (inputs(42)) and (inputs(6));
    layer0_outputs(632) <= not((inputs(188)) or (inputs(97)));
    layer0_outputs(633) <= not(inputs(193)) or (inputs(202));
    layer0_outputs(634) <= not(inputs(162)) or (inputs(123));
    layer0_outputs(635) <= (inputs(17)) or (inputs(39));
    layer0_outputs(636) <= (inputs(183)) and (inputs(178));
    layer0_outputs(637) <= not(inputs(162));
    layer0_outputs(638) <= '1';
    layer0_outputs(639) <= inputs(151);
    layer0_outputs(640) <= not(inputs(176));
    layer0_outputs(641) <= not(inputs(85));
    layer0_outputs(642) <= not(inputs(103));
    layer0_outputs(643) <= not(inputs(109)) or (inputs(62));
    layer0_outputs(644) <= '0';
    layer0_outputs(645) <= (inputs(243)) and (inputs(5));
    layer0_outputs(646) <= (inputs(159)) and (inputs(166));
    layer0_outputs(647) <= not(inputs(135));
    layer0_outputs(648) <= (inputs(53)) and (inputs(9));
    layer0_outputs(649) <= '0';
    layer0_outputs(650) <= not((inputs(86)) or (inputs(192)));
    layer0_outputs(651) <= not(inputs(155));
    layer0_outputs(652) <= not(inputs(186));
    layer0_outputs(653) <= not(inputs(126));
    layer0_outputs(654) <= inputs(129);
    layer0_outputs(655) <= '1';
    layer0_outputs(656) <= inputs(99);
    layer0_outputs(657) <= '1';
    layer0_outputs(658) <= not((inputs(149)) xor (inputs(252)));
    layer0_outputs(659) <= inputs(214);
    layer0_outputs(660) <= inputs(239);
    layer0_outputs(661) <= inputs(112);
    layer0_outputs(662) <= not(inputs(68));
    layer0_outputs(663) <= (inputs(84)) xor (inputs(252));
    layer0_outputs(664) <= not((inputs(41)) or (inputs(133)));
    layer0_outputs(665) <= '1';
    layer0_outputs(666) <= (inputs(124)) or (inputs(254));
    layer0_outputs(667) <= not(inputs(79)) or (inputs(51));
    layer0_outputs(668) <= (inputs(176)) or (inputs(149));
    layer0_outputs(669) <= not(inputs(61));
    layer0_outputs(670) <= (inputs(133)) and not (inputs(242));
    layer0_outputs(671) <= not((inputs(218)) or (inputs(6)));
    layer0_outputs(672) <= (inputs(68)) and not (inputs(202));
    layer0_outputs(673) <= not(inputs(165));
    layer0_outputs(674) <= not(inputs(88));
    layer0_outputs(675) <= (inputs(169)) or (inputs(86));
    layer0_outputs(676) <= (inputs(195)) or (inputs(254));
    layer0_outputs(677) <= not(inputs(69)) or (inputs(56));
    layer0_outputs(678) <= not((inputs(42)) or (inputs(62)));
    layer0_outputs(679) <= (inputs(144)) and (inputs(245));
    layer0_outputs(680) <= (inputs(180)) or (inputs(210));
    layer0_outputs(681) <= not(inputs(137)) or (inputs(80));
    layer0_outputs(682) <= not(inputs(161)) or (inputs(231));
    layer0_outputs(683) <= not(inputs(160));
    layer0_outputs(684) <= not(inputs(22)) or (inputs(190));
    layer0_outputs(685) <= (inputs(116)) or (inputs(155));
    layer0_outputs(686) <= not((inputs(164)) and (inputs(67)));
    layer0_outputs(687) <= (inputs(136)) and not (inputs(46));
    layer0_outputs(688) <= not((inputs(10)) and (inputs(122)));
    layer0_outputs(689) <= '0';
    layer0_outputs(690) <= (inputs(1)) and not (inputs(155));
    layer0_outputs(691) <= not((inputs(158)) xor (inputs(109)));
    layer0_outputs(692) <= inputs(192);
    layer0_outputs(693) <= (inputs(57)) and not (inputs(171));
    layer0_outputs(694) <= (inputs(207)) or (inputs(46));
    layer0_outputs(695) <= (inputs(214)) and (inputs(21));
    layer0_outputs(696) <= (inputs(252)) and (inputs(244));
    layer0_outputs(697) <= (inputs(34)) or (inputs(19));
    layer0_outputs(698) <= (inputs(47)) and not (inputs(212));
    layer0_outputs(699) <= (inputs(95)) and not (inputs(254));
    layer0_outputs(700) <= '0';
    layer0_outputs(701) <= (inputs(70)) and (inputs(183));
    layer0_outputs(702) <= (inputs(59)) and not (inputs(186));
    layer0_outputs(703) <= not(inputs(109)) or (inputs(153));
    layer0_outputs(704) <= '1';
    layer0_outputs(705) <= not((inputs(247)) and (inputs(210)));
    layer0_outputs(706) <= not(inputs(193));
    layer0_outputs(707) <= not(inputs(150)) or (inputs(241));
    layer0_outputs(708) <= not((inputs(134)) and (inputs(177)));
    layer0_outputs(709) <= not(inputs(127)) or (inputs(241));
    layer0_outputs(710) <= '0';
    layer0_outputs(711) <= '1';
    layer0_outputs(712) <= '0';
    layer0_outputs(713) <= not((inputs(129)) or (inputs(126)));
    layer0_outputs(714) <= (inputs(98)) or (inputs(83));
    layer0_outputs(715) <= not((inputs(11)) or (inputs(108)));
    layer0_outputs(716) <= (inputs(117)) or (inputs(77));
    layer0_outputs(717) <= '0';
    layer0_outputs(718) <= not((inputs(232)) and (inputs(113)));
    layer0_outputs(719) <= inputs(60);
    layer0_outputs(720) <= not(inputs(119)) or (inputs(82));
    layer0_outputs(721) <= not(inputs(100)) or (inputs(201));
    layer0_outputs(722) <= not(inputs(183));
    layer0_outputs(723) <= inputs(4);
    layer0_outputs(724) <= not(inputs(117));
    layer0_outputs(725) <= not(inputs(96)) or (inputs(199));
    layer0_outputs(726) <= '0';
    layer0_outputs(727) <= (inputs(131)) and not (inputs(250));
    layer0_outputs(728) <= not(inputs(188)) or (inputs(189));
    layer0_outputs(729) <= (inputs(28)) and (inputs(146));
    layer0_outputs(730) <= inputs(56);
    layer0_outputs(731) <= not(inputs(196)) or (inputs(128));
    layer0_outputs(732) <= '1';
    layer0_outputs(733) <= (inputs(83)) or (inputs(177));
    layer0_outputs(734) <= (inputs(31)) and (inputs(91));
    layer0_outputs(735) <= not(inputs(59));
    layer0_outputs(736) <= (inputs(136)) or (inputs(153));
    layer0_outputs(737) <= (inputs(45)) and (inputs(129));
    layer0_outputs(738) <= inputs(248);
    layer0_outputs(739) <= not(inputs(195));
    layer0_outputs(740) <= inputs(216);
    layer0_outputs(741) <= '1';
    layer0_outputs(742) <= not((inputs(171)) or (inputs(26)));
    layer0_outputs(743) <= inputs(175);
    layer0_outputs(744) <= '0';
    layer0_outputs(745) <= not((inputs(51)) or (inputs(212)));
    layer0_outputs(746) <= not((inputs(52)) and (inputs(209)));
    layer0_outputs(747) <= '1';
    layer0_outputs(748) <= not((inputs(137)) or (inputs(153)));
    layer0_outputs(749) <= inputs(177);
    layer0_outputs(750) <= inputs(122);
    layer0_outputs(751) <= not((inputs(22)) or (inputs(18)));
    layer0_outputs(752) <= (inputs(125)) and (inputs(228));
    layer0_outputs(753) <= (inputs(210)) and (inputs(72));
    layer0_outputs(754) <= not((inputs(40)) and (inputs(85)));
    layer0_outputs(755) <= '1';
    layer0_outputs(756) <= not((inputs(101)) and (inputs(61)));
    layer0_outputs(757) <= not(inputs(201));
    layer0_outputs(758) <= (inputs(2)) and not (inputs(104));
    layer0_outputs(759) <= '1';
    layer0_outputs(760) <= (inputs(2)) or (inputs(95));
    layer0_outputs(761) <= inputs(103);
    layer0_outputs(762) <= (inputs(172)) or (inputs(224));
    layer0_outputs(763) <= not((inputs(93)) xor (inputs(90)));
    layer0_outputs(764) <= not(inputs(85)) or (inputs(63));
    layer0_outputs(765) <= inputs(103);
    layer0_outputs(766) <= (inputs(96)) and not (inputs(175));
    layer0_outputs(767) <= (inputs(100)) and (inputs(158));
    layer0_outputs(768) <= not(inputs(222));
    layer0_outputs(769) <= not(inputs(109)) or (inputs(178));
    layer0_outputs(770) <= not(inputs(164));
    layer0_outputs(771) <= not(inputs(102));
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= inputs(136);
    layer0_outputs(774) <= not(inputs(169));
    layer0_outputs(775) <= not(inputs(88)) or (inputs(45));
    layer0_outputs(776) <= (inputs(91)) and (inputs(98));
    layer0_outputs(777) <= (inputs(210)) or (inputs(117));
    layer0_outputs(778) <= not((inputs(138)) and (inputs(26)));
    layer0_outputs(779) <= not(inputs(112));
    layer0_outputs(780) <= inputs(246);
    layer0_outputs(781) <= inputs(178);
    layer0_outputs(782) <= not(inputs(149)) or (inputs(111));
    layer0_outputs(783) <= (inputs(193)) or (inputs(220));
    layer0_outputs(784) <= (inputs(91)) and (inputs(74));
    layer0_outputs(785) <= inputs(111);
    layer0_outputs(786) <= not(inputs(69));
    layer0_outputs(787) <= (inputs(26)) and not (inputs(255));
    layer0_outputs(788) <= (inputs(117)) or (inputs(101));
    layer0_outputs(789) <= (inputs(44)) and (inputs(41));
    layer0_outputs(790) <= (inputs(31)) and not (inputs(184));
    layer0_outputs(791) <= inputs(210);
    layer0_outputs(792) <= not(inputs(203));
    layer0_outputs(793) <= not(inputs(99)) or (inputs(191));
    layer0_outputs(794) <= '0';
    layer0_outputs(795) <= (inputs(133)) or (inputs(37));
    layer0_outputs(796) <= (inputs(136)) and (inputs(128));
    layer0_outputs(797) <= not(inputs(10));
    layer0_outputs(798) <= not(inputs(135));
    layer0_outputs(799) <= (inputs(240)) and (inputs(147));
    layer0_outputs(800) <= not((inputs(164)) and (inputs(151)));
    layer0_outputs(801) <= not((inputs(113)) or (inputs(10)));
    layer0_outputs(802) <= '0';
    layer0_outputs(803) <= inputs(103);
    layer0_outputs(804) <= (inputs(142)) and not (inputs(187));
    layer0_outputs(805) <= not((inputs(158)) or (inputs(173)));
    layer0_outputs(806) <= '1';
    layer0_outputs(807) <= not(inputs(41)) or (inputs(205));
    layer0_outputs(808) <= '0';
    layer0_outputs(809) <= (inputs(177)) and (inputs(125));
    layer0_outputs(810) <= '1';
    layer0_outputs(811) <= (inputs(135)) and not (inputs(222));
    layer0_outputs(812) <= not((inputs(59)) or (inputs(30)));
    layer0_outputs(813) <= (inputs(223)) and not (inputs(71));
    layer0_outputs(814) <= inputs(8);
    layer0_outputs(815) <= not((inputs(236)) or (inputs(124)));
    layer0_outputs(816) <= not((inputs(56)) or (inputs(20)));
    layer0_outputs(817) <= not(inputs(195));
    layer0_outputs(818) <= '0';
    layer0_outputs(819) <= (inputs(104)) and not (inputs(25));
    layer0_outputs(820) <= not(inputs(104)) or (inputs(190));
    layer0_outputs(821) <= '0';
    layer0_outputs(822) <= not(inputs(164)) or (inputs(49));
    layer0_outputs(823) <= not(inputs(52)) or (inputs(22));
    layer0_outputs(824) <= (inputs(56)) and not (inputs(200));
    layer0_outputs(825) <= inputs(211);
    layer0_outputs(826) <= inputs(199);
    layer0_outputs(827) <= not((inputs(96)) xor (inputs(131)));
    layer0_outputs(828) <= (inputs(25)) or (inputs(46));
    layer0_outputs(829) <= (inputs(107)) and not (inputs(13));
    layer0_outputs(830) <= (inputs(140)) and not (inputs(66));
    layer0_outputs(831) <= (inputs(189)) and not (inputs(21));
    layer0_outputs(832) <= (inputs(133)) or (inputs(81));
    layer0_outputs(833) <= not((inputs(62)) or (inputs(158)));
    layer0_outputs(834) <= '0';
    layer0_outputs(835) <= not((inputs(0)) and (inputs(190)));
    layer0_outputs(836) <= not((inputs(80)) or (inputs(66)));
    layer0_outputs(837) <= not(inputs(231)) or (inputs(59));
    layer0_outputs(838) <= (inputs(203)) and (inputs(57));
    layer0_outputs(839) <= '1';
    layer0_outputs(840) <= (inputs(89)) and not (inputs(88));
    layer0_outputs(841) <= '0';
    layer0_outputs(842) <= not((inputs(142)) and (inputs(227)));
    layer0_outputs(843) <= not((inputs(111)) or (inputs(4)));
    layer0_outputs(844) <= inputs(56);
    layer0_outputs(845) <= not(inputs(137));
    layer0_outputs(846) <= not((inputs(193)) and (inputs(197)));
    layer0_outputs(847) <= (inputs(66)) and not (inputs(174));
    layer0_outputs(848) <= not(inputs(101));
    layer0_outputs(849) <= (inputs(225)) and not (inputs(49));
    layer0_outputs(850) <= not(inputs(126));
    layer0_outputs(851) <= '0';
    layer0_outputs(852) <= (inputs(151)) and not (inputs(83));
    layer0_outputs(853) <= inputs(51);
    layer0_outputs(854) <= (inputs(117)) or (inputs(196));
    layer0_outputs(855) <= not(inputs(105));
    layer0_outputs(856) <= '1';
    layer0_outputs(857) <= (inputs(15)) and not (inputs(182));
    layer0_outputs(858) <= inputs(56);
    layer0_outputs(859) <= (inputs(12)) and not (inputs(20));
    layer0_outputs(860) <= '1';
    layer0_outputs(861) <= (inputs(139)) and (inputs(126));
    layer0_outputs(862) <= not(inputs(44)) or (inputs(239));
    layer0_outputs(863) <= not(inputs(37)) or (inputs(190));
    layer0_outputs(864) <= not(inputs(113));
    layer0_outputs(865) <= '1';
    layer0_outputs(866) <= (inputs(209)) and not (inputs(148));
    layer0_outputs(867) <= (inputs(76)) and (inputs(103));
    layer0_outputs(868) <= '1';
    layer0_outputs(869) <= (inputs(201)) or (inputs(182));
    layer0_outputs(870) <= (inputs(134)) or (inputs(153));
    layer0_outputs(871) <= inputs(174);
    layer0_outputs(872) <= not(inputs(151)) or (inputs(48));
    layer0_outputs(873) <= not(inputs(69));
    layer0_outputs(874) <= (inputs(63)) and (inputs(108));
    layer0_outputs(875) <= '1';
    layer0_outputs(876) <= not(inputs(196));
    layer0_outputs(877) <= '0';
    layer0_outputs(878) <= not(inputs(102));
    layer0_outputs(879) <= '0';
    layer0_outputs(880) <= (inputs(220)) or (inputs(234));
    layer0_outputs(881) <= inputs(106);
    layer0_outputs(882) <= (inputs(180)) and (inputs(197));
    layer0_outputs(883) <= not(inputs(135));
    layer0_outputs(884) <= '0';
    layer0_outputs(885) <= not(inputs(201));
    layer0_outputs(886) <= not((inputs(164)) xor (inputs(160)));
    layer0_outputs(887) <= not(inputs(24));
    layer0_outputs(888) <= not(inputs(105));
    layer0_outputs(889) <= '1';
    layer0_outputs(890) <= not(inputs(4)) or (inputs(112));
    layer0_outputs(891) <= (inputs(14)) and not (inputs(54));
    layer0_outputs(892) <= not((inputs(27)) and (inputs(66)));
    layer0_outputs(893) <= '1';
    layer0_outputs(894) <= '1';
    layer0_outputs(895) <= not(inputs(254));
    layer0_outputs(896) <= not((inputs(144)) xor (inputs(163)));
    layer0_outputs(897) <= '1';
    layer0_outputs(898) <= not((inputs(123)) or (inputs(12)));
    layer0_outputs(899) <= '1';
    layer0_outputs(900) <= not((inputs(46)) and (inputs(212)));
    layer0_outputs(901) <= not(inputs(164));
    layer0_outputs(902) <= not(inputs(51));
    layer0_outputs(903) <= not((inputs(66)) or (inputs(109)));
    layer0_outputs(904) <= not((inputs(246)) or (inputs(225)));
    layer0_outputs(905) <= (inputs(79)) and not (inputs(10));
    layer0_outputs(906) <= not((inputs(98)) or (inputs(224)));
    layer0_outputs(907) <= inputs(228);
    layer0_outputs(908) <= not((inputs(215)) or (inputs(231)));
    layer0_outputs(909) <= (inputs(62)) and not (inputs(200));
    layer0_outputs(910) <= (inputs(207)) xor (inputs(67));
    layer0_outputs(911) <= not(inputs(158));
    layer0_outputs(912) <= inputs(196);
    layer0_outputs(913) <= not(inputs(103)) or (inputs(187));
    layer0_outputs(914) <= not((inputs(93)) or (inputs(24)));
    layer0_outputs(915) <= '0';
    layer0_outputs(916) <= '0';
    layer0_outputs(917) <= inputs(131);
    layer0_outputs(918) <= '1';
    layer0_outputs(919) <= (inputs(245)) xor (inputs(209));
    layer0_outputs(920) <= inputs(239);
    layer0_outputs(921) <= inputs(213);
    layer0_outputs(922) <= '1';
    layer0_outputs(923) <= not(inputs(76)) or (inputs(209));
    layer0_outputs(924) <= (inputs(57)) and not (inputs(0));
    layer0_outputs(925) <= (inputs(52)) or (inputs(20));
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= '0';
    layer0_outputs(928) <= not(inputs(211));
    layer0_outputs(929) <= not(inputs(171));
    layer0_outputs(930) <= not((inputs(130)) xor (inputs(47)));
    layer0_outputs(931) <= '0';
    layer0_outputs(932) <= not((inputs(124)) or (inputs(75)));
    layer0_outputs(933) <= inputs(147);
    layer0_outputs(934) <= not(inputs(33));
    layer0_outputs(935) <= (inputs(199)) and (inputs(156));
    layer0_outputs(936) <= not((inputs(111)) xor (inputs(223)));
    layer0_outputs(937) <= '0';
    layer0_outputs(938) <= not(inputs(158));
    layer0_outputs(939) <= not((inputs(111)) or (inputs(55)));
    layer0_outputs(940) <= inputs(151);
    layer0_outputs(941) <= '1';
    layer0_outputs(942) <= (inputs(175)) and (inputs(226));
    layer0_outputs(943) <= not(inputs(139)) or (inputs(140));
    layer0_outputs(944) <= inputs(102);
    layer0_outputs(945) <= inputs(166);
    layer0_outputs(946) <= not(inputs(187)) or (inputs(122));
    layer0_outputs(947) <= not(inputs(120)) or (inputs(84));
    layer0_outputs(948) <= (inputs(11)) and not (inputs(204));
    layer0_outputs(949) <= inputs(229);
    layer0_outputs(950) <= '1';
    layer0_outputs(951) <= not(inputs(82));
    layer0_outputs(952) <= (inputs(20)) and not (inputs(106));
    layer0_outputs(953) <= inputs(25);
    layer0_outputs(954) <= '0';
    layer0_outputs(955) <= (inputs(121)) and not (inputs(165));
    layer0_outputs(956) <= inputs(153);
    layer0_outputs(957) <= not((inputs(178)) or (inputs(83)));
    layer0_outputs(958) <= (inputs(2)) and not (inputs(76));
    layer0_outputs(959) <= not(inputs(73)) or (inputs(135));
    layer0_outputs(960) <= (inputs(234)) and (inputs(209));
    layer0_outputs(961) <= not(inputs(163));
    layer0_outputs(962) <= '0';
    layer0_outputs(963) <= (inputs(68)) and not (inputs(201));
    layer0_outputs(964) <= not((inputs(29)) and (inputs(6)));
    layer0_outputs(965) <= not((inputs(252)) and (inputs(84)));
    layer0_outputs(966) <= '1';
    layer0_outputs(967) <= (inputs(210)) or (inputs(178));
    layer0_outputs(968) <= (inputs(192)) and not (inputs(199));
    layer0_outputs(969) <= not(inputs(70)) or (inputs(108));
    layer0_outputs(970) <= '1';
    layer0_outputs(971) <= not(inputs(209)) or (inputs(125));
    layer0_outputs(972) <= (inputs(6)) and (inputs(20));
    layer0_outputs(973) <= not((inputs(148)) or (inputs(236)));
    layer0_outputs(974) <= (inputs(43)) or (inputs(192));
    layer0_outputs(975) <= (inputs(234)) and not (inputs(84));
    layer0_outputs(976) <= inputs(231);
    layer0_outputs(977) <= (inputs(32)) and not (inputs(11));
    layer0_outputs(978) <= '1';
    layer0_outputs(979) <= not((inputs(100)) and (inputs(108)));
    layer0_outputs(980) <= not(inputs(204));
    layer0_outputs(981) <= not(inputs(14));
    layer0_outputs(982) <= inputs(132);
    layer0_outputs(983) <= (inputs(84)) and not (inputs(58));
    layer0_outputs(984) <= (inputs(16)) and not (inputs(199));
    layer0_outputs(985) <= '0';
    layer0_outputs(986) <= not(inputs(98));
    layer0_outputs(987) <= (inputs(140)) or (inputs(172));
    layer0_outputs(988) <= '1';
    layer0_outputs(989) <= not((inputs(29)) or (inputs(167)));
    layer0_outputs(990) <= (inputs(16)) or (inputs(128));
    layer0_outputs(991) <= not((inputs(173)) xor (inputs(177)));
    layer0_outputs(992) <= inputs(44);
    layer0_outputs(993) <= not(inputs(228)) or (inputs(221));
    layer0_outputs(994) <= inputs(42);
    layer0_outputs(995) <= inputs(85);
    layer0_outputs(996) <= '1';
    layer0_outputs(997) <= (inputs(172)) or (inputs(122));
    layer0_outputs(998) <= (inputs(215)) and (inputs(127));
    layer0_outputs(999) <= '0';
    layer0_outputs(1000) <= inputs(178);
    layer0_outputs(1001) <= inputs(232);
    layer0_outputs(1002) <= '1';
    layer0_outputs(1003) <= '1';
    layer0_outputs(1004) <= '1';
    layer0_outputs(1005) <= (inputs(60)) or (inputs(30));
    layer0_outputs(1006) <= (inputs(30)) or (inputs(72));
    layer0_outputs(1007) <= '0';
    layer0_outputs(1008) <= (inputs(136)) and not (inputs(225));
    layer0_outputs(1009) <= (inputs(77)) and (inputs(54));
    layer0_outputs(1010) <= inputs(220);
    layer0_outputs(1011) <= (inputs(35)) or (inputs(0));
    layer0_outputs(1012) <= '1';
    layer0_outputs(1013) <= inputs(40);
    layer0_outputs(1014) <= (inputs(14)) and not (inputs(18));
    layer0_outputs(1015) <= not(inputs(59));
    layer0_outputs(1016) <= not(inputs(196));
    layer0_outputs(1017) <= not(inputs(0));
    layer0_outputs(1018) <= (inputs(242)) and not (inputs(112));
    layer0_outputs(1019) <= inputs(128);
    layer0_outputs(1020) <= (inputs(69)) or (inputs(114));
    layer0_outputs(1021) <= not(inputs(7)) or (inputs(14));
    layer0_outputs(1022) <= (inputs(127)) or (inputs(233));
    layer0_outputs(1023) <= inputs(97);
    layer0_outputs(1024) <= not((inputs(103)) and (inputs(226)));
    layer0_outputs(1025) <= (inputs(204)) or (inputs(76));
    layer0_outputs(1026) <= (inputs(236)) and not (inputs(165));
    layer0_outputs(1027) <= not(inputs(200));
    layer0_outputs(1028) <= not((inputs(239)) or (inputs(34)));
    layer0_outputs(1029) <= '0';
    layer0_outputs(1030) <= (inputs(20)) and not (inputs(212));
    layer0_outputs(1031) <= not((inputs(96)) xor (inputs(21)));
    layer0_outputs(1032) <= inputs(238);
    layer0_outputs(1033) <= (inputs(24)) or (inputs(171));
    layer0_outputs(1034) <= '0';
    layer0_outputs(1035) <= (inputs(227)) and not (inputs(246));
    layer0_outputs(1036) <= '1';
    layer0_outputs(1037) <= inputs(195);
    layer0_outputs(1038) <= (inputs(192)) xor (inputs(47));
    layer0_outputs(1039) <= (inputs(218)) and not (inputs(66));
    layer0_outputs(1040) <= (inputs(237)) and not (inputs(193));
    layer0_outputs(1041) <= '0';
    layer0_outputs(1042) <= not((inputs(22)) or (inputs(207)));
    layer0_outputs(1043) <= (inputs(223)) xor (inputs(229));
    layer0_outputs(1044) <= '1';
    layer0_outputs(1045) <= (inputs(101)) and not (inputs(124));
    layer0_outputs(1046) <= not((inputs(41)) or (inputs(151)));
    layer0_outputs(1047) <= not(inputs(233));
    layer0_outputs(1048) <= '0';
    layer0_outputs(1049) <= not(inputs(46)) or (inputs(182));
    layer0_outputs(1050) <= not(inputs(25));
    layer0_outputs(1051) <= not((inputs(102)) and (inputs(32)));
    layer0_outputs(1052) <= inputs(238);
    layer0_outputs(1053) <= (inputs(192)) and (inputs(192));
    layer0_outputs(1054) <= inputs(106);
    layer0_outputs(1055) <= (inputs(123)) and not (inputs(215));
    layer0_outputs(1056) <= '1';
    layer0_outputs(1057) <= '0';
    layer0_outputs(1058) <= inputs(14);
    layer0_outputs(1059) <= not(inputs(113));
    layer0_outputs(1060) <= not(inputs(187)) or (inputs(250));
    layer0_outputs(1061) <= inputs(137);
    layer0_outputs(1062) <= (inputs(70)) and not (inputs(0));
    layer0_outputs(1063) <= not(inputs(188));
    layer0_outputs(1064) <= inputs(188);
    layer0_outputs(1065) <= (inputs(36)) and not (inputs(231));
    layer0_outputs(1066) <= not(inputs(179));
    layer0_outputs(1067) <= inputs(180);
    layer0_outputs(1068) <= inputs(175);
    layer0_outputs(1069) <= (inputs(64)) and not (inputs(125));
    layer0_outputs(1070) <= not((inputs(230)) or (inputs(243)));
    layer0_outputs(1071) <= (inputs(179)) or (inputs(238));
    layer0_outputs(1072) <= '1';
    layer0_outputs(1073) <= '1';
    layer0_outputs(1074) <= inputs(149);
    layer0_outputs(1075) <= inputs(93);
    layer0_outputs(1076) <= inputs(123);
    layer0_outputs(1077) <= not(inputs(124)) or (inputs(183));
    layer0_outputs(1078) <= inputs(118);
    layer0_outputs(1079) <= inputs(13);
    layer0_outputs(1080) <= not(inputs(137)) or (inputs(220));
    layer0_outputs(1081) <= (inputs(76)) or (inputs(243));
    layer0_outputs(1082) <= not(inputs(228));
    layer0_outputs(1083) <= not(inputs(24));
    layer0_outputs(1084) <= not(inputs(237));
    layer0_outputs(1085) <= inputs(99);
    layer0_outputs(1086) <= inputs(231);
    layer0_outputs(1087) <= inputs(36);
    layer0_outputs(1088) <= not((inputs(144)) or (inputs(213)));
    layer0_outputs(1089) <= not((inputs(202)) xor (inputs(219)));
    layer0_outputs(1090) <= (inputs(78)) and not (inputs(17));
    layer0_outputs(1091) <= not(inputs(181));
    layer0_outputs(1092) <= (inputs(16)) xor (inputs(106));
    layer0_outputs(1093) <= not(inputs(135));
    layer0_outputs(1094) <= (inputs(42)) and (inputs(41));
    layer0_outputs(1095) <= '1';
    layer0_outputs(1096) <= (inputs(243)) or (inputs(213));
    layer0_outputs(1097) <= '1';
    layer0_outputs(1098) <= not(inputs(106));
    layer0_outputs(1099) <= (inputs(108)) or (inputs(207));
    layer0_outputs(1100) <= '1';
    layer0_outputs(1101) <= not((inputs(220)) or (inputs(30)));
    layer0_outputs(1102) <= not((inputs(207)) or (inputs(52)));
    layer0_outputs(1103) <= not((inputs(148)) or (inputs(60)));
    layer0_outputs(1104) <= not(inputs(184));
    layer0_outputs(1105) <= (inputs(178)) and not (inputs(250));
    layer0_outputs(1106) <= '1';
    layer0_outputs(1107) <= inputs(228);
    layer0_outputs(1108) <= not((inputs(6)) or (inputs(172)));
    layer0_outputs(1109) <= (inputs(119)) xor (inputs(88));
    layer0_outputs(1110) <= (inputs(252)) xor (inputs(156));
    layer0_outputs(1111) <= '1';
    layer0_outputs(1112) <= not(inputs(130));
    layer0_outputs(1113) <= not(inputs(146)) or (inputs(111));
    layer0_outputs(1114) <= '1';
    layer0_outputs(1115) <= inputs(60);
    layer0_outputs(1116) <= (inputs(194)) or (inputs(76));
    layer0_outputs(1117) <= (inputs(241)) and not (inputs(242));
    layer0_outputs(1118) <= not(inputs(251)) or (inputs(12));
    layer0_outputs(1119) <= not((inputs(241)) and (inputs(195)));
    layer0_outputs(1120) <= '1';
    layer0_outputs(1121) <= not((inputs(163)) or (inputs(117)));
    layer0_outputs(1122) <= not(inputs(196)) or (inputs(67));
    layer0_outputs(1123) <= inputs(49);
    layer0_outputs(1124) <= (inputs(22)) xor (inputs(39));
    layer0_outputs(1125) <= inputs(57);
    layer0_outputs(1126) <= not(inputs(191));
    layer0_outputs(1127) <= (inputs(136)) or (inputs(21));
    layer0_outputs(1128) <= (inputs(239)) or (inputs(68));
    layer0_outputs(1129) <= '1';
    layer0_outputs(1130) <= '1';
    layer0_outputs(1131) <= inputs(163);
    layer0_outputs(1132) <= not(inputs(54)) or (inputs(51));
    layer0_outputs(1133) <= not((inputs(83)) or (inputs(157)));
    layer0_outputs(1134) <= not(inputs(99));
    layer0_outputs(1135) <= not((inputs(83)) or (inputs(143)));
    layer0_outputs(1136) <= not((inputs(86)) and (inputs(130)));
    layer0_outputs(1137) <= (inputs(71)) or (inputs(215));
    layer0_outputs(1138) <= not(inputs(79)) or (inputs(89));
    layer0_outputs(1139) <= (inputs(18)) and not (inputs(38));
    layer0_outputs(1140) <= (inputs(252)) and not (inputs(239));
    layer0_outputs(1141) <= not(inputs(225));
    layer0_outputs(1142) <= not(inputs(114)) or (inputs(152));
    layer0_outputs(1143) <= '0';
    layer0_outputs(1144) <= (inputs(238)) and not (inputs(232));
    layer0_outputs(1145) <= inputs(55);
    layer0_outputs(1146) <= not((inputs(217)) xor (inputs(207)));
    layer0_outputs(1147) <= '1';
    layer0_outputs(1148) <= not((inputs(145)) or (inputs(208)));
    layer0_outputs(1149) <= not(inputs(75)) or (inputs(221));
    layer0_outputs(1150) <= not(inputs(131));
    layer0_outputs(1151) <= inputs(54);
    layer0_outputs(1152) <= (inputs(88)) xor (inputs(146));
    layer0_outputs(1153) <= inputs(180);
    layer0_outputs(1154) <= not((inputs(154)) and (inputs(81)));
    layer0_outputs(1155) <= (inputs(237)) and (inputs(167));
    layer0_outputs(1156) <= '0';
    layer0_outputs(1157) <= not(inputs(66));
    layer0_outputs(1158) <= not((inputs(238)) xor (inputs(234)));
    layer0_outputs(1159) <= '1';
    layer0_outputs(1160) <= inputs(179);
    layer0_outputs(1161) <= inputs(152);
    layer0_outputs(1162) <= inputs(161);
    layer0_outputs(1163) <= '1';
    layer0_outputs(1164) <= not((inputs(104)) or (inputs(161)));
    layer0_outputs(1165) <= not(inputs(252)) or (inputs(228));
    layer0_outputs(1166) <= '1';
    layer0_outputs(1167) <= (inputs(213)) or (inputs(169));
    layer0_outputs(1168) <= not((inputs(232)) and (inputs(245)));
    layer0_outputs(1169) <= '1';
    layer0_outputs(1170) <= not(inputs(117));
    layer0_outputs(1171) <= (inputs(112)) and not (inputs(90));
    layer0_outputs(1172) <= (inputs(119)) xor (inputs(170));
    layer0_outputs(1173) <= (inputs(216)) or (inputs(203));
    layer0_outputs(1174) <= not(inputs(213));
    layer0_outputs(1175) <= not(inputs(109)) or (inputs(106));
    layer0_outputs(1176) <= not((inputs(118)) and (inputs(225)));
    layer0_outputs(1177) <= (inputs(31)) and (inputs(23));
    layer0_outputs(1178) <= '0';
    layer0_outputs(1179) <= not((inputs(194)) or (inputs(194)));
    layer0_outputs(1180) <= inputs(99);
    layer0_outputs(1181) <= not(inputs(247)) or (inputs(64));
    layer0_outputs(1182) <= not(inputs(254));
    layer0_outputs(1183) <= '0';
    layer0_outputs(1184) <= not(inputs(18));
    layer0_outputs(1185) <= not(inputs(56));
    layer0_outputs(1186) <= not(inputs(218)) or (inputs(185));
    layer0_outputs(1187) <= (inputs(144)) or (inputs(82));
    layer0_outputs(1188) <= not(inputs(242)) or (inputs(242));
    layer0_outputs(1189) <= '1';
    layer0_outputs(1190) <= inputs(200);
    layer0_outputs(1191) <= not(inputs(110));
    layer0_outputs(1192) <= (inputs(191)) and not (inputs(235));
    layer0_outputs(1193) <= inputs(174);
    layer0_outputs(1194) <= (inputs(92)) or (inputs(255));
    layer0_outputs(1195) <= inputs(116);
    layer0_outputs(1196) <= (inputs(203)) or (inputs(88));
    layer0_outputs(1197) <= not((inputs(235)) xor (inputs(22)));
    layer0_outputs(1198) <= not(inputs(229));
    layer0_outputs(1199) <= (inputs(219)) and (inputs(117));
    layer0_outputs(1200) <= not(inputs(230));
    layer0_outputs(1201) <= '0';
    layer0_outputs(1202) <= not((inputs(204)) or (inputs(64)));
    layer0_outputs(1203) <= (inputs(6)) or (inputs(123));
    layer0_outputs(1204) <= not(inputs(110));
    layer0_outputs(1205) <= '1';
    layer0_outputs(1206) <= not(inputs(224));
    layer0_outputs(1207) <= inputs(159);
    layer0_outputs(1208) <= not((inputs(212)) or (inputs(127)));
    layer0_outputs(1209) <= '1';
    layer0_outputs(1210) <= (inputs(249)) and (inputs(9));
    layer0_outputs(1211) <= (inputs(231)) and not (inputs(61));
    layer0_outputs(1212) <= not(inputs(141));
    layer0_outputs(1213) <= '0';
    layer0_outputs(1214) <= not(inputs(175)) or (inputs(109));
    layer0_outputs(1215) <= (inputs(168)) and not (inputs(176));
    layer0_outputs(1216) <= not(inputs(135));
    layer0_outputs(1217) <= not(inputs(82)) or (inputs(39));
    layer0_outputs(1218) <= inputs(39);
    layer0_outputs(1219) <= '0';
    layer0_outputs(1220) <= inputs(236);
    layer0_outputs(1221) <= (inputs(95)) and (inputs(233));
    layer0_outputs(1222) <= not(inputs(226)) or (inputs(101));
    layer0_outputs(1223) <= inputs(186);
    layer0_outputs(1224) <= (inputs(14)) xor (inputs(233));
    layer0_outputs(1225) <= (inputs(70)) or (inputs(36));
    layer0_outputs(1226) <= inputs(89);
    layer0_outputs(1227) <= not(inputs(118));
    layer0_outputs(1228) <= (inputs(57)) and (inputs(85));
    layer0_outputs(1229) <= not(inputs(145)) or (inputs(13));
    layer0_outputs(1230) <= '1';
    layer0_outputs(1231) <= inputs(71);
    layer0_outputs(1232) <= not(inputs(52)) or (inputs(242));
    layer0_outputs(1233) <= not(inputs(51)) or (inputs(33));
    layer0_outputs(1234) <= not((inputs(3)) or (inputs(120)));
    layer0_outputs(1235) <= (inputs(69)) and not (inputs(11));
    layer0_outputs(1236) <= inputs(92);
    layer0_outputs(1237) <= (inputs(38)) and not (inputs(250));
    layer0_outputs(1238) <= inputs(45);
    layer0_outputs(1239) <= inputs(49);
    layer0_outputs(1240) <= '1';
    layer0_outputs(1241) <= not(inputs(114)) or (inputs(139));
    layer0_outputs(1242) <= (inputs(254)) or (inputs(105));
    layer0_outputs(1243) <= (inputs(158)) and not (inputs(6));
    layer0_outputs(1244) <= not(inputs(154)) or (inputs(20));
    layer0_outputs(1245) <= (inputs(43)) and not (inputs(187));
    layer0_outputs(1246) <= '1';
    layer0_outputs(1247) <= not(inputs(114));
    layer0_outputs(1248) <= not(inputs(228)) or (inputs(237));
    layer0_outputs(1249) <= inputs(91);
    layer0_outputs(1250) <= not(inputs(83)) or (inputs(59));
    layer0_outputs(1251) <= not(inputs(95));
    layer0_outputs(1252) <= inputs(48);
    layer0_outputs(1253) <= not(inputs(181)) or (inputs(114));
    layer0_outputs(1254) <= (inputs(17)) and not (inputs(69));
    layer0_outputs(1255) <= '1';
    layer0_outputs(1256) <= not(inputs(41));
    layer0_outputs(1257) <= not(inputs(114));
    layer0_outputs(1258) <= (inputs(90)) and not (inputs(173));
    layer0_outputs(1259) <= not(inputs(22)) or (inputs(99));
    layer0_outputs(1260) <= (inputs(69)) and not (inputs(138));
    layer0_outputs(1261) <= not((inputs(168)) or (inputs(166)));
    layer0_outputs(1262) <= '0';
    layer0_outputs(1263) <= not((inputs(188)) or (inputs(128)));
    layer0_outputs(1264) <= inputs(114);
    layer0_outputs(1265) <= not(inputs(219));
    layer0_outputs(1266) <= (inputs(64)) xor (inputs(165));
    layer0_outputs(1267) <= not((inputs(119)) and (inputs(165)));
    layer0_outputs(1268) <= not(inputs(132)) or (inputs(139));
    layer0_outputs(1269) <= (inputs(14)) or (inputs(211));
    layer0_outputs(1270) <= not((inputs(130)) xor (inputs(136)));
    layer0_outputs(1271) <= not(inputs(215));
    layer0_outputs(1272) <= not((inputs(153)) and (inputs(69)));
    layer0_outputs(1273) <= inputs(95);
    layer0_outputs(1274) <= not(inputs(163));
    layer0_outputs(1275) <= (inputs(127)) and (inputs(164));
    layer0_outputs(1276) <= (inputs(38)) or (inputs(74));
    layer0_outputs(1277) <= inputs(227);
    layer0_outputs(1278) <= (inputs(70)) and not (inputs(96));
    layer0_outputs(1279) <= not(inputs(169));
    layer0_outputs(1280) <= not(inputs(135));
    layer0_outputs(1281) <= (inputs(94)) and not (inputs(35));
    layer0_outputs(1282) <= not(inputs(61));
    layer0_outputs(1283) <= '1';
    layer0_outputs(1284) <= not(inputs(13));
    layer0_outputs(1285) <= (inputs(45)) and not (inputs(45));
    layer0_outputs(1286) <= (inputs(242)) or (inputs(7));
    layer0_outputs(1287) <= '1';
    layer0_outputs(1288) <= not(inputs(103));
    layer0_outputs(1289) <= '1';
    layer0_outputs(1290) <= '1';
    layer0_outputs(1291) <= (inputs(111)) or (inputs(85));
    layer0_outputs(1292) <= not(inputs(129));
    layer0_outputs(1293) <= inputs(8);
    layer0_outputs(1294) <= not(inputs(39)) or (inputs(134));
    layer0_outputs(1295) <= not((inputs(90)) and (inputs(38)));
    layer0_outputs(1296) <= inputs(155);
    layer0_outputs(1297) <= (inputs(173)) and not (inputs(167));
    layer0_outputs(1298) <= (inputs(239)) and (inputs(185));
    layer0_outputs(1299) <= (inputs(45)) and not (inputs(198));
    layer0_outputs(1300) <= not(inputs(129));
    layer0_outputs(1301) <= not(inputs(252)) or (inputs(97));
    layer0_outputs(1302) <= (inputs(218)) or (inputs(194));
    layer0_outputs(1303) <= (inputs(60)) or (inputs(108));
    layer0_outputs(1304) <= inputs(234);
    layer0_outputs(1305) <= (inputs(174)) and (inputs(198));
    layer0_outputs(1306) <= not((inputs(149)) and (inputs(140)));
    layer0_outputs(1307) <= not(inputs(87));
    layer0_outputs(1308) <= not(inputs(169));
    layer0_outputs(1309) <= (inputs(242)) xor (inputs(121));
    layer0_outputs(1310) <= (inputs(7)) and (inputs(89));
    layer0_outputs(1311) <= not(inputs(62));
    layer0_outputs(1312) <= not(inputs(230)) or (inputs(9));
    layer0_outputs(1313) <= not(inputs(255));
    layer0_outputs(1314) <= (inputs(205)) and not (inputs(209));
    layer0_outputs(1315) <= inputs(76);
    layer0_outputs(1316) <= not(inputs(238));
    layer0_outputs(1317) <= not(inputs(166)) or (inputs(31));
    layer0_outputs(1318) <= inputs(213);
    layer0_outputs(1319) <= (inputs(7)) and not (inputs(241));
    layer0_outputs(1320) <= not((inputs(215)) or (inputs(93)));
    layer0_outputs(1321) <= (inputs(2)) and (inputs(247));
    layer0_outputs(1322) <= not(inputs(119)) or (inputs(189));
    layer0_outputs(1323) <= inputs(122);
    layer0_outputs(1324) <= (inputs(245)) and not (inputs(33));
    layer0_outputs(1325) <= (inputs(236)) xor (inputs(187));
    layer0_outputs(1326) <= (inputs(29)) xor (inputs(96));
    layer0_outputs(1327) <= inputs(211);
    layer0_outputs(1328) <= not((inputs(218)) and (inputs(222)));
    layer0_outputs(1329) <= inputs(254);
    layer0_outputs(1330) <= inputs(77);
    layer0_outputs(1331) <= not((inputs(40)) and (inputs(28)));
    layer0_outputs(1332) <= (inputs(149)) or (inputs(139));
    layer0_outputs(1333) <= (inputs(117)) or (inputs(174));
    layer0_outputs(1334) <= (inputs(85)) and not (inputs(18));
    layer0_outputs(1335) <= (inputs(126)) and (inputs(205));
    layer0_outputs(1336) <= '0';
    layer0_outputs(1337) <= (inputs(136)) and not (inputs(123));
    layer0_outputs(1338) <= '0';
    layer0_outputs(1339) <= not((inputs(26)) or (inputs(79)));
    layer0_outputs(1340) <= '1';
    layer0_outputs(1341) <= (inputs(223)) xor (inputs(100));
    layer0_outputs(1342) <= (inputs(117)) and not (inputs(126));
    layer0_outputs(1343) <= not(inputs(201)) or (inputs(229));
    layer0_outputs(1344) <= (inputs(25)) or (inputs(5));
    layer0_outputs(1345) <= inputs(93);
    layer0_outputs(1346) <= not(inputs(166));
    layer0_outputs(1347) <= not(inputs(96)) or (inputs(99));
    layer0_outputs(1348) <= '1';
    layer0_outputs(1349) <= (inputs(53)) or (inputs(3));
    layer0_outputs(1350) <= not(inputs(80)) or (inputs(97));
    layer0_outputs(1351) <= not((inputs(59)) or (inputs(105)));
    layer0_outputs(1352) <= (inputs(193)) and not (inputs(251));
    layer0_outputs(1353) <= '1';
    layer0_outputs(1354) <= '0';
    layer0_outputs(1355) <= (inputs(118)) and not (inputs(110));
    layer0_outputs(1356) <= not(inputs(44));
    layer0_outputs(1357) <= inputs(244);
    layer0_outputs(1358) <= not(inputs(101));
    layer0_outputs(1359) <= (inputs(36)) and (inputs(175));
    layer0_outputs(1360) <= (inputs(221)) xor (inputs(190));
    layer0_outputs(1361) <= inputs(153);
    layer0_outputs(1362) <= (inputs(103)) and not (inputs(127));
    layer0_outputs(1363) <= inputs(110);
    layer0_outputs(1364) <= inputs(84);
    layer0_outputs(1365) <= not(inputs(113));
    layer0_outputs(1366) <= (inputs(139)) or (inputs(35));
    layer0_outputs(1367) <= not((inputs(147)) and (inputs(163)));
    layer0_outputs(1368) <= (inputs(117)) and not (inputs(217));
    layer0_outputs(1369) <= not(inputs(156)) or (inputs(237));
    layer0_outputs(1370) <= not(inputs(227));
    layer0_outputs(1371) <= not((inputs(22)) and (inputs(205)));
    layer0_outputs(1372) <= inputs(98);
    layer0_outputs(1373) <= inputs(104);
    layer0_outputs(1374) <= '1';
    layer0_outputs(1375) <= '0';
    layer0_outputs(1376) <= inputs(83);
    layer0_outputs(1377) <= not((inputs(48)) or (inputs(210)));
    layer0_outputs(1378) <= (inputs(164)) or (inputs(15));
    layer0_outputs(1379) <= not(inputs(25)) or (inputs(164));
    layer0_outputs(1380) <= not((inputs(188)) and (inputs(58)));
    layer0_outputs(1381) <= '1';
    layer0_outputs(1382) <= (inputs(221)) and not (inputs(40));
    layer0_outputs(1383) <= inputs(219);
    layer0_outputs(1384) <= (inputs(31)) or (inputs(229));
    layer0_outputs(1385) <= '1';
    layer0_outputs(1386) <= (inputs(233)) xor (inputs(202));
    layer0_outputs(1387) <= not((inputs(236)) or (inputs(159)));
    layer0_outputs(1388) <= not(inputs(18)) or (inputs(118));
    layer0_outputs(1389) <= (inputs(41)) and not (inputs(222));
    layer0_outputs(1390) <= '0';
    layer0_outputs(1391) <= '0';
    layer0_outputs(1392) <= not(inputs(253)) or (inputs(102));
    layer0_outputs(1393) <= not(inputs(89));
    layer0_outputs(1394) <= (inputs(253)) and not (inputs(113));
    layer0_outputs(1395) <= not(inputs(136)) or (inputs(0));
    layer0_outputs(1396) <= (inputs(16)) xor (inputs(161));
    layer0_outputs(1397) <= '1';
    layer0_outputs(1398) <= inputs(76);
    layer0_outputs(1399) <= not(inputs(181)) or (inputs(184));
    layer0_outputs(1400) <= not(inputs(97)) or (inputs(183));
    layer0_outputs(1401) <= not((inputs(68)) or (inputs(247)));
    layer0_outputs(1402) <= not((inputs(210)) or (inputs(38)));
    layer0_outputs(1403) <= (inputs(88)) and not (inputs(80));
    layer0_outputs(1404) <= inputs(244);
    layer0_outputs(1405) <= not((inputs(193)) and (inputs(111)));
    layer0_outputs(1406) <= (inputs(36)) and not (inputs(3));
    layer0_outputs(1407) <= inputs(46);
    layer0_outputs(1408) <= '1';
    layer0_outputs(1409) <= inputs(93);
    layer0_outputs(1410) <= inputs(187);
    layer0_outputs(1411) <= (inputs(46)) and (inputs(34));
    layer0_outputs(1412) <= '0';
    layer0_outputs(1413) <= (inputs(225)) and not (inputs(44));
    layer0_outputs(1414) <= (inputs(116)) xor (inputs(2));
    layer0_outputs(1415) <= '1';
    layer0_outputs(1416) <= not(inputs(115));
    layer0_outputs(1417) <= '0';
    layer0_outputs(1418) <= (inputs(148)) and not (inputs(240));
    layer0_outputs(1419) <= not(inputs(146)) or (inputs(174));
    layer0_outputs(1420) <= (inputs(66)) or (inputs(5));
    layer0_outputs(1421) <= not(inputs(163));
    layer0_outputs(1422) <= not((inputs(86)) and (inputs(28)));
    layer0_outputs(1423) <= (inputs(210)) or (inputs(247));
    layer0_outputs(1424) <= (inputs(113)) or (inputs(147));
    layer0_outputs(1425) <= not(inputs(180));
    layer0_outputs(1426) <= not(inputs(209));
    layer0_outputs(1427) <= not((inputs(253)) or (inputs(186)));
    layer0_outputs(1428) <= (inputs(188)) and (inputs(177));
    layer0_outputs(1429) <= (inputs(98)) or (inputs(43));
    layer0_outputs(1430) <= (inputs(96)) and (inputs(109));
    layer0_outputs(1431) <= (inputs(95)) xor (inputs(76));
    layer0_outputs(1432) <= '0';
    layer0_outputs(1433) <= (inputs(206)) or (inputs(123));
    layer0_outputs(1434) <= not((inputs(84)) or (inputs(94)));
    layer0_outputs(1435) <= not(inputs(169)) or (inputs(152));
    layer0_outputs(1436) <= '0';
    layer0_outputs(1437) <= (inputs(236)) or (inputs(172));
    layer0_outputs(1438) <= inputs(135);
    layer0_outputs(1439) <= not((inputs(54)) or (inputs(157)));
    layer0_outputs(1440) <= not(inputs(110));
    layer0_outputs(1441) <= not(inputs(138)) or (inputs(91));
    layer0_outputs(1442) <= '0';
    layer0_outputs(1443) <= (inputs(169)) and not (inputs(13));
    layer0_outputs(1444) <= '1';
    layer0_outputs(1445) <= '1';
    layer0_outputs(1446) <= not((inputs(131)) and (inputs(150)));
    layer0_outputs(1447) <= not((inputs(235)) xor (inputs(162)));
    layer0_outputs(1448) <= not(inputs(193)) or (inputs(34));
    layer0_outputs(1449) <= (inputs(168)) and not (inputs(107));
    layer0_outputs(1450) <= not(inputs(176)) or (inputs(70));
    layer0_outputs(1451) <= inputs(72);
    layer0_outputs(1452) <= '0';
    layer0_outputs(1453) <= (inputs(19)) and not (inputs(16));
    layer0_outputs(1454) <= not(inputs(23));
    layer0_outputs(1455) <= inputs(156);
    layer0_outputs(1456) <= inputs(108);
    layer0_outputs(1457) <= not((inputs(16)) and (inputs(65)));
    layer0_outputs(1458) <= '1';
    layer0_outputs(1459) <= not(inputs(197)) or (inputs(1));
    layer0_outputs(1460) <= not(inputs(43));
    layer0_outputs(1461) <= not(inputs(8));
    layer0_outputs(1462) <= not(inputs(37));
    layer0_outputs(1463) <= '1';
    layer0_outputs(1464) <= (inputs(14)) and (inputs(14));
    layer0_outputs(1465) <= inputs(48);
    layer0_outputs(1466) <= not(inputs(67)) or (inputs(245));
    layer0_outputs(1467) <= inputs(166);
    layer0_outputs(1468) <= (inputs(82)) and not (inputs(82));
    layer0_outputs(1469) <= '1';
    layer0_outputs(1470) <= (inputs(72)) and (inputs(144));
    layer0_outputs(1471) <= (inputs(85)) and not (inputs(124));
    layer0_outputs(1472) <= (inputs(196)) and not (inputs(105));
    layer0_outputs(1473) <= not(inputs(53)) or (inputs(181));
    layer0_outputs(1474) <= not(inputs(167));
    layer0_outputs(1475) <= inputs(121);
    layer0_outputs(1476) <= '1';
    layer0_outputs(1477) <= not((inputs(156)) or (inputs(9)));
    layer0_outputs(1478) <= inputs(7);
    layer0_outputs(1479) <= not((inputs(153)) or (inputs(165)));
    layer0_outputs(1480) <= inputs(24);
    layer0_outputs(1481) <= (inputs(49)) and not (inputs(17));
    layer0_outputs(1482) <= inputs(59);
    layer0_outputs(1483) <= not((inputs(61)) and (inputs(233)));
    layer0_outputs(1484) <= '1';
    layer0_outputs(1485) <= (inputs(33)) and (inputs(175));
    layer0_outputs(1486) <= (inputs(112)) and not (inputs(54));
    layer0_outputs(1487) <= not(inputs(168)) or (inputs(109));
    layer0_outputs(1488) <= inputs(232);
    layer0_outputs(1489) <= not((inputs(13)) or (inputs(169)));
    layer0_outputs(1490) <= '0';
    layer0_outputs(1491) <= not(inputs(7)) or (inputs(196));
    layer0_outputs(1492) <= not(inputs(52));
    layer0_outputs(1493) <= not(inputs(98));
    layer0_outputs(1494) <= (inputs(88)) and not (inputs(117));
    layer0_outputs(1495) <= '0';
    layer0_outputs(1496) <= (inputs(154)) or (inputs(173));
    layer0_outputs(1497) <= not(inputs(10));
    layer0_outputs(1498) <= (inputs(48)) or (inputs(54));
    layer0_outputs(1499) <= not(inputs(179)) or (inputs(14));
    layer0_outputs(1500) <= not((inputs(32)) or (inputs(134)));
    layer0_outputs(1501) <= '0';
    layer0_outputs(1502) <= (inputs(104)) or (inputs(151));
    layer0_outputs(1503) <= (inputs(50)) and (inputs(142));
    layer0_outputs(1504) <= not(inputs(197));
    layer0_outputs(1505) <= (inputs(84)) and (inputs(173));
    layer0_outputs(1506) <= inputs(61);
    layer0_outputs(1507) <= not(inputs(190)) or (inputs(13));
    layer0_outputs(1508) <= not(inputs(135));
    layer0_outputs(1509) <= '0';
    layer0_outputs(1510) <= not(inputs(199));
    layer0_outputs(1511) <= not(inputs(143)) or (inputs(205));
    layer0_outputs(1512) <= not(inputs(143));
    layer0_outputs(1513) <= not(inputs(226)) or (inputs(194));
    layer0_outputs(1514) <= (inputs(115)) and not (inputs(137));
    layer0_outputs(1515) <= inputs(77);
    layer0_outputs(1516) <= (inputs(194)) and (inputs(136));
    layer0_outputs(1517) <= '1';
    layer0_outputs(1518) <= not(inputs(4)) or (inputs(142));
    layer0_outputs(1519) <= not(inputs(112)) or (inputs(14));
    layer0_outputs(1520) <= not(inputs(163)) or (inputs(2));
    layer0_outputs(1521) <= (inputs(8)) or (inputs(206));
    layer0_outputs(1522) <= (inputs(86)) and not (inputs(191));
    layer0_outputs(1523) <= '1';
    layer0_outputs(1524) <= (inputs(230)) and not (inputs(225));
    layer0_outputs(1525) <= not(inputs(97));
    layer0_outputs(1526) <= not(inputs(103)) or (inputs(224));
    layer0_outputs(1527) <= not(inputs(100));
    layer0_outputs(1528) <= not((inputs(86)) and (inputs(247)));
    layer0_outputs(1529) <= '1';
    layer0_outputs(1530) <= inputs(75);
    layer0_outputs(1531) <= not((inputs(110)) or (inputs(127)));
    layer0_outputs(1532) <= '1';
    layer0_outputs(1533) <= not(inputs(188));
    layer0_outputs(1534) <= not((inputs(226)) and (inputs(216)));
    layer0_outputs(1535) <= not((inputs(125)) or (inputs(206)));
    layer0_outputs(1536) <= inputs(8);
    layer0_outputs(1537) <= not(inputs(240)) or (inputs(137));
    layer0_outputs(1538) <= inputs(111);
    layer0_outputs(1539) <= not(inputs(180));
    layer0_outputs(1540) <= '1';
    layer0_outputs(1541) <= not(inputs(89));
    layer0_outputs(1542) <= not(inputs(188)) or (inputs(201));
    layer0_outputs(1543) <= not(inputs(5)) or (inputs(52));
    layer0_outputs(1544) <= inputs(97);
    layer0_outputs(1545) <= inputs(200);
    layer0_outputs(1546) <= (inputs(81)) xor (inputs(30));
    layer0_outputs(1547) <= '1';
    layer0_outputs(1548) <= (inputs(156)) and not (inputs(252));
    layer0_outputs(1549) <= '0';
    layer0_outputs(1550) <= (inputs(255)) or (inputs(90));
    layer0_outputs(1551) <= (inputs(223)) and (inputs(68));
    layer0_outputs(1552) <= (inputs(4)) and not (inputs(10));
    layer0_outputs(1553) <= not(inputs(44));
    layer0_outputs(1554) <= (inputs(168)) and (inputs(251));
    layer0_outputs(1555) <= (inputs(214)) and not (inputs(74));
    layer0_outputs(1556) <= inputs(195);
    layer0_outputs(1557) <= not(inputs(113));
    layer0_outputs(1558) <= not(inputs(112));
    layer0_outputs(1559) <= '1';
    layer0_outputs(1560) <= '1';
    layer0_outputs(1561) <= (inputs(242)) and not (inputs(97));
    layer0_outputs(1562) <= (inputs(165)) or (inputs(2));
    layer0_outputs(1563) <= not(inputs(160)) or (inputs(157));
    layer0_outputs(1564) <= (inputs(208)) and (inputs(31));
    layer0_outputs(1565) <= inputs(140);
    layer0_outputs(1566) <= not(inputs(70));
    layer0_outputs(1567) <= (inputs(219)) and not (inputs(90));
    layer0_outputs(1568) <= '1';
    layer0_outputs(1569) <= '0';
    layer0_outputs(1570) <= '0';
    layer0_outputs(1571) <= (inputs(135)) and not (inputs(167));
    layer0_outputs(1572) <= '0';
    layer0_outputs(1573) <= inputs(161);
    layer0_outputs(1574) <= not(inputs(12));
    layer0_outputs(1575) <= (inputs(91)) and not (inputs(241));
    layer0_outputs(1576) <= inputs(20);
    layer0_outputs(1577) <= not((inputs(11)) or (inputs(250)));
    layer0_outputs(1578) <= inputs(10);
    layer0_outputs(1579) <= not(inputs(135));
    layer0_outputs(1580) <= not((inputs(109)) or (inputs(107)));
    layer0_outputs(1581) <= (inputs(226)) and not (inputs(168));
    layer0_outputs(1582) <= not((inputs(159)) and (inputs(6)));
    layer0_outputs(1583) <= not((inputs(219)) and (inputs(70)));
    layer0_outputs(1584) <= not(inputs(18));
    layer0_outputs(1585) <= not(inputs(116)) or (inputs(25));
    layer0_outputs(1586) <= '0';
    layer0_outputs(1587) <= inputs(120);
    layer0_outputs(1588) <= '0';
    layer0_outputs(1589) <= not((inputs(89)) and (inputs(97)));
    layer0_outputs(1590) <= (inputs(133)) and not (inputs(49));
    layer0_outputs(1591) <= (inputs(201)) xor (inputs(209));
    layer0_outputs(1592) <= '0';
    layer0_outputs(1593) <= (inputs(70)) and not (inputs(30));
    layer0_outputs(1594) <= (inputs(12)) and not (inputs(126));
    layer0_outputs(1595) <= not(inputs(169)) or (inputs(92));
    layer0_outputs(1596) <= not(inputs(27)) or (inputs(211));
    layer0_outputs(1597) <= not(inputs(19));
    layer0_outputs(1598) <= (inputs(230)) or (inputs(239));
    layer0_outputs(1599) <= (inputs(101)) or (inputs(190));
    layer0_outputs(1600) <= (inputs(75)) or (inputs(47));
    layer0_outputs(1601) <= not(inputs(149));
    layer0_outputs(1602) <= '0';
    layer0_outputs(1603) <= inputs(211);
    layer0_outputs(1604) <= not(inputs(164));
    layer0_outputs(1605) <= inputs(222);
    layer0_outputs(1606) <= '0';
    layer0_outputs(1607) <= (inputs(171)) and not (inputs(91));
    layer0_outputs(1608) <= not(inputs(162));
    layer0_outputs(1609) <= not(inputs(35));
    layer0_outputs(1610) <= (inputs(13)) and not (inputs(251));
    layer0_outputs(1611) <= inputs(196);
    layer0_outputs(1612) <= inputs(231);
    layer0_outputs(1613) <= not(inputs(153));
    layer0_outputs(1614) <= inputs(168);
    layer0_outputs(1615) <= not((inputs(188)) and (inputs(201)));
    layer0_outputs(1616) <= inputs(66);
    layer0_outputs(1617) <= not((inputs(157)) and (inputs(200)));
    layer0_outputs(1618) <= '1';
    layer0_outputs(1619) <= inputs(186);
    layer0_outputs(1620) <= '0';
    layer0_outputs(1621) <= inputs(255);
    layer0_outputs(1622) <= (inputs(21)) and not (inputs(211));
    layer0_outputs(1623) <= (inputs(41)) or (inputs(190));
    layer0_outputs(1624) <= '1';
    layer0_outputs(1625) <= inputs(192);
    layer0_outputs(1626) <= (inputs(44)) xor (inputs(159));
    layer0_outputs(1627) <= '0';
    layer0_outputs(1628) <= not(inputs(206)) or (inputs(175));
    layer0_outputs(1629) <= (inputs(12)) and not (inputs(62));
    layer0_outputs(1630) <= '0';
    layer0_outputs(1631) <= (inputs(249)) or (inputs(115));
    layer0_outputs(1632) <= (inputs(64)) xor (inputs(200));
    layer0_outputs(1633) <= not(inputs(135));
    layer0_outputs(1634) <= not(inputs(112));
    layer0_outputs(1635) <= inputs(121);
    layer0_outputs(1636) <= not(inputs(57)) or (inputs(237));
    layer0_outputs(1637) <= (inputs(160)) and not (inputs(155));
    layer0_outputs(1638) <= (inputs(105)) and (inputs(172));
    layer0_outputs(1639) <= (inputs(167)) and (inputs(138));
    layer0_outputs(1640) <= not(inputs(188)) or (inputs(199));
    layer0_outputs(1641) <= '0';
    layer0_outputs(1642) <= not(inputs(25));
    layer0_outputs(1643) <= (inputs(1)) and (inputs(198));
    layer0_outputs(1644) <= inputs(83);
    layer0_outputs(1645) <= inputs(81);
    layer0_outputs(1646) <= not((inputs(249)) or (inputs(168)));
    layer0_outputs(1647) <= '1';
    layer0_outputs(1648) <= not((inputs(159)) xor (inputs(53)));
    layer0_outputs(1649) <= (inputs(151)) and not (inputs(219));
    layer0_outputs(1650) <= not(inputs(96)) or (inputs(98));
    layer0_outputs(1651) <= '1';
    layer0_outputs(1652) <= not(inputs(47)) or (inputs(246));
    layer0_outputs(1653) <= not((inputs(78)) or (inputs(25)));
    layer0_outputs(1654) <= (inputs(32)) and not (inputs(248));
    layer0_outputs(1655) <= '1';
    layer0_outputs(1656) <= not((inputs(220)) or (inputs(33)));
    layer0_outputs(1657) <= not(inputs(105)) or (inputs(40));
    layer0_outputs(1658) <= inputs(208);
    layer0_outputs(1659) <= '0';
    layer0_outputs(1660) <= '0';
    layer0_outputs(1661) <= not(inputs(195));
    layer0_outputs(1662) <= (inputs(28)) and (inputs(215));
    layer0_outputs(1663) <= not((inputs(157)) or (inputs(13)));
    layer0_outputs(1664) <= (inputs(72)) or (inputs(106));
    layer0_outputs(1665) <= not(inputs(163)) or (inputs(147));
    layer0_outputs(1666) <= not((inputs(227)) and (inputs(232)));
    layer0_outputs(1667) <= not((inputs(253)) or (inputs(120)));
    layer0_outputs(1668) <= not(inputs(85)) or (inputs(4));
    layer0_outputs(1669) <= not((inputs(177)) or (inputs(197)));
    layer0_outputs(1670) <= not(inputs(131));
    layer0_outputs(1671) <= not(inputs(80));
    layer0_outputs(1672) <= not(inputs(227));
    layer0_outputs(1673) <= (inputs(158)) or (inputs(195));
    layer0_outputs(1674) <= not(inputs(114));
    layer0_outputs(1675) <= not(inputs(28)) or (inputs(197));
    layer0_outputs(1676) <= not((inputs(2)) or (inputs(2)));
    layer0_outputs(1677) <= (inputs(118)) xor (inputs(149));
    layer0_outputs(1678) <= not((inputs(95)) and (inputs(23)));
    layer0_outputs(1679) <= inputs(118);
    layer0_outputs(1680) <= '0';
    layer0_outputs(1681) <= not((inputs(214)) or (inputs(207)));
    layer0_outputs(1682) <= not(inputs(166)) or (inputs(222));
    layer0_outputs(1683) <= '1';
    layer0_outputs(1684) <= not(inputs(172)) or (inputs(97));
    layer0_outputs(1685) <= not(inputs(195));
    layer0_outputs(1686) <= '1';
    layer0_outputs(1687) <= '1';
    layer0_outputs(1688) <= not(inputs(15));
    layer0_outputs(1689) <= (inputs(128)) and not (inputs(61));
    layer0_outputs(1690) <= '0';
    layer0_outputs(1691) <= '1';
    layer0_outputs(1692) <= not(inputs(221));
    layer0_outputs(1693) <= not((inputs(71)) and (inputs(223)));
    layer0_outputs(1694) <= (inputs(226)) and (inputs(145));
    layer0_outputs(1695) <= inputs(162);
    layer0_outputs(1696) <= not(inputs(143));
    layer0_outputs(1697) <= '0';
    layer0_outputs(1698) <= not(inputs(200));
    layer0_outputs(1699) <= not(inputs(208)) or (inputs(223));
    layer0_outputs(1700) <= '0';
    layer0_outputs(1701) <= not((inputs(84)) and (inputs(23)));
    layer0_outputs(1702) <= (inputs(218)) or (inputs(10));
    layer0_outputs(1703) <= not(inputs(110)) or (inputs(171));
    layer0_outputs(1704) <= not((inputs(143)) or (inputs(165)));
    layer0_outputs(1705) <= inputs(122);
    layer0_outputs(1706) <= (inputs(86)) or (inputs(9));
    layer0_outputs(1707) <= not((inputs(212)) or (inputs(195)));
    layer0_outputs(1708) <= '0';
    layer0_outputs(1709) <= inputs(14);
    layer0_outputs(1710) <= inputs(245);
    layer0_outputs(1711) <= not(inputs(99));
    layer0_outputs(1712) <= (inputs(249)) or (inputs(146));
    layer0_outputs(1713) <= (inputs(237)) or (inputs(161));
    layer0_outputs(1714) <= not(inputs(48));
    layer0_outputs(1715) <= (inputs(148)) and not (inputs(11));
    layer0_outputs(1716) <= inputs(5);
    layer0_outputs(1717) <= '0';
    layer0_outputs(1718) <= inputs(150);
    layer0_outputs(1719) <= inputs(48);
    layer0_outputs(1720) <= (inputs(93)) and not (inputs(26));
    layer0_outputs(1721) <= (inputs(64)) and not (inputs(99));
    layer0_outputs(1722) <= not((inputs(122)) and (inputs(223)));
    layer0_outputs(1723) <= not(inputs(140));
    layer0_outputs(1724) <= (inputs(255)) and not (inputs(72));
    layer0_outputs(1725) <= inputs(205);
    layer0_outputs(1726) <= (inputs(150)) or (inputs(204));
    layer0_outputs(1727) <= (inputs(56)) and not (inputs(178));
    layer0_outputs(1728) <= '1';
    layer0_outputs(1729) <= not(inputs(11)) or (inputs(36));
    layer0_outputs(1730) <= inputs(222);
    layer0_outputs(1731) <= inputs(45);
    layer0_outputs(1732) <= inputs(181);
    layer0_outputs(1733) <= inputs(232);
    layer0_outputs(1734) <= not((inputs(33)) and (inputs(131)));
    layer0_outputs(1735) <= not((inputs(32)) or (inputs(170)));
    layer0_outputs(1736) <= (inputs(43)) and (inputs(83));
    layer0_outputs(1737) <= inputs(128);
    layer0_outputs(1738) <= not(inputs(237));
    layer0_outputs(1739) <= (inputs(178)) and (inputs(51));
    layer0_outputs(1740) <= '1';
    layer0_outputs(1741) <= '1';
    layer0_outputs(1742) <= not(inputs(246));
    layer0_outputs(1743) <= '0';
    layer0_outputs(1744) <= (inputs(106)) or (inputs(122));
    layer0_outputs(1745) <= not(inputs(94));
    layer0_outputs(1746) <= (inputs(193)) and (inputs(241));
    layer0_outputs(1747) <= not((inputs(66)) or (inputs(100)));
    layer0_outputs(1748) <= not((inputs(5)) and (inputs(61)));
    layer0_outputs(1749) <= inputs(37);
    layer0_outputs(1750) <= not((inputs(166)) or (inputs(165)));
    layer0_outputs(1751) <= not((inputs(233)) or (inputs(143)));
    layer0_outputs(1752) <= inputs(137);
    layer0_outputs(1753) <= (inputs(200)) and not (inputs(211));
    layer0_outputs(1754) <= '1';
    layer0_outputs(1755) <= (inputs(227)) or (inputs(165));
    layer0_outputs(1756) <= not(inputs(192));
    layer0_outputs(1757) <= not(inputs(69));
    layer0_outputs(1758) <= not((inputs(16)) or (inputs(15)));
    layer0_outputs(1759) <= not(inputs(72));
    layer0_outputs(1760) <= not((inputs(10)) or (inputs(142)));
    layer0_outputs(1761) <= inputs(167);
    layer0_outputs(1762) <= (inputs(72)) xor (inputs(210));
    layer0_outputs(1763) <= not((inputs(238)) and (inputs(227)));
    layer0_outputs(1764) <= not((inputs(129)) and (inputs(1)));
    layer0_outputs(1765) <= '0';
    layer0_outputs(1766) <= not((inputs(155)) and (inputs(184)));
    layer0_outputs(1767) <= '0';
    layer0_outputs(1768) <= '1';
    layer0_outputs(1769) <= (inputs(2)) and not (inputs(3));
    layer0_outputs(1770) <= inputs(17);
    layer0_outputs(1771) <= '1';
    layer0_outputs(1772) <= (inputs(245)) xor (inputs(194));
    layer0_outputs(1773) <= '1';
    layer0_outputs(1774) <= (inputs(255)) and not (inputs(57));
    layer0_outputs(1775) <= (inputs(26)) or (inputs(147));
    layer0_outputs(1776) <= not(inputs(252));
    layer0_outputs(1777) <= (inputs(16)) xor (inputs(205));
    layer0_outputs(1778) <= inputs(8);
    layer0_outputs(1779) <= not((inputs(63)) or (inputs(184)));
    layer0_outputs(1780) <= not(inputs(98));
    layer0_outputs(1781) <= '1';
    layer0_outputs(1782) <= not((inputs(176)) or (inputs(130)));
    layer0_outputs(1783) <= inputs(147);
    layer0_outputs(1784) <= not((inputs(202)) or (inputs(201)));
    layer0_outputs(1785) <= '0';
    layer0_outputs(1786) <= '0';
    layer0_outputs(1787) <= inputs(179);
    layer0_outputs(1788) <= inputs(69);
    layer0_outputs(1789) <= (inputs(177)) and not (inputs(148));
    layer0_outputs(1790) <= not(inputs(115));
    layer0_outputs(1791) <= '0';
    layer0_outputs(1792) <= inputs(183);
    layer0_outputs(1793) <= not(inputs(226));
    layer0_outputs(1794) <= (inputs(121)) and not (inputs(131));
    layer0_outputs(1795) <= not((inputs(58)) or (inputs(131)));
    layer0_outputs(1796) <= inputs(202);
    layer0_outputs(1797) <= not(inputs(189)) or (inputs(113));
    layer0_outputs(1798) <= inputs(141);
    layer0_outputs(1799) <= '0';
    layer0_outputs(1800) <= not(inputs(60));
    layer0_outputs(1801) <= (inputs(182)) or (inputs(178));
    layer0_outputs(1802) <= not((inputs(156)) or (inputs(28)));
    layer0_outputs(1803) <= not(inputs(207));
    layer0_outputs(1804) <= inputs(75);
    layer0_outputs(1805) <= not((inputs(189)) xor (inputs(18)));
    layer0_outputs(1806) <= not(inputs(140)) or (inputs(137));
    layer0_outputs(1807) <= inputs(144);
    layer0_outputs(1808) <= not(inputs(38));
    layer0_outputs(1809) <= not(inputs(66)) or (inputs(8));
    layer0_outputs(1810) <= not(inputs(107));
    layer0_outputs(1811) <= not((inputs(12)) or (inputs(8)));
    layer0_outputs(1812) <= inputs(47);
    layer0_outputs(1813) <= not(inputs(228));
    layer0_outputs(1814) <= '1';
    layer0_outputs(1815) <= '1';
    layer0_outputs(1816) <= not(inputs(14));
    layer0_outputs(1817) <= not((inputs(223)) and (inputs(87)));
    layer0_outputs(1818) <= '1';
    layer0_outputs(1819) <= not(inputs(104));
    layer0_outputs(1820) <= '0';
    layer0_outputs(1821) <= not((inputs(8)) or (inputs(214)));
    layer0_outputs(1822) <= not((inputs(221)) or (inputs(235)));
    layer0_outputs(1823) <= (inputs(53)) and not (inputs(217));
    layer0_outputs(1824) <= '0';
    layer0_outputs(1825) <= '1';
    layer0_outputs(1826) <= inputs(83);
    layer0_outputs(1827) <= (inputs(74)) and (inputs(55));
    layer0_outputs(1828) <= (inputs(16)) or (inputs(147));
    layer0_outputs(1829) <= not(inputs(222)) or (inputs(180));
    layer0_outputs(1830) <= '0';
    layer0_outputs(1831) <= (inputs(194)) or (inputs(182));
    layer0_outputs(1832) <= not(inputs(163));
    layer0_outputs(1833) <= not(inputs(29)) or (inputs(58));
    layer0_outputs(1834) <= not(inputs(27));
    layer0_outputs(1835) <= not(inputs(91));
    layer0_outputs(1836) <= not((inputs(163)) or (inputs(201)));
    layer0_outputs(1837) <= inputs(86);
    layer0_outputs(1838) <= inputs(207);
    layer0_outputs(1839) <= (inputs(84)) or (inputs(24));
    layer0_outputs(1840) <= '0';
    layer0_outputs(1841) <= not((inputs(253)) or (inputs(25)));
    layer0_outputs(1842) <= (inputs(46)) or (inputs(65));
    layer0_outputs(1843) <= inputs(218);
    layer0_outputs(1844) <= inputs(20);
    layer0_outputs(1845) <= not(inputs(178)) or (inputs(64));
    layer0_outputs(1846) <= not((inputs(108)) or (inputs(45)));
    layer0_outputs(1847) <= (inputs(192)) xor (inputs(223));
    layer0_outputs(1848) <= (inputs(236)) and (inputs(209));
    layer0_outputs(1849) <= '1';
    layer0_outputs(1850) <= not(inputs(240)) or (inputs(0));
    layer0_outputs(1851) <= '0';
    layer0_outputs(1852) <= (inputs(234)) or (inputs(107));
    layer0_outputs(1853) <= (inputs(143)) or (inputs(21));
    layer0_outputs(1854) <= inputs(203);
    layer0_outputs(1855) <= not((inputs(191)) or (inputs(173)));
    layer0_outputs(1856) <= not(inputs(234));
    layer0_outputs(1857) <= not(inputs(238));
    layer0_outputs(1858) <= not(inputs(168)) or (inputs(233));
    layer0_outputs(1859) <= not((inputs(246)) or (inputs(174)));
    layer0_outputs(1860) <= '0';
    layer0_outputs(1861) <= '1';
    layer0_outputs(1862) <= (inputs(200)) and not (inputs(37));
    layer0_outputs(1863) <= (inputs(149)) or (inputs(209));
    layer0_outputs(1864) <= not(inputs(99));
    layer0_outputs(1865) <= not((inputs(36)) and (inputs(169)));
    layer0_outputs(1866) <= (inputs(148)) or (inputs(131));
    layer0_outputs(1867) <= '1';
    layer0_outputs(1868) <= '0';
    layer0_outputs(1869) <= (inputs(110)) or (inputs(163));
    layer0_outputs(1870) <= (inputs(57)) and not (inputs(89));
    layer0_outputs(1871) <= not(inputs(168));
    layer0_outputs(1872) <= '1';
    layer0_outputs(1873) <= not((inputs(197)) and (inputs(45)));
    layer0_outputs(1874) <= not(inputs(22));
    layer0_outputs(1875) <= inputs(104);
    layer0_outputs(1876) <= not(inputs(146));
    layer0_outputs(1877) <= not((inputs(94)) and (inputs(203)));
    layer0_outputs(1878) <= inputs(78);
    layer0_outputs(1879) <= not(inputs(72));
    layer0_outputs(1880) <= inputs(241);
    layer0_outputs(1881) <= not((inputs(22)) or (inputs(17)));
    layer0_outputs(1882) <= (inputs(33)) and not (inputs(201));
    layer0_outputs(1883) <= not(inputs(221));
    layer0_outputs(1884) <= not(inputs(169)) or (inputs(101));
    layer0_outputs(1885) <= (inputs(120)) and (inputs(131));
    layer0_outputs(1886) <= '1';
    layer0_outputs(1887) <= not((inputs(74)) xor (inputs(255)));
    layer0_outputs(1888) <= (inputs(241)) or (inputs(7));
    layer0_outputs(1889) <= not((inputs(84)) or (inputs(63)));
    layer0_outputs(1890) <= not(inputs(80)) or (inputs(39));
    layer0_outputs(1891) <= not(inputs(161));
    layer0_outputs(1892) <= (inputs(165)) and (inputs(100));
    layer0_outputs(1893) <= not(inputs(152));
    layer0_outputs(1894) <= not((inputs(181)) or (inputs(137)));
    layer0_outputs(1895) <= not(inputs(162));
    layer0_outputs(1896) <= not(inputs(165));
    layer0_outputs(1897) <= '1';
    layer0_outputs(1898) <= not((inputs(144)) or (inputs(100)));
    layer0_outputs(1899) <= not(inputs(15));
    layer0_outputs(1900) <= not(inputs(251)) or (inputs(100));
    layer0_outputs(1901) <= not(inputs(218));
    layer0_outputs(1902) <= (inputs(201)) and not (inputs(122));
    layer0_outputs(1903) <= '0';
    layer0_outputs(1904) <= inputs(76);
    layer0_outputs(1905) <= (inputs(130)) or (inputs(165));
    layer0_outputs(1906) <= not(inputs(149));
    layer0_outputs(1907) <= not(inputs(67));
    layer0_outputs(1908) <= inputs(112);
    layer0_outputs(1909) <= (inputs(82)) and not (inputs(184));
    layer0_outputs(1910) <= '0';
    layer0_outputs(1911) <= '0';
    layer0_outputs(1912) <= '0';
    layer0_outputs(1913) <= not((inputs(191)) or (inputs(235)));
    layer0_outputs(1914) <= '1';
    layer0_outputs(1915) <= (inputs(249)) and (inputs(172));
    layer0_outputs(1916) <= inputs(93);
    layer0_outputs(1917) <= (inputs(213)) or (inputs(143));
    layer0_outputs(1918) <= not(inputs(202)) or (inputs(98));
    layer0_outputs(1919) <= (inputs(211)) and not (inputs(60));
    layer0_outputs(1920) <= not((inputs(84)) or (inputs(78)));
    layer0_outputs(1921) <= not(inputs(97));
    layer0_outputs(1922) <= (inputs(138)) xor (inputs(190));
    layer0_outputs(1923) <= (inputs(45)) and (inputs(131));
    layer0_outputs(1924) <= (inputs(176)) and (inputs(19));
    layer0_outputs(1925) <= not(inputs(151)) or (inputs(139));
    layer0_outputs(1926) <= not(inputs(218)) or (inputs(95));
    layer0_outputs(1927) <= not((inputs(41)) or (inputs(148)));
    layer0_outputs(1928) <= not(inputs(102)) or (inputs(109));
    layer0_outputs(1929) <= '0';
    layer0_outputs(1930) <= inputs(183);
    layer0_outputs(1931) <= (inputs(196)) or (inputs(148));
    layer0_outputs(1932) <= (inputs(79)) or (inputs(102));
    layer0_outputs(1933) <= inputs(105);
    layer0_outputs(1934) <= (inputs(0)) and not (inputs(115));
    layer0_outputs(1935) <= inputs(105);
    layer0_outputs(1936) <= inputs(244);
    layer0_outputs(1937) <= not(inputs(12)) or (inputs(245));
    layer0_outputs(1938) <= inputs(224);
    layer0_outputs(1939) <= '1';
    layer0_outputs(1940) <= not((inputs(51)) or (inputs(254)));
    layer0_outputs(1941) <= '0';
    layer0_outputs(1942) <= inputs(216);
    layer0_outputs(1943) <= inputs(103);
    layer0_outputs(1944) <= not(inputs(91)) or (inputs(70));
    layer0_outputs(1945) <= '1';
    layer0_outputs(1946) <= not(inputs(148));
    layer0_outputs(1947) <= inputs(131);
    layer0_outputs(1948) <= not((inputs(34)) or (inputs(92)));
    layer0_outputs(1949) <= '1';
    layer0_outputs(1950) <= not(inputs(103)) or (inputs(17));
    layer0_outputs(1951) <= (inputs(111)) or (inputs(179));
    layer0_outputs(1952) <= (inputs(141)) and not (inputs(253));
    layer0_outputs(1953) <= (inputs(79)) and not (inputs(225));
    layer0_outputs(1954) <= inputs(119);
    layer0_outputs(1955) <= (inputs(93)) and (inputs(42));
    layer0_outputs(1956) <= inputs(181);
    layer0_outputs(1957) <= (inputs(80)) xor (inputs(0));
    layer0_outputs(1958) <= '0';
    layer0_outputs(1959) <= '0';
    layer0_outputs(1960) <= (inputs(110)) xor (inputs(219));
    layer0_outputs(1961) <= not(inputs(84));
    layer0_outputs(1962) <= '1';
    layer0_outputs(1963) <= not(inputs(194)) or (inputs(235));
    layer0_outputs(1964) <= inputs(194);
    layer0_outputs(1965) <= not((inputs(21)) or (inputs(19)));
    layer0_outputs(1966) <= '1';
    layer0_outputs(1967) <= inputs(173);
    layer0_outputs(1968) <= not(inputs(51));
    layer0_outputs(1969) <= (inputs(114)) and not (inputs(218));
    layer0_outputs(1970) <= not((inputs(127)) or (inputs(194)));
    layer0_outputs(1971) <= not(inputs(146));
    layer0_outputs(1972) <= (inputs(6)) or (inputs(75));
    layer0_outputs(1973) <= (inputs(71)) and (inputs(40));
    layer0_outputs(1974) <= not(inputs(20)) or (inputs(65));
    layer0_outputs(1975) <= inputs(136);
    layer0_outputs(1976) <= not((inputs(116)) or (inputs(61)));
    layer0_outputs(1977) <= not(inputs(227)) or (inputs(239));
    layer0_outputs(1978) <= not(inputs(78)) or (inputs(24));
    layer0_outputs(1979) <= not((inputs(217)) or (inputs(116)));
    layer0_outputs(1980) <= not(inputs(228)) or (inputs(136));
    layer0_outputs(1981) <= not((inputs(95)) xor (inputs(181)));
    layer0_outputs(1982) <= (inputs(107)) and not (inputs(77));
    layer0_outputs(1983) <= not((inputs(110)) or (inputs(33)));
    layer0_outputs(1984) <= inputs(193);
    layer0_outputs(1985) <= inputs(138);
    layer0_outputs(1986) <= not(inputs(75)) or (inputs(134));
    layer0_outputs(1987) <= inputs(212);
    layer0_outputs(1988) <= inputs(171);
    layer0_outputs(1989) <= (inputs(231)) or (inputs(21));
    layer0_outputs(1990) <= not((inputs(52)) and (inputs(42)));
    layer0_outputs(1991) <= inputs(91);
    layer0_outputs(1992) <= (inputs(21)) and not (inputs(26));
    layer0_outputs(1993) <= (inputs(27)) or (inputs(80));
    layer0_outputs(1994) <= (inputs(176)) and not (inputs(207));
    layer0_outputs(1995) <= (inputs(87)) and not (inputs(103));
    layer0_outputs(1996) <= not(inputs(230));
    layer0_outputs(1997) <= (inputs(85)) and not (inputs(207));
    layer0_outputs(1998) <= '1';
    layer0_outputs(1999) <= inputs(95);
    layer0_outputs(2000) <= '1';
    layer0_outputs(2001) <= '0';
    layer0_outputs(2002) <= inputs(89);
    layer0_outputs(2003) <= not(inputs(83));
    layer0_outputs(2004) <= inputs(45);
    layer0_outputs(2005) <= '1';
    layer0_outputs(2006) <= not(inputs(117));
    layer0_outputs(2007) <= not(inputs(165));
    layer0_outputs(2008) <= not(inputs(108)) or (inputs(184));
    layer0_outputs(2009) <= (inputs(27)) or (inputs(143));
    layer0_outputs(2010) <= not(inputs(22));
    layer0_outputs(2011) <= (inputs(229)) and not (inputs(154));
    layer0_outputs(2012) <= (inputs(4)) or (inputs(20));
    layer0_outputs(2013) <= inputs(120);
    layer0_outputs(2014) <= '1';
    layer0_outputs(2015) <= '0';
    layer0_outputs(2016) <= '0';
    layer0_outputs(2017) <= not(inputs(9));
    layer0_outputs(2018) <= inputs(32);
    layer0_outputs(2019) <= inputs(178);
    layer0_outputs(2020) <= '0';
    layer0_outputs(2021) <= not((inputs(187)) or (inputs(210)));
    layer0_outputs(2022) <= (inputs(170)) and not (inputs(2));
    layer0_outputs(2023) <= '1';
    layer0_outputs(2024) <= inputs(164);
    layer0_outputs(2025) <= not((inputs(255)) xor (inputs(234)));
    layer0_outputs(2026) <= not(inputs(109)) or (inputs(4));
    layer0_outputs(2027) <= '1';
    layer0_outputs(2028) <= (inputs(255)) or (inputs(149));
    layer0_outputs(2029) <= (inputs(91)) and not (inputs(85));
    layer0_outputs(2030) <= not(inputs(171));
    layer0_outputs(2031) <= not((inputs(194)) or (inputs(187)));
    layer0_outputs(2032) <= not((inputs(139)) or (inputs(46)));
    layer0_outputs(2033) <= '0';
    layer0_outputs(2034) <= (inputs(181)) and not (inputs(132));
    layer0_outputs(2035) <= inputs(12);
    layer0_outputs(2036) <= (inputs(112)) xor (inputs(86));
    layer0_outputs(2037) <= not(inputs(118)) or (inputs(206));
    layer0_outputs(2038) <= not(inputs(99));
    layer0_outputs(2039) <= not(inputs(225)) or (inputs(34));
    layer0_outputs(2040) <= not(inputs(77));
    layer0_outputs(2041) <= not(inputs(52)) or (inputs(59));
    layer0_outputs(2042) <= '0';
    layer0_outputs(2043) <= not(inputs(157));
    layer0_outputs(2044) <= not(inputs(31));
    layer0_outputs(2045) <= not(inputs(153)) or (inputs(212));
    layer0_outputs(2046) <= '1';
    layer0_outputs(2047) <= not(inputs(232)) or (inputs(224));
    layer0_outputs(2048) <= '0';
    layer0_outputs(2049) <= (inputs(130)) and (inputs(19));
    layer0_outputs(2050) <= not((inputs(131)) or (inputs(129)));
    layer0_outputs(2051) <= not((inputs(205)) or (inputs(179)));
    layer0_outputs(2052) <= (inputs(63)) and not (inputs(13));
    layer0_outputs(2053) <= not(inputs(94)) or (inputs(223));
    layer0_outputs(2054) <= not((inputs(4)) or (inputs(206)));
    layer0_outputs(2055) <= not(inputs(124)) or (inputs(226));
    layer0_outputs(2056) <= not(inputs(90)) or (inputs(86));
    layer0_outputs(2057) <= inputs(13);
    layer0_outputs(2058) <= (inputs(95)) and not (inputs(19));
    layer0_outputs(2059) <= '0';
    layer0_outputs(2060) <= '0';
    layer0_outputs(2061) <= '0';
    layer0_outputs(2062) <= '0';
    layer0_outputs(2063) <= (inputs(213)) and not (inputs(242));
    layer0_outputs(2064) <= not(inputs(153));
    layer0_outputs(2065) <= not((inputs(7)) or (inputs(170)));
    layer0_outputs(2066) <= (inputs(99)) and (inputs(6));
    layer0_outputs(2067) <= '1';
    layer0_outputs(2068) <= not(inputs(196));
    layer0_outputs(2069) <= not(inputs(228));
    layer0_outputs(2070) <= '0';
    layer0_outputs(2071) <= inputs(132);
    layer0_outputs(2072) <= inputs(146);
    layer0_outputs(2073) <= (inputs(240)) and not (inputs(6));
    layer0_outputs(2074) <= (inputs(239)) and (inputs(136));
    layer0_outputs(2075) <= not((inputs(177)) or (inputs(148)));
    layer0_outputs(2076) <= not((inputs(116)) xor (inputs(225)));
    layer0_outputs(2077) <= inputs(149);
    layer0_outputs(2078) <= not(inputs(59));
    layer0_outputs(2079) <= (inputs(121)) or (inputs(29));
    layer0_outputs(2080) <= (inputs(39)) and (inputs(142));
    layer0_outputs(2081) <= '1';
    layer0_outputs(2082) <= '0';
    layer0_outputs(2083) <= (inputs(15)) xor (inputs(78));
    layer0_outputs(2084) <= inputs(164);
    layer0_outputs(2085) <= (inputs(243)) and not (inputs(64));
    layer0_outputs(2086) <= '0';
    layer0_outputs(2087) <= (inputs(51)) and (inputs(201));
    layer0_outputs(2088) <= not(inputs(89)) or (inputs(197));
    layer0_outputs(2089) <= not((inputs(16)) xor (inputs(139)));
    layer0_outputs(2090) <= (inputs(80)) or (inputs(168));
    layer0_outputs(2091) <= (inputs(69)) xor (inputs(173));
    layer0_outputs(2092) <= not(inputs(121));
    layer0_outputs(2093) <= inputs(60);
    layer0_outputs(2094) <= not((inputs(5)) or (inputs(92)));
    layer0_outputs(2095) <= inputs(241);
    layer0_outputs(2096) <= not((inputs(178)) xor (inputs(239)));
    layer0_outputs(2097) <= not((inputs(141)) or (inputs(158)));
    layer0_outputs(2098) <= (inputs(244)) and not (inputs(183));
    layer0_outputs(2099) <= inputs(90);
    layer0_outputs(2100) <= '1';
    layer0_outputs(2101) <= not((inputs(206)) and (inputs(124)));
    layer0_outputs(2102) <= inputs(57);
    layer0_outputs(2103) <= not((inputs(20)) and (inputs(12)));
    layer0_outputs(2104) <= (inputs(160)) or (inputs(33));
    layer0_outputs(2105) <= not(inputs(15)) or (inputs(71));
    layer0_outputs(2106) <= '0';
    layer0_outputs(2107) <= '0';
    layer0_outputs(2108) <= inputs(98);
    layer0_outputs(2109) <= (inputs(173)) and (inputs(102));
    layer0_outputs(2110) <= not(inputs(154));
    layer0_outputs(2111) <= (inputs(179)) and not (inputs(249));
    layer0_outputs(2112) <= (inputs(197)) and not (inputs(26));
    layer0_outputs(2113) <= not((inputs(148)) and (inputs(164)));
    layer0_outputs(2114) <= not(inputs(162));
    layer0_outputs(2115) <= '1';
    layer0_outputs(2116) <= '0';
    layer0_outputs(2117) <= inputs(121);
    layer0_outputs(2118) <= (inputs(138)) and (inputs(65));
    layer0_outputs(2119) <= (inputs(15)) xor (inputs(89));
    layer0_outputs(2120) <= (inputs(199)) xor (inputs(241));
    layer0_outputs(2121) <= not(inputs(163));
    layer0_outputs(2122) <= (inputs(239)) or (inputs(15));
    layer0_outputs(2123) <= (inputs(180)) and (inputs(186));
    layer0_outputs(2124) <= '1';
    layer0_outputs(2125) <= '1';
    layer0_outputs(2126) <= not((inputs(32)) or (inputs(176)));
    layer0_outputs(2127) <= not((inputs(113)) or (inputs(53)));
    layer0_outputs(2128) <= not((inputs(66)) and (inputs(130)));
    layer0_outputs(2129) <= '1';
    layer0_outputs(2130) <= (inputs(115)) or (inputs(96));
    layer0_outputs(2131) <= inputs(150);
    layer0_outputs(2132) <= inputs(89);
    layer0_outputs(2133) <= '1';
    layer0_outputs(2134) <= (inputs(119)) and not (inputs(143));
    layer0_outputs(2135) <= '1';
    layer0_outputs(2136) <= (inputs(126)) or (inputs(53));
    layer0_outputs(2137) <= (inputs(170)) or (inputs(57));
    layer0_outputs(2138) <= inputs(52);
    layer0_outputs(2139) <= inputs(118);
    layer0_outputs(2140) <= (inputs(176)) and not (inputs(136));
    layer0_outputs(2141) <= (inputs(41)) and (inputs(249));
    layer0_outputs(2142) <= not(inputs(90)) or (inputs(191));
    layer0_outputs(2143) <= '0';
    layer0_outputs(2144) <= (inputs(5)) and (inputs(228));
    layer0_outputs(2145) <= (inputs(144)) and (inputs(22));
    layer0_outputs(2146) <= inputs(250);
    layer0_outputs(2147) <= '1';
    layer0_outputs(2148) <= not(inputs(195)) or (inputs(115));
    layer0_outputs(2149) <= not(inputs(145)) or (inputs(155));
    layer0_outputs(2150) <= not(inputs(179));
    layer0_outputs(2151) <= (inputs(170)) and (inputs(245));
    layer0_outputs(2152) <= '1';
    layer0_outputs(2153) <= '0';
    layer0_outputs(2154) <= not(inputs(119));
    layer0_outputs(2155) <= (inputs(199)) or (inputs(105));
    layer0_outputs(2156) <= not((inputs(119)) and (inputs(3)));
    layer0_outputs(2157) <= not((inputs(37)) and (inputs(147)));
    layer0_outputs(2158) <= (inputs(94)) and not (inputs(100));
    layer0_outputs(2159) <= inputs(202);
    layer0_outputs(2160) <= (inputs(223)) xor (inputs(112));
    layer0_outputs(2161) <= not(inputs(61));
    layer0_outputs(2162) <= not((inputs(77)) and (inputs(222)));
    layer0_outputs(2163) <= not(inputs(12));
    layer0_outputs(2164) <= '0';
    layer0_outputs(2165) <= inputs(232);
    layer0_outputs(2166) <= not((inputs(198)) and (inputs(40)));
    layer0_outputs(2167) <= not((inputs(30)) or (inputs(32)));
    layer0_outputs(2168) <= not((inputs(231)) and (inputs(102)));
    layer0_outputs(2169) <= (inputs(105)) and (inputs(142));
    layer0_outputs(2170) <= inputs(205);
    layer0_outputs(2171) <= not((inputs(239)) and (inputs(236)));
    layer0_outputs(2172) <= (inputs(36)) or (inputs(139));
    layer0_outputs(2173) <= inputs(173);
    layer0_outputs(2174) <= not(inputs(34)) or (inputs(210));
    layer0_outputs(2175) <= not((inputs(172)) xor (inputs(204)));
    layer0_outputs(2176) <= not(inputs(55)) or (inputs(174));
    layer0_outputs(2177) <= not(inputs(16));
    layer0_outputs(2178) <= not(inputs(167));
    layer0_outputs(2179) <= (inputs(140)) and not (inputs(192));
    layer0_outputs(2180) <= inputs(57);
    layer0_outputs(2181) <= '0';
    layer0_outputs(2182) <= (inputs(208)) and (inputs(95));
    layer0_outputs(2183) <= not(inputs(161));
    layer0_outputs(2184) <= not(inputs(4));
    layer0_outputs(2185) <= '0';
    layer0_outputs(2186) <= not(inputs(51));
    layer0_outputs(2187) <= not(inputs(232)) or (inputs(233));
    layer0_outputs(2188) <= '0';
    layer0_outputs(2189) <= not((inputs(115)) and (inputs(84)));
    layer0_outputs(2190) <= not(inputs(199)) or (inputs(220));
    layer0_outputs(2191) <= not((inputs(209)) xor (inputs(161)));
    layer0_outputs(2192) <= (inputs(58)) or (inputs(203));
    layer0_outputs(2193) <= not((inputs(79)) or (inputs(38)));
    layer0_outputs(2194) <= (inputs(120)) and not (inputs(112));
    layer0_outputs(2195) <= (inputs(141)) and not (inputs(176));
    layer0_outputs(2196) <= '1';
    layer0_outputs(2197) <= not(inputs(60)) or (inputs(143));
    layer0_outputs(2198) <= '0';
    layer0_outputs(2199) <= not(inputs(118));
    layer0_outputs(2200) <= '0';
    layer0_outputs(2201) <= '0';
    layer0_outputs(2202) <= not((inputs(151)) or (inputs(165)));
    layer0_outputs(2203) <= '1';
    layer0_outputs(2204) <= not((inputs(100)) and (inputs(227)));
    layer0_outputs(2205) <= '1';
    layer0_outputs(2206) <= (inputs(188)) or (inputs(145));
    layer0_outputs(2207) <= inputs(40);
    layer0_outputs(2208) <= inputs(178);
    layer0_outputs(2209) <= '0';
    layer0_outputs(2210) <= not(inputs(134)) or (inputs(5));
    layer0_outputs(2211) <= not(inputs(16));
    layer0_outputs(2212) <= (inputs(56)) and (inputs(110));
    layer0_outputs(2213) <= not(inputs(176));
    layer0_outputs(2214) <= not((inputs(65)) and (inputs(218)));
    layer0_outputs(2215) <= '1';
    layer0_outputs(2216) <= (inputs(181)) and not (inputs(123));
    layer0_outputs(2217) <= not((inputs(229)) or (inputs(2)));
    layer0_outputs(2218) <= not((inputs(203)) or (inputs(220)));
    layer0_outputs(2219) <= inputs(130);
    layer0_outputs(2220) <= inputs(89);
    layer0_outputs(2221) <= inputs(219);
    layer0_outputs(2222) <= inputs(121);
    layer0_outputs(2223) <= (inputs(184)) and not (inputs(33));
    layer0_outputs(2224) <= not((inputs(107)) and (inputs(109)));
    layer0_outputs(2225) <= (inputs(48)) and not (inputs(231));
    layer0_outputs(2226) <= inputs(177);
    layer0_outputs(2227) <= inputs(250);
    layer0_outputs(2228) <= not(inputs(131));
    layer0_outputs(2229) <= not((inputs(157)) xor (inputs(234)));
    layer0_outputs(2230) <= (inputs(188)) and not (inputs(43));
    layer0_outputs(2231) <= not(inputs(103));
    layer0_outputs(2232) <= (inputs(239)) and not (inputs(225));
    layer0_outputs(2233) <= not(inputs(102));
    layer0_outputs(2234) <= not(inputs(172));
    layer0_outputs(2235) <= not(inputs(50));
    layer0_outputs(2236) <= not((inputs(247)) or (inputs(92)));
    layer0_outputs(2237) <= inputs(120);
    layer0_outputs(2238) <= '1';
    layer0_outputs(2239) <= '0';
    layer0_outputs(2240) <= inputs(67);
    layer0_outputs(2241) <= (inputs(254)) xor (inputs(86));
    layer0_outputs(2242) <= not(inputs(151)) or (inputs(140));
    layer0_outputs(2243) <= not(inputs(97));
    layer0_outputs(2244) <= not(inputs(82));
    layer0_outputs(2245) <= inputs(161);
    layer0_outputs(2246) <= '1';
    layer0_outputs(2247) <= not((inputs(170)) or (inputs(84)));
    layer0_outputs(2248) <= (inputs(216)) and not (inputs(49));
    layer0_outputs(2249) <= '0';
    layer0_outputs(2250) <= inputs(238);
    layer0_outputs(2251) <= (inputs(219)) or (inputs(154));
    layer0_outputs(2252) <= (inputs(76)) xor (inputs(204));
    layer0_outputs(2253) <= not((inputs(122)) or (inputs(138)));
    layer0_outputs(2254) <= '0';
    layer0_outputs(2255) <= not(inputs(29));
    layer0_outputs(2256) <= inputs(177);
    layer0_outputs(2257) <= not(inputs(31)) or (inputs(91));
    layer0_outputs(2258) <= not(inputs(169));
    layer0_outputs(2259) <= not((inputs(125)) and (inputs(152)));
    layer0_outputs(2260) <= (inputs(0)) or (inputs(143));
    layer0_outputs(2261) <= (inputs(56)) or (inputs(46));
    layer0_outputs(2262) <= '1';
    layer0_outputs(2263) <= not(inputs(205)) or (inputs(31));
    layer0_outputs(2264) <= (inputs(82)) or (inputs(147));
    layer0_outputs(2265) <= (inputs(115)) or (inputs(104));
    layer0_outputs(2266) <= not(inputs(117));
    layer0_outputs(2267) <= (inputs(190)) or (inputs(204));
    layer0_outputs(2268) <= not(inputs(198)) or (inputs(143));
    layer0_outputs(2269) <= not(inputs(166));
    layer0_outputs(2270) <= not((inputs(131)) xor (inputs(195)));
    layer0_outputs(2271) <= not(inputs(245)) or (inputs(114));
    layer0_outputs(2272) <= inputs(248);
    layer0_outputs(2273) <= (inputs(37)) or (inputs(126));
    layer0_outputs(2274) <= not(inputs(10)) or (inputs(157));
    layer0_outputs(2275) <= (inputs(80)) and not (inputs(215));
    layer0_outputs(2276) <= not(inputs(7)) or (inputs(108));
    layer0_outputs(2277) <= not((inputs(182)) or (inputs(185)));
    layer0_outputs(2278) <= not((inputs(22)) and (inputs(29)));
    layer0_outputs(2279) <= (inputs(243)) or (inputs(40));
    layer0_outputs(2280) <= not(inputs(205)) or (inputs(55));
    layer0_outputs(2281) <= inputs(230);
    layer0_outputs(2282) <= (inputs(150)) or (inputs(123));
    layer0_outputs(2283) <= not((inputs(178)) or (inputs(173)));
    layer0_outputs(2284) <= not((inputs(48)) or (inputs(250)));
    layer0_outputs(2285) <= not(inputs(207)) or (inputs(43));
    layer0_outputs(2286) <= not(inputs(164)) or (inputs(181));
    layer0_outputs(2287) <= (inputs(251)) xor (inputs(47));
    layer0_outputs(2288) <= '0';
    layer0_outputs(2289) <= '0';
    layer0_outputs(2290) <= '1';
    layer0_outputs(2291) <= '1';
    layer0_outputs(2292) <= not(inputs(210));
    layer0_outputs(2293) <= (inputs(143)) and not (inputs(35));
    layer0_outputs(2294) <= (inputs(42)) and not (inputs(184));
    layer0_outputs(2295) <= '0';
    layer0_outputs(2296) <= '1';
    layer0_outputs(2297) <= not(inputs(43));
    layer0_outputs(2298) <= '0';
    layer0_outputs(2299) <= inputs(182);
    layer0_outputs(2300) <= not(inputs(180));
    layer0_outputs(2301) <= (inputs(114)) and (inputs(195));
    layer0_outputs(2302) <= not((inputs(122)) or (inputs(2)));
    layer0_outputs(2303) <= (inputs(220)) or (inputs(14));
    layer0_outputs(2304) <= (inputs(250)) or (inputs(67));
    layer0_outputs(2305) <= (inputs(85)) and not (inputs(81));
    layer0_outputs(2306) <= (inputs(8)) and not (inputs(182));
    layer0_outputs(2307) <= (inputs(146)) or (inputs(161));
    layer0_outputs(2308) <= (inputs(190)) and not (inputs(63));
    layer0_outputs(2309) <= (inputs(1)) and not (inputs(110));
    layer0_outputs(2310) <= inputs(75);
    layer0_outputs(2311) <= not((inputs(210)) or (inputs(87)));
    layer0_outputs(2312) <= inputs(106);
    layer0_outputs(2313) <= (inputs(68)) or (inputs(53));
    layer0_outputs(2314) <= not(inputs(42)) or (inputs(76));
    layer0_outputs(2315) <= not(inputs(119)) or (inputs(47));
    layer0_outputs(2316) <= (inputs(48)) or (inputs(189));
    layer0_outputs(2317) <= inputs(90);
    layer0_outputs(2318) <= not(inputs(127)) or (inputs(92));
    layer0_outputs(2319) <= (inputs(244)) and not (inputs(162));
    layer0_outputs(2320) <= inputs(88);
    layer0_outputs(2321) <= inputs(92);
    layer0_outputs(2322) <= not(inputs(37));
    layer0_outputs(2323) <= '1';
    layer0_outputs(2324) <= not((inputs(33)) or (inputs(63)));
    layer0_outputs(2325) <= inputs(216);
    layer0_outputs(2326) <= not((inputs(152)) and (inputs(234)));
    layer0_outputs(2327) <= not(inputs(210)) or (inputs(65));
    layer0_outputs(2328) <= not(inputs(120));
    layer0_outputs(2329) <= not((inputs(66)) or (inputs(101)));
    layer0_outputs(2330) <= '0';
    layer0_outputs(2331) <= inputs(123);
    layer0_outputs(2332) <= not(inputs(127));
    layer0_outputs(2333) <= inputs(103);
    layer0_outputs(2334) <= (inputs(32)) and (inputs(238));
    layer0_outputs(2335) <= (inputs(156)) xor (inputs(181));
    layer0_outputs(2336) <= '1';
    layer0_outputs(2337) <= not(inputs(44));
    layer0_outputs(2338) <= inputs(164);
    layer0_outputs(2339) <= not((inputs(54)) and (inputs(96)));
    layer0_outputs(2340) <= inputs(154);
    layer0_outputs(2341) <= '0';
    layer0_outputs(2342) <= not((inputs(7)) or (inputs(132)));
    layer0_outputs(2343) <= (inputs(66)) and (inputs(153));
    layer0_outputs(2344) <= not((inputs(172)) or (inputs(132)));
    layer0_outputs(2345) <= (inputs(19)) and not (inputs(239));
    layer0_outputs(2346) <= '0';
    layer0_outputs(2347) <= not(inputs(226));
    layer0_outputs(2348) <= not(inputs(227)) or (inputs(144));
    layer0_outputs(2349) <= not((inputs(208)) and (inputs(49)));
    layer0_outputs(2350) <= inputs(140);
    layer0_outputs(2351) <= not(inputs(60)) or (inputs(236));
    layer0_outputs(2352) <= '0';
    layer0_outputs(2353) <= not(inputs(212));
    layer0_outputs(2354) <= (inputs(74)) xor (inputs(12));
    layer0_outputs(2355) <= not(inputs(9));
    layer0_outputs(2356) <= not((inputs(92)) or (inputs(130)));
    layer0_outputs(2357) <= (inputs(123)) and not (inputs(28));
    layer0_outputs(2358) <= not((inputs(151)) or (inputs(137)));
    layer0_outputs(2359) <= '0';
    layer0_outputs(2360) <= (inputs(45)) or (inputs(126));
    layer0_outputs(2361) <= not(inputs(195));
    layer0_outputs(2362) <= (inputs(224)) and (inputs(110));
    layer0_outputs(2363) <= not(inputs(106)) or (inputs(226));
    layer0_outputs(2364) <= not((inputs(174)) and (inputs(195)));
    layer0_outputs(2365) <= '1';
    layer0_outputs(2366) <= not(inputs(93));
    layer0_outputs(2367) <= not((inputs(146)) and (inputs(217)));
    layer0_outputs(2368) <= '1';
    layer0_outputs(2369) <= not(inputs(249)) or (inputs(44));
    layer0_outputs(2370) <= '0';
    layer0_outputs(2371) <= (inputs(70)) or (inputs(94));
    layer0_outputs(2372) <= (inputs(150)) or (inputs(49));
    layer0_outputs(2373) <= not(inputs(97)) or (inputs(79));
    layer0_outputs(2374) <= (inputs(146)) xor (inputs(208));
    layer0_outputs(2375) <= (inputs(95)) and not (inputs(255));
    layer0_outputs(2376) <= not(inputs(252)) or (inputs(51));
    layer0_outputs(2377) <= (inputs(86)) or (inputs(105));
    layer0_outputs(2378) <= inputs(112);
    layer0_outputs(2379) <= not((inputs(239)) and (inputs(13)));
    layer0_outputs(2380) <= not((inputs(231)) and (inputs(179)));
    layer0_outputs(2381) <= inputs(30);
    layer0_outputs(2382) <= not(inputs(84)) or (inputs(194));
    layer0_outputs(2383) <= '0';
    layer0_outputs(2384) <= '1';
    layer0_outputs(2385) <= (inputs(18)) or (inputs(102));
    layer0_outputs(2386) <= inputs(55);
    layer0_outputs(2387) <= (inputs(153)) and not (inputs(32));
    layer0_outputs(2388) <= inputs(79);
    layer0_outputs(2389) <= not(inputs(128));
    layer0_outputs(2390) <= (inputs(66)) or (inputs(191));
    layer0_outputs(2391) <= '0';
    layer0_outputs(2392) <= not(inputs(194));
    layer0_outputs(2393) <= '0';
    layer0_outputs(2394) <= '0';
    layer0_outputs(2395) <= not(inputs(58));
    layer0_outputs(2396) <= (inputs(63)) or (inputs(219));
    layer0_outputs(2397) <= (inputs(147)) and not (inputs(73));
    layer0_outputs(2398) <= (inputs(127)) xor (inputs(106));
    layer0_outputs(2399) <= not((inputs(132)) or (inputs(87)));
    layer0_outputs(2400) <= not(inputs(196));
    layer0_outputs(2401) <= not(inputs(139));
    layer0_outputs(2402) <= (inputs(254)) and not (inputs(239));
    layer0_outputs(2403) <= inputs(215);
    layer0_outputs(2404) <= inputs(233);
    layer0_outputs(2405) <= inputs(39);
    layer0_outputs(2406) <= '1';
    layer0_outputs(2407) <= inputs(136);
    layer0_outputs(2408) <= not((inputs(92)) or (inputs(40)));
    layer0_outputs(2409) <= '0';
    layer0_outputs(2410) <= not(inputs(1)) or (inputs(83));
    layer0_outputs(2411) <= inputs(245);
    layer0_outputs(2412) <= not(inputs(83));
    layer0_outputs(2413) <= inputs(146);
    layer0_outputs(2414) <= not((inputs(165)) xor (inputs(243)));
    layer0_outputs(2415) <= not((inputs(114)) and (inputs(187)));
    layer0_outputs(2416) <= not(inputs(129));
    layer0_outputs(2417) <= '0';
    layer0_outputs(2418) <= '1';
    layer0_outputs(2419) <= (inputs(214)) and (inputs(156));
    layer0_outputs(2420) <= inputs(124);
    layer0_outputs(2421) <= (inputs(76)) or (inputs(50));
    layer0_outputs(2422) <= not(inputs(93)) or (inputs(130));
    layer0_outputs(2423) <= not(inputs(221));
    layer0_outputs(2424) <= (inputs(27)) and not (inputs(174));
    layer0_outputs(2425) <= '0';
    layer0_outputs(2426) <= '0';
    layer0_outputs(2427) <= not(inputs(195));
    layer0_outputs(2428) <= inputs(80);
    layer0_outputs(2429) <= inputs(176);
    layer0_outputs(2430) <= (inputs(105)) and not (inputs(170));
    layer0_outputs(2431) <= not(inputs(94));
    layer0_outputs(2432) <= not(inputs(9));
    layer0_outputs(2433) <= not(inputs(178)) or (inputs(111));
    layer0_outputs(2434) <= inputs(252);
    layer0_outputs(2435) <= not((inputs(15)) and (inputs(22)));
    layer0_outputs(2436) <= '1';
    layer0_outputs(2437) <= (inputs(254)) or (inputs(206));
    layer0_outputs(2438) <= not((inputs(198)) or (inputs(195)));
    layer0_outputs(2439) <= (inputs(197)) or (inputs(232));
    layer0_outputs(2440) <= '0';
    layer0_outputs(2441) <= (inputs(139)) and not (inputs(19));
    layer0_outputs(2442) <= not(inputs(222));
    layer0_outputs(2443) <= (inputs(144)) or (inputs(131));
    layer0_outputs(2444) <= inputs(108);
    layer0_outputs(2445) <= (inputs(85)) or (inputs(245));
    layer0_outputs(2446) <= not(inputs(251)) or (inputs(78));
    layer0_outputs(2447) <= not(inputs(128));
    layer0_outputs(2448) <= not((inputs(14)) xor (inputs(52)));
    layer0_outputs(2449) <= (inputs(201)) or (inputs(62));
    layer0_outputs(2450) <= not((inputs(95)) and (inputs(43)));
    layer0_outputs(2451) <= '1';
    layer0_outputs(2452) <= (inputs(52)) and not (inputs(171));
    layer0_outputs(2453) <= inputs(230);
    layer0_outputs(2454) <= not((inputs(149)) or (inputs(69)));
    layer0_outputs(2455) <= (inputs(254)) xor (inputs(241));
    layer0_outputs(2456) <= not(inputs(204)) or (inputs(138));
    layer0_outputs(2457) <= '0';
    layer0_outputs(2458) <= inputs(195);
    layer0_outputs(2459) <= inputs(87);
    layer0_outputs(2460) <= (inputs(222)) and not (inputs(0));
    layer0_outputs(2461) <= not((inputs(176)) and (inputs(36)));
    layer0_outputs(2462) <= not(inputs(204)) or (inputs(202));
    layer0_outputs(2463) <= not(inputs(68));
    layer0_outputs(2464) <= (inputs(73)) and (inputs(171));
    layer0_outputs(2465) <= inputs(122);
    layer0_outputs(2466) <= inputs(80);
    layer0_outputs(2467) <= '0';
    layer0_outputs(2468) <= '1';
    layer0_outputs(2469) <= not(inputs(255)) or (inputs(124));
    layer0_outputs(2470) <= not(inputs(185));
    layer0_outputs(2471) <= '1';
    layer0_outputs(2472) <= '0';
    layer0_outputs(2473) <= not(inputs(145)) or (inputs(161));
    layer0_outputs(2474) <= not((inputs(17)) and (inputs(158)));
    layer0_outputs(2475) <= not((inputs(132)) xor (inputs(162)));
    layer0_outputs(2476) <= not(inputs(142));
    layer0_outputs(2477) <= (inputs(18)) or (inputs(126));
    layer0_outputs(2478) <= (inputs(5)) or (inputs(171));
    layer0_outputs(2479) <= not(inputs(131));
    layer0_outputs(2480) <= not(inputs(143));
    layer0_outputs(2481) <= not((inputs(225)) or (inputs(232)));
    layer0_outputs(2482) <= not(inputs(229));
    layer0_outputs(2483) <= not(inputs(50)) or (inputs(71));
    layer0_outputs(2484) <= (inputs(108)) or (inputs(103));
    layer0_outputs(2485) <= not(inputs(32)) or (inputs(235));
    layer0_outputs(2486) <= (inputs(253)) and not (inputs(248));
    layer0_outputs(2487) <= inputs(247);
    layer0_outputs(2488) <= '1';
    layer0_outputs(2489) <= (inputs(110)) or (inputs(181));
    layer0_outputs(2490) <= (inputs(33)) xor (inputs(30));
    layer0_outputs(2491) <= not(inputs(198));
    layer0_outputs(2492) <= inputs(148);
    layer0_outputs(2493) <= not((inputs(129)) or (inputs(205)));
    layer0_outputs(2494) <= (inputs(164)) and not (inputs(226));
    layer0_outputs(2495) <= inputs(135);
    layer0_outputs(2496) <= (inputs(227)) or (inputs(91));
    layer0_outputs(2497) <= (inputs(97)) and not (inputs(102));
    layer0_outputs(2498) <= '1';
    layer0_outputs(2499) <= inputs(189);
    layer0_outputs(2500) <= not(inputs(242)) or (inputs(211));
    layer0_outputs(2501) <= '1';
    layer0_outputs(2502) <= not(inputs(129));
    layer0_outputs(2503) <= not((inputs(17)) or (inputs(221)));
    layer0_outputs(2504) <= (inputs(189)) and not (inputs(204));
    layer0_outputs(2505) <= '1';
    layer0_outputs(2506) <= (inputs(12)) and not (inputs(146));
    layer0_outputs(2507) <= not((inputs(117)) xor (inputs(66)));
    layer0_outputs(2508) <= not(inputs(182));
    layer0_outputs(2509) <= not(inputs(45)) or (inputs(161));
    layer0_outputs(2510) <= not((inputs(218)) or (inputs(189)));
    layer0_outputs(2511) <= (inputs(82)) and not (inputs(91));
    layer0_outputs(2512) <= not(inputs(187));
    layer0_outputs(2513) <= not(inputs(238));
    layer0_outputs(2514) <= inputs(100);
    layer0_outputs(2515) <= not(inputs(68));
    layer0_outputs(2516) <= not((inputs(140)) xor (inputs(219)));
    layer0_outputs(2517) <= not(inputs(244));
    layer0_outputs(2518) <= not(inputs(135)) or (inputs(187));
    layer0_outputs(2519) <= (inputs(229)) and not (inputs(158));
    layer0_outputs(2520) <= inputs(204);
    layer0_outputs(2521) <= not(inputs(168));
    layer0_outputs(2522) <= not(inputs(192));
    layer0_outputs(2523) <= '0';
    layer0_outputs(2524) <= not((inputs(116)) or (inputs(99)));
    layer0_outputs(2525) <= not(inputs(113));
    layer0_outputs(2526) <= (inputs(253)) and not (inputs(140));
    layer0_outputs(2527) <= not((inputs(197)) or (inputs(182)));
    layer0_outputs(2528) <= '1';
    layer0_outputs(2529) <= (inputs(179)) and not (inputs(212));
    layer0_outputs(2530) <= (inputs(225)) or (inputs(199));
    layer0_outputs(2531) <= not(inputs(172)) or (inputs(159));
    layer0_outputs(2532) <= '0';
    layer0_outputs(2533) <= not((inputs(62)) and (inputs(142)));
    layer0_outputs(2534) <= inputs(231);
    layer0_outputs(2535) <= (inputs(143)) and not (inputs(43));
    layer0_outputs(2536) <= inputs(226);
    layer0_outputs(2537) <= not((inputs(119)) or (inputs(4)));
    layer0_outputs(2538) <= not(inputs(114));
    layer0_outputs(2539) <= (inputs(19)) and (inputs(53));
    layer0_outputs(2540) <= (inputs(174)) or (inputs(204));
    layer0_outputs(2541) <= not(inputs(212));
    layer0_outputs(2542) <= (inputs(132)) and not (inputs(240));
    layer0_outputs(2543) <= '1';
    layer0_outputs(2544) <= '1';
    layer0_outputs(2545) <= inputs(116);
    layer0_outputs(2546) <= '1';
    layer0_outputs(2547) <= '0';
    layer0_outputs(2548) <= not((inputs(173)) and (inputs(250)));
    layer0_outputs(2549) <= inputs(211);
    layer0_outputs(2550) <= (inputs(32)) and not (inputs(178));
    layer0_outputs(2551) <= inputs(171);
    layer0_outputs(2552) <= not((inputs(111)) or (inputs(175)));
    layer0_outputs(2553) <= not(inputs(197));
    layer0_outputs(2554) <= (inputs(112)) and not (inputs(2));
    layer0_outputs(2555) <= (inputs(157)) and not (inputs(31));
    layer0_outputs(2556) <= (inputs(66)) and not (inputs(52));
    layer0_outputs(2557) <= '1';
    layer0_outputs(2558) <= (inputs(20)) or (inputs(84));
    layer0_outputs(2559) <= '0';
    layer0_outputs(2560) <= (inputs(84)) and not (inputs(71));
    layer0_outputs(2561) <= not((inputs(35)) or (inputs(230)));
    layer0_outputs(2562) <= (inputs(83)) and not (inputs(15));
    layer0_outputs(2563) <= not(inputs(178));
    layer0_outputs(2564) <= (inputs(69)) and not (inputs(85));
    layer0_outputs(2565) <= '1';
    layer0_outputs(2566) <= inputs(222);
    layer0_outputs(2567) <= not(inputs(131)) or (inputs(253));
    layer0_outputs(2568) <= not(inputs(227));
    layer0_outputs(2569) <= not(inputs(97));
    layer0_outputs(2570) <= (inputs(17)) and (inputs(49));
    layer0_outputs(2571) <= (inputs(0)) and (inputs(144));
    layer0_outputs(2572) <= '0';
    layer0_outputs(2573) <= not(inputs(186)) or (inputs(161));
    layer0_outputs(2574) <= not((inputs(181)) and (inputs(169)));
    layer0_outputs(2575) <= '0';
    layer0_outputs(2576) <= inputs(207);
    layer0_outputs(2577) <= not((inputs(176)) and (inputs(86)));
    layer0_outputs(2578) <= not(inputs(172));
    layer0_outputs(2579) <= not(inputs(197));
    layer0_outputs(2580) <= (inputs(183)) xor (inputs(156));
    layer0_outputs(2581) <= '0';
    layer0_outputs(2582) <= '0';
    layer0_outputs(2583) <= (inputs(155)) or (inputs(124));
    layer0_outputs(2584) <= not(inputs(131)) or (inputs(251));
    layer0_outputs(2585) <= inputs(63);
    layer0_outputs(2586) <= not(inputs(140));
    layer0_outputs(2587) <= (inputs(162)) or (inputs(172));
    layer0_outputs(2588) <= not(inputs(72));
    layer0_outputs(2589) <= (inputs(22)) and (inputs(214));
    layer0_outputs(2590) <= '0';
    layer0_outputs(2591) <= not(inputs(255));
    layer0_outputs(2592) <= not((inputs(19)) and (inputs(118)));
    layer0_outputs(2593) <= '0';
    layer0_outputs(2594) <= not((inputs(50)) and (inputs(27)));
    layer0_outputs(2595) <= not(inputs(236)) or (inputs(78));
    layer0_outputs(2596) <= inputs(229);
    layer0_outputs(2597) <= not(inputs(44));
    layer0_outputs(2598) <= '1';
    layer0_outputs(2599) <= not((inputs(92)) and (inputs(8)));
    layer0_outputs(2600) <= (inputs(247)) and not (inputs(86));
    layer0_outputs(2601) <= not(inputs(198)) or (inputs(62));
    layer0_outputs(2602) <= not(inputs(177));
    layer0_outputs(2603) <= '0';
    layer0_outputs(2604) <= '0';
    layer0_outputs(2605) <= '0';
    layer0_outputs(2606) <= (inputs(94)) or (inputs(192));
    layer0_outputs(2607) <= not((inputs(248)) or (inputs(68)));
    layer0_outputs(2608) <= (inputs(249)) and (inputs(242));
    layer0_outputs(2609) <= (inputs(40)) or (inputs(121));
    layer0_outputs(2610) <= (inputs(54)) and not (inputs(217));
    layer0_outputs(2611) <= not(inputs(230)) or (inputs(16));
    layer0_outputs(2612) <= '1';
    layer0_outputs(2613) <= '0';
    layer0_outputs(2614) <= not((inputs(23)) or (inputs(108)));
    layer0_outputs(2615) <= not((inputs(43)) or (inputs(95)));
    layer0_outputs(2616) <= '1';
    layer0_outputs(2617) <= not(inputs(222));
    layer0_outputs(2618) <= '0';
    layer0_outputs(2619) <= (inputs(91)) or (inputs(73));
    layer0_outputs(2620) <= (inputs(198)) and not (inputs(85));
    layer0_outputs(2621) <= not(inputs(81));
    layer0_outputs(2622) <= not(inputs(113));
    layer0_outputs(2623) <= (inputs(52)) and not (inputs(88));
    layer0_outputs(2624) <= not(inputs(181)) or (inputs(113));
    layer0_outputs(2625) <= not((inputs(139)) or (inputs(103)));
    layer0_outputs(2626) <= (inputs(34)) xor (inputs(173));
    layer0_outputs(2627) <= (inputs(252)) and not (inputs(128));
    layer0_outputs(2628) <= not(inputs(67));
    layer0_outputs(2629) <= not(inputs(6));
    layer0_outputs(2630) <= (inputs(57)) and not (inputs(7));
    layer0_outputs(2631) <= not((inputs(61)) or (inputs(182)));
    layer0_outputs(2632) <= '0';
    layer0_outputs(2633) <= (inputs(145)) and (inputs(232));
    layer0_outputs(2634) <= not(inputs(167)) or (inputs(81));
    layer0_outputs(2635) <= not((inputs(255)) or (inputs(110)));
    layer0_outputs(2636) <= not((inputs(38)) or (inputs(116)));
    layer0_outputs(2637) <= (inputs(125)) xor (inputs(125));
    layer0_outputs(2638) <= not(inputs(132)) or (inputs(224));
    layer0_outputs(2639) <= inputs(142);
    layer0_outputs(2640) <= not(inputs(243)) or (inputs(143));
    layer0_outputs(2641) <= not((inputs(180)) or (inputs(253)));
    layer0_outputs(2642) <= inputs(122);
    layer0_outputs(2643) <= '1';
    layer0_outputs(2644) <= (inputs(230)) or (inputs(179));
    layer0_outputs(2645) <= not(inputs(208));
    layer0_outputs(2646) <= (inputs(107)) and (inputs(107));
    layer0_outputs(2647) <= (inputs(46)) or (inputs(195));
    layer0_outputs(2648) <= '1';
    layer0_outputs(2649) <= not((inputs(124)) or (inputs(101)));
    layer0_outputs(2650) <= not(inputs(160)) or (inputs(213));
    layer0_outputs(2651) <= not(inputs(121)) or (inputs(12));
    layer0_outputs(2652) <= '1';
    layer0_outputs(2653) <= '1';
    layer0_outputs(2654) <= (inputs(203)) and not (inputs(154));
    layer0_outputs(2655) <= '1';
    layer0_outputs(2656) <= not(inputs(118));
    layer0_outputs(2657) <= '0';
    layer0_outputs(2658) <= inputs(67);
    layer0_outputs(2659) <= not((inputs(250)) or (inputs(145)));
    layer0_outputs(2660) <= (inputs(48)) or (inputs(209));
    layer0_outputs(2661) <= (inputs(68)) or (inputs(53));
    layer0_outputs(2662) <= inputs(98);
    layer0_outputs(2663) <= (inputs(221)) and not (inputs(60));
    layer0_outputs(2664) <= not((inputs(62)) xor (inputs(123)));
    layer0_outputs(2665) <= (inputs(92)) xor (inputs(18));
    layer0_outputs(2666) <= (inputs(34)) or (inputs(216));
    layer0_outputs(2667) <= not(inputs(183));
    layer0_outputs(2668) <= '1';
    layer0_outputs(2669) <= '0';
    layer0_outputs(2670) <= (inputs(187)) or (inputs(204));
    layer0_outputs(2671) <= inputs(222);
    layer0_outputs(2672) <= inputs(60);
    layer0_outputs(2673) <= not((inputs(49)) or (inputs(237)));
    layer0_outputs(2674) <= not(inputs(101));
    layer0_outputs(2675) <= inputs(125);
    layer0_outputs(2676) <= not(inputs(221));
    layer0_outputs(2677) <= (inputs(167)) and not (inputs(233));
    layer0_outputs(2678) <= '1';
    layer0_outputs(2679) <= (inputs(100)) or (inputs(4));
    layer0_outputs(2680) <= '1';
    layer0_outputs(2681) <= inputs(198);
    layer0_outputs(2682) <= not(inputs(240));
    layer0_outputs(2683) <= '0';
    layer0_outputs(2684) <= not(inputs(13));
    layer0_outputs(2685) <= not(inputs(101)) or (inputs(212));
    layer0_outputs(2686) <= not((inputs(135)) or (inputs(206)));
    layer0_outputs(2687) <= '1';
    layer0_outputs(2688) <= '0';
    layer0_outputs(2689) <= inputs(150);
    layer0_outputs(2690) <= (inputs(127)) or (inputs(79));
    layer0_outputs(2691) <= not((inputs(162)) and (inputs(104)));
    layer0_outputs(2692) <= not((inputs(77)) or (inputs(75)));
    layer0_outputs(2693) <= (inputs(46)) and not (inputs(210));
    layer0_outputs(2694) <= not(inputs(203));
    layer0_outputs(2695) <= (inputs(159)) or (inputs(63));
    layer0_outputs(2696) <= not(inputs(162));
    layer0_outputs(2697) <= (inputs(73)) and (inputs(34));
    layer0_outputs(2698) <= not(inputs(135)) or (inputs(156));
    layer0_outputs(2699) <= (inputs(162)) and (inputs(30));
    layer0_outputs(2700) <= (inputs(209)) xor (inputs(149));
    layer0_outputs(2701) <= '0';
    layer0_outputs(2702) <= not((inputs(171)) and (inputs(128)));
    layer0_outputs(2703) <= not(inputs(130));
    layer0_outputs(2704) <= inputs(43);
    layer0_outputs(2705) <= not(inputs(151)) or (inputs(190));
    layer0_outputs(2706) <= '1';
    layer0_outputs(2707) <= (inputs(105)) or (inputs(254));
    layer0_outputs(2708) <= not(inputs(23));
    layer0_outputs(2709) <= (inputs(41)) and (inputs(139));
    layer0_outputs(2710) <= (inputs(53)) xor (inputs(222));
    layer0_outputs(2711) <= not(inputs(75)) or (inputs(157));
    layer0_outputs(2712) <= '1';
    layer0_outputs(2713) <= not(inputs(16));
    layer0_outputs(2714) <= (inputs(190)) and not (inputs(210));
    layer0_outputs(2715) <= inputs(234);
    layer0_outputs(2716) <= not(inputs(181)) or (inputs(47));
    layer0_outputs(2717) <= not(inputs(42));
    layer0_outputs(2718) <= inputs(121);
    layer0_outputs(2719) <= not(inputs(178));
    layer0_outputs(2720) <= not(inputs(223));
    layer0_outputs(2721) <= (inputs(177)) or (inputs(196));
    layer0_outputs(2722) <= not((inputs(221)) or (inputs(210)));
    layer0_outputs(2723) <= inputs(220);
    layer0_outputs(2724) <= (inputs(208)) and not (inputs(160));
    layer0_outputs(2725) <= not(inputs(26));
    layer0_outputs(2726) <= '1';
    layer0_outputs(2727) <= (inputs(224)) or (inputs(56));
    layer0_outputs(2728) <= not(inputs(12));
    layer0_outputs(2729) <= not(inputs(83));
    layer0_outputs(2730) <= '0';
    layer0_outputs(2731) <= not((inputs(119)) and (inputs(24)));
    layer0_outputs(2732) <= (inputs(176)) or (inputs(217));
    layer0_outputs(2733) <= inputs(190);
    layer0_outputs(2734) <= (inputs(25)) and not (inputs(153));
    layer0_outputs(2735) <= (inputs(160)) and (inputs(180));
    layer0_outputs(2736) <= not((inputs(77)) xor (inputs(51)));
    layer0_outputs(2737) <= not(inputs(168)) or (inputs(218));
    layer0_outputs(2738) <= '1';
    layer0_outputs(2739) <= '1';
    layer0_outputs(2740) <= (inputs(173)) and not (inputs(14));
    layer0_outputs(2741) <= not((inputs(98)) and (inputs(99)));
    layer0_outputs(2742) <= not(inputs(121));
    layer0_outputs(2743) <= not(inputs(230));
    layer0_outputs(2744) <= (inputs(161)) and not (inputs(65));
    layer0_outputs(2745) <= (inputs(223)) and (inputs(71));
    layer0_outputs(2746) <= not((inputs(254)) or (inputs(133)));
    layer0_outputs(2747) <= (inputs(19)) and not (inputs(94));
    layer0_outputs(2748) <= not(inputs(96));
    layer0_outputs(2749) <= (inputs(170)) and not (inputs(83));
    layer0_outputs(2750) <= not(inputs(181));
    layer0_outputs(2751) <= not(inputs(116)) or (inputs(49));
    layer0_outputs(2752) <= '0';
    layer0_outputs(2753) <= '0';
    layer0_outputs(2754) <= '0';
    layer0_outputs(2755) <= not(inputs(81));
    layer0_outputs(2756) <= not(inputs(238));
    layer0_outputs(2757) <= '0';
    layer0_outputs(2758) <= not(inputs(232));
    layer0_outputs(2759) <= inputs(126);
    layer0_outputs(2760) <= not(inputs(211));
    layer0_outputs(2761) <= '0';
    layer0_outputs(2762) <= not(inputs(76)) or (inputs(117));
    layer0_outputs(2763) <= '1';
    layer0_outputs(2764) <= not(inputs(47));
    layer0_outputs(2765) <= '1';
    layer0_outputs(2766) <= '0';
    layer0_outputs(2767) <= not((inputs(28)) and (inputs(173)));
    layer0_outputs(2768) <= not(inputs(189));
    layer0_outputs(2769) <= not(inputs(244)) or (inputs(128));
    layer0_outputs(2770) <= not((inputs(29)) and (inputs(79)));
    layer0_outputs(2771) <= not((inputs(166)) or (inputs(29)));
    layer0_outputs(2772) <= not(inputs(177));
    layer0_outputs(2773) <= inputs(128);
    layer0_outputs(2774) <= not(inputs(6)) or (inputs(96));
    layer0_outputs(2775) <= (inputs(190)) and not (inputs(72));
    layer0_outputs(2776) <= not(inputs(200)) or (inputs(152));
    layer0_outputs(2777) <= not(inputs(175)) or (inputs(87));
    layer0_outputs(2778) <= '1';
    layer0_outputs(2779) <= not((inputs(170)) or (inputs(85)));
    layer0_outputs(2780) <= inputs(198);
    layer0_outputs(2781) <= not((inputs(147)) xor (inputs(223)));
    layer0_outputs(2782) <= inputs(25);
    layer0_outputs(2783) <= inputs(194);
    layer0_outputs(2784) <= '1';
    layer0_outputs(2785) <= (inputs(160)) and not (inputs(228));
    layer0_outputs(2786) <= not(inputs(153));
    layer0_outputs(2787) <= not(inputs(78));
    layer0_outputs(2788) <= not(inputs(106)) or (inputs(250));
    layer0_outputs(2789) <= inputs(247);
    layer0_outputs(2790) <= inputs(231);
    layer0_outputs(2791) <= (inputs(154)) or (inputs(36));
    layer0_outputs(2792) <= (inputs(15)) and not (inputs(58));
    layer0_outputs(2793) <= not((inputs(191)) or (inputs(234)));
    layer0_outputs(2794) <= not(inputs(74));
    layer0_outputs(2795) <= '1';
    layer0_outputs(2796) <= not(inputs(154)) or (inputs(116));
    layer0_outputs(2797) <= not(inputs(50)) or (inputs(104));
    layer0_outputs(2798) <= '1';
    layer0_outputs(2799) <= (inputs(51)) or (inputs(185));
    layer0_outputs(2800) <= (inputs(210)) and not (inputs(179));
    layer0_outputs(2801) <= inputs(59);
    layer0_outputs(2802) <= not(inputs(142)) or (inputs(18));
    layer0_outputs(2803) <= not(inputs(3));
    layer0_outputs(2804) <= not((inputs(86)) or (inputs(67)));
    layer0_outputs(2805) <= (inputs(23)) or (inputs(189));
    layer0_outputs(2806) <= not(inputs(109)) or (inputs(164));
    layer0_outputs(2807) <= '0';
    layer0_outputs(2808) <= inputs(52);
    layer0_outputs(2809) <= not((inputs(251)) xor (inputs(137)));
    layer0_outputs(2810) <= not(inputs(221)) or (inputs(152));
    layer0_outputs(2811) <= inputs(107);
    layer0_outputs(2812) <= (inputs(204)) xor (inputs(65));
    layer0_outputs(2813) <= not(inputs(190)) or (inputs(246));
    layer0_outputs(2814) <= not((inputs(51)) and (inputs(34)));
    layer0_outputs(2815) <= inputs(102);
    layer0_outputs(2816) <= not(inputs(164));
    layer0_outputs(2817) <= inputs(164);
    layer0_outputs(2818) <= not(inputs(185)) or (inputs(25));
    layer0_outputs(2819) <= (inputs(123)) or (inputs(6));
    layer0_outputs(2820) <= '0';
    layer0_outputs(2821) <= (inputs(14)) and not (inputs(73));
    layer0_outputs(2822) <= inputs(148);
    layer0_outputs(2823) <= inputs(170);
    layer0_outputs(2824) <= (inputs(0)) and not (inputs(28));
    layer0_outputs(2825) <= not(inputs(193)) or (inputs(2));
    layer0_outputs(2826) <= (inputs(132)) or (inputs(220));
    layer0_outputs(2827) <= inputs(142);
    layer0_outputs(2828) <= inputs(255);
    layer0_outputs(2829) <= not(inputs(181)) or (inputs(27));
    layer0_outputs(2830) <= '0';
    layer0_outputs(2831) <= (inputs(104)) or (inputs(139));
    layer0_outputs(2832) <= '1';
    layer0_outputs(2833) <= inputs(16);
    layer0_outputs(2834) <= (inputs(141)) xor (inputs(190));
    layer0_outputs(2835) <= (inputs(214)) and not (inputs(28));
    layer0_outputs(2836) <= inputs(145);
    layer0_outputs(2837) <= not((inputs(233)) or (inputs(35)));
    layer0_outputs(2838) <= not((inputs(159)) xor (inputs(207)));
    layer0_outputs(2839) <= inputs(230);
    layer0_outputs(2840) <= inputs(119);
    layer0_outputs(2841) <= '1';
    layer0_outputs(2842) <= inputs(223);
    layer0_outputs(2843) <= not(inputs(120)) or (inputs(212));
    layer0_outputs(2844) <= (inputs(20)) or (inputs(182));
    layer0_outputs(2845) <= (inputs(26)) and not (inputs(172));
    layer0_outputs(2846) <= (inputs(17)) or (inputs(209));
    layer0_outputs(2847) <= not((inputs(191)) and (inputs(203)));
    layer0_outputs(2848) <= not(inputs(94)) or (inputs(24));
    layer0_outputs(2849) <= (inputs(174)) or (inputs(212));
    layer0_outputs(2850) <= not(inputs(24));
    layer0_outputs(2851) <= not((inputs(73)) and (inputs(234)));
    layer0_outputs(2852) <= not((inputs(167)) and (inputs(148)));
    layer0_outputs(2853) <= (inputs(30)) or (inputs(3));
    layer0_outputs(2854) <= not(inputs(135));
    layer0_outputs(2855) <= '1';
    layer0_outputs(2856) <= not(inputs(5)) or (inputs(103));
    layer0_outputs(2857) <= (inputs(108)) and not (inputs(237));
    layer0_outputs(2858) <= not((inputs(5)) and (inputs(71)));
    layer0_outputs(2859) <= '1';
    layer0_outputs(2860) <= (inputs(142)) and (inputs(41));
    layer0_outputs(2861) <= (inputs(158)) xor (inputs(82));
    layer0_outputs(2862) <= not(inputs(221)) or (inputs(61));
    layer0_outputs(2863) <= (inputs(104)) and not (inputs(65));
    layer0_outputs(2864) <= not((inputs(189)) or (inputs(47)));
    layer0_outputs(2865) <= '0';
    layer0_outputs(2866) <= (inputs(24)) and not (inputs(88));
    layer0_outputs(2867) <= not(inputs(176)) or (inputs(155));
    layer0_outputs(2868) <= not(inputs(90));
    layer0_outputs(2869) <= inputs(203);
    layer0_outputs(2870) <= inputs(167);
    layer0_outputs(2871) <= not(inputs(132));
    layer0_outputs(2872) <= inputs(17);
    layer0_outputs(2873) <= (inputs(129)) and (inputs(64));
    layer0_outputs(2874) <= '0';
    layer0_outputs(2875) <= (inputs(108)) and not (inputs(134));
    layer0_outputs(2876) <= '1';
    layer0_outputs(2877) <= (inputs(251)) and (inputs(189));
    layer0_outputs(2878) <= not((inputs(158)) and (inputs(113)));
    layer0_outputs(2879) <= not((inputs(27)) or (inputs(95)));
    layer0_outputs(2880) <= (inputs(234)) and not (inputs(30));
    layer0_outputs(2881) <= (inputs(87)) and (inputs(109));
    layer0_outputs(2882) <= '1';
    layer0_outputs(2883) <= (inputs(180)) and (inputs(38));
    layer0_outputs(2884) <= inputs(167);
    layer0_outputs(2885) <= (inputs(254)) and (inputs(208));
    layer0_outputs(2886) <= (inputs(138)) or (inputs(191));
    layer0_outputs(2887) <= inputs(16);
    layer0_outputs(2888) <= not(inputs(189));
    layer0_outputs(2889) <= '0';
    layer0_outputs(2890) <= not((inputs(19)) or (inputs(36)));
    layer0_outputs(2891) <= (inputs(219)) or (inputs(175));
    layer0_outputs(2892) <= not(inputs(115));
    layer0_outputs(2893) <= not(inputs(52)) or (inputs(249));
    layer0_outputs(2894) <= (inputs(149)) and (inputs(46));
    layer0_outputs(2895) <= inputs(76);
    layer0_outputs(2896) <= not(inputs(242)) or (inputs(55));
    layer0_outputs(2897) <= (inputs(69)) or (inputs(21));
    layer0_outputs(2898) <= '1';
    layer0_outputs(2899) <= (inputs(21)) or (inputs(22));
    layer0_outputs(2900) <= not((inputs(196)) xor (inputs(100)));
    layer0_outputs(2901) <= inputs(78);
    layer0_outputs(2902) <= not(inputs(212)) or (inputs(36));
    layer0_outputs(2903) <= not(inputs(166));
    layer0_outputs(2904) <= not(inputs(188)) or (inputs(140));
    layer0_outputs(2905) <= (inputs(169)) or (inputs(175));
    layer0_outputs(2906) <= not((inputs(30)) xor (inputs(75)));
    layer0_outputs(2907) <= (inputs(193)) xor (inputs(208));
    layer0_outputs(2908) <= inputs(250);
    layer0_outputs(2909) <= inputs(155);
    layer0_outputs(2910) <= not(inputs(127)) or (inputs(236));
    layer0_outputs(2911) <= not(inputs(127));
    layer0_outputs(2912) <= '1';
    layer0_outputs(2913) <= inputs(196);
    layer0_outputs(2914) <= not(inputs(189));
    layer0_outputs(2915) <= not(inputs(221)) or (inputs(47));
    layer0_outputs(2916) <= inputs(7);
    layer0_outputs(2917) <= (inputs(191)) or (inputs(73));
    layer0_outputs(2918) <= not(inputs(89)) or (inputs(8));
    layer0_outputs(2919) <= inputs(97);
    layer0_outputs(2920) <= not(inputs(190));
    layer0_outputs(2921) <= inputs(100);
    layer0_outputs(2922) <= (inputs(132)) and (inputs(207));
    layer0_outputs(2923) <= inputs(98);
    layer0_outputs(2924) <= '0';
    layer0_outputs(2925) <= (inputs(35)) or (inputs(73));
    layer0_outputs(2926) <= (inputs(205)) and (inputs(68));
    layer0_outputs(2927) <= not((inputs(108)) and (inputs(253)));
    layer0_outputs(2928) <= inputs(240);
    layer0_outputs(2929) <= (inputs(159)) and not (inputs(103));
    layer0_outputs(2930) <= not(inputs(180));
    layer0_outputs(2931) <= not(inputs(182)) or (inputs(93));
    layer0_outputs(2932) <= inputs(129);
    layer0_outputs(2933) <= (inputs(154)) and not (inputs(220));
    layer0_outputs(2934) <= not(inputs(17)) or (inputs(78));
    layer0_outputs(2935) <= inputs(118);
    layer0_outputs(2936) <= not(inputs(8));
    layer0_outputs(2937) <= not(inputs(148));
    layer0_outputs(2938) <= not(inputs(248)) or (inputs(44));
    layer0_outputs(2939) <= not(inputs(88));
    layer0_outputs(2940) <= inputs(101);
    layer0_outputs(2941) <= (inputs(86)) and not (inputs(206));
    layer0_outputs(2942) <= (inputs(72)) and not (inputs(177));
    layer0_outputs(2943) <= not((inputs(132)) xor (inputs(126)));
    layer0_outputs(2944) <= (inputs(37)) and (inputs(159));
    layer0_outputs(2945) <= inputs(170);
    layer0_outputs(2946) <= not(inputs(51)) or (inputs(167));
    layer0_outputs(2947) <= '1';
    layer0_outputs(2948) <= '1';
    layer0_outputs(2949) <= not(inputs(226));
    layer0_outputs(2950) <= '1';
    layer0_outputs(2951) <= '1';
    layer0_outputs(2952) <= not(inputs(227));
    layer0_outputs(2953) <= not(inputs(128));
    layer0_outputs(2954) <= (inputs(81)) and not (inputs(130));
    layer0_outputs(2955) <= not((inputs(252)) or (inputs(199)));
    layer0_outputs(2956) <= not(inputs(119));
    layer0_outputs(2957) <= inputs(64);
    layer0_outputs(2958) <= (inputs(209)) and not (inputs(103));
    layer0_outputs(2959) <= not(inputs(46)) or (inputs(87));
    layer0_outputs(2960) <= '1';
    layer0_outputs(2961) <= not((inputs(74)) or (inputs(92)));
    layer0_outputs(2962) <= not(inputs(226));
    layer0_outputs(2963) <= '1';
    layer0_outputs(2964) <= not(inputs(63));
    layer0_outputs(2965) <= inputs(240);
    layer0_outputs(2966) <= inputs(140);
    layer0_outputs(2967) <= inputs(159);
    layer0_outputs(2968) <= '1';
    layer0_outputs(2969) <= inputs(26);
    layer0_outputs(2970) <= not((inputs(4)) and (inputs(38)));
    layer0_outputs(2971) <= not((inputs(39)) or (inputs(191)));
    layer0_outputs(2972) <= '1';
    layer0_outputs(2973) <= '1';
    layer0_outputs(2974) <= not((inputs(249)) and (inputs(58)));
    layer0_outputs(2975) <= not((inputs(148)) or (inputs(147)));
    layer0_outputs(2976) <= not(inputs(21));
    layer0_outputs(2977) <= not(inputs(251));
    layer0_outputs(2978) <= '1';
    layer0_outputs(2979) <= (inputs(28)) and (inputs(120));
    layer0_outputs(2980) <= not((inputs(22)) or (inputs(105)));
    layer0_outputs(2981) <= not((inputs(224)) or (inputs(177)));
    layer0_outputs(2982) <= '1';
    layer0_outputs(2983) <= not((inputs(185)) or (inputs(118)));
    layer0_outputs(2984) <= not((inputs(98)) or (inputs(219)));
    layer0_outputs(2985) <= inputs(232);
    layer0_outputs(2986) <= '0';
    layer0_outputs(2987) <= not(inputs(116)) or (inputs(60));
    layer0_outputs(2988) <= inputs(74);
    layer0_outputs(2989) <= not(inputs(4)) or (inputs(97));
    layer0_outputs(2990) <= (inputs(150)) xor (inputs(252));
    layer0_outputs(2991) <= not((inputs(15)) or (inputs(95)));
    layer0_outputs(2992) <= inputs(117);
    layer0_outputs(2993) <= not(inputs(9)) or (inputs(180));
    layer0_outputs(2994) <= '1';
    layer0_outputs(2995) <= not(inputs(145));
    layer0_outputs(2996) <= inputs(105);
    layer0_outputs(2997) <= (inputs(3)) and not (inputs(67));
    layer0_outputs(2998) <= (inputs(116)) xor (inputs(34));
    layer0_outputs(2999) <= (inputs(88)) or (inputs(116));
    layer0_outputs(3000) <= not(inputs(17));
    layer0_outputs(3001) <= '0';
    layer0_outputs(3002) <= inputs(118);
    layer0_outputs(3003) <= '1';
    layer0_outputs(3004) <= inputs(96);
    layer0_outputs(3005) <= not(inputs(136));
    layer0_outputs(3006) <= not((inputs(74)) or (inputs(186)));
    layer0_outputs(3007) <= inputs(251);
    layer0_outputs(3008) <= (inputs(10)) or (inputs(203));
    layer0_outputs(3009) <= not(inputs(90)) or (inputs(81));
    layer0_outputs(3010) <= (inputs(95)) xor (inputs(198));
    layer0_outputs(3011) <= not(inputs(7));
    layer0_outputs(3012) <= not(inputs(187));
    layer0_outputs(3013) <= not((inputs(156)) or (inputs(37)));
    layer0_outputs(3014) <= inputs(187);
    layer0_outputs(3015) <= (inputs(111)) and not (inputs(17));
    layer0_outputs(3016) <= not(inputs(194));
    layer0_outputs(3017) <= (inputs(199)) or (inputs(125));
    layer0_outputs(3018) <= not(inputs(122)) or (inputs(158));
    layer0_outputs(3019) <= (inputs(206)) xor (inputs(206));
    layer0_outputs(3020) <= not(inputs(116)) or (inputs(11));
    layer0_outputs(3021) <= (inputs(125)) and not (inputs(155));
    layer0_outputs(3022) <= not((inputs(115)) or (inputs(125)));
    layer0_outputs(3023) <= not(inputs(146)) or (inputs(163));
    layer0_outputs(3024) <= (inputs(205)) xor (inputs(37));
    layer0_outputs(3025) <= not(inputs(167)) or (inputs(253));
    layer0_outputs(3026) <= not((inputs(87)) and (inputs(220)));
    layer0_outputs(3027) <= (inputs(87)) and not (inputs(204));
    layer0_outputs(3028) <= '0';
    layer0_outputs(3029) <= '0';
    layer0_outputs(3030) <= '1';
    layer0_outputs(3031) <= '1';
    layer0_outputs(3032) <= (inputs(106)) and (inputs(170));
    layer0_outputs(3033) <= inputs(59);
    layer0_outputs(3034) <= '0';
    layer0_outputs(3035) <= (inputs(47)) xor (inputs(207));
    layer0_outputs(3036) <= (inputs(232)) and not (inputs(151));
    layer0_outputs(3037) <= not((inputs(137)) xor (inputs(15)));
    layer0_outputs(3038) <= inputs(207);
    layer0_outputs(3039) <= (inputs(7)) and not (inputs(12));
    layer0_outputs(3040) <= '1';
    layer0_outputs(3041) <= not(inputs(210));
    layer0_outputs(3042) <= not(inputs(66));
    layer0_outputs(3043) <= inputs(69);
    layer0_outputs(3044) <= '0';
    layer0_outputs(3045) <= (inputs(135)) and not (inputs(155));
    layer0_outputs(3046) <= not(inputs(192)) or (inputs(73));
    layer0_outputs(3047) <= inputs(17);
    layer0_outputs(3048) <= (inputs(193)) and not (inputs(163));
    layer0_outputs(3049) <= (inputs(128)) and not (inputs(219));
    layer0_outputs(3050) <= (inputs(171)) xor (inputs(67));
    layer0_outputs(3051) <= not(inputs(204));
    layer0_outputs(3052) <= (inputs(179)) and not (inputs(224));
    layer0_outputs(3053) <= (inputs(5)) and not (inputs(160));
    layer0_outputs(3054) <= (inputs(70)) and not (inputs(62));
    layer0_outputs(3055) <= not(inputs(77));
    layer0_outputs(3056) <= not((inputs(202)) and (inputs(134)));
    layer0_outputs(3057) <= '1';
    layer0_outputs(3058) <= not(inputs(146));
    layer0_outputs(3059) <= (inputs(67)) or (inputs(116));
    layer0_outputs(3060) <= not(inputs(234));
    layer0_outputs(3061) <= inputs(202);
    layer0_outputs(3062) <= '0';
    layer0_outputs(3063) <= not((inputs(244)) and (inputs(143)));
    layer0_outputs(3064) <= not((inputs(147)) or (inputs(186)));
    layer0_outputs(3065) <= not(inputs(179)) or (inputs(49));
    layer0_outputs(3066) <= (inputs(246)) and (inputs(49));
    layer0_outputs(3067) <= not(inputs(176));
    layer0_outputs(3068) <= inputs(137);
    layer0_outputs(3069) <= not(inputs(136)) or (inputs(91));
    layer0_outputs(3070) <= (inputs(49)) and not (inputs(62));
    layer0_outputs(3071) <= not((inputs(101)) or (inputs(9)));
    layer0_outputs(3072) <= not(inputs(88)) or (inputs(140));
    layer0_outputs(3073) <= not((inputs(31)) or (inputs(35)));
    layer0_outputs(3074) <= '1';
    layer0_outputs(3075) <= '0';
    layer0_outputs(3076) <= not(inputs(217)) or (inputs(191));
    layer0_outputs(3077) <= (inputs(115)) xor (inputs(162));
    layer0_outputs(3078) <= not(inputs(48));
    layer0_outputs(3079) <= not(inputs(16)) or (inputs(247));
    layer0_outputs(3080) <= '0';
    layer0_outputs(3081) <= (inputs(154)) and not (inputs(77));
    layer0_outputs(3082) <= (inputs(4)) and not (inputs(241));
    layer0_outputs(3083) <= '0';
    layer0_outputs(3084) <= (inputs(193)) and not (inputs(150));
    layer0_outputs(3085) <= (inputs(235)) and (inputs(201));
    layer0_outputs(3086) <= (inputs(64)) and not (inputs(116));
    layer0_outputs(3087) <= not(inputs(255)) or (inputs(155));
    layer0_outputs(3088) <= not(inputs(18));
    layer0_outputs(3089) <= (inputs(62)) or (inputs(0));
    layer0_outputs(3090) <= (inputs(174)) or (inputs(34));
    layer0_outputs(3091) <= '1';
    layer0_outputs(3092) <= not((inputs(82)) or (inputs(38)));
    layer0_outputs(3093) <= not((inputs(100)) xor (inputs(103)));
    layer0_outputs(3094) <= inputs(71);
    layer0_outputs(3095) <= inputs(93);
    layer0_outputs(3096) <= '1';
    layer0_outputs(3097) <= not((inputs(64)) and (inputs(50)));
    layer0_outputs(3098) <= '1';
    layer0_outputs(3099) <= '0';
    layer0_outputs(3100) <= inputs(138);
    layer0_outputs(3101) <= not((inputs(63)) or (inputs(215)));
    layer0_outputs(3102) <= inputs(229);
    layer0_outputs(3103) <= not((inputs(29)) and (inputs(175)));
    layer0_outputs(3104) <= '0';
    layer0_outputs(3105) <= (inputs(67)) and (inputs(160));
    layer0_outputs(3106) <= not(inputs(64)) or (inputs(42));
    layer0_outputs(3107) <= not((inputs(153)) and (inputs(188)));
    layer0_outputs(3108) <= '0';
    layer0_outputs(3109) <= inputs(102);
    layer0_outputs(3110) <= (inputs(216)) and (inputs(117));
    layer0_outputs(3111) <= (inputs(127)) or (inputs(50));
    layer0_outputs(3112) <= not(inputs(168)) or (inputs(102));
    layer0_outputs(3113) <= (inputs(16)) and not (inputs(126));
    layer0_outputs(3114) <= not((inputs(239)) or (inputs(75)));
    layer0_outputs(3115) <= not(inputs(162));
    layer0_outputs(3116) <= '1';
    layer0_outputs(3117) <= (inputs(78)) and not (inputs(27));
    layer0_outputs(3118) <= (inputs(43)) and not (inputs(43));
    layer0_outputs(3119) <= not(inputs(220)) or (inputs(110));
    layer0_outputs(3120) <= '0';
    layer0_outputs(3121) <= not((inputs(201)) and (inputs(183)));
    layer0_outputs(3122) <= not((inputs(192)) or (inputs(202)));
    layer0_outputs(3123) <= not((inputs(222)) xor (inputs(209)));
    layer0_outputs(3124) <= '0';
    layer0_outputs(3125) <= (inputs(18)) or (inputs(109));
    layer0_outputs(3126) <= not(inputs(254)) or (inputs(124));
    layer0_outputs(3127) <= not(inputs(26));
    layer0_outputs(3128) <= inputs(20);
    layer0_outputs(3129) <= (inputs(217)) and not (inputs(128));
    layer0_outputs(3130) <= inputs(222);
    layer0_outputs(3131) <= (inputs(244)) or (inputs(91));
    layer0_outputs(3132) <= not((inputs(9)) or (inputs(120)));
    layer0_outputs(3133) <= not(inputs(122));
    layer0_outputs(3134) <= (inputs(75)) xor (inputs(63));
    layer0_outputs(3135) <= (inputs(74)) and not (inputs(32));
    layer0_outputs(3136) <= not(inputs(134));
    layer0_outputs(3137) <= '1';
    layer0_outputs(3138) <= not(inputs(92));
    layer0_outputs(3139) <= not(inputs(210));
    layer0_outputs(3140) <= not(inputs(93)) or (inputs(34));
    layer0_outputs(3141) <= '0';
    layer0_outputs(3142) <= not(inputs(28));
    layer0_outputs(3143) <= not(inputs(208)) or (inputs(107));
    layer0_outputs(3144) <= inputs(227);
    layer0_outputs(3145) <= (inputs(206)) and not (inputs(95));
    layer0_outputs(3146) <= '1';
    layer0_outputs(3147) <= '1';
    layer0_outputs(3148) <= not(inputs(45));
    layer0_outputs(3149) <= '1';
    layer0_outputs(3150) <= not(inputs(25));
    layer0_outputs(3151) <= not(inputs(80)) or (inputs(94));
    layer0_outputs(3152) <= not((inputs(206)) or (inputs(220)));
    layer0_outputs(3153) <= (inputs(249)) or (inputs(231));
    layer0_outputs(3154) <= '0';
    layer0_outputs(3155) <= (inputs(120)) and not (inputs(250));
    layer0_outputs(3156) <= (inputs(177)) or (inputs(216));
    layer0_outputs(3157) <= (inputs(239)) and (inputs(136));
    layer0_outputs(3158) <= (inputs(22)) or (inputs(3));
    layer0_outputs(3159) <= (inputs(193)) or (inputs(21));
    layer0_outputs(3160) <= not((inputs(0)) or (inputs(160)));
    layer0_outputs(3161) <= not(inputs(55));
    layer0_outputs(3162) <= '0';
    layer0_outputs(3163) <= not(inputs(135));
    layer0_outputs(3164) <= not((inputs(63)) or (inputs(95)));
    layer0_outputs(3165) <= (inputs(147)) or (inputs(162));
    layer0_outputs(3166) <= (inputs(243)) and not (inputs(81));
    layer0_outputs(3167) <= '0';
    layer0_outputs(3168) <= '0';
    layer0_outputs(3169) <= (inputs(98)) or (inputs(117));
    layer0_outputs(3170) <= '1';
    layer0_outputs(3171) <= not(inputs(247));
    layer0_outputs(3172) <= inputs(190);
    layer0_outputs(3173) <= not((inputs(246)) or (inputs(128)));
    layer0_outputs(3174) <= inputs(203);
    layer0_outputs(3175) <= '1';
    layer0_outputs(3176) <= not((inputs(211)) or (inputs(16)));
    layer0_outputs(3177) <= (inputs(139)) or (inputs(191));
    layer0_outputs(3178) <= not(inputs(117)) or (inputs(18));
    layer0_outputs(3179) <= (inputs(23)) and (inputs(75));
    layer0_outputs(3180) <= '1';
    layer0_outputs(3181) <= inputs(60);
    layer0_outputs(3182) <= (inputs(175)) or (inputs(233));
    layer0_outputs(3183) <= not(inputs(147)) or (inputs(10));
    layer0_outputs(3184) <= not(inputs(123));
    layer0_outputs(3185) <= (inputs(138)) and not (inputs(212));
    layer0_outputs(3186) <= not(inputs(240)) or (inputs(144));
    layer0_outputs(3187) <= not(inputs(113));
    layer0_outputs(3188) <= inputs(114);
    layer0_outputs(3189) <= not(inputs(0));
    layer0_outputs(3190) <= not(inputs(166));
    layer0_outputs(3191) <= (inputs(143)) or (inputs(92));
    layer0_outputs(3192) <= not(inputs(52)) or (inputs(32));
    layer0_outputs(3193) <= '1';
    layer0_outputs(3194) <= '1';
    layer0_outputs(3195) <= inputs(57);
    layer0_outputs(3196) <= not(inputs(169));
    layer0_outputs(3197) <= (inputs(166)) and not (inputs(101));
    layer0_outputs(3198) <= (inputs(73)) or (inputs(193));
    layer0_outputs(3199) <= '0';
    layer0_outputs(3200) <= inputs(225);
    layer0_outputs(3201) <= (inputs(110)) and (inputs(85));
    layer0_outputs(3202) <= inputs(106);
    layer0_outputs(3203) <= not(inputs(35));
    layer0_outputs(3204) <= not(inputs(114));
    layer0_outputs(3205) <= '0';
    layer0_outputs(3206) <= not((inputs(126)) and (inputs(82)));
    layer0_outputs(3207) <= '1';
    layer0_outputs(3208) <= inputs(227);
    layer0_outputs(3209) <= (inputs(162)) or (inputs(107));
    layer0_outputs(3210) <= inputs(192);
    layer0_outputs(3211) <= not(inputs(139)) or (inputs(34));
    layer0_outputs(3212) <= (inputs(253)) and not (inputs(113));
    layer0_outputs(3213) <= not((inputs(37)) or (inputs(193)));
    layer0_outputs(3214) <= (inputs(138)) or (inputs(84));
    layer0_outputs(3215) <= not(inputs(225)) or (inputs(129));
    layer0_outputs(3216) <= inputs(131);
    layer0_outputs(3217) <= not((inputs(215)) or (inputs(5)));
    layer0_outputs(3218) <= inputs(18);
    layer0_outputs(3219) <= inputs(175);
    layer0_outputs(3220) <= '0';
    layer0_outputs(3221) <= '1';
    layer0_outputs(3222) <= (inputs(28)) or (inputs(168));
    layer0_outputs(3223) <= not(inputs(142));
    layer0_outputs(3224) <= not((inputs(231)) or (inputs(232)));
    layer0_outputs(3225) <= not((inputs(153)) xor (inputs(128)));
    layer0_outputs(3226) <= (inputs(79)) or (inputs(67));
    layer0_outputs(3227) <= inputs(133);
    layer0_outputs(3228) <= (inputs(86)) and (inputs(51));
    layer0_outputs(3229) <= inputs(223);
    layer0_outputs(3230) <= not((inputs(18)) or (inputs(117)));
    layer0_outputs(3231) <= inputs(231);
    layer0_outputs(3232) <= (inputs(153)) xor (inputs(47));
    layer0_outputs(3233) <= not((inputs(211)) xor (inputs(174)));
    layer0_outputs(3234) <= (inputs(252)) or (inputs(213));
    layer0_outputs(3235) <= (inputs(1)) or (inputs(23));
    layer0_outputs(3236) <= not(inputs(111)) or (inputs(251));
    layer0_outputs(3237) <= not(inputs(176));
    layer0_outputs(3238) <= (inputs(86)) and (inputs(238));
    layer0_outputs(3239) <= not(inputs(208));
    layer0_outputs(3240) <= (inputs(210)) or (inputs(79));
    layer0_outputs(3241) <= '0';
    layer0_outputs(3242) <= (inputs(24)) or (inputs(239));
    layer0_outputs(3243) <= not((inputs(136)) and (inputs(124)));
    layer0_outputs(3244) <= '0';
    layer0_outputs(3245) <= '0';
    layer0_outputs(3246) <= '0';
    layer0_outputs(3247) <= '0';
    layer0_outputs(3248) <= not(inputs(151)) or (inputs(186));
    layer0_outputs(3249) <= not(inputs(206));
    layer0_outputs(3250) <= (inputs(198)) and (inputs(100));
    layer0_outputs(3251) <= '1';
    layer0_outputs(3252) <= inputs(113);
    layer0_outputs(3253) <= (inputs(18)) or (inputs(28));
    layer0_outputs(3254) <= not(inputs(104)) or (inputs(110));
    layer0_outputs(3255) <= (inputs(193)) and not (inputs(58));
    layer0_outputs(3256) <= not((inputs(142)) or (inputs(208)));
    layer0_outputs(3257) <= inputs(100);
    layer0_outputs(3258) <= (inputs(219)) or (inputs(254));
    layer0_outputs(3259) <= not(inputs(124)) or (inputs(54));
    layer0_outputs(3260) <= (inputs(48)) and not (inputs(151));
    layer0_outputs(3261) <= (inputs(19)) or (inputs(20));
    layer0_outputs(3262) <= (inputs(120)) and not (inputs(94));
    layer0_outputs(3263) <= not(inputs(184));
    layer0_outputs(3264) <= not((inputs(129)) or (inputs(55)));
    layer0_outputs(3265) <= inputs(231);
    layer0_outputs(3266) <= '1';
    layer0_outputs(3267) <= inputs(177);
    layer0_outputs(3268) <= '0';
    layer0_outputs(3269) <= (inputs(1)) or (inputs(34));
    layer0_outputs(3270) <= not(inputs(166)) or (inputs(63));
    layer0_outputs(3271) <= '1';
    layer0_outputs(3272) <= (inputs(72)) and not (inputs(188));
    layer0_outputs(3273) <= not(inputs(19));
    layer0_outputs(3274) <= not((inputs(167)) or (inputs(241)));
    layer0_outputs(3275) <= (inputs(69)) or (inputs(33));
    layer0_outputs(3276) <= '1';
    layer0_outputs(3277) <= not((inputs(93)) or (inputs(193)));
    layer0_outputs(3278) <= (inputs(82)) or (inputs(132));
    layer0_outputs(3279) <= not((inputs(187)) or (inputs(132)));
    layer0_outputs(3280) <= (inputs(176)) and not (inputs(240));
    layer0_outputs(3281) <= not(inputs(15));
    layer0_outputs(3282) <= (inputs(207)) xor (inputs(4));
    layer0_outputs(3283) <= inputs(111);
    layer0_outputs(3284) <= not((inputs(22)) xor (inputs(98)));
    layer0_outputs(3285) <= (inputs(7)) and not (inputs(159));
    layer0_outputs(3286) <= (inputs(72)) and not (inputs(94));
    layer0_outputs(3287) <= (inputs(0)) and not (inputs(83));
    layer0_outputs(3288) <= not(inputs(40));
    layer0_outputs(3289) <= (inputs(60)) and (inputs(73));
    layer0_outputs(3290) <= not(inputs(8)) or (inputs(246));
    layer0_outputs(3291) <= not(inputs(49));
    layer0_outputs(3292) <= not(inputs(206));
    layer0_outputs(3293) <= (inputs(182)) and not (inputs(132));
    layer0_outputs(3294) <= (inputs(184)) and not (inputs(88));
    layer0_outputs(3295) <= inputs(122);
    layer0_outputs(3296) <= not(inputs(241));
    layer0_outputs(3297) <= (inputs(110)) and not (inputs(200));
    layer0_outputs(3298) <= (inputs(180)) and not (inputs(3));
    layer0_outputs(3299) <= not(inputs(75)) or (inputs(255));
    layer0_outputs(3300) <= (inputs(48)) and not (inputs(61));
    layer0_outputs(3301) <= (inputs(247)) and not (inputs(92));
    layer0_outputs(3302) <= not(inputs(15));
    layer0_outputs(3303) <= not(inputs(217));
    layer0_outputs(3304) <= not(inputs(105)) or (inputs(14));
    layer0_outputs(3305) <= '0';
    layer0_outputs(3306) <= not((inputs(33)) or (inputs(247)));
    layer0_outputs(3307) <= (inputs(254)) or (inputs(215));
    layer0_outputs(3308) <= not(inputs(61));
    layer0_outputs(3309) <= not(inputs(17));
    layer0_outputs(3310) <= '1';
    layer0_outputs(3311) <= not(inputs(133));
    layer0_outputs(3312) <= (inputs(15)) or (inputs(105));
    layer0_outputs(3313) <= not(inputs(92)) or (inputs(217));
    layer0_outputs(3314) <= inputs(210);
    layer0_outputs(3315) <= (inputs(39)) xor (inputs(169));
    layer0_outputs(3316) <= not(inputs(97));
    layer0_outputs(3317) <= '1';
    layer0_outputs(3318) <= '1';
    layer0_outputs(3319) <= not((inputs(124)) or (inputs(144)));
    layer0_outputs(3320) <= inputs(171);
    layer0_outputs(3321) <= not(inputs(209)) or (inputs(112));
    layer0_outputs(3322) <= not((inputs(213)) and (inputs(168)));
    layer0_outputs(3323) <= inputs(63);
    layer0_outputs(3324) <= (inputs(121)) and not (inputs(249));
    layer0_outputs(3325) <= inputs(161);
    layer0_outputs(3326) <= not((inputs(60)) or (inputs(46)));
    layer0_outputs(3327) <= '1';
    layer0_outputs(3328) <= not((inputs(68)) xor (inputs(174)));
    layer0_outputs(3329) <= inputs(214);
    layer0_outputs(3330) <= inputs(221);
    layer0_outputs(3331) <= (inputs(138)) and not (inputs(246));
    layer0_outputs(3332) <= '0';
    layer0_outputs(3333) <= '0';
    layer0_outputs(3334) <= not((inputs(73)) or (inputs(70)));
    layer0_outputs(3335) <= inputs(184);
    layer0_outputs(3336) <= not(inputs(1)) or (inputs(198));
    layer0_outputs(3337) <= (inputs(71)) and (inputs(86));
    layer0_outputs(3338) <= (inputs(31)) and not (inputs(95));
    layer0_outputs(3339) <= not(inputs(96)) or (inputs(158));
    layer0_outputs(3340) <= (inputs(248)) xor (inputs(31));
    layer0_outputs(3341) <= inputs(104);
    layer0_outputs(3342) <= inputs(159);
    layer0_outputs(3343) <= '0';
    layer0_outputs(3344) <= inputs(6);
    layer0_outputs(3345) <= not((inputs(14)) or (inputs(172)));
    layer0_outputs(3346) <= (inputs(105)) and not (inputs(3));
    layer0_outputs(3347) <= (inputs(14)) and not (inputs(191));
    layer0_outputs(3348) <= (inputs(208)) and not (inputs(112));
    layer0_outputs(3349) <= not((inputs(88)) or (inputs(117)));
    layer0_outputs(3350) <= (inputs(246)) or (inputs(63));
    layer0_outputs(3351) <= (inputs(224)) and not (inputs(122));
    layer0_outputs(3352) <= (inputs(109)) and not (inputs(164));
    layer0_outputs(3353) <= '0';
    layer0_outputs(3354) <= not(inputs(102));
    layer0_outputs(3355) <= '1';
    layer0_outputs(3356) <= not((inputs(202)) or (inputs(207)));
    layer0_outputs(3357) <= not(inputs(179));
    layer0_outputs(3358) <= '1';
    layer0_outputs(3359) <= '0';
    layer0_outputs(3360) <= (inputs(133)) and not (inputs(186));
    layer0_outputs(3361) <= inputs(117);
    layer0_outputs(3362) <= (inputs(209)) and not (inputs(147));
    layer0_outputs(3363) <= '0';
    layer0_outputs(3364) <= inputs(222);
    layer0_outputs(3365) <= (inputs(104)) and not (inputs(209));
    layer0_outputs(3366) <= inputs(252);
    layer0_outputs(3367) <= (inputs(16)) xor (inputs(238));
    layer0_outputs(3368) <= inputs(230);
    layer0_outputs(3369) <= not((inputs(67)) or (inputs(187)));
    layer0_outputs(3370) <= (inputs(135)) and not (inputs(137));
    layer0_outputs(3371) <= (inputs(201)) or (inputs(214));
    layer0_outputs(3372) <= (inputs(92)) and (inputs(4));
    layer0_outputs(3373) <= not((inputs(60)) or (inputs(35)));
    layer0_outputs(3374) <= not((inputs(216)) or (inputs(76)));
    layer0_outputs(3375) <= inputs(213);
    layer0_outputs(3376) <= (inputs(31)) and (inputs(77));
    layer0_outputs(3377) <= inputs(231);
    layer0_outputs(3378) <= inputs(163);
    layer0_outputs(3379) <= (inputs(6)) or (inputs(21));
    layer0_outputs(3380) <= inputs(74);
    layer0_outputs(3381) <= (inputs(182)) xor (inputs(163));
    layer0_outputs(3382) <= (inputs(233)) and (inputs(148));
    layer0_outputs(3383) <= (inputs(178)) and (inputs(243));
    layer0_outputs(3384) <= not(inputs(197));
    layer0_outputs(3385) <= inputs(134);
    layer0_outputs(3386) <= not(inputs(107));
    layer0_outputs(3387) <= not((inputs(225)) xor (inputs(1)));
    layer0_outputs(3388) <= inputs(109);
    layer0_outputs(3389) <= (inputs(231)) and (inputs(126));
    layer0_outputs(3390) <= not(inputs(227));
    layer0_outputs(3391) <= inputs(32);
    layer0_outputs(3392) <= not(inputs(116)) or (inputs(123));
    layer0_outputs(3393) <= (inputs(183)) and not (inputs(36));
    layer0_outputs(3394) <= (inputs(226)) and (inputs(193));
    layer0_outputs(3395) <= (inputs(12)) and not (inputs(203));
    layer0_outputs(3396) <= not(inputs(68)) or (inputs(220));
    layer0_outputs(3397) <= inputs(61);
    layer0_outputs(3398) <= (inputs(27)) and not (inputs(198));
    layer0_outputs(3399) <= (inputs(138)) xor (inputs(36));
    layer0_outputs(3400) <= not(inputs(191));
    layer0_outputs(3401) <= inputs(22);
    layer0_outputs(3402) <= not((inputs(20)) and (inputs(197)));
    layer0_outputs(3403) <= not(inputs(178)) or (inputs(47));
    layer0_outputs(3404) <= (inputs(51)) and not (inputs(218));
    layer0_outputs(3405) <= '0';
    layer0_outputs(3406) <= (inputs(191)) xor (inputs(160));
    layer0_outputs(3407) <= not(inputs(178));
    layer0_outputs(3408) <= (inputs(142)) and not (inputs(135));
    layer0_outputs(3409) <= inputs(135);
    layer0_outputs(3410) <= not((inputs(115)) or (inputs(113)));
    layer0_outputs(3411) <= not(inputs(188));
    layer0_outputs(3412) <= (inputs(253)) xor (inputs(248));
    layer0_outputs(3413) <= (inputs(102)) and not (inputs(84));
    layer0_outputs(3414) <= '1';
    layer0_outputs(3415) <= not((inputs(52)) and (inputs(154)));
    layer0_outputs(3416) <= inputs(127);
    layer0_outputs(3417) <= (inputs(237)) or (inputs(208));
    layer0_outputs(3418) <= not((inputs(236)) and (inputs(74)));
    layer0_outputs(3419) <= '0';
    layer0_outputs(3420) <= not(inputs(35)) or (inputs(94));
    layer0_outputs(3421) <= inputs(6);
    layer0_outputs(3422) <= not(inputs(45));
    layer0_outputs(3423) <= not((inputs(141)) or (inputs(3)));
    layer0_outputs(3424) <= inputs(121);
    layer0_outputs(3425) <= (inputs(150)) and not (inputs(247));
    layer0_outputs(3426) <= not(inputs(92));
    layer0_outputs(3427) <= not(inputs(49));
    layer0_outputs(3428) <= not((inputs(229)) or (inputs(47)));
    layer0_outputs(3429) <= '1';
    layer0_outputs(3430) <= not(inputs(88)) or (inputs(59));
    layer0_outputs(3431) <= not(inputs(56)) or (inputs(85));
    layer0_outputs(3432) <= not(inputs(205));
    layer0_outputs(3433) <= not(inputs(189));
    layer0_outputs(3434) <= not(inputs(212));
    layer0_outputs(3435) <= '0';
    layer0_outputs(3436) <= (inputs(254)) and not (inputs(95));
    layer0_outputs(3437) <= not(inputs(139)) or (inputs(216));
    layer0_outputs(3438) <= not((inputs(70)) or (inputs(233)));
    layer0_outputs(3439) <= (inputs(35)) or (inputs(225));
    layer0_outputs(3440) <= '1';
    layer0_outputs(3441) <= not(inputs(180)) or (inputs(54));
    layer0_outputs(3442) <= inputs(55);
    layer0_outputs(3443) <= not(inputs(42));
    layer0_outputs(3444) <= (inputs(253)) or (inputs(193));
    layer0_outputs(3445) <= not(inputs(19)) or (inputs(192));
    layer0_outputs(3446) <= '0';
    layer0_outputs(3447) <= not(inputs(161)) or (inputs(108));
    layer0_outputs(3448) <= (inputs(251)) or (inputs(92));
    layer0_outputs(3449) <= not((inputs(221)) and (inputs(134)));
    layer0_outputs(3450) <= (inputs(66)) and not (inputs(77));
    layer0_outputs(3451) <= '1';
    layer0_outputs(3452) <= inputs(157);
    layer0_outputs(3453) <= '0';
    layer0_outputs(3454) <= not((inputs(2)) and (inputs(150)));
    layer0_outputs(3455) <= (inputs(82)) and not (inputs(213));
    layer0_outputs(3456) <= not((inputs(183)) or (inputs(200)));
    layer0_outputs(3457) <= (inputs(244)) or (inputs(47));
    layer0_outputs(3458) <= '1';
    layer0_outputs(3459) <= not(inputs(138));
    layer0_outputs(3460) <= '0';
    layer0_outputs(3461) <= not((inputs(87)) or (inputs(97)));
    layer0_outputs(3462) <= not(inputs(82)) or (inputs(207));
    layer0_outputs(3463) <= not(inputs(187)) or (inputs(130));
    layer0_outputs(3464) <= not(inputs(72));
    layer0_outputs(3465) <= '0';
    layer0_outputs(3466) <= not((inputs(188)) and (inputs(190)));
    layer0_outputs(3467) <= '0';
    layer0_outputs(3468) <= not(inputs(232)) or (inputs(50));
    layer0_outputs(3469) <= inputs(99);
    layer0_outputs(3470) <= not(inputs(171));
    layer0_outputs(3471) <= '1';
    layer0_outputs(3472) <= not(inputs(62)) or (inputs(170));
    layer0_outputs(3473) <= not((inputs(193)) or (inputs(196)));
    layer0_outputs(3474) <= '0';
    layer0_outputs(3475) <= not((inputs(141)) and (inputs(242)));
    layer0_outputs(3476) <= '1';
    layer0_outputs(3477) <= (inputs(247)) and not (inputs(141));
    layer0_outputs(3478) <= inputs(52);
    layer0_outputs(3479) <= not((inputs(61)) or (inputs(127)));
    layer0_outputs(3480) <= '0';
    layer0_outputs(3481) <= (inputs(75)) or (inputs(128));
    layer0_outputs(3482) <= not(inputs(210));
    layer0_outputs(3483) <= not((inputs(208)) and (inputs(65)));
    layer0_outputs(3484) <= (inputs(98)) or (inputs(249));
    layer0_outputs(3485) <= inputs(67);
    layer0_outputs(3486) <= (inputs(193)) and not (inputs(45));
    layer0_outputs(3487) <= '1';
    layer0_outputs(3488) <= not(inputs(61)) or (inputs(185));
    layer0_outputs(3489) <= not(inputs(133)) or (inputs(134));
    layer0_outputs(3490) <= (inputs(50)) and (inputs(162));
    layer0_outputs(3491) <= not(inputs(136)) or (inputs(160));
    layer0_outputs(3492) <= (inputs(51)) xor (inputs(95));
    layer0_outputs(3493) <= not((inputs(29)) or (inputs(82)));
    layer0_outputs(3494) <= (inputs(31)) and not (inputs(249));
    layer0_outputs(3495) <= inputs(7);
    layer0_outputs(3496) <= inputs(88);
    layer0_outputs(3497) <= inputs(173);
    layer0_outputs(3498) <= not((inputs(153)) and (inputs(183)));
    layer0_outputs(3499) <= not(inputs(133));
    layer0_outputs(3500) <= (inputs(176)) or (inputs(181));
    layer0_outputs(3501) <= not(inputs(133)) or (inputs(31));
    layer0_outputs(3502) <= (inputs(64)) or (inputs(84));
    layer0_outputs(3503) <= inputs(167);
    layer0_outputs(3504) <= (inputs(208)) and (inputs(102));
    layer0_outputs(3505) <= inputs(246);
    layer0_outputs(3506) <= not(inputs(127)) or (inputs(31));
    layer0_outputs(3507) <= '1';
    layer0_outputs(3508) <= (inputs(28)) or (inputs(197));
    layer0_outputs(3509) <= (inputs(69)) and not (inputs(250));
    layer0_outputs(3510) <= '0';
    layer0_outputs(3511) <= inputs(55);
    layer0_outputs(3512) <= not(inputs(55));
    layer0_outputs(3513) <= not(inputs(28)) or (inputs(132));
    layer0_outputs(3514) <= not((inputs(203)) or (inputs(144)));
    layer0_outputs(3515) <= '1';
    layer0_outputs(3516) <= (inputs(116)) and not (inputs(175));
    layer0_outputs(3517) <= '1';
    layer0_outputs(3518) <= not(inputs(214)) or (inputs(207));
    layer0_outputs(3519) <= not((inputs(59)) or (inputs(123)));
    layer0_outputs(3520) <= (inputs(66)) xor (inputs(115));
    layer0_outputs(3521) <= '0';
    layer0_outputs(3522) <= (inputs(36)) xor (inputs(124));
    layer0_outputs(3523) <= not((inputs(41)) xor (inputs(165)));
    layer0_outputs(3524) <= not((inputs(129)) xor (inputs(25)));
    layer0_outputs(3525) <= inputs(235);
    layer0_outputs(3526) <= '1';
    layer0_outputs(3527) <= '0';
    layer0_outputs(3528) <= not(inputs(217)) or (inputs(17));
    layer0_outputs(3529) <= (inputs(22)) and not (inputs(48));
    layer0_outputs(3530) <= not(inputs(126)) or (inputs(107));
    layer0_outputs(3531) <= (inputs(23)) or (inputs(1));
    layer0_outputs(3532) <= (inputs(207)) or (inputs(23));
    layer0_outputs(3533) <= not(inputs(107));
    layer0_outputs(3534) <= (inputs(124)) and (inputs(45));
    layer0_outputs(3535) <= inputs(19);
    layer0_outputs(3536) <= (inputs(85)) xor (inputs(157));
    layer0_outputs(3537) <= '1';
    layer0_outputs(3538) <= '1';
    layer0_outputs(3539) <= not((inputs(14)) or (inputs(215)));
    layer0_outputs(3540) <= (inputs(94)) and not (inputs(238));
    layer0_outputs(3541) <= (inputs(226)) and not (inputs(127));
    layer0_outputs(3542) <= '1';
    layer0_outputs(3543) <= not((inputs(144)) xor (inputs(149)));
    layer0_outputs(3544) <= '1';
    layer0_outputs(3545) <= (inputs(222)) and not (inputs(75));
    layer0_outputs(3546) <= '0';
    layer0_outputs(3547) <= not(inputs(24)) or (inputs(87));
    layer0_outputs(3548) <= (inputs(70)) and not (inputs(111));
    layer0_outputs(3549) <= not((inputs(191)) or (inputs(184)));
    layer0_outputs(3550) <= not((inputs(242)) and (inputs(23)));
    layer0_outputs(3551) <= not((inputs(204)) xor (inputs(92)));
    layer0_outputs(3552) <= '0';
    layer0_outputs(3553) <= '0';
    layer0_outputs(3554) <= not((inputs(61)) xor (inputs(161)));
    layer0_outputs(3555) <= (inputs(152)) and not (inputs(58));
    layer0_outputs(3556) <= '0';
    layer0_outputs(3557) <= (inputs(75)) and not (inputs(24));
    layer0_outputs(3558) <= not((inputs(84)) and (inputs(253)));
    layer0_outputs(3559) <= (inputs(97)) or (inputs(74));
    layer0_outputs(3560) <= (inputs(156)) or (inputs(160));
    layer0_outputs(3561) <= '1';
    layer0_outputs(3562) <= not(inputs(221));
    layer0_outputs(3563) <= inputs(104);
    layer0_outputs(3564) <= inputs(172);
    layer0_outputs(3565) <= '1';
    layer0_outputs(3566) <= not(inputs(30)) or (inputs(250));
    layer0_outputs(3567) <= inputs(245);
    layer0_outputs(3568) <= (inputs(245)) and not (inputs(32));
    layer0_outputs(3569) <= (inputs(27)) and not (inputs(221));
    layer0_outputs(3570) <= '0';
    layer0_outputs(3571) <= not(inputs(217));
    layer0_outputs(3572) <= not(inputs(129));
    layer0_outputs(3573) <= (inputs(245)) and not (inputs(182));
    layer0_outputs(3574) <= (inputs(119)) or (inputs(242));
    layer0_outputs(3575) <= (inputs(53)) or (inputs(112));
    layer0_outputs(3576) <= not(inputs(65)) or (inputs(177));
    layer0_outputs(3577) <= (inputs(115)) and not (inputs(217));
    layer0_outputs(3578) <= inputs(17);
    layer0_outputs(3579) <= inputs(247);
    layer0_outputs(3580) <= (inputs(202)) or (inputs(19));
    layer0_outputs(3581) <= (inputs(177)) xor (inputs(144));
    layer0_outputs(3582) <= '0';
    layer0_outputs(3583) <= inputs(158);
    layer0_outputs(3584) <= '0';
    layer0_outputs(3585) <= '0';
    layer0_outputs(3586) <= (inputs(157)) and (inputs(247));
    layer0_outputs(3587) <= not(inputs(215)) or (inputs(219));
    layer0_outputs(3588) <= not((inputs(78)) or (inputs(122)));
    layer0_outputs(3589) <= '0';
    layer0_outputs(3590) <= '1';
    layer0_outputs(3591) <= inputs(163);
    layer0_outputs(3592) <= not((inputs(58)) or (inputs(0)));
    layer0_outputs(3593) <= not((inputs(170)) or (inputs(79)));
    layer0_outputs(3594) <= '0';
    layer0_outputs(3595) <= (inputs(230)) or (inputs(128));
    layer0_outputs(3596) <= '1';
    layer0_outputs(3597) <= '0';
    layer0_outputs(3598) <= (inputs(118)) xor (inputs(176));
    layer0_outputs(3599) <= inputs(232);
    layer0_outputs(3600) <= not(inputs(253));
    layer0_outputs(3601) <= (inputs(167)) and (inputs(179));
    layer0_outputs(3602) <= (inputs(153)) and (inputs(63));
    layer0_outputs(3603) <= '1';
    layer0_outputs(3604) <= (inputs(239)) xor (inputs(121));
    layer0_outputs(3605) <= not(inputs(109)) or (inputs(16));
    layer0_outputs(3606) <= not((inputs(128)) xor (inputs(167)));
    layer0_outputs(3607) <= inputs(168);
    layer0_outputs(3608) <= '1';
    layer0_outputs(3609) <= (inputs(148)) and not (inputs(206));
    layer0_outputs(3610) <= inputs(126);
    layer0_outputs(3611) <= not((inputs(217)) and (inputs(220)));
    layer0_outputs(3612) <= (inputs(169)) xor (inputs(118));
    layer0_outputs(3613) <= not(inputs(216));
    layer0_outputs(3614) <= not((inputs(155)) and (inputs(231)));
    layer0_outputs(3615) <= not((inputs(236)) and (inputs(134)));
    layer0_outputs(3616) <= not(inputs(247));
    layer0_outputs(3617) <= '0';
    layer0_outputs(3618) <= not(inputs(241));
    layer0_outputs(3619) <= not(inputs(247));
    layer0_outputs(3620) <= '0';
    layer0_outputs(3621) <= (inputs(21)) and (inputs(137));
    layer0_outputs(3622) <= inputs(190);
    layer0_outputs(3623) <= (inputs(142)) or (inputs(154));
    layer0_outputs(3624) <= inputs(33);
    layer0_outputs(3625) <= not((inputs(247)) or (inputs(175)));
    layer0_outputs(3626) <= (inputs(158)) and (inputs(139));
    layer0_outputs(3627) <= '0';
    layer0_outputs(3628) <= (inputs(184)) or (inputs(144));
    layer0_outputs(3629) <= not(inputs(151));
    layer0_outputs(3630) <= inputs(151);
    layer0_outputs(3631) <= '0';
    layer0_outputs(3632) <= '1';
    layer0_outputs(3633) <= not(inputs(92)) or (inputs(213));
    layer0_outputs(3634) <= not((inputs(222)) or (inputs(91)));
    layer0_outputs(3635) <= '1';
    layer0_outputs(3636) <= (inputs(220)) and (inputs(82));
    layer0_outputs(3637) <= not(inputs(183));
    layer0_outputs(3638) <= inputs(189);
    layer0_outputs(3639) <= (inputs(78)) or (inputs(21));
    layer0_outputs(3640) <= not(inputs(229));
    layer0_outputs(3641) <= not((inputs(195)) or (inputs(197)));
    layer0_outputs(3642) <= inputs(166);
    layer0_outputs(3643) <= not(inputs(232)) or (inputs(10));
    layer0_outputs(3644) <= '0';
    layer0_outputs(3645) <= not(inputs(205));
    layer0_outputs(3646) <= inputs(197);
    layer0_outputs(3647) <= inputs(116);
    layer0_outputs(3648) <= inputs(245);
    layer0_outputs(3649) <= (inputs(123)) or (inputs(102));
    layer0_outputs(3650) <= not(inputs(204)) or (inputs(248));
    layer0_outputs(3651) <= (inputs(187)) and not (inputs(255));
    layer0_outputs(3652) <= not(inputs(91));
    layer0_outputs(3653) <= (inputs(241)) xor (inputs(61));
    layer0_outputs(3654) <= '1';
    layer0_outputs(3655) <= not((inputs(90)) and (inputs(234)));
    layer0_outputs(3656) <= '1';
    layer0_outputs(3657) <= not(inputs(116));
    layer0_outputs(3658) <= not((inputs(169)) or (inputs(74)));
    layer0_outputs(3659) <= inputs(108);
    layer0_outputs(3660) <= '0';
    layer0_outputs(3661) <= inputs(85);
    layer0_outputs(3662) <= inputs(182);
    layer0_outputs(3663) <= inputs(2);
    layer0_outputs(3664) <= (inputs(125)) and not (inputs(240));
    layer0_outputs(3665) <= (inputs(93)) or (inputs(138));
    layer0_outputs(3666) <= '1';
    layer0_outputs(3667) <= not((inputs(92)) and (inputs(121)));
    layer0_outputs(3668) <= not(inputs(156)) or (inputs(149));
    layer0_outputs(3669) <= inputs(219);
    layer0_outputs(3670) <= (inputs(173)) and (inputs(156));
    layer0_outputs(3671) <= not(inputs(18)) or (inputs(10));
    layer0_outputs(3672) <= '0';
    layer0_outputs(3673) <= (inputs(234)) and not (inputs(252));
    layer0_outputs(3674) <= inputs(104);
    layer0_outputs(3675) <= (inputs(169)) and not (inputs(6));
    layer0_outputs(3676) <= not(inputs(59));
    layer0_outputs(3677) <= not((inputs(212)) xor (inputs(12)));
    layer0_outputs(3678) <= inputs(127);
    layer0_outputs(3679) <= inputs(177);
    layer0_outputs(3680) <= not((inputs(35)) and (inputs(87)));
    layer0_outputs(3681) <= not(inputs(166));
    layer0_outputs(3682) <= not((inputs(184)) and (inputs(194)));
    layer0_outputs(3683) <= '0';
    layer0_outputs(3684) <= (inputs(131)) and not (inputs(212));
    layer0_outputs(3685) <= not((inputs(15)) or (inputs(209)));
    layer0_outputs(3686) <= '1';
    layer0_outputs(3687) <= not(inputs(106)) or (inputs(130));
    layer0_outputs(3688) <= not((inputs(223)) xor (inputs(116)));
    layer0_outputs(3689) <= inputs(228);
    layer0_outputs(3690) <= not((inputs(126)) or (inputs(77)));
    layer0_outputs(3691) <= '1';
    layer0_outputs(3692) <= not((inputs(196)) or (inputs(209)));
    layer0_outputs(3693) <= (inputs(196)) or (inputs(245));
    layer0_outputs(3694) <= inputs(212);
    layer0_outputs(3695) <= (inputs(229)) and not (inputs(240));
    layer0_outputs(3696) <= inputs(127);
    layer0_outputs(3697) <= not(inputs(0)) or (inputs(31));
    layer0_outputs(3698) <= '0';
    layer0_outputs(3699) <= '0';
    layer0_outputs(3700) <= not(inputs(217)) or (inputs(208));
    layer0_outputs(3701) <= inputs(49);
    layer0_outputs(3702) <= (inputs(60)) and (inputs(110));
    layer0_outputs(3703) <= not((inputs(110)) and (inputs(68)));
    layer0_outputs(3704) <= inputs(194);
    layer0_outputs(3705) <= not(inputs(166));
    layer0_outputs(3706) <= inputs(193);
    layer0_outputs(3707) <= not((inputs(169)) and (inputs(38)));
    layer0_outputs(3708) <= (inputs(41)) and not (inputs(183));
    layer0_outputs(3709) <= not(inputs(113)) or (inputs(92));
    layer0_outputs(3710) <= not(inputs(226)) or (inputs(63));
    layer0_outputs(3711) <= '0';
    layer0_outputs(3712) <= '0';
    layer0_outputs(3713) <= not(inputs(162)) or (inputs(222));
    layer0_outputs(3714) <= not((inputs(34)) or (inputs(160)));
    layer0_outputs(3715) <= not((inputs(208)) or (inputs(184)));
    layer0_outputs(3716) <= (inputs(173)) or (inputs(123));
    layer0_outputs(3717) <= (inputs(96)) and not (inputs(34));
    layer0_outputs(3718) <= (inputs(103)) and not (inputs(161));
    layer0_outputs(3719) <= not((inputs(71)) or (inputs(170)));
    layer0_outputs(3720) <= not(inputs(225)) or (inputs(30));
    layer0_outputs(3721) <= not(inputs(163));
    layer0_outputs(3722) <= (inputs(192)) and (inputs(242));
    layer0_outputs(3723) <= not(inputs(226)) or (inputs(40));
    layer0_outputs(3724) <= '1';
    layer0_outputs(3725) <= '1';
    layer0_outputs(3726) <= inputs(230);
    layer0_outputs(3727) <= not((inputs(151)) and (inputs(158)));
    layer0_outputs(3728) <= inputs(126);
    layer0_outputs(3729) <= inputs(230);
    layer0_outputs(3730) <= not((inputs(108)) or (inputs(172)));
    layer0_outputs(3731) <= (inputs(231)) and not (inputs(238));
    layer0_outputs(3732) <= not(inputs(83));
    layer0_outputs(3733) <= '1';
    layer0_outputs(3734) <= not((inputs(67)) and (inputs(125)));
    layer0_outputs(3735) <= not(inputs(209));
    layer0_outputs(3736) <= not(inputs(37));
    layer0_outputs(3737) <= not(inputs(79)) or (inputs(232));
    layer0_outputs(3738) <= not((inputs(158)) or (inputs(242)));
    layer0_outputs(3739) <= not((inputs(185)) or (inputs(18)));
    layer0_outputs(3740) <= '0';
    layer0_outputs(3741) <= inputs(141);
    layer0_outputs(3742) <= not((inputs(197)) or (inputs(197)));
    layer0_outputs(3743) <= (inputs(240)) xor (inputs(179));
    layer0_outputs(3744) <= inputs(177);
    layer0_outputs(3745) <= not((inputs(145)) and (inputs(55)));
    layer0_outputs(3746) <= not(inputs(68)) or (inputs(142));
    layer0_outputs(3747) <= '1';
    layer0_outputs(3748) <= '1';
    layer0_outputs(3749) <= inputs(216);
    layer0_outputs(3750) <= inputs(103);
    layer0_outputs(3751) <= (inputs(222)) and (inputs(43));
    layer0_outputs(3752) <= not(inputs(165));
    layer0_outputs(3753) <= (inputs(47)) or (inputs(14));
    layer0_outputs(3754) <= '0';
    layer0_outputs(3755) <= inputs(119);
    layer0_outputs(3756) <= not(inputs(114)) or (inputs(152));
    layer0_outputs(3757) <= not((inputs(214)) xor (inputs(238)));
    layer0_outputs(3758) <= (inputs(158)) or (inputs(186));
    layer0_outputs(3759) <= not(inputs(211)) or (inputs(13));
    layer0_outputs(3760) <= not((inputs(240)) and (inputs(119)));
    layer0_outputs(3761) <= inputs(134);
    layer0_outputs(3762) <= (inputs(90)) and not (inputs(189));
    layer0_outputs(3763) <= '1';
    layer0_outputs(3764) <= inputs(165);
    layer0_outputs(3765) <= not(inputs(68)) or (inputs(200));
    layer0_outputs(3766) <= inputs(214);
    layer0_outputs(3767) <= not(inputs(229)) or (inputs(166));
    layer0_outputs(3768) <= (inputs(157)) and not (inputs(56));
    layer0_outputs(3769) <= (inputs(130)) and not (inputs(188));
    layer0_outputs(3770) <= inputs(160);
    layer0_outputs(3771) <= inputs(20);
    layer0_outputs(3772) <= (inputs(190)) and not (inputs(12));
    layer0_outputs(3773) <= inputs(65);
    layer0_outputs(3774) <= not(inputs(4));
    layer0_outputs(3775) <= not((inputs(34)) xor (inputs(11)));
    layer0_outputs(3776) <= '0';
    layer0_outputs(3777) <= '0';
    layer0_outputs(3778) <= (inputs(4)) and not (inputs(127));
    layer0_outputs(3779) <= (inputs(159)) or (inputs(9));
    layer0_outputs(3780) <= '0';
    layer0_outputs(3781) <= not(inputs(44));
    layer0_outputs(3782) <= not((inputs(83)) or (inputs(182)));
    layer0_outputs(3783) <= not(inputs(204));
    layer0_outputs(3784) <= not(inputs(226));
    layer0_outputs(3785) <= not(inputs(135));
    layer0_outputs(3786) <= (inputs(194)) and (inputs(114));
    layer0_outputs(3787) <= (inputs(220)) xor (inputs(66));
    layer0_outputs(3788) <= (inputs(49)) or (inputs(64));
    layer0_outputs(3789) <= not(inputs(173)) or (inputs(166));
    layer0_outputs(3790) <= inputs(218);
    layer0_outputs(3791) <= not((inputs(18)) or (inputs(125)));
    layer0_outputs(3792) <= not(inputs(120));
    layer0_outputs(3793) <= (inputs(38)) and not (inputs(108));
    layer0_outputs(3794) <= (inputs(198)) xor (inputs(119));
    layer0_outputs(3795) <= '1';
    layer0_outputs(3796) <= not(inputs(104)) or (inputs(5));
    layer0_outputs(3797) <= inputs(130);
    layer0_outputs(3798) <= not(inputs(233));
    layer0_outputs(3799) <= (inputs(51)) and not (inputs(245));
    layer0_outputs(3800) <= not((inputs(155)) and (inputs(215)));
    layer0_outputs(3801) <= '1';
    layer0_outputs(3802) <= (inputs(104)) or (inputs(11));
    layer0_outputs(3803) <= (inputs(240)) xor (inputs(109));
    layer0_outputs(3804) <= not((inputs(112)) or (inputs(203)));
    layer0_outputs(3805) <= not((inputs(114)) or (inputs(217)));
    layer0_outputs(3806) <= not((inputs(215)) or (inputs(194)));
    layer0_outputs(3807) <= '0';
    layer0_outputs(3808) <= not(inputs(85)) or (inputs(178));
    layer0_outputs(3809) <= not(inputs(143));
    layer0_outputs(3810) <= (inputs(94)) or (inputs(239));
    layer0_outputs(3811) <= '0';
    layer0_outputs(3812) <= not(inputs(127));
    layer0_outputs(3813) <= '1';
    layer0_outputs(3814) <= inputs(94);
    layer0_outputs(3815) <= not(inputs(153));
    layer0_outputs(3816) <= not(inputs(219));
    layer0_outputs(3817) <= (inputs(16)) xor (inputs(252));
    layer0_outputs(3818) <= '1';
    layer0_outputs(3819) <= inputs(49);
    layer0_outputs(3820) <= '0';
    layer0_outputs(3821) <= (inputs(69)) and (inputs(152));
    layer0_outputs(3822) <= not(inputs(186));
    layer0_outputs(3823) <= (inputs(81)) and not (inputs(83));
    layer0_outputs(3824) <= not(inputs(51));
    layer0_outputs(3825) <= (inputs(8)) or (inputs(175));
    layer0_outputs(3826) <= not(inputs(144)) or (inputs(53));
    layer0_outputs(3827) <= (inputs(0)) and (inputs(111));
    layer0_outputs(3828) <= '1';
    layer0_outputs(3829) <= inputs(170);
    layer0_outputs(3830) <= not(inputs(50));
    layer0_outputs(3831) <= '0';
    layer0_outputs(3832) <= inputs(88);
    layer0_outputs(3833) <= (inputs(100)) xor (inputs(56));
    layer0_outputs(3834) <= not(inputs(10)) or (inputs(162));
    layer0_outputs(3835) <= not(inputs(122));
    layer0_outputs(3836) <= inputs(84);
    layer0_outputs(3837) <= not((inputs(201)) and (inputs(139)));
    layer0_outputs(3838) <= inputs(52);
    layer0_outputs(3839) <= (inputs(101)) and (inputs(7));
    layer0_outputs(3840) <= '0';
    layer0_outputs(3841) <= (inputs(100)) or (inputs(165));
    layer0_outputs(3842) <= (inputs(106)) and not (inputs(208));
    layer0_outputs(3843) <= not((inputs(224)) or (inputs(50)));
    layer0_outputs(3844) <= inputs(156);
    layer0_outputs(3845) <= not((inputs(11)) and (inputs(38)));
    layer0_outputs(3846) <= inputs(21);
    layer0_outputs(3847) <= inputs(219);
    layer0_outputs(3848) <= '1';
    layer0_outputs(3849) <= not((inputs(78)) and (inputs(175)));
    layer0_outputs(3850) <= '1';
    layer0_outputs(3851) <= '0';
    layer0_outputs(3852) <= not((inputs(78)) xor (inputs(129)));
    layer0_outputs(3853) <= not(inputs(9)) or (inputs(1));
    layer0_outputs(3854) <= inputs(164);
    layer0_outputs(3855) <= not(inputs(14));
    layer0_outputs(3856) <= inputs(37);
    layer0_outputs(3857) <= not(inputs(248));
    layer0_outputs(3858) <= (inputs(199)) and not (inputs(55));
    layer0_outputs(3859) <= inputs(211);
    layer0_outputs(3860) <= (inputs(15)) and not (inputs(137));
    layer0_outputs(3861) <= (inputs(65)) and (inputs(185));
    layer0_outputs(3862) <= (inputs(76)) and (inputs(160));
    layer0_outputs(3863) <= not(inputs(234));
    layer0_outputs(3864) <= not(inputs(113));
    layer0_outputs(3865) <= inputs(162);
    layer0_outputs(3866) <= (inputs(174)) and not (inputs(223));
    layer0_outputs(3867) <= not(inputs(153));
    layer0_outputs(3868) <= (inputs(15)) and (inputs(199));
    layer0_outputs(3869) <= '0';
    layer0_outputs(3870) <= not(inputs(15));
    layer0_outputs(3871) <= (inputs(167)) and not (inputs(132));
    layer0_outputs(3872) <= not(inputs(27));
    layer0_outputs(3873) <= not((inputs(93)) xor (inputs(63)));
    layer0_outputs(3874) <= (inputs(50)) and not (inputs(40));
    layer0_outputs(3875) <= '1';
    layer0_outputs(3876) <= (inputs(24)) and (inputs(98));
    layer0_outputs(3877) <= (inputs(58)) or (inputs(126));
    layer0_outputs(3878) <= (inputs(234)) and not (inputs(54));
    layer0_outputs(3879) <= not(inputs(65));
    layer0_outputs(3880) <= '1';
    layer0_outputs(3881) <= not(inputs(37)) or (inputs(209));
    layer0_outputs(3882) <= not(inputs(182));
    layer0_outputs(3883) <= (inputs(242)) and not (inputs(228));
    layer0_outputs(3884) <= inputs(222);
    layer0_outputs(3885) <= not(inputs(182));
    layer0_outputs(3886) <= (inputs(37)) xor (inputs(18));
    layer0_outputs(3887) <= inputs(24);
    layer0_outputs(3888) <= not(inputs(178)) or (inputs(105));
    layer0_outputs(3889) <= not(inputs(100));
    layer0_outputs(3890) <= not((inputs(242)) and (inputs(40)));
    layer0_outputs(3891) <= (inputs(231)) or (inputs(16));
    layer0_outputs(3892) <= not((inputs(21)) or (inputs(233)));
    layer0_outputs(3893) <= not(inputs(29));
    layer0_outputs(3894) <= not((inputs(40)) xor (inputs(95)));
    layer0_outputs(3895) <= (inputs(157)) and not (inputs(173));
    layer0_outputs(3896) <= (inputs(53)) and not (inputs(175));
    layer0_outputs(3897) <= not(inputs(74)) or (inputs(164));
    layer0_outputs(3898) <= not((inputs(219)) and (inputs(162)));
    layer0_outputs(3899) <= not(inputs(122)) or (inputs(32));
    layer0_outputs(3900) <= '0';
    layer0_outputs(3901) <= '1';
    layer0_outputs(3902) <= not(inputs(86));
    layer0_outputs(3903) <= '1';
    layer0_outputs(3904) <= not(inputs(160));
    layer0_outputs(3905) <= (inputs(81)) or (inputs(253));
    layer0_outputs(3906) <= not(inputs(70));
    layer0_outputs(3907) <= '0';
    layer0_outputs(3908) <= not(inputs(17)) or (inputs(75));
    layer0_outputs(3909) <= not(inputs(124)) or (inputs(81));
    layer0_outputs(3910) <= inputs(128);
    layer0_outputs(3911) <= not(inputs(134));
    layer0_outputs(3912) <= (inputs(123)) or (inputs(105));
    layer0_outputs(3913) <= '0';
    layer0_outputs(3914) <= inputs(240);
    layer0_outputs(3915) <= (inputs(243)) or (inputs(217));
    layer0_outputs(3916) <= (inputs(49)) and (inputs(13));
    layer0_outputs(3917) <= not((inputs(29)) or (inputs(67)));
    layer0_outputs(3918) <= not(inputs(201)) or (inputs(193));
    layer0_outputs(3919) <= not((inputs(60)) and (inputs(193)));
    layer0_outputs(3920) <= not(inputs(153)) or (inputs(43));
    layer0_outputs(3921) <= (inputs(181)) and not (inputs(182));
    layer0_outputs(3922) <= (inputs(156)) or (inputs(129));
    layer0_outputs(3923) <= not(inputs(176));
    layer0_outputs(3924) <= (inputs(72)) and not (inputs(221));
    layer0_outputs(3925) <= '0';
    layer0_outputs(3926) <= not(inputs(114)) or (inputs(37));
    layer0_outputs(3927) <= not(inputs(24)) or (inputs(120));
    layer0_outputs(3928) <= (inputs(30)) xor (inputs(20));
    layer0_outputs(3929) <= not(inputs(188)) or (inputs(217));
    layer0_outputs(3930) <= not(inputs(18));
    layer0_outputs(3931) <= not(inputs(50));
    layer0_outputs(3932) <= not((inputs(220)) or (inputs(172)));
    layer0_outputs(3933) <= '1';
    layer0_outputs(3934) <= not(inputs(160)) or (inputs(171));
    layer0_outputs(3935) <= not((inputs(117)) and (inputs(254)));
    layer0_outputs(3936) <= not((inputs(214)) and (inputs(237)));
    layer0_outputs(3937) <= not(inputs(92));
    layer0_outputs(3938) <= not((inputs(3)) or (inputs(228)));
    layer0_outputs(3939) <= inputs(25);
    layer0_outputs(3940) <= (inputs(132)) and not (inputs(223));
    layer0_outputs(3941) <= not((inputs(186)) or (inputs(81)));
    layer0_outputs(3942) <= not((inputs(79)) or (inputs(247)));
    layer0_outputs(3943) <= '0';
    layer0_outputs(3944) <= '1';
    layer0_outputs(3945) <= not(inputs(225));
    layer0_outputs(3946) <= not(inputs(239));
    layer0_outputs(3947) <= not((inputs(29)) or (inputs(77)));
    layer0_outputs(3948) <= '0';
    layer0_outputs(3949) <= (inputs(14)) and not (inputs(174));
    layer0_outputs(3950) <= '1';
    layer0_outputs(3951) <= not(inputs(232)) or (inputs(109));
    layer0_outputs(3952) <= not(inputs(243));
    layer0_outputs(3953) <= not(inputs(48));
    layer0_outputs(3954) <= '0';
    layer0_outputs(3955) <= (inputs(151)) and not (inputs(206));
    layer0_outputs(3956) <= not((inputs(14)) and (inputs(86)));
    layer0_outputs(3957) <= not((inputs(15)) or (inputs(35)));
    layer0_outputs(3958) <= not((inputs(34)) and (inputs(30)));
    layer0_outputs(3959) <= '0';
    layer0_outputs(3960) <= (inputs(61)) and not (inputs(73));
    layer0_outputs(3961) <= '1';
    layer0_outputs(3962) <= (inputs(177)) xor (inputs(132));
    layer0_outputs(3963) <= not((inputs(218)) or (inputs(227)));
    layer0_outputs(3964) <= not((inputs(80)) xor (inputs(20)));
    layer0_outputs(3965) <= not(inputs(143));
    layer0_outputs(3966) <= inputs(196);
    layer0_outputs(3967) <= (inputs(2)) or (inputs(93));
    layer0_outputs(3968) <= (inputs(120)) and not (inputs(139));
    layer0_outputs(3969) <= (inputs(21)) and not (inputs(223));
    layer0_outputs(3970) <= not((inputs(88)) or (inputs(28)));
    layer0_outputs(3971) <= (inputs(52)) xor (inputs(4));
    layer0_outputs(3972) <= inputs(172);
    layer0_outputs(3973) <= not((inputs(25)) or (inputs(102)));
    layer0_outputs(3974) <= (inputs(26)) and (inputs(50));
    layer0_outputs(3975) <= not(inputs(59));
    layer0_outputs(3976) <= (inputs(41)) and (inputs(162));
    layer0_outputs(3977) <= (inputs(128)) and (inputs(67));
    layer0_outputs(3978) <= not((inputs(27)) or (inputs(115)));
    layer0_outputs(3979) <= (inputs(102)) and (inputs(74));
    layer0_outputs(3980) <= not((inputs(0)) or (inputs(48)));
    layer0_outputs(3981) <= not((inputs(221)) or (inputs(188)));
    layer0_outputs(3982) <= inputs(196);
    layer0_outputs(3983) <= (inputs(223)) xor (inputs(148));
    layer0_outputs(3984) <= (inputs(14)) and (inputs(77));
    layer0_outputs(3985) <= '0';
    layer0_outputs(3986) <= '1';
    layer0_outputs(3987) <= (inputs(99)) or (inputs(115));
    layer0_outputs(3988) <= not((inputs(237)) and (inputs(107)));
    layer0_outputs(3989) <= inputs(62);
    layer0_outputs(3990) <= not((inputs(237)) or (inputs(251)));
    layer0_outputs(3991) <= '0';
    layer0_outputs(3992) <= inputs(178);
    layer0_outputs(3993) <= (inputs(226)) and (inputs(236));
    layer0_outputs(3994) <= not(inputs(146));
    layer0_outputs(3995) <= (inputs(173)) or (inputs(1));
    layer0_outputs(3996) <= '0';
    layer0_outputs(3997) <= not((inputs(187)) or (inputs(50)));
    layer0_outputs(3998) <= (inputs(168)) and not (inputs(207));
    layer0_outputs(3999) <= (inputs(177)) and not (inputs(173));
    layer0_outputs(4000) <= '0';
    layer0_outputs(4001) <= (inputs(205)) and not (inputs(141));
    layer0_outputs(4002) <= '0';
    layer0_outputs(4003) <= '0';
    layer0_outputs(4004) <= inputs(108);
    layer0_outputs(4005) <= inputs(52);
    layer0_outputs(4006) <= not(inputs(117));
    layer0_outputs(4007) <= '0';
    layer0_outputs(4008) <= not(inputs(178));
    layer0_outputs(4009) <= not((inputs(76)) and (inputs(11)));
    layer0_outputs(4010) <= (inputs(179)) and (inputs(245));
    layer0_outputs(4011) <= not(inputs(50)) or (inputs(182));
    layer0_outputs(4012) <= inputs(104);
    layer0_outputs(4013) <= not((inputs(211)) and (inputs(37)));
    layer0_outputs(4014) <= (inputs(1)) or (inputs(140));
    layer0_outputs(4015) <= '0';
    layer0_outputs(4016) <= inputs(191);
    layer0_outputs(4017) <= '0';
    layer0_outputs(4018) <= not(inputs(167)) or (inputs(10));
    layer0_outputs(4019) <= not(inputs(168));
    layer0_outputs(4020) <= not(inputs(18));
    layer0_outputs(4021) <= (inputs(248)) and not (inputs(46));
    layer0_outputs(4022) <= (inputs(185)) and (inputs(54));
    layer0_outputs(4023) <= (inputs(9)) and (inputs(126));
    layer0_outputs(4024) <= not(inputs(199));
    layer0_outputs(4025) <= inputs(128);
    layer0_outputs(4026) <= '1';
    layer0_outputs(4027) <= '1';
    layer0_outputs(4028) <= not(inputs(97)) or (inputs(13));
    layer0_outputs(4029) <= '1';
    layer0_outputs(4030) <= (inputs(48)) or (inputs(253));
    layer0_outputs(4031) <= '1';
    layer0_outputs(4032) <= not((inputs(191)) or (inputs(182)));
    layer0_outputs(4033) <= (inputs(141)) and not (inputs(21));
    layer0_outputs(4034) <= not(inputs(55)) or (inputs(150));
    layer0_outputs(4035) <= inputs(121);
    layer0_outputs(4036) <= inputs(103);
    layer0_outputs(4037) <= not((inputs(76)) xor (inputs(1)));
    layer0_outputs(4038) <= inputs(141);
    layer0_outputs(4039) <= not(inputs(218)) or (inputs(99));
    layer0_outputs(4040) <= not((inputs(158)) or (inputs(131)));
    layer0_outputs(4041) <= not(inputs(205));
    layer0_outputs(4042) <= (inputs(12)) and (inputs(30));
    layer0_outputs(4043) <= inputs(35);
    layer0_outputs(4044) <= (inputs(82)) and not (inputs(216));
    layer0_outputs(4045) <= (inputs(132)) or (inputs(27));
    layer0_outputs(4046) <= inputs(99);
    layer0_outputs(4047) <= '1';
    layer0_outputs(4048) <= '0';
    layer0_outputs(4049) <= (inputs(75)) xor (inputs(17));
    layer0_outputs(4050) <= (inputs(109)) and (inputs(251));
    layer0_outputs(4051) <= '1';
    layer0_outputs(4052) <= (inputs(253)) or (inputs(122));
    layer0_outputs(4053) <= not(inputs(254));
    layer0_outputs(4054) <= '1';
    layer0_outputs(4055) <= not(inputs(66)) or (inputs(159));
    layer0_outputs(4056) <= not(inputs(236)) or (inputs(7));
    layer0_outputs(4057) <= inputs(68);
    layer0_outputs(4058) <= (inputs(8)) or (inputs(122));
    layer0_outputs(4059) <= (inputs(233)) or (inputs(224));
    layer0_outputs(4060) <= not(inputs(122));
    layer0_outputs(4061) <= not(inputs(143));
    layer0_outputs(4062) <= inputs(148);
    layer0_outputs(4063) <= inputs(201);
    layer0_outputs(4064) <= (inputs(31)) and (inputs(178));
    layer0_outputs(4065) <= inputs(128);
    layer0_outputs(4066) <= inputs(38);
    layer0_outputs(4067) <= not(inputs(168)) or (inputs(111));
    layer0_outputs(4068) <= (inputs(75)) and not (inputs(177));
    layer0_outputs(4069) <= not((inputs(213)) and (inputs(34)));
    layer0_outputs(4070) <= not(inputs(151)) or (inputs(207));
    layer0_outputs(4071) <= not((inputs(89)) or (inputs(42)));
    layer0_outputs(4072) <= (inputs(138)) xor (inputs(191));
    layer0_outputs(4073) <= not(inputs(206)) or (inputs(164));
    layer0_outputs(4074) <= not(inputs(165)) or (inputs(107));
    layer0_outputs(4075) <= not(inputs(32));
    layer0_outputs(4076) <= '1';
    layer0_outputs(4077) <= (inputs(117)) and not (inputs(43));
    layer0_outputs(4078) <= inputs(199);
    layer0_outputs(4079) <= '1';
    layer0_outputs(4080) <= (inputs(213)) and not (inputs(108));
    layer0_outputs(4081) <= not(inputs(174)) or (inputs(170));
    layer0_outputs(4082) <= inputs(63);
    layer0_outputs(4083) <= inputs(141);
    layer0_outputs(4084) <= not(inputs(140));
    layer0_outputs(4085) <= not((inputs(136)) and (inputs(18)));
    layer0_outputs(4086) <= not(inputs(224)) or (inputs(216));
    layer0_outputs(4087) <= '1';
    layer0_outputs(4088) <= '1';
    layer0_outputs(4089) <= '0';
    layer0_outputs(4090) <= (inputs(66)) or (inputs(129));
    layer0_outputs(4091) <= not(inputs(47)) or (inputs(121));
    layer0_outputs(4092) <= not(inputs(134));
    layer0_outputs(4093) <= (inputs(205)) or (inputs(146));
    layer0_outputs(4094) <= not((inputs(226)) or (inputs(89)));
    layer0_outputs(4095) <= not(inputs(25));
    layer0_outputs(4096) <= inputs(165);
    layer0_outputs(4097) <= not(inputs(162)) or (inputs(146));
    layer0_outputs(4098) <= '1';
    layer0_outputs(4099) <= '0';
    layer0_outputs(4100) <= '0';
    layer0_outputs(4101) <= (inputs(176)) and not (inputs(39));
    layer0_outputs(4102) <= not(inputs(55)) or (inputs(63));
    layer0_outputs(4103) <= not(inputs(165)) or (inputs(46));
    layer0_outputs(4104) <= not(inputs(4));
    layer0_outputs(4105) <= inputs(210);
    layer0_outputs(4106) <= not((inputs(138)) and (inputs(237)));
    layer0_outputs(4107) <= inputs(148);
    layer0_outputs(4108) <= inputs(189);
    layer0_outputs(4109) <= not(inputs(26));
    layer0_outputs(4110) <= (inputs(211)) and not (inputs(182));
    layer0_outputs(4111) <= not(inputs(234));
    layer0_outputs(4112) <= not(inputs(97));
    layer0_outputs(4113) <= (inputs(107)) or (inputs(59));
    layer0_outputs(4114) <= not(inputs(169));
    layer0_outputs(4115) <= inputs(90);
    layer0_outputs(4116) <= not(inputs(48));
    layer0_outputs(4117) <= '1';
    layer0_outputs(4118) <= '0';
    layer0_outputs(4119) <= inputs(249);
    layer0_outputs(4120) <= not(inputs(133)) or (inputs(121));
    layer0_outputs(4121) <= (inputs(127)) and not (inputs(56));
    layer0_outputs(4122) <= '0';
    layer0_outputs(4123) <= not(inputs(141));
    layer0_outputs(4124) <= (inputs(174)) and not (inputs(17));
    layer0_outputs(4125) <= (inputs(58)) and not (inputs(183));
    layer0_outputs(4126) <= not((inputs(227)) or (inputs(181)));
    layer0_outputs(4127) <= not(inputs(228));
    layer0_outputs(4128) <= (inputs(125)) and not (inputs(217));
    layer0_outputs(4129) <= not(inputs(80));
    layer0_outputs(4130) <= (inputs(83)) or (inputs(49));
    layer0_outputs(4131) <= (inputs(33)) or (inputs(17));
    layer0_outputs(4132) <= (inputs(175)) xor (inputs(61));
    layer0_outputs(4133) <= '0';
    layer0_outputs(4134) <= (inputs(56)) and (inputs(154));
    layer0_outputs(4135) <= not(inputs(23));
    layer0_outputs(4136) <= not((inputs(192)) or (inputs(183)));
    layer0_outputs(4137) <= (inputs(71)) and not (inputs(90));
    layer0_outputs(4138) <= (inputs(140)) and (inputs(130));
    layer0_outputs(4139) <= inputs(79);
    layer0_outputs(4140) <= not((inputs(237)) xor (inputs(191)));
    layer0_outputs(4141) <= not(inputs(158));
    layer0_outputs(4142) <= (inputs(77)) or (inputs(0));
    layer0_outputs(4143) <= (inputs(99)) or (inputs(69));
    layer0_outputs(4144) <= not(inputs(76));
    layer0_outputs(4145) <= (inputs(96)) and not (inputs(218));
    layer0_outputs(4146) <= not((inputs(177)) or (inputs(208)));
    layer0_outputs(4147) <= inputs(84);
    layer0_outputs(4148) <= inputs(125);
    layer0_outputs(4149) <= not((inputs(75)) or (inputs(57)));
    layer0_outputs(4150) <= inputs(227);
    layer0_outputs(4151) <= '1';
    layer0_outputs(4152) <= (inputs(156)) or (inputs(2));
    layer0_outputs(4153) <= (inputs(174)) and not (inputs(222));
    layer0_outputs(4154) <= (inputs(74)) and not (inputs(247));
    layer0_outputs(4155) <= not(inputs(11)) or (inputs(150));
    layer0_outputs(4156) <= not(inputs(120));
    layer0_outputs(4157) <= '1';
    layer0_outputs(4158) <= inputs(252);
    layer0_outputs(4159) <= (inputs(194)) and not (inputs(118));
    layer0_outputs(4160) <= not(inputs(163));
    layer0_outputs(4161) <= '1';
    layer0_outputs(4162) <= not(inputs(17));
    layer0_outputs(4163) <= (inputs(161)) and not (inputs(128));
    layer0_outputs(4164) <= not((inputs(52)) or (inputs(54)));
    layer0_outputs(4165) <= '0';
    layer0_outputs(4166) <= not(inputs(24));
    layer0_outputs(4167) <= not(inputs(93));
    layer0_outputs(4168) <= not(inputs(57));
    layer0_outputs(4169) <= not(inputs(223));
    layer0_outputs(4170) <= (inputs(189)) and (inputs(35));
    layer0_outputs(4171) <= '0';
    layer0_outputs(4172) <= (inputs(15)) xor (inputs(152));
    layer0_outputs(4173) <= inputs(210);
    layer0_outputs(4174) <= inputs(100);
    layer0_outputs(4175) <= inputs(161);
    layer0_outputs(4176) <= inputs(55);
    layer0_outputs(4177) <= not(inputs(236)) or (inputs(114));
    layer0_outputs(4178) <= not(inputs(201)) or (inputs(131));
    layer0_outputs(4179) <= not(inputs(187)) or (inputs(145));
    layer0_outputs(4180) <= '0';
    layer0_outputs(4181) <= inputs(114);
    layer0_outputs(4182) <= (inputs(202)) and (inputs(202));
    layer0_outputs(4183) <= inputs(59);
    layer0_outputs(4184) <= not(inputs(180));
    layer0_outputs(4185) <= not((inputs(184)) xor (inputs(27)));
    layer0_outputs(4186) <= inputs(194);
    layer0_outputs(4187) <= not((inputs(95)) and (inputs(191)));
    layer0_outputs(4188) <= not(inputs(150));
    layer0_outputs(4189) <= (inputs(151)) and not (inputs(146));
    layer0_outputs(4190) <= '0';
    layer0_outputs(4191) <= not(inputs(72));
    layer0_outputs(4192) <= (inputs(85)) or (inputs(38));
    layer0_outputs(4193) <= '0';
    layer0_outputs(4194) <= not((inputs(67)) or (inputs(157)));
    layer0_outputs(4195) <= not((inputs(207)) or (inputs(51)));
    layer0_outputs(4196) <= inputs(238);
    layer0_outputs(4197) <= not(inputs(143)) or (inputs(93));
    layer0_outputs(4198) <= (inputs(160)) or (inputs(85));
    layer0_outputs(4199) <= inputs(253);
    layer0_outputs(4200) <= inputs(156);
    layer0_outputs(4201) <= (inputs(133)) and not (inputs(40));
    layer0_outputs(4202) <= not(inputs(172));
    layer0_outputs(4203) <= (inputs(159)) and (inputs(41));
    layer0_outputs(4204) <= inputs(248);
    layer0_outputs(4205) <= (inputs(77)) or (inputs(62));
    layer0_outputs(4206) <= not(inputs(127));
    layer0_outputs(4207) <= not((inputs(164)) or (inputs(160)));
    layer0_outputs(4208) <= not((inputs(244)) or (inputs(27)));
    layer0_outputs(4209) <= (inputs(87)) or (inputs(89));
    layer0_outputs(4210) <= inputs(222);
    layer0_outputs(4211) <= '1';
    layer0_outputs(4212) <= not(inputs(37)) or (inputs(141));
    layer0_outputs(4213) <= (inputs(104)) and not (inputs(189));
    layer0_outputs(4214) <= not(inputs(36));
    layer0_outputs(4215) <= not(inputs(155));
    layer0_outputs(4216) <= inputs(250);
    layer0_outputs(4217) <= not(inputs(110));
    layer0_outputs(4218) <= not(inputs(118));
    layer0_outputs(4219) <= not(inputs(46)) or (inputs(174));
    layer0_outputs(4220) <= not(inputs(93));
    layer0_outputs(4221) <= not(inputs(217)) or (inputs(27));
    layer0_outputs(4222) <= (inputs(135)) or (inputs(30));
    layer0_outputs(4223) <= '1';
    layer0_outputs(4224) <= not(inputs(148));
    layer0_outputs(4225) <= (inputs(130)) and not (inputs(54));
    layer0_outputs(4226) <= (inputs(231)) and not (inputs(238));
    layer0_outputs(4227) <= inputs(72);
    layer0_outputs(4228) <= (inputs(190)) or (inputs(195));
    layer0_outputs(4229) <= '1';
    layer0_outputs(4230) <= '0';
    layer0_outputs(4231) <= (inputs(119)) and not (inputs(156));
    layer0_outputs(4232) <= (inputs(240)) or (inputs(215));
    layer0_outputs(4233) <= '0';
    layer0_outputs(4234) <= (inputs(157)) and not (inputs(152));
    layer0_outputs(4235) <= '1';
    layer0_outputs(4236) <= not((inputs(198)) or (inputs(23)));
    layer0_outputs(4237) <= not((inputs(236)) and (inputs(65)));
    layer0_outputs(4238) <= not(inputs(97));
    layer0_outputs(4239) <= '0';
    layer0_outputs(4240) <= not(inputs(198)) or (inputs(144));
    layer0_outputs(4241) <= (inputs(247)) or (inputs(238));
    layer0_outputs(4242) <= not(inputs(75));
    layer0_outputs(4243) <= not((inputs(50)) or (inputs(248)));
    layer0_outputs(4244) <= not((inputs(179)) or (inputs(235)));
    layer0_outputs(4245) <= (inputs(120)) and not (inputs(230));
    layer0_outputs(4246) <= not((inputs(109)) or (inputs(219)));
    layer0_outputs(4247) <= not(inputs(136)) or (inputs(219));
    layer0_outputs(4248) <= (inputs(107)) and not (inputs(79));
    layer0_outputs(4249) <= (inputs(38)) or (inputs(60));
    layer0_outputs(4250) <= (inputs(34)) xor (inputs(140));
    layer0_outputs(4251) <= not(inputs(46)) or (inputs(17));
    layer0_outputs(4252) <= inputs(113);
    layer0_outputs(4253) <= '0';
    layer0_outputs(4254) <= (inputs(159)) xor (inputs(1));
    layer0_outputs(4255) <= not((inputs(181)) or (inputs(161)));
    layer0_outputs(4256) <= '1';
    layer0_outputs(4257) <= (inputs(137)) and not (inputs(172));
    layer0_outputs(4258) <= not(inputs(198));
    layer0_outputs(4259) <= (inputs(155)) or (inputs(50));
    layer0_outputs(4260) <= not((inputs(47)) and (inputs(185)));
    layer0_outputs(4261) <= (inputs(126)) and not (inputs(217));
    layer0_outputs(4262) <= '1';
    layer0_outputs(4263) <= (inputs(103)) or (inputs(120));
    layer0_outputs(4264) <= (inputs(91)) xor (inputs(66));
    layer0_outputs(4265) <= not(inputs(182));
    layer0_outputs(4266) <= (inputs(227)) or (inputs(241));
    layer0_outputs(4267) <= '0';
    layer0_outputs(4268) <= not(inputs(68));
    layer0_outputs(4269) <= not(inputs(82));
    layer0_outputs(4270) <= inputs(125);
    layer0_outputs(4271) <= (inputs(98)) and not (inputs(228));
    layer0_outputs(4272) <= '1';
    layer0_outputs(4273) <= not((inputs(106)) and (inputs(127)));
    layer0_outputs(4274) <= '0';
    layer0_outputs(4275) <= not(inputs(167)) or (inputs(127));
    layer0_outputs(4276) <= (inputs(19)) and not (inputs(245));
    layer0_outputs(4277) <= inputs(246);
    layer0_outputs(4278) <= not(inputs(99)) or (inputs(47));
    layer0_outputs(4279) <= not(inputs(139));
    layer0_outputs(4280) <= not((inputs(22)) or (inputs(156)));
    layer0_outputs(4281) <= '0';
    layer0_outputs(4282) <= '1';
    layer0_outputs(4283) <= not((inputs(200)) and (inputs(98)));
    layer0_outputs(4284) <= inputs(93);
    layer0_outputs(4285) <= (inputs(21)) and not (inputs(169));
    layer0_outputs(4286) <= '0';
    layer0_outputs(4287) <= (inputs(176)) or (inputs(147));
    layer0_outputs(4288) <= not(inputs(74));
    layer0_outputs(4289) <= not((inputs(138)) xor (inputs(17)));
    layer0_outputs(4290) <= (inputs(211)) or (inputs(180));
    layer0_outputs(4291) <= '1';
    layer0_outputs(4292) <= (inputs(65)) and (inputs(185));
    layer0_outputs(4293) <= '0';
    layer0_outputs(4294) <= (inputs(152)) and (inputs(26));
    layer0_outputs(4295) <= not((inputs(44)) and (inputs(11)));
    layer0_outputs(4296) <= inputs(164);
    layer0_outputs(4297) <= (inputs(208)) and not (inputs(114));
    layer0_outputs(4298) <= not(inputs(253)) or (inputs(50));
    layer0_outputs(4299) <= (inputs(101)) xor (inputs(10));
    layer0_outputs(4300) <= not((inputs(154)) or (inputs(152)));
    layer0_outputs(4301) <= '0';
    layer0_outputs(4302) <= not((inputs(164)) or (inputs(195)));
    layer0_outputs(4303) <= (inputs(25)) and not (inputs(163));
    layer0_outputs(4304) <= not((inputs(64)) or (inputs(63)));
    layer0_outputs(4305) <= inputs(137);
    layer0_outputs(4306) <= not(inputs(26)) or (inputs(157));
    layer0_outputs(4307) <= not(inputs(176));
    layer0_outputs(4308) <= (inputs(32)) xor (inputs(246));
    layer0_outputs(4309) <= not((inputs(56)) or (inputs(244)));
    layer0_outputs(4310) <= (inputs(79)) xor (inputs(72));
    layer0_outputs(4311) <= (inputs(243)) and (inputs(155));
    layer0_outputs(4312) <= not((inputs(81)) and (inputs(180)));
    layer0_outputs(4313) <= not(inputs(118)) or (inputs(17));
    layer0_outputs(4314) <= not((inputs(47)) xor (inputs(109)));
    layer0_outputs(4315) <= inputs(74);
    layer0_outputs(4316) <= not((inputs(107)) or (inputs(175)));
    layer0_outputs(4317) <= '0';
    layer0_outputs(4318) <= not((inputs(194)) xor (inputs(189)));
    layer0_outputs(4319) <= not((inputs(82)) or (inputs(128)));
    layer0_outputs(4320) <= (inputs(151)) and not (inputs(5));
    layer0_outputs(4321) <= '1';
    layer0_outputs(4322) <= not((inputs(119)) and (inputs(38)));
    layer0_outputs(4323) <= inputs(0);
    layer0_outputs(4324) <= (inputs(20)) and not (inputs(249));
    layer0_outputs(4325) <= not((inputs(145)) xor (inputs(37)));
    layer0_outputs(4326) <= (inputs(165)) or (inputs(196));
    layer0_outputs(4327) <= not((inputs(43)) or (inputs(64)));
    layer0_outputs(4328) <= '1';
    layer0_outputs(4329) <= '0';
    layer0_outputs(4330) <= inputs(146);
    layer0_outputs(4331) <= not(inputs(77));
    layer0_outputs(4332) <= (inputs(48)) or (inputs(58));
    layer0_outputs(4333) <= not((inputs(167)) or (inputs(240)));
    layer0_outputs(4334) <= (inputs(93)) or (inputs(71));
    layer0_outputs(4335) <= not(inputs(99));
    layer0_outputs(4336) <= not(inputs(230));
    layer0_outputs(4337) <= not(inputs(167));
    layer0_outputs(4338) <= '0';
    layer0_outputs(4339) <= (inputs(229)) or (inputs(208));
    layer0_outputs(4340) <= not((inputs(32)) or (inputs(137)));
    layer0_outputs(4341) <= '1';
    layer0_outputs(4342) <= inputs(129);
    layer0_outputs(4343) <= not(inputs(10)) or (inputs(0));
    layer0_outputs(4344) <= '1';
    layer0_outputs(4345) <= '1';
    layer0_outputs(4346) <= (inputs(223)) or (inputs(242));
    layer0_outputs(4347) <= not(inputs(141));
    layer0_outputs(4348) <= not(inputs(12));
    layer0_outputs(4349) <= not(inputs(233));
    layer0_outputs(4350) <= not(inputs(55)) or (inputs(250));
    layer0_outputs(4351) <= not(inputs(217));
    layer0_outputs(4352) <= inputs(0);
    layer0_outputs(4353) <= not((inputs(154)) xor (inputs(171)));
    layer0_outputs(4354) <= not(inputs(130));
    layer0_outputs(4355) <= inputs(153);
    layer0_outputs(4356) <= (inputs(220)) and not (inputs(151));
    layer0_outputs(4357) <= not((inputs(204)) or (inputs(216)));
    layer0_outputs(4358) <= inputs(73);
    layer0_outputs(4359) <= not(inputs(151));
    layer0_outputs(4360) <= (inputs(143)) or (inputs(87));
    layer0_outputs(4361) <= not(inputs(169)) or (inputs(100));
    layer0_outputs(4362) <= (inputs(210)) or (inputs(233));
    layer0_outputs(4363) <= (inputs(123)) and (inputs(179));
    layer0_outputs(4364) <= not(inputs(87));
    layer0_outputs(4365) <= not(inputs(229)) or (inputs(59));
    layer0_outputs(4366) <= '0';
    layer0_outputs(4367) <= '1';
    layer0_outputs(4368) <= not(inputs(176));
    layer0_outputs(4369) <= not(inputs(67));
    layer0_outputs(4370) <= (inputs(81)) or (inputs(172));
    layer0_outputs(4371) <= not((inputs(195)) or (inputs(75)));
    layer0_outputs(4372) <= not(inputs(135));
    layer0_outputs(4373) <= not(inputs(206));
    layer0_outputs(4374) <= (inputs(116)) or (inputs(158));
    layer0_outputs(4375) <= not(inputs(105));
    layer0_outputs(4376) <= not((inputs(176)) and (inputs(28)));
    layer0_outputs(4377) <= not(inputs(64)) or (inputs(79));
    layer0_outputs(4378) <= (inputs(208)) or (inputs(27));
    layer0_outputs(4379) <= (inputs(218)) and not (inputs(31));
    layer0_outputs(4380) <= not(inputs(212)) or (inputs(1));
    layer0_outputs(4381) <= (inputs(206)) or (inputs(245));
    layer0_outputs(4382) <= inputs(16);
    layer0_outputs(4383) <= (inputs(11)) and not (inputs(149));
    layer0_outputs(4384) <= (inputs(158)) and not (inputs(64));
    layer0_outputs(4385) <= inputs(130);
    layer0_outputs(4386) <= not(inputs(147)) or (inputs(4));
    layer0_outputs(4387) <= (inputs(21)) or (inputs(33));
    layer0_outputs(4388) <= not(inputs(169));
    layer0_outputs(4389) <= not(inputs(181));
    layer0_outputs(4390) <= (inputs(49)) xor (inputs(18));
    layer0_outputs(4391) <= not(inputs(79));
    layer0_outputs(4392) <= not(inputs(252));
    layer0_outputs(4393) <= '0';
    layer0_outputs(4394) <= (inputs(227)) and not (inputs(5));
    layer0_outputs(4395) <= '1';
    layer0_outputs(4396) <= not((inputs(83)) xor (inputs(71)));
    layer0_outputs(4397) <= inputs(160);
    layer0_outputs(4398) <= '0';
    layer0_outputs(4399) <= not(inputs(194));
    layer0_outputs(4400) <= not(inputs(78));
    layer0_outputs(4401) <= not(inputs(213)) or (inputs(7));
    layer0_outputs(4402) <= (inputs(157)) or (inputs(239));
    layer0_outputs(4403) <= '1';
    layer0_outputs(4404) <= inputs(163);
    layer0_outputs(4405) <= not(inputs(231));
    layer0_outputs(4406) <= (inputs(255)) and not (inputs(69));
    layer0_outputs(4407) <= inputs(39);
    layer0_outputs(4408) <= (inputs(174)) and (inputs(181));
    layer0_outputs(4409) <= not((inputs(44)) and (inputs(78)));
    layer0_outputs(4410) <= not((inputs(214)) xor (inputs(231)));
    layer0_outputs(4411) <= inputs(123);
    layer0_outputs(4412) <= not((inputs(213)) or (inputs(56)));
    layer0_outputs(4413) <= '0';
    layer0_outputs(4414) <= (inputs(63)) or (inputs(31));
    layer0_outputs(4415) <= '1';
    layer0_outputs(4416) <= inputs(109);
    layer0_outputs(4417) <= inputs(2);
    layer0_outputs(4418) <= inputs(23);
    layer0_outputs(4419) <= '0';
    layer0_outputs(4420) <= '0';
    layer0_outputs(4421) <= '1';
    layer0_outputs(4422) <= not((inputs(188)) or (inputs(71)));
    layer0_outputs(4423) <= '1';
    layer0_outputs(4424) <= not(inputs(188));
    layer0_outputs(4425) <= not(inputs(170));
    layer0_outputs(4426) <= inputs(67);
    layer0_outputs(4427) <= (inputs(62)) and not (inputs(111));
    layer0_outputs(4428) <= not(inputs(97));
    layer0_outputs(4429) <= (inputs(89)) or (inputs(224));
    layer0_outputs(4430) <= (inputs(146)) and not (inputs(90));
    layer0_outputs(4431) <= '1';
    layer0_outputs(4432) <= inputs(253);
    layer0_outputs(4433) <= not(inputs(144));
    layer0_outputs(4434) <= '1';
    layer0_outputs(4435) <= '1';
    layer0_outputs(4436) <= not(inputs(167));
    layer0_outputs(4437) <= not(inputs(155));
    layer0_outputs(4438) <= (inputs(201)) and (inputs(189));
    layer0_outputs(4439) <= not((inputs(98)) and (inputs(96)));
    layer0_outputs(4440) <= (inputs(29)) or (inputs(254));
    layer0_outputs(4441) <= '0';
    layer0_outputs(4442) <= not((inputs(51)) and (inputs(207)));
    layer0_outputs(4443) <= inputs(68);
    layer0_outputs(4444) <= (inputs(230)) and not (inputs(108));
    layer0_outputs(4445) <= (inputs(67)) xor (inputs(53));
    layer0_outputs(4446) <= not((inputs(119)) xor (inputs(142)));
    layer0_outputs(4447) <= '1';
    layer0_outputs(4448) <= '0';
    layer0_outputs(4449) <= not(inputs(30));
    layer0_outputs(4450) <= (inputs(59)) and (inputs(78));
    layer0_outputs(4451) <= not(inputs(146)) or (inputs(139));
    layer0_outputs(4452) <= inputs(25);
    layer0_outputs(4453) <= inputs(200);
    layer0_outputs(4454) <= '0';
    layer0_outputs(4455) <= '1';
    layer0_outputs(4456) <= inputs(85);
    layer0_outputs(4457) <= inputs(112);
    layer0_outputs(4458) <= not(inputs(178));
    layer0_outputs(4459) <= not((inputs(98)) or (inputs(81)));
    layer0_outputs(4460) <= '0';
    layer0_outputs(4461) <= (inputs(163)) or (inputs(115));
    layer0_outputs(4462) <= not(inputs(81));
    layer0_outputs(4463) <= (inputs(224)) xor (inputs(145));
    layer0_outputs(4464) <= (inputs(192)) or (inputs(26));
    layer0_outputs(4465) <= '1';
    layer0_outputs(4466) <= (inputs(62)) and not (inputs(98));
    layer0_outputs(4467) <= '0';
    layer0_outputs(4468) <= (inputs(236)) or (inputs(48));
    layer0_outputs(4469) <= not(inputs(152)) or (inputs(205));
    layer0_outputs(4470) <= (inputs(202)) or (inputs(175));
    layer0_outputs(4471) <= not((inputs(184)) xor (inputs(215)));
    layer0_outputs(4472) <= '1';
    layer0_outputs(4473) <= (inputs(253)) and (inputs(25));
    layer0_outputs(4474) <= not((inputs(199)) and (inputs(60)));
    layer0_outputs(4475) <= inputs(228);
    layer0_outputs(4476) <= (inputs(112)) and not (inputs(83));
    layer0_outputs(4477) <= not((inputs(211)) and (inputs(59)));
    layer0_outputs(4478) <= (inputs(14)) and (inputs(82));
    layer0_outputs(4479) <= not(inputs(125));
    layer0_outputs(4480) <= not(inputs(145));
    layer0_outputs(4481) <= not(inputs(102));
    layer0_outputs(4482) <= (inputs(219)) and (inputs(212));
    layer0_outputs(4483) <= not((inputs(172)) or (inputs(44)));
    layer0_outputs(4484) <= not(inputs(83));
    layer0_outputs(4485) <= '1';
    layer0_outputs(4486) <= not(inputs(223));
    layer0_outputs(4487) <= '0';
    layer0_outputs(4488) <= not((inputs(250)) and (inputs(246)));
    layer0_outputs(4489) <= (inputs(224)) and (inputs(1));
    layer0_outputs(4490) <= not(inputs(43));
    layer0_outputs(4491) <= not((inputs(44)) or (inputs(253)));
    layer0_outputs(4492) <= not((inputs(65)) and (inputs(141)));
    layer0_outputs(4493) <= not((inputs(66)) or (inputs(122)));
    layer0_outputs(4494) <= (inputs(138)) or (inputs(237));
    layer0_outputs(4495) <= '1';
    layer0_outputs(4496) <= not(inputs(47));
    layer0_outputs(4497) <= not(inputs(227)) or (inputs(106));
    layer0_outputs(4498) <= (inputs(74)) or (inputs(50));
    layer0_outputs(4499) <= not(inputs(100));
    layer0_outputs(4500) <= not(inputs(126)) or (inputs(104));
    layer0_outputs(4501) <= (inputs(80)) and (inputs(130));
    layer0_outputs(4502) <= '1';
    layer0_outputs(4503) <= inputs(31);
    layer0_outputs(4504) <= '1';
    layer0_outputs(4505) <= inputs(150);
    layer0_outputs(4506) <= (inputs(109)) or (inputs(59));
    layer0_outputs(4507) <= (inputs(229)) and not (inputs(207));
    layer0_outputs(4508) <= not((inputs(232)) and (inputs(214)));
    layer0_outputs(4509) <= not(inputs(118));
    layer0_outputs(4510) <= not(inputs(189));
    layer0_outputs(4511) <= '0';
    layer0_outputs(4512) <= (inputs(73)) and not (inputs(147));
    layer0_outputs(4513) <= (inputs(119)) and not (inputs(103));
    layer0_outputs(4514) <= not((inputs(147)) and (inputs(126)));
    layer0_outputs(4515) <= not((inputs(111)) or (inputs(62)));
    layer0_outputs(4516) <= (inputs(188)) and not (inputs(7));
    layer0_outputs(4517) <= not((inputs(70)) and (inputs(9)));
    layer0_outputs(4518) <= not(inputs(193));
    layer0_outputs(4519) <= (inputs(233)) and (inputs(92));
    layer0_outputs(4520) <= not(inputs(17));
    layer0_outputs(4521) <= not(inputs(118)) or (inputs(135));
    layer0_outputs(4522) <= not(inputs(71)) or (inputs(206));
    layer0_outputs(4523) <= not(inputs(81));
    layer0_outputs(4524) <= (inputs(48)) and not (inputs(217));
    layer0_outputs(4525) <= not((inputs(37)) and (inputs(8)));
    layer0_outputs(4526) <= not((inputs(137)) or (inputs(222)));
    layer0_outputs(4527) <= not((inputs(78)) and (inputs(43)));
    layer0_outputs(4528) <= not(inputs(107));
    layer0_outputs(4529) <= inputs(220);
    layer0_outputs(4530) <= not(inputs(65));
    layer0_outputs(4531) <= not((inputs(234)) or (inputs(238)));
    layer0_outputs(4532) <= '1';
    layer0_outputs(4533) <= (inputs(217)) or (inputs(211));
    layer0_outputs(4534) <= not(inputs(177));
    layer0_outputs(4535) <= (inputs(235)) or (inputs(49));
    layer0_outputs(4536) <= not(inputs(232));
    layer0_outputs(4537) <= not(inputs(212));
    layer0_outputs(4538) <= '1';
    layer0_outputs(4539) <= not(inputs(229));
    layer0_outputs(4540) <= '1';
    layer0_outputs(4541) <= inputs(13);
    layer0_outputs(4542) <= '0';
    layer0_outputs(4543) <= not((inputs(145)) and (inputs(158)));
    layer0_outputs(4544) <= (inputs(4)) and not (inputs(17));
    layer0_outputs(4545) <= not(inputs(129));
    layer0_outputs(4546) <= not((inputs(102)) or (inputs(249)));
    layer0_outputs(4547) <= not(inputs(167)) or (inputs(192));
    layer0_outputs(4548) <= (inputs(253)) and not (inputs(244));
    layer0_outputs(4549) <= not((inputs(3)) and (inputs(153)));
    layer0_outputs(4550) <= not((inputs(71)) xor (inputs(145)));
    layer0_outputs(4551) <= inputs(195);
    layer0_outputs(4552) <= not(inputs(104)) or (inputs(135));
    layer0_outputs(4553) <= (inputs(186)) and not (inputs(212));
    layer0_outputs(4554) <= (inputs(14)) and not (inputs(49));
    layer0_outputs(4555) <= not(inputs(145));
    layer0_outputs(4556) <= (inputs(108)) and (inputs(186));
    layer0_outputs(4557) <= not((inputs(48)) or (inputs(36)));
    layer0_outputs(4558) <= not(inputs(232));
    layer0_outputs(4559) <= not(inputs(61)) or (inputs(206));
    layer0_outputs(4560) <= (inputs(105)) or (inputs(82));
    layer0_outputs(4561) <= not(inputs(198)) or (inputs(171));
    layer0_outputs(4562) <= not(inputs(88));
    layer0_outputs(4563) <= inputs(82);
    layer0_outputs(4564) <= '0';
    layer0_outputs(4565) <= (inputs(105)) and (inputs(85));
    layer0_outputs(4566) <= not(inputs(216));
    layer0_outputs(4567) <= not(inputs(157));
    layer0_outputs(4568) <= (inputs(238)) and not (inputs(62));
    layer0_outputs(4569) <= '1';
    layer0_outputs(4570) <= not(inputs(25));
    layer0_outputs(4571) <= not((inputs(29)) or (inputs(72)));
    layer0_outputs(4572) <= (inputs(154)) or (inputs(117));
    layer0_outputs(4573) <= inputs(115);
    layer0_outputs(4574) <= inputs(7);
    layer0_outputs(4575) <= inputs(114);
    layer0_outputs(4576) <= (inputs(182)) and (inputs(253));
    layer0_outputs(4577) <= (inputs(23)) and (inputs(212));
    layer0_outputs(4578) <= '0';
    layer0_outputs(4579) <= '0';
    layer0_outputs(4580) <= not(inputs(230)) or (inputs(60));
    layer0_outputs(4581) <= not((inputs(64)) or (inputs(196)));
    layer0_outputs(4582) <= inputs(226);
    layer0_outputs(4583) <= not(inputs(38));
    layer0_outputs(4584) <= '1';
    layer0_outputs(4585) <= not(inputs(247)) or (inputs(76));
    layer0_outputs(4586) <= (inputs(68)) xor (inputs(239));
    layer0_outputs(4587) <= '0';
    layer0_outputs(4588) <= inputs(149);
    layer0_outputs(4589) <= not(inputs(148));
    layer0_outputs(4590) <= inputs(196);
    layer0_outputs(4591) <= '0';
    layer0_outputs(4592) <= '1';
    layer0_outputs(4593) <= inputs(203);
    layer0_outputs(4594) <= not((inputs(140)) xor (inputs(249)));
    layer0_outputs(4595) <= (inputs(151)) and not (inputs(46));
    layer0_outputs(4596) <= not(inputs(196)) or (inputs(91));
    layer0_outputs(4597) <= '1';
    layer0_outputs(4598) <= '0';
    layer0_outputs(4599) <= not(inputs(95)) or (inputs(91));
    layer0_outputs(4600) <= '1';
    layer0_outputs(4601) <= not(inputs(211));
    layer0_outputs(4602) <= not(inputs(193)) or (inputs(165));
    layer0_outputs(4603) <= '1';
    layer0_outputs(4604) <= (inputs(199)) and (inputs(190));
    layer0_outputs(4605) <= (inputs(118)) xor (inputs(131));
    layer0_outputs(4606) <= '1';
    layer0_outputs(4607) <= inputs(106);
    layer0_outputs(4608) <= (inputs(41)) and (inputs(113));
    layer0_outputs(4609) <= not((inputs(195)) or (inputs(236)));
    layer0_outputs(4610) <= inputs(195);
    layer0_outputs(4611) <= (inputs(31)) and (inputs(32));
    layer0_outputs(4612) <= not((inputs(88)) and (inputs(122)));
    layer0_outputs(4613) <= inputs(213);
    layer0_outputs(4614) <= '0';
    layer0_outputs(4615) <= (inputs(61)) and not (inputs(105));
    layer0_outputs(4616) <= not(inputs(150));
    layer0_outputs(4617) <= '0';
    layer0_outputs(4618) <= not((inputs(113)) or (inputs(121)));
    layer0_outputs(4619) <= not(inputs(196));
    layer0_outputs(4620) <= not((inputs(79)) xor (inputs(26)));
    layer0_outputs(4621) <= not(inputs(175));
    layer0_outputs(4622) <= (inputs(254)) and (inputs(48));
    layer0_outputs(4623) <= (inputs(15)) and (inputs(3));
    layer0_outputs(4624) <= (inputs(116)) and (inputs(65));
    layer0_outputs(4625) <= (inputs(109)) or (inputs(235));
    layer0_outputs(4626) <= inputs(246);
    layer0_outputs(4627) <= not(inputs(19));
    layer0_outputs(4628) <= not((inputs(18)) or (inputs(63)));
    layer0_outputs(4629) <= not(inputs(167)) or (inputs(238));
    layer0_outputs(4630) <= (inputs(199)) xor (inputs(240));
    layer0_outputs(4631) <= '1';
    layer0_outputs(4632) <= '1';
    layer0_outputs(4633) <= not(inputs(23));
    layer0_outputs(4634) <= not((inputs(225)) or (inputs(178)));
    layer0_outputs(4635) <= not(inputs(198));
    layer0_outputs(4636) <= not((inputs(177)) or (inputs(207)));
    layer0_outputs(4637) <= not(inputs(9)) or (inputs(241));
    layer0_outputs(4638) <= '1';
    layer0_outputs(4639) <= (inputs(125)) and not (inputs(37));
    layer0_outputs(4640) <= not((inputs(6)) or (inputs(196)));
    layer0_outputs(4641) <= inputs(186);
    layer0_outputs(4642) <= inputs(150);
    layer0_outputs(4643) <= not(inputs(187)) or (inputs(1));
    layer0_outputs(4644) <= not((inputs(111)) or (inputs(21)));
    layer0_outputs(4645) <= (inputs(232)) and not (inputs(198));
    layer0_outputs(4646) <= '1';
    layer0_outputs(4647) <= not(inputs(242)) or (inputs(185));
    layer0_outputs(4648) <= inputs(180);
    layer0_outputs(4649) <= '1';
    layer0_outputs(4650) <= inputs(33);
    layer0_outputs(4651) <= not((inputs(192)) xor (inputs(152)));
    layer0_outputs(4652) <= not(inputs(52));
    layer0_outputs(4653) <= inputs(103);
    layer0_outputs(4654) <= (inputs(76)) or (inputs(43));
    layer0_outputs(4655) <= (inputs(120)) and not (inputs(63));
    layer0_outputs(4656) <= not(inputs(6));
    layer0_outputs(4657) <= not(inputs(127));
    layer0_outputs(4658) <= not((inputs(111)) xor (inputs(9)));
    layer0_outputs(4659) <= '0';
    layer0_outputs(4660) <= '1';
    layer0_outputs(4661) <= inputs(76);
    layer0_outputs(4662) <= not(inputs(111));
    layer0_outputs(4663) <= not(inputs(43)) or (inputs(89));
    layer0_outputs(4664) <= not(inputs(246));
    layer0_outputs(4665) <= '0';
    layer0_outputs(4666) <= inputs(58);
    layer0_outputs(4667) <= (inputs(228)) and not (inputs(158));
    layer0_outputs(4668) <= not(inputs(72));
    layer0_outputs(4669) <= (inputs(135)) and (inputs(131));
    layer0_outputs(4670) <= (inputs(160)) and not (inputs(239));
    layer0_outputs(4671) <= not((inputs(81)) or (inputs(184)));
    layer0_outputs(4672) <= inputs(211);
    layer0_outputs(4673) <= not((inputs(226)) or (inputs(174)));
    layer0_outputs(4674) <= (inputs(134)) or (inputs(154));
    layer0_outputs(4675) <= (inputs(28)) xor (inputs(196));
    layer0_outputs(4676) <= '1';
    layer0_outputs(4677) <= not(inputs(0));
    layer0_outputs(4678) <= not(inputs(180)) or (inputs(13));
    layer0_outputs(4679) <= not((inputs(162)) or (inputs(47)));
    layer0_outputs(4680) <= not(inputs(158));
    layer0_outputs(4681) <= not(inputs(172));
    layer0_outputs(4682) <= (inputs(11)) and not (inputs(165));
    layer0_outputs(4683) <= (inputs(81)) or (inputs(182));
    layer0_outputs(4684) <= (inputs(1)) or (inputs(91));
    layer0_outputs(4685) <= inputs(95);
    layer0_outputs(4686) <= (inputs(189)) and not (inputs(169));
    layer0_outputs(4687) <= (inputs(38)) and (inputs(105));
    layer0_outputs(4688) <= inputs(74);
    layer0_outputs(4689) <= not(inputs(206)) or (inputs(10));
    layer0_outputs(4690) <= inputs(66);
    layer0_outputs(4691) <= not(inputs(84));
    layer0_outputs(4692) <= inputs(10);
    layer0_outputs(4693) <= not(inputs(214)) or (inputs(39));
    layer0_outputs(4694) <= '0';
    layer0_outputs(4695) <= inputs(25);
    layer0_outputs(4696) <= not((inputs(89)) or (inputs(53)));
    layer0_outputs(4697) <= not((inputs(94)) or (inputs(22)));
    layer0_outputs(4698) <= not((inputs(205)) and (inputs(185)));
    layer0_outputs(4699) <= inputs(189);
    layer0_outputs(4700) <= not(inputs(167)) or (inputs(133));
    layer0_outputs(4701) <= not(inputs(147));
    layer0_outputs(4702) <= not((inputs(87)) xor (inputs(79)));
    layer0_outputs(4703) <= (inputs(27)) and not (inputs(251));
    layer0_outputs(4704) <= '1';
    layer0_outputs(4705) <= inputs(167);
    layer0_outputs(4706) <= inputs(138);
    layer0_outputs(4707) <= not(inputs(219));
    layer0_outputs(4708) <= (inputs(83)) or (inputs(144));
    layer0_outputs(4709) <= (inputs(117)) or (inputs(155));
    layer0_outputs(4710) <= inputs(178);
    layer0_outputs(4711) <= '0';
    layer0_outputs(4712) <= (inputs(33)) and not (inputs(129));
    layer0_outputs(4713) <= inputs(255);
    layer0_outputs(4714) <= '0';
    layer0_outputs(4715) <= not((inputs(249)) or (inputs(3)));
    layer0_outputs(4716) <= not(inputs(129)) or (inputs(75));
    layer0_outputs(4717) <= not(inputs(97));
    layer0_outputs(4718) <= '1';
    layer0_outputs(4719) <= (inputs(104)) or (inputs(31));
    layer0_outputs(4720) <= not(inputs(138));
    layer0_outputs(4721) <= (inputs(62)) xor (inputs(232));
    layer0_outputs(4722) <= inputs(33);
    layer0_outputs(4723) <= not(inputs(1));
    layer0_outputs(4724) <= (inputs(239)) or (inputs(167));
    layer0_outputs(4725) <= not((inputs(57)) and (inputs(41)));
    layer0_outputs(4726) <= not(inputs(164));
    layer0_outputs(4727) <= not(inputs(152)) or (inputs(79));
    layer0_outputs(4728) <= '0';
    layer0_outputs(4729) <= (inputs(142)) and not (inputs(46));
    layer0_outputs(4730) <= '0';
    layer0_outputs(4731) <= not((inputs(119)) and (inputs(137)));
    layer0_outputs(4732) <= not((inputs(216)) and (inputs(145)));
    layer0_outputs(4733) <= (inputs(6)) and not (inputs(132));
    layer0_outputs(4734) <= not((inputs(180)) or (inputs(147)));
    layer0_outputs(4735) <= '0';
    layer0_outputs(4736) <= (inputs(13)) xor (inputs(124));
    layer0_outputs(4737) <= (inputs(242)) and (inputs(159));
    layer0_outputs(4738) <= not(inputs(145));
    layer0_outputs(4739) <= not(inputs(251)) or (inputs(10));
    layer0_outputs(4740) <= not(inputs(133)) or (inputs(213));
    layer0_outputs(4741) <= (inputs(103)) and not (inputs(4));
    layer0_outputs(4742) <= (inputs(230)) and (inputs(45));
    layer0_outputs(4743) <= (inputs(173)) and not (inputs(36));
    layer0_outputs(4744) <= not((inputs(255)) xor (inputs(98)));
    layer0_outputs(4745) <= '1';
    layer0_outputs(4746) <= not(inputs(248));
    layer0_outputs(4747) <= '0';
    layer0_outputs(4748) <= '0';
    layer0_outputs(4749) <= not(inputs(42));
    layer0_outputs(4750) <= not(inputs(172));
    layer0_outputs(4751) <= not(inputs(57)) or (inputs(172));
    layer0_outputs(4752) <= not(inputs(204));
    layer0_outputs(4753) <= not((inputs(195)) and (inputs(229)));
    layer0_outputs(4754) <= not(inputs(247));
    layer0_outputs(4755) <= (inputs(74)) or (inputs(24));
    layer0_outputs(4756) <= not(inputs(188));
    layer0_outputs(4757) <= '0';
    layer0_outputs(4758) <= (inputs(70)) and not (inputs(36));
    layer0_outputs(4759) <= not(inputs(96));
    layer0_outputs(4760) <= not(inputs(54)) or (inputs(154));
    layer0_outputs(4761) <= inputs(137);
    layer0_outputs(4762) <= (inputs(30)) and not (inputs(105));
    layer0_outputs(4763) <= not((inputs(140)) or (inputs(131)));
    layer0_outputs(4764) <= not(inputs(35)) or (inputs(203));
    layer0_outputs(4765) <= not(inputs(91));
    layer0_outputs(4766) <= not((inputs(237)) or (inputs(107)));
    layer0_outputs(4767) <= '0';
    layer0_outputs(4768) <= (inputs(13)) and not (inputs(96));
    layer0_outputs(4769) <= not(inputs(182)) or (inputs(27));
    layer0_outputs(4770) <= not(inputs(197)) or (inputs(107));
    layer0_outputs(4771) <= not(inputs(124)) or (inputs(56));
    layer0_outputs(4772) <= '0';
    layer0_outputs(4773) <= not(inputs(123));
    layer0_outputs(4774) <= '0';
    layer0_outputs(4775) <= not((inputs(38)) or (inputs(203)));
    layer0_outputs(4776) <= inputs(160);
    layer0_outputs(4777) <= '0';
    layer0_outputs(4778) <= '1';
    layer0_outputs(4779) <= (inputs(43)) or (inputs(44));
    layer0_outputs(4780) <= not((inputs(170)) or (inputs(100)));
    layer0_outputs(4781) <= inputs(138);
    layer0_outputs(4782) <= '1';
    layer0_outputs(4783) <= (inputs(192)) and not (inputs(205));
    layer0_outputs(4784) <= inputs(154);
    layer0_outputs(4785) <= (inputs(123)) or (inputs(140));
    layer0_outputs(4786) <= not(inputs(110)) or (inputs(171));
    layer0_outputs(4787) <= not(inputs(45));
    layer0_outputs(4788) <= not(inputs(94));
    layer0_outputs(4789) <= (inputs(39)) and (inputs(88));
    layer0_outputs(4790) <= not(inputs(221));
    layer0_outputs(4791) <= '0';
    layer0_outputs(4792) <= (inputs(123)) and not (inputs(242));
    layer0_outputs(4793) <= not(inputs(101));
    layer0_outputs(4794) <= (inputs(253)) or (inputs(52));
    layer0_outputs(4795) <= not(inputs(102)) or (inputs(139));
    layer0_outputs(4796) <= not(inputs(177)) or (inputs(89));
    layer0_outputs(4797) <= (inputs(5)) or (inputs(127));
    layer0_outputs(4798) <= not(inputs(94));
    layer0_outputs(4799) <= '0';
    layer0_outputs(4800) <= inputs(150);
    layer0_outputs(4801) <= not(inputs(27)) or (inputs(106));
    layer0_outputs(4802) <= (inputs(157)) and not (inputs(85));
    layer0_outputs(4803) <= not((inputs(156)) or (inputs(187)));
    layer0_outputs(4804) <= (inputs(115)) and (inputs(129));
    layer0_outputs(4805) <= not((inputs(196)) and (inputs(154)));
    layer0_outputs(4806) <= inputs(120);
    layer0_outputs(4807) <= (inputs(235)) and (inputs(20));
    layer0_outputs(4808) <= not(inputs(16)) or (inputs(100));
    layer0_outputs(4809) <= (inputs(2)) or (inputs(22));
    layer0_outputs(4810) <= not((inputs(6)) xor (inputs(11)));
    layer0_outputs(4811) <= not((inputs(204)) and (inputs(30)));
    layer0_outputs(4812) <= (inputs(228)) xor (inputs(198));
    layer0_outputs(4813) <= '1';
    layer0_outputs(4814) <= (inputs(189)) and not (inputs(118));
    layer0_outputs(4815) <= not(inputs(245)) or (inputs(1));
    layer0_outputs(4816) <= inputs(144);
    layer0_outputs(4817) <= (inputs(73)) or (inputs(91));
    layer0_outputs(4818) <= '0';
    layer0_outputs(4819) <= '1';
    layer0_outputs(4820) <= not(inputs(200)) or (inputs(141));
    layer0_outputs(4821) <= not(inputs(108));
    layer0_outputs(4822) <= (inputs(14)) and not (inputs(134));
    layer0_outputs(4823) <= not((inputs(85)) and (inputs(216)));
    layer0_outputs(4824) <= '1';
    layer0_outputs(4825) <= (inputs(219)) and not (inputs(51));
    layer0_outputs(4826) <= '1';
    layer0_outputs(4827) <= not(inputs(118));
    layer0_outputs(4828) <= not((inputs(6)) or (inputs(73)));
    layer0_outputs(4829) <= (inputs(181)) and not (inputs(244));
    layer0_outputs(4830) <= (inputs(42)) xor (inputs(44));
    layer0_outputs(4831) <= inputs(180);
    layer0_outputs(4832) <= inputs(78);
    layer0_outputs(4833) <= not((inputs(228)) or (inputs(234)));
    layer0_outputs(4834) <= not((inputs(208)) or (inputs(221)));
    layer0_outputs(4835) <= not(inputs(101)) or (inputs(35));
    layer0_outputs(4836) <= (inputs(164)) or (inputs(171));
    layer0_outputs(4837) <= (inputs(5)) or (inputs(130));
    layer0_outputs(4838) <= '0';
    layer0_outputs(4839) <= '1';
    layer0_outputs(4840) <= (inputs(121)) or (inputs(19));
    layer0_outputs(4841) <= not((inputs(213)) or (inputs(209)));
    layer0_outputs(4842) <= not((inputs(243)) or (inputs(214)));
    layer0_outputs(4843) <= not(inputs(18)) or (inputs(156));
    layer0_outputs(4844) <= not(inputs(139)) or (inputs(222));
    layer0_outputs(4845) <= not((inputs(190)) or (inputs(110)));
    layer0_outputs(4846) <= inputs(162);
    layer0_outputs(4847) <= (inputs(204)) or (inputs(56));
    layer0_outputs(4848) <= (inputs(7)) or (inputs(20));
    layer0_outputs(4849) <= not(inputs(231));
    layer0_outputs(4850) <= not(inputs(24));
    layer0_outputs(4851) <= inputs(150);
    layer0_outputs(4852) <= not(inputs(183)) or (inputs(147));
    layer0_outputs(4853) <= (inputs(216)) or (inputs(234));
    layer0_outputs(4854) <= not(inputs(173));
    layer0_outputs(4855) <= inputs(53);
    layer0_outputs(4856) <= '0';
    layer0_outputs(4857) <= not(inputs(111));
    layer0_outputs(4858) <= not(inputs(124));
    layer0_outputs(4859) <= not((inputs(54)) and (inputs(29)));
    layer0_outputs(4860) <= not(inputs(119)) or (inputs(49));
    layer0_outputs(4861) <= (inputs(143)) and not (inputs(96));
    layer0_outputs(4862) <= not(inputs(115));
    layer0_outputs(4863) <= (inputs(81)) and (inputs(186));
    layer0_outputs(4864) <= inputs(181);
    layer0_outputs(4865) <= '1';
    layer0_outputs(4866) <= (inputs(224)) and (inputs(2));
    layer0_outputs(4867) <= inputs(192);
    layer0_outputs(4868) <= not(inputs(94));
    layer0_outputs(4869) <= (inputs(211)) and not (inputs(59));
    layer0_outputs(4870) <= not(inputs(89)) or (inputs(203));
    layer0_outputs(4871) <= not(inputs(205)) or (inputs(212));
    layer0_outputs(4872) <= not((inputs(38)) and (inputs(20)));
    layer0_outputs(4873) <= '0';
    layer0_outputs(4874) <= not(inputs(62));
    layer0_outputs(4875) <= '0';
    layer0_outputs(4876) <= not(inputs(145));
    layer0_outputs(4877) <= inputs(235);
    layer0_outputs(4878) <= not(inputs(202)) or (inputs(205));
    layer0_outputs(4879) <= inputs(181);
    layer0_outputs(4880) <= not((inputs(168)) and (inputs(205)));
    layer0_outputs(4881) <= inputs(23);
    layer0_outputs(4882) <= '0';
    layer0_outputs(4883) <= '1';
    layer0_outputs(4884) <= (inputs(99)) and not (inputs(198));
    layer0_outputs(4885) <= (inputs(53)) and (inputs(25));
    layer0_outputs(4886) <= not((inputs(216)) and (inputs(78)));
    layer0_outputs(4887) <= (inputs(255)) or (inputs(179));
    layer0_outputs(4888) <= not((inputs(32)) xor (inputs(248)));
    layer0_outputs(4889) <= inputs(120);
    layer0_outputs(4890) <= inputs(146);
    layer0_outputs(4891) <= inputs(26);
    layer0_outputs(4892) <= not((inputs(55)) or (inputs(93)));
    layer0_outputs(4893) <= not(inputs(17)) or (inputs(238));
    layer0_outputs(4894) <= not((inputs(131)) or (inputs(132)));
    layer0_outputs(4895) <= (inputs(157)) and not (inputs(155));
    layer0_outputs(4896) <= not(inputs(73));
    layer0_outputs(4897) <= not((inputs(229)) or (inputs(126)));
    layer0_outputs(4898) <= not(inputs(34)) or (inputs(142));
    layer0_outputs(4899) <= not(inputs(120));
    layer0_outputs(4900) <= '0';
    layer0_outputs(4901) <= not((inputs(175)) or (inputs(30)));
    layer0_outputs(4902) <= inputs(5);
    layer0_outputs(4903) <= inputs(23);
    layer0_outputs(4904) <= not((inputs(3)) or (inputs(33)));
    layer0_outputs(4905) <= not((inputs(108)) or (inputs(113)));
    layer0_outputs(4906) <= (inputs(11)) xor (inputs(94));
    layer0_outputs(4907) <= not(inputs(54)) or (inputs(48));
    layer0_outputs(4908) <= (inputs(73)) and not (inputs(133));
    layer0_outputs(4909) <= inputs(1);
    layer0_outputs(4910) <= not(inputs(163));
    layer0_outputs(4911) <= not(inputs(69));
    layer0_outputs(4912) <= '1';
    layer0_outputs(4913) <= not((inputs(109)) or (inputs(20)));
    layer0_outputs(4914) <= not((inputs(214)) and (inputs(250)));
    layer0_outputs(4915) <= not(inputs(102));
    layer0_outputs(4916) <= (inputs(9)) or (inputs(155));
    layer0_outputs(4917) <= not(inputs(66));
    layer0_outputs(4918) <= not((inputs(56)) or (inputs(87)));
    layer0_outputs(4919) <= '0';
    layer0_outputs(4920) <= '0';
    layer0_outputs(4921) <= '0';
    layer0_outputs(4922) <= inputs(89);
    layer0_outputs(4923) <= inputs(109);
    layer0_outputs(4924) <= inputs(45);
    layer0_outputs(4925) <= not(inputs(19)) or (inputs(207));
    layer0_outputs(4926) <= not(inputs(190)) or (inputs(104));
    layer0_outputs(4927) <= not(inputs(74));
    layer0_outputs(4928) <= not(inputs(24)) or (inputs(85));
    layer0_outputs(4929) <= (inputs(23)) and not (inputs(213));
    layer0_outputs(4930) <= inputs(93);
    layer0_outputs(4931) <= '0';
    layer0_outputs(4932) <= '1';
    layer0_outputs(4933) <= not(inputs(135));
    layer0_outputs(4934) <= not(inputs(45)) or (inputs(237));
    layer0_outputs(4935) <= not(inputs(84));
    layer0_outputs(4936) <= not(inputs(25));
    layer0_outputs(4937) <= inputs(86);
    layer0_outputs(4938) <= not((inputs(140)) and (inputs(229)));
    layer0_outputs(4939) <= not((inputs(195)) or (inputs(142)));
    layer0_outputs(4940) <= not(inputs(64));
    layer0_outputs(4941) <= (inputs(222)) or (inputs(225));
    layer0_outputs(4942) <= not(inputs(181));
    layer0_outputs(4943) <= '0';
    layer0_outputs(4944) <= not((inputs(49)) and (inputs(126)));
    layer0_outputs(4945) <= (inputs(115)) and not (inputs(18));
    layer0_outputs(4946) <= not(inputs(248));
    layer0_outputs(4947) <= '1';
    layer0_outputs(4948) <= (inputs(71)) and not (inputs(188));
    layer0_outputs(4949) <= not(inputs(51)) or (inputs(146));
    layer0_outputs(4950) <= not(inputs(127));
    layer0_outputs(4951) <= inputs(212);
    layer0_outputs(4952) <= inputs(140);
    layer0_outputs(4953) <= (inputs(159)) and (inputs(172));
    layer0_outputs(4954) <= (inputs(167)) or (inputs(107));
    layer0_outputs(4955) <= not(inputs(24));
    layer0_outputs(4956) <= (inputs(110)) or (inputs(231));
    layer0_outputs(4957) <= inputs(143);
    layer0_outputs(4958) <= inputs(227);
    layer0_outputs(4959) <= '1';
    layer0_outputs(4960) <= '1';
    layer0_outputs(4961) <= inputs(8);
    layer0_outputs(4962) <= (inputs(210)) or (inputs(227));
    layer0_outputs(4963) <= inputs(213);
    layer0_outputs(4964) <= not((inputs(180)) xor (inputs(176)));
    layer0_outputs(4965) <= (inputs(19)) and not (inputs(36));
    layer0_outputs(4966) <= (inputs(17)) or (inputs(169));
    layer0_outputs(4967) <= inputs(5);
    layer0_outputs(4968) <= not((inputs(9)) and (inputs(212)));
    layer0_outputs(4969) <= (inputs(215)) xor (inputs(159));
    layer0_outputs(4970) <= not(inputs(104));
    layer0_outputs(4971) <= (inputs(80)) and not (inputs(235));
    layer0_outputs(4972) <= inputs(15);
    layer0_outputs(4973) <= inputs(85);
    layer0_outputs(4974) <= '0';
    layer0_outputs(4975) <= not(inputs(29));
    layer0_outputs(4976) <= '0';
    layer0_outputs(4977) <= inputs(140);
    layer0_outputs(4978) <= (inputs(210)) or (inputs(96));
    layer0_outputs(4979) <= not(inputs(95));
    layer0_outputs(4980) <= not((inputs(52)) xor (inputs(72)));
    layer0_outputs(4981) <= not(inputs(129));
    layer0_outputs(4982) <= not(inputs(246)) or (inputs(251));
    layer0_outputs(4983) <= '1';
    layer0_outputs(4984) <= not(inputs(200)) or (inputs(134));
    layer0_outputs(4985) <= (inputs(244)) and (inputs(199));
    layer0_outputs(4986) <= '0';
    layer0_outputs(4987) <= (inputs(129)) and not (inputs(3));
    layer0_outputs(4988) <= not((inputs(177)) or (inputs(71)));
    layer0_outputs(4989) <= inputs(134);
    layer0_outputs(4990) <= (inputs(216)) or (inputs(163));
    layer0_outputs(4991) <= inputs(60);
    layer0_outputs(4992) <= '0';
    layer0_outputs(4993) <= (inputs(101)) and (inputs(250));
    layer0_outputs(4994) <= not((inputs(11)) and (inputs(162)));
    layer0_outputs(4995) <= not(inputs(232));
    layer0_outputs(4996) <= '1';
    layer0_outputs(4997) <= (inputs(100)) and not (inputs(143));
    layer0_outputs(4998) <= (inputs(161)) and (inputs(201));
    layer0_outputs(4999) <= (inputs(45)) and (inputs(148));
    layer0_outputs(5000) <= '0';
    layer0_outputs(5001) <= not(inputs(209));
    layer0_outputs(5002) <= not(inputs(106));
    layer0_outputs(5003) <= not(inputs(219));
    layer0_outputs(5004) <= inputs(77);
    layer0_outputs(5005) <= '0';
    layer0_outputs(5006) <= not((inputs(121)) or (inputs(20)));
    layer0_outputs(5007) <= '1';
    layer0_outputs(5008) <= (inputs(228)) or (inputs(243));
    layer0_outputs(5009) <= not(inputs(24)) or (inputs(116));
    layer0_outputs(5010) <= (inputs(13)) and not (inputs(11));
    layer0_outputs(5011) <= (inputs(186)) and not (inputs(26));
    layer0_outputs(5012) <= '1';
    layer0_outputs(5013) <= not(inputs(90));
    layer0_outputs(5014) <= (inputs(146)) or (inputs(65));
    layer0_outputs(5015) <= not((inputs(175)) or (inputs(129)));
    layer0_outputs(5016) <= inputs(54);
    layer0_outputs(5017) <= inputs(78);
    layer0_outputs(5018) <= not(inputs(147));
    layer0_outputs(5019) <= not(inputs(48)) or (inputs(12));
    layer0_outputs(5020) <= '1';
    layer0_outputs(5021) <= '0';
    layer0_outputs(5022) <= not((inputs(134)) and (inputs(44)));
    layer0_outputs(5023) <= (inputs(111)) or (inputs(123));
    layer0_outputs(5024) <= (inputs(68)) and not (inputs(32));
    layer0_outputs(5025) <= inputs(238);
    layer0_outputs(5026) <= (inputs(145)) and (inputs(251));
    layer0_outputs(5027) <= (inputs(104)) and (inputs(45));
    layer0_outputs(5028) <= (inputs(245)) or (inputs(189));
    layer0_outputs(5029) <= '1';
    layer0_outputs(5030) <= not((inputs(102)) or (inputs(18)));
    layer0_outputs(5031) <= not(inputs(6)) or (inputs(182));
    layer0_outputs(5032) <= not(inputs(232));
    layer0_outputs(5033) <= (inputs(91)) or (inputs(252));
    layer0_outputs(5034) <= not((inputs(221)) or (inputs(170)));
    layer0_outputs(5035) <= not(inputs(184));
    layer0_outputs(5036) <= not(inputs(60)) or (inputs(132));
    layer0_outputs(5037) <= (inputs(38)) and not (inputs(249));
    layer0_outputs(5038) <= inputs(226);
    layer0_outputs(5039) <= not((inputs(26)) and (inputs(94)));
    layer0_outputs(5040) <= not((inputs(23)) xor (inputs(33)));
    layer0_outputs(5041) <= '0';
    layer0_outputs(5042) <= (inputs(99)) and not (inputs(42));
    layer0_outputs(5043) <= (inputs(228)) or (inputs(200));
    layer0_outputs(5044) <= inputs(103);
    layer0_outputs(5045) <= inputs(231);
    layer0_outputs(5046) <= inputs(101);
    layer0_outputs(5047) <= not((inputs(80)) xor (inputs(217)));
    layer0_outputs(5048) <= (inputs(61)) and not (inputs(121));
    layer0_outputs(5049) <= not((inputs(141)) or (inputs(142)));
    layer0_outputs(5050) <= not((inputs(46)) or (inputs(92)));
    layer0_outputs(5051) <= inputs(112);
    layer0_outputs(5052) <= (inputs(244)) and not (inputs(78));
    layer0_outputs(5053) <= inputs(141);
    layer0_outputs(5054) <= (inputs(175)) and not (inputs(244));
    layer0_outputs(5055) <= '0';
    layer0_outputs(5056) <= not((inputs(117)) and (inputs(197)));
    layer0_outputs(5057) <= inputs(43);
    layer0_outputs(5058) <= '0';
    layer0_outputs(5059) <= not((inputs(40)) or (inputs(95)));
    layer0_outputs(5060) <= inputs(40);
    layer0_outputs(5061) <= not((inputs(36)) and (inputs(125)));
    layer0_outputs(5062) <= (inputs(183)) and not (inputs(81));
    layer0_outputs(5063) <= not(inputs(101)) or (inputs(116));
    layer0_outputs(5064) <= (inputs(117)) and not (inputs(126));
    layer0_outputs(5065) <= not(inputs(230)) or (inputs(152));
    layer0_outputs(5066) <= (inputs(125)) or (inputs(119));
    layer0_outputs(5067) <= not(inputs(89)) or (inputs(132));
    layer0_outputs(5068) <= (inputs(126)) xor (inputs(35));
    layer0_outputs(5069) <= (inputs(155)) and (inputs(41));
    layer0_outputs(5070) <= not((inputs(147)) and (inputs(74)));
    layer0_outputs(5071) <= not(inputs(98)) or (inputs(77));
    layer0_outputs(5072) <= not((inputs(60)) and (inputs(7)));
    layer0_outputs(5073) <= inputs(136);
    layer0_outputs(5074) <= (inputs(46)) or (inputs(29));
    layer0_outputs(5075) <= not(inputs(84)) or (inputs(158));
    layer0_outputs(5076) <= not(inputs(71));
    layer0_outputs(5077) <= not(inputs(59));
    layer0_outputs(5078) <= not(inputs(8)) or (inputs(52));
    layer0_outputs(5079) <= (inputs(69)) or (inputs(178));
    layer0_outputs(5080) <= not((inputs(235)) or (inputs(45)));
    layer0_outputs(5081) <= not(inputs(60));
    layer0_outputs(5082) <= not(inputs(108));
    layer0_outputs(5083) <= (inputs(184)) and not (inputs(114));
    layer0_outputs(5084) <= (inputs(19)) and (inputs(126));
    layer0_outputs(5085) <= not(inputs(80)) or (inputs(125));
    layer0_outputs(5086) <= not(inputs(130)) or (inputs(95));
    layer0_outputs(5087) <= (inputs(115)) or (inputs(59));
    layer0_outputs(5088) <= not((inputs(189)) xor (inputs(81)));
    layer0_outputs(5089) <= not((inputs(121)) and (inputs(31)));
    layer0_outputs(5090) <= inputs(209);
    layer0_outputs(5091) <= (inputs(22)) or (inputs(96));
    layer0_outputs(5092) <= '0';
    layer0_outputs(5093) <= not((inputs(161)) and (inputs(48)));
    layer0_outputs(5094) <= not(inputs(9));
    layer0_outputs(5095) <= not(inputs(180));
    layer0_outputs(5096) <= (inputs(97)) and not (inputs(206));
    layer0_outputs(5097) <= not(inputs(122));
    layer0_outputs(5098) <= not(inputs(108)) or (inputs(128));
    layer0_outputs(5099) <= not(inputs(2));
    layer0_outputs(5100) <= '0';
    layer0_outputs(5101) <= inputs(39);
    layer0_outputs(5102) <= not(inputs(150));
    layer0_outputs(5103) <= '1';
    layer0_outputs(5104) <= not((inputs(6)) and (inputs(58)));
    layer0_outputs(5105) <= not(inputs(253));
    layer0_outputs(5106) <= inputs(42);
    layer0_outputs(5107) <= (inputs(188)) or (inputs(122));
    layer0_outputs(5108) <= not((inputs(90)) and (inputs(170)));
    layer0_outputs(5109) <= (inputs(239)) and (inputs(91));
    layer0_outputs(5110) <= (inputs(21)) or (inputs(97));
    layer0_outputs(5111) <= not(inputs(245));
    layer0_outputs(5112) <= inputs(252);
    layer0_outputs(5113) <= (inputs(60)) and not (inputs(234));
    layer0_outputs(5114) <= (inputs(225)) and not (inputs(205));
    layer0_outputs(5115) <= inputs(173);
    layer0_outputs(5116) <= not(inputs(207)) or (inputs(192));
    layer0_outputs(5117) <= not(inputs(77));
    layer0_outputs(5118) <= (inputs(133)) and (inputs(22));
    layer0_outputs(5119) <= not(inputs(38)) or (inputs(219));
    layer1_outputs(0) <= layer0_outputs(3866);
    layer1_outputs(1) <= not((layer0_outputs(3056)) and (layer0_outputs(911)));
    layer1_outputs(2) <= (layer0_outputs(3954)) and not (layer0_outputs(2064));
    layer1_outputs(3) <= not(layer0_outputs(2494));
    layer1_outputs(4) <= (layer0_outputs(4962)) or (layer0_outputs(3113));
    layer1_outputs(5) <= not(layer0_outputs(3427)) or (layer0_outputs(48));
    layer1_outputs(6) <= not((layer0_outputs(4614)) and (layer0_outputs(2464)));
    layer1_outputs(7) <= (layer0_outputs(1053)) or (layer0_outputs(3966));
    layer1_outputs(8) <= not(layer0_outputs(4795));
    layer1_outputs(9) <= '0';
    layer1_outputs(10) <= '0';
    layer1_outputs(11) <= '0';
    layer1_outputs(12) <= not(layer0_outputs(412)) or (layer0_outputs(1426));
    layer1_outputs(13) <= not((layer0_outputs(1204)) xor (layer0_outputs(829)));
    layer1_outputs(14) <= layer0_outputs(3705);
    layer1_outputs(15) <= layer0_outputs(3045);
    layer1_outputs(16) <= (layer0_outputs(1700)) or (layer0_outputs(3532));
    layer1_outputs(17) <= (layer0_outputs(4456)) and not (layer0_outputs(1827));
    layer1_outputs(18) <= not(layer0_outputs(4779)) or (layer0_outputs(1566));
    layer1_outputs(19) <= not((layer0_outputs(3119)) and (layer0_outputs(4245)));
    layer1_outputs(20) <= (layer0_outputs(3982)) or (layer0_outputs(2375));
    layer1_outputs(21) <= not(layer0_outputs(426));
    layer1_outputs(22) <= not((layer0_outputs(4589)) and (layer0_outputs(2659)));
    layer1_outputs(23) <= layer0_outputs(3073);
    layer1_outputs(24) <= layer0_outputs(3687);
    layer1_outputs(25) <= not(layer0_outputs(569)) or (layer0_outputs(193));
    layer1_outputs(26) <= (layer0_outputs(4052)) and not (layer0_outputs(3646));
    layer1_outputs(27) <= not(layer0_outputs(1891));
    layer1_outputs(28) <= (layer0_outputs(1148)) and not (layer0_outputs(138));
    layer1_outputs(29) <= (layer0_outputs(1797)) and not (layer0_outputs(206));
    layer1_outputs(30) <= layer0_outputs(332);
    layer1_outputs(31) <= not((layer0_outputs(29)) and (layer0_outputs(903)));
    layer1_outputs(32) <= not((layer0_outputs(4075)) and (layer0_outputs(3509)));
    layer1_outputs(33) <= (layer0_outputs(2533)) and not (layer0_outputs(2283));
    layer1_outputs(34) <= '1';
    layer1_outputs(35) <= layer0_outputs(1760);
    layer1_outputs(36) <= not((layer0_outputs(1922)) or (layer0_outputs(1182)));
    layer1_outputs(37) <= not(layer0_outputs(4278));
    layer1_outputs(38) <= '1';
    layer1_outputs(39) <= not(layer0_outputs(4017));
    layer1_outputs(40) <= not(layer0_outputs(1902));
    layer1_outputs(41) <= (layer0_outputs(3504)) and (layer0_outputs(1957));
    layer1_outputs(42) <= layer0_outputs(2825);
    layer1_outputs(43) <= (layer0_outputs(4210)) or (layer0_outputs(2300));
    layer1_outputs(44) <= not(layer0_outputs(4360));
    layer1_outputs(45) <= not(layer0_outputs(4129)) or (layer0_outputs(3979));
    layer1_outputs(46) <= not((layer0_outputs(4314)) and (layer0_outputs(3844)));
    layer1_outputs(47) <= (layer0_outputs(1038)) or (layer0_outputs(281));
    layer1_outputs(48) <= '1';
    layer1_outputs(49) <= (layer0_outputs(2792)) and not (layer0_outputs(1691));
    layer1_outputs(50) <= (layer0_outputs(4549)) and (layer0_outputs(5052));
    layer1_outputs(51) <= not(layer0_outputs(3203));
    layer1_outputs(52) <= not((layer0_outputs(1614)) or (layer0_outputs(3588)));
    layer1_outputs(53) <= layer0_outputs(5086);
    layer1_outputs(54) <= (layer0_outputs(4770)) xor (layer0_outputs(3734));
    layer1_outputs(55) <= '0';
    layer1_outputs(56) <= not(layer0_outputs(2874)) or (layer0_outputs(1825));
    layer1_outputs(57) <= (layer0_outputs(333)) or (layer0_outputs(3325));
    layer1_outputs(58) <= not(layer0_outputs(1843));
    layer1_outputs(59) <= not((layer0_outputs(4765)) and (layer0_outputs(3132)));
    layer1_outputs(60) <= '0';
    layer1_outputs(61) <= not((layer0_outputs(2759)) or (layer0_outputs(2325)));
    layer1_outputs(62) <= not(layer0_outputs(2842)) or (layer0_outputs(2730));
    layer1_outputs(63) <= (layer0_outputs(285)) xor (layer0_outputs(2802));
    layer1_outputs(64) <= not((layer0_outputs(872)) xor (layer0_outputs(3455)));
    layer1_outputs(65) <= '0';
    layer1_outputs(66) <= not(layer0_outputs(4330));
    layer1_outputs(67) <= '0';
    layer1_outputs(68) <= (layer0_outputs(377)) and (layer0_outputs(1988));
    layer1_outputs(69) <= (layer0_outputs(4762)) and (layer0_outputs(4192));
    layer1_outputs(70) <= not(layer0_outputs(2480));
    layer1_outputs(71) <= not((layer0_outputs(1669)) and (layer0_outputs(1542)));
    layer1_outputs(72) <= layer0_outputs(1448);
    layer1_outputs(73) <= not(layer0_outputs(3927));
    layer1_outputs(74) <= layer0_outputs(1805);
    layer1_outputs(75) <= (layer0_outputs(2138)) or (layer0_outputs(525));
    layer1_outputs(76) <= (layer0_outputs(3227)) and not (layer0_outputs(2062));
    layer1_outputs(77) <= not((layer0_outputs(3464)) and (layer0_outputs(4355)));
    layer1_outputs(78) <= '1';
    layer1_outputs(79) <= not((layer0_outputs(4425)) and (layer0_outputs(2374)));
    layer1_outputs(80) <= '0';
    layer1_outputs(81) <= not(layer0_outputs(4528)) or (layer0_outputs(1052));
    layer1_outputs(82) <= not(layer0_outputs(1170));
    layer1_outputs(83) <= layer0_outputs(3739);
    layer1_outputs(84) <= not(layer0_outputs(78));
    layer1_outputs(85) <= '0';
    layer1_outputs(86) <= '0';
    layer1_outputs(87) <= not((layer0_outputs(4576)) and (layer0_outputs(2709)));
    layer1_outputs(88) <= '0';
    layer1_outputs(89) <= not(layer0_outputs(3740)) or (layer0_outputs(3327));
    layer1_outputs(90) <= not((layer0_outputs(370)) and (layer0_outputs(4016)));
    layer1_outputs(91) <= (layer0_outputs(1915)) or (layer0_outputs(3709));
    layer1_outputs(92) <= not(layer0_outputs(4691));
    layer1_outputs(93) <= not(layer0_outputs(1695)) or (layer0_outputs(1511));
    layer1_outputs(94) <= layer0_outputs(2208);
    layer1_outputs(95) <= not(layer0_outputs(1846)) or (layer0_outputs(3181));
    layer1_outputs(96) <= layer0_outputs(1859);
    layer1_outputs(97) <= (layer0_outputs(3304)) and (layer0_outputs(2947));
    layer1_outputs(98) <= not(layer0_outputs(1591));
    layer1_outputs(99) <= (layer0_outputs(2416)) and not (layer0_outputs(2792));
    layer1_outputs(100) <= not(layer0_outputs(1104));
    layer1_outputs(101) <= not((layer0_outputs(3668)) or (layer0_outputs(542)));
    layer1_outputs(102) <= not(layer0_outputs(1178)) or (layer0_outputs(4034));
    layer1_outputs(103) <= not((layer0_outputs(928)) or (layer0_outputs(2633)));
    layer1_outputs(104) <= not(layer0_outputs(5087)) or (layer0_outputs(2786));
    layer1_outputs(105) <= (layer0_outputs(1711)) or (layer0_outputs(1675));
    layer1_outputs(106) <= not((layer0_outputs(4508)) or (layer0_outputs(2612)));
    layer1_outputs(107) <= '0';
    layer1_outputs(108) <= not(layer0_outputs(2940));
    layer1_outputs(109) <= not(layer0_outputs(3390)) or (layer0_outputs(2594));
    layer1_outputs(110) <= not((layer0_outputs(2488)) and (layer0_outputs(648)));
    layer1_outputs(111) <= (layer0_outputs(3582)) and (layer0_outputs(990));
    layer1_outputs(112) <= not(layer0_outputs(3778));
    layer1_outputs(113) <= not(layer0_outputs(3360));
    layer1_outputs(114) <= not((layer0_outputs(283)) or (layer0_outputs(3860)));
    layer1_outputs(115) <= not(layer0_outputs(1552));
    layer1_outputs(116) <= (layer0_outputs(2056)) or (layer0_outputs(4240));
    layer1_outputs(117) <= not((layer0_outputs(4571)) or (layer0_outputs(4021)));
    layer1_outputs(118) <= '1';
    layer1_outputs(119) <= not((layer0_outputs(519)) and (layer0_outputs(915)));
    layer1_outputs(120) <= (layer0_outputs(3249)) or (layer0_outputs(3352));
    layer1_outputs(121) <= '0';
    layer1_outputs(122) <= (layer0_outputs(4206)) and not (layer0_outputs(3564));
    layer1_outputs(123) <= not(layer0_outputs(1297));
    layer1_outputs(124) <= '0';
    layer1_outputs(125) <= not(layer0_outputs(1929)) or (layer0_outputs(3610));
    layer1_outputs(126) <= '0';
    layer1_outputs(127) <= '0';
    layer1_outputs(128) <= '0';
    layer1_outputs(129) <= layer0_outputs(1638);
    layer1_outputs(130) <= '1';
    layer1_outputs(131) <= not((layer0_outputs(4100)) and (layer0_outputs(5090)));
    layer1_outputs(132) <= not(layer0_outputs(1558));
    layer1_outputs(133) <= layer0_outputs(789);
    layer1_outputs(134) <= (layer0_outputs(4643)) and (layer0_outputs(2935));
    layer1_outputs(135) <= not(layer0_outputs(1369)) or (layer0_outputs(2836));
    layer1_outputs(136) <= (layer0_outputs(319)) and not (layer0_outputs(809));
    layer1_outputs(137) <= not((layer0_outputs(602)) or (layer0_outputs(1303)));
    layer1_outputs(138) <= not((layer0_outputs(98)) or (layer0_outputs(4299)));
    layer1_outputs(139) <= (layer0_outputs(1082)) or (layer0_outputs(4677));
    layer1_outputs(140) <= not(layer0_outputs(107)) or (layer0_outputs(736));
    layer1_outputs(141) <= layer0_outputs(4641);
    layer1_outputs(142) <= layer0_outputs(5106);
    layer1_outputs(143) <= (layer0_outputs(431)) and (layer0_outputs(4860));
    layer1_outputs(144) <= not(layer0_outputs(2587));
    layer1_outputs(145) <= '1';
    layer1_outputs(146) <= layer0_outputs(2071);
    layer1_outputs(147) <= layer0_outputs(1835);
    layer1_outputs(148) <= not(layer0_outputs(4099)) or (layer0_outputs(996));
    layer1_outputs(149) <= layer0_outputs(83);
    layer1_outputs(150) <= not((layer0_outputs(3544)) or (layer0_outputs(3645)));
    layer1_outputs(151) <= layer0_outputs(4284);
    layer1_outputs(152) <= (layer0_outputs(307)) and (layer0_outputs(967));
    layer1_outputs(153) <= layer0_outputs(120);
    layer1_outputs(154) <= (layer0_outputs(3)) and not (layer0_outputs(4537));
    layer1_outputs(155) <= (layer0_outputs(2718)) xor (layer0_outputs(2702));
    layer1_outputs(156) <= not((layer0_outputs(4412)) xor (layer0_outputs(274)));
    layer1_outputs(157) <= (layer0_outputs(3228)) and (layer0_outputs(2396));
    layer1_outputs(158) <= (layer0_outputs(4302)) and (layer0_outputs(232));
    layer1_outputs(159) <= not(layer0_outputs(4803));
    layer1_outputs(160) <= '1';
    layer1_outputs(161) <= (layer0_outputs(2970)) and not (layer0_outputs(5111));
    layer1_outputs(162) <= not((layer0_outputs(4950)) or (layer0_outputs(121)));
    layer1_outputs(163) <= (layer0_outputs(3376)) and not (layer0_outputs(1113));
    layer1_outputs(164) <= not(layer0_outputs(3502));
    layer1_outputs(165) <= not(layer0_outputs(2866));
    layer1_outputs(166) <= not((layer0_outputs(3867)) and (layer0_outputs(1279)));
    layer1_outputs(167) <= '0';
    layer1_outputs(168) <= '1';
    layer1_outputs(169) <= layer0_outputs(1429);
    layer1_outputs(170) <= layer0_outputs(1669);
    layer1_outputs(171) <= (layer0_outputs(532)) and not (layer0_outputs(2869));
    layer1_outputs(172) <= not(layer0_outputs(1437));
    layer1_outputs(173) <= layer0_outputs(4389);
    layer1_outputs(174) <= (layer0_outputs(4416)) and not (layer0_outputs(678));
    layer1_outputs(175) <= not(layer0_outputs(4919)) or (layer0_outputs(3354));
    layer1_outputs(176) <= (layer0_outputs(429)) and not (layer0_outputs(311));
    layer1_outputs(177) <= '1';
    layer1_outputs(178) <= '0';
    layer1_outputs(179) <= not((layer0_outputs(3034)) and (layer0_outputs(3029)));
    layer1_outputs(180) <= not(layer0_outputs(1723)) or (layer0_outputs(4243));
    layer1_outputs(181) <= not((layer0_outputs(4406)) or (layer0_outputs(934)));
    layer1_outputs(182) <= not(layer0_outputs(1286));
    layer1_outputs(183) <= not((layer0_outputs(2140)) or (layer0_outputs(2302)));
    layer1_outputs(184) <= (layer0_outputs(4922)) and (layer0_outputs(4082));
    layer1_outputs(185) <= not(layer0_outputs(2740));
    layer1_outputs(186) <= (layer0_outputs(2871)) and (layer0_outputs(2748));
    layer1_outputs(187) <= '1';
    layer1_outputs(188) <= '1';
    layer1_outputs(189) <= not(layer0_outputs(1947));
    layer1_outputs(190) <= (layer0_outputs(4019)) and not (layer0_outputs(740));
    layer1_outputs(191) <= not((layer0_outputs(520)) or (layer0_outputs(746)));
    layer1_outputs(192) <= not((layer0_outputs(3474)) and (layer0_outputs(82)));
    layer1_outputs(193) <= not(layer0_outputs(1653));
    layer1_outputs(194) <= not(layer0_outputs(1951));
    layer1_outputs(195) <= not(layer0_outputs(2956)) or (layer0_outputs(3031));
    layer1_outputs(196) <= not((layer0_outputs(3524)) and (layer0_outputs(2027)));
    layer1_outputs(197) <= not((layer0_outputs(1408)) and (layer0_outputs(1987)));
    layer1_outputs(198) <= (layer0_outputs(5094)) and not (layer0_outputs(3125));
    layer1_outputs(199) <= not(layer0_outputs(4460)) or (layer0_outputs(375));
    layer1_outputs(200) <= (layer0_outputs(2053)) and not (layer0_outputs(3532));
    layer1_outputs(201) <= (layer0_outputs(3753)) and not (layer0_outputs(903));
    layer1_outputs(202) <= (layer0_outputs(3768)) and not (layer0_outputs(677));
    layer1_outputs(203) <= not((layer0_outputs(548)) and (layer0_outputs(3627)));
    layer1_outputs(204) <= (layer0_outputs(4806)) or (layer0_outputs(885));
    layer1_outputs(205) <= not(layer0_outputs(3173));
    layer1_outputs(206) <= layer0_outputs(3790);
    layer1_outputs(207) <= layer0_outputs(1342);
    layer1_outputs(208) <= '1';
    layer1_outputs(209) <= (layer0_outputs(4713)) and not (layer0_outputs(1104));
    layer1_outputs(210) <= not(layer0_outputs(2577));
    layer1_outputs(211) <= layer0_outputs(260);
    layer1_outputs(212) <= (layer0_outputs(2633)) and not (layer0_outputs(1197));
    layer1_outputs(213) <= '0';
    layer1_outputs(214) <= '0';
    layer1_outputs(215) <= layer0_outputs(2464);
    layer1_outputs(216) <= '0';
    layer1_outputs(217) <= (layer0_outputs(3750)) or (layer0_outputs(1871));
    layer1_outputs(218) <= not((layer0_outputs(4743)) or (layer0_outputs(317)));
    layer1_outputs(219) <= '0';
    layer1_outputs(220) <= not((layer0_outputs(2404)) and (layer0_outputs(5069)));
    layer1_outputs(221) <= layer0_outputs(493);
    layer1_outputs(222) <= (layer0_outputs(1824)) or (layer0_outputs(925));
    layer1_outputs(223) <= not(layer0_outputs(1434));
    layer1_outputs(224) <= (layer0_outputs(3050)) and (layer0_outputs(1973));
    layer1_outputs(225) <= (layer0_outputs(2906)) xor (layer0_outputs(3432));
    layer1_outputs(226) <= not(layer0_outputs(2186)) or (layer0_outputs(216));
    layer1_outputs(227) <= '0';
    layer1_outputs(228) <= not((layer0_outputs(931)) and (layer0_outputs(1789)));
    layer1_outputs(229) <= layer0_outputs(2899);
    layer1_outputs(230) <= '1';
    layer1_outputs(231) <= not((layer0_outputs(3100)) or (layer0_outputs(3248)));
    layer1_outputs(232) <= not(layer0_outputs(4327)) or (layer0_outputs(2122));
    layer1_outputs(233) <= not((layer0_outputs(4868)) or (layer0_outputs(103)));
    layer1_outputs(234) <= (layer0_outputs(3847)) and (layer0_outputs(2173));
    layer1_outputs(235) <= (layer0_outputs(660)) and (layer0_outputs(1563));
    layer1_outputs(236) <= (layer0_outputs(4652)) and not (layer0_outputs(580));
    layer1_outputs(237) <= '1';
    layer1_outputs(238) <= not((layer0_outputs(20)) and (layer0_outputs(1864)));
    layer1_outputs(239) <= (layer0_outputs(890)) and not (layer0_outputs(3065));
    layer1_outputs(240) <= (layer0_outputs(2614)) and not (layer0_outputs(3810));
    layer1_outputs(241) <= not(layer0_outputs(256)) or (layer0_outputs(4853));
    layer1_outputs(242) <= not(layer0_outputs(1696)) or (layer0_outputs(1548));
    layer1_outputs(243) <= not(layer0_outputs(2308)) or (layer0_outputs(764));
    layer1_outputs(244) <= (layer0_outputs(2885)) and (layer0_outputs(1774));
    layer1_outputs(245) <= not(layer0_outputs(4731)) or (layer0_outputs(892));
    layer1_outputs(246) <= '0';
    layer1_outputs(247) <= not((layer0_outputs(350)) or (layer0_outputs(2581)));
    layer1_outputs(248) <= not((layer0_outputs(2576)) and (layer0_outputs(4883)));
    layer1_outputs(249) <= layer0_outputs(4965);
    layer1_outputs(250) <= not((layer0_outputs(42)) and (layer0_outputs(2874)));
    layer1_outputs(251) <= not(layer0_outputs(2834));
    layer1_outputs(252) <= not(layer0_outputs(1262)) or (layer0_outputs(4408));
    layer1_outputs(253) <= (layer0_outputs(980)) and (layer0_outputs(3859));
    layer1_outputs(254) <= '1';
    layer1_outputs(255) <= not(layer0_outputs(3654)) or (layer0_outputs(1433));
    layer1_outputs(256) <= (layer0_outputs(3264)) and not (layer0_outputs(2560));
    layer1_outputs(257) <= (layer0_outputs(1086)) or (layer0_outputs(3290));
    layer1_outputs(258) <= layer0_outputs(2202);
    layer1_outputs(259) <= layer0_outputs(421);
    layer1_outputs(260) <= '0';
    layer1_outputs(261) <= '1';
    layer1_outputs(262) <= not((layer0_outputs(2637)) and (layer0_outputs(102)));
    layer1_outputs(263) <= '1';
    layer1_outputs(264) <= (layer0_outputs(343)) and not (layer0_outputs(5000));
    layer1_outputs(265) <= (layer0_outputs(3144)) and not (layer0_outputs(1782));
    layer1_outputs(266) <= layer0_outputs(1496);
    layer1_outputs(267) <= layer0_outputs(4337);
    layer1_outputs(268) <= not(layer0_outputs(3556)) or (layer0_outputs(2666));
    layer1_outputs(269) <= not((layer0_outputs(4479)) or (layer0_outputs(128)));
    layer1_outputs(270) <= (layer0_outputs(4979)) and (layer0_outputs(3605));
    layer1_outputs(271) <= not((layer0_outputs(471)) and (layer0_outputs(4892)));
    layer1_outputs(272) <= (layer0_outputs(1386)) and (layer0_outputs(1124));
    layer1_outputs(273) <= layer0_outputs(5087);
    layer1_outputs(274) <= layer0_outputs(3190);
    layer1_outputs(275) <= (layer0_outputs(344)) and not (layer0_outputs(2849));
    layer1_outputs(276) <= layer0_outputs(5117);
    layer1_outputs(277) <= '1';
    layer1_outputs(278) <= (layer0_outputs(878)) and not (layer0_outputs(4046));
    layer1_outputs(279) <= (layer0_outputs(507)) and (layer0_outputs(2789));
    layer1_outputs(280) <= not(layer0_outputs(17));
    layer1_outputs(281) <= (layer0_outputs(1466)) and not (layer0_outputs(4309));
    layer1_outputs(282) <= (layer0_outputs(3082)) xor (layer0_outputs(489));
    layer1_outputs(283) <= layer0_outputs(4887);
    layer1_outputs(284) <= not((layer0_outputs(1185)) and (layer0_outputs(2178)));
    layer1_outputs(285) <= (layer0_outputs(793)) and not (layer0_outputs(561));
    layer1_outputs(286) <= not((layer0_outputs(4183)) and (layer0_outputs(558)));
    layer1_outputs(287) <= not(layer0_outputs(4287));
    layer1_outputs(288) <= layer0_outputs(1207);
    layer1_outputs(289) <= not(layer0_outputs(478)) or (layer0_outputs(1614));
    layer1_outputs(290) <= not((layer0_outputs(4233)) and (layer0_outputs(4287)));
    layer1_outputs(291) <= not((layer0_outputs(1026)) or (layer0_outputs(2220)));
    layer1_outputs(292) <= (layer0_outputs(4782)) or (layer0_outputs(2648));
    layer1_outputs(293) <= (layer0_outputs(2868)) and not (layer0_outputs(4445));
    layer1_outputs(294) <= not(layer0_outputs(1035));
    layer1_outputs(295) <= layer0_outputs(222);
    layer1_outputs(296) <= not(layer0_outputs(3580)) or (layer0_outputs(1509));
    layer1_outputs(297) <= not((layer0_outputs(1339)) or (layer0_outputs(4857)));
    layer1_outputs(298) <= '1';
    layer1_outputs(299) <= not(layer0_outputs(3055));
    layer1_outputs(300) <= (layer0_outputs(5004)) or (layer0_outputs(2047));
    layer1_outputs(301) <= (layer0_outputs(921)) and not (layer0_outputs(1414));
    layer1_outputs(302) <= not(layer0_outputs(3514)) or (layer0_outputs(3819));
    layer1_outputs(303) <= not((layer0_outputs(1837)) or (layer0_outputs(3092)));
    layer1_outputs(304) <= (layer0_outputs(916)) and (layer0_outputs(1377));
    layer1_outputs(305) <= '0';
    layer1_outputs(306) <= '1';
    layer1_outputs(307) <= layer0_outputs(224);
    layer1_outputs(308) <= layer0_outputs(2750);
    layer1_outputs(309) <= '1';
    layer1_outputs(310) <= not(layer0_outputs(3566)) or (layer0_outputs(4665));
    layer1_outputs(311) <= not(layer0_outputs(3363)) or (layer0_outputs(213));
    layer1_outputs(312) <= not(layer0_outputs(421));
    layer1_outputs(313) <= '1';
    layer1_outputs(314) <= not(layer0_outputs(4432));
    layer1_outputs(315) <= not((layer0_outputs(2078)) and (layer0_outputs(4144)));
    layer1_outputs(316) <= '0';
    layer1_outputs(317) <= (layer0_outputs(4779)) and not (layer0_outputs(2457));
    layer1_outputs(318) <= not(layer0_outputs(1472));
    layer1_outputs(319) <= layer0_outputs(319);
    layer1_outputs(320) <= (layer0_outputs(623)) and not (layer0_outputs(61));
    layer1_outputs(321) <= '1';
    layer1_outputs(322) <= layer0_outputs(2361);
    layer1_outputs(323) <= not(layer0_outputs(797));
    layer1_outputs(324) <= '0';
    layer1_outputs(325) <= (layer0_outputs(3850)) and not (layer0_outputs(3946));
    layer1_outputs(326) <= layer0_outputs(4551);
    layer1_outputs(327) <= not((layer0_outputs(409)) and (layer0_outputs(2400)));
    layer1_outputs(328) <= (layer0_outputs(2524)) or (layer0_outputs(4346));
    layer1_outputs(329) <= not(layer0_outputs(2050)) or (layer0_outputs(2107));
    layer1_outputs(330) <= not(layer0_outputs(1068)) or (layer0_outputs(1184));
    layer1_outputs(331) <= layer0_outputs(1198);
    layer1_outputs(332) <= (layer0_outputs(4271)) and (layer0_outputs(3914));
    layer1_outputs(333) <= (layer0_outputs(2670)) and not (layer0_outputs(3365));
    layer1_outputs(334) <= (layer0_outputs(1578)) or (layer0_outputs(1344));
    layer1_outputs(335) <= not(layer0_outputs(2159));
    layer1_outputs(336) <= not((layer0_outputs(1136)) or (layer0_outputs(4680)));
    layer1_outputs(337) <= '1';
    layer1_outputs(338) <= '0';
    layer1_outputs(339) <= (layer0_outputs(4815)) and (layer0_outputs(1543));
    layer1_outputs(340) <= not(layer0_outputs(4800));
    layer1_outputs(341) <= layer0_outputs(2055);
    layer1_outputs(342) <= not((layer0_outputs(3051)) and (layer0_outputs(1242)));
    layer1_outputs(343) <= '1';
    layer1_outputs(344) <= (layer0_outputs(261)) xor (layer0_outputs(3963));
    layer1_outputs(345) <= not(layer0_outputs(1820)) or (layer0_outputs(4182));
    layer1_outputs(346) <= '0';
    layer1_outputs(347) <= '1';
    layer1_outputs(348) <= not(layer0_outputs(3102));
    layer1_outputs(349) <= not(layer0_outputs(3283));
    layer1_outputs(350) <= not(layer0_outputs(3616));
    layer1_outputs(351) <= not((layer0_outputs(2945)) or (layer0_outputs(2998)));
    layer1_outputs(352) <= (layer0_outputs(4620)) and not (layer0_outputs(1616));
    layer1_outputs(353) <= '0';
    layer1_outputs(354) <= (layer0_outputs(4563)) and not (layer0_outputs(4927));
    layer1_outputs(355) <= layer0_outputs(3512);
    layer1_outputs(356) <= not(layer0_outputs(4570)) or (layer0_outputs(3219));
    layer1_outputs(357) <= not(layer0_outputs(2827)) or (layer0_outputs(4304));
    layer1_outputs(358) <= not(layer0_outputs(1668)) or (layer0_outputs(5046));
    layer1_outputs(359) <= '0';
    layer1_outputs(360) <= not(layer0_outputs(247));
    layer1_outputs(361) <= '1';
    layer1_outputs(362) <= not((layer0_outputs(18)) or (layer0_outputs(3823)));
    layer1_outputs(363) <= layer0_outputs(3727);
    layer1_outputs(364) <= (layer0_outputs(5056)) or (layer0_outputs(3226));
    layer1_outputs(365) <= not((layer0_outputs(941)) or (layer0_outputs(741)));
    layer1_outputs(366) <= not(layer0_outputs(2118));
    layer1_outputs(367) <= (layer0_outputs(2930)) and not (layer0_outputs(1605));
    layer1_outputs(368) <= layer0_outputs(2318);
    layer1_outputs(369) <= (layer0_outputs(4294)) and (layer0_outputs(5074));
    layer1_outputs(370) <= not(layer0_outputs(1127));
    layer1_outputs(371) <= not(layer0_outputs(3278));
    layer1_outputs(372) <= (layer0_outputs(1258)) and not (layer0_outputs(4550));
    layer1_outputs(373) <= '1';
    layer1_outputs(374) <= (layer0_outputs(1956)) and (layer0_outputs(3609));
    layer1_outputs(375) <= layer0_outputs(1477);
    layer1_outputs(376) <= '0';
    layer1_outputs(377) <= layer0_outputs(4506);
    layer1_outputs(378) <= (layer0_outputs(3910)) or (layer0_outputs(2148));
    layer1_outputs(379) <= (layer0_outputs(1627)) and not (layer0_outputs(1136));
    layer1_outputs(380) <= not(layer0_outputs(1489));
    layer1_outputs(381) <= not(layer0_outputs(1152)) or (layer0_outputs(132));
    layer1_outputs(382) <= not((layer0_outputs(1646)) or (layer0_outputs(709)));
    layer1_outputs(383) <= (layer0_outputs(4486)) and (layer0_outputs(2453));
    layer1_outputs(384) <= (layer0_outputs(4336)) and (layer0_outputs(1916));
    layer1_outputs(385) <= not(layer0_outputs(2744));
    layer1_outputs(386) <= not(layer0_outputs(873)) or (layer0_outputs(2162));
    layer1_outputs(387) <= not(layer0_outputs(2961));
    layer1_outputs(388) <= layer0_outputs(4419);
    layer1_outputs(389) <= '1';
    layer1_outputs(390) <= layer0_outputs(2853);
    layer1_outputs(391) <= '0';
    layer1_outputs(392) <= layer0_outputs(5014);
    layer1_outputs(393) <= not(layer0_outputs(3663)) or (layer0_outputs(2395));
    layer1_outputs(394) <= layer0_outputs(3151);
    layer1_outputs(395) <= (layer0_outputs(3602)) or (layer0_outputs(1855));
    layer1_outputs(396) <= not(layer0_outputs(2225)) or (layer0_outputs(4199));
    layer1_outputs(397) <= layer0_outputs(785);
    layer1_outputs(398) <= not(layer0_outputs(3265));
    layer1_outputs(399) <= (layer0_outputs(1361)) and not (layer0_outputs(2821));
    layer1_outputs(400) <= not(layer0_outputs(3139));
    layer1_outputs(401) <= not(layer0_outputs(1384)) or (layer0_outputs(1046));
    layer1_outputs(402) <= not((layer0_outputs(3525)) and (layer0_outputs(2928)));
    layer1_outputs(403) <= (layer0_outputs(1609)) and not (layer0_outputs(5057));
    layer1_outputs(404) <= layer0_outputs(1078);
    layer1_outputs(405) <= not(layer0_outputs(4749)) or (layer0_outputs(727));
    layer1_outputs(406) <= (layer0_outputs(4530)) and not (layer0_outputs(1334));
    layer1_outputs(407) <= not(layer0_outputs(4298)) or (layer0_outputs(35));
    layer1_outputs(408) <= layer0_outputs(250);
    layer1_outputs(409) <= '0';
    layer1_outputs(410) <= (layer0_outputs(3338)) xor (layer0_outputs(2795));
    layer1_outputs(411) <= not((layer0_outputs(337)) or (layer0_outputs(3691)));
    layer1_outputs(412) <= not((layer0_outputs(2782)) or (layer0_outputs(439)));
    layer1_outputs(413) <= layer0_outputs(114);
    layer1_outputs(414) <= not(layer0_outputs(2817)) or (layer0_outputs(4504));
    layer1_outputs(415) <= '1';
    layer1_outputs(416) <= layer0_outputs(1464);
    layer1_outputs(417) <= (layer0_outputs(1257)) and (layer0_outputs(485));
    layer1_outputs(418) <= (layer0_outputs(1288)) and (layer0_outputs(1858));
    layer1_outputs(419) <= not(layer0_outputs(4585));
    layer1_outputs(420) <= '0';
    layer1_outputs(421) <= layer0_outputs(4719);
    layer1_outputs(422) <= layer0_outputs(4215);
    layer1_outputs(423) <= (layer0_outputs(1254)) and not (layer0_outputs(1385));
    layer1_outputs(424) <= (layer0_outputs(2886)) and not (layer0_outputs(1824));
    layer1_outputs(425) <= (layer0_outputs(1986)) or (layer0_outputs(1576));
    layer1_outputs(426) <= (layer0_outputs(1461)) or (layer0_outputs(4289));
    layer1_outputs(427) <= (layer0_outputs(3059)) and (layer0_outputs(1393));
    layer1_outputs(428) <= not(layer0_outputs(3715));
    layer1_outputs(429) <= '0';
    layer1_outputs(430) <= layer0_outputs(4125);
    layer1_outputs(431) <= (layer0_outputs(4139)) and (layer0_outputs(2772));
    layer1_outputs(432) <= not(layer0_outputs(715));
    layer1_outputs(433) <= (layer0_outputs(2012)) or (layer0_outputs(492));
    layer1_outputs(434) <= not((layer0_outputs(713)) and (layer0_outputs(3535)));
    layer1_outputs(435) <= '1';
    layer1_outputs(436) <= '0';
    layer1_outputs(437) <= '0';
    layer1_outputs(438) <= '1';
    layer1_outputs(439) <= (layer0_outputs(364)) or (layer0_outputs(1162));
    layer1_outputs(440) <= not(layer0_outputs(4101));
    layer1_outputs(441) <= '1';
    layer1_outputs(442) <= '1';
    layer1_outputs(443) <= layer0_outputs(698);
    layer1_outputs(444) <= (layer0_outputs(2535)) or (layer0_outputs(4724));
    layer1_outputs(445) <= not((layer0_outputs(2039)) or (layer0_outputs(1371)));
    layer1_outputs(446) <= '1';
    layer1_outputs(447) <= (layer0_outputs(1952)) and (layer0_outputs(3958));
    layer1_outputs(448) <= (layer0_outputs(2888)) and not (layer0_outputs(1978));
    layer1_outputs(449) <= not((layer0_outputs(4815)) or (layer0_outputs(3856)));
    layer1_outputs(450) <= '1';
    layer1_outputs(451) <= not((layer0_outputs(2370)) and (layer0_outputs(3175)));
    layer1_outputs(452) <= (layer0_outputs(3355)) and (layer0_outputs(3401));
    layer1_outputs(453) <= (layer0_outputs(2054)) and (layer0_outputs(1507));
    layer1_outputs(454) <= not(layer0_outputs(3179));
    layer1_outputs(455) <= layer0_outputs(4402);
    layer1_outputs(456) <= not(layer0_outputs(4558)) or (layer0_outputs(4668));
    layer1_outputs(457) <= not(layer0_outputs(1034)) or (layer0_outputs(2468));
    layer1_outputs(458) <= (layer0_outputs(4111)) and (layer0_outputs(3144));
    layer1_outputs(459) <= not(layer0_outputs(642));
    layer1_outputs(460) <= not(layer0_outputs(3992));
    layer1_outputs(461) <= not(layer0_outputs(774));
    layer1_outputs(462) <= not((layer0_outputs(1780)) and (layer0_outputs(3657)));
    layer1_outputs(463) <= layer0_outputs(2551);
    layer1_outputs(464) <= (layer0_outputs(1404)) and not (layer0_outputs(260));
    layer1_outputs(465) <= '0';
    layer1_outputs(466) <= not(layer0_outputs(659)) or (layer0_outputs(3626));
    layer1_outputs(467) <= '1';
    layer1_outputs(468) <= (layer0_outputs(2437)) and not (layer0_outputs(3794));
    layer1_outputs(469) <= (layer0_outputs(2008)) or (layer0_outputs(2978));
    layer1_outputs(470) <= not(layer0_outputs(4292)) or (layer0_outputs(1779));
    layer1_outputs(471) <= not(layer0_outputs(4340)) or (layer0_outputs(3940));
    layer1_outputs(472) <= not((layer0_outputs(2780)) or (layer0_outputs(1131)));
    layer1_outputs(473) <= '0';
    layer1_outputs(474) <= not(layer0_outputs(2388));
    layer1_outputs(475) <= not(layer0_outputs(154));
    layer1_outputs(476) <= (layer0_outputs(4251)) xor (layer0_outputs(2917));
    layer1_outputs(477) <= (layer0_outputs(2069)) or (layer0_outputs(3403));
    layer1_outputs(478) <= '0';
    layer1_outputs(479) <= '0';
    layer1_outputs(480) <= layer0_outputs(3258);
    layer1_outputs(481) <= layer0_outputs(2984);
    layer1_outputs(482) <= '1';
    layer1_outputs(483) <= (layer0_outputs(968)) and not (layer0_outputs(4893));
    layer1_outputs(484) <= '0';
    layer1_outputs(485) <= not(layer0_outputs(2024));
    layer1_outputs(486) <= not((layer0_outputs(5089)) xor (layer0_outputs(2430)));
    layer1_outputs(487) <= (layer0_outputs(2916)) and (layer0_outputs(2697));
    layer1_outputs(488) <= (layer0_outputs(4178)) and (layer0_outputs(881));
    layer1_outputs(489) <= (layer0_outputs(3923)) or (layer0_outputs(352));
    layer1_outputs(490) <= layer0_outputs(4241);
    layer1_outputs(491) <= not(layer0_outputs(1066));
    layer1_outputs(492) <= not(layer0_outputs(2364)) or (layer0_outputs(1628));
    layer1_outputs(493) <= '0';
    layer1_outputs(494) <= not(layer0_outputs(2071)) or (layer0_outputs(1756));
    layer1_outputs(495) <= (layer0_outputs(1113)) or (layer0_outputs(1006));
    layer1_outputs(496) <= '1';
    layer1_outputs(497) <= not((layer0_outputs(1566)) and (layer0_outputs(3477)));
    layer1_outputs(498) <= (layer0_outputs(2222)) and not (layer0_outputs(2088));
    layer1_outputs(499) <= '0';
    layer1_outputs(500) <= '0';
    layer1_outputs(501) <= layer0_outputs(3595);
    layer1_outputs(502) <= not((layer0_outputs(877)) and (layer0_outputs(3881)));
    layer1_outputs(503) <= (layer0_outputs(2841)) or (layer0_outputs(3848));
    layer1_outputs(504) <= '0';
    layer1_outputs(505) <= '0';
    layer1_outputs(506) <= (layer0_outputs(1010)) or (layer0_outputs(854));
    layer1_outputs(507) <= layer0_outputs(2442);
    layer1_outputs(508) <= (layer0_outputs(2231)) and (layer0_outputs(3484));
    layer1_outputs(509) <= not(layer0_outputs(2243)) or (layer0_outputs(4045));
    layer1_outputs(510) <= not(layer0_outputs(2691));
    layer1_outputs(511) <= (layer0_outputs(3050)) and not (layer0_outputs(2100));
    layer1_outputs(512) <= not(layer0_outputs(2377)) or (layer0_outputs(598));
    layer1_outputs(513) <= not(layer0_outputs(2981));
    layer1_outputs(514) <= '0';
    layer1_outputs(515) <= not(layer0_outputs(2075));
    layer1_outputs(516) <= layer0_outputs(3265);
    layer1_outputs(517) <= layer0_outputs(2721);
    layer1_outputs(518) <= not(layer0_outputs(3213)) or (layer0_outputs(1033));
    layer1_outputs(519) <= not(layer0_outputs(1971)) or (layer0_outputs(1472));
    layer1_outputs(520) <= layer0_outputs(756);
    layer1_outputs(521) <= '0';
    layer1_outputs(522) <= layer0_outputs(408);
    layer1_outputs(523) <= '0';
    layer1_outputs(524) <= '0';
    layer1_outputs(525) <= '1';
    layer1_outputs(526) <= '0';
    layer1_outputs(527) <= (layer0_outputs(1405)) and not (layer0_outputs(2485));
    layer1_outputs(528) <= (layer0_outputs(4462)) xor (layer0_outputs(1470));
    layer1_outputs(529) <= '0';
    layer1_outputs(530) <= (layer0_outputs(3891)) and not (layer0_outputs(1981));
    layer1_outputs(531) <= layer0_outputs(2921);
    layer1_outputs(532) <= '0';
    layer1_outputs(533) <= (layer0_outputs(3572)) and (layer0_outputs(3780));
    layer1_outputs(534) <= '1';
    layer1_outputs(535) <= not(layer0_outputs(1567));
    layer1_outputs(536) <= not(layer0_outputs(2057)) or (layer0_outputs(1012));
    layer1_outputs(537) <= (layer0_outputs(4967)) or (layer0_outputs(3134));
    layer1_outputs(538) <= not(layer0_outputs(4834));
    layer1_outputs(539) <= not(layer0_outputs(2866));
    layer1_outputs(540) <= not(layer0_outputs(2355));
    layer1_outputs(541) <= layer0_outputs(940);
    layer1_outputs(542) <= '1';
    layer1_outputs(543) <= not(layer0_outputs(1278));
    layer1_outputs(544) <= not(layer0_outputs(2083));
    layer1_outputs(545) <= layer0_outputs(4191);
    layer1_outputs(546) <= not((layer0_outputs(1071)) and (layer0_outputs(2455)));
    layer1_outputs(547) <= '0';
    layer1_outputs(548) <= (layer0_outputs(839)) and not (layer0_outputs(4618));
    layer1_outputs(549) <= '1';
    layer1_outputs(550) <= not(layer0_outputs(3573)) or (layer0_outputs(1248));
    layer1_outputs(551) <= layer0_outputs(3280);
    layer1_outputs(552) <= not(layer0_outputs(2017)) or (layer0_outputs(4020));
    layer1_outputs(553) <= not(layer0_outputs(2312));
    layer1_outputs(554) <= (layer0_outputs(4386)) and (layer0_outputs(190));
    layer1_outputs(555) <= (layer0_outputs(238)) and (layer0_outputs(3659));
    layer1_outputs(556) <= layer0_outputs(2778);
    layer1_outputs(557) <= not((layer0_outputs(4645)) xor (layer0_outputs(2843)));
    layer1_outputs(558) <= layer0_outputs(3808);
    layer1_outputs(559) <= not((layer0_outputs(4874)) or (layer0_outputs(524)));
    layer1_outputs(560) <= not(layer0_outputs(1144));
    layer1_outputs(561) <= layer0_outputs(4653);
    layer1_outputs(562) <= layer0_outputs(1409);
    layer1_outputs(563) <= (layer0_outputs(2035)) and (layer0_outputs(0));
    layer1_outputs(564) <= '0';
    layer1_outputs(565) <= (layer0_outputs(4685)) or (layer0_outputs(4596));
    layer1_outputs(566) <= '1';
    layer1_outputs(567) <= layer0_outputs(3854);
    layer1_outputs(568) <= not(layer0_outputs(2549));
    layer1_outputs(569) <= not(layer0_outputs(4427));
    layer1_outputs(570) <= not((layer0_outputs(2881)) and (layer0_outputs(1732)));
    layer1_outputs(571) <= not((layer0_outputs(2384)) or (layer0_outputs(4962)));
    layer1_outputs(572) <= not(layer0_outputs(1244));
    layer1_outputs(573) <= layer0_outputs(11);
    layer1_outputs(574) <= not(layer0_outputs(1505)) or (layer0_outputs(3884));
    layer1_outputs(575) <= not((layer0_outputs(3205)) and (layer0_outputs(634)));
    layer1_outputs(576) <= not((layer0_outputs(3676)) xor (layer0_outputs(4646)));
    layer1_outputs(577) <= layer0_outputs(3839);
    layer1_outputs(578) <= not((layer0_outputs(3439)) or (layer0_outputs(271)));
    layer1_outputs(579) <= not(layer0_outputs(1607));
    layer1_outputs(580) <= '0';
    layer1_outputs(581) <= (layer0_outputs(894)) or (layer0_outputs(3263));
    layer1_outputs(582) <= '1';
    layer1_outputs(583) <= '0';
    layer1_outputs(584) <= (layer0_outputs(624)) and not (layer0_outputs(231));
    layer1_outputs(585) <= layer0_outputs(914);
    layer1_outputs(586) <= not(layer0_outputs(2122));
    layer1_outputs(587) <= not((layer0_outputs(1300)) and (layer0_outputs(5018)));
    layer1_outputs(588) <= not(layer0_outputs(1731));
    layer1_outputs(589) <= (layer0_outputs(2488)) and not (layer0_outputs(1192));
    layer1_outputs(590) <= (layer0_outputs(2883)) and not (layer0_outputs(1809));
    layer1_outputs(591) <= not((layer0_outputs(3789)) or (layer0_outputs(53)));
    layer1_outputs(592) <= not(layer0_outputs(1885)) or (layer0_outputs(208));
    layer1_outputs(593) <= (layer0_outputs(362)) and not (layer0_outputs(1323));
    layer1_outputs(594) <= (layer0_outputs(4002)) and not (layer0_outputs(3204));
    layer1_outputs(595) <= not(layer0_outputs(2731));
    layer1_outputs(596) <= (layer0_outputs(2979)) and (layer0_outputs(4438));
    layer1_outputs(597) <= (layer0_outputs(3067)) and not (layer0_outputs(777));
    layer1_outputs(598) <= not(layer0_outputs(641));
    layer1_outputs(599) <= (layer0_outputs(671)) and (layer0_outputs(2331));
    layer1_outputs(600) <= (layer0_outputs(2059)) and not (layer0_outputs(2000));
    layer1_outputs(601) <= layer0_outputs(1520);
    layer1_outputs(602) <= layer0_outputs(1306);
    layer1_outputs(603) <= (layer0_outputs(2349)) or (layer0_outputs(3686));
    layer1_outputs(604) <= not((layer0_outputs(2867)) or (layer0_outputs(2502)));
    layer1_outputs(605) <= (layer0_outputs(451)) and not (layer0_outputs(786));
    layer1_outputs(606) <= (layer0_outputs(1528)) or (layer0_outputs(1476));
    layer1_outputs(607) <= '1';
    layer1_outputs(608) <= '1';
    layer1_outputs(609) <= not(layer0_outputs(4602)) or (layer0_outputs(2109));
    layer1_outputs(610) <= not(layer0_outputs(2840));
    layer1_outputs(611) <= not(layer0_outputs(652)) or (layer0_outputs(2647));
    layer1_outputs(612) <= (layer0_outputs(2236)) and not (layer0_outputs(2714));
    layer1_outputs(613) <= layer0_outputs(825);
    layer1_outputs(614) <= (layer0_outputs(765)) and not (layer0_outputs(4811));
    layer1_outputs(615) <= not(layer0_outputs(508));
    layer1_outputs(616) <= layer0_outputs(3435);
    layer1_outputs(617) <= (layer0_outputs(251)) and not (layer0_outputs(4063));
    layer1_outputs(618) <= not(layer0_outputs(3770)) or (layer0_outputs(920));
    layer1_outputs(619) <= (layer0_outputs(4607)) and (layer0_outputs(3934));
    layer1_outputs(620) <= not((layer0_outputs(4903)) or (layer0_outputs(4716)));
    layer1_outputs(621) <= not((layer0_outputs(4335)) xor (layer0_outputs(3450)));
    layer1_outputs(622) <= '0';
    layer1_outputs(623) <= '1';
    layer1_outputs(624) <= not((layer0_outputs(2575)) and (layer0_outputs(2508)));
    layer1_outputs(625) <= (layer0_outputs(3444)) and not (layer0_outputs(2326));
    layer1_outputs(626) <= (layer0_outputs(3085)) and (layer0_outputs(1242));
    layer1_outputs(627) <= (layer0_outputs(3149)) and not (layer0_outputs(2642));
    layer1_outputs(628) <= not(layer0_outputs(1923)) or (layer0_outputs(3498));
    layer1_outputs(629) <= not(layer0_outputs(660)) or (layer0_outputs(978));
    layer1_outputs(630) <= layer0_outputs(2123);
    layer1_outputs(631) <= not((layer0_outputs(4005)) xor (layer0_outputs(870)));
    layer1_outputs(632) <= not((layer0_outputs(5036)) and (layer0_outputs(562)));
    layer1_outputs(633) <= (layer0_outputs(3737)) and (layer0_outputs(3554));
    layer1_outputs(634) <= not(layer0_outputs(5109)) or (layer0_outputs(2629));
    layer1_outputs(635) <= not(layer0_outputs(4371)) or (layer0_outputs(488));
    layer1_outputs(636) <= (layer0_outputs(1361)) and (layer0_outputs(1805));
    layer1_outputs(637) <= (layer0_outputs(2500)) and (layer0_outputs(1030));
    layer1_outputs(638) <= '1';
    layer1_outputs(639) <= layer0_outputs(2520);
    layer1_outputs(640) <= not(layer0_outputs(4960)) or (layer0_outputs(1668));
    layer1_outputs(641) <= '1';
    layer1_outputs(642) <= layer0_outputs(5030);
    layer1_outputs(643) <= not(layer0_outputs(4923));
    layer1_outputs(644) <= not((layer0_outputs(4112)) and (layer0_outputs(3470)));
    layer1_outputs(645) <= '0';
    layer1_outputs(646) <= layer0_outputs(1751);
    layer1_outputs(647) <= not(layer0_outputs(2607));
    layer1_outputs(648) <= layer0_outputs(4592);
    layer1_outputs(649) <= not(layer0_outputs(743));
    layer1_outputs(650) <= not(layer0_outputs(775)) or (layer0_outputs(1738));
    layer1_outputs(651) <= (layer0_outputs(4498)) xor (layer0_outputs(3537));
    layer1_outputs(652) <= not((layer0_outputs(1148)) and (layer0_outputs(5111)));
    layer1_outputs(653) <= not(layer0_outputs(4359));
    layer1_outputs(654) <= not((layer0_outputs(3888)) and (layer0_outputs(2106)));
    layer1_outputs(655) <= (layer0_outputs(161)) and not (layer0_outputs(3882));
    layer1_outputs(656) <= not(layer0_outputs(3165)) or (layer0_outputs(1571));
    layer1_outputs(657) <= (layer0_outputs(2773)) and (layer0_outputs(802));
    layer1_outputs(658) <= '0';
    layer1_outputs(659) <= not((layer0_outputs(3163)) and (layer0_outputs(5102)));
    layer1_outputs(660) <= not(layer0_outputs(258));
    layer1_outputs(661) <= not((layer0_outputs(5045)) and (layer0_outputs(1590)));
    layer1_outputs(662) <= not((layer0_outputs(3502)) xor (layer0_outputs(3258)));
    layer1_outputs(663) <= (layer0_outputs(3962)) and not (layer0_outputs(2691));
    layer1_outputs(664) <= not(layer0_outputs(1598));
    layer1_outputs(665) <= not((layer0_outputs(1938)) and (layer0_outputs(3510)));
    layer1_outputs(666) <= '1';
    layer1_outputs(667) <= not(layer0_outputs(836)) or (layer0_outputs(4104));
    layer1_outputs(668) <= not(layer0_outputs(4263));
    layer1_outputs(669) <= (layer0_outputs(156)) or (layer0_outputs(3063));
    layer1_outputs(670) <= not((layer0_outputs(2974)) or (layer0_outputs(4606)));
    layer1_outputs(671) <= layer0_outputs(41);
    layer1_outputs(672) <= '0';
    layer1_outputs(673) <= layer0_outputs(4110);
    layer1_outputs(674) <= layer0_outputs(4428);
    layer1_outputs(675) <= (layer0_outputs(2610)) and not (layer0_outputs(3289));
    layer1_outputs(676) <= not(layer0_outputs(5035));
    layer1_outputs(677) <= not(layer0_outputs(3022)) or (layer0_outputs(814));
    layer1_outputs(678) <= (layer0_outputs(621)) and (layer0_outputs(312));
    layer1_outputs(679) <= not(layer0_outputs(3391)) or (layer0_outputs(2810));
    layer1_outputs(680) <= not(layer0_outputs(4387));
    layer1_outputs(681) <= (layer0_outputs(2630)) or (layer0_outputs(1480));
    layer1_outputs(682) <= not(layer0_outputs(605)) or (layer0_outputs(2626));
    layer1_outputs(683) <= '1';
    layer1_outputs(684) <= (layer0_outputs(273)) and not (layer0_outputs(4878));
    layer1_outputs(685) <= '1';
    layer1_outputs(686) <= not(layer0_outputs(4332));
    layer1_outputs(687) <= '1';
    layer1_outputs(688) <= layer0_outputs(2307);
    layer1_outputs(689) <= not(layer0_outputs(3543));
    layer1_outputs(690) <= not(layer0_outputs(1790)) or (layer0_outputs(4053));
    layer1_outputs(691) <= '0';
    layer1_outputs(692) <= not(layer0_outputs(716));
    layer1_outputs(693) <= (layer0_outputs(838)) and not (layer0_outputs(4495));
    layer1_outputs(694) <= (layer0_outputs(1664)) and (layer0_outputs(4471));
    layer1_outputs(695) <= (layer0_outputs(2017)) and not (layer0_outputs(2108));
    layer1_outputs(696) <= layer0_outputs(3485);
    layer1_outputs(697) <= not(layer0_outputs(3894));
    layer1_outputs(698) <= layer0_outputs(3909);
    layer1_outputs(699) <= not(layer0_outputs(1103));
    layer1_outputs(700) <= (layer0_outputs(3049)) and (layer0_outputs(108));
    layer1_outputs(701) <= '1';
    layer1_outputs(702) <= not((layer0_outputs(4040)) and (layer0_outputs(3503)));
    layer1_outputs(703) <= (layer0_outputs(3190)) and not (layer0_outputs(3871));
    layer1_outputs(704) <= (layer0_outputs(1207)) and (layer0_outputs(4254));
    layer1_outputs(705) <= not(layer0_outputs(499)) or (layer0_outputs(119));
    layer1_outputs(706) <= '0';
    layer1_outputs(707) <= (layer0_outputs(1634)) and (layer0_outputs(3782));
    layer1_outputs(708) <= not(layer0_outputs(1394)) or (layer0_outputs(4323));
    layer1_outputs(709) <= not(layer0_outputs(3275)) or (layer0_outputs(2351));
    layer1_outputs(710) <= not(layer0_outputs(4226));
    layer1_outputs(711) <= not(layer0_outputs(3884));
    layer1_outputs(712) <= not(layer0_outputs(1812)) or (layer0_outputs(2552));
    layer1_outputs(713) <= not((layer0_outputs(1441)) or (layer0_outputs(1619)));
    layer1_outputs(714) <= '1';
    layer1_outputs(715) <= '0';
    layer1_outputs(716) <= '1';
    layer1_outputs(717) <= (layer0_outputs(1576)) or (layer0_outputs(1819));
    layer1_outputs(718) <= not((layer0_outputs(1194)) and (layer0_outputs(1488)));
    layer1_outputs(719) <= not((layer0_outputs(3128)) and (layer0_outputs(4404)));
    layer1_outputs(720) <= '1';
    layer1_outputs(721) <= not(layer0_outputs(3969)) or (layer0_outputs(3377));
    layer1_outputs(722) <= (layer0_outputs(3078)) and not (layer0_outputs(2191));
    layer1_outputs(723) <= not(layer0_outputs(4658)) or (layer0_outputs(1999));
    layer1_outputs(724) <= '0';
    layer1_outputs(725) <= (layer0_outputs(3578)) and (layer0_outputs(3324));
    layer1_outputs(726) <= not((layer0_outputs(4354)) or (layer0_outputs(1167)));
    layer1_outputs(727) <= (layer0_outputs(278)) and (layer0_outputs(3248));
    layer1_outputs(728) <= not((layer0_outputs(3386)) or (layer0_outputs(298)));
    layer1_outputs(729) <= '1';
    layer1_outputs(730) <= layer0_outputs(387);
    layer1_outputs(731) <= (layer0_outputs(3670)) and not (layer0_outputs(3623));
    layer1_outputs(732) <= (layer0_outputs(4458)) and not (layer0_outputs(4812));
    layer1_outputs(733) <= (layer0_outputs(3911)) and not (layer0_outputs(114));
    layer1_outputs(734) <= '0';
    layer1_outputs(735) <= not(layer0_outputs(2734)) or (layer0_outputs(2628));
    layer1_outputs(736) <= not(layer0_outputs(1425));
    layer1_outputs(737) <= not(layer0_outputs(585));
    layer1_outputs(738) <= (layer0_outputs(5083)) and not (layer0_outputs(4496));
    layer1_outputs(739) <= (layer0_outputs(2695)) and (layer0_outputs(1139));
    layer1_outputs(740) <= layer0_outputs(1839);
    layer1_outputs(741) <= layer0_outputs(2903);
    layer1_outputs(742) <= not(layer0_outputs(449));
    layer1_outputs(743) <= layer0_outputs(2983);
    layer1_outputs(744) <= layer0_outputs(4862);
    layer1_outputs(745) <= layer0_outputs(4872);
    layer1_outputs(746) <= layer0_outputs(845);
    layer1_outputs(747) <= not(layer0_outputs(32));
    layer1_outputs(748) <= (layer0_outputs(3773)) or (layer0_outputs(4316));
    layer1_outputs(749) <= layer0_outputs(1942);
    layer1_outputs(750) <= not(layer0_outputs(2980));
    layer1_outputs(751) <= '0';
    layer1_outputs(752) <= layer0_outputs(3040);
    layer1_outputs(753) <= not(layer0_outputs(3250));
    layer1_outputs(754) <= layer0_outputs(2264);
    layer1_outputs(755) <= (layer0_outputs(2964)) or (layer0_outputs(3442));
    layer1_outputs(756) <= layer0_outputs(993);
    layer1_outputs(757) <= not(layer0_outputs(3348));
    layer1_outputs(758) <= not(layer0_outputs(2910)) or (layer0_outputs(847));
    layer1_outputs(759) <= '1';
    layer1_outputs(760) <= '1';
    layer1_outputs(761) <= not(layer0_outputs(1500));
    layer1_outputs(762) <= (layer0_outputs(4935)) and not (layer0_outputs(1081));
    layer1_outputs(763) <= not(layer0_outputs(4248));
    layer1_outputs(764) <= '0';
    layer1_outputs(765) <= not((layer0_outputs(4041)) or (layer0_outputs(3557)));
    layer1_outputs(766) <= '0';
    layer1_outputs(767) <= layer0_outputs(3940);
    layer1_outputs(768) <= layer0_outputs(1268);
    layer1_outputs(769) <= not(layer0_outputs(1019)) or (layer0_outputs(1943));
    layer1_outputs(770) <= not(layer0_outputs(889));
    layer1_outputs(771) <= '0';
    layer1_outputs(772) <= '0';
    layer1_outputs(773) <= (layer0_outputs(2413)) or (layer0_outputs(1342));
    layer1_outputs(774) <= '0';
    layer1_outputs(775) <= layer0_outputs(4615);
    layer1_outputs(776) <= (layer0_outputs(3345)) and not (layer0_outputs(3404));
    layer1_outputs(777) <= (layer0_outputs(3723)) and (layer0_outputs(2146));
    layer1_outputs(778) <= not(layer0_outputs(1338)) or (layer0_outputs(5007));
    layer1_outputs(779) <= not(layer0_outputs(4389)) or (layer0_outputs(2278));
    layer1_outputs(780) <= (layer0_outputs(1500)) and not (layer0_outputs(4191));
    layer1_outputs(781) <= not(layer0_outputs(189));
    layer1_outputs(782) <= (layer0_outputs(2588)) and (layer0_outputs(1088));
    layer1_outputs(783) <= '0';
    layer1_outputs(784) <= '1';
    layer1_outputs(785) <= not(layer0_outputs(1745));
    layer1_outputs(786) <= not(layer0_outputs(1534));
    layer1_outputs(787) <= '1';
    layer1_outputs(788) <= layer0_outputs(2407);
    layer1_outputs(789) <= '1';
    layer1_outputs(790) <= not(layer0_outputs(3996));
    layer1_outputs(791) <= not((layer0_outputs(3037)) and (layer0_outputs(4333)));
    layer1_outputs(792) <= layer0_outputs(4681);
    layer1_outputs(793) <= not(layer0_outputs(1557));
    layer1_outputs(794) <= not((layer0_outputs(2021)) and (layer0_outputs(2962)));
    layer1_outputs(795) <= '0';
    layer1_outputs(796) <= not((layer0_outputs(3020)) or (layer0_outputs(356)));
    layer1_outputs(797) <= (layer0_outputs(3938)) or (layer0_outputs(2770));
    layer1_outputs(798) <= not(layer0_outputs(3391)) or (layer0_outputs(4119));
    layer1_outputs(799) <= '1';
    layer1_outputs(800) <= (layer0_outputs(4617)) and not (layer0_outputs(3189));
    layer1_outputs(801) <= '1';
    layer1_outputs(802) <= (layer0_outputs(49)) and not (layer0_outputs(4649));
    layer1_outputs(803) <= (layer0_outputs(773)) or (layer0_outputs(3942));
    layer1_outputs(804) <= layer0_outputs(4637);
    layer1_outputs(805) <= (layer0_outputs(3334)) and (layer0_outputs(2332));
    layer1_outputs(806) <= not((layer0_outputs(1609)) or (layer0_outputs(1937)));
    layer1_outputs(807) <= layer0_outputs(4030);
    layer1_outputs(808) <= layer0_outputs(1928);
    layer1_outputs(809) <= (layer0_outputs(618)) and not (layer0_outputs(1708));
    layer1_outputs(810) <= not((layer0_outputs(835)) and (layer0_outputs(2826)));
    layer1_outputs(811) <= (layer0_outputs(2995)) and (layer0_outputs(4957));
    layer1_outputs(812) <= layer0_outputs(2387);
    layer1_outputs(813) <= not(layer0_outputs(4315));
    layer1_outputs(814) <= (layer0_outputs(2248)) and not (layer0_outputs(2786));
    layer1_outputs(815) <= '0';
    layer1_outputs(816) <= not((layer0_outputs(4650)) and (layer0_outputs(1041)));
    layer1_outputs(817) <= (layer0_outputs(286)) and not (layer0_outputs(5023));
    layer1_outputs(818) <= '0';
    layer1_outputs(819) <= not(layer0_outputs(4349)) or (layer0_outputs(4852));
    layer1_outputs(820) <= (layer0_outputs(2018)) and (layer0_outputs(3617));
    layer1_outputs(821) <= (layer0_outputs(594)) and not (layer0_outputs(4755));
    layer1_outputs(822) <= (layer0_outputs(693)) xor (layer0_outputs(2197));
    layer1_outputs(823) <= not(layer0_outputs(4130)) or (layer0_outputs(1513));
    layer1_outputs(824) <= (layer0_outputs(477)) and not (layer0_outputs(3434));
    layer1_outputs(825) <= (layer0_outputs(239)) and not (layer0_outputs(715));
    layer1_outputs(826) <= (layer0_outputs(1731)) and not (layer0_outputs(1015));
    layer1_outputs(827) <= '0';
    layer1_outputs(828) <= not(layer0_outputs(473));
    layer1_outputs(829) <= layer0_outputs(3109);
    layer1_outputs(830) <= '0';
    layer1_outputs(831) <= (layer0_outputs(2939)) and not (layer0_outputs(4867));
    layer1_outputs(832) <= '0';
    layer1_outputs(833) <= '1';
    layer1_outputs(834) <= (layer0_outputs(1527)) or (layer0_outputs(1803));
    layer1_outputs(835) <= (layer0_outputs(3304)) and not (layer0_outputs(650));
    layer1_outputs(836) <= (layer0_outputs(220)) and not (layer0_outputs(1332));
    layer1_outputs(837) <= (layer0_outputs(952)) and not (layer0_outputs(3928));
    layer1_outputs(838) <= not(layer0_outputs(3572));
    layer1_outputs(839) <= not(layer0_outputs(4879));
    layer1_outputs(840) <= not((layer0_outputs(5119)) and (layer0_outputs(2797)));
    layer1_outputs(841) <= not(layer0_outputs(4460)) or (layer0_outputs(1713));
    layer1_outputs(842) <= '0';
    layer1_outputs(843) <= '0';
    layer1_outputs(844) <= (layer0_outputs(2645)) and not (layer0_outputs(4812));
    layer1_outputs(845) <= not(layer0_outputs(4525));
    layer1_outputs(846) <= not(layer0_outputs(2717));
    layer1_outputs(847) <= '0';
    layer1_outputs(848) <= (layer0_outputs(4918)) and (layer0_outputs(1330));
    layer1_outputs(849) <= '0';
    layer1_outputs(850) <= not((layer0_outputs(558)) and (layer0_outputs(1912)));
    layer1_outputs(851) <= (layer0_outputs(3905)) and (layer0_outputs(581));
    layer1_outputs(852) <= (layer0_outputs(1154)) or (layer0_outputs(4996));
    layer1_outputs(853) <= (layer0_outputs(2942)) and not (layer0_outputs(3328));
    layer1_outputs(854) <= not(layer0_outputs(2174)) or (layer0_outputs(158));
    layer1_outputs(855) <= (layer0_outputs(3744)) and not (layer0_outputs(3121));
    layer1_outputs(856) <= '1';
    layer1_outputs(857) <= layer0_outputs(4846);
    layer1_outputs(858) <= (layer0_outputs(5072)) or (layer0_outputs(12));
    layer1_outputs(859) <= (layer0_outputs(2769)) and not (layer0_outputs(2260));
    layer1_outputs(860) <= not(layer0_outputs(1911)) or (layer0_outputs(2327));
    layer1_outputs(861) <= layer0_outputs(2424);
    layer1_outputs(862) <= '1';
    layer1_outputs(863) <= layer0_outputs(2394);
    layer1_outputs(864) <= not((layer0_outputs(4754)) or (layer0_outputs(4452)));
    layer1_outputs(865) <= not(layer0_outputs(1697)) or (layer0_outputs(4731));
    layer1_outputs(866) <= not(layer0_outputs(1257)) or (layer0_outputs(4351));
    layer1_outputs(867) <= '1';
    layer1_outputs(868) <= not(layer0_outputs(1875));
    layer1_outputs(869) <= layer0_outputs(4565);
    layer1_outputs(870) <= not(layer0_outputs(3116)) or (layer0_outputs(2466));
    layer1_outputs(871) <= not(layer0_outputs(879)) or (layer0_outputs(2509));
    layer1_outputs(872) <= not((layer0_outputs(2223)) or (layer0_outputs(736)));
    layer1_outputs(873) <= not((layer0_outputs(1192)) or (layer0_outputs(5033)));
    layer1_outputs(874) <= '1';
    layer1_outputs(875) <= not(layer0_outputs(3731)) or (layer0_outputs(2016));
    layer1_outputs(876) <= layer0_outputs(4671);
    layer1_outputs(877) <= (layer0_outputs(1804)) and not (layer0_outputs(2764));
    layer1_outputs(878) <= not((layer0_outputs(670)) or (layer0_outputs(3059)));
    layer1_outputs(879) <= '1';
    layer1_outputs(880) <= (layer0_outputs(4966)) and not (layer0_outputs(4209));
    layer1_outputs(881) <= layer0_outputs(4268);
    layer1_outputs(882) <= layer0_outputs(3396);
    layer1_outputs(883) <= (layer0_outputs(2986)) and (layer0_outputs(2025));
    layer1_outputs(884) <= not((layer0_outputs(2389)) and (layer0_outputs(90)));
    layer1_outputs(885) <= (layer0_outputs(1071)) and not (layer0_outputs(4707));
    layer1_outputs(886) <= (layer0_outputs(1370)) and (layer0_outputs(2051));
    layer1_outputs(887) <= not((layer0_outputs(4899)) and (layer0_outputs(3278)));
    layer1_outputs(888) <= not(layer0_outputs(2747)) or (layer0_outputs(2827));
    layer1_outputs(889) <= (layer0_outputs(3287)) and not (layer0_outputs(4636));
    layer1_outputs(890) <= (layer0_outputs(93)) and (layer0_outputs(1564));
    layer1_outputs(891) <= (layer0_outputs(804)) and (layer0_outputs(1902));
    layer1_outputs(892) <= not(layer0_outputs(2927)) or (layer0_outputs(1679));
    layer1_outputs(893) <= not((layer0_outputs(945)) and (layer0_outputs(2640)));
    layer1_outputs(894) <= layer0_outputs(4418);
    layer1_outputs(895) <= not((layer0_outputs(2543)) or (layer0_outputs(2290)));
    layer1_outputs(896) <= '0';
    layer1_outputs(897) <= not(layer0_outputs(4720));
    layer1_outputs(898) <= '1';
    layer1_outputs(899) <= '1';
    layer1_outputs(900) <= not((layer0_outputs(2791)) and (layer0_outputs(4943)));
    layer1_outputs(901) <= (layer0_outputs(29)) and not (layer0_outputs(1093));
    layer1_outputs(902) <= not((layer0_outputs(619)) and (layer0_outputs(1418)));
    layer1_outputs(903) <= '1';
    layer1_outputs(904) <= '0';
    layer1_outputs(905) <= (layer0_outputs(4467)) and not (layer0_outputs(4620));
    layer1_outputs(906) <= (layer0_outputs(3375)) and not (layer0_outputs(3759));
    layer1_outputs(907) <= (layer0_outputs(4395)) or (layer0_outputs(3680));
    layer1_outputs(908) <= not(layer0_outputs(479));
    layer1_outputs(909) <= '1';
    layer1_outputs(910) <= not(layer0_outputs(1499)) or (layer0_outputs(3368));
    layer1_outputs(911) <= not(layer0_outputs(5));
    layer1_outputs(912) <= not(layer0_outputs(3392));
    layer1_outputs(913) <= layer0_outputs(3242);
    layer1_outputs(914) <= layer0_outputs(1560);
    layer1_outputs(915) <= not(layer0_outputs(3684));
    layer1_outputs(916) <= not((layer0_outputs(4448)) and (layer0_outputs(505)));
    layer1_outputs(917) <= not(layer0_outputs(4228));
    layer1_outputs(918) <= layer0_outputs(455);
    layer1_outputs(919) <= '0';
    layer1_outputs(920) <= (layer0_outputs(4913)) and not (layer0_outputs(5115));
    layer1_outputs(921) <= not(layer0_outputs(4304));
    layer1_outputs(922) <= '0';
    layer1_outputs(923) <= layer0_outputs(1248);
    layer1_outputs(924) <= (layer0_outputs(2694)) and not (layer0_outputs(3848));
    layer1_outputs(925) <= not((layer0_outputs(2438)) and (layer0_outputs(1421)));
    layer1_outputs(926) <= '1';
    layer1_outputs(927) <= (layer0_outputs(2420)) and not (layer0_outputs(3900));
    layer1_outputs(928) <= (layer0_outputs(2750)) and (layer0_outputs(1926));
    layer1_outputs(929) <= not(layer0_outputs(607)) or (layer0_outputs(1271));
    layer1_outputs(930) <= (layer0_outputs(2567)) and not (layer0_outputs(5110));
    layer1_outputs(931) <= not((layer0_outputs(2912)) xor (layer0_outputs(4181)));
    layer1_outputs(932) <= not(layer0_outputs(3455)) or (layer0_outputs(1094));
    layer1_outputs(933) <= '1';
    layer1_outputs(934) <= '0';
    layer1_outputs(935) <= layer0_outputs(4132);
    layer1_outputs(936) <= layer0_outputs(203);
    layer1_outputs(937) <= not(layer0_outputs(1358));
    layer1_outputs(938) <= '1';
    layer1_outputs(939) <= layer0_outputs(4089);
    layer1_outputs(940) <= layer0_outputs(5054);
    layer1_outputs(941) <= not(layer0_outputs(2130));
    layer1_outputs(942) <= not(layer0_outputs(4809)) or (layer0_outputs(2286));
    layer1_outputs(943) <= (layer0_outputs(2761)) and not (layer0_outputs(1222));
    layer1_outputs(944) <= not(layer0_outputs(1091));
    layer1_outputs(945) <= '1';
    layer1_outputs(946) <= layer0_outputs(2038);
    layer1_outputs(947) <= (layer0_outputs(1335)) and (layer0_outputs(726));
    layer1_outputs(948) <= (layer0_outputs(8)) and not (layer0_outputs(4160));
    layer1_outputs(949) <= (layer0_outputs(2714)) and not (layer0_outputs(2505));
    layer1_outputs(950) <= layer0_outputs(2836);
    layer1_outputs(951) <= '0';
    layer1_outputs(952) <= not((layer0_outputs(2273)) or (layer0_outputs(2569)));
    layer1_outputs(953) <= layer0_outputs(383);
    layer1_outputs(954) <= (layer0_outputs(3330)) and (layer0_outputs(2359));
    layer1_outputs(955) <= not(layer0_outputs(3708)) or (layer0_outputs(1277));
    layer1_outputs(956) <= (layer0_outputs(3120)) and not (layer0_outputs(2596));
    layer1_outputs(957) <= (layer0_outputs(3759)) and (layer0_outputs(4760));
    layer1_outputs(958) <= not(layer0_outputs(4590));
    layer1_outputs(959) <= not(layer0_outputs(647));
    layer1_outputs(960) <= not((layer0_outputs(1100)) or (layer0_outputs(369)));
    layer1_outputs(961) <= not((layer0_outputs(4997)) xor (layer0_outputs(1801)));
    layer1_outputs(962) <= layer0_outputs(412);
    layer1_outputs(963) <= '0';
    layer1_outputs(964) <= '1';
    layer1_outputs(965) <= (layer0_outputs(2916)) and (layer0_outputs(1674));
    layer1_outputs(966) <= not(layer0_outputs(5017)) or (layer0_outputs(3806));
    layer1_outputs(967) <= not(layer0_outputs(3393));
    layer1_outputs(968) <= not(layer0_outputs(707));
    layer1_outputs(969) <= (layer0_outputs(3504)) and not (layer0_outputs(3141));
    layer1_outputs(970) <= not(layer0_outputs(4768));
    layer1_outputs(971) <= not(layer0_outputs(2988));
    layer1_outputs(972) <= not((layer0_outputs(617)) or (layer0_outputs(4907)));
    layer1_outputs(973) <= (layer0_outputs(1710)) and (layer0_outputs(2804));
    layer1_outputs(974) <= not(layer0_outputs(277));
    layer1_outputs(975) <= (layer0_outputs(2028)) or (layer0_outputs(732));
    layer1_outputs(976) <= (layer0_outputs(679)) or (layer0_outputs(1858));
    layer1_outputs(977) <= (layer0_outputs(853)) and not (layer0_outputs(5004));
    layer1_outputs(978) <= not(layer0_outputs(1189));
    layer1_outputs(979) <= (layer0_outputs(790)) and not (layer0_outputs(3106));
    layer1_outputs(980) <= '0';
    layer1_outputs(981) <= (layer0_outputs(4542)) and not (layer0_outputs(526));
    layer1_outputs(982) <= '0';
    layer1_outputs(983) <= not(layer0_outputs(4473)) or (layer0_outputs(2687));
    layer1_outputs(984) <= layer0_outputs(204);
    layer1_outputs(985) <= (layer0_outputs(1739)) and not (layer0_outputs(36));
    layer1_outputs(986) <= layer0_outputs(2216);
    layer1_outputs(987) <= layer0_outputs(3920);
    layer1_outputs(988) <= not(layer0_outputs(536));
    layer1_outputs(989) <= layer0_outputs(2069);
    layer1_outputs(990) <= layer0_outputs(165);
    layer1_outputs(991) <= not(layer0_outputs(4359));
    layer1_outputs(992) <= not(layer0_outputs(2817)) or (layer0_outputs(1227));
    layer1_outputs(993) <= (layer0_outputs(4297)) and not (layer0_outputs(2978));
    layer1_outputs(994) <= (layer0_outputs(2141)) and (layer0_outputs(2974));
    layer1_outputs(995) <= not(layer0_outputs(3775)) or (layer0_outputs(1650));
    layer1_outputs(996) <= not(layer0_outputs(976)) or (layer0_outputs(3886));
    layer1_outputs(997) <= '1';
    layer1_outputs(998) <= not(layer0_outputs(2673));
    layer1_outputs(999) <= (layer0_outputs(2708)) and not (layer0_outputs(3035));
    layer1_outputs(1000) <= not(layer0_outputs(1177)) or (layer0_outputs(3758));
    layer1_outputs(1001) <= (layer0_outputs(3569)) and not (layer0_outputs(735));
    layer1_outputs(1002) <= not((layer0_outputs(4212)) or (layer0_outputs(4227)));
    layer1_outputs(1003) <= (layer0_outputs(430)) and (layer0_outputs(1777));
    layer1_outputs(1004) <= not(layer0_outputs(2324)) or (layer0_outputs(4311));
    layer1_outputs(1005) <= (layer0_outputs(2297)) and not (layer0_outputs(2211));
    layer1_outputs(1006) <= not(layer0_outputs(1321));
    layer1_outputs(1007) <= (layer0_outputs(3092)) and not (layer0_outputs(795));
    layer1_outputs(1008) <= not(layer0_outputs(503));
    layer1_outputs(1009) <= not(layer0_outputs(502)) or (layer0_outputs(1449));
    layer1_outputs(1010) <= not(layer0_outputs(3410));
    layer1_outputs(1011) <= '1';
    layer1_outputs(1012) <= '1';
    layer1_outputs(1013) <= layer0_outputs(779);
    layer1_outputs(1014) <= (layer0_outputs(3656)) and not (layer0_outputs(3394));
    layer1_outputs(1015) <= layer0_outputs(4057);
    layer1_outputs(1016) <= layer0_outputs(564);
    layer1_outputs(1017) <= not(layer0_outputs(170));
    layer1_outputs(1018) <= (layer0_outputs(805)) and not (layer0_outputs(3466));
    layer1_outputs(1019) <= not((layer0_outputs(3459)) xor (layer0_outputs(2012)));
    layer1_outputs(1020) <= not(layer0_outputs(2165)) or (layer0_outputs(1100));
    layer1_outputs(1021) <= (layer0_outputs(288)) and (layer0_outputs(4818));
    layer1_outputs(1022) <= (layer0_outputs(1151)) or (layer0_outputs(2304));
    layer1_outputs(1023) <= not(layer0_outputs(3613));
    layer1_outputs(1024) <= '0';
    layer1_outputs(1025) <= (layer0_outputs(136)) and not (layer0_outputs(3445));
    layer1_outputs(1026) <= (layer0_outputs(987)) and (layer0_outputs(3881));
    layer1_outputs(1027) <= not(layer0_outputs(3925)) or (layer0_outputs(4481));
    layer1_outputs(1028) <= (layer0_outputs(89)) or (layer0_outputs(3774));
    layer1_outputs(1029) <= '0';
    layer1_outputs(1030) <= (layer0_outputs(4278)) or (layer0_outputs(1231));
    layer1_outputs(1031) <= layer0_outputs(1434);
    layer1_outputs(1032) <= not((layer0_outputs(4597)) and (layer0_outputs(4981)));
    layer1_outputs(1033) <= not(layer0_outputs(2762)) or (layer0_outputs(1814));
    layer1_outputs(1034) <= (layer0_outputs(1004)) or (layer0_outputs(1539));
    layer1_outputs(1035) <= layer0_outputs(792);
    layer1_outputs(1036) <= '1';
    layer1_outputs(1037) <= (layer0_outputs(4018)) and not (layer0_outputs(3393));
    layer1_outputs(1038) <= not(layer0_outputs(25)) or (layer0_outputs(277));
    layer1_outputs(1039) <= not(layer0_outputs(3614)) or (layer0_outputs(3872));
    layer1_outputs(1040) <= not(layer0_outputs(3753)) or (layer0_outputs(77));
    layer1_outputs(1041) <= (layer0_outputs(3598)) or (layer0_outputs(2764));
    layer1_outputs(1042) <= '0';
    layer1_outputs(1043) <= not((layer0_outputs(3869)) and (layer0_outputs(1497)));
    layer1_outputs(1044) <= not(layer0_outputs(5080)) or (layer0_outputs(4079));
    layer1_outputs(1045) <= (layer0_outputs(199)) and (layer0_outputs(818));
    layer1_outputs(1046) <= not(layer0_outputs(706)) or (layer0_outputs(3588));
    layer1_outputs(1047) <= not(layer0_outputs(2676)) or (layer0_outputs(3219));
    layer1_outputs(1048) <= layer0_outputs(191);
    layer1_outputs(1049) <= '0';
    layer1_outputs(1050) <= not(layer0_outputs(2131));
    layer1_outputs(1051) <= not(layer0_outputs(4958));
    layer1_outputs(1052) <= not(layer0_outputs(1905)) or (layer0_outputs(1982));
    layer1_outputs(1053) <= not(layer0_outputs(1917));
    layer1_outputs(1054) <= not(layer0_outputs(1108)) or (layer0_outputs(4593));
    layer1_outputs(1055) <= not((layer0_outputs(3507)) and (layer0_outputs(2151)));
    layer1_outputs(1056) <= (layer0_outputs(2683)) and (layer0_outputs(3657));
    layer1_outputs(1057) <= not((layer0_outputs(2617)) xor (layer0_outputs(4232)));
    layer1_outputs(1058) <= not(layer0_outputs(2308)) or (layer0_outputs(1276));
    layer1_outputs(1059) <= layer0_outputs(4692);
    layer1_outputs(1060) <= (layer0_outputs(3319)) and (layer0_outputs(383));
    layer1_outputs(1061) <= not((layer0_outputs(2063)) and (layer0_outputs(3729)));
    layer1_outputs(1062) <= '1';
    layer1_outputs(1063) <= (layer0_outputs(942)) and not (layer0_outputs(2228));
    layer1_outputs(1064) <= (layer0_outputs(4476)) and (layer0_outputs(3364));
    layer1_outputs(1065) <= '1';
    layer1_outputs(1066) <= not((layer0_outputs(2492)) xor (layer0_outputs(1435)));
    layer1_outputs(1067) <= (layer0_outputs(4022)) or (layer0_outputs(3901));
    layer1_outputs(1068) <= '1';
    layer1_outputs(1069) <= '1';
    layer1_outputs(1070) <= (layer0_outputs(4172)) and not (layer0_outputs(3250));
    layer1_outputs(1071) <= (layer0_outputs(2066)) and (layer0_outputs(3142));
    layer1_outputs(1072) <= not(layer0_outputs(2684));
    layer1_outputs(1073) <= (layer0_outputs(3661)) and (layer0_outputs(34));
    layer1_outputs(1074) <= (layer0_outputs(1123)) or (layer0_outputs(3041));
    layer1_outputs(1075) <= '1';
    layer1_outputs(1076) <= '0';
    layer1_outputs(1077) <= not(layer0_outputs(4526)) or (layer0_outputs(2217));
    layer1_outputs(1078) <= '1';
    layer1_outputs(1079) <= (layer0_outputs(141)) and (layer0_outputs(506));
    layer1_outputs(1080) <= layer0_outputs(608);
    layer1_outputs(1081) <= (layer0_outputs(4742)) and not (layer0_outputs(2067));
    layer1_outputs(1082) <= not((layer0_outputs(3766)) or (layer0_outputs(4969)));
    layer1_outputs(1083) <= not((layer0_outputs(3359)) and (layer0_outputs(3075)));
    layer1_outputs(1084) <= not((layer0_outputs(1477)) and (layer0_outputs(462)));
    layer1_outputs(1085) <= (layer0_outputs(1776)) and (layer0_outputs(3427));
    layer1_outputs(1086) <= (layer0_outputs(2745)) and (layer0_outputs(3268));
    layer1_outputs(1087) <= layer0_outputs(443);
    layer1_outputs(1088) <= not(layer0_outputs(1471)) or (layer0_outputs(2253));
    layer1_outputs(1089) <= not(layer0_outputs(2009));
    layer1_outputs(1090) <= not((layer0_outputs(2458)) or (layer0_outputs(1961)));
    layer1_outputs(1091) <= '0';
    layer1_outputs(1092) <= (layer0_outputs(2554)) xor (layer0_outputs(2936));
    layer1_outputs(1093) <= not(layer0_outputs(3101)) or (layer0_outputs(3184));
    layer1_outputs(1094) <= '1';
    layer1_outputs(1095) <= not(layer0_outputs(2019));
    layer1_outputs(1096) <= '0';
    layer1_outputs(1097) <= '1';
    layer1_outputs(1098) <= not(layer0_outputs(3767));
    layer1_outputs(1099) <= layer0_outputs(1088);
    layer1_outputs(1100) <= '0';
    layer1_outputs(1101) <= not(layer0_outputs(1309)) or (layer0_outputs(2270));
    layer1_outputs(1102) <= (layer0_outputs(4693)) and not (layer0_outputs(3214));
    layer1_outputs(1103) <= '0';
    layer1_outputs(1104) <= '1';
    layer1_outputs(1105) <= layer0_outputs(4914);
    layer1_outputs(1106) <= not(layer0_outputs(2884));
    layer1_outputs(1107) <= layer0_outputs(1237);
    layer1_outputs(1108) <= not(layer0_outputs(3842));
    layer1_outputs(1109) <= '1';
    layer1_outputs(1110) <= not(layer0_outputs(4176)) or (layer0_outputs(476));
    layer1_outputs(1111) <= not((layer0_outputs(4440)) or (layer0_outputs(557)));
    layer1_outputs(1112) <= '0';
    layer1_outputs(1113) <= (layer0_outputs(3287)) and not (layer0_outputs(3079));
    layer1_outputs(1114) <= not((layer0_outputs(4414)) and (layer0_outputs(4647)));
    layer1_outputs(1115) <= '0';
    layer1_outputs(1116) <= layer0_outputs(89);
    layer1_outputs(1117) <= layer0_outputs(3151);
    layer1_outputs(1118) <= layer0_outputs(1208);
    layer1_outputs(1119) <= not((layer0_outputs(3389)) or (layer0_outputs(3506)));
    layer1_outputs(1120) <= not(layer0_outputs(283)) or (layer0_outputs(3286));
    layer1_outputs(1121) <= (layer0_outputs(3422)) and not (layer0_outputs(2310));
    layer1_outputs(1122) <= not((layer0_outputs(1282)) and (layer0_outputs(2213)));
    layer1_outputs(1123) <= (layer0_outputs(3744)) and (layer0_outputs(1106));
    layer1_outputs(1124) <= not(layer0_outputs(1819)) or (layer0_outputs(2969));
    layer1_outputs(1125) <= (layer0_outputs(3722)) and not (layer0_outputs(2736));
    layer1_outputs(1126) <= (layer0_outputs(552)) and (layer0_outputs(222));
    layer1_outputs(1127) <= not((layer0_outputs(4708)) and (layer0_outputs(3454)));
    layer1_outputs(1128) <= (layer0_outputs(4712)) or (layer0_outputs(3253));
    layer1_outputs(1129) <= not((layer0_outputs(575)) or (layer0_outputs(4229)));
    layer1_outputs(1130) <= not(layer0_outputs(1084));
    layer1_outputs(1131) <= '0';
    layer1_outputs(1132) <= (layer0_outputs(3667)) and not (layer0_outputs(598));
    layer1_outputs(1133) <= (layer0_outputs(3357)) and not (layer0_outputs(535));
    layer1_outputs(1134) <= (layer0_outputs(3223)) and not (layer0_outputs(142));
    layer1_outputs(1135) <= not(layer0_outputs(2329));
    layer1_outputs(1136) <= '1';
    layer1_outputs(1137) <= not((layer0_outputs(4136)) or (layer0_outputs(4744)));
    layer1_outputs(1138) <= '0';
    layer1_outputs(1139) <= (layer0_outputs(2161)) and not (layer0_outputs(2091));
    layer1_outputs(1140) <= not((layer0_outputs(2457)) and (layer0_outputs(4124)));
    layer1_outputs(1141) <= not(layer0_outputs(4633)) or (layer0_outputs(3106));
    layer1_outputs(1142) <= not((layer0_outputs(2814)) or (layer0_outputs(2)));
    layer1_outputs(1143) <= not(layer0_outputs(4260)) or (layer0_outputs(4619));
    layer1_outputs(1144) <= (layer0_outputs(3346)) and not (layer0_outputs(1176));
    layer1_outputs(1145) <= (layer0_outputs(4503)) or (layer0_outputs(4244));
    layer1_outputs(1146) <= not(layer0_outputs(975)) or (layer0_outputs(4397));
    layer1_outputs(1147) <= layer0_outputs(2646);
    layer1_outputs(1148) <= not(layer0_outputs(547));
    layer1_outputs(1149) <= not(layer0_outputs(521)) or (layer0_outputs(2725));
    layer1_outputs(1150) <= not(layer0_outputs(1237)) or (layer0_outputs(2609));
    layer1_outputs(1151) <= not(layer0_outputs(4301)) or (layer0_outputs(3448));
    layer1_outputs(1152) <= (layer0_outputs(4529)) and not (layer0_outputs(4700));
    layer1_outputs(1153) <= not((layer0_outputs(999)) or (layer0_outputs(1259)));
    layer1_outputs(1154) <= (layer0_outputs(2333)) or (layer0_outputs(1870));
    layer1_outputs(1155) <= (layer0_outputs(2500)) xor (layer0_outputs(1518));
    layer1_outputs(1156) <= (layer0_outputs(1788)) and not (layer0_outputs(1989));
    layer1_outputs(1157) <= (layer0_outputs(3481)) xor (layer0_outputs(2585));
    layer1_outputs(1158) <= not(layer0_outputs(3590));
    layer1_outputs(1159) <= '0';
    layer1_outputs(1160) <= not(layer0_outputs(4149));
    layer1_outputs(1161) <= layer0_outputs(88);
    layer1_outputs(1162) <= (layer0_outputs(1943)) or (layer0_outputs(495));
    layer1_outputs(1163) <= '0';
    layer1_outputs(1164) <= not((layer0_outputs(3321)) and (layer0_outputs(2157)));
    layer1_outputs(1165) <= '0';
    layer1_outputs(1166) <= '1';
    layer1_outputs(1167) <= '0';
    layer1_outputs(1168) <= (layer0_outputs(973)) and not (layer0_outputs(4258));
    layer1_outputs(1169) <= '1';
    layer1_outputs(1170) <= (layer0_outputs(1482)) or (layer0_outputs(3380));
    layer1_outputs(1171) <= layer0_outputs(2903);
    layer1_outputs(1172) <= layer0_outputs(3752);
    layer1_outputs(1173) <= (layer0_outputs(2176)) and not (layer0_outputs(4890));
    layer1_outputs(1174) <= not(layer0_outputs(4975));
    layer1_outputs(1175) <= not(layer0_outputs(1947));
    layer1_outputs(1176) <= not(layer0_outputs(4955)) or (layer0_outputs(1939));
    layer1_outputs(1177) <= '1';
    layer1_outputs(1178) <= '1';
    layer1_outputs(1179) <= (layer0_outputs(4383)) and not (layer0_outputs(1729));
    layer1_outputs(1180) <= not(layer0_outputs(1930));
    layer1_outputs(1181) <= not(layer0_outputs(3964));
    layer1_outputs(1182) <= layer0_outputs(1520);
    layer1_outputs(1183) <= '0';
    layer1_outputs(1184) <= '1';
    layer1_outputs(1185) <= not(layer0_outputs(361));
    layer1_outputs(1186) <= not((layer0_outputs(902)) or (layer0_outputs(4273)));
    layer1_outputs(1187) <= (layer0_outputs(1693)) and not (layer0_outputs(4014));
    layer1_outputs(1188) <= (layer0_outputs(2132)) and not (layer0_outputs(2276));
    layer1_outputs(1189) <= not((layer0_outputs(1189)) or (layer0_outputs(4720)));
    layer1_outputs(1190) <= (layer0_outputs(1784)) or (layer0_outputs(2305));
    layer1_outputs(1191) <= not((layer0_outputs(1161)) and (layer0_outputs(4854)));
    layer1_outputs(1192) <= (layer0_outputs(2358)) or (layer0_outputs(1673));
    layer1_outputs(1193) <= layer0_outputs(4142);
    layer1_outputs(1194) <= layer0_outputs(46);
    layer1_outputs(1195) <= layer0_outputs(3479);
    layer1_outputs(1196) <= '0';
    layer1_outputs(1197) <= not((layer0_outputs(3634)) and (layer0_outputs(4930)));
    layer1_outputs(1198) <= layer0_outputs(4773);
    layer1_outputs(1199) <= (layer0_outputs(3513)) xor (layer0_outputs(988));
    layer1_outputs(1200) <= (layer0_outputs(4270)) and (layer0_outputs(2257));
    layer1_outputs(1201) <= not(layer0_outputs(4781));
    layer1_outputs(1202) <= not(layer0_outputs(4108)) or (layer0_outputs(225));
    layer1_outputs(1203) <= not((layer0_outputs(2899)) or (layer0_outputs(3814)));
    layer1_outputs(1204) <= '1';
    layer1_outputs(1205) <= layer0_outputs(3872);
    layer1_outputs(1206) <= not((layer0_outputs(1878)) or (layer0_outputs(1154)));
    layer1_outputs(1207) <= '1';
    layer1_outputs(1208) <= (layer0_outputs(3780)) and (layer0_outputs(3773));
    layer1_outputs(1209) <= layer0_outputs(1603);
    layer1_outputs(1210) <= (layer0_outputs(2860)) or (layer0_outputs(4452));
    layer1_outputs(1211) <= (layer0_outputs(1306)) or (layer0_outputs(895));
    layer1_outputs(1212) <= (layer0_outputs(1157)) and not (layer0_outputs(2240));
    layer1_outputs(1213) <= (layer0_outputs(463)) or (layer0_outputs(345));
    layer1_outputs(1214) <= not((layer0_outputs(4512)) or (layer0_outputs(4518)));
    layer1_outputs(1215) <= (layer0_outputs(5051)) or (layer0_outputs(1672));
    layer1_outputs(1216) <= layer0_outputs(110);
    layer1_outputs(1217) <= (layer0_outputs(3930)) and (layer0_outputs(4201));
    layer1_outputs(1218) <= layer0_outputs(2002);
    layer1_outputs(1219) <= layer0_outputs(3587);
    layer1_outputs(1220) <= not((layer0_outputs(1621)) and (layer0_outputs(2032)));
    layer1_outputs(1221) <= '1';
    layer1_outputs(1222) <= layer0_outputs(3574);
    layer1_outputs(1223) <= not(layer0_outputs(1263));
    layer1_outputs(1224) <= layer0_outputs(3714);
    layer1_outputs(1225) <= '1';
    layer1_outputs(1226) <= not(layer0_outputs(2168)) or (layer0_outputs(4509));
    layer1_outputs(1227) <= layer0_outputs(4672);
    layer1_outputs(1228) <= (layer0_outputs(3688)) and not (layer0_outputs(3408));
    layer1_outputs(1229) <= (layer0_outputs(1933)) and not (layer0_outputs(522));
    layer1_outputs(1230) <= not(layer0_outputs(4964));
    layer1_outputs(1231) <= not(layer0_outputs(2381)) or (layer0_outputs(3739));
    layer1_outputs(1232) <= not(layer0_outputs(3562));
    layer1_outputs(1233) <= (layer0_outputs(2540)) and not (layer0_outputs(1279));
    layer1_outputs(1234) <= not(layer0_outputs(2932));
    layer1_outputs(1235) <= layer0_outputs(4607);
    layer1_outputs(1236) <= layer0_outputs(1620);
    layer1_outputs(1237) <= not(layer0_outputs(3609));
    layer1_outputs(1238) <= layer0_outputs(695);
    layer1_outputs(1239) <= '1';
    layer1_outputs(1240) <= (layer0_outputs(1590)) xor (layer0_outputs(3843));
    layer1_outputs(1241) <= not((layer0_outputs(1115)) and (layer0_outputs(2426)));
    layer1_outputs(1242) <= not(layer0_outputs(4492));
    layer1_outputs(1243) <= not((layer0_outputs(1670)) xor (layer0_outputs(3927)));
    layer1_outputs(1244) <= not((layer0_outputs(4038)) and (layer0_outputs(1147)));
    layer1_outputs(1245) <= not((layer0_outputs(3876)) or (layer0_outputs(1387)));
    layer1_outputs(1246) <= (layer0_outputs(3899)) and (layer0_outputs(1080));
    layer1_outputs(1247) <= not((layer0_outputs(245)) and (layer0_outputs(391)));
    layer1_outputs(1248) <= not((layer0_outputs(2190)) or (layer0_outputs(1734)));
    layer1_outputs(1249) <= not(layer0_outputs(1439)) or (layer0_outputs(1395));
    layer1_outputs(1250) <= '1';
    layer1_outputs(1251) <= not(layer0_outputs(4203)) or (layer0_outputs(2367));
    layer1_outputs(1252) <= not(layer0_outputs(1850));
    layer1_outputs(1253) <= not((layer0_outputs(606)) xor (layer0_outputs(4838)));
    layer1_outputs(1254) <= (layer0_outputs(3043)) or (layer0_outputs(2700));
    layer1_outputs(1255) <= (layer0_outputs(1442)) and not (layer0_outputs(1461));
    layer1_outputs(1256) <= not((layer0_outputs(2331)) or (layer0_outputs(3610)));
    layer1_outputs(1257) <= '1';
    layer1_outputs(1258) <= not(layer0_outputs(1881));
    layer1_outputs(1259) <= (layer0_outputs(3028)) xor (layer0_outputs(262));
    layer1_outputs(1260) <= not(layer0_outputs(1833)) or (layer0_outputs(2172));
    layer1_outputs(1261) <= layer0_outputs(3208);
    layer1_outputs(1262) <= (layer0_outputs(429)) and not (layer0_outputs(541));
    layer1_outputs(1263) <= not(layer0_outputs(4644)) or (layer0_outputs(787));
    layer1_outputs(1264) <= not((layer0_outputs(943)) and (layer0_outputs(167)));
    layer1_outputs(1265) <= layer0_outputs(714);
    layer1_outputs(1266) <= not(layer0_outputs(4234));
    layer1_outputs(1267) <= '1';
    layer1_outputs(1268) <= (layer0_outputs(4982)) and (layer0_outputs(2263));
    layer1_outputs(1269) <= not(layer0_outputs(1649));
    layer1_outputs(1270) <= not(layer0_outputs(852));
    layer1_outputs(1271) <= not(layer0_outputs(147));
    layer1_outputs(1272) <= '0';
    layer1_outputs(1273) <= not(layer0_outputs(153)) or (layer0_outputs(4649));
    layer1_outputs(1274) <= (layer0_outputs(1743)) and (layer0_outputs(2855));
    layer1_outputs(1275) <= layer0_outputs(2008);
    layer1_outputs(1276) <= (layer0_outputs(1130)) and not (layer0_outputs(270));
    layer1_outputs(1277) <= not(layer0_outputs(2119)) or (layer0_outputs(4999));
    layer1_outputs(1278) <= (layer0_outputs(2339)) xor (layer0_outputs(1622));
    layer1_outputs(1279) <= layer0_outputs(3569);
    layer1_outputs(1280) <= not(layer0_outputs(4491));
    layer1_outputs(1281) <= (layer0_outputs(5092)) and (layer0_outputs(2467));
    layer1_outputs(1282) <= '0';
    layer1_outputs(1283) <= layer0_outputs(144);
    layer1_outputs(1284) <= not((layer0_outputs(4918)) and (layer0_outputs(3398)));
    layer1_outputs(1285) <= not(layer0_outputs(1132)) or (layer0_outputs(4824));
    layer1_outputs(1286) <= (layer0_outputs(1663)) and not (layer0_outputs(2677));
    layer1_outputs(1287) <= (layer0_outputs(1199)) and not (layer0_outputs(257));
    layer1_outputs(1288) <= not(layer0_outputs(3145));
    layer1_outputs(1289) <= '0';
    layer1_outputs(1290) <= layer0_outputs(1955);
    layer1_outputs(1291) <= not((layer0_outputs(3955)) or (layer0_outputs(2463)));
    layer1_outputs(1292) <= layer0_outputs(3109);
    layer1_outputs(1293) <= not((layer0_outputs(3584)) and (layer0_outputs(5010)));
    layer1_outputs(1294) <= layer0_outputs(1724);
    layer1_outputs(1295) <= layer0_outputs(3021);
    layer1_outputs(1296) <= not((layer0_outputs(2915)) or (layer0_outputs(3492)));
    layer1_outputs(1297) <= '1';
    layer1_outputs(1298) <= not(layer0_outputs(4913));
    layer1_outputs(1299) <= not(layer0_outputs(1323));
    layer1_outputs(1300) <= layer0_outputs(1905);
    layer1_outputs(1301) <= not(layer0_outputs(1402));
    layer1_outputs(1302) <= not(layer0_outputs(4152));
    layer1_outputs(1303) <= '1';
    layer1_outputs(1304) <= not((layer0_outputs(380)) and (layer0_outputs(3267)));
    layer1_outputs(1305) <= '0';
    layer1_outputs(1306) <= (layer0_outputs(931)) or (layer0_outputs(4992));
    layer1_outputs(1307) <= layer0_outputs(3820);
    layer1_outputs(1308) <= not(layer0_outputs(4019));
    layer1_outputs(1309) <= (layer0_outputs(4114)) and not (layer0_outputs(626));
    layer1_outputs(1310) <= '1';
    layer1_outputs(1311) <= (layer0_outputs(498)) and not (layer0_outputs(2639));
    layer1_outputs(1312) <= '1';
    layer1_outputs(1313) <= not(layer0_outputs(2319));
    layer1_outputs(1314) <= not((layer0_outputs(1519)) or (layer0_outputs(2777)));
    layer1_outputs(1315) <= not((layer0_outputs(195)) and (layer0_outputs(3108)));
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= (layer0_outputs(3761)) and not (layer0_outputs(3047));
    layer1_outputs(1318) <= (layer0_outputs(2187)) or (layer0_outputs(3103));
    layer1_outputs(1319) <= '0';
    layer1_outputs(1320) <= not(layer0_outputs(2843));
    layer1_outputs(1321) <= '1';
    layer1_outputs(1322) <= not(layer0_outputs(4798));
    layer1_outputs(1323) <= '1';
    layer1_outputs(1324) <= not(layer0_outputs(3282));
    layer1_outputs(1325) <= not((layer0_outputs(936)) and (layer0_outputs(1191)));
    layer1_outputs(1326) <= '1';
    layer1_outputs(1327) <= (layer0_outputs(4285)) and not (layer0_outputs(3443));
    layer1_outputs(1328) <= not(layer0_outputs(2975));
    layer1_outputs(1329) <= layer0_outputs(4409);
    layer1_outputs(1330) <= (layer0_outputs(1480)) or (layer0_outputs(445));
    layer1_outputs(1331) <= not(layer0_outputs(679)) or (layer0_outputs(1601));
    layer1_outputs(1332) <= layer0_outputs(2891);
    layer1_outputs(1333) <= layer0_outputs(3090);
    layer1_outputs(1334) <= layer0_outputs(533);
    layer1_outputs(1335) <= '1';
    layer1_outputs(1336) <= '1';
    layer1_outputs(1337) <= not((layer0_outputs(1719)) xor (layer0_outputs(3520)));
    layer1_outputs(1338) <= not(layer0_outputs(2513)) or (layer0_outputs(1725));
    layer1_outputs(1339) <= layer0_outputs(3396);
    layer1_outputs(1340) <= not(layer0_outputs(4057));
    layer1_outputs(1341) <= not(layer0_outputs(4746));
    layer1_outputs(1342) <= layer0_outputs(2918);
    layer1_outputs(1343) <= layer0_outputs(1567);
    layer1_outputs(1344) <= not(layer0_outputs(3599));
    layer1_outputs(1345) <= (layer0_outputs(4365)) and (layer0_outputs(880));
    layer1_outputs(1346) <= (layer0_outputs(2791)) and not (layer0_outputs(2812));
    layer1_outputs(1347) <= not((layer0_outputs(990)) or (layer0_outputs(4369)));
    layer1_outputs(1348) <= layer0_outputs(1261);
    layer1_outputs(1349) <= (layer0_outputs(4941)) and not (layer0_outputs(340));
    layer1_outputs(1350) <= not(layer0_outputs(3445));
    layer1_outputs(1351) <= not(layer0_outputs(2407));
    layer1_outputs(1352) <= not(layer0_outputs(267));
    layer1_outputs(1353) <= (layer0_outputs(1927)) and not (layer0_outputs(3053));
    layer1_outputs(1354) <= not(layer0_outputs(2816));
    layer1_outputs(1355) <= (layer0_outputs(2115)) and not (layer0_outputs(1269));
    layer1_outputs(1356) <= (layer0_outputs(1165)) and not (layer0_outputs(4873));
    layer1_outputs(1357) <= (layer0_outputs(3822)) xor (layer0_outputs(104));
    layer1_outputs(1358) <= (layer0_outputs(340)) or (layer0_outputs(2041));
    layer1_outputs(1359) <= '0';
    layer1_outputs(1360) <= layer0_outputs(5081);
    layer1_outputs(1361) <= layer0_outputs(1234);
    layer1_outputs(1362) <= not(layer0_outputs(4143));
    layer1_outputs(1363) <= layer0_outputs(590);
    layer1_outputs(1364) <= (layer0_outputs(3102)) and not (layer0_outputs(2578));
    layer1_outputs(1365) <= not((layer0_outputs(3860)) and (layer0_outputs(742)));
    layer1_outputs(1366) <= '0';
    layer1_outputs(1367) <= not(layer0_outputs(4193)) or (layer0_outputs(544));
    layer1_outputs(1368) <= not(layer0_outputs(734)) or (layer0_outputs(1655));
    layer1_outputs(1369) <= (layer0_outputs(4169)) or (layer0_outputs(1715));
    layer1_outputs(1370) <= not((layer0_outputs(1473)) xor (layer0_outputs(315)));
    layer1_outputs(1371) <= layer0_outputs(739);
    layer1_outputs(1372) <= '0';
    layer1_outputs(1373) <= '1';
    layer1_outputs(1374) <= (layer0_outputs(4261)) and (layer0_outputs(5052));
    layer1_outputs(1375) <= (layer0_outputs(4621)) or (layer0_outputs(2744));
    layer1_outputs(1376) <= (layer0_outputs(4579)) and (layer0_outputs(1452));
    layer1_outputs(1377) <= '1';
    layer1_outputs(1378) <= '0';
    layer1_outputs(1379) <= '0';
    layer1_outputs(1380) <= (layer0_outputs(3743)) and (layer0_outputs(3953));
    layer1_outputs(1381) <= not(layer0_outputs(983)) or (layer0_outputs(2466));
    layer1_outputs(1382) <= not(layer0_outputs(3012)) or (layer0_outputs(4825));
    layer1_outputs(1383) <= layer0_outputs(4427);
    layer1_outputs(1384) <= not(layer0_outputs(3371)) or (layer0_outputs(4682));
    layer1_outputs(1385) <= layer0_outputs(3179);
    layer1_outputs(1386) <= not(layer0_outputs(3403));
    layer1_outputs(1387) <= layer0_outputs(1776);
    layer1_outputs(1388) <= not(layer0_outputs(3811)) or (layer0_outputs(2113));
    layer1_outputs(1389) <= layer0_outputs(1853);
    layer1_outputs(1390) <= not((layer0_outputs(3932)) or (layer0_outputs(2565)));
    layer1_outputs(1391) <= not(layer0_outputs(1410)) or (layer0_outputs(3971));
    layer1_outputs(1392) <= '0';
    layer1_outputs(1393) <= layer0_outputs(5065);
    layer1_outputs(1394) <= (layer0_outputs(3706)) and not (layer0_outputs(3476));
    layer1_outputs(1395) <= not(layer0_outputs(1090)) or (layer0_outputs(4757));
    layer1_outputs(1396) <= not(layer0_outputs(1103));
    layer1_outputs(1397) <= (layer0_outputs(66)) and (layer0_outputs(4813));
    layer1_outputs(1398) <= not(layer0_outputs(442)) or (layer0_outputs(4610));
    layer1_outputs(1399) <= '1';
    layer1_outputs(1400) <= '0';
    layer1_outputs(1401) <= layer0_outputs(515);
    layer1_outputs(1402) <= layer0_outputs(2443);
    layer1_outputs(1403) <= not(layer0_outputs(761));
    layer1_outputs(1404) <= not(layer0_outputs(848));
    layer1_outputs(1405) <= not(layer0_outputs(1451));
    layer1_outputs(1406) <= not(layer0_outputs(4384)) or (layer0_outputs(1125));
    layer1_outputs(1407) <= not(layer0_outputs(331));
    layer1_outputs(1408) <= not((layer0_outputs(4538)) xor (layer0_outputs(2688)));
    layer1_outputs(1409) <= not(layer0_outputs(684));
    layer1_outputs(1410) <= '0';
    layer1_outputs(1411) <= not(layer0_outputs(2635));
    layer1_outputs(1412) <= layer0_outputs(837);
    layer1_outputs(1413) <= layer0_outputs(4207);
    layer1_outputs(1414) <= (layer0_outputs(1986)) or (layer0_outputs(2043));
    layer1_outputs(1415) <= not((layer0_outputs(4840)) and (layer0_outputs(658)));
    layer1_outputs(1416) <= '1';
    layer1_outputs(1417) <= not((layer0_outputs(15)) or (layer0_outputs(3800)));
    layer1_outputs(1418) <= '1';
    layer1_outputs(1419) <= (layer0_outputs(3387)) and (layer0_outputs(151));
    layer1_outputs(1420) <= layer0_outputs(1762);
    layer1_outputs(1421) <= not(layer0_outputs(3989)) or (layer0_outputs(1374));
    layer1_outputs(1422) <= '1';
    layer1_outputs(1423) <= (layer0_outputs(3770)) and not (layer0_outputs(4637));
    layer1_outputs(1424) <= not((layer0_outputs(653)) or (layer0_outputs(496)));
    layer1_outputs(1425) <= '0';
    layer1_outputs(1426) <= '1';
    layer1_outputs(1427) <= not(layer0_outputs(1362));
    layer1_outputs(1428) <= not(layer0_outputs(654));
    layer1_outputs(1429) <= '1';
    layer1_outputs(1430) <= (layer0_outputs(556)) and (layer0_outputs(2493));
    layer1_outputs(1431) <= not(layer0_outputs(5011)) or (layer0_outputs(2483));
    layer1_outputs(1432) <= not(layer0_outputs(1561));
    layer1_outputs(1433) <= '0';
    layer1_outputs(1434) <= not(layer0_outputs(717)) or (layer0_outputs(4410));
    layer1_outputs(1435) <= (layer0_outputs(957)) and not (layer0_outputs(3801));
    layer1_outputs(1436) <= (layer0_outputs(3236)) and (layer0_outputs(4273));
    layer1_outputs(1437) <= not(layer0_outputs(3277));
    layer1_outputs(1438) <= (layer0_outputs(4617)) and not (layer0_outputs(3221));
    layer1_outputs(1439) <= layer0_outputs(150);
    layer1_outputs(1440) <= layer0_outputs(1832);
    layer1_outputs(1441) <= not(layer0_outputs(2240));
    layer1_outputs(1442) <= layer0_outputs(1446);
    layer1_outputs(1443) <= not((layer0_outputs(3437)) and (layer0_outputs(613)));
    layer1_outputs(1444) <= not(layer0_outputs(682)) or (layer0_outputs(3971));
    layer1_outputs(1445) <= layer0_outputs(1760);
    layer1_outputs(1446) <= (layer0_outputs(971)) and not (layer0_outputs(3904));
    layer1_outputs(1447) <= '0';
    layer1_outputs(1448) <= '0';
    layer1_outputs(1449) <= not(layer0_outputs(1326));
    layer1_outputs(1450) <= not(layer0_outputs(1667));
    layer1_outputs(1451) <= not(layer0_outputs(187)) or (layer0_outputs(3939));
    layer1_outputs(1452) <= not(layer0_outputs(2652)) or (layer0_outputs(4876));
    layer1_outputs(1453) <= not(layer0_outputs(4466)) or (layer0_outputs(4303));
    layer1_outputs(1454) <= not(layer0_outputs(4834)) or (layer0_outputs(147));
    layer1_outputs(1455) <= (layer0_outputs(3902)) and not (layer0_outputs(4563));
    layer1_outputs(1456) <= '0';
    layer1_outputs(1457) <= not((layer0_outputs(4151)) or (layer0_outputs(4447)));
    layer1_outputs(1458) <= (layer0_outputs(4550)) xor (layer0_outputs(59));
    layer1_outputs(1459) <= not((layer0_outputs(3173)) or (layer0_outputs(2645)));
    layer1_outputs(1460) <= layer0_outputs(703);
    layer1_outputs(1461) <= (layer0_outputs(2760)) and (layer0_outputs(2096));
    layer1_outputs(1462) <= (layer0_outputs(4677)) xor (layer0_outputs(2433));
    layer1_outputs(1463) <= (layer0_outputs(1631)) or (layer0_outputs(177));
    layer1_outputs(1464) <= '1';
    layer1_outputs(1465) <= '1';
    layer1_outputs(1466) <= not(layer0_outputs(1750));
    layer1_outputs(1467) <= '0';
    layer1_outputs(1468) <= '1';
    layer1_outputs(1469) <= layer0_outputs(2127);
    layer1_outputs(1470) <= not(layer0_outputs(4328)) or (layer0_outputs(1956));
    layer1_outputs(1471) <= '1';
    layer1_outputs(1472) <= '1';
    layer1_outputs(1473) <= '0';
    layer1_outputs(1474) <= '0';
    layer1_outputs(1475) <= (layer0_outputs(1811)) and (layer0_outputs(3576));
    layer1_outputs(1476) <= '1';
    layer1_outputs(1477) <= layer0_outputs(384);
    layer1_outputs(1478) <= not(layer0_outputs(1806));
    layer1_outputs(1479) <= not((layer0_outputs(2613)) and (layer0_outputs(3979)));
    layer1_outputs(1480) <= not(layer0_outputs(1717)) or (layer0_outputs(1901));
    layer1_outputs(1481) <= '1';
    layer1_outputs(1482) <= layer0_outputs(2244);
    layer1_outputs(1483) <= not((layer0_outputs(2076)) and (layer0_outputs(4314)));
    layer1_outputs(1484) <= '0';
    layer1_outputs(1485) <= (layer0_outputs(528)) and (layer0_outputs(3372));
    layer1_outputs(1486) <= not(layer0_outputs(968));
    layer1_outputs(1487) <= layer0_outputs(1150);
    layer1_outputs(1488) <= (layer0_outputs(3379)) and not (layer0_outputs(4820));
    layer1_outputs(1489) <= not(layer0_outputs(3185));
    layer1_outputs(1490) <= '0';
    layer1_outputs(1491) <= not((layer0_outputs(2202)) or (layer0_outputs(4629)));
    layer1_outputs(1492) <= not(layer0_outputs(4869)) or (layer0_outputs(4178));
    layer1_outputs(1493) <= (layer0_outputs(2335)) and (layer0_outputs(2060));
    layer1_outputs(1494) <= not(layer0_outputs(2550));
    layer1_outputs(1495) <= (layer0_outputs(1723)) or (layer0_outputs(1828));
    layer1_outputs(1496) <= not(layer0_outputs(1761));
    layer1_outputs(1497) <= layer0_outputs(1643);
    layer1_outputs(1498) <= not(layer0_outputs(4516)) or (layer0_outputs(150));
    layer1_outputs(1499) <= '1';
    layer1_outputs(1500) <= layer0_outputs(2992);
    layer1_outputs(1501) <= not((layer0_outputs(4008)) and (layer0_outputs(4012)));
    layer1_outputs(1502) <= (layer0_outputs(2930)) and (layer0_outputs(4115));
    layer1_outputs(1503) <= (layer0_outputs(2741)) and (layer0_outputs(242));
    layer1_outputs(1504) <= not((layer0_outputs(1649)) xor (layer0_outputs(1187)));
    layer1_outputs(1505) <= not(layer0_outputs(5));
    layer1_outputs(1506) <= not(layer0_outputs(4725)) or (layer0_outputs(2085));
    layer1_outputs(1507) <= (layer0_outputs(1135)) or (layer0_outputs(1722));
    layer1_outputs(1508) <= (layer0_outputs(2105)) and (layer0_outputs(8));
    layer1_outputs(1509) <= '0';
    layer1_outputs(1510) <= '0';
    layer1_outputs(1511) <= not(layer0_outputs(4130)) or (layer0_outputs(76));
    layer1_outputs(1512) <= '0';
    layer1_outputs(1513) <= '0';
    layer1_outputs(1514) <= not(layer0_outputs(2244));
    layer1_outputs(1515) <= not(layer0_outputs(842));
    layer1_outputs(1516) <= layer0_outputs(2521);
    layer1_outputs(1517) <= not(layer0_outputs(205)) or (layer0_outputs(4940));
    layer1_outputs(1518) <= '0';
    layer1_outputs(1519) <= not(layer0_outputs(2265)) or (layer0_outputs(4691));
    layer1_outputs(1520) <= not(layer0_outputs(1036));
    layer1_outputs(1521) <= '0';
    layer1_outputs(1522) <= '0';
    layer1_outputs(1523) <= not((layer0_outputs(3294)) and (layer0_outputs(2551)));
    layer1_outputs(1524) <= (layer0_outputs(3225)) and not (layer0_outputs(1823));
    layer1_outputs(1525) <= layer0_outputs(420);
    layer1_outputs(1526) <= layer0_outputs(293);
    layer1_outputs(1527) <= (layer0_outputs(1684)) and (layer0_outputs(2283));
    layer1_outputs(1528) <= not(layer0_outputs(2521));
    layer1_outputs(1529) <= not(layer0_outputs(4591)) or (layer0_outputs(1294));
    layer1_outputs(1530) <= not(layer0_outputs(3068));
    layer1_outputs(1531) <= '1';
    layer1_outputs(1532) <= '1';
    layer1_outputs(1533) <= (layer0_outputs(3786)) and (layer0_outputs(3364));
    layer1_outputs(1534) <= not(layer0_outputs(3216));
    layer1_outputs(1535) <= '0';
    layer1_outputs(1536) <= (layer0_outputs(2446)) and not (layer0_outputs(3129));
    layer1_outputs(1537) <= (layer0_outputs(2350)) and not (layer0_outputs(747));
    layer1_outputs(1538) <= not(layer0_outputs(4640));
    layer1_outputs(1539) <= not((layer0_outputs(436)) xor (layer0_outputs(3893)));
    layer1_outputs(1540) <= not((layer0_outputs(3519)) and (layer0_outputs(1494)));
    layer1_outputs(1541) <= not(layer0_outputs(1366));
    layer1_outputs(1542) <= not((layer0_outputs(1415)) or (layer0_outputs(1087)));
    layer1_outputs(1543) <= (layer0_outputs(3097)) or (layer0_outputs(2546));
    layer1_outputs(1544) <= '1';
    layer1_outputs(1545) <= '1';
    layer1_outputs(1546) <= not(layer0_outputs(2196)) or (layer0_outputs(5001));
    layer1_outputs(1547) <= not(layer0_outputs(5058)) or (layer0_outputs(3875));
    layer1_outputs(1548) <= not(layer0_outputs(3473)) or (layer0_outputs(4879));
    layer1_outputs(1549) <= not(layer0_outputs(1013));
    layer1_outputs(1550) <= layer0_outputs(673);
    layer1_outputs(1551) <= not(layer0_outputs(1898)) or (layer0_outputs(4003));
    layer1_outputs(1552) <= '1';
    layer1_outputs(1553) <= (layer0_outputs(1899)) and (layer0_outputs(2976));
    layer1_outputs(1554) <= (layer0_outputs(4559)) and (layer0_outputs(3371));
    layer1_outputs(1555) <= (layer0_outputs(4276)) and (layer0_outputs(3984));
    layer1_outputs(1556) <= (layer0_outputs(1879)) and not (layer0_outputs(3534));
    layer1_outputs(1557) <= (layer0_outputs(394)) and not (layer0_outputs(2321));
    layer1_outputs(1558) <= '0';
    layer1_outputs(1559) <= layer0_outputs(51);
    layer1_outputs(1560) <= not((layer0_outputs(527)) or (layer0_outputs(5049)));
    layer1_outputs(1561) <= (layer0_outputs(3912)) and not (layer0_outputs(3444));
    layer1_outputs(1562) <= not((layer0_outputs(1995)) or (layer0_outputs(2679)));
    layer1_outputs(1563) <= (layer0_outputs(1016)) or (layer0_outputs(3363));
    layer1_outputs(1564) <= (layer0_outputs(386)) and (layer0_outputs(949));
    layer1_outputs(1565) <= not((layer0_outputs(3024)) or (layer0_outputs(1378)));
    layer1_outputs(1566) <= '0';
    layer1_outputs(1567) <= not((layer0_outputs(2751)) and (layer0_outputs(4827)));
    layer1_outputs(1568) <= '1';
    layer1_outputs(1569) <= not((layer0_outputs(2960)) or (layer0_outputs(3096)));
    layer1_outputs(1570) <= not(layer0_outputs(214));
    layer1_outputs(1571) <= layer0_outputs(1780);
    layer1_outputs(1572) <= not(layer0_outputs(961));
    layer1_outputs(1573) <= not(layer0_outputs(4446)) or (layer0_outputs(2169));
    layer1_outputs(1574) <= not(layer0_outputs(2479));
    layer1_outputs(1575) <= '0';
    layer1_outputs(1576) <= not(layer0_outputs(1595));
    layer1_outputs(1577) <= not((layer0_outputs(4158)) and (layer0_outputs(3817)));
    layer1_outputs(1578) <= not(layer0_outputs(2677));
    layer1_outputs(1579) <= not((layer0_outputs(2351)) or (layer0_outputs(2622)));
    layer1_outputs(1580) <= not(layer0_outputs(2139)) or (layer0_outputs(398));
    layer1_outputs(1581) <= not((layer0_outputs(3064)) or (layer0_outputs(1270)));
    layer1_outputs(1582) <= (layer0_outputs(1909)) or (layer0_outputs(363));
    layer1_outputs(1583) <= not(layer0_outputs(2413));
    layer1_outputs(1584) <= not((layer0_outputs(730)) or (layer0_outputs(3094)));
    layer1_outputs(1585) <= not((layer0_outputs(4128)) and (layer0_outputs(3812)));
    layer1_outputs(1586) <= not((layer0_outputs(4153)) or (layer0_outputs(2804)));
    layer1_outputs(1587) <= not((layer0_outputs(3308)) or (layer0_outputs(3366)));
    layer1_outputs(1588) <= not(layer0_outputs(1508));
    layer1_outputs(1589) <= not(layer0_outputs(2258));
    layer1_outputs(1590) <= '0';
    layer1_outputs(1591) <= '0';
    layer1_outputs(1592) <= layer0_outputs(5015);
    layer1_outputs(1593) <= '1';
    layer1_outputs(1594) <= layer0_outputs(1964);
    layer1_outputs(1595) <= not(layer0_outputs(5119));
    layer1_outputs(1596) <= '0';
    layer1_outputs(1597) <= (layer0_outputs(3107)) or (layer0_outputs(2515));
    layer1_outputs(1598) <= not((layer0_outputs(4174)) and (layer0_outputs(686)));
    layer1_outputs(1599) <= not((layer0_outputs(1785)) and (layer0_outputs(998)));
    layer1_outputs(1600) <= layer0_outputs(1403);
    layer1_outputs(1601) <= (layer0_outputs(1717)) and not (layer0_outputs(687));
    layer1_outputs(1602) <= '0';
    layer1_outputs(1603) <= not((layer0_outputs(2121)) and (layer0_outputs(3213)));
    layer1_outputs(1604) <= layer0_outputs(3385);
    layer1_outputs(1605) <= not((layer0_outputs(1514)) and (layer0_outputs(1992)));
    layer1_outputs(1606) <= '0';
    layer1_outputs(1607) <= '0';
    layer1_outputs(1608) <= '1';
    layer1_outputs(1609) <= not(layer0_outputs(3682)) or (layer0_outputs(1216));
    layer1_outputs(1610) <= layer0_outputs(124);
    layer1_outputs(1611) <= not(layer0_outputs(2251));
    layer1_outputs(1612) <= layer0_outputs(4685);
    layer1_outputs(1613) <= '0';
    layer1_outputs(1614) <= (layer0_outputs(4096)) and not (layer0_outputs(4562));
    layer1_outputs(1615) <= (layer0_outputs(3140)) and not (layer0_outputs(2954));
    layer1_outputs(1616) <= not(layer0_outputs(1692));
    layer1_outputs(1617) <= not(layer0_outputs(4454)) or (layer0_outputs(1563));
    layer1_outputs(1618) <= '1';
    layer1_outputs(1619) <= not(layer0_outputs(2179)) or (layer0_outputs(4744));
    layer1_outputs(1620) <= '0';
    layer1_outputs(1621) <= not(layer0_outputs(2513));
    layer1_outputs(1622) <= (layer0_outputs(3925)) or (layer0_outputs(2920));
    layer1_outputs(1623) <= (layer0_outputs(57)) or (layer0_outputs(3207));
    layer1_outputs(1624) <= not(layer0_outputs(3516));
    layer1_outputs(1625) <= layer0_outputs(3295);
    layer1_outputs(1626) <= layer0_outputs(1354);
    layer1_outputs(1627) <= (layer0_outputs(1580)) and not (layer0_outputs(707));
    layer1_outputs(1628) <= (layer0_outputs(2003)) and not (layer0_outputs(4670));
    layer1_outputs(1629) <= not(layer0_outputs(4246)) or (layer0_outputs(1695));
    layer1_outputs(1630) <= '1';
    layer1_outputs(1631) <= not((layer0_outputs(62)) and (layer0_outputs(2034)));
    layer1_outputs(1632) <= not((layer0_outputs(4168)) or (layer0_outputs(440)));
    layer1_outputs(1633) <= not((layer0_outputs(4401)) and (layer0_outputs(794)));
    layer1_outputs(1634) <= (layer0_outputs(4771)) and (layer0_outputs(3209));
    layer1_outputs(1635) <= not(layer0_outputs(302));
    layer1_outputs(1636) <= not((layer0_outputs(3025)) and (layer0_outputs(1270)));
    layer1_outputs(1637) <= not(layer0_outputs(4536));
    layer1_outputs(1638) <= '0';
    layer1_outputs(1639) <= layer0_outputs(2649);
    layer1_outputs(1640) <= not((layer0_outputs(3021)) or (layer0_outputs(2806)));
    layer1_outputs(1641) <= (layer0_outputs(1029)) and not (layer0_outputs(3415));
    layer1_outputs(1642) <= not(layer0_outputs(3827));
    layer1_outputs(1643) <= not((layer0_outputs(901)) and (layer0_outputs(2781)));
    layer1_outputs(1644) <= (layer0_outputs(5023)) and not (layer0_outputs(259));
    layer1_outputs(1645) <= not(layer0_outputs(680));
    layer1_outputs(1646) <= '1';
    layer1_outputs(1647) <= layer0_outputs(2363);
    layer1_outputs(1648) <= (layer0_outputs(1512)) and not (layer0_outputs(1283));
    layer1_outputs(1649) <= (layer0_outputs(444)) or (layer0_outputs(2754));
    layer1_outputs(1650) <= not((layer0_outputs(834)) and (layer0_outputs(5101)));
    layer1_outputs(1651) <= not(layer0_outputs(4793)) or (layer0_outputs(867));
    layer1_outputs(1652) <= not((layer0_outputs(2919)) or (layer0_outputs(4362)));
    layer1_outputs(1653) <= not(layer0_outputs(3515));
    layer1_outputs(1654) <= not(layer0_outputs(4977)) or (layer0_outputs(80));
    layer1_outputs(1655) <= not(layer0_outputs(1604));
    layer1_outputs(1656) <= (layer0_outputs(655)) and (layer0_outputs(242));
    layer1_outputs(1657) <= not(layer0_outputs(2501));
    layer1_outputs(1658) <= not((layer0_outputs(5006)) and (layer0_outputs(2893)));
    layer1_outputs(1659) <= (layer0_outputs(4895)) and not (layer0_outputs(3469));
    layer1_outputs(1660) <= not(layer0_outputs(2183)) or (layer0_outputs(3285));
    layer1_outputs(1661) <= layer0_outputs(662);
    layer1_outputs(1662) <= not((layer0_outputs(3600)) and (layer0_outputs(1102)));
    layer1_outputs(1663) <= (layer0_outputs(1687)) and not (layer0_outputs(3640));
    layer1_outputs(1664) <= layer0_outputs(1701);
    layer1_outputs(1665) <= not(layer0_outputs(434));
    layer1_outputs(1666) <= not(layer0_outputs(4482));
    layer1_outputs(1667) <= layer0_outputs(486);
    layer1_outputs(1668) <= '1';
    layer1_outputs(1669) <= not(layer0_outputs(1333));
    layer1_outputs(1670) <= not((layer0_outputs(402)) or (layer0_outputs(45)));
    layer1_outputs(1671) <= not((layer0_outputs(3677)) and (layer0_outputs(1883)));
    layer1_outputs(1672) <= (layer0_outputs(4629)) and (layer0_outputs(4396));
    layer1_outputs(1673) <= (layer0_outputs(4373)) and not (layer0_outputs(940));
    layer1_outputs(1674) <= layer0_outputs(365);
    layer1_outputs(1675) <= not(layer0_outputs(2248)) or (layer0_outputs(2024));
    layer1_outputs(1676) <= (layer0_outputs(624)) and (layer0_outputs(1606));
    layer1_outputs(1677) <= layer0_outputs(4136);
    layer1_outputs(1678) <= not(layer0_outputs(382)) or (layer0_outputs(964));
    layer1_outputs(1679) <= not(layer0_outputs(401)) or (layer0_outputs(1796));
    layer1_outputs(1680) <= not(layer0_outputs(896));
    layer1_outputs(1681) <= (layer0_outputs(4939)) and not (layer0_outputs(325));
    layer1_outputs(1682) <= not(layer0_outputs(2114));
    layer1_outputs(1683) <= '0';
    layer1_outputs(1684) <= not((layer0_outputs(5008)) and (layer0_outputs(3730)));
    layer1_outputs(1685) <= (layer0_outputs(4257)) and (layer0_outputs(2013));
    layer1_outputs(1686) <= layer0_outputs(1629);
    layer1_outputs(1687) <= (layer0_outputs(5009)) and not (layer0_outputs(1719));
    layer1_outputs(1688) <= not(layer0_outputs(4401)) or (layer0_outputs(4242));
    layer1_outputs(1689) <= layer0_outputs(487);
    layer1_outputs(1690) <= (layer0_outputs(3078)) or (layer0_outputs(3429));
    layer1_outputs(1691) <= not(layer0_outputs(3017));
    layer1_outputs(1692) <= '0';
    layer1_outputs(1693) <= (layer0_outputs(4437)) and not (layer0_outputs(4998));
    layer1_outputs(1694) <= not(layer0_outputs(5100)) or (layer0_outputs(4134));
    layer1_outputs(1695) <= (layer0_outputs(2392)) and (layer0_outputs(4373));
    layer1_outputs(1696) <= layer0_outputs(3694);
    layer1_outputs(1697) <= (layer0_outputs(1877)) and not (layer0_outputs(422));
    layer1_outputs(1698) <= '0';
    layer1_outputs(1699) <= not((layer0_outputs(134)) and (layer0_outputs(2509)));
    layer1_outputs(1700) <= layer0_outputs(4392);
    layer1_outputs(1701) <= not((layer0_outputs(517)) or (layer0_outputs(3434)));
    layer1_outputs(1702) <= '1';
    layer1_outputs(1703) <= '1';
    layer1_outputs(1704) <= '1';
    layer1_outputs(1705) <= not(layer0_outputs(4564));
    layer1_outputs(1706) <= (layer0_outputs(4783)) and not (layer0_outputs(950));
    layer1_outputs(1707) <= (layer0_outputs(1798)) and not (layer0_outputs(3367));
    layer1_outputs(1708) <= '1';
    layer1_outputs(1709) <= '1';
    layer1_outputs(1710) <= not((layer0_outputs(1225)) and (layer0_outputs(2146)));
    layer1_outputs(1711) <= not((layer0_outputs(4697)) or (layer0_outputs(3313)));
    layer1_outputs(1712) <= not((layer0_outputs(3430)) or (layer0_outputs(574)));
    layer1_outputs(1713) <= '1';
    layer1_outputs(1714) <= '0';
    layer1_outputs(1715) <= '0';
    layer1_outputs(1716) <= (layer0_outputs(2470)) and (layer0_outputs(2732));
    layer1_outputs(1717) <= (layer0_outputs(3405)) and (layer0_outputs(4330));
    layer1_outputs(1718) <= not(layer0_outputs(4056)) or (layer0_outputs(1725));
    layer1_outputs(1719) <= '0';
    layer1_outputs(1720) <= '0';
    layer1_outputs(1721) <= not(layer0_outputs(1793)) or (layer0_outputs(4590));
    layer1_outputs(1722) <= not((layer0_outputs(2489)) and (layer0_outputs(1372)));
    layer1_outputs(1723) <= '0';
    layer1_outputs(1724) <= '0';
    layer1_outputs(1725) <= (layer0_outputs(975)) or (layer0_outputs(303));
    layer1_outputs(1726) <= (layer0_outputs(1083)) or (layer0_outputs(2967));
    layer1_outputs(1727) <= not(layer0_outputs(696)) or (layer0_outputs(1027));
    layer1_outputs(1728) <= '0';
    layer1_outputs(1729) <= not(layer0_outputs(1007));
    layer1_outputs(1730) <= not(layer0_outputs(351)) or (layer0_outputs(3240));
    layer1_outputs(1731) <= not(layer0_outputs(677)) or (layer0_outputs(2078));
    layer1_outputs(1732) <= not((layer0_outputs(1444)) or (layer0_outputs(592)));
    layer1_outputs(1733) <= layer0_outputs(3983);
    layer1_outputs(1734) <= (layer0_outputs(127)) or (layer0_outputs(3458));
    layer1_outputs(1735) <= (layer0_outputs(1671)) or (layer0_outputs(4716));
    layer1_outputs(1736) <= (layer0_outputs(4916)) and not (layer0_outputs(3515));
    layer1_outputs(1737) <= not((layer0_outputs(909)) or (layer0_outputs(3039)));
    layer1_outputs(1738) <= layer0_outputs(3802);
    layer1_outputs(1739) <= '1';
    layer1_outputs(1740) <= layer0_outputs(904);
    layer1_outputs(1741) <= not(layer0_outputs(2658));
    layer1_outputs(1742) <= '0';
    layer1_outputs(1743) <= '0';
    layer1_outputs(1744) <= not(layer0_outputs(620)) or (layer0_outputs(4585));
    layer1_outputs(1745) <= layer0_outputs(1613);
    layer1_outputs(1746) <= not(layer0_outputs(2338));
    layer1_outputs(1747) <= '0';
    layer1_outputs(1748) <= not((layer0_outputs(1206)) and (layer0_outputs(3799)));
    layer1_outputs(1749) <= not(layer0_outputs(295));
    layer1_outputs(1750) <= (layer0_outputs(4870)) and (layer0_outputs(4721));
    layer1_outputs(1751) <= layer0_outputs(72);
    layer1_outputs(1752) <= not(layer0_outputs(3034)) or (layer0_outputs(374));
    layer1_outputs(1753) <= not(layer0_outputs(3665));
    layer1_outputs(1754) <= (layer0_outputs(4387)) and not (layer0_outputs(3025));
    layer1_outputs(1755) <= not(layer0_outputs(2858));
    layer1_outputs(1756) <= '0';
    layer1_outputs(1757) <= (layer0_outputs(4611)) xor (layer0_outputs(4678));
    layer1_outputs(1758) <= '0';
    layer1_outputs(1759) <= not(layer0_outputs(3037));
    layer1_outputs(1760) <= '1';
    layer1_outputs(1761) <= layer0_outputs(3679);
    layer1_outputs(1762) <= not(layer0_outputs(1825)) or (layer0_outputs(4946));
    layer1_outputs(1763) <= layer0_outputs(3718);
    layer1_outputs(1764) <= '0';
    layer1_outputs(1765) <= layer0_outputs(4342);
    layer1_outputs(1766) <= not(layer0_outputs(3943)) or (layer0_outputs(2436));
    layer1_outputs(1767) <= (layer0_outputs(3299)) and (layer0_outputs(2356));
    layer1_outputs(1768) <= not(layer0_outputs(3256)) or (layer0_outputs(2284));
    layer1_outputs(1769) <= '0';
    layer1_outputs(1770) <= not(layer0_outputs(3983)) or (layer0_outputs(2245));
    layer1_outputs(1771) <= '0';
    layer1_outputs(1772) <= (layer0_outputs(3875)) and not (layer0_outputs(4966));
    layer1_outputs(1773) <= layer0_outputs(2944);
    layer1_outputs(1774) <= '0';
    layer1_outputs(1775) <= not(layer0_outputs(3697)) or (layer0_outputs(1393));
    layer1_outputs(1776) <= (layer0_outputs(2755)) and not (layer0_outputs(115));
    layer1_outputs(1777) <= layer0_outputs(3172);
    layer1_outputs(1778) <= (layer0_outputs(5050)) and (layer0_outputs(4803));
    layer1_outputs(1779) <= layer0_outputs(3607);
    layer1_outputs(1780) <= (layer0_outputs(763)) and not (layer0_outputs(1315));
    layer1_outputs(1781) <= not((layer0_outputs(3762)) and (layer0_outputs(2547)));
    layer1_outputs(1782) <= layer0_outputs(566);
    layer1_outputs(1783) <= not(layer0_outputs(73)) or (layer0_outputs(1874));
    layer1_outputs(1784) <= (layer0_outputs(1934)) and not (layer0_outputs(3010));
    layer1_outputs(1785) <= not(layer0_outputs(3804));
    layer1_outputs(1786) <= '1';
    layer1_outputs(1787) <= layer0_outputs(400);
    layer1_outputs(1788) <= not((layer0_outputs(1498)) or (layer0_outputs(5078)));
    layer1_outputs(1789) <= layer0_outputs(812);
    layer1_outputs(1790) <= not(layer0_outputs(4095)) or (layer0_outputs(2913));
    layer1_outputs(1791) <= not(layer0_outputs(10)) or (layer0_outputs(473));
    layer1_outputs(1792) <= '1';
    layer1_outputs(1793) <= (layer0_outputs(2525)) and not (layer0_outputs(1638));
    layer1_outputs(1794) <= (layer0_outputs(341)) and (layer0_outputs(3138));
    layer1_outputs(1795) <= not(layer0_outputs(304)) or (layer0_outputs(4633));
    layer1_outputs(1796) <= layer0_outputs(460);
    layer1_outputs(1797) <= '0';
    layer1_outputs(1798) <= not(layer0_outputs(4210)) or (layer0_outputs(4932));
    layer1_outputs(1799) <= (layer0_outputs(2719)) and (layer0_outputs(1666));
    layer1_outputs(1800) <= '0';
    layer1_outputs(1801) <= layer0_outputs(2685);
    layer1_outputs(1802) <= '1';
    layer1_outputs(1803) <= not((layer0_outputs(2534)) and (layer0_outputs(1936)));
    layer1_outputs(1804) <= (layer0_outputs(4318)) and (layer0_outputs(1632));
    layer1_outputs(1805) <= '0';
    layer1_outputs(1806) <= layer0_outputs(4830);
    layer1_outputs(1807) <= layer0_outputs(382);
    layer1_outputs(1808) <= not(layer0_outputs(1134));
    layer1_outputs(1809) <= (layer0_outputs(1110)) and not (layer0_outputs(2311));
    layer1_outputs(1810) <= (layer0_outputs(3511)) xor (layer0_outputs(3647));
    layer1_outputs(1811) <= layer0_outputs(1236);
    layer1_outputs(1812) <= not(layer0_outputs(4388)) or (layer0_outputs(1639));
    layer1_outputs(1813) <= not((layer0_outputs(284)) and (layer0_outputs(2494)));
    layer1_outputs(1814) <= '0';
    layer1_outputs(1815) <= (layer0_outputs(2506)) and not (layer0_outputs(3544));
    layer1_outputs(1816) <= '1';
    layer1_outputs(1817) <= not(layer0_outputs(3915)) or (layer0_outputs(551));
    layer1_outputs(1818) <= not((layer0_outputs(2846)) and (layer0_outputs(2204)));
    layer1_outputs(1819) <= '0';
    layer1_outputs(1820) <= (layer0_outputs(4203)) and not (layer0_outputs(5099));
    layer1_outputs(1821) <= not((layer0_outputs(3650)) or (layer0_outputs(887)));
    layer1_outputs(1822) <= not(layer0_outputs(3297));
    layer1_outputs(1823) <= not(layer0_outputs(335));
    layer1_outputs(1824) <= '1';
    layer1_outputs(1825) <= (layer0_outputs(3792)) and not (layer0_outputs(2280));
    layer1_outputs(1826) <= not(layer0_outputs(994));
    layer1_outputs(1827) <= (layer0_outputs(4306)) and (layer0_outputs(4928));
    layer1_outputs(1828) <= (layer0_outputs(3312)) and not (layer0_outputs(4390));
    layer1_outputs(1829) <= '1';
    layer1_outputs(1830) <= (layer0_outputs(4250)) and not (layer0_outputs(377));
    layer1_outputs(1831) <= not((layer0_outputs(2221)) and (layer0_outputs(985)));
    layer1_outputs(1832) <= (layer0_outputs(4712)) and not (layer0_outputs(4588));
    layer1_outputs(1833) <= not((layer0_outputs(3479)) and (layer0_outputs(3957)));
    layer1_outputs(1834) <= (layer0_outputs(1873)) and (layer0_outputs(269));
    layer1_outputs(1835) <= (layer0_outputs(3517)) and not (layer0_outputs(1456));
    layer1_outputs(1836) <= (layer0_outputs(309)) and (layer0_outputs(2233));
    layer1_outputs(1837) <= (layer0_outputs(4900)) and (layer0_outputs(1561));
    layer1_outputs(1838) <= (layer0_outputs(1769)) and (layer0_outputs(2600));
    layer1_outputs(1839) <= not((layer0_outputs(944)) or (layer0_outputs(1608)));
    layer1_outputs(1840) <= not(layer0_outputs(1380)) or (layer0_outputs(3738));
    layer1_outputs(1841) <= (layer0_outputs(4559)) and not (layer0_outputs(186));
    layer1_outputs(1842) <= '1';
    layer1_outputs(1843) <= not((layer0_outputs(3642)) and (layer0_outputs(4823)));
    layer1_outputs(1844) <= not(layer0_outputs(557)) or (layer0_outputs(3054));
    layer1_outputs(1845) <= not(layer0_outputs(3500));
    layer1_outputs(1846) <= (layer0_outputs(654)) or (layer0_outputs(2563));
    layer1_outputs(1847) <= not((layer0_outputs(456)) and (layer0_outputs(1682)));
    layer1_outputs(1848) <= (layer0_outputs(2501)) or (layer0_outputs(583));
    layer1_outputs(1849) <= layer0_outputs(2365);
    layer1_outputs(1850) <= not(layer0_outputs(3246)) or (layer0_outputs(3615));
    layer1_outputs(1851) <= '0';
    layer1_outputs(1852) <= not(layer0_outputs(2759)) or (layer0_outputs(323));
    layer1_outputs(1853) <= (layer0_outputs(3673)) and not (layer0_outputs(4027));
    layer1_outputs(1854) <= not((layer0_outputs(1870)) or (layer0_outputs(2949)));
    layer1_outputs(1855) <= layer0_outputs(1736);
    layer1_outputs(1856) <= layer0_outputs(1704);
    layer1_outputs(1857) <= (layer0_outputs(3685)) or (layer0_outputs(221));
    layer1_outputs(1858) <= not((layer0_outputs(3620)) and (layer0_outputs(2711)));
    layer1_outputs(1859) <= '1';
    layer1_outputs(1860) <= (layer0_outputs(1179)) and not (layer0_outputs(237));
    layer1_outputs(1861) <= layer0_outputs(4218);
    layer1_outputs(1862) <= '0';
    layer1_outputs(1863) <= (layer0_outputs(3732)) or (layer0_outputs(4732));
    layer1_outputs(1864) <= layer0_outputs(2198);
    layer1_outputs(1865) <= (layer0_outputs(4993)) and not (layer0_outputs(780));
    layer1_outputs(1866) <= '0';
    layer1_outputs(1867) <= layer0_outputs(4577);
    layer1_outputs(1868) <= (layer0_outputs(4419)) and not (layer0_outputs(609));
    layer1_outputs(1869) <= (layer0_outputs(2462)) and not (layer0_outputs(4259));
    layer1_outputs(1870) <= (layer0_outputs(3553)) and not (layer0_outputs(1431));
    layer1_outputs(1871) <= not((layer0_outputs(768)) or (layer0_outputs(2547)));
    layer1_outputs(1872) <= not(layer0_outputs(2463));
    layer1_outputs(1873) <= (layer0_outputs(4143)) and (layer0_outputs(3837));
    layer1_outputs(1874) <= '1';
    layer1_outputs(1875) <= layer0_outputs(2160);
    layer1_outputs(1876) <= (layer0_outputs(2984)) or (layer0_outputs(466));
    layer1_outputs(1877) <= '0';
    layer1_outputs(1878) <= not(layer0_outputs(3423));
    layer1_outputs(1879) <= '1';
    layer1_outputs(1880) <= '0';
    layer1_outputs(1881) <= '0';
    layer1_outputs(1882) <= not(layer0_outputs(4494));
    layer1_outputs(1883) <= '0';
    layer1_outputs(1884) <= not(layer0_outputs(1834));
    layer1_outputs(1885) <= not(layer0_outputs(419));
    layer1_outputs(1886) <= not((layer0_outputs(4897)) or (layer0_outputs(2222)));
    layer1_outputs(1887) <= (layer0_outputs(1440)) or (layer0_outputs(2828));
    layer1_outputs(1888) <= layer0_outputs(551);
    layer1_outputs(1889) <= (layer0_outputs(4772)) xor (layer0_outputs(2399));
    layer1_outputs(1890) <= not(layer0_outputs(1316)) or (layer0_outputs(2886));
    layer1_outputs(1891) <= '0';
    layer1_outputs(1892) <= not(layer0_outputs(991)) or (layer0_outputs(4544));
    layer1_outputs(1893) <= not(layer0_outputs(5037));
    layer1_outputs(1894) <= not(layer0_outputs(55)) or (layer0_outputs(4153));
    layer1_outputs(1895) <= layer0_outputs(1424);
    layer1_outputs(1896) <= layer0_outputs(1909);
    layer1_outputs(1897) <= '0';
    layer1_outputs(1898) <= not((layer0_outputs(683)) or (layer0_outputs(1842)));
    layer1_outputs(1899) <= not((layer0_outputs(23)) or (layer0_outputs(1815)));
    layer1_outputs(1900) <= (layer0_outputs(2504)) and (layer0_outputs(3945));
    layer1_outputs(1901) <= (layer0_outputs(819)) and not (layer0_outputs(2529));
    layer1_outputs(1902) <= '0';
    layer1_outputs(1903) <= not(layer0_outputs(266));
    layer1_outputs(1904) <= (layer0_outputs(3930)) xor (layer0_outputs(2104));
    layer1_outputs(1905) <= not(layer0_outputs(176));
    layer1_outputs(1906) <= '0';
    layer1_outputs(1907) <= not(layer0_outputs(4219));
    layer1_outputs(1908) <= '1';
    layer1_outputs(1909) <= not((layer0_outputs(3904)) and (layer0_outputs(2779)));
    layer1_outputs(1910) <= (layer0_outputs(2889)) and not (layer0_outputs(4506));
    layer1_outputs(1911) <= not((layer0_outputs(3342)) or (layer0_outputs(2371)));
    layer1_outputs(1912) <= not(layer0_outputs(4548));
    layer1_outputs(1913) <= not(layer0_outputs(831)) or (layer0_outputs(1312));
    layer1_outputs(1914) <= (layer0_outputs(273)) or (layer0_outputs(2558));
    layer1_outputs(1915) <= '1';
    layer1_outputs(1916) <= (layer0_outputs(1553)) and not (layer0_outputs(3024));
    layer1_outputs(1917) <= not(layer0_outputs(2860));
    layer1_outputs(1918) <= '0';
    layer1_outputs(1919) <= layer0_outputs(991);
    layer1_outputs(1920) <= not(layer0_outputs(172));
    layer1_outputs(1921) <= '0';
    layer1_outputs(1922) <= layer0_outputs(98);
    layer1_outputs(1923) <= '0';
    layer1_outputs(1924) <= not(layer0_outputs(4696));
    layer1_outputs(1925) <= not(layer0_outputs(714));
    layer1_outputs(1926) <= (layer0_outputs(4616)) or (layer0_outputs(2601));
    layer1_outputs(1927) <= '0';
    layer1_outputs(1928) <= (layer0_outputs(4216)) and (layer0_outputs(4030));
    layer1_outputs(1929) <= not(layer0_outputs(4070));
    layer1_outputs(1930) <= not(layer0_outputs(2964)) or (layer0_outputs(3664));
    layer1_outputs(1931) <= '1';
    layer1_outputs(1932) <= (layer0_outputs(4949)) and not (layer0_outputs(1572));
    layer1_outputs(1933) <= layer0_outputs(616);
    layer1_outputs(1934) <= '0';
    layer1_outputs(1935) <= layer0_outputs(3193);
    layer1_outputs(1936) <= (layer0_outputs(3785)) and not (layer0_outputs(2996));
    layer1_outputs(1937) <= not((layer0_outputs(5098)) and (layer0_outputs(440)));
    layer1_outputs(1938) <= (layer0_outputs(4006)) or (layer0_outputs(681));
    layer1_outputs(1939) <= not(layer0_outputs(3571)) or (layer0_outputs(2692));
    layer1_outputs(1940) <= '1';
    layer1_outputs(1941) <= layer0_outputs(1005);
    layer1_outputs(1942) <= (layer0_outputs(2191)) and not (layer0_outputs(2303));
    layer1_outputs(1943) <= layer0_outputs(315);
    layer1_outputs(1944) <= not((layer0_outputs(4173)) and (layer0_outputs(3081)));
    layer1_outputs(1945) <= '1';
    layer1_outputs(1946) <= (layer0_outputs(2344)) and (layer0_outputs(4908));
    layer1_outputs(1947) <= not(layer0_outputs(1982)) or (layer0_outputs(4192));
    layer1_outputs(1948) <= not((layer0_outputs(1688)) or (layer0_outputs(5019)));
    layer1_outputs(1949) <= layer0_outputs(2698);
    layer1_outputs(1950) <= not(layer0_outputs(5096)) or (layer0_outputs(1419));
    layer1_outputs(1951) <= (layer0_outputs(4181)) and (layer0_outputs(2882));
    layer1_outputs(1952) <= '0';
    layer1_outputs(1953) <= not(layer0_outputs(226)) or (layer0_outputs(3932));
    layer1_outputs(1954) <= (layer0_outputs(2123)) and not (layer0_outputs(3895));
    layer1_outputs(1955) <= not(layer0_outputs(1681));
    layer1_outputs(1956) <= not(layer0_outputs(5036));
    layer1_outputs(1957) <= layer0_outputs(2897);
    layer1_outputs(1958) <= not(layer0_outputs(5076));
    layer1_outputs(1959) <= not((layer0_outputs(2523)) and (layer0_outputs(914)));
    layer1_outputs(1960) <= (layer0_outputs(334)) and not (layer0_outputs(4115));
    layer1_outputs(1961) <= not(layer0_outputs(767)) or (layer0_outputs(4184));
    layer1_outputs(1962) <= not(layer0_outputs(3520));
    layer1_outputs(1963) <= not(layer0_outputs(1311));
    layer1_outputs(1964) <= not(layer0_outputs(2249)) or (layer0_outputs(602));
    layer1_outputs(1965) <= (layer0_outputs(1047)) xor (layer0_outputs(5012));
    layer1_outputs(1966) <= not(layer0_outputs(1931));
    layer1_outputs(1967) <= (layer0_outputs(845)) and not (layer0_outputs(4909));
    layer1_outputs(1968) <= (layer0_outputs(2163)) or (layer0_outputs(4955));
    layer1_outputs(1969) <= '0';
    layer1_outputs(1970) <= '1';
    layer1_outputs(1971) <= layer0_outputs(2092);
    layer1_outputs(1972) <= '0';
    layer1_outputs(1973) <= not(layer0_outputs(1035));
    layer1_outputs(1974) <= not(layer0_outputs(4613)) or (layer0_outputs(2085));
    layer1_outputs(1975) <= '1';
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= layer0_outputs(125);
    layer1_outputs(1978) <= (layer0_outputs(2894)) and not (layer0_outputs(369));
    layer1_outputs(1979) <= '1';
    layer1_outputs(1980) <= '1';
    layer1_outputs(1981) <= (layer0_outputs(3907)) and (layer0_outputs(999));
    layer1_outputs(1982) <= (layer0_outputs(3644)) xor (layer0_outputs(99));
    layer1_outputs(1983) <= not((layer0_outputs(2048)) or (layer0_outputs(4908)));
    layer1_outputs(1984) <= not(layer0_outputs(2856));
    layer1_outputs(1985) <= not(layer0_outputs(2737));
    layer1_outputs(1986) <= not(layer0_outputs(621)) or (layer0_outputs(2345));
    layer1_outputs(1987) <= not((layer0_outputs(2967)) and (layer0_outputs(4266)));
    layer1_outputs(1988) <= '1';
    layer1_outputs(1989) <= not(layer0_outputs(4091));
    layer1_outputs(1990) <= layer0_outputs(4859);
    layer1_outputs(1991) <= (layer0_outputs(2054)) and not (layer0_outputs(5073));
    layer1_outputs(1992) <= not((layer0_outputs(631)) or (layer0_outputs(3014)));
    layer1_outputs(1993) <= (layer0_outputs(3117)) and not (layer0_outputs(682));
    layer1_outputs(1994) <= not(layer0_outputs(4290));
    layer1_outputs(1995) <= not((layer0_outputs(2878)) and (layer0_outputs(4105)));
    layer1_outputs(1996) <= (layer0_outputs(2251)) and not (layer0_outputs(1764));
    layer1_outputs(1997) <= layer0_outputs(432);
    layer1_outputs(1998) <= not(layer0_outputs(4443));
    layer1_outputs(1999) <= layer0_outputs(509);
    layer1_outputs(2000) <= (layer0_outputs(413)) and not (layer0_outputs(2712));
    layer1_outputs(2001) <= '0';
    layer1_outputs(2002) <= not(layer0_outputs(1150));
    layer1_outputs(2003) <= (layer0_outputs(4337)) and (layer0_outputs(70));
    layer1_outputs(2004) <= (layer0_outputs(1133)) and not (layer0_outputs(1610));
    layer1_outputs(2005) <= not((layer0_outputs(3401)) or (layer0_outputs(4437)));
    layer1_outputs(2006) <= layer0_outputs(2779);
    layer1_outputs(2007) <= layer0_outputs(3518);
    layer1_outputs(2008) <= (layer0_outputs(1752)) and not (layer0_outputs(4871));
    layer1_outputs(2009) <= (layer0_outputs(3701)) or (layer0_outputs(1129));
    layer1_outputs(2010) <= '1';
    layer1_outputs(2011) <= not(layer0_outputs(3054)) or (layer0_outputs(478));
    layer1_outputs(2012) <= '1';
    layer1_outputs(2013) <= (layer0_outputs(3156)) and not (layer0_outputs(1531));
    layer1_outputs(2014) <= (layer0_outputs(6)) or (layer0_outputs(705));
    layer1_outputs(2015) <= (layer0_outputs(290)) and (layer0_outputs(1063));
    layer1_outputs(2016) <= (layer0_outputs(851)) and not (layer0_outputs(3756));
    layer1_outputs(2017) <= (layer0_outputs(1331)) and not (layer0_outputs(4929));
    layer1_outputs(2018) <= layer0_outputs(4322);
    layer1_outputs(2019) <= (layer0_outputs(2788)) and not (layer0_outputs(1565));
    layer1_outputs(2020) <= (layer0_outputs(1069)) and not (layer0_outputs(1487));
    layer1_outputs(2021) <= layer0_outputs(3838);
    layer1_outputs(2022) <= not(layer0_outputs(2837)) or (layer0_outputs(1715));
    layer1_outputs(2023) <= (layer0_outputs(1546)) or (layer0_outputs(4673));
    layer1_outputs(2024) <= layer0_outputs(3949);
    layer1_outputs(2025) <= not(layer0_outputs(4213)) or (layer0_outputs(397));
    layer1_outputs(2026) <= not(layer0_outputs(111)) or (layer0_outputs(3929));
    layer1_outputs(2027) <= (layer0_outputs(1704)) and not (layer0_outputs(4296));
    layer1_outputs(2028) <= not(layer0_outputs(3856));
    layer1_outputs(2029) <= not(layer0_outputs(2700)) or (layer0_outputs(3212));
    layer1_outputs(2030) <= (layer0_outputs(2089)) or (layer0_outputs(723));
    layer1_outputs(2031) <= layer0_outputs(1554);
    layer1_outputs(2032) <= not((layer0_outputs(3685)) or (layer0_outputs(1584)));
    layer1_outputs(2033) <= '1';
    layer1_outputs(2034) <= '1';
    layer1_outputs(2035) <= '0';
    layer1_outputs(2036) <= (layer0_outputs(1264)) and not (layer0_outputs(1945));
    layer1_outputs(2037) <= '0';
    layer1_outputs(2038) <= not(layer0_outputs(4254));
    layer1_outputs(2039) <= not(layer0_outputs(3007)) or (layer0_outputs(4182));
    layer1_outputs(2040) <= not((layer0_outputs(721)) and (layer0_outputs(3171)));
    layer1_outputs(2041) <= not((layer0_outputs(4224)) or (layer0_outputs(2829)));
    layer1_outputs(2042) <= not(layer0_outputs(1269)) or (layer0_outputs(1464));
    layer1_outputs(2043) <= not(layer0_outputs(2347));
    layer1_outputs(2044) <= (layer0_outputs(3554)) and (layer0_outputs(2105));
    layer1_outputs(2045) <= layer0_outputs(3598);
    layer1_outputs(2046) <= not(layer0_outputs(943));
    layer1_outputs(2047) <= (layer0_outputs(2082)) and not (layer0_outputs(2726));
    layer1_outputs(2048) <= '1';
    layer1_outputs(2049) <= '0';
    layer1_outputs(2050) <= not(layer0_outputs(4060));
    layer1_outputs(2051) <= layer0_outputs(4436);
    layer1_outputs(2052) <= layer0_outputs(5099);
    layer1_outputs(2053) <= not(layer0_outputs(3623));
    layer1_outputs(2054) <= (layer0_outputs(697)) and not (layer0_outputs(3303));
    layer1_outputs(2055) <= not(layer0_outputs(3105)) or (layer0_outputs(3290));
    layer1_outputs(2056) <= (layer0_outputs(5082)) and not (layer0_outputs(264));
    layer1_outputs(2057) <= not(layer0_outputs(4412));
    layer1_outputs(2058) <= (layer0_outputs(3798)) xor (layer0_outputs(1617));
    layer1_outputs(2059) <= not(layer0_outputs(2107));
    layer1_outputs(2060) <= not((layer0_outputs(4522)) and (layer0_outputs(4265)));
    layer1_outputs(2061) <= not(layer0_outputs(4268));
    layer1_outputs(2062) <= not(layer0_outputs(1575)) or (layer0_outputs(2241));
    layer1_outputs(2063) <= not(layer0_outputs(3349));
    layer1_outputs(2064) <= not((layer0_outputs(1808)) and (layer0_outputs(4009)));
    layer1_outputs(2065) <= '1';
    layer1_outputs(2066) <= (layer0_outputs(3375)) and (layer0_outputs(3069));
    layer1_outputs(2067) <= (layer0_outputs(185)) and not (layer0_outputs(979));
    layer1_outputs(2068) <= not((layer0_outputs(1656)) and (layer0_outputs(4954)));
    layer1_outputs(2069) <= not(layer0_outputs(393));
    layer1_outputs(2070) <= (layer0_outputs(3548)) or (layer0_outputs(1406));
    layer1_outputs(2071) <= not((layer0_outputs(3473)) and (layer0_outputs(1422)));
    layer1_outputs(2072) <= '1';
    layer1_outputs(2073) <= not((layer0_outputs(1619)) or (layer0_outputs(3717)));
    layer1_outputs(2074) <= (layer0_outputs(1550)) or (layer0_outputs(2004));
    layer1_outputs(2075) <= not(layer0_outputs(3378));
    layer1_outputs(2076) <= not(layer0_outputs(4241));
    layer1_outputs(2077) <= (layer0_outputs(3757)) and not (layer0_outputs(3164));
    layer1_outputs(2078) <= (layer0_outputs(1735)) or (layer0_outputs(2989));
    layer1_outputs(2079) <= '0';
    layer1_outputs(2080) <= layer0_outputs(2879);
    layer1_outputs(2081) <= '1';
    layer1_outputs(2082) <= not((layer0_outputs(2736)) and (layer0_outputs(2840)));
    layer1_outputs(2083) <= not(layer0_outputs(4279)) or (layer0_outputs(1383));
    layer1_outputs(2084) <= (layer0_outputs(3834)) and not (layer0_outputs(3873));
    layer1_outputs(2085) <= layer0_outputs(1954);
    layer1_outputs(2086) <= not(layer0_outputs(690));
    layer1_outputs(2087) <= '0';
    layer1_outputs(2088) <= layer0_outputs(4580);
    layer1_outputs(2089) <= not(layer0_outputs(4741)) or (layer0_outputs(425));
    layer1_outputs(2090) <= (layer0_outputs(1831)) and not (layer0_outputs(2067));
    layer1_outputs(2091) <= (layer0_outputs(1181)) and not (layer0_outputs(4764));
    layer1_outputs(2092) <= '1';
    layer1_outputs(2093) <= not(layer0_outputs(3156));
    layer1_outputs(2094) <= (layer0_outputs(781)) and not (layer0_outputs(2503));
    layer1_outputs(2095) <= layer0_outputs(3803);
    layer1_outputs(2096) <= '0';
    layer1_outputs(2097) <= not(layer0_outputs(3160));
    layer1_outputs(2098) <= '0';
    layer1_outputs(2099) <= not(layer0_outputs(2129));
    layer1_outputs(2100) <= not((layer0_outputs(1718)) and (layer0_outputs(1822)));
    layer1_outputs(2101) <= '1';
    layer1_outputs(2102) <= (layer0_outputs(2702)) or (layer0_outputs(71));
    layer1_outputs(2103) <= not((layer0_outputs(2144)) and (layer0_outputs(2170)));
    layer1_outputs(2104) <= layer0_outputs(4582);
    layer1_outputs(2105) <= '1';
    layer1_outputs(2106) <= not(layer0_outputs(4475));
    layer1_outputs(2107) <= not(layer0_outputs(1672)) or (layer0_outputs(645));
    layer1_outputs(2108) <= '1';
    layer1_outputs(2109) <= not(layer0_outputs(650)) or (layer0_outputs(2820));
    layer1_outputs(2110) <= not(layer0_outputs(3492)) or (layer0_outputs(1746));
    layer1_outputs(2111) <= (layer0_outputs(5113)) or (layer0_outputs(3481));
    layer1_outputs(2112) <= not((layer0_outputs(2641)) or (layer0_outputs(1470)));
    layer1_outputs(2113) <= '1';
    layer1_outputs(2114) <= not(layer0_outputs(4329)) or (layer0_outputs(1476));
    layer1_outputs(2115) <= not((layer0_outputs(3198)) and (layer0_outputs(4577)));
    layer1_outputs(2116) <= not(layer0_outputs(4274)) or (layer0_outputs(1416));
    layer1_outputs(2117) <= not(layer0_outputs(2524));
    layer1_outputs(2118) <= '1';
    layer1_outputs(2119) <= not((layer0_outputs(2334)) or (layer0_outputs(4656)));
    layer1_outputs(2120) <= not(layer0_outputs(4648));
    layer1_outputs(2121) <= not(layer0_outputs(3845)) or (layer0_outputs(833));
    layer1_outputs(2122) <= not(layer0_outputs(2943));
    layer1_outputs(2123) <= layer0_outputs(3354);
    layer1_outputs(2124) <= layer0_outputs(4887);
    layer1_outputs(2125) <= not(layer0_outputs(744)) or (layer0_outputs(376));
    layer1_outputs(2126) <= '1';
    layer1_outputs(2127) <= not(layer0_outputs(3273)) or (layer0_outputs(347));
    layer1_outputs(2128) <= not(layer0_outputs(4989)) or (layer0_outputs(5084));
    layer1_outputs(2129) <= not(layer0_outputs(4217));
    layer1_outputs(2130) <= (layer0_outputs(4499)) and not (layer0_outputs(3663));
    layer1_outputs(2131) <= (layer0_outputs(4126)) and not (layer0_outputs(569));
    layer1_outputs(2132) <= layer0_outputs(4113);
    layer1_outputs(2133) <= (layer0_outputs(4980)) and not (layer0_outputs(24));
    layer1_outputs(2134) <= layer0_outputs(2414);
    layer1_outputs(2135) <= (layer0_outputs(469)) and not (layer0_outputs(3887));
    layer1_outputs(2136) <= not(layer0_outputs(4751));
    layer1_outputs(2137) <= not(layer0_outputs(901));
    layer1_outputs(2138) <= not(layer0_outputs(3126));
    layer1_outputs(2139) <= not((layer0_outputs(3568)) and (layer0_outputs(3606)));
    layer1_outputs(2140) <= (layer0_outputs(1057)) and (layer0_outputs(3883));
    layer1_outputs(2141) <= not((layer0_outputs(826)) xor (layer0_outputs(2156)));
    layer1_outputs(2142) <= '0';
    layer1_outputs(2143) <= not(layer0_outputs(1501));
    layer1_outputs(2144) <= not((layer0_outputs(331)) or (layer0_outputs(1077)));
    layer1_outputs(2145) <= '1';
    layer1_outputs(2146) <= not(layer0_outputs(4509));
    layer1_outputs(2147) <= (layer0_outputs(5035)) and not (layer0_outputs(888));
    layer1_outputs(2148) <= '1';
    layer1_outputs(2149) <= not((layer0_outputs(4004)) or (layer0_outputs(2931)));
    layer1_outputs(2150) <= '1';
    layer1_outputs(2151) <= (layer0_outputs(2844)) and (layer0_outputs(574));
    layer1_outputs(2152) <= not((layer0_outputs(133)) and (layer0_outputs(810)));
    layer1_outputs(2153) <= not(layer0_outputs(2393)) or (layer0_outputs(2946));
    layer1_outputs(2154) <= not((layer0_outputs(3098)) or (layer0_outputs(2364)));
    layer1_outputs(2155) <= (layer0_outputs(5092)) and not (layer0_outputs(2450));
    layer1_outputs(2156) <= layer0_outputs(5071);
    layer1_outputs(2157) <= not(layer0_outputs(3693)) or (layer0_outputs(4315));
    layer1_outputs(2158) <= '0';
    layer1_outputs(2159) <= not(layer0_outputs(2718));
    layer1_outputs(2160) <= (layer0_outputs(1054)) and not (layer0_outputs(464));
    layer1_outputs(2161) <= '0';
    layer1_outputs(2162) <= '1';
    layer1_outputs(2163) <= (layer0_outputs(2574)) and not (layer0_outputs(2486));
    layer1_outputs(2164) <= (layer0_outputs(2467)) and not (layer0_outputs(4855));
    layer1_outputs(2165) <= not(layer0_outputs(2195));
    layer1_outputs(2166) <= (layer0_outputs(930)) and not (layer0_outputs(4729));
    layer1_outputs(2167) <= not(layer0_outputs(3048));
    layer1_outputs(2168) <= not((layer0_outputs(3624)) and (layer0_outputs(1699)));
    layer1_outputs(2169) <= layer0_outputs(687);
    layer1_outputs(2170) <= '1';
    layer1_outputs(2171) <= not(layer0_outputs(1782));
    layer1_outputs(2172) <= not((layer0_outputs(1263)) xor (layer0_outputs(1176)));
    layer1_outputs(2173) <= (layer0_outputs(55)) and not (layer0_outputs(513));
    layer1_outputs(2174) <= layer0_outputs(2969);
    layer1_outputs(2175) <= '1';
    layer1_outputs(2176) <= not(layer0_outputs(753)) or (layer0_outputs(3845));
    layer1_outputs(2177) <= '1';
    layer1_outputs(2178) <= not(layer0_outputs(632)) or (layer0_outputs(520));
    layer1_outputs(2179) <= (layer0_outputs(4076)) or (layer0_outputs(1340));
    layer1_outputs(2180) <= not((layer0_outputs(4049)) or (layer0_outputs(320)));
    layer1_outputs(2181) <= not((layer0_outputs(5102)) or (layer0_outputs(5024)));
    layer1_outputs(2182) <= not(layer0_outputs(5009));
    layer1_outputs(2183) <= not((layer0_outputs(4740)) or (layer0_outputs(1623)));
    layer1_outputs(2184) <= not((layer0_outputs(1796)) or (layer0_outputs(2385)));
    layer1_outputs(2185) <= '1';
    layer1_outputs(2186) <= (layer0_outputs(2911)) and (layer0_outputs(2561));
    layer1_outputs(2187) <= layer0_outputs(2350);
    layer1_outputs(2188) <= not(layer0_outputs(362));
    layer1_outputs(2189) <= layer0_outputs(1942);
    layer1_outputs(2190) <= (layer0_outputs(4545)) and not (layer0_outputs(2662));
    layer1_outputs(2191) <= not((layer0_outputs(4679)) and (layer0_outputs(3324)));
    layer1_outputs(2192) <= not(layer0_outputs(4109));
    layer1_outputs(2193) <= (layer0_outputs(4138)) or (layer0_outputs(3459));
    layer1_outputs(2194) <= not(layer0_outputs(1065)) or (layer0_outputs(1624));
    layer1_outputs(2195) <= (layer0_outputs(3970)) and not (layer0_outputs(1991));
    layer1_outputs(2196) <= '1';
    layer1_outputs(2197) <= (layer0_outputs(4699)) or (layer0_outputs(3796));
    layer1_outputs(2198) <= (layer0_outputs(2281)) or (layer0_outputs(1573));
    layer1_outputs(2199) <= '1';
    layer1_outputs(2200) <= '0';
    layer1_outputs(2201) <= (layer0_outputs(3994)) or (layer0_outputs(5096));
    layer1_outputs(2202) <= not(layer0_outputs(2038));
    layer1_outputs(2203) <= layer0_outputs(1996);
    layer1_outputs(2204) <= layer0_outputs(1141);
    layer1_outputs(2205) <= '1';
    layer1_outputs(2206) <= layer0_outputs(2918);
    layer1_outputs(2207) <= not(layer0_outputs(2564)) or (layer0_outputs(2357));
    layer1_outputs(2208) <= not(layer0_outputs(801));
    layer1_outputs(2209) <= not(layer0_outputs(4799)) or (layer0_outputs(3986));
    layer1_outputs(2210) <= layer0_outputs(2611);
    layer1_outputs(2211) <= not(layer0_outputs(1175));
    layer1_outputs(2212) <= not(layer0_outputs(2333));
    layer1_outputs(2213) <= (layer0_outputs(926)) and not (layer0_outputs(1460));
    layer1_outputs(2214) <= not((layer0_outputs(1045)) or (layer0_outputs(796)));
    layer1_outputs(2215) <= not((layer0_outputs(604)) or (layer0_outputs(2029)));
    layer1_outputs(2216) <= not(layer0_outputs(3558)) or (layer0_outputs(4059));
    layer1_outputs(2217) <= not((layer0_outputs(3115)) and (layer0_outputs(3497)));
    layer1_outputs(2218) <= '0';
    layer1_outputs(2219) <= (layer0_outputs(1026)) and (layer0_outputs(2173));
    layer1_outputs(2220) <= not((layer0_outputs(349)) and (layer0_outputs(2397)));
    layer1_outputs(2221) <= (layer0_outputs(3870)) and not (layer0_outputs(3890));
    layer1_outputs(2222) <= not(layer0_outputs(3967));
    layer1_outputs(2223) <= not((layer0_outputs(2951)) or (layer0_outputs(4169)));
    layer1_outputs(2224) <= not((layer0_outputs(3326)) and (layer0_outputs(3488)));
    layer1_outputs(2225) <= '0';
    layer1_outputs(2226) <= not(layer0_outputs(843));
    layer1_outputs(2227) <= not(layer0_outputs(653));
    layer1_outputs(2228) <= '0';
    layer1_outputs(2229) <= (layer0_outputs(1536)) and not (layer0_outputs(2345));
    layer1_outputs(2230) <= not(layer0_outputs(3273)) or (layer0_outputs(4697));
    layer1_outputs(2231) <= not((layer0_outputs(345)) or (layer0_outputs(1337)));
    layer1_outputs(2232) <= layer0_outputs(4827);
    layer1_outputs(2233) <= layer0_outputs(4208);
    layer1_outputs(2234) <= (layer0_outputs(1335)) and not (layer0_outputs(868));
    layer1_outputs(2235) <= not(layer0_outputs(378)) or (layer0_outputs(4468));
    layer1_outputs(2236) <= not(layer0_outputs(727)) or (layer0_outputs(2372));
    layer1_outputs(2237) <= not(layer0_outputs(3317)) or (layer0_outputs(1421));
    layer1_outputs(2238) <= (layer0_outputs(3196)) and not (layer0_outputs(2655));
    layer1_outputs(2239) <= (layer0_outputs(2087)) and not (layer0_outputs(4364));
    layer1_outputs(2240) <= not(layer0_outputs(1430));
    layer1_outputs(2241) <= not(layer0_outputs(1977)) or (layer0_outputs(2883));
    layer1_outputs(2242) <= not(layer0_outputs(3634));
    layer1_outputs(2243) <= '1';
    layer1_outputs(2244) <= (layer0_outputs(1721)) or (layer0_outputs(3380));
    layer1_outputs(2245) <= layer0_outputs(2538);
    layer1_outputs(2246) <= layer0_outputs(3335);
    layer1_outputs(2247) <= not(layer0_outputs(838)) or (layer0_outputs(3389));
    layer1_outputs(2248) <= not(layer0_outputs(3227)) or (layer0_outputs(3720));
    layer1_outputs(2249) <= '1';
    layer1_outputs(2250) <= (layer0_outputs(905)) or (layer0_outputs(4560));
    layer1_outputs(2251) <= not(layer0_outputs(1794)) or (layer0_outputs(3669));
    layer1_outputs(2252) <= not((layer0_outputs(858)) and (layer0_outputs(4854)));
    layer1_outputs(2253) <= not((layer0_outputs(2771)) and (layer0_outputs(2115)));
    layer1_outputs(2254) <= '0';
    layer1_outputs(2255) <= (layer0_outputs(2621)) and not (layer0_outputs(2631));
    layer1_outputs(2256) <= not(layer0_outputs(4823));
    layer1_outputs(2257) <= '0';
    layer1_outputs(2258) <= not((layer0_outputs(1043)) and (layer0_outputs(902)));
    layer1_outputs(2259) <= not(layer0_outputs(3787));
    layer1_outputs(2260) <= not((layer0_outputs(4091)) and (layer0_outputs(3272)));
    layer1_outputs(2261) <= layer0_outputs(2880);
    layer1_outputs(2262) <= (layer0_outputs(804)) or (layer0_outputs(3710));
    layer1_outputs(2263) <= '1';
    layer1_outputs(2264) <= layer0_outputs(3288);
    layer1_outputs(2265) <= not(layer0_outputs(299)) or (layer0_outputs(4431));
    layer1_outputs(2266) <= (layer0_outputs(3895)) and (layer0_outputs(4372));
    layer1_outputs(2267) <= '0';
    layer1_outputs(2268) <= not((layer0_outputs(840)) or (layer0_outputs(3498)));
    layer1_outputs(2269) <= not((layer0_outputs(2302)) and (layer0_outputs(3957)));
    layer1_outputs(2270) <= not(layer0_outputs(1371));
    layer1_outputs(2271) <= (layer0_outputs(1622)) xor (layer0_outputs(4905));
    layer1_outputs(2272) <= not((layer0_outputs(1468)) or (layer0_outputs(1158)));
    layer1_outputs(2273) <= not(layer0_outputs(1370));
    layer1_outputs(2274) <= '1';
    layer1_outputs(2275) <= not(layer0_outputs(1849)) or (layer0_outputs(2095));
    layer1_outputs(2276) <= '0';
    layer1_outputs(2277) <= layer0_outputs(4715);
    layer1_outputs(2278) <= layer0_outputs(1009);
    layer1_outputs(2279) <= (layer0_outputs(4345)) or (layer0_outputs(769));
    layer1_outputs(2280) <= (layer0_outputs(2431)) or (layer0_outputs(3542));
    layer1_outputs(2281) <= layer0_outputs(4202);
    layer1_outputs(2282) <= '1';
    layer1_outputs(2283) <= not(layer0_outputs(2733));
    layer1_outputs(2284) <= not(layer0_outputs(2376));
    layer1_outputs(2285) <= (layer0_outputs(1443)) and not (layer0_outputs(3643));
    layer1_outputs(2286) <= not(layer0_outputs(4555)) or (layer0_outputs(3892));
    layer1_outputs(2287) <= '1';
    layer1_outputs(2288) <= '1';
    layer1_outputs(2289) <= not(layer0_outputs(2152));
    layer1_outputs(2290) <= not(layer0_outputs(977));
    layer1_outputs(2291) <= (layer0_outputs(3781)) and not (layer0_outputs(1533));
    layer1_outputs(2292) <= not(layer0_outputs(4933));
    layer1_outputs(2293) <= not(layer0_outputs(138));
    layer1_outputs(2294) <= not((layer0_outputs(3811)) xor (layer0_outputs(4379)));
    layer1_outputs(2295) <= not(layer0_outputs(1467));
    layer1_outputs(2296) <= not(layer0_outputs(2214)) or (layer0_outputs(5040));
    layer1_outputs(2297) <= (layer0_outputs(1613)) xor (layer0_outputs(1239));
    layer1_outputs(2298) <= not((layer0_outputs(4848)) and (layer0_outputs(2465)));
    layer1_outputs(2299) <= (layer0_outputs(3077)) and not (layer0_outputs(3741));
    layer1_outputs(2300) <= (layer0_outputs(3118)) and not (layer0_outputs(3789));
    layer1_outputs(2301) <= layer0_outputs(3148);
    layer1_outputs(2302) <= (layer0_outputs(3409)) xor (layer0_outputs(4608));
    layer1_outputs(2303) <= layer0_outputs(2163);
    layer1_outputs(2304) <= not(layer0_outputs(2454));
    layer1_outputs(2305) <= (layer0_outputs(3580)) and (layer0_outputs(910));
    layer1_outputs(2306) <= not(layer0_outputs(354));
    layer1_outputs(2307) <= '1';
    layer1_outputs(2308) <= not(layer0_outputs(2642));
    layer1_outputs(2309) <= (layer0_outputs(882)) and not (layer0_outputs(5085));
    layer1_outputs(2310) <= (layer0_outputs(307)) and not (layer0_outputs(4463));
    layer1_outputs(2311) <= (layer0_outputs(842)) and not (layer0_outputs(1742));
    layer1_outputs(2312) <= not((layer0_outputs(59)) and (layer0_outputs(658)));
    layer1_outputs(2313) <= (layer0_outputs(4747)) and (layer0_outputs(2070));
    layer1_outputs(2314) <= not(layer0_outputs(3306)) or (layer0_outputs(634));
    layer1_outputs(2315) <= (layer0_outputs(3217)) and not (layer0_outputs(3486));
    layer1_outputs(2316) <= not(layer0_outputs(2316));
    layer1_outputs(2317) <= (layer0_outputs(3413)) and not (layer0_outputs(704));
    layer1_outputs(2318) <= layer0_outputs(5079);
    layer1_outputs(2319) <= not(layer0_outputs(512)) or (layer0_outputs(2250));
    layer1_outputs(2320) <= (layer0_outputs(861)) and not (layer0_outputs(4011));
    layer1_outputs(2321) <= (layer0_outputs(2829)) and not (layer0_outputs(938));
    layer1_outputs(2322) <= not(layer0_outputs(1045));
    layer1_outputs(2323) <= '1';
    layer1_outputs(2324) <= layer0_outputs(1848);
    layer1_outputs(2325) <= not((layer0_outputs(4188)) and (layer0_outputs(494)));
    layer1_outputs(2326) <= not(layer0_outputs(728)) or (layer0_outputs(2297));
    layer1_outputs(2327) <= '0';
    layer1_outputs(2328) <= (layer0_outputs(1266)) and not (layer0_outputs(1686));
    layer1_outputs(2329) <= (layer0_outputs(754)) and not (layer0_outputs(1453));
    layer1_outputs(2330) <= (layer0_outputs(3797)) or (layer0_outputs(1291));
    layer1_outputs(2331) <= not((layer0_outputs(4904)) or (layer0_outputs(5044)));
    layer1_outputs(2332) <= not(layer0_outputs(365));
    layer1_outputs(2333) <= not(layer0_outputs(874)) or (layer0_outputs(4634));
    layer1_outputs(2334) <= not((layer0_outputs(919)) or (layer0_outputs(2309)));
    layer1_outputs(2335) <= layer0_outputs(1775);
    layer1_outputs(2336) <= layer0_outputs(3301);
    layer1_outputs(2337) <= layer0_outputs(4612);
    layer1_outputs(2338) <= layer0_outputs(1006);
    layer1_outputs(2339) <= not((layer0_outputs(3751)) and (layer0_outputs(3362)));
    layer1_outputs(2340) <= (layer0_outputs(3295)) or (layer0_outputs(385));
    layer1_outputs(2341) <= layer0_outputs(4288);
    layer1_outputs(2342) <= not(layer0_outputs(3296)) or (layer0_outputs(516));
    layer1_outputs(2343) <= not(layer0_outputs(3077));
    layer1_outputs(2344) <= not(layer0_outputs(4787));
    layer1_outputs(2345) <= (layer0_outputs(267)) and not (layer0_outputs(1878));
    layer1_outputs(2346) <= not(layer0_outputs(399));
    layer1_outputs(2347) <= not(layer0_outputs(3260));
    layer1_outputs(2348) <= not(layer0_outputs(4995)) or (layer0_outputs(2245));
    layer1_outputs(2349) <= '1';
    layer1_outputs(2350) <= (layer0_outputs(3834)) and not (layer0_outputs(4802));
    layer1_outputs(2351) <= not((layer0_outputs(3322)) and (layer0_outputs(539)));
    layer1_outputs(2352) <= not(layer0_outputs(1935));
    layer1_outputs(2353) <= not(layer0_outputs(3428));
    layer1_outputs(2354) <= (layer0_outputs(2623)) xor (layer0_outputs(3549));
    layer1_outputs(2355) <= layer0_outputs(2793);
    layer1_outputs(2356) <= '1';
    layer1_outputs(2357) <= not(layer0_outputs(1224));
    layer1_outputs(2358) <= layer0_outputs(1866);
    layer1_outputs(2359) <= (layer0_outputs(3432)) and not (layer0_outputs(3174));
    layer1_outputs(2360) <= not((layer0_outputs(746)) or (layer0_outputs(1513)));
    layer1_outputs(2361) <= not(layer0_outputs(2540));
    layer1_outputs(2362) <= (layer0_outputs(2288)) and not (layer0_outputs(1069));
    layer1_outputs(2363) <= not((layer0_outputs(3522)) or (layer0_outputs(1702)));
    layer1_outputs(2364) <= layer0_outputs(306);
    layer1_outputs(2365) <= '0';
    layer1_outputs(2366) <= not(layer0_outputs(1234));
    layer1_outputs(2367) <= not((layer0_outputs(2798)) and (layer0_outputs(1000)));
    layer1_outputs(2368) <= layer0_outputs(2134);
    layer1_outputs(2369) <= (layer0_outputs(1771)) and not (layer0_outputs(4368));
    layer1_outputs(2370) <= (layer0_outputs(4866)) or (layer0_outputs(647));
    layer1_outputs(2371) <= not((layer0_outputs(355)) and (layer0_outputs(4730)));
    layer1_outputs(2372) <= (layer0_outputs(1198)) and (layer0_outputs(4914));
    layer1_outputs(2373) <= '1';
    layer1_outputs(2374) <= not((layer0_outputs(5117)) and (layer0_outputs(3651)));
    layer1_outputs(2375) <= (layer0_outputs(2299)) and not (layer0_outputs(3323));
    layer1_outputs(2376) <= not(layer0_outputs(4068));
    layer1_outputs(2377) <= (layer0_outputs(601)) or (layer0_outputs(657));
    layer1_outputs(2378) <= not(layer0_outputs(1572)) or (layer0_outputs(1764));
    layer1_outputs(2379) <= (layer0_outputs(4751)) or (layer0_outputs(452));
    layer1_outputs(2380) <= (layer0_outputs(1970)) and not (layer0_outputs(1001));
    layer1_outputs(2381) <= (layer0_outputs(4081)) and (layer0_outputs(4361));
    layer1_outputs(2382) <= layer0_outputs(2097);
    layer1_outputs(2383) <= layer0_outputs(731);
    layer1_outputs(2384) <= (layer0_outputs(3269)) and not (layer0_outputs(4942));
    layer1_outputs(2385) <= '1';
    layer1_outputs(2386) <= not((layer0_outputs(1059)) and (layer0_outputs(26)));
    layer1_outputs(2387) <= not((layer0_outputs(4582)) or (layer0_outputs(4568)));
    layer1_outputs(2388) <= not((layer0_outputs(4858)) and (layer0_outputs(2227)));
    layer1_outputs(2389) <= (layer0_outputs(4062)) and not (layer0_outputs(2846));
    layer1_outputs(2390) <= not(layer0_outputs(5022));
    layer1_outputs(2391) <= not(layer0_outputs(533)) or (layer0_outputs(2335));
    layer1_outputs(2392) <= not(layer0_outputs(1585)) or (layer0_outputs(818));
    layer1_outputs(2393) <= not((layer0_outputs(3513)) and (layer0_outputs(4186)));
    layer1_outputs(2394) <= not(layer0_outputs(4519)) or (layer0_outputs(1114));
    layer1_outputs(2395) <= (layer0_outputs(2559)) and not (layer0_outputs(1490));
    layer1_outputs(2396) <= not((layer0_outputs(3058)) xor (layer0_outputs(109)));
    layer1_outputs(2397) <= not(layer0_outputs(3978));
    layer1_outputs(2398) <= not(layer0_outputs(2628));
    layer1_outputs(2399) <= layer0_outputs(3208);
    layer1_outputs(2400) <= not(layer0_outputs(4973));
    layer1_outputs(2401) <= not(layer0_outputs(4385));
    layer1_outputs(2402) <= not((layer0_outputs(4906)) and (layer0_outputs(42)));
    layer1_outputs(2403) <= not(layer0_outputs(1253));
    layer1_outputs(2404) <= not(layer0_outputs(3555));
    layer1_outputs(2405) <= '1';
    layer1_outputs(2406) <= not(layer0_outputs(2490)) or (layer0_outputs(2557));
    layer1_outputs(2407) <= (layer0_outputs(2304)) xor (layer0_outputs(3742));
    layer1_outputs(2408) <= layer0_outputs(1435);
    layer1_outputs(2409) <= not((layer0_outputs(3843)) or (layer0_outputs(770)));
    layer1_outputs(2410) <= '0';
    layer1_outputs(2411) <= (layer0_outputs(4426)) and not (layer0_outputs(2674));
    layer1_outputs(2412) <= not(layer0_outputs(3833));
    layer1_outputs(2413) <= layer0_outputs(3407);
    layer1_outputs(2414) <= (layer0_outputs(4275)) or (layer0_outputs(948));
    layer1_outputs(2415) <= not(layer0_outputs(2562)) or (layer0_outputs(994));
    layer1_outputs(2416) <= '0';
    layer1_outputs(2417) <= not((layer0_outputs(3570)) and (layer0_outputs(4624)));
    layer1_outputs(2418) <= not((layer0_outputs(308)) or (layer0_outputs(2816)));
    layer1_outputs(2419) <= '0';
    layer1_outputs(2420) <= not(layer0_outputs(1510)) or (layer0_outputs(4829));
    layer1_outputs(2421) <= not((layer0_outputs(4152)) xor (layer0_outputs(1028)));
    layer1_outputs(2422) <= '1';
    layer1_outputs(2423) <= (layer0_outputs(2808)) and not (layer0_outputs(4310));
    layer1_outputs(2424) <= layer0_outputs(1384);
    layer1_outputs(2425) <= not(layer0_outputs(1534)) or (layer0_outputs(3735));
    layer1_outputs(2426) <= not(layer0_outputs(4595));
    layer1_outputs(2427) <= not(layer0_outputs(4358));
    layer1_outputs(2428) <= not(layer0_outputs(353)) or (layer0_outputs(5056));
    layer1_outputs(2429) <= (layer0_outputs(1296)) or (layer0_outputs(171));
    layer1_outputs(2430) <= '0';
    layer1_outputs(2431) <= (layer0_outputs(3642)) and not (layer0_outputs(4405));
    layer1_outputs(2432) <= (layer0_outputs(776)) or (layer0_outputs(241));
    layer1_outputs(2433) <= (layer0_outputs(3157)) and not (layer0_outputs(2990));
    layer1_outputs(2434) <= (layer0_outputs(1373)) and not (layer0_outputs(2869));
    layer1_outputs(2435) <= layer0_outputs(207);
    layer1_outputs(2436) <= (layer0_outputs(1729)) and (layer0_outputs(1079));
    layer1_outputs(2437) <= (layer0_outputs(2965)) or (layer0_outputs(3018));
    layer1_outputs(2438) <= (layer0_outputs(353)) xor (layer0_outputs(516));
    layer1_outputs(2439) <= '0';
    layer1_outputs(2440) <= '1';
    layer1_outputs(2441) <= (layer0_outputs(3670)) and not (layer0_outputs(898));
    layer1_outputs(2442) <= (layer0_outputs(3900)) and not (layer0_outputs(3251));
    layer1_outputs(2443) <= (layer0_outputs(3185)) or (layer0_outputs(101));
    layer1_outputs(2444) <= layer0_outputs(1925);
    layer1_outputs(2445) <= (layer0_outputs(2848)) or (layer0_outputs(4625));
    layer1_outputs(2446) <= not(layer0_outputs(3954));
    layer1_outputs(2447) <= (layer0_outputs(1662)) and not (layer0_outputs(4599));
    layer1_outputs(2448) <= (layer0_outputs(3906)) and not (layer0_outputs(2127));
    layer1_outputs(2449) <= not(layer0_outputs(304));
    layer1_outputs(2450) <= not((layer0_outputs(2018)) or (layer0_outputs(4988)));
    layer1_outputs(2451) <= not((layer0_outputs(4564)) or (layer0_outputs(22)));
    layer1_outputs(2452) <= not(layer0_outputs(4875)) or (layer0_outputs(3978));
    layer1_outputs(2453) <= not(layer0_outputs(3468));
    layer1_outputs(2454) <= not((layer0_outputs(4250)) or (layer0_outputs(3435)));
    layer1_outputs(2455) <= '0';
    layer1_outputs(2456) <= not(layer0_outputs(2636));
    layer1_outputs(2457) <= (layer0_outputs(4326)) and not (layer0_outputs(3019));
    layer1_outputs(2458) <= not((layer0_outputs(628)) or (layer0_outputs(3772)));
    layer1_outputs(2459) <= '1';
    layer1_outputs(2460) <= (layer0_outputs(3798)) and not (layer0_outputs(2690));
    layer1_outputs(2461) <= not(layer0_outputs(3700)) or (layer0_outputs(3675));
    layer1_outputs(2462) <= not(layer0_outputs(1795));
    layer1_outputs(2463) <= (layer0_outputs(4529)) and not (layer0_outputs(4884));
    layer1_outputs(2464) <= not(layer0_outputs(2379));
    layer1_outputs(2465) <= not(layer0_outputs(4263)) or (layer0_outputs(2684));
    layer1_outputs(2466) <= (layer0_outputs(963)) and not (layer0_outputs(3584));
    layer1_outputs(2467) <= not((layer0_outputs(2228)) and (layer0_outputs(2370)));
    layer1_outputs(2468) <= not(layer0_outputs(483));
    layer1_outputs(2469) <= (layer0_outputs(3361)) and not (layer0_outputs(3447));
    layer1_outputs(2470) <= layer0_outputs(3783);
    layer1_outputs(2471) <= layer0_outputs(508);
    layer1_outputs(2472) <= not((layer0_outputs(862)) and (layer0_outputs(709)));
    layer1_outputs(2473) <= (layer0_outputs(4236)) and not (layer0_outputs(706));
    layer1_outputs(2474) <= (layer0_outputs(5098)) and not (layer0_outputs(1857));
    layer1_outputs(2475) <= '1';
    layer1_outputs(2476) <= (layer0_outputs(3105)) and not (layer0_outputs(2753));
    layer1_outputs(2477) <= not(layer0_outputs(4103));
    layer1_outputs(2478) <= (layer0_outputs(1018)) or (layer0_outputs(2386));
    layer1_outputs(2479) <= (layer0_outputs(1522)) or (layer0_outputs(917));
    layer1_outputs(2480) <= layer0_outputs(4094);
    layer1_outputs(2481) <= (layer0_outputs(223)) and (layer0_outputs(3452));
    layer1_outputs(2482) <= (layer0_outputs(3976)) and not (layer0_outputs(3215));
    layer1_outputs(2483) <= not((layer0_outputs(529)) and (layer0_outputs(2922)));
    layer1_outputs(2484) <= '1';
    layer1_outputs(2485) <= layer0_outputs(3732);
    layer1_outputs(2486) <= layer0_outputs(1345);
    layer1_outputs(2487) <= (layer0_outputs(2199)) and (layer0_outputs(2892));
    layer1_outputs(2488) <= (layer0_outputs(81)) xor (layer0_outputs(3332));
    layer1_outputs(2489) <= layer0_outputs(2506);
    layer1_outputs(2490) <= '1';
    layer1_outputs(2491) <= not((layer0_outputs(5005)) and (layer0_outputs(2474)));
    layer1_outputs(2492) <= (layer0_outputs(3865)) and (layer0_outputs(3542));
    layer1_outputs(2493) <= (layer0_outputs(2596)) and (layer0_outputs(1423));
    layer1_outputs(2494) <= not(layer0_outputs(1047)) or (layer0_outputs(135));
    layer1_outputs(2495) <= (layer0_outputs(1501)) and (layer0_outputs(4199));
    layer1_outputs(2496) <= layer0_outputs(279);
    layer1_outputs(2497) <= '0';
    layer1_outputs(2498) <= layer0_outputs(2380);
    layer1_outputs(2499) <= not(layer0_outputs(1390));
    layer1_outputs(2500) <= not((layer0_outputs(4766)) and (layer0_outputs(4162)));
    layer1_outputs(2501) <= not((layer0_outputs(775)) and (layer0_outputs(4531)));
    layer1_outputs(2502) <= not((layer0_outputs(3736)) or (layer0_outputs(1252)));
    layer1_outputs(2503) <= '1';
    layer1_outputs(2504) <= not(layer0_outputs(2667));
    layer1_outputs(2505) <= (layer0_outputs(391)) and not (layer0_outputs(3239));
    layer1_outputs(2506) <= (layer0_outputs(1098)) and not (layer0_outputs(3130));
    layer1_outputs(2507) <= (layer0_outputs(4733)) and not (layer0_outputs(2768));
    layer1_outputs(2508) <= not(layer0_outputs(1826));
    layer1_outputs(2509) <= '1';
    layer1_outputs(2510) <= (layer0_outputs(587)) xor (layer0_outputs(2415));
    layer1_outputs(2511) <= (layer0_outputs(762)) xor (layer0_outputs(1560));
    layer1_outputs(2512) <= not(layer0_outputs(2987)) or (layer0_outputs(2043));
    layer1_outputs(2513) <= not(layer0_outputs(2850));
    layer1_outputs(2514) <= (layer0_outputs(815)) and (layer0_outputs(1313));
    layer1_outputs(2515) <= (layer0_outputs(3889)) and not (layer0_outputs(4360));
    layer1_outputs(2516) <= layer0_outputs(1229);
    layer1_outputs(2517) <= '0';
    layer1_outputs(2518) <= (layer0_outputs(4888)) and not (layer0_outputs(4796));
    layer1_outputs(2519) <= not((layer0_outputs(2218)) xor (layer0_outputs(446)));
    layer1_outputs(2520) <= not((layer0_outputs(1324)) and (layer0_outputs(5008)));
    layer1_outputs(2521) <= (layer0_outputs(1506)) and not (layer0_outputs(1497));
    layer1_outputs(2522) <= not(layer0_outputs(1755));
    layer1_outputs(2523) <= '1';
    layer1_outputs(2524) <= not((layer0_outputs(2523)) and (layer0_outputs(3182)));
    layer1_outputs(2525) <= not((layer0_outputs(733)) xor (layer0_outputs(2763)));
    layer1_outputs(2526) <= (layer0_outputs(2287)) or (layer0_outputs(1526));
    layer1_outputs(2527) <= (layer0_outputs(303)) and (layer0_outputs(612));
    layer1_outputs(2528) <= (layer0_outputs(614)) and not (layer0_outputs(2868));
    layer1_outputs(2529) <= (layer0_outputs(545)) xor (layer0_outputs(188));
    layer1_outputs(2530) <= (layer0_outputs(1379)) and not (layer0_outputs(3089));
    layer1_outputs(2531) <= not(layer0_outputs(4442));
    layer1_outputs(2532) <= (layer0_outputs(2161)) and not (layer0_outputs(4844));
    layer1_outputs(2533) <= not(layer0_outputs(2913));
    layer1_outputs(2534) <= '1';
    layer1_outputs(2535) <= not(layer0_outputs(2110));
    layer1_outputs(2536) <= (layer0_outputs(4939)) and not (layer0_outputs(871));
    layer1_outputs(2537) <= (layer0_outputs(2559)) or (layer0_outputs(355));
    layer1_outputs(2538) <= not(layer0_outputs(523)) or (layer0_outputs(4047));
    layer1_outputs(2539) <= not(layer0_outputs(3094)) or (layer0_outputs(1204));
    layer1_outputs(2540) <= (layer0_outputs(409)) and not (layer0_outputs(1044));
    layer1_outputs(2541) <= not(layer0_outputs(3587)) or (layer0_outputs(3298));
    layer1_outputs(2542) <= not(layer0_outputs(907)) or (layer0_outputs(2991));
    layer1_outputs(2543) <= '1';
    layer1_outputs(2544) <= not(layer0_outputs(2401));
    layer1_outputs(2545) <= not(layer0_outputs(4709));
    layer1_outputs(2546) <= not(layer0_outputs(1616));
    layer1_outputs(2547) <= '0';
    layer1_outputs(2548) <= (layer0_outputs(2880)) and not (layer0_outputs(3420));
    layer1_outputs(2549) <= (layer0_outputs(855)) and (layer0_outputs(3005));
    layer1_outputs(2550) <= '0';
    layer1_outputs(2551) <= '0';
    layer1_outputs(2552) <= not(layer0_outputs(2955));
    layer1_outputs(2553) <= not((layer0_outputs(2117)) xor (layer0_outputs(3330)));
    layer1_outputs(2554) <= (layer0_outputs(3150)) and not (layer0_outputs(2733));
    layer1_outputs(2555) <= layer0_outputs(4084);
    layer1_outputs(2556) <= not(layer0_outputs(2330));
    layer1_outputs(2557) <= not(layer0_outputs(4339));
    layer1_outputs(2558) <= layer0_outputs(496);
    layer1_outputs(2559) <= not((layer0_outputs(2822)) or (layer0_outputs(1643)));
    layer1_outputs(2560) <= layer0_outputs(4634);
    layer1_outputs(2561) <= not(layer0_outputs(2989)) or (layer0_outputs(4635));
    layer1_outputs(2562) <= '0';
    layer1_outputs(2563) <= (layer0_outputs(817)) and not (layer0_outputs(1195));
    layer1_outputs(2564) <= layer0_outputs(3551);
    layer1_outputs(2565) <= (layer0_outputs(1349)) and not (layer0_outputs(1205));
    layer1_outputs(2566) <= not((layer0_outputs(2314)) or (layer0_outputs(1240)));
    layer1_outputs(2567) <= (layer0_outputs(4129)) or (layer0_outputs(1033));
    layer1_outputs(2568) <= (layer0_outputs(4158)) and not (layer0_outputs(4739));
    layer1_outputs(2569) <= (layer0_outputs(142)) and (layer0_outputs(2946));
    layer1_outputs(2570) <= not(layer0_outputs(70));
    layer1_outputs(2571) <= (layer0_outputs(4344)) or (layer0_outputs(2382));
    layer1_outputs(2572) <= layer0_outputs(3992);
    layer1_outputs(2573) <= not((layer0_outputs(1214)) or (layer0_outputs(597)));
    layer1_outputs(2574) <= not((layer0_outputs(1032)) xor (layer0_outputs(2839)));
    layer1_outputs(2575) <= layer0_outputs(898);
    layer1_outputs(2576) <= not((layer0_outputs(4750)) xor (layer0_outputs(4839)));
    layer1_outputs(2577) <= layer0_outputs(3968);
    layer1_outputs(2578) <= '0';
    layer1_outputs(2579) <= not((layer0_outputs(1720)) and (layer0_outputs(3503)));
    layer1_outputs(2580) <= layer0_outputs(416);
    layer1_outputs(2581) <= not(layer0_outputs(2497)) or (layer0_outputs(160));
    layer1_outputs(2582) <= not(layer0_outputs(2564));
    layer1_outputs(2583) <= not((layer0_outputs(2790)) and (layer0_outputs(2873)));
    layer1_outputs(2584) <= layer0_outputs(4941);
    layer1_outputs(2585) <= '0';
    layer1_outputs(2586) <= not(layer0_outputs(1522));
    layer1_outputs(2587) <= layer0_outputs(3664);
    layer1_outputs(2588) <= not(layer0_outputs(1747));
    layer1_outputs(2589) <= (layer0_outputs(224)) and (layer0_outputs(184));
    layer1_outputs(2590) <= not(layer0_outputs(1376));
    layer1_outputs(2591) <= (layer0_outputs(4077)) and (layer0_outputs(318));
    layer1_outputs(2592) <= not(layer0_outputs(1980));
    layer1_outputs(2593) <= (layer0_outputs(1536)) and (layer0_outputs(361));
    layer1_outputs(2594) <= (layer0_outputs(756)) and (layer0_outputs(388));
    layer1_outputs(2595) <= not((layer0_outputs(742)) or (layer0_outputs(2068)));
    layer1_outputs(2596) <= layer0_outputs(4308);
    layer1_outputs(2597) <= '1';
    layer1_outputs(2598) <= '1';
    layer1_outputs(2599) <= not(layer0_outputs(3836));
    layer1_outputs(2600) <= not((layer0_outputs(2481)) or (layer0_outputs(3591)));
    layer1_outputs(2601) <= (layer0_outputs(2571)) and (layer0_outputs(1485));
    layer1_outputs(2602) <= '1';
    layer1_outputs(2603) <= not(layer0_outputs(1778));
    layer1_outputs(2604) <= '1';
    layer1_outputs(2605) <= not(layer0_outputs(576));
    layer1_outputs(2606) <= not(layer0_outputs(843));
    layer1_outputs(2607) <= not(layer0_outputs(2182)) or (layer0_outputs(2997));
    layer1_outputs(2608) <= layer0_outputs(2453);
    layer1_outputs(2609) <= '1';
    layer1_outputs(2610) <= not(layer0_outputs(3832));
    layer1_outputs(2611) <= layer0_outputs(5011);
    layer1_outputs(2612) <= layer0_outputs(2952);
    layer1_outputs(2613) <= '1';
    layer1_outputs(2614) <= layer0_outputs(4536);
    layer1_outputs(2615) <= (layer0_outputs(466)) and not (layer0_outputs(402));
    layer1_outputs(2616) <= (layer0_outputs(1773)) and not (layer0_outputs(4435));
    layer1_outputs(2617) <= not(layer0_outputs(2136));
    layer1_outputs(2618) <= '1';
    layer1_outputs(2619) <= '1';
    layer1_outputs(2620) <= not(layer0_outputs(3348)) or (layer0_outputs(4392));
    layer1_outputs(2621) <= (layer0_outputs(4701)) and not (layer0_outputs(1250));
    layer1_outputs(2622) <= (layer0_outputs(3136)) and not (layer0_outputs(976));
    layer1_outputs(2623) <= (layer0_outputs(4753)) and not (layer0_outputs(3011));
    layer1_outputs(2624) <= layer0_outputs(4893);
    layer1_outputs(2625) <= not(layer0_outputs(3962)) or (layer0_outputs(2505));
    layer1_outputs(2626) <= not(layer0_outputs(2205)) or (layer0_outputs(3835));
    layer1_outputs(2627) <= layer0_outputs(4242);
    layer1_outputs(2628) <= (layer0_outputs(1319)) or (layer0_outputs(1835));
    layer1_outputs(2629) <= not(layer0_outputs(3545)) or (layer0_outputs(511));
    layer1_outputs(2630) <= not(layer0_outputs(1896));
    layer1_outputs(2631) <= not(layer0_outputs(3494)) or (layer0_outputs(1308));
    layer1_outputs(2632) <= not(layer0_outputs(2579)) or (layer0_outputs(2709));
    layer1_outputs(2633) <= not(layer0_outputs(1946));
    layer1_outputs(2634) <= (layer0_outputs(3497)) and (layer0_outputs(1128));
    layer1_outputs(2635) <= not(layer0_outputs(2639));
    layer1_outputs(2636) <= layer0_outputs(2825);
    layer1_outputs(2637) <= (layer0_outputs(4154)) and (layer0_outputs(4215));
    layer1_outputs(2638) <= (layer0_outputs(306)) and not (layer0_outputs(1458));
    layer1_outputs(2639) <= (layer0_outputs(9)) and not (layer0_outputs(2767));
    layer1_outputs(2640) <= (layer0_outputs(1160)) or (layer0_outputs(3669));
    layer1_outputs(2641) <= '1';
    layer1_outputs(2642) <= (layer0_outputs(4666)) and not (layer0_outputs(4320));
    layer1_outputs(2643) <= not(layer0_outputs(3682)) or (layer0_outputs(4896));
    layer1_outputs(2644) <= (layer0_outputs(1585)) or (layer0_outputs(4922));
    layer1_outputs(2645) <= not((layer0_outputs(1017)) and (layer0_outputs(2772)));
    layer1_outputs(2646) <= (layer0_outputs(1867)) and not (layer0_outputs(4034));
    layer1_outputs(2647) <= not((layer0_outputs(1802)) or (layer0_outputs(1856)));
    layer1_outputs(2648) <= layer0_outputs(874);
    layer1_outputs(2649) <= layer0_outputs(2938);
    layer1_outputs(2650) <= (layer0_outputs(3114)) and (layer0_outputs(3091));
    layer1_outputs(2651) <= '1';
    layer1_outputs(2652) <= '1';
    layer1_outputs(2653) <= '1';
    layer1_outputs(2654) <= not((layer0_outputs(3533)) and (layer0_outputs(1524)));
    layer1_outputs(2655) <= '0';
    layer1_outputs(2656) <= not(layer0_outputs(4105));
    layer1_outputs(2657) <= layer0_outputs(1482);
    layer1_outputs(2658) <= (layer0_outputs(1129)) or (layer0_outputs(4328));
    layer1_outputs(2659) <= not((layer0_outputs(4839)) and (layer0_outputs(2298)));
    layer1_outputs(2660) <= not((layer0_outputs(2214)) or (layer0_outputs(2728)));
    layer1_outputs(2661) <= '0';
    layer1_outputs(2662) <= (layer0_outputs(1056)) and not (layer0_outputs(3508));
    layer1_outputs(2663) <= not((layer0_outputs(125)) or (layer0_outputs(2893)));
    layer1_outputs(2664) <= (layer0_outputs(4743)) and (layer0_outputs(1771));
    layer1_outputs(2665) <= not(layer0_outputs(2510));
    layer1_outputs(2666) <= layer0_outputs(5114);
    layer1_outputs(2667) <= layer0_outputs(4797);
    layer1_outputs(2668) <= layer0_outputs(4396);
    layer1_outputs(2669) <= not((layer0_outputs(3511)) or (layer0_outputs(953)));
    layer1_outputs(2670) <= not(layer0_outputs(3339)) or (layer0_outputs(5030));
    layer1_outputs(2671) <= not(layer0_outputs(888));
    layer1_outputs(2672) <= not(layer0_outputs(4788));
    layer1_outputs(2673) <= not(layer0_outputs(2209)) or (layer0_outputs(3441));
    layer1_outputs(2674) <= (layer0_outputs(969)) and (layer0_outputs(662));
    layer1_outputs(2675) <= not(layer0_outputs(777));
    layer1_outputs(2676) <= not(layer0_outputs(3132));
    layer1_outputs(2677) <= (layer0_outputs(705)) and not (layer0_outputs(1367));
    layer1_outputs(2678) <= (layer0_outputs(4505)) and not (layer0_outputs(3776));
    layer1_outputs(2679) <= not((layer0_outputs(1479)) or (layer0_outputs(849)));
    layer1_outputs(2680) <= not((layer0_outputs(2985)) and (layer0_outputs(4348)));
    layer1_outputs(2681) <= not((layer0_outputs(880)) xor (layer0_outputs(2428)));
    layer1_outputs(2682) <= '0';
    layer1_outputs(2683) <= (layer0_outputs(4635)) and not (layer0_outputs(823));
    layer1_outputs(2684) <= (layer0_outputs(2435)) or (layer0_outputs(2271));
    layer1_outputs(2685) <= layer0_outputs(346);
    layer1_outputs(2686) <= not(layer0_outputs(5066)) or (layer0_outputs(4172));
    layer1_outputs(2687) <= not(layer0_outputs(1836)) or (layer0_outputs(4975));
    layer1_outputs(2688) <= '1';
    layer1_outputs(2689) <= '1';
    layer1_outputs(2690) <= not((layer0_outputs(635)) and (layer0_outputs(4735)));
    layer1_outputs(2691) <= not(layer0_outputs(3583));
    layer1_outputs(2692) <= '0';
    layer1_outputs(2693) <= not(layer0_outputs(730));
    layer1_outputs(2694) <= not((layer0_outputs(2097)) and (layer0_outputs(2531)));
    layer1_outputs(2695) <= (layer0_outputs(2486)) and not (layer0_outputs(5094));
    layer1_outputs(2696) <= layer0_outputs(3703);
    layer1_outputs(2697) <= '0';
    layer1_outputs(2698) <= not(layer0_outputs(4205));
    layer1_outputs(2699) <= (layer0_outputs(3858)) and not (layer0_outputs(3368));
    layer1_outputs(2700) <= '1';
    layer1_outputs(2701) <= (layer0_outputs(4581)) and not (layer0_outputs(617));
    layer1_outputs(2702) <= (layer0_outputs(4523)) and not (layer0_outputs(2219));
    layer1_outputs(2703) <= (layer0_outputs(4230)) and not (layer0_outputs(2644));
    layer1_outputs(2704) <= not((layer0_outputs(4991)) and (layer0_outputs(1432)));
    layer1_outputs(2705) <= (layer0_outputs(4078)) or (layer0_outputs(467));
    layer1_outputs(2706) <= not(layer0_outputs(2805)) or (layer0_outputs(1196));
    layer1_outputs(2707) <= '0';
    layer1_outputs(2708) <= not(layer0_outputs(1273));
    layer1_outputs(2709) <= (layer0_outputs(2255)) and (layer0_outputs(5043));
    layer1_outputs(2710) <= not((layer0_outputs(1660)) or (layer0_outputs(3919)));
    layer1_outputs(2711) <= layer0_outputs(2310);
    layer1_outputs(2712) <= '1';
    layer1_outputs(2713) <= (layer0_outputs(4566)) and (layer0_outputs(578));
    layer1_outputs(2714) <= (layer0_outputs(3995)) or (layer0_outputs(1039));
    layer1_outputs(2715) <= not((layer0_outputs(3829)) or (layer0_outputs(5053)));
    layer1_outputs(2716) <= not(layer0_outputs(2075));
    layer1_outputs(2717) <= not(layer0_outputs(1891)) or (layer0_outputs(3781));
    layer1_outputs(2718) <= (layer0_outputs(3889)) and not (layer0_outputs(4221));
    layer1_outputs(2719) <= not(layer0_outputs(181)) or (layer0_outputs(4754));
    layer1_outputs(2720) <= (layer0_outputs(3163)) and not (layer0_outputs(3296));
    layer1_outputs(2721) <= not(layer0_outputs(105));
    layer1_outputs(2722) <= '1';
    layer1_outputs(2723) <= (layer0_outputs(2560)) and (layer0_outputs(2403));
    layer1_outputs(2724) <= '1';
    layer1_outputs(2725) <= not((layer0_outputs(1115)) or (layer0_outputs(2707)));
    layer1_outputs(2726) <= layer0_outputs(1364);
    layer1_outputs(2727) <= '1';
    layer1_outputs(2728) <= layer0_outputs(4470);
    layer1_outputs(2729) <= '0';
    layer1_outputs(2730) <= not((layer0_outputs(3769)) or (layer0_outputs(2268)));
    layer1_outputs(2731) <= layer0_outputs(143);
    layer1_outputs(2732) <= (layer0_outputs(549)) and (layer0_outputs(189));
    layer1_outputs(2733) <= (layer0_outputs(1665)) or (layer0_outputs(543));
    layer1_outputs(2734) <= not(layer0_outputs(4097)) or (layer0_outputs(3242));
    layer1_outputs(2735) <= not(layer0_outputs(3536));
    layer1_outputs(2736) <= not(layer0_outputs(916));
    layer1_outputs(2737) <= not((layer0_outputs(495)) or (layer0_outputs(2563)));
    layer1_outputs(2738) <= layer0_outputs(2742);
    layer1_outputs(2739) <= (layer0_outputs(1727)) and not (layer0_outputs(4865));
    layer1_outputs(2740) <= '0';
    layer1_outputs(2741) <= '0';
    layer1_outputs(2742) <= not((layer0_outputs(1577)) and (layer0_outputs(4906)));
    layer1_outputs(2743) <= layer0_outputs(3373);
    layer1_outputs(2744) <= layer0_outputs(4537);
    layer1_outputs(2745) <= not(layer0_outputs(669)) or (layer0_outputs(1926));
    layer1_outputs(2746) <= layer0_outputs(2536);
    layer1_outputs(2747) <= not(layer0_outputs(611)) or (layer0_outputs(263));
    layer1_outputs(2748) <= '1';
    layer1_outputs(2749) <= layer0_outputs(2382);
    layer1_outputs(2750) <= not(layer0_outputs(606)) or (layer0_outputs(39));
    layer1_outputs(2751) <= (layer0_outputs(2033)) and not (layer0_outputs(2348));
    layer1_outputs(2752) <= (layer0_outputs(2803)) and not (layer0_outputs(3967));
    layer1_outputs(2753) <= (layer0_outputs(2390)) and not (layer0_outputs(1744));
    layer1_outputs(2754) <= (layer0_outputs(4917)) and (layer0_outputs(2556));
    layer1_outputs(2755) <= (layer0_outputs(1064)) xor (layer0_outputs(2480));
    layer1_outputs(2756) <= '1';
    layer1_outputs(2757) <= not(layer0_outputs(4994)) or (layer0_outputs(2852));
    layer1_outputs(2758) <= not((layer0_outputs(2618)) and (layer0_outputs(608)));
    layer1_outputs(2759) <= not((layer0_outputs(2170)) xor (layer0_outputs(4643)));
    layer1_outputs(2760) <= (layer0_outputs(2784)) or (layer0_outputs(4920));
    layer1_outputs(2761) <= not((layer0_outputs(3562)) or (layer0_outputs(1524)));
    layer1_outputs(2762) <= '0';
    layer1_outputs(2763) <= '0';
    layer1_outputs(2764) <= not(layer0_outputs(3706));
    layer1_outputs(2765) <= '0';
    layer1_outputs(2766) <= not((layer0_outputs(823)) and (layer0_outputs(4255)));
    layer1_outputs(2767) <= not(layer0_outputs(4015)) or (layer0_outputs(1290));
    layer1_outputs(2768) <= (layer0_outputs(691)) and not (layer0_outputs(2441));
    layer1_outputs(2769) <= '0';
    layer1_outputs(2770) <= (layer0_outputs(373)) and not (layer0_outputs(1552));
    layer1_outputs(2771) <= not((layer0_outputs(3988)) or (layer0_outputs(1981)));
    layer1_outputs(2772) <= '1';
    layer1_outputs(2773) <= (layer0_outputs(1975)) and not (layer0_outputs(426));
    layer1_outputs(2774) <= (layer0_outputs(3381)) and not (layer0_outputs(1708));
    layer1_outputs(2775) <= (layer0_outputs(1968)) and (layer0_outputs(4247));
    layer1_outputs(2776) <= (layer0_outputs(1586)) and not (layer0_outputs(759));
    layer1_outputs(2777) <= '1';
    layer1_outputs(2778) <= (layer0_outputs(4561)) and not (layer0_outputs(3336));
    layer1_outputs(2779) <= not((layer0_outputs(3808)) or (layer0_outputs(676)));
    layer1_outputs(2780) <= not(layer0_outputs(2634));
    layer1_outputs(2781) <= not(layer0_outputs(4255)) or (layer0_outputs(5042));
    layer1_outputs(2782) <= '0';
    layer1_outputs(2783) <= layer0_outputs(1884);
    layer1_outputs(2784) <= layer0_outputs(2358);
    layer1_outputs(2785) <= not(layer0_outputs(2661));
    layer1_outputs(2786) <= (layer0_outputs(1698)) xor (layer0_outputs(3231));
    layer1_outputs(2787) <= not(layer0_outputs(3574)) or (layer0_outputs(25));
    layer1_outputs(2788) <= not(layer0_outputs(485)) or (layer0_outputs(4284));
    layer1_outputs(2789) <= layer0_outputs(554);
    layer1_outputs(2790) <= (layer0_outputs(3830)) or (layer0_outputs(3277));
    layer1_outputs(2791) <= (layer0_outputs(4910)) and (layer0_outputs(4502));
    layer1_outputs(2792) <= (layer0_outputs(1032)) and not (layer0_outputs(4513));
    layer1_outputs(2793) <= '0';
    layer1_outputs(2794) <= (layer0_outputs(2672)) and (layer0_outputs(1105));
    layer1_outputs(2795) <= not((layer0_outputs(472)) and (layer0_outputs(3038)));
    layer1_outputs(2796) <= '0';
    layer1_outputs(2797) <= layer0_outputs(3027);
    layer1_outputs(2798) <= layer0_outputs(4379);
    layer1_outputs(2799) <= not(layer0_outputs(1223));
    layer1_outputs(2800) <= not(layer0_outputs(4588));
    layer1_outputs(2801) <= (layer0_outputs(892)) and not (layer0_outputs(4849));
    layer1_outputs(2802) <= '1';
    layer1_outputs(2803) <= '1';
    layer1_outputs(2804) <= not(layer0_outputs(3757)) or (layer0_outputs(2566));
    layer1_outputs(2805) <= not(layer0_outputs(3360));
    layer1_outputs(2806) <= (layer0_outputs(762)) and (layer0_outputs(1339));
    layer1_outputs(2807) <= (layer0_outputs(164)) and (layer0_outputs(297));
    layer1_outputs(2808) <= '0';
    layer1_outputs(2809) <= not(layer0_outputs(2928)) or (layer0_outputs(3336));
    layer1_outputs(2810) <= (layer0_outputs(3311)) and (layer0_outputs(4238));
    layer1_outputs(2811) <= layer0_outputs(2716);
    layer1_outputs(2812) <= not((layer0_outputs(4627)) and (layer0_outputs(4628)));
    layer1_outputs(2813) <= layer0_outputs(2660);
    layer1_outputs(2814) <= not(layer0_outputs(1284)) or (layer0_outputs(2569));
    layer1_outputs(2815) <= layer0_outputs(2697);
    layer1_outputs(2816) <= layer0_outputs(1573);
    layer1_outputs(2817) <= (layer0_outputs(676)) and not (layer0_outputs(4414));
    layer1_outputs(2818) <= layer0_outputs(908);
    layer1_outputs(2819) <= not(layer0_outputs(3493)) or (layer0_outputs(1429));
    layer1_outputs(2820) <= (layer0_outputs(481)) and (layer0_outputs(1142));
    layer1_outputs(2821) <= layer0_outputs(3499);
    layer1_outputs(2822) <= '0';
    layer1_outputs(2823) <= not(layer0_outputs(4978));
    layer1_outputs(2824) <= (layer0_outputs(4116)) and (layer0_outputs(531));
    layer1_outputs(2825) <= not((layer0_outputs(4380)) and (layer0_outputs(1685)));
    layer1_outputs(2826) <= layer0_outputs(3032);
    layer1_outputs(2827) <= not(layer0_outputs(519));
    layer1_outputs(2828) <= not(layer0_outputs(366));
    layer1_outputs(2829) <= (layer0_outputs(1592)) or (layer0_outputs(1181));
    layer1_outputs(2830) <= not(layer0_outputs(1317)) or (layer0_outputs(3807));
    layer1_outputs(2831) <= not(layer0_outputs(1149));
    layer1_outputs(2832) <= not(layer0_outputs(2606));
    layer1_outputs(2833) <= layer0_outputs(571);
    layer1_outputs(2834) <= not((layer0_outputs(900)) and (layer0_outputs(2074)));
    layer1_outputs(2835) <= not(layer0_outputs(1250));
    layer1_outputs(2836) <= not((layer0_outputs(954)) or (layer0_outputs(2183)));
    layer1_outputs(2837) <= (layer0_outputs(3530)) and (layer0_outputs(2996));
    layer1_outputs(2838) <= not(layer0_outputs(3127));
    layer1_outputs(2839) <= (layer0_outputs(2491)) and (layer0_outputs(4534));
    layer1_outputs(2840) <= (layer0_outputs(4863)) and not (layer0_outputs(2157));
    layer1_outputs(2841) <= not(layer0_outputs(2790));
    layer1_outputs(2842) <= not(layer0_outputs(3192));
    layer1_outputs(2843) <= not((layer0_outputs(3726)) and (layer0_outputs(3394)));
    layer1_outputs(2844) <= (layer0_outputs(832)) and not (layer0_outputs(3177));
    layer1_outputs(2845) <= (layer0_outputs(2932)) or (layer0_outputs(3309));
    layer1_outputs(2846) <= not(layer0_outputs(987));
    layer1_outputs(2847) <= (layer0_outputs(2688)) and not (layer0_outputs(1185));
    layer1_outputs(2848) <= '0';
    layer1_outputs(2849) <= not(layer0_outputs(4738));
    layer1_outputs(2850) <= '0';
    layer1_outputs(2851) <= layer0_outputs(3158);
    layer1_outputs(2852) <= not((layer0_outputs(1865)) or (layer0_outputs(425)));
    layer1_outputs(2853) <= not(layer0_outputs(3539));
    layer1_outputs(2854) <= not(layer0_outputs(3949)) or (layer0_outputs(640));
    layer1_outputs(2855) <= layer0_outputs(1635);
    layer1_outputs(2856) <= layer0_outputs(1024);
    layer1_outputs(2857) <= not(layer0_outputs(4164)) or (layer0_outputs(152));
    layer1_outputs(2858) <= not((layer0_outputs(4027)) or (layer0_outputs(3879)));
    layer1_outputs(2859) <= (layer0_outputs(4216)) and not (layer0_outputs(4488));
    layer1_outputs(2860) <= (layer0_outputs(3451)) and not (layer0_outputs(2793));
    layer1_outputs(2861) <= (layer0_outputs(3120)) and not (layer0_outputs(4558));
    layer1_outputs(2862) <= not((layer0_outputs(2497)) and (layer0_outputs(37)));
    layer1_outputs(2863) <= not((layer0_outputs(2929)) or (layer0_outputs(4521)));
    layer1_outputs(2864) <= layer0_outputs(4024);
    layer1_outputs(2865) <= '1';
    layer1_outputs(2866) <= not((layer0_outputs(1617)) or (layer0_outputs(4031)));
    layer1_outputs(2867) <= not((layer0_outputs(471)) or (layer0_outputs(4877)));
    layer1_outputs(2868) <= not(layer0_outputs(3245)) or (layer0_outputs(146));
    layer1_outputs(2869) <= '0';
    layer1_outputs(2870) <= (layer0_outputs(1121)) and not (layer0_outputs(4997));
    layer1_outputs(2871) <= layer0_outputs(443);
    layer1_outputs(2872) <= '0';
    layer1_outputs(2873) <= (layer0_outputs(4940)) and not (layer0_outputs(2446));
    layer1_outputs(2874) <= (layer0_outputs(636)) and not (layer0_outputs(1628));
    layer1_outputs(2875) <= (layer0_outputs(1831)) or (layer0_outputs(1907));
    layer1_outputs(2876) <= not(layer0_outputs(3936));
    layer1_outputs(2877) <= not(layer0_outputs(1844)) or (layer0_outputs(2983));
    layer1_outputs(2878) <= not(layer0_outputs(1413)) or (layer0_outputs(3221));
    layer1_outputs(2879) <= not((layer0_outputs(2319)) and (layer0_outputs(4142)));
    layer1_outputs(2880) <= layer0_outputs(289);
    layer1_outputs(2881) <= '0';
    layer1_outputs(2882) <= not(layer0_outputs(1648)) or (layer0_outputs(3797));
    layer1_outputs(2883) <= layer0_outputs(1203);
    layer1_outputs(2884) <= not((layer0_outputs(850)) and (layer0_outputs(359)));
    layer1_outputs(2885) <= not((layer0_outputs(3960)) or (layer0_outputs(3540)));
    layer1_outputs(2886) <= layer0_outputs(326);
    layer1_outputs(2887) <= '0';
    layer1_outputs(2888) <= not(layer0_outputs(162));
    layer1_outputs(2889) <= (layer0_outputs(3172)) or (layer0_outputs(1124));
    layer1_outputs(2890) <= not((layer0_outputs(4690)) or (layer0_outputs(116)));
    layer1_outputs(2891) <= '1';
    layer1_outputs(2892) <= not((layer0_outputs(2061)) or (layer0_outputs(5006)));
    layer1_outputs(2893) <= '0';
    layer1_outputs(2894) <= '0';
    layer1_outputs(2895) <= '0';
    layer1_outputs(2896) <= layer0_outputs(3966);
    layer1_outputs(2897) <= not((layer0_outputs(220)) or (layer0_outputs(3127)));
    layer1_outputs(2898) <= (layer0_outputs(2408)) and not (layer0_outputs(1373));
    layer1_outputs(2899) <= '0';
    layer1_outputs(2900) <= '1';
    layer1_outputs(2901) <= not(layer0_outputs(4670)) or (layer0_outputs(3568));
    layer1_outputs(2902) <= (layer0_outputs(1983)) xor (layer0_outputs(4528));
    layer1_outputs(2903) <= not(layer0_outputs(3786)) or (layer0_outputs(2739));
    layer1_outputs(2904) <= (layer0_outputs(2266)) or (layer0_outputs(3559));
    layer1_outputs(2905) <= (layer0_outputs(4843)) or (layer0_outputs(3066));
    layer1_outputs(2906) <= not(layer0_outputs(637));
    layer1_outputs(2907) <= (layer0_outputs(4901)) and not (layer0_outputs(876));
    layer1_outputs(2908) <= not(layer0_outputs(3862));
    layer1_outputs(2909) <= layer0_outputs(3052);
    layer1_outputs(2910) <= layer0_outputs(2478);
    layer1_outputs(2911) <= layer0_outputs(1645);
    layer1_outputs(2912) <= '1';
    layer1_outputs(2913) <= not(layer0_outputs(2419));
    layer1_outputs(2914) <= not(layer0_outputs(3469));
    layer1_outputs(2915) <= '1';
    layer1_outputs(2916) <= '0';
    layer1_outputs(2917) <= (layer0_outputs(1387)) and not (layer0_outputs(4683));
    layer1_outputs(2918) <= not((layer0_outputs(4995)) and (layer0_outputs(3489)));
    layer1_outputs(2919) <= (layer0_outputs(4068)) and not (layer0_outputs(2458));
    layer1_outputs(2920) <= layer0_outputs(3254);
    layer1_outputs(2921) <= not(layer0_outputs(1420));
    layer1_outputs(2922) <= not((layer0_outputs(1663)) and (layer0_outputs(1401)));
    layer1_outputs(2923) <= not(layer0_outputs(2576)) or (layer0_outputs(1415));
    layer1_outputs(2924) <= not((layer0_outputs(1186)) or (layer0_outputs(1090)));
    layer1_outputs(2925) <= not((layer0_outputs(2118)) or (layer0_outputs(2077)));
    layer1_outputs(2926) <= not(layer0_outputs(4276));
    layer1_outputs(2927) <= (layer0_outputs(4534)) or (layer0_outputs(4262));
    layer1_outputs(2928) <= not(layer0_outputs(2588));
    layer1_outputs(2929) <= (layer0_outputs(4411)) and not (layer0_outputs(1165));
    layer1_outputs(2930) <= not((layer0_outputs(4833)) and (layer0_outputs(3934)));
    layer1_outputs(2931) <= (layer0_outputs(4978)) and not (layer0_outputs(4234));
    layer1_outputs(2932) <= not(layer0_outputs(5062));
    layer1_outputs(2933) <= '0';
    layer1_outputs(2934) <= '0';
    layer1_outputs(2935) <= '1';
    layer1_outputs(2936) <= (layer0_outputs(4465)) xor (layer0_outputs(1286));
    layer1_outputs(2937) <= '1';
    layer1_outputs(2938) <= not((layer0_outputs(1716)) or (layer0_outputs(4687)));
    layer1_outputs(2939) <= layer0_outputs(1744);
    layer1_outputs(2940) <= not(layer0_outputs(2369));
    layer1_outputs(2941) <= layer0_outputs(4496);
    layer1_outputs(2942) <= not(layer0_outputs(2971)) or (layer0_outputs(4990));
    layer1_outputs(2943) <= '1';
    layer1_outputs(2944) <= (layer0_outputs(3337)) and not (layer0_outputs(2132));
    layer1_outputs(2945) <= not(layer0_outputs(3367));
    layer1_outputs(2946) <= '1';
    layer1_outputs(2947) <= (layer0_outputs(3674)) and not (layer0_outputs(148));
    layer1_outputs(2948) <= '0';
    layer1_outputs(2949) <= layer0_outputs(4972);
    layer1_outputs(2950) <= layer0_outputs(4286);
    layer1_outputs(2951) <= (layer0_outputs(3929)) and not (layer0_outputs(5075));
    layer1_outputs(2952) <= '0';
    layer1_outputs(2953) <= (layer0_outputs(3990)) and (layer0_outputs(4096));
    layer1_outputs(2954) <= not((layer0_outputs(2101)) or (layer0_outputs(2254)));
    layer1_outputs(2955) <= (layer0_outputs(3475)) and not (layer0_outputs(1283));
    layer1_outputs(2956) <= not(layer0_outputs(2555)) or (layer0_outputs(970));
    layer1_outputs(2957) <= '1';
    layer1_outputs(2958) <= (layer0_outputs(2851)) and not (layer0_outputs(4092));
    layer1_outputs(2959) <= layer0_outputs(586);
    layer1_outputs(2960) <= (layer0_outputs(4989)) and not (layer0_outputs(3612));
    layer1_outputs(2961) <= (layer0_outputs(3517)) and not (layer0_outputs(3468));
    layer1_outputs(2962) <= '0';
    layer1_outputs(2963) <= (layer0_outputs(4259)) or (layer0_outputs(4111));
    layer1_outputs(2964) <= layer0_outputs(1362);
    layer1_outputs(2965) <= (layer0_outputs(5057)) and (layer0_outputs(2897));
    layer1_outputs(2966) <= (layer0_outputs(7)) and (layer0_outputs(4897));
    layer1_outputs(2967) <= (layer0_outputs(1789)) and not (layer0_outputs(2908));
    layer1_outputs(2968) <= layer0_outputs(1935);
    layer1_outputs(2969) <= (layer0_outputs(2476)) or (layer0_outputs(2558));
    layer1_outputs(2970) <= '1';
    layer1_outputs(2971) <= layer0_outputs(4436);
    layer1_outputs(2972) <= not(layer0_outputs(1253));
    layer1_outputs(2973) <= (layer0_outputs(5047)) xor (layer0_outputs(3918));
    layer1_outputs(2974) <= '1';
    layer1_outputs(2975) <= (layer0_outputs(2859)) or (layer0_outputs(134));
    layer1_outputs(2976) <= (layer0_outputs(771)) and (layer0_outputs(538));
    layer1_outputs(2977) <= not(layer0_outputs(1140)) or (layer0_outputs(475));
    layer1_outputs(2978) <= (layer0_outputs(4660)) and not (layer0_outputs(1145));
    layer1_outputs(2979) <= layer0_outputs(4717);
    layer1_outputs(2980) <= not(layer0_outputs(2514));
    layer1_outputs(2981) <= not(layer0_outputs(1940));
    layer1_outputs(2982) <= not(layer0_outputs(1705));
    layer1_outputs(2983) <= not(layer0_outputs(4166));
    layer1_outputs(2984) <= not((layer0_outputs(2811)) or (layer0_outputs(446)));
    layer1_outputs(2985) <= not(layer0_outputs(4037));
    layer1_outputs(2986) <= not(layer0_outputs(5073));
    layer1_outputs(2987) <= not((layer0_outputs(1428)) and (layer0_outputs(2670)));
    layer1_outputs(2988) <= '1';
    layer1_outputs(2989) <= not((layer0_outputs(4672)) xor (layer0_outputs(4829)));
    layer1_outputs(2990) <= not((layer0_outputs(3625)) or (layer0_outputs(1904)));
    layer1_outputs(2991) <= (layer0_outputs(2169)) and not (layer0_outputs(4445));
    layer1_outputs(2992) <= (layer0_outputs(3069)) or (layer0_outputs(3581));
    layer1_outputs(2993) <= layer0_outputs(3690);
    layer1_outputs(2994) <= not(layer0_outputs(3158)) or (layer0_outputs(2437));
    layer1_outputs(2995) <= layer0_outputs(4123);
    layer1_outputs(2996) <= layer0_outputs(3855);
    layer1_outputs(2997) <= not((layer0_outputs(420)) and (layer0_outputs(2045)));
    layer1_outputs(2998) <= not((layer0_outputs(168)) or (layer0_outputs(447)));
    layer1_outputs(2999) <= layer0_outputs(4059);
    layer1_outputs(3000) <= (layer0_outputs(3621)) and not (layer0_outputs(2313));
    layer1_outputs(3001) <= not(layer0_outputs(347)) or (layer0_outputs(3424));
    layer1_outputs(3002) <= (layer0_outputs(3565)) or (layer0_outputs(5113));
    layer1_outputs(3003) <= layer0_outputs(112);
    layer1_outputs(3004) <= not(layer0_outputs(619)) or (layer0_outputs(2256));
    layer1_outputs(3005) <= layer0_outputs(2338);
    layer1_outputs(3006) <= '1';
    layer1_outputs(3007) <= layer0_outputs(4374);
    layer1_outputs(3008) <= '0';
    layer1_outputs(3009) <= not(layer0_outputs(392));
    layer1_outputs(3010) <= not(layer0_outputs(3433));
    layer1_outputs(3011) <= layer0_outputs(3708);
    layer1_outputs(3012) <= layer0_outputs(4543);
    layer1_outputs(3013) <= not(layer0_outputs(3559));
    layer1_outputs(3014) <= not(layer0_outputs(2176)) or (layer0_outputs(47));
    layer1_outputs(3015) <= (layer0_outputs(949)) and not (layer0_outputs(1655));
    layer1_outputs(3016) <= '0';
    layer1_outputs(3017) <= layer0_outputs(2890);
    layer1_outputs(3018) <= '0';
    layer1_outputs(3019) <= layer0_outputs(4892);
    layer1_outputs(3020) <= (layer0_outputs(2813)) and not (layer0_outputs(3748));
    layer1_outputs(3021) <= (layer0_outputs(4669)) and not (layer0_outputs(2432));
    layer1_outputs(3022) <= layer0_outputs(1525);
    layer1_outputs(3023) <= not(layer0_outputs(3964)) or (layer0_outputs(1431));
    layer1_outputs(3024) <= not(layer0_outputs(4374));
    layer1_outputs(3025) <= not(layer0_outputs(2160)) or (layer0_outputs(1120));
    layer1_outputs(3026) <= (layer0_outputs(2267)) and not (layer0_outputs(4693));
    layer1_outputs(3027) <= layer0_outputs(1753);
    layer1_outputs(3028) <= '0';
    layer1_outputs(3029) <= (layer0_outputs(1652)) and (layer0_outputs(1318));
    layer1_outputs(3030) <= (layer0_outputs(1883)) and (layer0_outputs(3411));
    layer1_outputs(3031) <= (layer0_outputs(5093)) or (layer0_outputs(3906));
    layer1_outputs(3032) <= (layer0_outputs(2721)) and not (layer0_outputs(2896));
    layer1_outputs(3033) <= not(layer0_outputs(1)) or (layer0_outputs(1243));
    layer1_outputs(3034) <= (layer0_outputs(958)) and not (layer0_outputs(699));
    layer1_outputs(3035) <= not((layer0_outputs(1693)) and (layer0_outputs(381)));
    layer1_outputs(3036) <= layer0_outputs(586);
    layer1_outputs(3037) <= (layer0_outputs(312)) and (layer0_outputs(4798));
    layer1_outputs(3038) <= layer0_outputs(2597);
    layer1_outputs(3039) <= layer0_outputs(3734);
    layer1_outputs(3040) <= not((layer0_outputs(1608)) and (layer0_outputs(1101)));
    layer1_outputs(3041) <= not(layer0_outputs(1707));
    layer1_outputs(3042) <= not(layer0_outputs(2194)) or (layer0_outputs(1239));
    layer1_outputs(3043) <= not(layer0_outputs(4400));
    layer1_outputs(3044) <= '1';
    layer1_outputs(3045) <= layer0_outputs(844);
    layer1_outputs(3046) <= '0';
    layer1_outputs(3047) <= not(layer0_outputs(540)) or (layer0_outputs(5088));
    layer1_outputs(3048) <= not(layer0_outputs(2898));
    layer1_outputs(3049) <= layer0_outputs(1030);
    layer1_outputs(3050) <= not(layer0_outputs(275)) or (layer0_outputs(3174));
    layer1_outputs(3051) <= (layer0_outputs(126)) or (layer0_outputs(2904));
    layer1_outputs(3052) <= (layer0_outputs(1350)) or (layer0_outputs(981));
    layer1_outputs(3053) <= layer0_outputs(633);
    layer1_outputs(3054) <= not(layer0_outputs(3351)) or (layer0_outputs(4609));
    layer1_outputs(3055) <= not((layer0_outputs(4324)) or (layer0_outputs(4810)));
    layer1_outputs(3056) <= not(layer0_outputs(2647));
    layer1_outputs(3057) <= (layer0_outputs(66)) and not (layer0_outputs(559));
    layer1_outputs(3058) <= (layer0_outputs(3297)) and (layer0_outputs(1714));
    layer1_outputs(3059) <= not(layer0_outputs(4867)) or (layer0_outputs(1072));
    layer1_outputs(3060) <= not((layer0_outputs(1997)) or (layer0_outputs(2267)));
    layer1_outputs(3061) <= layer0_outputs(3911);
    layer1_outputs(3062) <= '1';
    layer1_outputs(3063) <= layer0_outputs(314);
    layer1_outputs(3064) <= not(layer0_outputs(3678)) or (layer0_outputs(2681));
    layer1_outputs(3065) <= not((layer0_outputs(4746)) or (layer0_outputs(1200)));
    layer1_outputs(3066) <= not(layer0_outputs(1320)) or (layer0_outputs(1658));
    layer1_outputs(3067) <= (layer0_outputs(448)) and not (layer0_outputs(4600));
    layer1_outputs(3068) <= not(layer0_outputs(2831));
    layer1_outputs(3069) <= '1';
    layer1_outputs(3070) <= (layer0_outputs(4399)) and not (layer0_outputs(680));
    layer1_outputs(3071) <= '1';
    layer1_outputs(3072) <= not(layer0_outputs(4894)) or (layer0_outputs(1645));
    layer1_outputs(3073) <= (layer0_outputs(3244)) or (layer0_outputs(20));
    layer1_outputs(3074) <= not(layer0_outputs(2472)) or (layer0_outputs(2093));
    layer1_outputs(3075) <= not(layer0_outputs(4311));
    layer1_outputs(3076) <= (layer0_outputs(2503)) and not (layer0_outputs(4911));
    layer1_outputs(3077) <= not(layer0_outputs(525)) or (layer0_outputs(3809));
    layer1_outputs(3078) <= not(layer0_outputs(862));
    layer1_outputs(3079) <= not(layer0_outputs(4394));
    layer1_outputs(3080) <= (layer0_outputs(107)) xor (layer0_outputs(3057));
    layer1_outputs(3081) <= not(layer0_outputs(3449)) or (layer0_outputs(967));
    layer1_outputs(3082) <= not(layer0_outputs(4222)) or (layer0_outputs(4569));
    layer1_outputs(3083) <= (layer0_outputs(4813)) and not (layer0_outputs(579));
    layer1_outputs(3084) <= (layer0_outputs(4961)) and (layer0_outputs(814));
    layer1_outputs(3085) <= '1';
    layer1_outputs(3086) <= '1';
    layer1_outputs(3087) <= not((layer0_outputs(3253)) or (layer0_outputs(509)));
    layer1_outputs(3088) <= not((layer0_outputs(4952)) or (layer0_outputs(414)));
    layer1_outputs(3089) <= layer0_outputs(2808);
    layer1_outputs(3090) <= (layer0_outputs(1885)) and not (layer0_outputs(5103));
    layer1_outputs(3091) <= '0';
    layer1_outputs(3092) <= not((layer0_outputs(1180)) or (layer0_outputs(4794)));
    layer1_outputs(3093) <= (layer0_outputs(282)) and not (layer0_outputs(4110));
    layer1_outputs(3094) <= not(layer0_outputs(3662)) or (layer0_outputs(4762));
    layer1_outputs(3095) <= not(layer0_outputs(4407));
    layer1_outputs(3096) <= not(layer0_outputs(539));
    layer1_outputs(3097) <= (layer0_outputs(1290)) or (layer0_outputs(2692));
    layer1_outputs(3098) <= not((layer0_outputs(430)) and (layer0_outputs(1876)));
    layer1_outputs(3099) <= not(layer0_outputs(4119)) or (layer0_outputs(3478));
    layer1_outputs(3100) <= (layer0_outputs(3001)) and not (layer0_outputs(3116));
    layer1_outputs(3101) <= (layer0_outputs(4861)) and (layer0_outputs(2944));
    layer1_outputs(3102) <= (layer0_outputs(4749)) and (layer0_outputs(956));
    layer1_outputs(3103) <= layer0_outputs(2545);
    layer1_outputs(3104) <= not(layer0_outputs(2343)) or (layer0_outputs(2166));
    layer1_outputs(3105) <= (layer0_outputs(3426)) and not (layer0_outputs(984));
    layer1_outputs(3106) <= not(layer0_outputs(1287));
    layer1_outputs(3107) <= '0';
    layer1_outputs(3108) <= (layer0_outputs(2924)) and (layer0_outputs(933));
    layer1_outputs(3109) <= (layer0_outputs(2011)) or (layer0_outputs(924));
    layer1_outputs(3110) <= (layer0_outputs(4915)) and not (layer0_outputs(193));
    layer1_outputs(3111) <= (layer0_outputs(4961)) or (layer0_outputs(2562));
    layer1_outputs(3112) <= '1';
    layer1_outputs(3113) <= not(layer0_outputs(1075)) or (layer0_outputs(2366));
    layer1_outputs(3114) <= not((layer0_outputs(4028)) and (layer0_outputs(2477)));
    layer1_outputs(3115) <= layer0_outputs(2725);
    layer1_outputs(3116) <= not((layer0_outputs(2794)) or (layer0_outputs(2839)));
    layer1_outputs(3117) <= (layer0_outputs(2689)) or (layer0_outputs(2519));
    layer1_outputs(3118) <= '1';
    layer1_outputs(3119) <= layer0_outputs(3630);
    layer1_outputs(3120) <= not(layer0_outputs(2735)) or (layer0_outputs(253));
    layer1_outputs(3121) <= (layer0_outputs(1217)) and (layer0_outputs(4719));
    layer1_outputs(3122) <= (layer0_outputs(858)) and not (layer0_outputs(4613));
    layer1_outputs(3123) <= (layer0_outputs(1856)) xor (layer0_outputs(3994));
    layer1_outputs(3124) <= not((layer0_outputs(4441)) or (layer0_outputs(4616)));
    layer1_outputs(3125) <= not((layer0_outputs(4194)) and (layer0_outputs(3977)));
    layer1_outputs(3126) <= not(layer0_outputs(4625)) or (layer0_outputs(196));
    layer1_outputs(3127) <= (layer0_outputs(1091)) or (layer0_outputs(178));
    layer1_outputs(3128) <= (layer0_outputs(2873)) and not (layer0_outputs(2771));
    layer1_outputs(3129) <= not(layer0_outputs(2815));
    layer1_outputs(3130) <= '0';
    layer1_outputs(3131) <= (layer0_outputs(3718)) or (layer0_outputs(497));
    layer1_outputs(3132) <= layer0_outputs(3665);
    layer1_outputs(3133) <= layer0_outputs(498);
    layer1_outputs(3134) <= '1';
    layer1_outputs(3135) <= (layer0_outputs(2599)) or (layer0_outputs(2632));
    layer1_outputs(3136) <= (layer0_outputs(4338)) and not (layer0_outputs(4398));
    layer1_outputs(3137) <= layer0_outputs(2586);
    layer1_outputs(3138) <= (layer0_outputs(3298)) and not (layer0_outputs(576));
    layer1_outputs(3139) <= not(layer0_outputs(1391));
    layer1_outputs(3140) <= not((layer0_outputs(4197)) and (layer0_outputs(433)));
    layer1_outputs(3141) <= not((layer0_outputs(2340)) or (layer0_outputs(3138)));
    layer1_outputs(3142) <= layer0_outputs(1690);
    layer1_outputs(3143) <= not(layer0_outputs(2892)) or (layer0_outputs(1122));
    layer1_outputs(3144) <= not(layer0_outputs(2591)) or (layer0_outputs(1022));
    layer1_outputs(3145) <= (layer0_outputs(1597)) or (layer0_outputs(4264));
    layer1_outputs(3146) <= '1';
    layer1_outputs(3147) <= not(layer0_outputs(4093));
    layer1_outputs(3148) <= not(layer0_outputs(1581)) or (layer0_outputs(592));
    layer1_outputs(3149) <= not(layer0_outputs(3885));
    layer1_outputs(3150) <= '1';
    layer1_outputs(3151) <= not((layer0_outputs(1699)) xor (layer0_outputs(3026)));
    layer1_outputs(3152) <= '0';
    layer1_outputs(3153) <= '1';
    layer1_outputs(3154) <= '1';
    layer1_outputs(3155) <= layer0_outputs(532);
    layer1_outputs(3156) <= (layer0_outputs(2091)) or (layer0_outputs(2875));
    layer1_outputs(3157) <= '1';
    layer1_outputs(3158) <= not(layer0_outputs(1360));
    layer1_outputs(3159) <= (layer0_outputs(2966)) and not (layer0_outputs(1601));
    layer1_outputs(3160) <= not(layer0_outputs(668));
    layer1_outputs(3161) <= (layer0_outputs(960)) and not (layer0_outputs(4664));
    layer1_outputs(3162) <= not((layer0_outputs(692)) or (layer0_outputs(1350)));
    layer1_outputs(3163) <= not((layer0_outputs(1062)) or (layer0_outputs(863)));
    layer1_outputs(3164) <= not(layer0_outputs(4183)) or (layer0_outputs(5080));
    layer1_outputs(3165) <= '0';
    layer1_outputs(3166) <= '0';
    layer1_outputs(3167) <= not(layer0_outputs(4310));
    layer1_outputs(3168) <= layer0_outputs(3386);
    layer1_outputs(3169) <= not(layer0_outputs(2084));
    layer1_outputs(3170) <= (layer0_outputs(3320)) and not (layer0_outputs(844));
    layer1_outputs(3171) <= layer0_outputs(1264);
    layer1_outputs(3172) <= not(layer0_outputs(1842));
    layer1_outputs(3173) <= '0';
    layer1_outputs(3174) <= '0';
    layer1_outputs(3175) <= (layer0_outputs(2372)) and not (layer0_outputs(2847));
    layer1_outputs(3176) <= layer0_outputs(4126);
    layer1_outputs(3177) <= layer0_outputs(3410);
    layer1_outputs(3178) <= layer0_outputs(3841);
    layer1_outputs(3179) <= (layer0_outputs(3411)) and not (layer0_outputs(40));
    layer1_outputs(3180) <= (layer0_outputs(1459)) and not (layer0_outputs(1327));
    layer1_outputs(3181) <= (layer0_outputs(1983)) and not (layer0_outputs(1315));
    layer1_outputs(3182) <= not(layer0_outputs(4726));
    layer1_outputs(3183) <= layer0_outputs(3176);
    layer1_outputs(3184) <= '1';
    layer1_outputs(3185) <= not(layer0_outputs(2493)) or (layer0_outputs(694));
    layer1_outputs(3186) <= (layer0_outputs(4741)) and not (layer0_outputs(240));
    layer1_outputs(3187) <= not(layer0_outputs(2722));
    layer1_outputs(3188) <= layer0_outputs(906);
    layer1_outputs(3189) <= not(layer0_outputs(230)) or (layer0_outputs(3252));
    layer1_outputs(3190) <= not((layer0_outputs(4562)) or (layer0_outputs(1866)));
    layer1_outputs(3191) <= not(layer0_outputs(2015));
    layer1_outputs(3192) <= not(layer0_outputs(2324));
    layer1_outputs(3193) <= (layer0_outputs(3409)) or (layer0_outputs(965));
    layer1_outputs(3194) <= '1';
    layer1_outputs(3195) <= (layer0_outputs(1734)) or (layer0_outputs(290));
    layer1_outputs(3196) <= (layer0_outputs(329)) and not (layer0_outputs(2259));
    layer1_outputs(3197) <= not((layer0_outputs(148)) or (layer0_outputs(1211)));
    layer1_outputs(3198) <= (layer0_outputs(40)) or (layer0_outputs(827));
    layer1_outputs(3199) <= '1';
    layer1_outputs(3200) <= not(layer0_outputs(3595));
    layer1_outputs(3201) <= '0';
    layer1_outputs(3202) <= layer0_outputs(1332);
    layer1_outputs(3203) <= not((layer0_outputs(2704)) xor (layer0_outputs(4934)));
    layer1_outputs(3204) <= '1';
    layer1_outputs(3205) <= not(layer0_outputs(788));
    layer1_outputs(3206) <= layer0_outputs(2519);
    layer1_outputs(3207) <= (layer0_outputs(1372)) and (layer0_outputs(1313));
    layer1_outputs(3208) <= not(layer0_outputs(3625));
    layer1_outputs(3209) <= not(layer0_outputs(4219)) or (layer0_outputs(1716));
    layer1_outputs(3210) <= not((layer0_outputs(2230)) or (layer0_outputs(3991)));
    layer1_outputs(3211) <= '1';
    layer1_outputs(3212) <= '0';
    layer1_outputs(3213) <= (layer0_outputs(952)) and not (layer0_outputs(721));
    layer1_outputs(3214) <= (layer0_outputs(4951)) or (layer0_outputs(2951));
    layer1_outputs(3215) <= (layer0_outputs(4870)) or (layer0_outputs(4098));
    layer1_outputs(3216) <= not(layer0_outputs(2705)) or (layer0_outputs(3938));
    layer1_outputs(3217) <= layer0_outputs(3987);
    layer1_outputs(3218) <= not(layer0_outputs(610)) or (layer0_outputs(2474));
    layer1_outputs(3219) <= layer0_outputs(651);
    layer1_outputs(3220) <= '1';
    layer1_outputs(3221) <= not((layer0_outputs(4936)) and (layer0_outputs(4459)));
    layer1_outputs(3222) <= not(layer0_outputs(4609));
    layer1_outputs(3223) <= layer0_outputs(3201);
    layer1_outputs(3224) <= (layer0_outputs(2668)) or (layer0_outputs(1212));
    layer1_outputs(3225) <= not(layer0_outputs(1049));
    layer1_outputs(3226) <= '0';
    layer1_outputs(3227) <= '1';
    layer1_outputs(3228) <= layer0_outputs(1020);
    layer1_outputs(3229) <= (layer0_outputs(1998)) and (layer0_outputs(1888));
    layer1_outputs(3230) <= not(layer0_outputs(803));
    layer1_outputs(3231) <= not(layer0_outputs(1416)) or (layer0_outputs(571));
    layer1_outputs(3232) <= '1';
    layer1_outputs(3233) <= not(layer0_outputs(2109)) or (layer0_outputs(2269));
    layer1_outputs(3234) <= (layer0_outputs(1886)) or (layer0_outputs(1427));
    layer1_outputs(3235) <= (layer0_outputs(2377)) or (layer0_outputs(1675));
    layer1_outputs(3236) <= '0';
    layer1_outputs(3237) <= layer0_outputs(2690);
    layer1_outputs(3238) <= (layer0_outputs(1736)) or (layer0_outputs(4127));
    layer1_outputs(3239) <= not((layer0_outputs(105)) and (layer0_outputs(2352)));
    layer1_outputs(3240) <= layer0_outputs(3426);
    layer1_outputs(3241) <= (layer0_outputs(3915)) or (layer0_outputs(4005));
    layer1_outputs(3242) <= (layer0_outputs(4761)) or (layer0_outputs(3262));
    layer1_outputs(3243) <= '0';
    layer1_outputs(3244) <= not((layer0_outputs(1241)) and (layer0_outputs(4347)));
    layer1_outputs(3245) <= '0';
    layer1_outputs(3246) <= (layer0_outputs(2565)) or (layer0_outputs(996));
    layer1_outputs(3247) <= not(layer0_outputs(2269));
    layer1_outputs(3248) <= not(layer0_outputs(4575));
    layer1_outputs(3249) <= layer0_outputs(1772);
    layer1_outputs(3250) <= not((layer0_outputs(4368)) xor (layer0_outputs(923)));
    layer1_outputs(3251) <= (layer0_outputs(4424)) and not (layer0_outputs(2905));
    layer1_outputs(3252) <= not(layer0_outputs(1813)) or (layer0_outputs(4807));
    layer1_outputs(3253) <= (layer0_outputs(512)) and not (layer0_outputs(816));
    layer1_outputs(3254) <= (layer0_outputs(3509)) or (layer0_outputs(3873));
    layer1_outputs(3255) <= not(layer0_outputs(765));
    layer1_outputs(3256) <= layer0_outputs(1064);
    layer1_outputs(3257) <= not(layer0_outputs(1673));
    layer1_outputs(3258) <= not(layer0_outputs(60));
    layer1_outputs(3259) <= '1';
    layer1_outputs(3260) <= not(layer0_outputs(4548)) or (layer0_outputs(3381));
    layer1_outputs(3261) <= layer0_outputs(2007);
    layer1_outputs(3262) <= not(layer0_outputs(1767)) or (layer0_outputs(4739));
    layer1_outputs(3263) <= layer0_outputs(4457);
    layer1_outputs(3264) <= not((layer0_outputs(983)) or (layer0_outputs(1800)));
    layer1_outputs(3265) <= '1';
    layer1_outputs(3266) <= layer0_outputs(3547);
    layer1_outputs(3267) <= not((layer0_outputs(4233)) and (layer0_outputs(4931)));
    layer1_outputs(3268) <= (layer0_outputs(5112)) and not (layer0_outputs(4331));
    layer1_outputs(3269) <= not((layer0_outputs(2887)) and (layer0_outputs(3923)));
    layer1_outputs(3270) <= not(layer0_outputs(588)) or (layer0_outputs(3778));
    layer1_outputs(3271) <= not((layer0_outputs(2430)) or (layer0_outputs(2388)));
    layer1_outputs(3272) <= not(layer0_outputs(1341));
    layer1_outputs(3273) <= (layer0_outputs(3431)) and (layer0_outputs(2541));
    layer1_outputs(3274) <= not(layer0_outputs(375));
    layer1_outputs(3275) <= (layer0_outputs(1990)) and not (layer0_outputs(458));
    layer1_outputs(3276) <= not((layer0_outputs(4832)) xor (layer0_outputs(2619)));
    layer1_outputs(3277) <= not(layer0_outputs(4735)) or (layer0_outputs(4589));
    layer1_outputs(3278) <= not(layer0_outputs(793));
    layer1_outputs(3279) <= not((layer0_outputs(4546)) or (layer0_outputs(3416)));
    layer1_outputs(3280) <= layer0_outputs(1931);
    layer1_outputs(3281) <= (layer0_outputs(235)) and not (layer0_outputs(457));
    layer1_outputs(3282) <= '1';
    layer1_outputs(3283) <= '0';
    layer1_outputs(3284) <= layer0_outputs(981);
    layer1_outputs(3285) <= not(layer0_outputs(207)) or (layer0_outputs(737));
    layer1_outputs(3286) <= not((layer0_outputs(3472)) or (layer0_outputs(2498)));
    layer1_outputs(3287) <= '0';
    layer1_outputs(3288) <= (layer0_outputs(1080)) and not (layer0_outputs(895));
    layer1_outputs(3289) <= layer0_outputs(982);
    layer1_outputs(3290) <= (layer0_outputs(1626)) xor (layer0_outputs(1462));
    layer1_outputs(3291) <= not(layer0_outputs(4519)) or (layer0_outputs(3456));
    layer1_outputs(3292) <= not(layer0_outputs(4540)) or (layer0_outputs(913));
    layer1_outputs(3293) <= (layer0_outputs(800)) and (layer0_outputs(1882));
    layer1_outputs(3294) <= not(layer0_outputs(3784)) or (layer0_outputs(4082));
    layer1_outputs(3295) <= (layer0_outputs(689)) and (layer0_outputs(2953));
    layer1_outputs(3296) <= '0';
    layer1_outputs(3297) <= not(layer0_outputs(4737)) or (layer0_outputs(2424));
    layer1_outputs(3298) <= (layer0_outputs(77)) and (layer0_outputs(1251));
    layer1_outputs(3299) <= '1';
    layer1_outputs(3300) <= not(layer0_outputs(2010)) or (layer0_outputs(4107));
    layer1_outputs(3301) <= not(layer0_outputs(2113));
    layer1_outputs(3302) <= layer0_outputs(4706);
    layer1_outputs(3303) <= '0';
    layer1_outputs(3304) <= layer0_outputs(595);
    layer1_outputs(3305) <= (layer0_outputs(2355)) and not (layer0_outputs(1479));
    layer1_outputs(3306) <= (layer0_outputs(3384)) and (layer0_outputs(4755));
    layer1_outputs(3307) <= not(layer0_outputs(2972));
    layer1_outputs(3308) <= (layer0_outputs(3952)) and (layer0_outputs(156));
    layer1_outputs(3309) <= not(layer0_outputs(2746)) or (layer0_outputs(5064));
    layer1_outputs(3310) <= layer0_outputs(5055);
    layer1_outputs(3311) <= not((layer0_outputs(774)) or (layer0_outputs(1454)));
    layer1_outputs(3312) <= not((layer0_outputs(616)) or (layer0_outputs(2745)));
    layer1_outputs(3313) <= not((layer0_outputs(674)) or (layer0_outputs(5040)));
    layer1_outputs(3314) <= not(layer0_outputs(1667));
    layer1_outputs(3315) <= not(layer0_outputs(556));
    layer1_outputs(3316) <= not(layer0_outputs(3631)) or (layer0_outputs(2346));
    layer1_outputs(3317) <= layer0_outputs(3299);
    layer1_outputs(3318) <= (layer0_outputs(2970)) and (layer0_outputs(5026));
    layer1_outputs(3319) <= '0';
    layer1_outputs(3320) <= '0';
    layer1_outputs(3321) <= '1';
    layer1_outputs(3322) <= '0';
    layer1_outputs(3323) <= (layer0_outputs(3436)) and (layer0_outputs(56));
    layer1_outputs(3324) <= not(layer0_outputs(1498)) or (layer0_outputs(3062));
    layer1_outputs(3325) <= (layer0_outputs(2796)) or (layer0_outputs(208));
    layer1_outputs(3326) <= (layer0_outputs(3743)) or (layer0_outputs(3175));
    layer1_outputs(3327) <= '1';
    layer1_outputs(3328) <= (layer0_outputs(3134)) and not (layer0_outputs(389));
    layer1_outputs(3329) <= '0';
    layer1_outputs(3330) <= (layer0_outputs(5002)) or (layer0_outputs(1395));
    layer1_outputs(3331) <= layer0_outputs(154);
    layer1_outputs(3332) <= (layer0_outputs(1544)) and (layer0_outputs(1221));
    layer1_outputs(3333) <= layer0_outputs(244);
    layer1_outputs(3334) <= layer0_outputs(3755);
    layer1_outputs(3335) <= '0';
    layer1_outputs(3336) <= (layer0_outputs(4530)) and not (layer0_outputs(3041));
    layer1_outputs(3337) <= (layer0_outputs(1293)) and not (layer0_outputs(1928));
    layer1_outputs(3338) <= not(layer0_outputs(4547)) or (layer0_outputs(202));
    layer1_outputs(3339) <= '0';
    layer1_outputs(3340) <= not((layer0_outputs(5097)) or (layer0_outputs(4352)));
    layer1_outputs(3341) <= not((layer0_outputs(3489)) or (layer0_outputs(3271)));
    layer1_outputs(3342) <= not(layer0_outputs(1876)) or (layer0_outputs(1984));
    layer1_outputs(3343) <= not(layer0_outputs(3184));
    layer1_outputs(3344) <= not(layer0_outputs(530));
    layer1_outputs(3345) <= layer0_outputs(831);
    layer1_outputs(3346) <= '0';
    layer1_outputs(3347) <= not(layer0_outputs(572));
    layer1_outputs(3348) <= '0';
    layer1_outputs(3349) <= (layer0_outputs(3857)) and not (layer0_outputs(1228));
    layer1_outputs(3350) <= '0';
    layer1_outputs(3351) <= (layer0_outputs(3274)) and (layer0_outputs(2491));
    layer1_outputs(3352) <= not((layer0_outputs(4371)) and (layer0_outputs(1887)));
    layer1_outputs(3353) <= layer0_outputs(3716);
    layer1_outputs(3354) <= '1';
    layer1_outputs(3355) <= not((layer0_outputs(3384)) or (layer0_outputs(3315)));
    layer1_outputs(3356) <= not(layer0_outputs(4161)) or (layer0_outputs(81));
    layer1_outputs(3357) <= not(layer0_outputs(2211));
    layer1_outputs(3358) <= layer0_outputs(4052);
    layer1_outputs(3359) <= not(layer0_outputs(3629));
    layer1_outputs(3360) <= layer0_outputs(1612);
    layer1_outputs(3361) <= layer0_outputs(3472);
    layer1_outputs(3362) <= (layer0_outputs(3339)) and not (layer0_outputs(477));
    layer1_outputs(3363) <= not(layer0_outputs(2074)) or (layer0_outputs(4028));
    layer1_outputs(3364) <= '1';
    layer1_outputs(3365) <= not((layer0_outputs(1247)) or (layer0_outputs(1594)));
    layer1_outputs(3366) <= (layer0_outputs(4557)) and not (layer0_outputs(3893));
    layer1_outputs(3367) <= not((layer0_outputs(758)) or (layer0_outputs(438)));
    layer1_outputs(3368) <= '0';
    layer1_outputs(3369) <= layer0_outputs(1527);
    layer1_outputs(3370) <= not((layer0_outputs(3262)) and (layer0_outputs(3180)));
    layer1_outputs(3371) <= not(layer0_outputs(2117)) or (layer0_outputs(4267));
    layer1_outputs(3372) <= layer0_outputs(199);
    layer1_outputs(3373) <= not(layer0_outputs(2473)) or (layer0_outputs(1788));
    layer1_outputs(3374) <= not(layer0_outputs(2751)) or (layer0_outputs(588));
    layer1_outputs(3375) <= layer0_outputs(2030);
    layer1_outputs(3376) <= not(layer0_outputs(4846));
    layer1_outputs(3377) <= (layer0_outputs(4702)) xor (layer0_outputs(1125));
    layer1_outputs(3378) <= not(layer0_outputs(3537));
    layer1_outputs(3379) <= not(layer0_outputs(3269));
    layer1_outputs(3380) <= not(layer0_outputs(3676)) or (layer0_outputs(4131));
    layer1_outputs(3381) <= layer0_outputs(1756);
    layer1_outputs(3382) <= not((layer0_outputs(2535)) or (layer0_outputs(4535)));
    layer1_outputs(3383) <= '1';
    layer1_outputs(3384) <= layer0_outputs(2011);
    layer1_outputs(3385) <= not(layer0_outputs(139));
    layer1_outputs(3386) <= layer0_outputs(3499);
    layer1_outputs(3387) <= '0';
    layer1_outputs(3388) <= layer0_outputs(4062);
    layer1_outputs(3389) <= not((layer0_outputs(1053)) or (layer0_outputs(549)));
    layer1_outputs(3390) <= (layer0_outputs(2422)) and (layer0_outputs(4763));
    layer1_outputs(3391) <= layer0_outputs(4000);
    layer1_outputs(3392) <= '0';
    layer1_outputs(3393) <= '1';
    layer1_outputs(3394) <= (layer0_outputs(298)) and (layer0_outputs(4356));
    layer1_outputs(3395) <= not((layer0_outputs(1681)) or (layer0_outputs(3661)));
    layer1_outputs(3396) <= not(layer0_outputs(4228));
    layer1_outputs(3397) <= (layer0_outputs(4799)) and (layer0_outputs(2411));
    layer1_outputs(3398) <= '1';
    layer1_outputs(3399) <= '0';
    layer1_outputs(3400) <= layer0_outputs(4853);
    layer1_outputs(3401) <= (layer0_outputs(3093)) and (layer0_outputs(5058));
    layer1_outputs(3402) <= not((layer0_outputs(631)) or (layer0_outputs(3518)));
    layer1_outputs(3403) <= '0';
    layer1_outputs(3404) <= not(layer0_outputs(3736)) or (layer0_outputs(43));
    layer1_outputs(3405) <= not(layer0_outputs(5014)) or (layer0_outputs(1817));
    layer1_outputs(3406) <= (layer0_outputs(3952)) xor (layer0_outputs(3613));
    layer1_outputs(3407) <= layer0_outputs(2925);
    layer1_outputs(3408) <= (layer0_outputs(5034)) and not (layer0_outputs(1936));
    layer1_outputs(3409) <= '0';
    layer1_outputs(3410) <= not((layer0_outputs(3406)) and (layer0_outputs(248)));
    layer1_outputs(3411) <= layer0_outputs(2922);
    layer1_outputs(3412) <= (layer0_outputs(3990)) and (layer0_outputs(305));
    layer1_outputs(3413) <= layer0_outputs(3951);
    layer1_outputs(3414) <= layer0_outputs(630);
    layer1_outputs(3415) <= not(layer0_outputs(2399)) or (layer0_outputs(2528));
    layer1_outputs(3416) <= '0';
    layer1_outputs(3417) <= not(layer0_outputs(1575)) or (layer0_outputs(2958));
    layer1_outputs(3418) <= (layer0_outputs(3731)) and (layer0_outputs(776));
    layer1_outputs(3419) <= not((layer0_outputs(1229)) and (layer0_outputs(1901)));
    layer1_outputs(3420) <= not(layer0_outputs(2073)) or (layer0_outputs(231));
    layer1_outputs(3421) <= layer0_outputs(711);
    layer1_outputs(3422) <= not(layer0_outputs(3238)) or (layer0_outputs(78));
    layer1_outputs(3423) <= layer0_outputs(1238);
    layer1_outputs(3424) <= not((layer0_outputs(3194)) and (layer0_outputs(2402)));
    layer1_outputs(3425) <= (layer0_outputs(2273)) and (layer0_outputs(4104));
    layer1_outputs(3426) <= layer0_outputs(2937);
    layer1_outputs(3427) <= not((layer0_outputs(3931)) xor (layer0_outputs(4001)));
    layer1_outputs(3428) <= '0';
    layer1_outputs(3429) <= not(layer0_outputs(3487));
    layer1_outputs(3430) <= (layer0_outputs(4397)) and not (layer0_outputs(1795));
    layer1_outputs(3431) <= (layer0_outputs(3390)) and (layer0_outputs(1208));
    layer1_outputs(3432) <= layer0_outputs(3126);
    layer1_outputs(3433) <= (layer0_outputs(2036)) and not (layer0_outputs(1910));
    layer1_outputs(3434) <= '1';
    layer1_outputs(3435) <= not(layer0_outputs(2780));
    layer1_outputs(3436) <= (layer0_outputs(666)) or (layer0_outputs(4810));
    layer1_outputs(3437) <= '0';
    layer1_outputs(3438) <= (layer0_outputs(123)) and not (layer0_outputs(2178));
    layer1_outputs(3439) <= (layer0_outputs(5076)) or (layer0_outputs(3667));
    layer1_outputs(3440) <= '1';
    layer1_outputs(3441) <= layer0_outputs(3098);
    layer1_outputs(3442) <= not(layer0_outputs(368));
    layer1_outputs(3443) <= not(layer0_outputs(1696));
    layer1_outputs(3444) <= not(layer0_outputs(2966)) or (layer0_outputs(3876));
    layer1_outputs(3445) <= '0';
    layer1_outputs(3446) <= (layer0_outputs(2531)) and (layer0_outputs(3847));
    layer1_outputs(3447) <= not(layer0_outputs(484)) or (layer0_outputs(3228));
    layer1_outputs(3448) <= not((layer0_outputs(2708)) or (layer0_outputs(2809)));
    layer1_outputs(3449) <= '1';
    layer1_outputs(3450) <= (layer0_outputs(3741)) and not (layer0_outputs(30));
    layer1_outputs(3451) <= layer0_outputs(1146);
    layer1_outputs(3452) <= '0';
    layer1_outputs(3453) <= not(layer0_outputs(3485));
    layer1_outputs(3454) <= not((layer0_outputs(1894)) or (layer0_outputs(615)));
    layer1_outputs(3455) <= layer0_outputs(1530);
    layer1_outputs(3456) <= layer0_outputs(2150);
    layer1_outputs(3457) <= (layer0_outputs(351)) and not (layer0_outputs(4722));
    layer1_outputs(3458) <= (layer0_outputs(4164)) and not (layer0_outputs(4024));
    layer1_outputs(3459) <= not(layer0_outputs(2375));
    layer1_outputs(3460) <= layer0_outputs(661);
    layer1_outputs(3461) <= not((layer0_outputs(1641)) and (layer0_outputs(4141)));
    layer1_outputs(3462) <= '0';
    layer1_outputs(3463) <= layer0_outputs(2036);
    layer1_outputs(3464) <= not(layer0_outputs(472)) or (layer0_outputs(343));
    layer1_outputs(3465) <= (layer0_outputs(2179)) and (layer0_outputs(1299));
    layer1_outputs(3466) <= layer0_outputs(1838);
    layer1_outputs(3467) <= not((layer0_outputs(1950)) and (layer0_outputs(2993)));
    layer1_outputs(3468) <= layer0_outputs(820);
    layer1_outputs(3469) <= (layer0_outputs(1528)) and not (layer0_outputs(4750));
    layer1_outputs(3470) <= (layer0_outputs(1145)) and not (layer0_outputs(1266));
    layer1_outputs(3471) <= not((layer0_outputs(2556)) and (layer0_outputs(4556)));
    layer1_outputs(3472) <= '1';
    layer1_outputs(3473) <= '0';
    layer1_outputs(3474) <= not(layer0_outputs(1392)) or (layer0_outputs(3218));
    layer1_outputs(3475) <= not(layer0_outputs(1443));
    layer1_outputs(3476) <= '0';
    layer1_outputs(3477) <= layer0_outputs(1533);
    layer1_outputs(3478) <= layer0_outputs(1249);
    layer1_outputs(3479) <= not(layer0_outputs(1284));
    layer1_outputs(3480) <= not(layer0_outputs(226)) or (layer0_outputs(2477));
    layer1_outputs(3481) <= not((layer0_outputs(4299)) or (layer0_outputs(3897)));
    layer1_outputs(3482) <= '0';
    layer1_outputs(3483) <= not((layer0_outputs(643)) and (layer0_outputs(4518)));
    layer1_outputs(3484) <= not(layer0_outputs(1367));
    layer1_outputs(3485) <= '0';
    layer1_outputs(3486) <= not(layer0_outputs(4148));
    layer1_outputs(3487) <= '0';
    layer1_outputs(3488) <= (layer0_outputs(3880)) and (layer0_outputs(3177));
    layer1_outputs(3489) <= layer0_outputs(2805);
    layer1_outputs(3490) <= '0';
    layer1_outputs(3491) <= (layer0_outputs(4074)) or (layer0_outputs(3752));
    layer1_outputs(3492) <= (layer0_outputs(4202)) and not (layer0_outputs(3716));
    layer1_outputs(3493) <= (layer0_outputs(3506)) and (layer0_outputs(3505));
    layer1_outputs(3494) <= '1';
    layer1_outputs(3495) <= (layer0_outputs(1085)) xor (layer0_outputs(3746));
    layer1_outputs(3496) <= '1';
    layer1_outputs(3497) <= not(layer0_outputs(4372));
    layer1_outputs(3498) <= (layer0_outputs(4095)) and not (layer0_outputs(2550));
    layer1_outputs(3499) <= not(layer0_outputs(1360));
    layer1_outputs(3500) <= not(layer0_outputs(1402)) or (layer0_outputs(1976));
    layer1_outputs(3501) <= (layer0_outputs(506)) and not (layer0_outputs(1078));
    layer1_outputs(3502) <= not((layer0_outputs(2826)) or (layer0_outputs(1281)));
    layer1_outputs(3503) <= not(layer0_outputs(3414));
    layer1_outputs(3504) <= (layer0_outputs(2586)) and not (layer0_outputs(1289));
    layer1_outputs(3505) <= (layer0_outputs(2514)) and (layer0_outputs(5012));
    layer1_outputs(3506) <= not(layer0_outputs(2954)) or (layer0_outputs(2640));
    layer1_outputs(3507) <= (layer0_outputs(423)) and (layer0_outputs(470));
    layer1_outputs(3508) <= '1';
    layer1_outputs(3509) <= not(layer0_outputs(3307));
    layer1_outputs(3510) <= not((layer0_outputs(1044)) xor (layer0_outputs(4015)));
    layer1_outputs(3511) <= not(layer0_outputs(929));
    layer1_outputs(3512) <= (layer0_outputs(2593)) and not (layer0_outputs(1484));
    layer1_outputs(3513) <= not(layer0_outputs(3352)) or (layer0_outputs(21));
    layer1_outputs(3514) <= (layer0_outputs(2327)) and not (layer0_outputs(2272));
    layer1_outputs(3515) <= not(layer0_outputs(795)) or (layer0_outputs(3704));
    layer1_outputs(3516) <= not((layer0_outputs(4375)) or (layer0_outputs(49)));
    layer1_outputs(3517) <= (layer0_outputs(2627)) and (layer0_outputs(1321));
    layer1_outputs(3518) <= not(layer0_outputs(396)) or (layer0_outputs(1863));
    layer1_outputs(3519) <= not((layer0_outputs(5101)) and (layer0_outputs(2680)));
    layer1_outputs(3520) <= '0';
    layer1_outputs(3521) <= not(layer0_outputs(4748)) or (layer0_outputs(3471));
    layer1_outputs(3522) <= '0';
    layer1_outputs(3523) <= '0';
    layer1_outputs(3524) <= layer0_outputs(4837);
    layer1_outputs(3525) <= not(layer0_outputs(2052)) or (layer0_outputs(3814));
    layer1_outputs(3526) <= layer0_outputs(1844);
    layer1_outputs(3527) <= layer0_outputs(3130);
    layer1_outputs(3528) <= (layer0_outputs(3256)) and not (layer0_outputs(1305));
    layer1_outputs(3529) <= '0';
    layer1_outputs(3530) <= not((layer0_outputs(2845)) or (layer0_outputs(4114)));
    layer1_outputs(3531) <= layer0_outputs(1168);
    layer1_outputs(3532) <= (layer0_outputs(2908)) and not (layer0_outputs(3988));
    layer1_outputs(3533) <= '0';
    layer1_outputs(3534) <= layer0_outputs(1880);
    layer1_outputs(3535) <= not(layer0_outputs(1294));
    layer1_outputs(3536) <= layer0_outputs(75);
    layer1_outputs(3537) <= not(layer0_outputs(2154));
    layer1_outputs(3538) <= '0';
    layer1_outputs(3539) <= not(layer0_outputs(2881));
    layer1_outputs(3540) <= layer0_outputs(203);
    layer1_outputs(3541) <= '1';
    layer1_outputs(3542) <= not(layer0_outputs(3159));
    layer1_outputs(3543) <= not(layer0_outputs(2431)) or (layer0_outputs(3095));
    layer1_outputs(3544) <= not((layer0_outputs(3398)) or (layer0_outputs(4069)));
    layer1_outputs(3545) <= '1';
    layer1_outputs(3546) <= not((layer0_outputs(1987)) xor (layer0_outputs(1405)));
    layer1_outputs(3547) <= '0';
    layer1_outputs(3548) <= (layer0_outputs(281)) and not (layer0_outputs(3003));
    layer1_outputs(3549) <= '0';
    layer1_outputs(3550) <= not(layer0_outputs(904)) or (layer0_outputs(462));
    layer1_outputs(3551) <= (layer0_outputs(1861)) and not (layer0_outputs(4734));
    layer1_outputs(3552) <= (layer0_outputs(3372)) and (layer0_outputs(2363));
    layer1_outputs(3553) <= layer0_outputs(2134);
    layer1_outputs(3554) <= (layer0_outputs(322)) and (layer0_outputs(1618));
    layer1_outputs(3555) <= '0';
    layer1_outputs(3556) <= (layer0_outputs(5027)) and not (layer0_outputs(197));
    layer1_outputs(3557) <= '0';
    layer1_outputs(3558) <= not((layer0_outputs(3055)) xor (layer0_outputs(4365)));
    layer1_outputs(3559) <= (layer0_outputs(3998)) and not (layer0_outputs(1516));
    layer1_outputs(3560) <= '1';
    layer1_outputs(3561) <= '0';
    layer1_outputs(3562) <= (layer0_outputs(2605)) and not (layer0_outputs(2415));
    layer1_outputs(3563) <= layer0_outputs(1562);
    layer1_outputs(3564) <= not(layer0_outputs(4469));
    layer1_outputs(3565) <= not((layer0_outputs(1388)) or (layer0_outputs(4417)));
    layer1_outputs(3566) <= (layer0_outputs(3161)) and not (layer0_outputs(2459));
    layer1_outputs(3567) <= not((layer0_outputs(2727)) and (layer0_outputs(826)));
    layer1_outputs(3568) <= layer0_outputs(470);
    layer1_outputs(3569) <= not((layer0_outputs(3284)) and (layer0_outputs(244)));
    layer1_outputs(3570) <= (layer0_outputs(1648)) and not (layer0_outputs(3491));
    layer1_outputs(3571) <= layer0_outputs(45);
    layer1_outputs(3572) <= not(layer0_outputs(2552)) or (layer0_outputs(642));
    layer1_outputs(3573) <= not(layer0_outputs(4924));
    layer1_outputs(3574) <= not((layer0_outputs(3068)) and (layer0_outputs(4980)));
    layer1_outputs(3575) <= (layer0_outputs(3648)) and (layer0_outputs(419));
    layer1_outputs(3576) <= '0';
    layer1_outputs(3577) <= not((layer0_outputs(1965)) and (layer0_outputs(2032)));
    layer1_outputs(3578) <= '0';
    layer1_outputs(3579) <= not(layer0_outputs(2312));
    layer1_outputs(3580) <= '0';
    layer1_outputs(3581) <= not((layer0_outputs(2909)) or (layer0_outputs(28)));
    layer1_outputs(3582) <= not((layer0_outputs(2862)) and (layer0_outputs(4987)));
    layer1_outputs(3583) <= '0';
    layer1_outputs(3584) <= (layer0_outputs(1627)) and not (layer0_outputs(3853));
    layer1_outputs(3585) <= (layer0_outputs(1190)) xor (layer0_outputs(2577));
    layer1_outputs(3586) <= layer0_outputs(1364);
    layer1_outputs(3587) <= not(layer0_outputs(1733)) or (layer0_outputs(96));
    layer1_outputs(3588) <= '0';
    layer1_outputs(3589) <= not((layer0_outputs(3260)) and (layer0_outputs(612)));
    layer1_outputs(3590) <= not(layer0_outputs(2287));
    layer1_outputs(3591) <= '0';
    layer1_outputs(3592) <= not(layer0_outputs(4618));
    layer1_outputs(3593) <= layer0_outputs(982);
    layer1_outputs(3594) <= '1';
    layer1_outputs(3595) <= layer0_outputs(4574);
    layer1_outputs(3596) <= not(layer0_outputs(2875)) or (layer0_outputs(3117));
    layer1_outputs(3597) <= '0';
    layer1_outputs(3598) <= (layer0_outputs(4598)) and not (layer0_outputs(1205));
    layer1_outputs(3599) <= layer0_outputs(1733);
    layer1_outputs(3600) <= not((layer0_outputs(1301)) and (layer0_outputs(3861)));
    layer1_outputs(3601) <= (layer0_outputs(2126)) and not (layer0_outputs(2567));
    layer1_outputs(3602) <= (layer0_outputs(300)) and not (layer0_outputs(4859));
    layer1_outputs(3603) <= not(layer0_outputs(3197));
    layer1_outputs(3604) <= layer0_outputs(4982);
    layer1_outputs(3605) <= '0';
    layer1_outputs(3606) <= not(layer0_outputs(3202)) or (layer0_outputs(3907));
    layer1_outputs(3607) <= '0';
    layer1_outputs(3608) <= not(layer0_outputs(1620)) or (layer0_outputs(3719));
    layer1_outputs(3609) <= '0';
    layer1_outputs(3610) <= layer0_outputs(3342);
    layer1_outputs(3611) <= (layer0_outputs(3679)) or (layer0_outputs(4283));
    layer1_outputs(3612) <= (layer0_outputs(603)) or (layer0_outputs(3960));
    layer1_outputs(3613) <= (layer0_outputs(4999)) or (layer0_outputs(2785));
    layer1_outputs(3614) <= not((layer0_outputs(3624)) and (layer0_outputs(1260)));
    layer1_outputs(3615) <= '1';
    layer1_outputs(3616) <= (layer0_outputs(3145)) and (layer0_outputs(4733));
    layer1_outputs(3617) <= (layer0_outputs(1783)) or (layer0_outputs(1792));
    layer1_outputs(3618) <= '0';
    layer1_outputs(3619) <= not(layer0_outputs(2855)) or (layer0_outputs(3791));
    layer1_outputs(3620) <= layer0_outputs(1153);
    layer1_outputs(3621) <= not(layer0_outputs(1280)) or (layer0_outputs(1849));
    layer1_outputs(3622) <= not(layer0_outputs(5049)) or (layer0_outputs(4128));
    layer1_outputs(3623) <= '1';
    layer1_outputs(3624) <= '1';
    layer1_outputs(3625) <= not(layer0_outputs(2753)) or (layer0_outputs(4009));
    layer1_outputs(3626) <= layer0_outputs(3200);
    layer1_outputs(3627) <= layer0_outputs(337);
    layer1_outputs(3628) <= not(layer0_outputs(2729)) or (layer0_outputs(68));
    layer1_outputs(3629) <= not(layer0_outputs(2694)) or (layer0_outputs(367));
    layer1_outputs(3630) <= not(layer0_outputs(1580));
    layer1_outputs(3631) <= (layer0_outputs(167)) and not (layer0_outputs(3747));
    layer1_outputs(3632) <= layer0_outputs(1757);
    layer1_outputs(3633) <= not(layer0_outputs(291)) or (layer0_outputs(2055));
    layer1_outputs(3634) <= '1';
    layer1_outputs(3635) <= not(layer0_outputs(3608)) or (layer0_outputs(1217));
    layer1_outputs(3636) <= not((layer0_outputs(526)) or (layer0_outputs(272)));
    layer1_outputs(3637) <= (layer0_outputs(3486)) and (layer0_outputs(3825));
    layer1_outputs(3638) <= not(layer0_outputs(1908));
    layer1_outputs(3639) <= (layer0_outputs(4932)) or (layer0_outputs(922));
    layer1_outputs(3640) <= (layer0_outputs(4774)) and not (layer0_outputs(1962));
    layer1_outputs(3641) <= '1';
    layer1_outputs(3642) <= not(layer0_outputs(4195));
    layer1_outputs(3643) <= (layer0_outputs(4943)) and (layer0_outputs(1538));
    layer1_outputs(3644) <= layer0_outputs(3601);
    layer1_outputs(3645) <= '1';
    layer1_outputs(3646) <= not((layer0_outputs(313)) and (layer0_outputs(2756)));
    layer1_outputs(3647) <= not(layer0_outputs(699)) or (layer0_outputs(3279));
    layer1_outputs(3648) <= layer0_outputs(537);
    layer1_outputs(3649) <= not(layer0_outputs(4705));
    layer1_outputs(3650) <= layer0_outputs(4926);
    layer1_outputs(3651) <= not(layer0_outputs(4632));
    layer1_outputs(3652) <= layer0_outputs(1066);
    layer1_outputs(3653) <= not(layer0_outputs(4636)) or (layer0_outputs(1107));
    layer1_outputs(3654) <= not(layer0_outputs(3830));
    layer1_outputs(3655) <= '0';
    layer1_outputs(3656) <= (layer0_outputs(4526)) and not (layer0_outputs(4429));
    layer1_outputs(3657) <= not((layer0_outputs(869)) and (layer0_outputs(1010)));
    layer1_outputs(3658) <= '1';
    layer1_outputs(3659) <= not(layer0_outputs(4787)) or (layer0_outputs(3619));
    layer1_outputs(3660) <= (layer0_outputs(1592)) and not (layer0_outputs(4698));
    layer1_outputs(3661) <= not(layer0_outputs(3576));
    layer1_outputs(3662) <= '0';
    layer1_outputs(3663) <= not(layer0_outputs(1167)) or (layer0_outputs(3946));
    layer1_outputs(3664) <= not(layer0_outputs(1200)) or (layer0_outputs(2987));
    layer1_outputs(3665) <= (layer0_outputs(2682)) or (layer0_outputs(2731));
    layer1_outputs(3666) <= not(layer0_outputs(3919));
    layer1_outputs(3667) <= (layer0_outputs(438)) or (layer0_outputs(1352));
    layer1_outputs(3668) <= layer0_outputs(1017);
    layer1_outputs(3669) <= not(layer0_outputs(3065));
    layer1_outputs(3670) <= layer0_outputs(2629);
    layer1_outputs(3671) <= (layer0_outputs(3316)) and not (layer0_outputs(4694));
    layer1_outputs(3672) <= not((layer0_outputs(1540)) or (layer0_outputs(454)));
    layer1_outputs(3673) <= (layer0_outputs(3764)) and not (layer0_outputs(2092));
    layer1_outputs(3674) <= not(layer0_outputs(1333)) or (layer0_outputs(4292));
    layer1_outputs(3675) <= (layer0_outputs(4937)) and not (layer0_outputs(2555));
    layer1_outputs(3676) <= not((layer0_outputs(789)) and (layer0_outputs(3901)));
    layer1_outputs(3677) <= (layer0_outputs(1599)) and not (layer0_outputs(3764));
    layer1_outputs(3678) <= not((layer0_outputs(3234)) and (layer0_outputs(4232)));
    layer1_outputs(3679) <= '0';
    layer1_outputs(3680) <= not(layer0_outputs(2058));
    layer1_outputs(3681) <= (layer0_outputs(1327)) and (layer0_outputs(4657));
    layer1_outputs(3682) <= not((layer0_outputs(960)) or (layer0_outputs(3331)));
    layer1_outputs(3683) <= not((layer0_outputs(211)) or (layer0_outputs(4753)));
    layer1_outputs(3684) <= not((layer0_outputs(3104)) and (layer0_outputs(2962)));
    layer1_outputs(3685) <= not((layer0_outputs(82)) and (layer0_outputs(4825)));
    layer1_outputs(3686) <= '0';
    layer1_outputs(3687) <= not(layer0_outputs(4067)) or (layer0_outputs(3042));
    layer1_outputs(3688) <= not(layer0_outputs(3437)) or (layer0_outputs(3640));
    layer1_outputs(3689) <= not((layer0_outputs(1714)) and (layer0_outputs(4403)));
    layer1_outputs(3690) <= not(layer0_outputs(918));
    layer1_outputs(3691) <= layer0_outputs(3464);
    layer1_outputs(3692) <= layer0_outputs(3101);
    layer1_outputs(3693) <= not((layer0_outputs(2317)) or (layer0_outputs(2444)));
    layer1_outputs(3694) <= not((layer0_outputs(2434)) and (layer0_outputs(1685)));
    layer1_outputs(3695) <= (layer0_outputs(2823)) and not (layer0_outputs(2439));
    layer1_outputs(3696) <= (layer0_outputs(3332)) and (layer0_outputs(5068));
    layer1_outputs(3697) <= '1';
    layer1_outputs(3698) <= not((layer0_outputs(3696)) or (layer0_outputs(2774)));
    layer1_outputs(3699) <= not(layer0_outputs(4201)) or (layer0_outputs(3965));
    layer1_outputs(3700) <= '0';
    layer1_outputs(3701) <= (layer0_outputs(5032)) or (layer0_outputs(3951));
    layer1_outputs(3702) <= '1';
    layer1_outputs(3703) <= not(layer0_outputs(87));
    layer1_outputs(3704) <= (layer0_outputs(4604)) or (layer0_outputs(857));
    layer1_outputs(3705) <= '1';
    layer1_outputs(3706) <= layer0_outputs(4727);
    layer1_outputs(3707) <= not(layer0_outputs(179));
    layer1_outputs(3708) <= '0';
    layer1_outputs(3709) <= (layer0_outputs(1846)) and not (layer0_outputs(4090));
    layer1_outputs(3710) <= '1';
    layer1_outputs(3711) <= not((layer0_outputs(1890)) or (layer0_outputs(3956)));
    layer1_outputs(3712) <= (layer0_outputs(4189)) and not (layer0_outputs(4064));
    layer1_outputs(3713) <= not(layer0_outputs(4073)) or (layer0_outputs(2028));
    layer1_outputs(3714) <= not((layer0_outputs(1521)) and (layer0_outputs(4901)));
    layer1_outputs(3715) <= (layer0_outputs(4043)) and not (layer0_outputs(3135));
    layer1_outputs(3716) <= not(layer0_outputs(2693));
    layer1_outputs(3717) <= not(layer0_outputs(2282));
    layer1_outputs(3718) <= '0';
    layer1_outputs(3719) <= '1';
    layer1_outputs(3720) <= layer0_outputs(4539);
    layer1_outputs(3721) <= '1';
    layer1_outputs(3722) <= layer0_outputs(2136);
    layer1_outputs(3723) <= '1';
    layer1_outputs(3724) <= not(layer0_outputs(1437));
    layer1_outputs(3725) <= not((layer0_outputs(2872)) and (layer0_outputs(1785)));
    layer1_outputs(3726) <= '0';
    layer1_outputs(3727) <= not(layer0_outputs(2719));
    layer1_outputs(3728) <= not(layer0_outputs(1556));
    layer1_outputs(3729) <= not(layer0_outputs(3534));
    layer1_outputs(3730) <= not(layer0_outputs(1041)) or (layer0_outputs(2832));
    layer1_outputs(3731) <= '0';
    layer1_outputs(3732) <= not((layer0_outputs(4845)) and (layer0_outputs(628)));
    layer1_outputs(3733) <= (layer0_outputs(3583)) and not (layer0_outputs(1989));
    layer1_outputs(3734) <= not((layer0_outputs(1676)) or (layer0_outputs(1219)));
    layer1_outputs(3735) <= (layer0_outputs(1209)) xor (layer0_outputs(4520));
    layer1_outputs(3736) <= layer0_outputs(1274);
    layer1_outputs(3737) <= not(layer0_outputs(2095)) or (layer0_outputs(1900));
    layer1_outputs(3738) <= not(layer0_outputs(3672)) or (layer0_outputs(1106));
    layer1_outputs(3739) <= not((layer0_outputs(4108)) or (layer0_outputs(2145)));
    layer1_outputs(3740) <= not(layer0_outputs(4222));
    layer1_outputs(3741) <= layer0_outputs(282);
    layer1_outputs(3742) <= not(layer0_outputs(577)) or (layer0_outputs(3999));
    layer1_outputs(3743) <= (layer0_outputs(2184)) and (layer0_outputs(4160));
    layer1_outputs(3744) <= layer0_outputs(4381);
    layer1_outputs(3745) <= not((layer0_outputs(3148)) and (layer0_outputs(1612)));
    layer1_outputs(3746) <= '0';
    layer1_outputs(3747) <= not(layer0_outputs(1921)) or (layer0_outputs(94));
    layer1_outputs(3748) <= not((layer0_outputs(4135)) or (layer0_outputs(2948)));
    layer1_outputs(3749) <= not((layer0_outputs(4726)) or (layer0_outputs(4623)));
    layer1_outputs(3750) <= (layer0_outputs(4593)) and not (layer0_outputs(2094));
    layer1_outputs(3751) <= not(layer0_outputs(2462)) or (layer0_outputs(4277));
    layer1_outputs(3752) <= not(layer0_outputs(913)) or (layer0_outputs(4678));
    layer1_outputs(3753) <= layer0_outputs(752);
    layer1_outputs(3754) <= not(layer0_outputs(380)) or (layer0_outputs(2864));
    layer1_outputs(3755) <= '0';
    layer1_outputs(3756) <= '0';
    layer1_outputs(3757) <= not((layer0_outputs(3152)) or (layer0_outputs(3793)));
    layer1_outputs(3758) <= (layer0_outputs(2601)) and not (layer0_outputs(2145));
    layer1_outputs(3759) <= '0';
    layer1_outputs(3760) <= not(layer0_outputs(4340));
    layer1_outputs(3761) <= (layer0_outputs(4878)) and not (layer0_outputs(34));
    layer1_outputs(3762) <= (layer0_outputs(1574)) or (layer0_outputs(1967));
    layer1_outputs(3763) <= not(layer0_outputs(3341));
    layer1_outputs(3764) <= not(layer0_outputs(1810));
    layer1_outputs(3765) <= not(layer0_outputs(4780));
    layer1_outputs(3766) <= not((layer0_outputs(1230)) or (layer0_outputs(1324)));
    layer1_outputs(3767) <= '0';
    layer1_outputs(3768) <= layer0_outputs(479);
    layer1_outputs(3769) <= not((layer0_outputs(3315)) xor (layer0_outputs(3067)));
    layer1_outputs(3770) <= layer0_outputs(2322);
    layer1_outputs(3771) <= not((layer0_outputs(1662)) and (layer0_outputs(1297)));
    layer1_outputs(3772) <= '1';
    layer1_outputs(3773) <= not(layer0_outputs(875));
    layer1_outputs(3774) <= not((layer0_outputs(246)) or (layer0_outputs(2666)));
    layer1_outputs(3775) <= not(layer0_outputs(1932));
    layer1_outputs(3776) <= '0';
    layer1_outputs(3777) <= not(layer0_outputs(4701));
    layer1_outputs(3778) <= (layer0_outputs(4444)) and (layer0_outputs(1491));
    layer1_outputs(3779) <= not(layer0_outputs(927)) or (layer0_outputs(1817));
    layer1_outputs(3780) <= (layer0_outputs(2618)) and not (layer0_outputs(1400));
    layer1_outputs(3781) <= not(layer0_outputs(1034)) or (layer0_outputs(685));
    layer1_outputs(3782) <= not(layer0_outputs(1098));
    layer1_outputs(3783) <= (layer0_outputs(4393)) and not (layer0_outputs(497));
    layer1_outputs(3784) <= (layer0_outputs(4134)) and (layer0_outputs(3563));
    layer1_outputs(3785) <= '0';
    layer1_outputs(3786) <= '1';
    layer1_outputs(3787) <= (layer0_outputs(1855)) and (layer0_outputs(2234));
    layer1_outputs(3788) <= not(layer0_outputs(4072)) or (layer0_outputs(1096));
    layer1_outputs(3789) <= not((layer0_outputs(1623)) and (layer0_outputs(717)));
    layer1_outputs(3790) <= (layer0_outputs(10)) or (layer0_outputs(672));
    layer1_outputs(3791) <= (layer0_outputs(3383)) and (layer0_outputs(1583));
    layer1_outputs(3792) <= layer0_outputs(656);
    layer1_outputs(3793) <= (layer0_outputs(401)) and not (layer0_outputs(2919));
    layer1_outputs(3794) <= '1';
    layer1_outputs(3795) <= not(layer0_outputs(2638));
    layer1_outputs(3796) <= layer0_outputs(2465);
    layer1_outputs(3797) <= not(layer0_outputs(912));
    layer1_outputs(3798) <= not(layer0_outputs(4573));
    layer1_outputs(3799) <= not(layer0_outputs(2676));
    layer1_outputs(3800) <= layer0_outputs(1653);
    layer1_outputs(3801) <= layer0_outputs(3329);
    layer1_outputs(3802) <= '0';
    layer1_outputs(3803) <= layer0_outputs(1011);
    layer1_outputs(3804) <= not(layer0_outputs(4159));
    layer1_outputs(3805) <= layer0_outputs(3211);
    layer1_outputs(3806) <= '0';
    layer1_outputs(3807) <= not((layer0_outputs(4902)) and (layer0_outputs(4462)));
    layer1_outputs(3808) <= (layer0_outputs(58)) and (layer0_outputs(4611));
    layer1_outputs(3809) <= (layer0_outputs(2968)) xor (layer0_outputs(2484));
    layer1_outputs(3810) <= layer0_outputs(4102);
    layer1_outputs(3811) <= not((layer0_outputs(3602)) and (layer0_outputs(1644)));
    layer1_outputs(3812) <= not((layer0_outputs(841)) and (layer0_outputs(761)));
    layer1_outputs(3813) <= not(layer0_outputs(4874)) or (layer0_outputs(1122));
    layer1_outputs(3814) <= layer0_outputs(2701);
    layer1_outputs(3815) <= (layer0_outputs(3066)) xor (layer0_outputs(2293));
    layer1_outputs(3816) <= (layer0_outputs(1050)) and (layer0_outputs(3086));
    layer1_outputs(3817) <= not((layer0_outputs(1075)) or (layer0_outputs(2099)));
    layer1_outputs(3818) <= not(layer0_outputs(4331));
    layer1_outputs(3819) <= not(layer0_outputs(1908)) or (layer0_outputs(1392));
    layer1_outputs(3820) <= (layer0_outputs(501)) or (layer0_outputs(126));
    layer1_outputs(3821) <= not(layer0_outputs(1749));
    layer1_outputs(3822) <= (layer0_outputs(3863)) and not (layer0_outputs(2221));
    layer1_outputs(3823) <= not((layer0_outputs(2669)) and (layer0_outputs(3162)));
    layer1_outputs(3824) <= '0';
    layer1_outputs(3825) <= (layer0_outputs(866)) and not (layer0_outputs(1024));
    layer1_outputs(3826) <= not(layer0_outputs(2834));
    layer1_outputs(3827) <= (layer0_outputs(3826)) and not (layer0_outputs(830));
    layer1_outputs(3828) <= not((layer0_outputs(5065)) or (layer0_outputs(1889)));
    layer1_outputs(3829) <= '0';
    layer1_outputs(3830) <= layer0_outputs(2247);
    layer1_outputs(3831) <= layer0_outputs(3011);
    layer1_outputs(3832) <= layer0_outputs(4339);
    layer1_outputs(3833) <= not((layer0_outputs(4204)) or (layer0_outputs(3859)));
    layer1_outputs(3834) <= (layer0_outputs(4973)) or (layer0_outputs(1596));
    layer1_outputs(3835) <= layer0_outputs(2602);
    layer1_outputs(3836) <= '1';
    layer1_outputs(3837) <= (layer0_outputs(278)) and not (layer0_outputs(2608));
    layer1_outputs(3838) <= not(layer0_outputs(4483)) or (layer0_outputs(2353));
    layer1_outputs(3839) <= '1';
    layer1_outputs(3840) <= not((layer0_outputs(3323)) or (layer0_outputs(4418)));
    layer1_outputs(3841) <= not((layer0_outputs(453)) and (layer0_outputs(95)));
    layer1_outputs(3842) <= '1';
    layer1_outputs(3843) <= '1';
    layer1_outputs(3844) <= (layer0_outputs(2232)) and (layer0_outputs(160));
    layer1_outputs(3845) <= not(layer0_outputs(17));
    layer1_outputs(3846) <= not(layer0_outputs(2553));
    layer1_outputs(3847) <= not((layer0_outputs(1132)) and (layer0_outputs(1996)));
    layer1_outputs(3848) <= (layer0_outputs(5032)) and (layer0_outputs(493));
    layer1_outputs(3849) <= (layer0_outputs(2603)) and (layer0_outputs(268));
    layer1_outputs(3850) <= not(layer0_outputs(4252));
    layer1_outputs(3851) <= '1';
    layer1_outputs(3852) <= layer0_outputs(3370);
    layer1_outputs(3853) <= not((layer0_outputs(2237)) and (layer0_outputs(4433)));
    layer1_outputs(3854) <= layer0_outputs(534);
    layer1_outputs(3855) <= '1';
    layer1_outputs(3856) <= '1';
    layer1_outputs(3857) <= layer0_outputs(2831);
    layer1_outputs(3858) <= (layer0_outputs(2062)) and not (layer0_outputs(1112));
    layer1_outputs(3859) <= '1';
    layer1_outputs(3860) <= (layer0_outputs(182)) and not (layer0_outputs(1640));
    layer1_outputs(3861) <= not(layer0_outputs(4137)) or (layer0_outputs(3760));
    layer1_outputs(3862) <= (layer0_outputs(4956)) or (layer0_outputs(4571));
    layer1_outputs(3863) <= '1';
    layer1_outputs(3864) <= '1';
    layer1_outputs(3865) <= not(layer0_outputs(1184)) or (layer0_outputs(3981));
    layer1_outputs(3866) <= '0';
    layer1_outputs(3867) <= layer0_outputs(935);
    layer1_outputs(3868) <= (layer0_outputs(1745)) and not (layer0_outputs(561));
    layer1_outputs(3869) <= '1';
    layer1_outputs(3870) <= (layer0_outputs(3842)) and not (layer0_outputs(3658));
    layer1_outputs(3871) <= not((layer0_outputs(1531)) xor (layer0_outputs(453)));
    layer1_outputs(3872) <= layer0_outputs(4775);
    layer1_outputs(3873) <= not((layer0_outputs(3431)) and (layer0_outputs(4240)));
    layer1_outputs(3874) <= not(layer0_outputs(2654)) or (layer0_outputs(3774));
    layer1_outputs(3875) <= '1';
    layer1_outputs(3876) <= layer0_outputs(3214);
    layer1_outputs(3877) <= (layer0_outputs(4885)) and not (layer0_outputs(5054));
    layer1_outputs(3878) <= layer0_outputs(4006);
    layer1_outputs(3879) <= layer0_outputs(1593);
    layer1_outputs(3880) <= not(layer0_outputs(381));
    layer1_outputs(3881) <= not((layer0_outputs(4383)) and (layer0_outputs(2833)));
    layer1_outputs(3882) <= not((layer0_outputs(3977)) or (layer0_outputs(1837)));
    layer1_outputs(3883) <= '1';
    layer1_outputs(3884) <= not((layer0_outputs(4510)) and (layer0_outputs(46)));
    layer1_outputs(3885) <= layer0_outputs(1750);
    layer1_outputs(3886) <= layer0_outputs(2663);
    layer1_outputs(3887) <= (layer0_outputs(1586)) and not (layer0_outputs(229));
    layer1_outputs(3888) <= '0';
    layer1_outputs(3889) <= not(layer0_outputs(3100)) or (layer0_outputs(2812));
    layer1_outputs(3890) <= (layer0_outputs(2165)) and not (layer0_outputs(2121));
    layer1_outputs(3891) <= layer0_outputs(4792);
    layer1_outputs(3892) <= (layer0_outputs(640)) xor (layer0_outputs(2936));
    layer1_outputs(3893) <= not(layer0_outputs(567));
    layer1_outputs(3894) <= (layer0_outputs(3647)) or (layer0_outputs(2060));
    layer1_outputs(3895) <= '1';
    layer1_outputs(3896) <= (layer0_outputs(2325)) and not (layer0_outputs(2527));
    layer1_outputs(3897) <= (layer0_outputs(3593)) and not (layer0_outputs(926));
    layer1_outputs(3898) <= layer0_outputs(2667);
    layer1_outputs(3899) <= not((layer0_outputs(848)) or (layer0_outputs(3621)));
    layer1_outputs(3900) <= (layer0_outputs(772)) and (layer0_outputs(4791));
    layer1_outputs(3901) <= (layer0_outputs(3593)) and (layer0_outputs(1101));
    layer1_outputs(3902) <= layer0_outputs(3701);
    layer1_outputs(3903) <= (layer0_outputs(4555)) or (layer0_outputs(3809));
    layer1_outputs(3904) <= not(layer0_outputs(1582)) or (layer0_outputs(3965));
    layer1_outputs(3905) <= not(layer0_outputs(2775));
    layer1_outputs(3906) <= not(layer0_outputs(1895)) or (layer0_outputs(1869));
    layer1_outputs(3907) <= not((layer0_outputs(750)) and (layer0_outputs(2734)));
    layer1_outputs(3908) <= layer0_outputs(3340);
    layer1_outputs(3909) <= not(layer0_outputs(973)) or (layer0_outputs(1265));
    layer1_outputs(3910) <= not((layer0_outputs(2137)) and (layer0_outputs(90)));
    layer1_outputs(3911) <= not((layer0_outputs(2022)) or (layer0_outputs(794)));
    layer1_outputs(3912) <= (layer0_outputs(725)) and (layer0_outputs(4194));
    layer1_outputs(3913) <= (layer0_outputs(434)) and not (layer0_outputs(418));
    layer1_outputs(3914) <= not(layer0_outputs(3810)) or (layer0_outputs(4976));
    layer1_outputs(3915) <= layer0_outputs(1418);
    layer1_outputs(3916) <= not(layer0_outputs(2422));
    layer1_outputs(3917) <= not((layer0_outputs(4974)) or (layer0_outputs(4500)));
    layer1_outputs(3918) <= layer0_outputs(5038);
    layer1_outputs(3919) <= '0';
    layer1_outputs(3920) <= (layer0_outputs(141)) or (layer0_outputs(2643));
    layer1_outputs(3921) <= not(layer0_outputs(4075)) or (layer0_outputs(2621));
    layer1_outputs(3922) <= not((layer0_outputs(4732)) or (layer0_outputs(810)));
    layer1_outputs(3923) <= (layer0_outputs(4584)) and not (layer0_outputs(2538));
    layer1_outputs(3924) <= layer0_outputs(1545);
    layer1_outputs(3925) <= (layer0_outputs(4007)) and not (layer0_outputs(806));
    layer1_outputs(3926) <= not(layer0_outputs(817)) or (layer0_outputs(371));
    layer1_outputs(3927) <= (layer0_outputs(1626)) and not (layer0_outputs(4480));
    layer1_outputs(3928) <= layer0_outputs(1960);
    layer1_outputs(3929) <= '1';
    layer1_outputs(3930) <= (layer0_outputs(395)) and (layer0_outputs(3968));
    layer1_outputs(3931) <= '1';
    layer1_outputs(3932) <= (layer0_outputs(504)) or (layer0_outputs(1092));
    layer1_outputs(3933) <= '0';
    layer1_outputs(3934) <= '0';
    layer1_outputs(3935) <= layer0_outputs(3362);
    layer1_outputs(3936) <= (layer0_outputs(1972)) and not (layer0_outputs(4543));
    layer1_outputs(3937) <= not(layer0_outputs(4333)) or (layer0_outputs(4938));
    layer1_outputs(3938) <= (layer0_outputs(1730)) or (layer0_outputs(332));
    layer1_outputs(3939) <= '1';
    layer1_outputs(3940) <= not(layer0_outputs(3452)) or (layer0_outputs(560));
    layer1_outputs(3941) <= not(layer0_outputs(3702)) or (layer0_outputs(2920));
    layer1_outputs(3942) <= not((layer0_outputs(2447)) xor (layer0_outputs(2006)));
    layer1_outputs(3943) <= layer0_outputs(792);
    layer1_outputs(3944) <= not(layer0_outputs(4710)) or (layer0_outputs(573));
    layer1_outputs(3945) <= layer0_outputs(2624);
    layer1_outputs(3946) <= '1';
    layer1_outputs(3947) <= layer0_outputs(4124);
    layer1_outputs(3948) <= not(layer0_outputs(1637)) or (layer0_outputs(3374));
    layer1_outputs(3949) <= not(layer0_outputs(2887)) or (layer0_outputs(597));
    layer1_outputs(3950) <= not((layer0_outputs(4930)) or (layer0_outputs(3852)));
    layer1_outputs(3951) <= not((layer0_outputs(1630)) and (layer0_outputs(1414)));
    layer1_outputs(3952) <= not((layer0_outputs(2007)) and (layer0_outputs(3594)));
    layer1_outputs(3953) <= not((layer0_outputs(2448)) or (layer0_outputs(4032)));
    layer1_outputs(3954) <= not((layer0_outputs(3220)) and (layer0_outputs(3421)));
    layer1_outputs(3955) <= not((layer0_outputs(529)) or (layer0_outputs(4851)));
    layer1_outputs(3956) <= (layer0_outputs(593)) and not (layer0_outputs(69));
    layer1_outputs(3957) <= not(layer0_outputs(339));
    layer1_outputs(3958) <= not((layer0_outputs(2857)) xor (layer0_outputs(732)));
    layer1_outputs(3959) <= layer0_outputs(2412);
    layer1_outputs(3960) <= not((layer0_outputs(2206)) and (layer0_outputs(4226)));
    layer1_outputs(3961) <= '0';
    layer1_outputs(3962) <= not(layer0_outputs(1889)) or (layer0_outputs(652));
    layer1_outputs(3963) <= '0';
    layer1_outputs(3964) <= not(layer0_outputs(1042)) or (layer0_outputs(159));
    layer1_outputs(3965) <= '0';
    layer1_outputs(3966) <= (layer0_outputs(4246)) and not (layer0_outputs(1838));
    layer1_outputs(3967) <= (layer0_outputs(3720)) and (layer0_outputs(4404));
    layer1_outputs(3968) <= not(layer0_outputs(3433));
    layer1_outputs(3969) <= (layer0_outputs(1555)) or (layer0_outputs(1197));
    layer1_outputs(3970) <= layer0_outputs(3630);
    layer1_outputs(3971) <= (layer0_outputs(1345)) and not (layer0_outputs(293));
    layer1_outputs(3972) <= not(layer0_outputs(1848)) or (layer0_outputs(1391));
    layer1_outputs(3973) <= layer0_outputs(1317);
    layer1_outputs(3974) <= '1';
    layer1_outputs(3975) <= layer0_outputs(2548);
    layer1_outputs(3976) <= (layer0_outputs(390)) or (layer0_outputs(872));
    layer1_outputs(3977) <= layer0_outputs(1076);
    layer1_outputs(3978) <= (layer0_outputs(4689)) or (layer0_outputs(1301));
    layer1_outputs(3979) <= (layer0_outputs(4200)) and not (layer0_outputs(2876));
    layer1_outputs(3980) <= (layer0_outputs(3176)) and not (layer0_outputs(1038));
    layer1_outputs(3981) <= (layer0_outputs(2516)) and not (layer0_outputs(4150));
    layer1_outputs(3982) <= layer0_outputs(2353);
    layer1_outputs(3983) <= layer0_outputs(305);
    layer1_outputs(3984) <= layer0_outputs(4705);
    layer1_outputs(3985) <= not((layer0_outputs(1919)) and (layer0_outputs(1014)));
    layer1_outputs(3986) <= '0';
    layer1_outputs(3987) <= not(layer0_outputs(2080)) or (layer0_outputs(2471));
    layer1_outputs(3988) <= (layer0_outputs(3908)) and not (layer0_outputs(4684));
    layer1_outputs(3989) <= (layer0_outputs(3861)) and not (layer0_outputs(600));
    layer1_outputs(3990) <= not(layer0_outputs(1879)) or (layer0_outputs(1119));
    layer1_outputs(3991) <= (layer0_outputs(3799)) and (layer0_outputs(3556));
    layer1_outputs(3992) <= not(layer0_outputs(1212));
    layer1_outputs(3993) <= not((layer0_outputs(3989)) or (layer0_outputs(2300)));
    layer1_outputs(3994) <= (layer0_outputs(4684)) xor (layer0_outputs(3935));
    layer1_outputs(3995) <= not(layer0_outputs(2870)) or (layer0_outputs(4309));
    layer1_outputs(3996) <= not((layer0_outputs(92)) and (layer0_outputs(2236)));
    layer1_outputs(3997) <= not((layer0_outputs(1389)) or (layer0_outputs(1119)));
    layer1_outputs(3998) <= layer0_outputs(1603);
    layer1_outputs(3999) <= (layer0_outputs(4615)) or (layer0_outputs(1105));
    layer1_outputs(4000) <= not((layer0_outputs(2742)) or (layer0_outputs(752)));
    layer1_outputs(4001) <= (layer0_outputs(4695)) and not (layer0_outputs(3570));
    layer1_outputs(4002) <= not((layer0_outputs(4622)) xor (layer0_outputs(2490)));
    layer1_outputs(4003) <= not(layer0_outputs(4067)) or (layer0_outputs(3462));
    layer1_outputs(4004) <= '1';
    layer1_outputs(4005) <= (layer0_outputs(1995)) and (layer0_outputs(3124));
    layer1_outputs(4006) <= (layer0_outputs(2156)) and not (layer0_outputs(2814));
    layer1_outputs(4007) <= not(layer0_outputs(3417));
    layer1_outputs(4008) <= '0';
    layer1_outputs(4009) <= not(layer0_outputs(2429));
    layer1_outputs(4010) <= layer0_outputs(685);
    layer1_outputs(4011) <= not(layer0_outputs(2934));
    layer1_outputs(4012) <= not((layer0_outputs(1758)) or (layer0_outputs(1698)));
    layer1_outputs(4013) <= not(layer0_outputs(3428));
    layer1_outputs(4014) <= '0';
    layer1_outputs(4015) <= not(layer0_outputs(849)) or (layer0_outputs(4231));
    layer1_outputs(4016) <= (layer0_outputs(1465)) or (layer0_outputs(5107));
    layer1_outputs(4017) <= '0';
    layer1_outputs(4018) <= not(layer0_outputs(1288)) or (layer0_outputs(4186));
    layer1_outputs(4019) <= not((layer0_outputs(3462)) and (layer0_outputs(4167)));
    layer1_outputs(4020) <= (layer0_outputs(2617)) and (layer0_outputs(1380));
    layer1_outputs(4021) <= not(layer0_outputs(783)) or (layer0_outputs(4147));
    layer1_outputs(4022) <= '0';
    layer1_outputs(4023) <= not((layer0_outputs(284)) or (layer0_outputs(2539)));
    layer1_outputs(4024) <= '0';
    layer1_outputs(4025) <= (layer0_outputs(3980)) and not (layer0_outputs(567));
    layer1_outputs(4026) <= not((layer0_outputs(523)) and (layer0_outputs(827)));
    layer1_outputs(4027) <= (layer0_outputs(587)) and (layer0_outputs(3088));
    layer1_outputs(4028) <= '1';
    layer1_outputs(4029) <= not((layer0_outputs(2757)) or (layer0_outputs(4375)));
    layer1_outputs(4030) <= (layer0_outputs(1749)) or (layer0_outputs(1523));
    layer1_outputs(4031) <= layer0_outputs(1892);
    layer1_outputs(4032) <= layer0_outputs(164);
    layer1_outputs(4033) <= layer0_outputs(3782);
    layer1_outputs(4034) <= layer0_outputs(3047);
    layer1_outputs(4035) <= layer0_outputs(1922);
    layer1_outputs(4036) <= (layer0_outputs(2993)) and not (layer0_outputs(4085));
    layer1_outputs(4037) <= (layer0_outputs(2114)) and (layer0_outputs(2646));
    layer1_outputs(4038) <= (layer0_outputs(1357)) and not (layer0_outputs(3730));
    layer1_outputs(4039) <= layer0_outputs(1226);
    layer1_outputs(4040) <= layer0_outputs(3033);
    layer1_outputs(4041) <= not(layer0_outputs(2189));
    layer1_outputs(4042) <= not(layer0_outputs(791)) or (layer0_outputs(1399));
    layer1_outputs(4043) <= not(layer0_outputs(1893));
    layer1_outputs(4044) <= not(layer0_outputs(1291));
    layer1_outputs(4045) <= layer0_outputs(3266);
    layer1_outputs(4046) <= not((layer0_outputs(3975)) and (layer0_outputs(2094)));
    layer1_outputs(4047) <= (layer0_outputs(1900)) or (layer0_outputs(4539));
    layer1_outputs(4048) <= not((layer0_outputs(1389)) and (layer0_outputs(1013)));
    layer1_outputs(4049) <= '1';
    layer1_outputs(4050) <= '0';
    layer1_outputs(4051) <= not((layer0_outputs(3692)) and (layer0_outputs(4377)));
    layer1_outputs(4052) <= not((layer0_outputs(837)) or (layer0_outputs(2100)));
    layer1_outputs(4053) <= not(layer0_outputs(2861)) or (layer0_outputs(753));
    layer1_outputs(4054) <= not(layer0_outputs(2568)) or (layer0_outputs(4266));
    layer1_outputs(4055) <= (layer0_outputs(2813)) and not (layer0_outputs(4915));
    layer1_outputs(4056) <= layer0_outputs(3603);
    layer1_outputs(4057) <= '1';
    layer1_outputs(4058) <= '0';
    layer1_outputs(4059) <= layer0_outputs(1074);
    layer1_outputs(4060) <= (layer0_outputs(3443)) and not (layer0_outputs(4692));
    layer1_outputs(4061) <= not(layer0_outputs(4942));
    layer1_outputs(4062) <= (layer0_outputs(4366)) and (layer0_outputs(4591));
    layer1_outputs(4063) <= layer0_outputs(1359);
    layer1_outputs(4064) <= '1';
    layer1_outputs(4065) <= layer0_outputs(1325);
    layer1_outputs(4066) <= not(layer0_outputs(1061)) or (layer0_outputs(2266));
    layer1_outputs(4067) <= layer0_outputs(3815);
    layer1_outputs(4068) <= (layer0_outputs(1383)) and (layer0_outputs(2975));
    layer1_outputs(4069) <= not(layer0_outputs(4847)) or (layer0_outputs(346));
    layer1_outputs(4070) <= layer0_outputs(461);
    layer1_outputs(4071) <= not((layer0_outputs(2416)) or (layer0_outputs(2761)));
    layer1_outputs(4072) <= not((layer0_outputs(4662)) xor (layer0_outputs(3300)));
    layer1_outputs(4073) <= (layer0_outputs(644)) or (layer0_outputs(1256));
    layer1_outputs(4074) <= not((layer0_outputs(4899)) and (layer0_outputs(1757)));
    layer1_outputs(4075) <= layer0_outputs(2998);
    layer1_outputs(4076) <= not(layer0_outputs(3378)) or (layer0_outputs(860));
    layer1_outputs(4077) <= not((layer0_outputs(641)) or (layer0_outputs(4033)));
    layer1_outputs(4078) <= '1';
    layer1_outputs(4079) <= not(layer0_outputs(2758));
    layer1_outputs(4080) <= (layer0_outputs(1777)) and not (layer0_outputs(3862));
    layer1_outputs(4081) <= layer0_outputs(1235);
    layer1_outputs(4082) <= (layer0_outputs(120)) and not (layer0_outputs(4848));
    layer1_outputs(4083) <= layer0_outputs(4198);
    layer1_outputs(4084) <= (layer0_outputs(861)) and not (layer0_outputs(725));
    layer1_outputs(4085) <= layer0_outputs(327);
    layer1_outputs(4086) <= not((layer0_outputs(2508)) and (layer0_outputs(651)));
    layer1_outputs(4087) <= not((layer0_outputs(3317)) xor (layer0_outputs(1596)));
    layer1_outputs(4088) <= (layer0_outputs(2724)) or (layer0_outputs(4601));
    layer1_outputs(4089) <= '0';
    layer1_outputs(4090) <= not(layer0_outputs(3382)) or (layer0_outputs(2934));
    layer1_outputs(4091) <= not(layer0_outputs(4785));
    layer1_outputs(4092) <= not(layer0_outputs(2885)) or (layer0_outputs(2));
    layer1_outputs(4093) <= not(layer0_outputs(584));
    layer1_outputs(4094) <= not(layer0_outputs(1471)) or (layer0_outputs(1687));
    layer1_outputs(4095) <= (layer0_outputs(1246)) or (layer0_outputs(5029));
    layer1_outputs(4096) <= '0';
    layer1_outputs(4097) <= (layer0_outputs(3463)) and not (layer0_outputs(2715));
    layer1_outputs(4098) <= not((layer0_outputs(291)) and (layer0_outputs(4781)));
    layer1_outputs(4099) <= (layer0_outputs(2448)) and not (layer0_outputs(4770));
    layer1_outputs(4100) <= not(layer0_outputs(106));
    layer1_outputs(4101) <= (layer0_outputs(1746)) and not (layer0_outputs(3259));
    layer1_outputs(4102) <= (layer0_outputs(2290)) or (layer0_outputs(4100));
    layer1_outputs(4103) <= '0';
    layer1_outputs(4104) <= '1';
    layer1_outputs(4105) <= (layer0_outputs(2434)) and not (layer0_outputs(3897));
    layer1_outputs(4106) <= layer0_outputs(3004);
    layer1_outputs(4107) <= layer0_outputs(2696);
    layer1_outputs(4108) <= '0';
    layer1_outputs(4109) <= not(layer0_outputs(1841));
    layer1_outputs(4110) <= (layer0_outputs(3261)) or (layer0_outputs(4837));
    layer1_outputs(4111) <= not(layer0_outputs(4148));
    layer1_outputs(4112) <= not((layer0_outputs(4288)) and (layer0_outputs(1052)));
    layer1_outputs(4113) <= (layer0_outputs(12)) and (layer0_outputs(4695));
    layer1_outputs(4114) <= (layer0_outputs(4850)) and not (layer0_outputs(4574));
    layer1_outputs(4115) <= layer0_outputs(2499);
    layer1_outputs(4116) <= layer0_outputs(1657);
    layer1_outputs(4117) <= '0';
    layer1_outputs(4118) <= not(layer0_outputs(3652));
    layer1_outputs(4119) <= not((layer0_outputs(2031)) and (layer0_outputs(1678)));
    layer1_outputs(4120) <= not(layer0_outputs(3771));
    layer1_outputs(4121) <= layer0_outputs(1502);
    layer1_outputs(4122) <= not((layer0_outputs(3237)) and (layer0_outputs(1054)));
    layer1_outputs(4123) <= (layer0_outputs(1040)) and (layer0_outputs(2197));
    layer1_outputs(4124) <= not((layer0_outputs(3917)) or (layer0_outputs(1713)));
    layer1_outputs(4125) <= not((layer0_outputs(2789)) and (layer0_outputs(3740)));
    layer1_outputs(4126) <= layer0_outputs(4785);
    layer1_outputs(4127) <= not((layer0_outputs(378)) or (layer0_outputs(4318)));
    layer1_outputs(4128) <= (layer0_outputs(3131)) and not (layer0_outputs(1227));
    layer1_outputs(4129) <= not((layer0_outputs(3475)) xor (layer0_outputs(4752)));
    layer1_outputs(4130) <= layer0_outputs(1841);
    layer1_outputs(4131) <= not(layer0_outputs(830)) or (layer0_outputs(2367));
    layer1_outputs(4132) <= not(layer0_outputs(4515)) or (layer0_outputs(4043));
    layer1_outputs(4133) <= (layer0_outputs(3831)) or (layer0_outputs(3257));
    layer1_outputs(4134) <= (layer0_outputs(3038)) and (layer0_outputs(4118));
    layer1_outputs(4135) <= (layer0_outputs(2623)) and not (layer0_outputs(4947));
    layer1_outputs(4136) <= (layer0_outputs(3111)) and not (layer0_outputs(2542));
    layer1_outputs(4137) <= not((layer0_outputs(3425)) and (layer0_outputs(2924)));
    layer1_outputs(4138) <= (layer0_outputs(233)) or (layer0_outputs(2941));
    layer1_outputs(4139) <= (layer0_outputs(3846)) or (layer0_outputs(3788));
    layer1_outputs(4140) <= (layer0_outputs(2583)) or (layer0_outputs(223));
    layer1_outputs(4141) <= not(layer0_outputs(4727));
    layer1_outputs(4142) <= not(layer0_outputs(2406));
    layer1_outputs(4143) <= layer0_outputs(367);
    layer1_outputs(4144) <= layer0_outputs(5095);
    layer1_outputs(4145) <= not((layer0_outputs(978)) xor (layer0_outputs(1514)));
    layer1_outputs(4146) <= not((layer0_outputs(2799)) or (layer0_outputs(2187)));
    layer1_outputs(4147) <= (layer0_outputs(4349)) and not (layer0_outputs(1037));
    layer1_outputs(4148) <= not(layer0_outputs(308));
    layer1_outputs(4149) <= not((layer0_outputs(4605)) and (layer0_outputs(33)));
    layer1_outputs(4150) <= (layer0_outputs(1407)) and not (layer0_outputs(3660));
    layer1_outputs(4151) <= not(layer0_outputs(4271)) or (layer0_outputs(2972));
    layer1_outputs(4152) <= not(layer0_outputs(4841)) or (layer0_outputs(1121));
    layer1_outputs(4153) <= (layer0_outputs(2154)) and not (layer0_outputs(4573));
    layer1_outputs(4154) <= '1';
    layer1_outputs(4155) <= '1';
    layer1_outputs(4156) <= (layer0_outputs(3805)) or (layer0_outputs(3135));
    layer1_outputs(4157) <= not(layer0_outputs(2306));
    layer1_outputs(4158) <= (layer0_outputs(4022)) or (layer0_outputs(3591));
    layer1_outputs(4159) <= (layer0_outputs(3325)) and not (layer0_outputs(195));
    layer1_outputs(4160) <= '0';
    layer1_outputs(4161) <= (layer0_outputs(1904)) and (layer0_outputs(4789));
    layer1_outputs(4162) <= not(layer0_outputs(1055));
    layer1_outputs(4163) <= layer0_outputs(998);
    layer1_outputs(4164) <= (layer0_outputs(1574)) or (layer0_outputs(183));
    layer1_outputs(4165) <= layer0_outputs(2518);
    layer1_outputs(4166) <= not(layer0_outputs(4552));
    layer1_outputs(4167) <= '0';
    layer1_outputs(4168) <= (layer0_outputs(180)) or (layer0_outputs(2101));
    layer1_outputs(4169) <= layer0_outputs(3641);
    layer1_outputs(4170) <= layer0_outputs(3189);
    layer1_outputs(4171) <= layer0_outputs(4231);
    layer1_outputs(4172) <= '1';
    layer1_outputs(4173) <= layer0_outputs(2292);
    layer1_outputs(4174) <= '1';
    layer1_outputs(4175) <= layer0_outputs(1595);
    layer1_outputs(4176) <= '0';
    layer1_outputs(4177) <= not(layer0_outputs(4688));
    layer1_outputs(4178) <= not((layer0_outputs(1549)) and (layer0_outputs(3959)));
    layer1_outputs(4179) <= (layer0_outputs(4560)) or (layer0_outputs(893));
    layer1_outputs(4180) <= not(layer0_outputs(2664)) or (layer0_outputs(86));
    layer1_outputs(4181) <= (layer0_outputs(1413)) and not (layer0_outputs(573));
    layer1_outputs(4182) <= '1';
    layer1_outputs(4183) <= '1';
    layer1_outputs(4184) <= not(layer0_outputs(2653));
    layer1_outputs(4185) <= (layer0_outputs(2590)) and not (layer0_outputs(3888));
    layer1_outputs(4186) <= not((layer0_outputs(928)) or (layer0_outputs(4354)));
    layer1_outputs(4187) <= not(layer0_outputs(1755));
    layer1_outputs(4188) <= layer0_outputs(527);
    layer1_outputs(4189) <= (layer0_outputs(3115)) and not (layer0_outputs(364));
    layer1_outputs(4190) <= not(layer0_outputs(404)) or (layer0_outputs(728));
    layer1_outputs(4191) <= (layer0_outputs(1235)) and not (layer0_outputs(1741));
    layer1_outputs(4192) <= (layer0_outputs(1930)) or (layer0_outputs(1109));
    layer1_outputs(4193) <= layer0_outputs(4856);
    layer1_outputs(4194) <= not((layer0_outputs(2522)) and (layer0_outputs(1920)));
    layer1_outputs(4195) <= not(layer0_outputs(1462)) or (layer0_outputs(1433));
    layer1_outputs(4196) <= not(layer0_outputs(2037)) or (layer0_outputs(939));
    layer1_outputs(4197) <= not((layer0_outputs(780)) or (layer0_outputs(1398)));
    layer1_outputs(4198) <= (layer0_outputs(487)) or (layer0_outputs(1025));
    layer1_outputs(4199) <= (layer0_outputs(2499)) or (layer0_outputs(1579));
    layer1_outputs(4200) <= layer0_outputs(2935);
    layer1_outputs(4201) <= not(layer0_outputs(507)) or (layer0_outputs(4490));
    layer1_outputs(4202) <= layer0_outputs(2534);
    layer1_outputs(4203) <= not((layer0_outputs(553)) and (layer0_outputs(1022)));
    layer1_outputs(4204) <= (layer0_outputs(3546)) and not (layer0_outputs(646));
    layer1_outputs(4205) <= not(layer0_outputs(505)) or (layer0_outputs(4595));
    layer1_outputs(4206) <= '1';
    layer1_outputs(4207) <= (layer0_outputs(2783)) or (layer0_outputs(83));
    layer1_outputs(4208) <= not(layer0_outputs(511));
    layer1_outputs(4209) <= not(layer0_outputs(1215));
    layer1_outputs(4210) <= not((layer0_outputs(4717)) or (layer0_outputs(2180)));
    layer1_outputs(4211) <= not((layer0_outputs(2286)) and (layer0_outputs(91)));
    layer1_outputs(4212) <= (layer0_outputs(3963)) and not (layer0_outputs(4395));
    layer1_outputs(4213) <= '0';
    layer1_outputs(4214) <= not((layer0_outputs(2004)) or (layer0_outputs(4409)));
    layer1_outputs(4215) <= not((layer0_outputs(3210)) and (layer0_outputs(1082)));
    layer1_outputs(4216) <= not((layer0_outputs(330)) or (layer0_outputs(2937)));
    layer1_outputs(4217) <= '0';
    layer1_outputs(4218) <= not(layer0_outputs(3815));
    layer1_outputs(4219) <= layer0_outputs(4416);
    layer1_outputs(4220) <= (layer0_outputs(4855)) and not (layer0_outputs(57));
    layer1_outputs(4221) <= '0';
    layer1_outputs(4222) <= layer0_outputs(2398);
    layer1_outputs(4223) <= layer0_outputs(5001);
    layer1_outputs(4224) <= (layer0_outputs(4357)) and not (layer0_outputs(292));
    layer1_outputs(4225) <= not(layer0_outputs(3552)) or (layer0_outputs(2580));
    layer1_outputs(4226) <= layer0_outputs(4544);
    layer1_outputs(4227) <= '0';
    layer1_outputs(4228) <= '1';
    layer1_outputs(4229) <= (layer0_outputs(3064)) or (layer0_outputs(3974));
    layer1_outputs(4230) <= not(layer0_outputs(611));
    layer1_outputs(4231) <= (layer0_outputs(568)) and not (layer0_outputs(2614));
    layer1_outputs(4232) <= not(layer0_outputs(248)) or (layer0_outputs(921));
    layer1_outputs(4233) <= (layer0_outputs(3821)) and not (layer0_outputs(635));
    layer1_outputs(4234) <= '0';
    layer1_outputs(4235) <= not((layer0_outputs(4493)) and (layer0_outputs(3980)));
    layer1_outputs(4236) <= '1';
    layer1_outputs(4237) <= layer0_outputs(3046);
    layer1_outputs(4238) <= layer0_outputs(1050);
    layer1_outputs(4239) <= (layer0_outputs(4481)) or (layer0_outputs(4449));
    layer1_outputs(4240) <= '0';
    layer1_outputs(4241) <= not(layer0_outputs(604));
    layer1_outputs(4242) <= '0';
    layer1_outputs(4243) <= (layer0_outputs(2159)) or (layer0_outputs(3765));
    layer1_outputs(4244) <= '1';
    layer1_outputs(4245) <= not((layer0_outputs(4422)) xor (layer0_outputs(1807)));
    layer1_outputs(4246) <= not(layer0_outputs(1970)) or (layer0_outputs(3531));
    layer1_outputs(4247) <= layer0_outputs(65);
    layer1_outputs(4248) <= not(layer0_outputs(2212));
    layer1_outputs(4249) <= not(layer0_outputs(1548));
    layer1_outputs(4250) <= layer0_outputs(1067);
    layer1_outputs(4251) <= not((layer0_outputs(3291)) and (layer0_outputs(263)));
    layer1_outputs(4252) <= not(layer0_outputs(4956));
    layer1_outputs(4253) <= not(layer0_outputs(2064)) or (layer0_outputs(3548));
    layer1_outputs(4254) <= '1';
    layer1_outputs(4255) <= (layer0_outputs(2445)) or (layer0_outputs(4890));
    layer1_outputs(4256) <= (layer0_outputs(5048)) and (layer0_outputs(4131));
    layer1_outputs(4257) <= (layer0_outputs(2001)) and not (layer0_outputs(1172));
    layer1_outputs(4258) <= not(layer0_outputs(4752));
    layer1_outputs(4259) <= (layer0_outputs(1521)) and not (layer0_outputs(4912));
    layer1_outputs(4260) <= not((layer0_outputs(1557)) or (layer0_outputs(3083)));
    layer1_outputs(4261) <= not(layer0_outputs(4332)) or (layer0_outputs(3655));
    layer1_outputs(4262) <= (layer0_outputs(490)) and (layer0_outputs(528));
    layer1_outputs(4263) <= '1';
    layer1_outputs(4264) <= (layer0_outputs(1979)) and not (layer0_outputs(1839));
    layer1_outputs(4265) <= not((layer0_outputs(76)) or (layer0_outputs(2811)));
    layer1_outputs(4266) <= '1';
    layer1_outputs(4267) <= layer0_outputs(3311);
    layer1_outputs(4268) <= (layer0_outputs(2410)) and not (layer0_outputs(4619));
    layer1_outputs(4269) <= (layer0_outputs(2158)) and not (layer0_outputs(2953));
    layer1_outputs(4270) <= '1';
    layer1_outputs(4271) <= layer0_outputs(175);
    layer1_outputs(4272) <= not(layer0_outputs(701)) or (layer0_outputs(1969));
    layer1_outputs(4273) <= (layer0_outputs(4)) and (layer0_outputs(100));
    layer1_outputs(4274) <= not(layer0_outputs(2356)) or (layer0_outputs(1374));
    layer1_outputs(4275) <= (layer0_outputs(3607)) and (layer0_outputs(2526));
    layer1_outputs(4276) <= not(layer0_outputs(632));
    layer1_outputs(4277) <= '1';
    layer1_outputs(4278) <= not((layer0_outputs(1985)) and (layer0_outputs(3225)));
    layer1_outputs(4279) <= (layer0_outputs(2250)) or (layer0_outputs(2729));
    layer1_outputs(4280) <= layer0_outputs(4177);
    layer1_outputs(4281) <= (layer0_outputs(4)) and (layer0_outputs(4302));
    layer1_outputs(4282) <= (layer0_outputs(4058)) and not (layer0_outputs(2530));
    layer1_outputs(4283) <= not(layer0_outputs(2177)) or (layer0_outputs(2606));
    layer1_outputs(4284) <= (layer0_outputs(2383)) or (layer0_outputs(1787));
    layer1_outputs(4285) <= not((layer0_outputs(757)) and (layer0_outputs(1019)));
    layer1_outputs(4286) <= (layer0_outputs(3864)) and not (layer0_outputs(4206));
    layer1_outputs(4287) <= (layer0_outputs(53)) and not (layer0_outputs(1625));
    layer1_outputs(4288) <= (layer0_outputs(197)) and not (layer0_outputs(4447));
    layer1_outputs(4289) <= not((layer0_outputs(19)) and (layer0_outputs(3474)));
    layer1_outputs(4290) <= (layer0_outputs(1410)) and (layer0_outputs(4135));
    layer1_outputs(4291) <= layer0_outputs(3319);
    layer1_outputs(4292) <= not((layer0_outputs(4469)) and (layer0_outputs(69)));
    layer1_outputs(4293) <= not((layer0_outputs(75)) and (layer0_outputs(4889)));
    layer1_outputs(4294) <= '1';
    layer1_outputs(4295) <= (layer0_outputs(227)) and not (layer0_outputs(4459));
    layer1_outputs(4296) <= not(layer0_outputs(2420));
    layer1_outputs(4297) <= not((layer0_outputs(2260)) or (layer0_outputs(622)));
    layer1_outputs(4298) <= layer0_outputs(855);
    layer1_outputs(4299) <= not(layer0_outputs(3293));
    layer1_outputs(4300) <= '1';
    layer1_outputs(4301) <= not(layer0_outputs(1202));
    layer1_outputs(4302) <= '1';
    layer1_outputs(4303) <= not(layer0_outputs(4784));
    layer1_outputs(4304) <= not((layer0_outputs(2824)) and (layer0_outputs(1860)));
    layer1_outputs(4305) <= not((layer0_outputs(4185)) and (layer0_outputs(4089)));
    layer1_outputs(4306) <= not(layer0_outputs(1008)) or (layer0_outputs(3237));
    layer1_outputs(4307) <= not(layer0_outputs(2660));
    layer1_outputs(4308) <= (layer0_outputs(643)) and not (layer0_outputs(3879));
    layer1_outputs(4309) <= not((layer0_outputs(2864)) or (layer0_outputs(1710)));
    layer1_outputs(4310) <= not(layer0_outputs(1946));
    layer1_outputs(4311) <= not((layer0_outputs(3626)) and (layer0_outputs(1703)));
    layer1_outputs(4312) <= (layer0_outputs(3114)) and not (layer0_outputs(2776));
    layer1_outputs(4313) <= '0';
    layer1_outputs(4314) <= not(layer0_outputs(3761));
    layer1_outputs(4315) <= not((layer0_outputs(1427)) xor (layer0_outputs(4243)));
    layer1_outputs(4316) <= '0';
    layer1_outputs(4317) <= not(layer0_outputs(2459)) or (layer0_outputs(1097));
    layer1_outputs(4318) <= (layer0_outputs(1786)) and not (layer0_outputs(2376));
    layer1_outputs(4319) <= not(layer0_outputs(1738)) or (layer0_outputs(3153));
    layer1_outputs(4320) <= not(layer0_outputs(2061)) or (layer0_outputs(4377));
    layer1_outputs(4321) <= '0';
    layer1_outputs(4322) <= not(layer0_outputs(2081));
    layer1_outputs(4323) <= not((layer0_outputs(4274)) and (layer0_outputs(1298)));
    layer1_outputs(4324) <= '0';
    layer1_outputs(4325) <= (layer0_outputs(3300)) or (layer0_outputs(2112));
    layer1_outputs(4326) <= (layer0_outputs(1141)) xor (layer0_outputs(3181));
    layer1_outputs(4327) <= not((layer0_outputs(1661)) or (layer0_outputs(4599)));
    layer1_outputs(4328) <= layer0_outputs(1869);
    layer1_outputs(4329) <= not(layer0_outputs(97));
    layer1_outputs(4330) <= not(layer0_outputs(4709));
    layer1_outputs(4331) <= not(layer0_outputs(4946));
    layer1_outputs(4332) <= (layer0_outputs(342)) and not (layer0_outputs(2042));
    layer1_outputs(4333) <= not(layer0_outputs(3369));
    layer1_outputs(4334) <= '0';
    layer1_outputs(4335) <= layer0_outputs(3122);
    layer1_outputs(4336) <= not(layer0_outputs(4517)) or (layer0_outputs(2554));
    layer1_outputs(4337) <= not((layer0_outputs(932)) or (layer0_outputs(693)));
    layer1_outputs(4338) <= not((layer0_outputs(1539)) and (layer0_outputs(1832)));
    layer1_outputs(4339) <= not(layer0_outputs(4430)) or (layer0_outputs(2595));
    layer1_outputs(4340) <= not((layer0_outputs(4493)) and (layer0_outputs(3133)));
    layer1_outputs(4341) <= (layer0_outputs(4783)) and (layer0_outputs(2393));
    layer1_outputs(4342) <= not((layer0_outputs(152)) or (layer0_outputs(1182)));
    layer1_outputs(4343) <= (layer0_outputs(4468)) or (layer0_outputs(1589));
    layer1_outputs(4344) <= not(layer0_outputs(3681)) or (layer0_outputs(2224));
    layer1_outputs(4345) <= (layer0_outputs(179)) and not (layer0_outputs(2058));
    layer1_outputs(4346) <= '1';
    layer1_outputs(4347) <= not(layer0_outputs(3346));
    layer1_outputs(4348) <= not(layer0_outputs(4305)) or (layer0_outputs(1813));
    layer1_outputs(4349) <= '1';
    layer1_outputs(4350) <= (layer0_outputs(3571)) and (layer0_outputs(1913));
    layer1_outputs(4351) <= not(layer0_outputs(4971)) or (layer0_outputs(2737));
    layer1_outputs(4352) <= '1';
    layer1_outputs(4353) <= not(layer0_outputs(1874)) or (layer0_outputs(3649));
    layer1_outputs(4354) <= '0';
    layer1_outputs(4355) <= '0';
    layer1_outputs(4356) <= layer0_outputs(935);
    layer1_outputs(4357) <= (layer0_outputs(2801)) or (layer0_outputs(3719));
    layer1_outputs(4358) <= (layer0_outputs(1256)) or (layer0_outputs(1322));
    layer1_outputs(4359) <= (layer0_outputs(3643)) and (layer0_outputs(13));
    layer1_outputs(4360) <= not(layer0_outputs(6)) or (layer0_outputs(770));
    layer1_outputs(4361) <= not((layer0_outputs(2580)) and (layer0_outputs(3351)));
    layer1_outputs(4362) <= not(layer0_outputs(2289));
    layer1_outputs(4363) <= (layer0_outputs(3477)) and not (layer0_outputs(2347));
    layer1_outputs(4364) <= not((layer0_outputs(1543)) and (layer0_outputs(4532)));
    layer1_outputs(4365) <= (layer0_outputs(326)) and (layer0_outputs(1913));
    layer1_outputs(4366) <= (layer0_outputs(2276)) and not (layer0_outputs(760));
    layer1_outputs(4367) <= '0';
    layer1_outputs(4368) <= (layer0_outputs(4816)) and not (layer0_outputs(4308));
    layer1_outputs(4369) <= '1';
    layer1_outputs(4370) <= not((layer0_outputs(2548)) or (layer0_outputs(2650)));
    layer1_outputs(4371) <= '1';
    layer1_outputs(4372) <= '0';
    layer1_outputs(4373) <= '0';
    layer1_outputs(4374) <= not(layer0_outputs(72)) or (layer0_outputs(3813));
    layer1_outputs(4375) <= not(layer0_outputs(4167));
    layer1_outputs(4376) <= '0';
    layer1_outputs(4377) <= '1';
    layer1_outputs(4378) <= '1';
    layer1_outputs(4379) <= layer0_outputs(234);
    layer1_outputs(4380) <= (layer0_outputs(1343)) or (layer0_outputs(2432));
    layer1_outputs(4381) <= '0';
    layer1_outputs(4382) <= not(layer0_outputs(683));
    layer1_outputs(4383) <= '1';
    layer1_outputs(4384) <= layer0_outputs(4390);
    layer1_outputs(4385) <= not((layer0_outputs(3650)) xor (layer0_outputs(1063)));
    layer1_outputs(4386) <= '0';
    layer1_outputs(4387) <= not(layer0_outputs(2445));
    layer1_outputs(4388) <= not((layer0_outputs(2876)) and (layer0_outputs(3171)));
    layer1_outputs(4389) <= (layer0_outputs(2914)) or (layer0_outputs(600));
    layer1_outputs(4390) <= '1';
    layer1_outputs(4391) <= not(layer0_outputs(833));
    layer1_outputs(4392) <= not((layer0_outputs(454)) or (layer0_outputs(2279)));
    layer1_outputs(4393) <= '0';
    layer1_outputs(4394) <= not((layer0_outputs(1830)) and (layer0_outputs(2475)));
    layer1_outputs(4395) <= layer0_outputs(4860);
    layer1_outputs(4396) <= (layer0_outputs(4507)) and (layer0_outputs(3689));
    layer1_outputs(4397) <= '1';
    layer1_outputs(4398) <= layer0_outputs(2010);
    layer1_outputs(4399) <= not(layer0_outputs(630));
    layer1_outputs(4400) <= not((layer0_outputs(3495)) and (layer0_outputs(109)));
    layer1_outputs(4401) <= not((layer0_outputs(3042)) or (layer0_outputs(2030)));
    layer1_outputs(4402) <= (layer0_outputs(2545)) and not (layer0_outputs(4004));
    layer1_outputs(4403) <= not(layer0_outputs(4036));
    layer1_outputs(4404) <= not((layer0_outputs(4977)) xor (layer0_outputs(4319)));
    layer1_outputs(4405) <= not(layer0_outputs(3447)) or (layer0_outputs(712));
    layer1_outputs(4406) <= not(layer0_outputs(3165)) or (layer0_outputs(4858));
    layer1_outputs(4407) <= '1';
    layer1_outputs(4408) <= not(layer0_outputs(488));
    layer1_outputs(4409) <= not(layer0_outputs(3370));
    layer1_outputs(4410) <= layer0_outputs(3270);
    layer1_outputs(4411) <= '1';
    layer1_outputs(4412) <= (layer0_outputs(1062)) or (layer0_outputs(2098));
    layer1_outputs(4413) <= not((layer0_outputs(4464)) or (layer0_outputs(3586)));
    layer1_outputs(4414) <= (layer0_outputs(1455)) and (layer0_outputs(1232));
    layer1_outputs(4415) <= (layer0_outputs(4655)) and not (layer0_outputs(171));
    layer1_outputs(4416) <= not((layer0_outputs(1957)) xor (layer0_outputs(4042)));
    layer1_outputs(4417) <= layer0_outputs(545);
    layer1_outputs(4418) <= (layer0_outputs(1029)) and (layer0_outputs(1411));
    layer1_outputs(4419) <= (layer0_outputs(309)) xor (layer0_outputs(1486));
    layer1_outputs(4420) <= (layer0_outputs(2218)) and (layer0_outputs(3279));
    layer1_outputs(4421) <= (layer0_outputs(1598)) or (layer0_outputs(85));
    layer1_outputs(4422) <= not(layer0_outputs(2510)) or (layer0_outputs(5028));
    layer1_outputs(4423) <= not((layer0_outputs(2184)) or (layer0_outputs(2423)));
    layer1_outputs(4424) <= '0';
    layer1_outputs(4425) <= layer0_outputs(4567);
    layer1_outputs(4426) <= layer0_outputs(1985);
    layer1_outputs(4427) <= layer0_outputs(155);
    layer1_outputs(4428) <= (layer0_outputs(4808)) and not (layer0_outputs(4291));
    layer1_outputs(4429) <= not(layer0_outputs(4275));
    layer1_outputs(4430) <= not(layer0_outputs(4489)) or (layer0_outputs(4845));
    layer1_outputs(4431) <= not((layer0_outputs(3223)) and (layer0_outputs(1355)));
    layer1_outputs(4432) <= layer0_outputs(1003);
    layer1_outputs(4433) <= (layer0_outputs(1007)) and not (layer0_outputs(1974));
    layer1_outputs(4434) <= not(layer0_outputs(4778));
    layer1_outputs(4435) <= '0';
    layer1_outputs(4436) <= not((layer0_outputs(2502)) and (layer0_outputs(591)));
    layer1_outputs(4437) <= layer0_outputs(3397);
    layer1_outputs(4438) <= (layer0_outputs(4979)) and not (layer0_outputs(4312));
    layer1_outputs(4439) <= '1';
    layer1_outputs(4440) <= not(layer0_outputs(4868));
    layer1_outputs(4441) <= (layer0_outputs(3635)) and not (layer0_outputs(3924));
    layer1_outputs(4442) <= not(layer0_outputs(4313)) or (layer0_outputs(3631));
    layer1_outputs(4443) <= not(layer0_outputs(788));
    layer1_outputs(4444) <= not((layer0_outputs(5095)) and (layer0_outputs(2479)));
    layer1_outputs(4445) <= (layer0_outputs(934)) or (layer0_outputs(1118));
    layer1_outputs(4446) <= not(layer0_outputs(5112)) or (layer0_outputs(5083));
    layer1_outputs(4447) <= (layer0_outputs(2630)) and (layer0_outputs(3400));
    layer1_outputs(4448) <= layer0_outputs(4439);
    layer1_outputs(4449) <= '0';
    layer1_outputs(4450) <= layer0_outputs(1310);
    layer1_outputs(4451) <= (layer0_outputs(3195)) xor (layer0_outputs(4936));
    layer1_outputs(4452) <= (layer0_outputs(3896)) and (layer0_outputs(2180));
    layer1_outputs(4453) <= not(layer0_outputs(3681)) or (layer0_outputs(1244));
    layer1_outputs(4454) <= layer0_outputs(2307);
    layer1_outputs(4455) <= layer0_outputs(3308);
    layer1_outputs(4456) <= not(layer0_outputs(1236));
    layer1_outputs(4457) <= (layer0_outputs(4706)) and not (layer0_outputs(4935));
    layer1_outputs(4458) <= not(layer0_outputs(2047)) or (layer0_outputs(1964));
    layer1_outputs(4459) <= not((layer0_outputs(3061)) or (layer0_outputs(219)));
    layer1_outputs(4460) <= '0';
    layer1_outputs(4461) <= not(layer0_outputs(749));
    layer1_outputs(4462) <= (layer0_outputs(3611)) and not (layer0_outputs(749));
    layer1_outputs(4463) <= not(layer0_outputs(2299)) or (layer0_outputs(4687));
    layer1_outputs(4464) <= layer0_outputs(4325);
    layer1_outputs(4465) <= (layer0_outputs(209)) and not (layer0_outputs(1249));
    layer1_outputs(4466) <= (layer0_outputs(4514)) or (layer0_outputs(1615));
    layer1_outputs(4467) <= layer0_outputs(1625);
    layer1_outputs(4468) <= '1';
    layer1_outputs(4469) <= (layer0_outputs(4601)) and not (layer0_outputs(1097));
    layer1_outputs(4470) <= (layer0_outputs(3713)) or (layer0_outputs(4342));
    layer1_outputs(4471) <= '1';
    layer1_outputs(4472) <= layer0_outputs(4554);
    layer1_outputs(4473) <= (layer0_outputs(2014)) and not (layer0_outputs(2285));
    layer1_outputs(4474) <= layer0_outputs(896);
    layer1_outputs(4475) <= not(layer0_outputs(3334)) or (layer0_outputs(2720));
    layer1_outputs(4476) <= not(layer0_outputs(5090));
    layer1_outputs(4477) <= layer0_outputs(1351);
    layer1_outputs(4478) <= not(layer0_outputs(1328));
    layer1_outputs(4479) <= layer0_outputs(1195);
    layer1_outputs(4480) <= not((layer0_outputs(2272)) or (layer0_outputs(4507)));
    layer1_outputs(4481) <= not(layer0_outputs(4064));
    layer1_outputs(4482) <= (layer0_outputs(301)) and (layer0_outputs(4902));
    layer1_outputs(4483) <= not((layer0_outputs(4512)) and (layer0_outputs(48)));
    layer1_outputs(4484) <= (layer0_outputs(27)) and (layer0_outputs(3327));
    layer1_outputs(4485) <= '1';
    layer1_outputs(4486) <= (layer0_outputs(3733)) and (layer0_outputs(3070));
    layer1_outputs(4487) <= layer0_outputs(2495);
    layer1_outputs(4488) <= (layer0_outputs(4622)) and not (layer0_outputs(4644));
    layer1_outputs(4489) <= (layer0_outputs(4972)) and not (layer0_outputs(2848));
    layer1_outputs(4490) <= layer0_outputs(1972);
    layer1_outputs(4491) <= (layer0_outputs(1709)) and not (layer0_outputs(4341));
    layer1_outputs(4492) <= not((layer0_outputs(172)) and (layer0_outputs(481)));
    layer1_outputs(4493) <= not(layer0_outputs(1732));
    layer1_outputs(4494) <= (layer0_outputs(733)) and not (layer0_outputs(1790));
    layer1_outputs(4495) <= (layer0_outputs(1812)) and not (layer0_outputs(4133));
    layer1_outputs(4496) <= layer0_outputs(44);
    layer1_outputs(4497) <= layer0_outputs(3112);
    layer1_outputs(4498) <= not((layer0_outputs(988)) or (layer0_outputs(3745)));
    layer1_outputs(4499) <= (layer0_outputs(581)) and (layer0_outputs(3494));
    layer1_outputs(4500) <= layer0_outputs(4905);
    layer1_outputs(4501) <= (layer0_outputs(3196)) and (layer0_outputs(4074));
    layer1_outputs(4502) <= (layer0_outputs(408)) and not (layer0_outputs(1953));
    layer1_outputs(4503) <= not(layer0_outputs(3558)) or (layer0_outputs(3216));
    layer1_outputs(4504) <= not(layer0_outputs(3243)) or (layer0_outputs(3423));
    layer1_outputs(4505) <= layer0_outputs(2863);
    layer1_outputs(4506) <= (layer0_outputs(4385)) and not (layer0_outputs(3567));
    layer1_outputs(4507) <= layer0_outputs(1466);
    layer1_outputs(4508) <= layer0_outputs(1833);
    layer1_outputs(4509) <= (layer0_outputs(1218)) or (layer0_outputs(212));
    layer1_outputs(4510) <= not(layer0_outputs(692)) or (layer0_outputs(4090));
    layer1_outputs(4511) <= layer0_outputs(1821);
    layer1_outputs(4512) <= not(layer0_outputs(354)) or (layer0_outputs(4106));
    layer1_outputs(4513) <= not(layer0_outputs(3779));
    layer1_outputs(4514) <= not(layer0_outputs(535));
    layer1_outputs(4515) <= layer0_outputs(4669);
    layer1_outputs(4516) <= not(layer0_outputs(4145)) or (layer0_outputs(127));
    layer1_outputs(4517) <= not((layer0_outputs(627)) and (layer0_outputs(1809)));
    layer1_outputs(4518) <= not(layer0_outputs(3183)) or (layer0_outputs(4101));
    layer1_outputs(4519) <= (layer0_outputs(4984)) and (layer0_outputs(458));
    layer1_outputs(4520) <= (layer0_outputs(117)) and not (layer0_outputs(4334));
    layer1_outputs(4521) <= (layer0_outputs(887)) and (layer0_outputs(3710));
    layer1_outputs(4522) <= '0';
    layer1_outputs(4523) <= not((layer0_outputs(1076)) xor (layer0_outputs(1914)));
    layer1_outputs(4524) <= not((layer0_outputs(565)) and (layer0_outputs(957)));
    layer1_outputs(4525) <= layer0_outputs(5017);
    layer1_outputs(4526) <= not(layer0_outputs(1822));
    layer1_outputs(4527) <= (layer0_outputs(4323)) and not (layer0_outputs(1604));
    layer1_outputs(4528) <= (layer0_outputs(2570)) xor (layer0_outputs(5107));
    layer1_outputs(4529) <= layer0_outputs(3093);
    layer1_outputs(4530) <= layer0_outputs(4156);
    layer1_outputs(4531) <= (layer0_outputs(1216)) or (layer0_outputs(2659));
    layer1_outputs(4532) <= (layer0_outputs(1933)) and not (layer0_outputs(2661));
    layer1_outputs(4533) <= not(layer0_outputs(56));
    layer1_outputs(4534) <= not((layer0_outputs(4641)) or (layer0_outputs(1671)));
    layer1_outputs(4535) <= not((layer0_outputs(1852)) or (layer0_outputs(85)));
    layer1_outputs(4536) <= layer0_outputs(3272);
    layer1_outputs(4537) <= not(layer0_outputs(1428));
    layer1_outputs(4538) <= (layer0_outputs(3916)) or (layer0_outputs(3140));
    layer1_outputs(4539) <= '0';
    layer1_outputs(4540) <= (layer0_outputs(2111)) and not (layer0_outputs(4384));
    layer1_outputs(4541) <= not(layer0_outputs(2220));
    layer1_outputs(4542) <= (layer0_outputs(4223)) and not (layer0_outputs(997));
    layer1_outputs(4543) <= layer0_outputs(1438);
    layer1_outputs(4544) <= not(layer0_outputs(3560));
    layer1_outputs(4545) <= (layer0_outputs(417)) and not (layer0_outputs(2806));
    layer1_outputs(4546) <= (layer0_outputs(3166)) and not (layer0_outputs(4258));
    layer1_outputs(4547) <= '0';
    layer1_outputs(4548) <= '1';
    layer1_outputs(4549) <= layer0_outputs(368);
    layer1_outputs(4550) <= (layer0_outputs(3612)) and not (layer0_outputs(2000));
    layer1_outputs(4551) <= '1';
    layer1_outputs(4552) <= '1';
    layer1_outputs(4553) <= not(layer0_outputs(476));
    layer1_outputs(4554) <= not(layer0_outputs(2053));
    layer1_outputs(4555) <= not((layer0_outputs(3849)) or (layer0_outputs(1945)));
    layer1_outputs(4556) <= not(layer0_outputs(3013));
    layer1_outputs(4557) <= layer0_outputs(1963);
    layer1_outputs(4558) <= (layer0_outputs(2037)) xor (layer0_outputs(3188));
    layer1_outputs(4559) <= not(layer0_outputs(2925)) or (layer0_outputs(907));
    layer1_outputs(4560) <= (layer0_outputs(3060)) or (layer0_outputs(700));
    layer1_outputs(4561) <= (layer0_outputs(2296)) and not (layer0_outputs(4723));
    layer1_outputs(4562) <= layer0_outputs(1787);
    layer1_outputs(4563) <= layer0_outputs(3866);
    layer1_outputs(4564) <= (layer0_outputs(759)) or (layer0_outputs(4495));
    layer1_outputs(4565) <= not(layer0_outputs(3541)) or (layer0_outputs(1382));
    layer1_outputs(4566) <= not(layer0_outputs(1676)) or (layer0_outputs(5053));
    layer1_outputs(4567) <= '0';
    layer1_outputs(4568) <= not((layer0_outputs(1475)) and (layer0_outputs(407)));
    layer1_outputs(4569) <= not((layer0_outputs(3076)) xor (layer0_outputs(4738)));
    layer1_outputs(4570) <= not((layer0_outputs(1278)) or (layer0_outputs(490)));
    layer1_outputs(4571) <= (layer0_outputs(613)) and not (layer0_outputs(669));
    layer1_outputs(4572) <= (layer0_outputs(1177)) and not (layer0_outputs(1137));
    layer1_outputs(4573) <= not(layer0_outputs(696)) or (layer0_outputs(2282));
    layer1_outputs(4574) <= '0';
    layer1_outputs(4575) <= (layer0_outputs(4184)) and not (layer0_outputs(1998));
    layer1_outputs(4576) <= not((layer0_outputs(5082)) or (layer0_outputs(2485)));
    layer1_outputs(4577) <= not((layer0_outputs(1126)) xor (layer0_outputs(3209)));
    layer1_outputs(4578) <= not(layer0_outputs(4159));
    layer1_outputs(4579) <= '1';
    layer1_outputs(4580) <= not((layer0_outputs(3159)) or (layer0_outputs(2374)));
    layer1_outputs(4581) <= (layer0_outputs(1164)) and not (layer0_outputs(1400));
    layer1_outputs(4582) <= not(layer0_outputs(4658)) or (layer0_outputs(2421));
    layer1_outputs(4583) <= not(layer0_outputs(1688));
    layer1_outputs(4584) <= not(layer0_outputs(751)) or (layer0_outputs(3619));
    layer1_outputs(4585) <= not(layer0_outputs(2408));
    layer1_outputs(4586) <= not(layer0_outputs(2895)) or (layer0_outputs(4864));
    layer1_outputs(4587) <= not(layer0_outputs(1845));
    layer1_outputs(4588) <= not(layer0_outputs(3705));
    layer1_outputs(4589) <= not(layer0_outputs(2378)) or (layer0_outputs(2752));
    layer1_outputs(4590) <= not(layer0_outputs(158));
    layer1_outputs(4591) <= (layer0_outputs(5105)) and not (layer0_outputs(3762));
    layer1_outputs(4592) <= not(layer0_outputs(2337)) or (layer0_outputs(74));
    layer1_outputs(4593) <= '1';
    layer1_outputs(4594) <= layer0_outputs(5016);
    layer1_outputs(4595) <= layer0_outputs(4895);
    layer1_outputs(4596) <= not((layer0_outputs(3855)) and (layer0_outputs(2835)));
    layer1_outputs(4597) <= (layer0_outputs(4639)) or (layer0_outputs(1541));
    layer1_outputs(4598) <= '0';
    layer1_outputs(4599) <= (layer0_outputs(2701)) or (layer0_outputs(461));
    layer1_outputs(4600) <= not(layer0_outputs(1545));
    layer1_outputs(4601) <= not(layer0_outputs(2716)) or (layer0_outputs(589));
    layer1_outputs(4602) <= not(layer0_outputs(4763));
    layer1_outputs(4603) <= not(layer0_outputs(1872)) or (layer0_outputs(3224));
    layer1_outputs(4604) <= (layer0_outputs(3945)) and (layer0_outputs(675));
    layer1_outputs(4605) <= layer0_outputs(513);
    layer1_outputs(4606) <= '0';
    layer1_outputs(4607) <= (layer0_outputs(1000)) or (layer0_outputs(4831));
    layer1_outputs(4608) <= layer0_outputs(4198);
    layer1_outputs(4609) <= not(layer0_outputs(3084)) or (layer0_outputs(3514));
    layer1_outputs(4610) <= not(layer0_outputs(1173));
    layer1_outputs(4611) <= not(layer0_outputs(3350)) or (layer0_outputs(518));
    layer1_outputs(4612) <= (layer0_outputs(4125)) and (layer0_outputs(3107));
    layer1_outputs(4613) <= (layer0_outputs(4213)) and (layer0_outputs(3639));
    layer1_outputs(4614) <= not(layer0_outputs(2065));
    layer1_outputs(4615) <= not((layer0_outputs(4700)) or (layer0_outputs(798)));
    layer1_outputs(4616) <= not(layer0_outputs(2939));
    layer1_outputs(4617) <= (layer0_outputs(3712)) and not (layer0_outputs(966));
    layer1_outputs(4618) <= '1';
    layer1_outputs(4619) <= layer0_outputs(100);
    layer1_outputs(4620) <= not(layer0_outputs(2110)) or (layer0_outputs(3529));
    layer1_outputs(4621) <= not((layer0_outputs(3014)) and (layer0_outputs(328)));
    layer1_outputs(4622) <= layer0_outputs(2213);
    layer1_outputs(4623) <= not(layer0_outputs(2452)) or (layer0_outputs(4256));
    layer1_outputs(4624) <= not(layer0_outputs(1133)) or (layer0_outputs(4651));
    layer1_outputs(4625) <= not((layer0_outputs(2870)) or (layer0_outputs(3407)));
    layer1_outputs(4626) <= (layer0_outputs(3087)) or (layer0_outputs(3606));
    layer1_outputs(4627) <= layer0_outputs(1950);
    layer1_outputs(4628) <= (layer0_outputs(4063)) and not (layer0_outputs(3119));
    layer1_outputs(4629) <= not(layer0_outputs(2871)) or (layer0_outputs(589));
    layer1_outputs(4630) <= '0';
    layer1_outputs(4631) <= not(layer0_outputs(5027));
    layer1_outputs(4632) <= (layer0_outputs(1503)) and not (layer0_outputs(2322));
    layer1_outputs(4633) <= not(layer0_outputs(99)) or (layer0_outputs(3725));
    layer1_outputs(4634) <= (layer0_outputs(3972)) and not (layer0_outputs(2517));
    layer1_outputs(4635) <= layer0_outputs(1359);
    layer1_outputs(4636) <= (layer0_outputs(4776)) and not (layer0_outputs(1357));
    layer1_outputs(4637) <= (layer0_outputs(4343)) and (layer0_outputs(5031));
    layer1_outputs(4638) <= not(layer0_outputs(2405));
    layer1_outputs(4639) <= (layer0_outputs(951)) and not (layer0_outputs(2443));
    layer1_outputs(4640) <= (layer0_outputs(4842)) and not (layer0_outputs(214));
    layer1_outputs(4641) <= not(layer0_outputs(4171)) or (layer0_outputs(2149));
    layer1_outputs(4642) <= (layer0_outputs(2275)) or (layer0_outputs(3072));
    layer1_outputs(4643) <= not(layer0_outputs(2785)) or (layer0_outputs(3953));
    layer1_outputs(4644) <= (layer0_outputs(1023)) and not (layer0_outputs(3755));
    layer1_outputs(4645) <= not(layer0_outputs(1379));
    layer1_outputs(4646) <= not(layer0_outputs(1356));
    layer1_outputs(4647) <= (layer0_outputs(1859)) and not (layer0_outputs(3522));
    layer1_outputs(4648) <= (layer0_outputs(582)) and (layer0_outputs(877));
    layer1_outputs(4649) <= (layer0_outputs(4981)) and not (layer0_outputs(2079));
    layer1_outputs(4650) <= (layer0_outputs(1273)) and not (layer0_outputs(358));
    layer1_outputs(4651) <= not((layer0_outputs(2227)) or (layer0_outputs(911)));
    layer1_outputs(4652) <= (layer0_outputs(4317)) and (layer0_outputs(4851));
    layer1_outputs(4653) <= not(layer0_outputs(116));
    layer1_outputs(4654) <= (layer0_outputs(3178)) or (layer0_outputs(3397));
    layer1_outputs(4655) <= not((layer0_outputs(2343)) xor (layer0_outputs(800)));
    layer1_outputs(4656) <= not((layer0_outputs(555)) and (layer0_outputs(4456)));
    layer1_outputs(4657) <= not((layer0_outputs(4380)) and (layer0_outputs(4120)));
    layer1_outputs(4658) <= not(layer0_outputs(4179)) or (layer0_outputs(1916));
    layer1_outputs(4659) <= '0';
    layer1_outputs(4660) <= not((layer0_outputs(3169)) or (layer0_outputs(151)));
    layer1_outputs(4661) <= (layer0_outputs(4703)) and (layer0_outputs(568));
    layer1_outputs(4662) <= layer0_outputs(668);
    layer1_outputs(4663) <= (layer0_outputs(2627)) and (layer0_outputs(4420));
    layer1_outputs(4664) <= layer0_outputs(3997);
    layer1_outputs(4665) <= not(layer0_outputs(1929)) or (layer0_outputs(3170));
    layer1_outputs(4666) <= (layer0_outputs(3871)) or (layer0_outputs(2034));
    layer1_outputs(4667) <= layer0_outputs(104);
    layer1_outputs(4668) <= '1';
    layer1_outputs(4669) <= not(layer0_outputs(3505)) or (layer0_outputs(2758));
    layer1_outputs(4670) <= '0';
    layer1_outputs(4671) <= (layer0_outputs(1424)) or (layer0_outputs(4847));
    layer1_outputs(4672) <= (layer0_outputs(181)) and not (layer0_outputs(3886));
    layer1_outputs(4673) <= not(layer0_outputs(763));
    layer1_outputs(4674) <= layer0_outputs(4430);
    layer1_outputs(4675) <= not(layer0_outputs(2141)) or (layer0_outputs(4425));
    layer1_outputs(4676) <= not(layer0_outputs(4109));
    layer1_outputs(4677) <= (layer0_outputs(5024)) or (layer0_outputs(5064));
    layer1_outputs(4678) <= '1';
    layer1_outputs(4679) <= (layer0_outputs(1924)) and not (layer0_outputs(3654));
    layer1_outputs(4680) <= '0';
    layer1_outputs(4681) <= not((layer0_outputs(2783)) and (layer0_outputs(2309)));
    layer1_outputs(4682) <= (layer0_outputs(3779)) and not (layer0_outputs(1459));
    layer1_outputs(4683) <= (layer0_outputs(2689)) or (layer0_outputs(3541));
    layer1_outputs(4684) <= (layer0_outputs(4857)) and not (layer0_outputs(2921));
    layer1_outputs(4685) <= not(layer0_outputs(3526));
    layer1_outputs(4686) <= not((layer0_outputs(1285)) and (layer0_outputs(3083)));
    layer1_outputs(4687) <= not(layer0_outputs(1488)) or (layer0_outputs(1661));
    layer1_outputs(4688) <= layer0_outputs(3874);
    layer1_outputs(4689) <= not(layer0_outputs(4477)) or (layer0_outputs(3072));
    layer1_outputs(4690) <= not(layer0_outputs(2277)) or (layer0_outputs(3017));
    layer1_outputs(4691) <= (layer0_outputs(3695)) and not (layer0_outputs(3312));
    layer1_outputs(4692) <= layer0_outputs(3314);
    layer1_outputs(4693) <= (layer0_outputs(691)) and not (layer0_outputs(1530));
    layer1_outputs(4694) <= not(layer0_outputs(4093));
    layer1_outputs(4695) <= not(layer0_outputs(2723));
    layer1_outputs(4696) <= '1';
    layer1_outputs(4697) <= '1';
    layer1_outputs(4698) <= layer0_outputs(1493);
    layer1_outputs(4699) <= '0';
    layer1_outputs(4700) <= layer0_outputs(3153);
    layer1_outputs(4701) <= '0';
    layer1_outputs(4702) <= not((layer0_outputs(2766)) and (layer0_outputs(3585)));
    layer1_outputs(4703) <= layer0_outputs(3628);
    layer1_outputs(4704) <= not((layer0_outputs(1172)) or (layer0_outputs(4341)));
    layer1_outputs(4705) <= (layer0_outputs(4307)) and not (layer0_outputs(3653));
    layer1_outputs(4706) <= '0';
    layer1_outputs(4707) <= layer0_outputs(3027);
    layer1_outputs(4708) <= (layer0_outputs(3823)) and (layer0_outputs(175));
    layer1_outputs(4709) <= '1';
    layer1_outputs(4710) <= not((layer0_outputs(786)) and (layer0_outputs(1308)));
    layer1_outputs(4711) <= not(layer0_outputs(2611));
    layer1_outputs(4712) <= not(layer0_outputs(2561)) or (layer0_outputs(1938));
    layer1_outputs(4713) <= not(layer0_outputs(3218)) or (layer0_outputs(1358));
    layer1_outputs(4714) <= '1';
    layer1_outputs(4715) <= layer0_outputs(5077);
    layer1_outputs(4716) <= '1';
    layer1_outputs(4717) <= not(layer0_outputs(1525)) or (layer0_outputs(638));
    layer1_outputs(4718) <= not(layer0_outputs(44));
    layer1_outputs(4719) <= (layer0_outputs(4769)) and (layer0_outputs(3235));
    layer1_outputs(4720) <= '0';
    layer1_outputs(4721) <= (layer0_outputs(4393)) and not (layer0_outputs(2339));
    layer1_outputs(4722) <= (layer0_outputs(3006)) and not (layer0_outputs(3470));
    layer1_outputs(4723) <= not((layer0_outputs(1403)) or (layer0_outputs(1677)));
    layer1_outputs(4724) <= not((layer0_outputs(2289)) and (layer0_outputs(1449)));
    layer1_outputs(4725) <= not((layer0_outputs(2402)) xor (layer0_outputs(4790)));
    layer1_outputs(4726) <= not(layer0_outputs(4828));
    layer1_outputs(4727) <= not(layer0_outputs(4071));
    layer1_outputs(4728) <= not((layer0_outputs(4508)) or (layer0_outputs(4805)));
    layer1_outputs(4729) <= '1';
    layer1_outputs(4730) <= layer0_outputs(1092);
    layer1_outputs(4731) <= layer0_outputs(4547);
    layer1_outputs(4732) <= layer0_outputs(4458);
    layer1_outputs(4733) <= layer0_outputs(416);
    layer1_outputs(4734) <= (layer0_outputs(1816)) and not (layer0_outputs(5043));
    layer1_outputs(4735) <= not(layer0_outputs(2489));
    layer1_outputs(4736) <= not(layer0_outputs(1504)) or (layer0_outputs(480));
    layer1_outputs(4737) <= layer0_outputs(2003);
    layer1_outputs(4738) <= (layer0_outputs(1758)) xor (layer0_outputs(1654));
    layer1_outputs(4739) <= not(layer0_outputs(656));
    layer1_outputs(4740) <= not(layer0_outputs(1917));
    layer1_outputs(4741) <= (layer0_outputs(3012)) and not (layer0_outputs(1366));
    layer1_outputs(4742) <= (layer0_outputs(2658)) or (layer0_outputs(1193));
    layer1_outputs(4743) <= not(layer0_outputs(4686));
    layer1_outputs(4744) <= '0';
    layer1_outputs(4745) <= (layer0_outputs(4832)) and not (layer0_outputs(2957));
    layer1_outputs(4746) <= layer0_outputs(162);
    layer1_outputs(4747) <= layer0_outputs(3229);
    layer1_outputs(4748) <= not(layer0_outputs(2301));
    layer1_outputs(4749) <= not(layer0_outputs(3337)) or (layer0_outputs(4106));
    layer1_outputs(4750) <= not(layer0_outputs(3000)) or (layer0_outputs(387));
    layer1_outputs(4751) <= not((layer0_outputs(1829)) or (layer0_outputs(4245)));
    layer1_outputs(4752) <= not((layer0_outputs(211)) or (layer0_outputs(2705)));
    layer1_outputs(4753) <= '0';
    layer1_outputs(4754) <= (layer0_outputs(2635)) xor (layer0_outputs(2842));
    layer1_outputs(4755) <= not(layer0_outputs(424));
    layer1_outputs(4756) <= '1';
    layer1_outputs(4757) <= '1';
    layer1_outputs(4758) <= (layer0_outputs(3405)) and (layer0_outputs(3836));
    layer1_outputs(4759) <= layer0_outputs(811);
    layer1_outputs(4760) <= layer0_outputs(4766);
    layer1_outputs(4761) <= layer0_outputs(4673);
    layer1_outputs(4762) <= '0';
    layer1_outputs(4763) <= not(layer0_outputs(1555)) or (layer0_outputs(570));
    layer1_outputs(4764) <= layer0_outputs(1881);
    layer1_outputs(4765) <= layer0_outputs(1726);
    layer1_outputs(4766) <= not(layer0_outputs(1158));
    layer1_outputs(4767) <= not(layer0_outputs(622)) or (layer0_outputs(3131));
    layer1_outputs(4768) <= layer0_outputs(190);
    layer1_outputs(4769) <= '1';
    layer1_outputs(4770) <= not((layer0_outputs(3438)) and (layer0_outputs(1089)));
    layer1_outputs(4771) <= (layer0_outputs(3291)) and (layer0_outputs(4084));
    layer1_outputs(4772) <= not(layer0_outputs(108));
    layer1_outputs(4773) <= not(layer0_outputs(3152));
    layer1_outputs(4774) <= layer0_outputs(4353);
    layer1_outputs(4775) <= not((layer0_outputs(1988)) or (layer0_outputs(2072)));
    layer1_outputs(4776) <= layer0_outputs(702);
    layer1_outputs(4777) <= not((layer0_outputs(4163)) or (layer0_outputs(254)));
    layer1_outputs(4778) <= '1';
    layer1_outputs(4779) <= '0';
    layer1_outputs(4780) <= not((layer0_outputs(4782)) or (layer0_outputs(2257)));
    layer1_outputs(4781) <= (layer0_outputs(989)) and (layer0_outputs(3577));
    layer1_outputs(4782) <= not(layer0_outputs(995));
    layer1_outputs(4783) <= not((layer0_outputs(4586)) or (layer0_outputs(1368)));
    layer1_outputs(4784) <= not(layer0_outputs(2602));
    layer1_outputs(4785) <= not(layer0_outputs(1312));
    layer1_outputs(4786) <= not(layer0_outputs(3638));
    layer1_outputs(4787) <= '1';
    layer1_outputs(4788) <= not((layer0_outputs(4180)) xor (layer0_outputs(1303)));
    layer1_outputs(4789) <= '0';
    layer1_outputs(4790) <= not((layer0_outputs(2328)) or (layer0_outputs(1011)));
    layer1_outputs(4791) <= not(layer0_outputs(2057)) or (layer0_outputs(3382));
    layer1_outputs(4792) <= (layer0_outputs(1016)) or (layer0_outputs(3356));
    layer1_outputs(4793) <= (layer0_outputs(1228)) and (layer0_outputs(1847));
    layer1_outputs(4794) <= not(layer0_outputs(335)) or (layer0_outputs(860));
    layer1_outputs(4795) <= (layer0_outputs(3461)) and not (layer0_outputs(4370));
    layer1_outputs(4796) <= not(layer0_outputs(4236)) or (layer0_outputs(3804));
    layer1_outputs(4797) <= '0';
    layer1_outputs(4798) <= not(layer0_outputs(1642)) or (layer0_outputs(3846));
    layer1_outputs(4799) <= '0';
    layer1_outputs(4800) <= not(layer0_outputs(2203)) or (layer0_outputs(1481));
    layer1_outputs(4801) <= not(layer0_outputs(4335));
    layer1_outputs(4802) <= '1';
    layer1_outputs(4803) <= '0';
    layer1_outputs(4804) <= '1';
    layer1_outputs(4805) <= layer0_outputs(4391);
    layer1_outputs(4806) <= not(layer0_outputs(339));
    layer1_outputs(4807) <= '1';
    layer1_outputs(4808) <= not(layer0_outputs(4501)) or (layer0_outputs(4523));
    layer1_outputs(4809) <= (layer0_outputs(2914)) and not (layer0_outputs(4821));
    layer1_outputs(4810) <= not(layer0_outputs(3203)) or (layer0_outputs(2867));
    layer1_outputs(4811) <= '1';
    layer1_outputs(4812) <= layer0_outputs(3578);
    layer1_outputs(4813) <= layer0_outputs(1085);
    layer1_outputs(4814) <= '1';
    layer1_outputs(4815) <= not(layer0_outputs(3052));
    layer1_outputs(4816) <= (layer0_outputs(4655)) xor (layer0_outputs(2832));
    layer1_outputs(4817) <= '1';
    layer1_outputs(4818) <= not((layer0_outputs(1965)) and (layer0_outputs(3937)));
    layer1_outputs(4819) <= not(layer0_outputs(4415));
    layer1_outputs(4820) <= not((layer0_outputs(3527)) or (layer0_outputs(3674)));
    layer1_outputs(4821) <= '0';
    layer1_outputs(4822) <= '0';
    layer1_outputs(4823) <= not(layer0_outputs(4040));
    layer1_outputs(4824) <= layer0_outputs(5013);
    layer1_outputs(4825) <= not(layer0_outputs(2087)) or (layer0_outputs(3301));
    layer1_outputs(4826) <= (layer0_outputs(149)) and not (layer0_outputs(1803));
    layer1_outputs(4827) <= layer0_outputs(1600);
    layer1_outputs(4828) <= (layer0_outputs(236)) or (layer0_outputs(969));
    layer1_outputs(4829) <= (layer0_outputs(31)) and (layer0_outputs(4487));
    layer1_outputs(4830) <= not((layer0_outputs(959)) or (layer0_outputs(2135)));
    layer1_outputs(4831) <= layer0_outputs(2068);
    layer1_outputs(4832) <= '0';
    layer1_outputs(4833) <= (layer0_outputs(1252)) and (layer0_outputs(1060));
    layer1_outputs(4834) <= (layer0_outputs(2895)) and (layer0_outputs(328));
    layer1_outputs(4835) <= (layer0_outputs(1157)) and (layer0_outputs(1781));
    layer1_outputs(4836) <= (layer0_outputs(3402)) or (layer0_outputs(3671));
    layer1_outputs(4837) <= not(layer0_outputs(724));
    layer1_outputs(4838) <= (layer0_outputs(807)) and not (layer0_outputs(2277));
    layer1_outputs(4839) <= '0';
    layer1_outputs(4840) <= layer0_outputs(2249);
    layer1_outputs(4841) <= '0';
    layer1_outputs(4842) <= layer0_outputs(3853);
    layer1_outputs(4843) <= layer0_outputs(2703);
    layer1_outputs(4844) <= (layer0_outputs(4541)) and (layer0_outputs(3329));
    layer1_outputs(4845) <= layer0_outputs(2762);
    layer1_outputs(4846) <= not(layer0_outputs(585));
    layer1_outputs(4847) <= layer0_outputs(1440);
    layer1_outputs(4848) <= '0';
    layer1_outputs(4849) <= not((layer0_outputs(1978)) or (layer0_outputs(3766)));
    layer1_outputs(4850) <= '0';
    layer1_outputs(4851) <= layer0_outputs(3921);
    layer1_outputs(4852) <= not(layer0_outputs(4985)) or (layer0_outputs(3818));
    layer1_outputs(4853) <= not((layer0_outputs(4795)) or (layer0_outputs(4175)));
    layer1_outputs(4854) <= '1';
    layer1_outputs(4855) <= not(layer0_outputs(1944)) or (layer0_outputs(3496));
    layer1_outputs(4856) <= not(layer0_outputs(3608)) or (layer0_outputs(2907));
    layer1_outputs(4857) <= (layer0_outputs(3036)) and not (layer0_outputs(4988));
    layer1_outputs(4858) <= not(layer0_outputs(4174));
    layer1_outputs(4859) <= '1';
    layer1_outputs(4860) <= not(layer0_outputs(2428)) or (layer0_outputs(3015));
    layer1_outputs(4861) <= not((layer0_outputs(4116)) or (layer0_outputs(3835)));
    layer1_outputs(4862) <= (layer0_outputs(2585)) or (layer0_outputs(4927));
    layer1_outputs(4863) <= (layer0_outputs(3627)) and not (layer0_outputs(3512));
    layer1_outputs(4864) <= (layer0_outputs(4156)) and not (layer0_outputs(2901));
    layer1_outputs(4865) <= (layer0_outputs(4661)) or (layer0_outputs(4197));
    layer1_outputs(4866) <= not(layer0_outputs(3942)) or (layer0_outputs(124));
    layer1_outputs(4867) <= not(layer0_outputs(2636)) or (layer0_outputs(657));
    layer1_outputs(4868) <= not(layer0_outputs(1707));
    layer1_outputs(4869) <= not((layer0_outputs(1143)) and (layer0_outputs(4363)));
    layer1_outputs(4870) <= '0';
    layer1_outputs(4871) <= '0';
    layer1_outputs(4872) <= not(layer0_outputs(4132)) or (layer0_outputs(603));
    layer1_outputs(4873) <= '0';
    layer1_outputs(4874) <= not(layer0_outputs(4674));
    layer1_outputs(4875) <= not(layer0_outputs(1475));
    layer1_outputs(4876) <= not(layer0_outputs(4688));
    layer1_outputs(4877) <= (layer0_outputs(500)) xor (layer0_outputs(1474));
    layer1_outputs(4878) <= not(layer0_outputs(813)) or (layer0_outputs(4381));
    layer1_outputs(4879) <= not(layer0_outputs(1923));
    layer1_outputs(4880) <= not((layer0_outputs(1823)) xor (layer0_outputs(2769)));
    layer1_outputs(4881) <= (layer0_outputs(1700)) and not (layer0_outputs(724));
    layer1_outputs(4882) <= (layer0_outputs(3222)) and (layer0_outputs(1587));
    layer1_outputs(4883) <= layer0_outputs(4480);
    layer1_outputs(4884) <= not((layer0_outputs(3341)) or (layer0_outputs(2040)));
    layer1_outputs(4885) <= (layer0_outputs(2460)) and (layer0_outputs(1955));
    layer1_outputs(4886) <= not(layer0_outputs(1276)) or (layer0_outputs(4531));
    layer1_outputs(4887) <= (layer0_outputs(36)) and (layer0_outputs(1199));
    layer1_outputs(4888) <= '0';
    layer1_outputs(4889) <= layer0_outputs(5074);
    layer1_outputs(4890) <= '1';
    layer1_outputs(4891) <= '0';
    layer1_outputs(4892) <= '0';
    layer1_outputs(4893) <= not(layer0_outputs(1058)) or (layer0_outputs(667));
    layer1_outputs(4894) <= (layer0_outputs(5038)) and not (layer0_outputs(2571));
    layer1_outputs(4895) <= layer0_outputs(4280);
    layer1_outputs(4896) <= (layer0_outputs(915)) and not (layer0_outputs(2285));
    layer1_outputs(4897) <= not(layer0_outputs(1203));
    layer1_outputs(4898) <= not(layer0_outputs(3575)) or (layer0_outputs(1591));
    layer1_outputs(4899) <= not(layer0_outputs(3579));
    layer1_outputs(4900) <= layer0_outputs(995);
    layer1_outputs(4901) <= not(layer0_outputs(4400)) or (layer0_outputs(3460));
    layer1_outputs(4902) <= not(layer0_outputs(3645)) or (layer0_outputs(4970));
    layer1_outputs(4903) <= (layer0_outputs(1175)) and not (layer0_outputs(2656));
    layer1_outputs(4904) <= not(layer0_outputs(484));
    layer1_outputs(4905) <= '0';
    layer1_outputs(4906) <= layer0_outputs(1329);
    layer1_outputs(4907) <= '1';
    layer1_outputs(4908) <= (layer0_outputs(2615)) and (layer0_outputs(3154));
    layer1_outputs(4909) <= not(layer0_outputs(773));
    layer1_outputs(4910) <= not(layer0_outputs(1804)) or (layer0_outputs(5028));
    layer1_outputs(4911) <= '1';
    layer1_outputs(4912) <= not(layer0_outputs(3508));
    layer1_outputs(4913) <= (layer0_outputs(201)) and not (layer0_outputs(1811));
    layer1_outputs(4914) <= not((layer0_outputs(3133)) and (layer0_outputs(1871)));
    layer1_outputs(4915) <= not(layer0_outputs(1292)) or (layer0_outputs(2077));
    layer1_outputs(4916) <= not(layer0_outputs(1579)) or (layer0_outputs(2193));
    layer1_outputs(4917) <= (layer0_outputs(4904)) and not (layer0_outputs(636));
    layer1_outputs(4918) <= not(layer0_outputs(4012)) or (layer0_outputs(2851));
    layer1_outputs(4919) <= not(layer0_outputs(2674)) or (layer0_outputs(1679));
    layer1_outputs(4920) <= not((layer0_outputs(1179)) xor (layer0_outputs(3913)));
    layer1_outputs(4921) <= not(layer0_outputs(2102)) or (layer0_outputs(3062));
    layer1_outputs(4922) <= layer0_outputs(4586);
    layer1_outputs(4923) <= (layer0_outputs(1829)) xor (layer0_outputs(1407));
    layer1_outputs(4924) <= layer0_outputs(1862);
    layer1_outputs(4925) <= not(layer0_outputs(2988));
    layer1_outputs(4926) <= not(layer0_outputs(2181)) or (layer0_outputs(1980));
    layer1_outputs(4927) <= not(layer0_outputs(3800));
    layer1_outputs(4928) <= '0';
    layer1_outputs(4929) <= '0';
    layer1_outputs(4930) <= not(layer0_outputs(1261));
    layer1_outputs(4931) <= not((layer0_outputs(3529)) or (layer0_outputs(3870)));
    layer1_outputs(4932) <= not(layer0_outputs(1840));
    layer1_outputs(4933) <= (layer0_outputs(531)) and (layer0_outputs(5106));
    layer1_outputs(4934) <= not((layer0_outputs(3366)) or (layer0_outputs(2541)));
    layer1_outputs(4935) <= not(layer0_outputs(4891));
    layer1_outputs(4936) <= '0';
    layer1_outputs(4937) <= (layer0_outputs(2900)) or (layer0_outputs(2665));
    layer1_outputs(4938) <= '0';
    layer1_outputs(4939) <= (layer0_outputs(4800)) and not (layer0_outputs(918));
    layer1_outputs(4940) <= not(layer0_outputs(3383));
    layer1_outputs(4941) <= not((layer0_outputs(1211)) or (layer0_outputs(3656)));
    layer1_outputs(4942) <= layer0_outputs(3555);
    layer1_outputs(4943) <= '0';
    layer1_outputs(4944) <= not(layer0_outputs(2961)) or (layer0_outputs(2625));
    layer1_outputs(4945) <= not((layer0_outputs(2579)) xor (layer0_outputs(4121)));
    layer1_outputs(4946) <= (layer0_outputs(4844)) xor (layer0_outputs(864));
    layer1_outputs(4947) <= (layer0_outputs(2368)) or (layer0_outputs(188));
    layer1_outputs(4948) <= layer0_outputs(4704);
    layer1_outputs(4949) <= not(layer0_outputs(521));
    layer1_outputs(4950) <= not((layer0_outputs(4713)) and (layer0_outputs(503)));
    layer1_outputs(4951) <= not(layer0_outputs(2104)) or (layer0_outputs(4654));
    layer1_outputs(4952) <= not(layer0_outputs(2727)) or (layer0_outputs(4472));
    layer1_outputs(4953) <= not((layer0_outputs(5013)) or (layer0_outputs(1808)));
    layer1_outputs(4954) <= (layer0_outputs(2384)) xor (layer0_outputs(3076));
    layer1_outputs(4955) <= not(layer0_outputs(1551)) or (layer0_outputs(629));
    layer1_outputs(4956) <= layer0_outputs(2162);
    layer1_outputs(4957) <= not(layer0_outputs(67));
    layer1_outputs(4958) <= '0';
    layer1_outputs(4959) <= layer0_outputs(5029);
    layer1_outputs(4960) <= (layer0_outputs(3361)) or (layer0_outputs(336));
    layer1_outputs(4961) <= (layer0_outputs(2243)) and not (layer0_outputs(908));
    layer1_outputs(4962) <= not(layer0_outputs(2782));
    layer1_outputs(4963) <= not((layer0_outputs(2194)) and (layer0_outputs(295)));
    layer1_outputs(4964) <= (layer0_outputs(1993)) and not (layer0_outputs(489));
    layer1_outputs(4965) <= layer0_outputs(3727);
    layer1_outputs(4966) <= (layer0_outputs(1356)) and (layer0_outputs(3286));
    layer1_outputs(4967) <= (layer0_outputs(4303)) and not (layer0_outputs(2773));
    layer1_outputs(4968) <= '1';
    layer1_outputs(4969) <= layer0_outputs(1274);
    layer1_outputs(4970) <= '1';
    layer1_outputs(4971) <= layer0_outputs(4187);
    layer1_outputs(4972) <= (layer0_outputs(1)) and not (layer0_outputs(14));
    layer1_outputs(4973) <= not((layer0_outputs(2235)) or (layer0_outputs(2447)));
    layer1_outputs(4974) <= not((layer0_outputs(1976)) and (layer0_outputs(1031)));
    layer1_outputs(4975) <= layer0_outputs(1277);
    layer1_outputs(4976) <= not((layer0_outputs(92)) and (layer0_outputs(2425)));
    layer1_outputs(4977) <= not(layer0_outputs(5042)) or (layer0_outputs(3191));
    layer1_outputs(4978) <= '1';
    layer1_outputs(4979) <= '1';
    layer1_outputs(4980) <= '1';
    layer1_outputs(4981) <= '1';
    layer1_outputs(4982) <= layer0_outputs(785);
    layer1_outputs(4983) <= not(layer0_outputs(1611));
    layer1_outputs(4984) <= layer0_outputs(2854);
    layer1_outputs(4985) <= not(layer0_outputs(1631));
    layer1_outputs(4986) <= '1';
    layer1_outputs(4987) <= not(layer0_outputs(128)) or (layer0_outputs(2511));
    layer1_outputs(4988) <= layer0_outputs(1142);
    layer1_outputs(4989) <= not(layer0_outputs(1894)) or (layer0_outputs(4533));
    layer1_outputs(4990) <= not(layer0_outputs(4945));
    layer1_outputs(4991) <= not((layer0_outputs(963)) xor (layer0_outputs(4269)));
    layer1_outputs(4992) <= not(layer0_outputs(2662)) or (layer0_outputs(2654));
    layer1_outputs(4993) <= not((layer0_outputs(4204)) or (layer0_outputs(2487)));
    layer1_outputs(4994) <= '1';
    layer1_outputs(4995) <= not(layer0_outputs(4218));
    layer1_outputs(4996) <= not(layer0_outputs(3689));
    layer1_outputs(4997) <= '0';
    layer1_outputs(4998) <= not(layer0_outputs(555)) or (layer0_outputs(2280));
    layer1_outputs(4999) <= (layer0_outputs(1337)) and not (layer0_outputs(2496));
    layer1_outputs(5000) <= layer0_outputs(4442);
    layer1_outputs(5001) <= (layer0_outputs(4253)) and (layer0_outputs(16));
    layer1_outputs(5002) <= not((layer0_outputs(4041)) and (layer0_outputs(2999)));
    layer1_outputs(5003) <= not((layer0_outputs(1408)) and (layer0_outputs(4200)));
    layer1_outputs(5004) <= '0';
    layer1_outputs(5005) <= (layer0_outputs(437)) and (layer0_outputs(3166));
    layer1_outputs(5006) <= not(layer0_outputs(4910)) or (layer0_outputs(2397));
    layer1_outputs(5007) <= not((layer0_outputs(3388)) and (layer0_outputs(3071)));
    layer1_outputs(5008) <= '0';
    layer1_outputs(5009) <= layer0_outputs(4881);
    layer1_outputs(5010) <= layer0_outputs(1138);
    layer1_outputs(5011) <= not(layer0_outputs(3257)) or (layer0_outputs(415));
    layer1_outputs(5012) <= layer0_outputs(4249);
    layer1_outputs(5013) <= layer0_outputs(1059);
    layer1_outputs(5014) <= (layer0_outputs(2784)) or (layer0_outputs(3763));
    layer1_outputs(5015) <= not(layer0_outputs(93)) or (layer0_outputs(2739));
    layer1_outputs(5016) <= layer0_outputs(678);
    layer1_outputs(5017) <= (layer0_outputs(5116)) and (layer0_outputs(1633));
    layer1_outputs(5018) <= not(layer0_outputs(1845)) or (layer0_outputs(3944));
    layer1_outputs(5019) <= (layer0_outputs(2167)) and (layer0_outputs(2615));
    layer1_outputs(5020) <= (layer0_outputs(748)) and not (layer0_outputs(2442));
    layer1_outputs(5021) <= not(layer0_outputs(2743)) or (layer0_outputs(4809));
    layer1_outputs(5022) <= not((layer0_outputs(289)) and (layer0_outputs(442)));
    layer1_outputs(5023) <= not(layer0_outputs(2009));
    layer1_outputs(5024) <= layer0_outputs(1346);
    layer1_outputs(5025) <= layer0_outputs(3270);
    layer1_outputs(5026) <= '0';
    layer1_outputs(5027) <= layer0_outputs(1853);
    layer1_outputs(5028) <= not(layer0_outputs(1977)) or (layer0_outputs(2403));
    layer1_outputs(5029) <= not((layer0_outputs(1152)) or (layer0_outputs(3547)));
    layer1_outputs(5030) <= not(layer0_outputs(4220));
    layer1_outputs(5031) <= (layer0_outputs(1712)) and (layer0_outputs(748));
    layer1_outputs(5032) <= (layer0_outputs(3482)) and not (layer0_outputs(2985));
    layer1_outputs(5033) <= (layer0_outputs(2837)) and (layer0_outputs(3801));
    layer1_outputs(5034) <= (layer0_outputs(3941)) and not (layer0_outputs(1599));
    layer1_outputs(5035) <= not(layer0_outputs(1099)) or (layer0_outputs(376));
    layer1_outputs(5036) <= (layer0_outputs(1689)) and not (layer0_outputs(2686));
    layer1_outputs(5037) <= not(layer0_outputs(1450)) or (layer0_outputs(1307));
    layer1_outputs(5038) <= '1';
    layer1_outputs(5039) <= (layer0_outputs(1213)) and not (layer0_outputs(4474));
    layer1_outputs(5040) <= (layer0_outputs(900)) and not (layer0_outputs(811));
    layer1_outputs(5041) <= (layer0_outputs(3696)) xor (layer0_outputs(2142));
    layer1_outputs(5042) <= '1';
    layer1_outputs(5043) <= not(layer0_outputs(5002));
    layer1_outputs(5044) <= '0';
    layer1_outputs(5045) <= '0';
    layer1_outputs(5046) <= not(layer0_outputs(3637));
    layer1_outputs(5047) <= not(layer0_outputs(243)) or (layer0_outputs(2215));
    layer1_outputs(5048) <= '0';
    layer1_outputs(5049) <= (layer0_outputs(212)) xor (layer0_outputs(2912));
    layer1_outputs(5050) <= not(layer0_outputs(4207));
    layer1_outputs(5051) <= not(layer0_outputs(601));
    layer1_outputs(5052) <= '0';
    layer1_outputs(5053) <= not(layer0_outputs(2476));
    layer1_outputs(5054) <= not(layer0_outputs(4974)) or (layer0_outputs(744));
    layer1_outputs(5055) <= not((layer0_outputs(2478)) or (layer0_outputs(3921)));
    layer1_outputs(5056) <= not(layer0_outputs(2838)) or (layer0_outputs(1994));
    layer1_outputs(5057) <= (layer0_outputs(269)) or (layer0_outputs(1854));
    layer1_outputs(5058) <= '0';
    layer1_outputs(5059) <= not(layer0_outputs(246));
    layer1_outputs(5060) <= not((layer0_outputs(3912)) and (layer0_outputs(4524)));
    layer1_outputs(5061) <= not((layer0_outputs(4220)) and (layer0_outputs(1241)));
    layer1_outputs(5062) <= '1';
    layer1_outputs(5063) <= (layer0_outputs(196)) and not (layer0_outputs(2072));
    layer1_outputs(5064) <= '0';
    layer1_outputs(5065) <= not(layer0_outputs(3948));
    layer1_outputs(5066) <= '1';
    layer1_outputs(5067) <= not((layer0_outputs(1223)) or (layer0_outputs(268)));
    layer1_outputs(5068) <= not(layer0_outputs(194));
    layer1_outputs(5069) <= not(layer0_outputs(2366)) or (layer0_outputs(4035));
    layer1_outputs(5070) <= (layer0_outputs(1225)) or (layer0_outputs(395));
    layer1_outputs(5071) <= not(layer0_outputs(4239)) or (layer0_outputs(3898));
    layer1_outputs(5072) <= (layer0_outputs(4295)) and not (layer0_outputs(4964));
    layer1_outputs(5073) <= (layer0_outputs(1151)) xor (layer0_outputs(5005));
    layer1_outputs(5074) <= layer0_outputs(1948);
    layer1_outputs(5075) <= '0';
    layer1_outputs(5076) <= layer0_outputs(3699);
    layer1_outputs(5077) <= not((layer0_outputs(2387)) or (layer0_outputs(1411)));
    layer1_outputs(5078) <= not(layer0_outputs(4120));
    layer1_outputs(5079) <= not((layer0_outputs(4177)) or (layer0_outputs(1652)));
    layer1_outputs(5080) <= '1';
    layer1_outputs(5081) <= '0';
    layer1_outputs(5082) <= not((layer0_outputs(5091)) or (layer0_outputs(4327)));
    layer1_outputs(5083) <= not(layer0_outputs(2090)) or (layer0_outputs(3090));
    layer1_outputs(5084) <= layer0_outputs(4718);
    layer1_outputs(5085) <= layer0_outputs(4127);
    layer1_outputs(5086) <= (layer0_outputs(1191)) or (layer0_outputs(52));
    layer1_outputs(5087) <= not((layer0_outputs(54)) or (layer0_outputs(2168)));
    layer1_outputs(5088) <= not((layer0_outputs(1639)) and (layer0_outputs(3465)));
    layer1_outputs(5089) <= (layer0_outputs(1664)) or (layer0_outputs(2189));
    layer1_outputs(5090) <= '1';
    layer1_outputs(5091) <= layer0_outputs(757);
    layer1_outputs(5092) <= (layer0_outputs(2620)) or (layer0_outputs(799));
    layer1_outputs(5093) <= not(layer0_outputs(3231));
    layer1_outputs(5094) <= not(layer0_outputs(955));
    layer1_outputs(5095) <= (layer0_outputs(4632)) or (layer0_outputs(3864));
    layer1_outputs(5096) <= not(layer0_outputs(3646)) or (layer0_outputs(1326));
    layer1_outputs(5097) <= not(layer0_outputs(3894)) or (layer0_outputs(923));
    layer1_outputs(5098) <= not(layer0_outputs(2760));
    layer1_outputs(5099) <= '0';
    layer1_outputs(5100) <= layer0_outputs(1377);
    layer1_outputs(5101) <= not((layer0_outputs(4113)) or (layer0_outputs(245)));
    layer1_outputs(5102) <= (layer0_outputs(91)) and not (layer0_outputs(719));
    layer1_outputs(5103) <= not((layer0_outputs(4657)) and (layer0_outputs(703)));
    layer1_outputs(5104) <= layer0_outputs(4708);
    layer1_outputs(5105) <= '1';
    layer1_outputs(5106) <= not(layer0_outputs(3824));
    layer1_outputs(5107) <= not(layer0_outputs(1496));
    layer1_outputs(5108) <= '1';
    layer1_outputs(5109) <= not((layer0_outputs(546)) xor (layer0_outputs(1558)));
    layer1_outputs(5110) <= not(layer0_outputs(2229)) or (layer0_outputs(1571));
    layer1_outputs(5111) <= (layer0_outputs(824)) and not (layer0_outputs(1454));
    layer1_outputs(5112) <= not(layer0_outputs(4924));
    layer1_outputs(5113) <= not((layer0_outputs(738)) and (layer0_outputs(321)));
    layer1_outputs(5114) <= not(layer0_outputs(4758)) or (layer0_outputs(2720));
    layer1_outputs(5115) <= (layer0_outputs(790)) and not (layer0_outputs(889));
    layer1_outputs(5116) <= not(layer0_outputs(1794));
    layer1_outputs(5117) <= layer0_outputs(4723);
    layer1_outputs(5118) <= not((layer0_outputs(4916)) and (layer0_outputs(3877)));
    layer1_outputs(5119) <= (layer0_outputs(2311)) and not (layer0_outputs(451));
    layer2_outputs(0) <= '1';
    layer2_outputs(1) <= layer1_outputs(3800);
    layer2_outputs(2) <= not(layer1_outputs(4636));
    layer2_outputs(3) <= not((layer1_outputs(3970)) or (layer1_outputs(380)));
    layer2_outputs(4) <= layer1_outputs(4079);
    layer2_outputs(5) <= layer1_outputs(2335);
    layer2_outputs(6) <= not(layer1_outputs(2859));
    layer2_outputs(7) <= not((layer1_outputs(4205)) or (layer1_outputs(4662)));
    layer2_outputs(8) <= layer1_outputs(1516);
    layer2_outputs(9) <= not(layer1_outputs(4499)) or (layer1_outputs(3705));
    layer2_outputs(10) <= layer1_outputs(1107);
    layer2_outputs(11) <= (layer1_outputs(3450)) and (layer1_outputs(2807));
    layer2_outputs(12) <= (layer1_outputs(3159)) and (layer1_outputs(1165));
    layer2_outputs(13) <= not(layer1_outputs(4204)) or (layer1_outputs(1310));
    layer2_outputs(14) <= not(layer1_outputs(4842));
    layer2_outputs(15) <= not(layer1_outputs(4966));
    layer2_outputs(16) <= (layer1_outputs(3614)) and not (layer1_outputs(2845));
    layer2_outputs(17) <= layer1_outputs(5106);
    layer2_outputs(18) <= (layer1_outputs(5020)) or (layer1_outputs(1757));
    layer2_outputs(19) <= (layer1_outputs(2995)) and not (layer1_outputs(3144));
    layer2_outputs(20) <= (layer1_outputs(1055)) and not (layer1_outputs(5098));
    layer2_outputs(21) <= '1';
    layer2_outputs(22) <= (layer1_outputs(1902)) and (layer1_outputs(1236));
    layer2_outputs(23) <= not((layer1_outputs(3747)) and (layer1_outputs(2852)));
    layer2_outputs(24) <= (layer1_outputs(1081)) or (layer1_outputs(3693));
    layer2_outputs(25) <= not(layer1_outputs(4686));
    layer2_outputs(26) <= layer1_outputs(2319);
    layer2_outputs(27) <= (layer1_outputs(766)) or (layer1_outputs(5098));
    layer2_outputs(28) <= not((layer1_outputs(3323)) xor (layer1_outputs(2658)));
    layer2_outputs(29) <= not((layer1_outputs(3685)) and (layer1_outputs(1374)));
    layer2_outputs(30) <= layer1_outputs(2774);
    layer2_outputs(31) <= not(layer1_outputs(459)) or (layer1_outputs(1179));
    layer2_outputs(32) <= '1';
    layer2_outputs(33) <= (layer1_outputs(921)) or (layer1_outputs(1232));
    layer2_outputs(34) <= (layer1_outputs(3611)) and (layer1_outputs(4711));
    layer2_outputs(35) <= '1';
    layer2_outputs(36) <= not(layer1_outputs(1399));
    layer2_outputs(37) <= '1';
    layer2_outputs(38) <= not((layer1_outputs(261)) and (layer1_outputs(1614)));
    layer2_outputs(39) <= (layer1_outputs(3097)) and not (layer1_outputs(784));
    layer2_outputs(40) <= (layer1_outputs(3233)) or (layer1_outputs(4376));
    layer2_outputs(41) <= not(layer1_outputs(1928)) or (layer1_outputs(4602));
    layer2_outputs(42) <= not((layer1_outputs(2260)) xor (layer1_outputs(4552)));
    layer2_outputs(43) <= layer1_outputs(3546);
    layer2_outputs(44) <= not(layer1_outputs(4329));
    layer2_outputs(45) <= not((layer1_outputs(4924)) or (layer1_outputs(4526)));
    layer2_outputs(46) <= not(layer1_outputs(4380));
    layer2_outputs(47) <= (layer1_outputs(4715)) and not (layer1_outputs(758));
    layer2_outputs(48) <= '1';
    layer2_outputs(49) <= '0';
    layer2_outputs(50) <= layer1_outputs(841);
    layer2_outputs(51) <= not((layer1_outputs(4235)) or (layer1_outputs(2241)));
    layer2_outputs(52) <= not((layer1_outputs(4194)) or (layer1_outputs(2022)));
    layer2_outputs(53) <= (layer1_outputs(1449)) or (layer1_outputs(3921));
    layer2_outputs(54) <= not(layer1_outputs(1338));
    layer2_outputs(55) <= (layer1_outputs(1354)) and not (layer1_outputs(2265));
    layer2_outputs(56) <= '1';
    layer2_outputs(57) <= (layer1_outputs(3830)) and (layer1_outputs(3985));
    layer2_outputs(58) <= not((layer1_outputs(2151)) and (layer1_outputs(1269)));
    layer2_outputs(59) <= not(layer1_outputs(400)) or (layer1_outputs(746));
    layer2_outputs(60) <= not((layer1_outputs(4577)) or (layer1_outputs(2569)));
    layer2_outputs(61) <= layer1_outputs(4074);
    layer2_outputs(62) <= not(layer1_outputs(1170)) or (layer1_outputs(1714));
    layer2_outputs(63) <= not(layer1_outputs(4965)) or (layer1_outputs(3114));
    layer2_outputs(64) <= not(layer1_outputs(3458)) or (layer1_outputs(2543));
    layer2_outputs(65) <= not(layer1_outputs(3898)) or (layer1_outputs(1942));
    layer2_outputs(66) <= '0';
    layer2_outputs(67) <= layer1_outputs(4114);
    layer2_outputs(68) <= not(layer1_outputs(5027));
    layer2_outputs(69) <= (layer1_outputs(2822)) and not (layer1_outputs(2190));
    layer2_outputs(70) <= '0';
    layer2_outputs(71) <= '0';
    layer2_outputs(72) <= not(layer1_outputs(3341)) or (layer1_outputs(1646));
    layer2_outputs(73) <= not(layer1_outputs(3001)) or (layer1_outputs(2421));
    layer2_outputs(74) <= layer1_outputs(923);
    layer2_outputs(75) <= (layer1_outputs(1230)) and not (layer1_outputs(1446));
    layer2_outputs(76) <= not((layer1_outputs(1950)) xor (layer1_outputs(1417)));
    layer2_outputs(77) <= not(layer1_outputs(3956)) or (layer1_outputs(766));
    layer2_outputs(78) <= not(layer1_outputs(3827)) or (layer1_outputs(4633));
    layer2_outputs(79) <= not((layer1_outputs(4679)) or (layer1_outputs(314)));
    layer2_outputs(80) <= (layer1_outputs(3814)) and not (layer1_outputs(624));
    layer2_outputs(81) <= '1';
    layer2_outputs(82) <= layer1_outputs(2500);
    layer2_outputs(83) <= layer1_outputs(5109);
    layer2_outputs(84) <= '0';
    layer2_outputs(85) <= not((layer1_outputs(1669)) and (layer1_outputs(4682)));
    layer2_outputs(86) <= (layer1_outputs(1233)) or (layer1_outputs(4268));
    layer2_outputs(87) <= not(layer1_outputs(4280));
    layer2_outputs(88) <= (layer1_outputs(5096)) and not (layer1_outputs(103));
    layer2_outputs(89) <= (layer1_outputs(4806)) and not (layer1_outputs(1699));
    layer2_outputs(90) <= layer1_outputs(1302);
    layer2_outputs(91) <= '1';
    layer2_outputs(92) <= not(layer1_outputs(2086)) or (layer1_outputs(1216));
    layer2_outputs(93) <= (layer1_outputs(2098)) and not (layer1_outputs(368));
    layer2_outputs(94) <= not((layer1_outputs(3301)) or (layer1_outputs(2163)));
    layer2_outputs(95) <= not(layer1_outputs(659));
    layer2_outputs(96) <= (layer1_outputs(3248)) and (layer1_outputs(1105));
    layer2_outputs(97) <= not(layer1_outputs(3773)) or (layer1_outputs(4500));
    layer2_outputs(98) <= '1';
    layer2_outputs(99) <= not((layer1_outputs(4016)) or (layer1_outputs(3876)));
    layer2_outputs(100) <= (layer1_outputs(496)) and not (layer1_outputs(4590));
    layer2_outputs(101) <= (layer1_outputs(4115)) and (layer1_outputs(4482));
    layer2_outputs(102) <= not((layer1_outputs(320)) and (layer1_outputs(4557)));
    layer2_outputs(103) <= '0';
    layer2_outputs(104) <= not(layer1_outputs(738)) or (layer1_outputs(1852));
    layer2_outputs(105) <= (layer1_outputs(4448)) and not (layer1_outputs(1278));
    layer2_outputs(106) <= layer1_outputs(2921);
    layer2_outputs(107) <= (layer1_outputs(2557)) and not (layer1_outputs(3464));
    layer2_outputs(108) <= '1';
    layer2_outputs(109) <= not(layer1_outputs(91));
    layer2_outputs(110) <= not(layer1_outputs(4079)) or (layer1_outputs(599));
    layer2_outputs(111) <= layer1_outputs(4639);
    layer2_outputs(112) <= not((layer1_outputs(740)) or (layer1_outputs(3448)));
    layer2_outputs(113) <= not(layer1_outputs(2539)) or (layer1_outputs(4953));
    layer2_outputs(114) <= '0';
    layer2_outputs(115) <= (layer1_outputs(3706)) and not (layer1_outputs(195));
    layer2_outputs(116) <= not(layer1_outputs(2908)) or (layer1_outputs(4439));
    layer2_outputs(117) <= layer1_outputs(2571);
    layer2_outputs(118) <= (layer1_outputs(2645)) or (layer1_outputs(2374));
    layer2_outputs(119) <= layer1_outputs(3277);
    layer2_outputs(120) <= (layer1_outputs(4219)) and (layer1_outputs(1341));
    layer2_outputs(121) <= not(layer1_outputs(4688));
    layer2_outputs(122) <= '1';
    layer2_outputs(123) <= '0';
    layer2_outputs(124) <= (layer1_outputs(2414)) or (layer1_outputs(1193));
    layer2_outputs(125) <= not(layer1_outputs(2277));
    layer2_outputs(126) <= not(layer1_outputs(1666));
    layer2_outputs(127) <= not(layer1_outputs(3709));
    layer2_outputs(128) <= (layer1_outputs(3473)) and (layer1_outputs(2384));
    layer2_outputs(129) <= (layer1_outputs(340)) or (layer1_outputs(1943));
    layer2_outputs(130) <= not((layer1_outputs(5048)) and (layer1_outputs(5039)));
    layer2_outputs(131) <= not(layer1_outputs(2600)) or (layer1_outputs(899));
    layer2_outputs(132) <= (layer1_outputs(4739)) and not (layer1_outputs(612));
    layer2_outputs(133) <= not((layer1_outputs(2923)) xor (layer1_outputs(1891)));
    layer2_outputs(134) <= (layer1_outputs(846)) and not (layer1_outputs(4003));
    layer2_outputs(135) <= not((layer1_outputs(3665)) or (layer1_outputs(1365)));
    layer2_outputs(136) <= '1';
    layer2_outputs(137) <= (layer1_outputs(2608)) and not (layer1_outputs(790));
    layer2_outputs(138) <= '0';
    layer2_outputs(139) <= layer1_outputs(1227);
    layer2_outputs(140) <= not(layer1_outputs(4713));
    layer2_outputs(141) <= not((layer1_outputs(3343)) or (layer1_outputs(562)));
    layer2_outputs(142) <= not((layer1_outputs(876)) and (layer1_outputs(2757)));
    layer2_outputs(143) <= (layer1_outputs(3328)) or (layer1_outputs(3764));
    layer2_outputs(144) <= layer1_outputs(2063);
    layer2_outputs(145) <= layer1_outputs(2882);
    layer2_outputs(146) <= not(layer1_outputs(1308));
    layer2_outputs(147) <= layer1_outputs(4000);
    layer2_outputs(148) <= layer1_outputs(5105);
    layer2_outputs(149) <= layer1_outputs(1854);
    layer2_outputs(150) <= '0';
    layer2_outputs(151) <= not((layer1_outputs(74)) and (layer1_outputs(2770)));
    layer2_outputs(152) <= not(layer1_outputs(3966));
    layer2_outputs(153) <= (layer1_outputs(4517)) or (layer1_outputs(4180));
    layer2_outputs(154) <= (layer1_outputs(3216)) or (layer1_outputs(3771));
    layer2_outputs(155) <= '1';
    layer2_outputs(156) <= (layer1_outputs(3252)) and not (layer1_outputs(1421));
    layer2_outputs(157) <= layer1_outputs(1208);
    layer2_outputs(158) <= not((layer1_outputs(1019)) or (layer1_outputs(250)));
    layer2_outputs(159) <= not(layer1_outputs(3338)) or (layer1_outputs(4601));
    layer2_outputs(160) <= not(layer1_outputs(5055));
    layer2_outputs(161) <= layer1_outputs(1330);
    layer2_outputs(162) <= layer1_outputs(2857);
    layer2_outputs(163) <= '1';
    layer2_outputs(164) <= not(layer1_outputs(2210));
    layer2_outputs(165) <= not(layer1_outputs(2412)) or (layer1_outputs(252));
    layer2_outputs(166) <= '1';
    layer2_outputs(167) <= layer1_outputs(4034);
    layer2_outputs(168) <= (layer1_outputs(1446)) or (layer1_outputs(4304));
    layer2_outputs(169) <= layer1_outputs(1809);
    layer2_outputs(170) <= layer1_outputs(1667);
    layer2_outputs(171) <= layer1_outputs(2227);
    layer2_outputs(172) <= (layer1_outputs(2820)) and not (layer1_outputs(2044));
    layer2_outputs(173) <= not(layer1_outputs(965)) or (layer1_outputs(4753));
    layer2_outputs(174) <= (layer1_outputs(3989)) or (layer1_outputs(494));
    layer2_outputs(175) <= (layer1_outputs(1932)) or (layer1_outputs(4742));
    layer2_outputs(176) <= not(layer1_outputs(4093));
    layer2_outputs(177) <= '1';
    layer2_outputs(178) <= not((layer1_outputs(904)) and (layer1_outputs(4480)));
    layer2_outputs(179) <= not(layer1_outputs(4670));
    layer2_outputs(180) <= not((layer1_outputs(3970)) or (layer1_outputs(4024)));
    layer2_outputs(181) <= (layer1_outputs(4317)) xor (layer1_outputs(1313));
    layer2_outputs(182) <= not((layer1_outputs(2214)) or (layer1_outputs(1481)));
    layer2_outputs(183) <= layer1_outputs(3337);
    layer2_outputs(184) <= (layer1_outputs(2306)) and not (layer1_outputs(3258));
    layer2_outputs(185) <= layer1_outputs(2509);
    layer2_outputs(186) <= (layer1_outputs(2445)) and not (layer1_outputs(4957));
    layer2_outputs(187) <= not(layer1_outputs(295)) or (layer1_outputs(822));
    layer2_outputs(188) <= layer1_outputs(1138);
    layer2_outputs(189) <= not(layer1_outputs(4771));
    layer2_outputs(190) <= layer1_outputs(4930);
    layer2_outputs(191) <= (layer1_outputs(3836)) and not (layer1_outputs(1741));
    layer2_outputs(192) <= (layer1_outputs(651)) or (layer1_outputs(4056));
    layer2_outputs(193) <= '1';
    layer2_outputs(194) <= not(layer1_outputs(2394));
    layer2_outputs(195) <= layer1_outputs(3818);
    layer2_outputs(196) <= not(layer1_outputs(2157)) or (layer1_outputs(4195));
    layer2_outputs(197) <= (layer1_outputs(2030)) and not (layer1_outputs(2154));
    layer2_outputs(198) <= not((layer1_outputs(3797)) and (layer1_outputs(1845)));
    layer2_outputs(199) <= (layer1_outputs(3794)) and not (layer1_outputs(1406));
    layer2_outputs(200) <= not(layer1_outputs(2697)) or (layer1_outputs(3975));
    layer2_outputs(201) <= (layer1_outputs(133)) or (layer1_outputs(2240));
    layer2_outputs(202) <= '1';
    layer2_outputs(203) <= (layer1_outputs(3542)) and not (layer1_outputs(4479));
    layer2_outputs(204) <= not(layer1_outputs(4542));
    layer2_outputs(205) <= '0';
    layer2_outputs(206) <= '1';
    layer2_outputs(207) <= (layer1_outputs(1298)) and not (layer1_outputs(2905));
    layer2_outputs(208) <= not((layer1_outputs(428)) or (layer1_outputs(5022)));
    layer2_outputs(209) <= not(layer1_outputs(4364));
    layer2_outputs(210) <= '1';
    layer2_outputs(211) <= layer1_outputs(773);
    layer2_outputs(212) <= (layer1_outputs(3903)) and (layer1_outputs(2585));
    layer2_outputs(213) <= layer1_outputs(5070);
    layer2_outputs(214) <= not(layer1_outputs(3208)) or (layer1_outputs(4275));
    layer2_outputs(215) <= '1';
    layer2_outputs(216) <= not(layer1_outputs(4522)) or (layer1_outputs(669));
    layer2_outputs(217) <= not(layer1_outputs(1502));
    layer2_outputs(218) <= not(layer1_outputs(1275));
    layer2_outputs(219) <= layer1_outputs(3916);
    layer2_outputs(220) <= not((layer1_outputs(4958)) xor (layer1_outputs(2549)));
    layer2_outputs(221) <= layer1_outputs(1635);
    layer2_outputs(222) <= not(layer1_outputs(4407));
    layer2_outputs(223) <= (layer1_outputs(2232)) and not (layer1_outputs(2117));
    layer2_outputs(224) <= (layer1_outputs(3095)) and not (layer1_outputs(1358));
    layer2_outputs(225) <= not((layer1_outputs(4987)) and (layer1_outputs(48)));
    layer2_outputs(226) <= '0';
    layer2_outputs(227) <= layer1_outputs(4614);
    layer2_outputs(228) <= not(layer1_outputs(4141)) or (layer1_outputs(1677));
    layer2_outputs(229) <= layer1_outputs(1237);
    layer2_outputs(230) <= (layer1_outputs(3822)) and not (layer1_outputs(3469));
    layer2_outputs(231) <= (layer1_outputs(2141)) or (layer1_outputs(2803));
    layer2_outputs(232) <= not(layer1_outputs(556));
    layer2_outputs(233) <= '0';
    layer2_outputs(234) <= '0';
    layer2_outputs(235) <= (layer1_outputs(3394)) and (layer1_outputs(1056));
    layer2_outputs(236) <= '0';
    layer2_outputs(237) <= (layer1_outputs(3860)) and not (layer1_outputs(3280));
    layer2_outputs(238) <= (layer1_outputs(2614)) and not (layer1_outputs(3599));
    layer2_outputs(239) <= not(layer1_outputs(1976)) or (layer1_outputs(4064));
    layer2_outputs(240) <= '0';
    layer2_outputs(241) <= not((layer1_outputs(797)) or (layer1_outputs(632)));
    layer2_outputs(242) <= not((layer1_outputs(2337)) xor (layer1_outputs(1673)));
    layer2_outputs(243) <= layer1_outputs(3222);
    layer2_outputs(244) <= layer1_outputs(2383);
    layer2_outputs(245) <= not(layer1_outputs(2641)) or (layer1_outputs(4239));
    layer2_outputs(246) <= (layer1_outputs(2293)) and not (layer1_outputs(3066));
    layer2_outputs(247) <= not(layer1_outputs(4640));
    layer2_outputs(248) <= layer1_outputs(135);
    layer2_outputs(249) <= not(layer1_outputs(4520)) or (layer1_outputs(2570));
    layer2_outputs(250) <= not(layer1_outputs(3317));
    layer2_outputs(251) <= not(layer1_outputs(4353));
    layer2_outputs(252) <= (layer1_outputs(2748)) xor (layer1_outputs(2265));
    layer2_outputs(253) <= not(layer1_outputs(552)) or (layer1_outputs(2160));
    layer2_outputs(254) <= (layer1_outputs(481)) and not (layer1_outputs(830));
    layer2_outputs(255) <= layer1_outputs(2271);
    layer2_outputs(256) <= '0';
    layer2_outputs(257) <= (layer1_outputs(1772)) and not (layer1_outputs(3558));
    layer2_outputs(258) <= not((layer1_outputs(695)) and (layer1_outputs(3041)));
    layer2_outputs(259) <= not(layer1_outputs(809));
    layer2_outputs(260) <= '1';
    layer2_outputs(261) <= not(layer1_outputs(833));
    layer2_outputs(262) <= not((layer1_outputs(491)) or (layer1_outputs(1332)));
    layer2_outputs(263) <= layer1_outputs(902);
    layer2_outputs(264) <= not((layer1_outputs(2775)) and (layer1_outputs(3029)));
    layer2_outputs(265) <= not((layer1_outputs(3641)) or (layer1_outputs(3191)));
    layer2_outputs(266) <= (layer1_outputs(2514)) and (layer1_outputs(3382));
    layer2_outputs(267) <= (layer1_outputs(2464)) and not (layer1_outputs(4890));
    layer2_outputs(268) <= '0';
    layer2_outputs(269) <= not((layer1_outputs(223)) xor (layer1_outputs(4594)));
    layer2_outputs(270) <= (layer1_outputs(1702)) and (layer1_outputs(498));
    layer2_outputs(271) <= '1';
    layer2_outputs(272) <= not(layer1_outputs(270));
    layer2_outputs(273) <= not((layer1_outputs(850)) and (layer1_outputs(2364)));
    layer2_outputs(274) <= (layer1_outputs(2393)) and not (layer1_outputs(2741));
    layer2_outputs(275) <= not(layer1_outputs(3986));
    layer2_outputs(276) <= not(layer1_outputs(1165)) or (layer1_outputs(3869));
    layer2_outputs(277) <= (layer1_outputs(1335)) and not (layer1_outputs(3693));
    layer2_outputs(278) <= not((layer1_outputs(138)) and (layer1_outputs(1276)));
    layer2_outputs(279) <= not(layer1_outputs(4502));
    layer2_outputs(280) <= not((layer1_outputs(725)) xor (layer1_outputs(1966)));
    layer2_outputs(281) <= not(layer1_outputs(1841));
    layer2_outputs(282) <= not(layer1_outputs(4863));
    layer2_outputs(283) <= not(layer1_outputs(3164));
    layer2_outputs(284) <= not((layer1_outputs(5053)) and (layer1_outputs(2475)));
    layer2_outputs(285) <= (layer1_outputs(940)) and not (layer1_outputs(1696));
    layer2_outputs(286) <= not(layer1_outputs(3892));
    layer2_outputs(287) <= layer1_outputs(1778);
    layer2_outputs(288) <= not(layer1_outputs(1559));
    layer2_outputs(289) <= layer1_outputs(364);
    layer2_outputs(290) <= not(layer1_outputs(1769)) or (layer1_outputs(1221));
    layer2_outputs(291) <= (layer1_outputs(3403)) or (layer1_outputs(1405));
    layer2_outputs(292) <= not(layer1_outputs(3846));
    layer2_outputs(293) <= layer1_outputs(1750);
    layer2_outputs(294) <= layer1_outputs(2766);
    layer2_outputs(295) <= not(layer1_outputs(1826));
    layer2_outputs(296) <= not(layer1_outputs(184)) or (layer1_outputs(2628));
    layer2_outputs(297) <= (layer1_outputs(2883)) xor (layer1_outputs(626));
    layer2_outputs(298) <= (layer1_outputs(597)) and (layer1_outputs(2755));
    layer2_outputs(299) <= (layer1_outputs(883)) and not (layer1_outputs(1529));
    layer2_outputs(300) <= (layer1_outputs(2168)) or (layer1_outputs(196));
    layer2_outputs(301) <= '0';
    layer2_outputs(302) <= (layer1_outputs(2683)) or (layer1_outputs(2243));
    layer2_outputs(303) <= not(layer1_outputs(3927));
    layer2_outputs(304) <= '1';
    layer2_outputs(305) <= layer1_outputs(2799);
    layer2_outputs(306) <= (layer1_outputs(4643)) or (layer1_outputs(721));
    layer2_outputs(307) <= not(layer1_outputs(3891));
    layer2_outputs(308) <= (layer1_outputs(1134)) or (layer1_outputs(3995));
    layer2_outputs(309) <= not(layer1_outputs(3679)) or (layer1_outputs(2124));
    layer2_outputs(310) <= (layer1_outputs(915)) and not (layer1_outputs(3264));
    layer2_outputs(311) <= (layer1_outputs(2452)) and not (layer1_outputs(1926));
    layer2_outputs(312) <= layer1_outputs(4790);
    layer2_outputs(313) <= layer1_outputs(910);
    layer2_outputs(314) <= not((layer1_outputs(1551)) or (layer1_outputs(3491)));
    layer2_outputs(315) <= layer1_outputs(4364);
    layer2_outputs(316) <= not(layer1_outputs(1844));
    layer2_outputs(317) <= (layer1_outputs(1290)) xor (layer1_outputs(2948));
    layer2_outputs(318) <= (layer1_outputs(2703)) and (layer1_outputs(2299));
    layer2_outputs(319) <= '1';
    layer2_outputs(320) <= not((layer1_outputs(2839)) and (layer1_outputs(2892)));
    layer2_outputs(321) <= (layer1_outputs(173)) and (layer1_outputs(5037));
    layer2_outputs(322) <= (layer1_outputs(1155)) and not (layer1_outputs(3259));
    layer2_outputs(323) <= not(layer1_outputs(539));
    layer2_outputs(324) <= (layer1_outputs(1152)) and (layer1_outputs(3929));
    layer2_outputs(325) <= (layer1_outputs(2008)) and (layer1_outputs(3773));
    layer2_outputs(326) <= (layer1_outputs(1674)) and (layer1_outputs(211));
    layer2_outputs(327) <= '1';
    layer2_outputs(328) <= not((layer1_outputs(2790)) or (layer1_outputs(1647)));
    layer2_outputs(329) <= layer1_outputs(2435);
    layer2_outputs(330) <= layer1_outputs(730);
    layer2_outputs(331) <= layer1_outputs(2517);
    layer2_outputs(332) <= (layer1_outputs(4563)) and not (layer1_outputs(919));
    layer2_outputs(333) <= (layer1_outputs(4975)) and not (layer1_outputs(2039));
    layer2_outputs(334) <= '0';
    layer2_outputs(335) <= layer1_outputs(4627);
    layer2_outputs(336) <= '1';
    layer2_outputs(337) <= layer1_outputs(119);
    layer2_outputs(338) <= '0';
    layer2_outputs(339) <= '0';
    layer2_outputs(340) <= '0';
    layer2_outputs(341) <= (layer1_outputs(1014)) and (layer1_outputs(1699));
    layer2_outputs(342) <= (layer1_outputs(3075)) or (layer1_outputs(4291));
    layer2_outputs(343) <= not(layer1_outputs(741));
    layer2_outputs(344) <= layer1_outputs(3962);
    layer2_outputs(345) <= not((layer1_outputs(1642)) or (layer1_outputs(665)));
    layer2_outputs(346) <= not(layer1_outputs(3178));
    layer2_outputs(347) <= not(layer1_outputs(3262)) or (layer1_outputs(3171));
    layer2_outputs(348) <= not(layer1_outputs(3832));
    layer2_outputs(349) <= not((layer1_outputs(1487)) and (layer1_outputs(2702)));
    layer2_outputs(350) <= not(layer1_outputs(4584));
    layer2_outputs(351) <= layer1_outputs(950);
    layer2_outputs(352) <= not(layer1_outputs(480));
    layer2_outputs(353) <= '1';
    layer2_outputs(354) <= layer1_outputs(2280);
    layer2_outputs(355) <= '1';
    layer2_outputs(356) <= not(layer1_outputs(1514)) or (layer1_outputs(660));
    layer2_outputs(357) <= (layer1_outputs(431)) and (layer1_outputs(1821));
    layer2_outputs(358) <= (layer1_outputs(4223)) or (layer1_outputs(1675));
    layer2_outputs(359) <= not(layer1_outputs(222));
    layer2_outputs(360) <= not((layer1_outputs(5101)) and (layer1_outputs(214)));
    layer2_outputs(361) <= '1';
    layer2_outputs(362) <= not(layer1_outputs(2925));
    layer2_outputs(363) <= not(layer1_outputs(4425)) or (layer1_outputs(878));
    layer2_outputs(364) <= not(layer1_outputs(112));
    layer2_outputs(365) <= not((layer1_outputs(4089)) and (layer1_outputs(1892)));
    layer2_outputs(366) <= not((layer1_outputs(663)) and (layer1_outputs(3770)));
    layer2_outputs(367) <= not(layer1_outputs(2854));
    layer2_outputs(368) <= not(layer1_outputs(4759));
    layer2_outputs(369) <= not(layer1_outputs(2058)) or (layer1_outputs(3518));
    layer2_outputs(370) <= not(layer1_outputs(1972)) or (layer1_outputs(566));
    layer2_outputs(371) <= not((layer1_outputs(1513)) or (layer1_outputs(1994)));
    layer2_outputs(372) <= '0';
    layer2_outputs(373) <= not((layer1_outputs(953)) and (layer1_outputs(3994)));
    layer2_outputs(374) <= not(layer1_outputs(4549));
    layer2_outputs(375) <= not(layer1_outputs(1970)) or (layer1_outputs(4462));
    layer2_outputs(376) <= '1';
    layer2_outputs(377) <= layer1_outputs(1384);
    layer2_outputs(378) <= (layer1_outputs(4039)) and not (layer1_outputs(1648));
    layer2_outputs(379) <= not(layer1_outputs(1780)) or (layer1_outputs(4869));
    layer2_outputs(380) <= '1';
    layer2_outputs(381) <= (layer1_outputs(2196)) and not (layer1_outputs(996));
    layer2_outputs(382) <= (layer1_outputs(2646)) and (layer1_outputs(2498));
    layer2_outputs(383) <= not(layer1_outputs(2825));
    layer2_outputs(384) <= not((layer1_outputs(1527)) and (layer1_outputs(4538)));
    layer2_outputs(385) <= not(layer1_outputs(644));
    layer2_outputs(386) <= '1';
    layer2_outputs(387) <= '0';
    layer2_outputs(388) <= '0';
    layer2_outputs(389) <= (layer1_outputs(3583)) and not (layer1_outputs(1422));
    layer2_outputs(390) <= '1';
    layer2_outputs(391) <= layer1_outputs(367);
    layer2_outputs(392) <= layer1_outputs(4638);
    layer2_outputs(393) <= not(layer1_outputs(2437)) or (layer1_outputs(2510));
    layer2_outputs(394) <= layer1_outputs(4215);
    layer2_outputs(395) <= layer1_outputs(2032);
    layer2_outputs(396) <= (layer1_outputs(333)) or (layer1_outputs(2674));
    layer2_outputs(397) <= not(layer1_outputs(4030));
    layer2_outputs(398) <= '1';
    layer2_outputs(399) <= not(layer1_outputs(3775));
    layer2_outputs(400) <= not(layer1_outputs(2404)) or (layer1_outputs(4599));
    layer2_outputs(401) <= not((layer1_outputs(2911)) and (layer1_outputs(2291)));
    layer2_outputs(402) <= not(layer1_outputs(1861));
    layer2_outputs(403) <= (layer1_outputs(1220)) and not (layer1_outputs(2246));
    layer2_outputs(404) <= not((layer1_outputs(2982)) or (layer1_outputs(4651)));
    layer2_outputs(405) <= not(layer1_outputs(4838)) or (layer1_outputs(2624));
    layer2_outputs(406) <= not((layer1_outputs(3497)) and (layer1_outputs(781)));
    layer2_outputs(407) <= (layer1_outputs(1402)) and not (layer1_outputs(1396));
    layer2_outputs(408) <= not((layer1_outputs(4327)) or (layer1_outputs(1962)));
    layer2_outputs(409) <= '0';
    layer2_outputs(410) <= not((layer1_outputs(4333)) and (layer1_outputs(3958)));
    layer2_outputs(411) <= (layer1_outputs(2588)) or (layer1_outputs(4664));
    layer2_outputs(412) <= not((layer1_outputs(3222)) or (layer1_outputs(1399)));
    layer2_outputs(413) <= not(layer1_outputs(3749)) or (layer1_outputs(2791));
    layer2_outputs(414) <= (layer1_outputs(555)) or (layer1_outputs(2759));
    layer2_outputs(415) <= (layer1_outputs(4826)) and not (layer1_outputs(3295));
    layer2_outputs(416) <= not(layer1_outputs(1971));
    layer2_outputs(417) <= not((layer1_outputs(3392)) and (layer1_outputs(2140)));
    layer2_outputs(418) <= layer1_outputs(3532);
    layer2_outputs(419) <= not(layer1_outputs(3958));
    layer2_outputs(420) <= layer1_outputs(1965);
    layer2_outputs(421) <= not(layer1_outputs(2614)) or (layer1_outputs(777));
    layer2_outputs(422) <= '0';
    layer2_outputs(423) <= (layer1_outputs(2827)) or (layer1_outputs(2097));
    layer2_outputs(424) <= '0';
    layer2_outputs(425) <= layer1_outputs(1742);
    layer2_outputs(426) <= not(layer1_outputs(4161)) or (layer1_outputs(1190));
    layer2_outputs(427) <= layer1_outputs(4930);
    layer2_outputs(428) <= not((layer1_outputs(1352)) xor (layer1_outputs(3256)));
    layer2_outputs(429) <= (layer1_outputs(2992)) and not (layer1_outputs(5011));
    layer2_outputs(430) <= not(layer1_outputs(185));
    layer2_outputs(431) <= (layer1_outputs(1035)) or (layer1_outputs(1116));
    layer2_outputs(432) <= not((layer1_outputs(1061)) or (layer1_outputs(2637)));
    layer2_outputs(433) <= not((layer1_outputs(316)) and (layer1_outputs(5093)));
    layer2_outputs(434) <= '1';
    layer2_outputs(435) <= layer1_outputs(3004);
    layer2_outputs(436) <= '0';
    layer2_outputs(437) <= (layer1_outputs(4848)) and not (layer1_outputs(408));
    layer2_outputs(438) <= not(layer1_outputs(3197));
    layer2_outputs(439) <= (layer1_outputs(2155)) and (layer1_outputs(2513));
    layer2_outputs(440) <= not((layer1_outputs(3161)) and (layer1_outputs(1484)));
    layer2_outputs(441) <= not(layer1_outputs(312)) or (layer1_outputs(4674));
    layer2_outputs(442) <= (layer1_outputs(4165)) and not (layer1_outputs(4549));
    layer2_outputs(443) <= (layer1_outputs(1262)) and (layer1_outputs(1195));
    layer2_outputs(444) <= (layer1_outputs(2474)) and not (layer1_outputs(4921));
    layer2_outputs(445) <= '1';
    layer2_outputs(446) <= layer1_outputs(1205);
    layer2_outputs(447) <= '0';
    layer2_outputs(448) <= layer1_outputs(1223);
    layer2_outputs(449) <= '0';
    layer2_outputs(450) <= (layer1_outputs(2846)) or (layer1_outputs(4767));
    layer2_outputs(451) <= (layer1_outputs(73)) and (layer1_outputs(1524));
    layer2_outputs(452) <= (layer1_outputs(1016)) or (layer1_outputs(806));
    layer2_outputs(453) <= (layer1_outputs(3099)) and (layer1_outputs(4307));
    layer2_outputs(454) <= (layer1_outputs(2102)) and not (layer1_outputs(1185));
    layer2_outputs(455) <= not((layer1_outputs(4351)) or (layer1_outputs(4265)));
    layer2_outputs(456) <= (layer1_outputs(2085)) xor (layer1_outputs(2696));
    layer2_outputs(457) <= (layer1_outputs(4008)) or (layer1_outputs(2726));
    layer2_outputs(458) <= not(layer1_outputs(1559));
    layer2_outputs(459) <= not((layer1_outputs(895)) or (layer1_outputs(5088)));
    layer2_outputs(460) <= '1';
    layer2_outputs(461) <= not(layer1_outputs(4975)) or (layer1_outputs(3567));
    layer2_outputs(462) <= not(layer1_outputs(1026));
    layer2_outputs(463) <= not((layer1_outputs(2850)) or (layer1_outputs(3261)));
    layer2_outputs(464) <= not(layer1_outputs(707));
    layer2_outputs(465) <= '1';
    layer2_outputs(466) <= (layer1_outputs(74)) and not (layer1_outputs(333));
    layer2_outputs(467) <= not(layer1_outputs(3577)) or (layer1_outputs(989));
    layer2_outputs(468) <= (layer1_outputs(1478)) and not (layer1_outputs(2501));
    layer2_outputs(469) <= (layer1_outputs(4237)) and (layer1_outputs(2963));
    layer2_outputs(470) <= not(layer1_outputs(297));
    layer2_outputs(471) <= not((layer1_outputs(2914)) and (layer1_outputs(4207)));
    layer2_outputs(472) <= not(layer1_outputs(4323)) or (layer1_outputs(4713));
    layer2_outputs(473) <= not(layer1_outputs(3057));
    layer2_outputs(474) <= not(layer1_outputs(2591)) or (layer1_outputs(2684));
    layer2_outputs(475) <= (layer1_outputs(3096)) or (layer1_outputs(4488));
    layer2_outputs(476) <= layer1_outputs(283);
    layer2_outputs(477) <= not(layer1_outputs(2260));
    layer2_outputs(478) <= (layer1_outputs(203)) and not (layer1_outputs(232));
    layer2_outputs(479) <= not(layer1_outputs(1461));
    layer2_outputs(480) <= not((layer1_outputs(1768)) and (layer1_outputs(274)));
    layer2_outputs(481) <= not(layer1_outputs(645)) or (layer1_outputs(3636));
    layer2_outputs(482) <= (layer1_outputs(4358)) or (layer1_outputs(3506));
    layer2_outputs(483) <= not(layer1_outputs(1192)) or (layer1_outputs(300));
    layer2_outputs(484) <= not(layer1_outputs(943)) or (layer1_outputs(909));
    layer2_outputs(485) <= layer1_outputs(466);
    layer2_outputs(486) <= layer1_outputs(3347);
    layer2_outputs(487) <= not(layer1_outputs(4337));
    layer2_outputs(488) <= (layer1_outputs(3211)) and not (layer1_outputs(5010));
    layer2_outputs(489) <= (layer1_outputs(3580)) and not (layer1_outputs(977));
    layer2_outputs(490) <= not((layer1_outputs(572)) or (layer1_outputs(3777)));
    layer2_outputs(491) <= (layer1_outputs(5077)) and not (layer1_outputs(4298));
    layer2_outputs(492) <= (layer1_outputs(2945)) and not (layer1_outputs(941));
    layer2_outputs(493) <= '1';
    layer2_outputs(494) <= (layer1_outputs(4421)) and not (layer1_outputs(4795));
    layer2_outputs(495) <= not(layer1_outputs(2448));
    layer2_outputs(496) <= not(layer1_outputs(872));
    layer2_outputs(497) <= not(layer1_outputs(4098));
    layer2_outputs(498) <= (layer1_outputs(1805)) and not (layer1_outputs(1492));
    layer2_outputs(499) <= (layer1_outputs(4120)) xor (layer1_outputs(2153));
    layer2_outputs(500) <= (layer1_outputs(503)) or (layer1_outputs(905));
    layer2_outputs(501) <= '0';
    layer2_outputs(502) <= layer1_outputs(568);
    layer2_outputs(503) <= not((layer1_outputs(322)) or (layer1_outputs(1651)));
    layer2_outputs(504) <= layer1_outputs(803);
    layer2_outputs(505) <= layer1_outputs(4345);
    layer2_outputs(506) <= not((layer1_outputs(1042)) and (layer1_outputs(2228)));
    layer2_outputs(507) <= layer1_outputs(1651);
    layer2_outputs(508) <= not(layer1_outputs(4755));
    layer2_outputs(509) <= (layer1_outputs(2245)) and (layer1_outputs(615));
    layer2_outputs(510) <= not((layer1_outputs(545)) and (layer1_outputs(2822)));
    layer2_outputs(511) <= not(layer1_outputs(3525)) or (layer1_outputs(2152));
    layer2_outputs(512) <= not((layer1_outputs(1630)) and (layer1_outputs(911)));
    layer2_outputs(513) <= not(layer1_outputs(5047)) or (layer1_outputs(1940));
    layer2_outputs(514) <= layer1_outputs(2633);
    layer2_outputs(515) <= (layer1_outputs(4973)) or (layer1_outputs(97));
    layer2_outputs(516) <= not(layer1_outputs(3056));
    layer2_outputs(517) <= (layer1_outputs(1151)) and (layer1_outputs(4025));
    layer2_outputs(518) <= '1';
    layer2_outputs(519) <= layer1_outputs(676);
    layer2_outputs(520) <= '0';
    layer2_outputs(521) <= not((layer1_outputs(3429)) and (layer1_outputs(191)));
    layer2_outputs(522) <= (layer1_outputs(482)) or (layer1_outputs(2557));
    layer2_outputs(523) <= '1';
    layer2_outputs(524) <= not(layer1_outputs(2090)) or (layer1_outputs(188));
    layer2_outputs(525) <= layer1_outputs(4375);
    layer2_outputs(526) <= '0';
    layer2_outputs(527) <= not(layer1_outputs(240));
    layer2_outputs(528) <= not(layer1_outputs(1457)) or (layer1_outputs(3052));
    layer2_outputs(529) <= (layer1_outputs(4613)) and not (layer1_outputs(1475));
    layer2_outputs(530) <= layer1_outputs(3534);
    layer2_outputs(531) <= '0';
    layer2_outputs(532) <= not((layer1_outputs(1864)) or (layer1_outputs(1483)));
    layer2_outputs(533) <= (layer1_outputs(4211)) or (layer1_outputs(4982));
    layer2_outputs(534) <= (layer1_outputs(981)) and not (layer1_outputs(4157));
    layer2_outputs(535) <= not(layer1_outputs(4773)) or (layer1_outputs(4188));
    layer2_outputs(536) <= layer1_outputs(3498);
    layer2_outputs(537) <= '1';
    layer2_outputs(538) <= layer1_outputs(1226);
    layer2_outputs(539) <= (layer1_outputs(3678)) or (layer1_outputs(4203));
    layer2_outputs(540) <= '1';
    layer2_outputs(541) <= '0';
    layer2_outputs(542) <= layer1_outputs(3844);
    layer2_outputs(543) <= (layer1_outputs(3087)) and not (layer1_outputs(3104));
    layer2_outputs(544) <= (layer1_outputs(4067)) and not (layer1_outputs(141));
    layer2_outputs(545) <= '0';
    layer2_outputs(546) <= (layer1_outputs(2899)) and (layer1_outputs(990));
    layer2_outputs(547) <= not((layer1_outputs(3681)) and (layer1_outputs(2488)));
    layer2_outputs(548) <= not((layer1_outputs(1460)) and (layer1_outputs(4249)));
    layer2_outputs(549) <= not(layer1_outputs(76));
    layer2_outputs(550) <= (layer1_outputs(4678)) and not (layer1_outputs(3238));
    layer2_outputs(551) <= not(layer1_outputs(2284)) or (layer1_outputs(4272));
    layer2_outputs(552) <= not(layer1_outputs(4187));
    layer2_outputs(553) <= not(layer1_outputs(1783));
    layer2_outputs(554) <= not(layer1_outputs(3247));
    layer2_outputs(555) <= layer1_outputs(2201);
    layer2_outputs(556) <= not(layer1_outputs(1680));
    layer2_outputs(557) <= layer1_outputs(3753);
    layer2_outputs(558) <= layer1_outputs(4084);
    layer2_outputs(559) <= not((layer1_outputs(4830)) and (layer1_outputs(3557)));
    layer2_outputs(560) <= (layer1_outputs(2366)) and (layer1_outputs(62));
    layer2_outputs(561) <= not(layer1_outputs(3688));
    layer2_outputs(562) <= (layer1_outputs(2856)) and (layer1_outputs(2867));
    layer2_outputs(563) <= layer1_outputs(5037);
    layer2_outputs(564) <= layer1_outputs(4739);
    layer2_outputs(565) <= not(layer1_outputs(3586));
    layer2_outputs(566) <= layer1_outputs(4949);
    layer2_outputs(567) <= layer1_outputs(2544);
    layer2_outputs(568) <= not((layer1_outputs(4638)) and (layer1_outputs(2076)));
    layer2_outputs(569) <= not(layer1_outputs(16)) or (layer1_outputs(4749));
    layer2_outputs(570) <= (layer1_outputs(2918)) and not (layer1_outputs(747));
    layer2_outputs(571) <= layer1_outputs(3111);
    layer2_outputs(572) <= not(layer1_outputs(285));
    layer2_outputs(573) <= not((layer1_outputs(319)) or (layer1_outputs(3602)));
    layer2_outputs(574) <= not(layer1_outputs(1372));
    layer2_outputs(575) <= not((layer1_outputs(4601)) or (layer1_outputs(2673)));
    layer2_outputs(576) <= (layer1_outputs(3072)) and not (layer1_outputs(3213));
    layer2_outputs(577) <= (layer1_outputs(2134)) and not (layer1_outputs(2737));
    layer2_outputs(578) <= not((layer1_outputs(1019)) and (layer1_outputs(1526)));
    layer2_outputs(579) <= not(layer1_outputs(1979));
    layer2_outputs(580) <= not((layer1_outputs(3956)) and (layer1_outputs(2794)));
    layer2_outputs(581) <= not(layer1_outputs(4326));
    layer2_outputs(582) <= '0';
    layer2_outputs(583) <= (layer1_outputs(4963)) and not (layer1_outputs(1095));
    layer2_outputs(584) <= not(layer1_outputs(2075));
    layer2_outputs(585) <= (layer1_outputs(1726)) and not (layer1_outputs(3810));
    layer2_outputs(586) <= '0';
    layer2_outputs(587) <= (layer1_outputs(4244)) or (layer1_outputs(2891));
    layer2_outputs(588) <= '0';
    layer2_outputs(589) <= not(layer1_outputs(4394)) or (layer1_outputs(1110));
    layer2_outputs(590) <= layer1_outputs(882);
    layer2_outputs(591) <= layer1_outputs(3108);
    layer2_outputs(592) <= not((layer1_outputs(1134)) and (layer1_outputs(2075)));
    layer2_outputs(593) <= '0';
    layer2_outputs(594) <= '1';
    layer2_outputs(595) <= (layer1_outputs(632)) and not (layer1_outputs(4272));
    layer2_outputs(596) <= not(layer1_outputs(2219)) or (layer1_outputs(1460));
    layer2_outputs(597) <= not(layer1_outputs(3718));
    layer2_outputs(598) <= not(layer1_outputs(2309)) or (layer1_outputs(272));
    layer2_outputs(599) <= not((layer1_outputs(2480)) and (layer1_outputs(1097)));
    layer2_outputs(600) <= (layer1_outputs(3980)) and not (layer1_outputs(1209));
    layer2_outputs(601) <= '0';
    layer2_outputs(602) <= '0';
    layer2_outputs(603) <= (layer1_outputs(2141)) and not (layer1_outputs(5089));
    layer2_outputs(604) <= (layer1_outputs(900)) and not (layer1_outputs(4219));
    layer2_outputs(605) <= not(layer1_outputs(1145)) or (layer1_outputs(2466));
    layer2_outputs(606) <= layer1_outputs(4259);
    layer2_outputs(607) <= layer1_outputs(5056);
    layer2_outputs(608) <= (layer1_outputs(3793)) and (layer1_outputs(1940));
    layer2_outputs(609) <= (layer1_outputs(1423)) and not (layer1_outputs(2819));
    layer2_outputs(610) <= not((layer1_outputs(2891)) or (layer1_outputs(432)));
    layer2_outputs(611) <= '1';
    layer2_outputs(612) <= not(layer1_outputs(2610));
    layer2_outputs(613) <= '1';
    layer2_outputs(614) <= '0';
    layer2_outputs(615) <= '1';
    layer2_outputs(616) <= '0';
    layer2_outputs(617) <= not(layer1_outputs(4653));
    layer2_outputs(618) <= layer1_outputs(3351);
    layer2_outputs(619) <= '1';
    layer2_outputs(620) <= layer1_outputs(588);
    layer2_outputs(621) <= '1';
    layer2_outputs(622) <= (layer1_outputs(4092)) and not (layer1_outputs(3040));
    layer2_outputs(623) <= not(layer1_outputs(1512)) or (layer1_outputs(3383));
    layer2_outputs(624) <= not((layer1_outputs(3087)) and (layer1_outputs(4859)));
    layer2_outputs(625) <= '0';
    layer2_outputs(626) <= not(layer1_outputs(3386));
    layer2_outputs(627) <= not(layer1_outputs(4927)) or (layer1_outputs(3856));
    layer2_outputs(628) <= '0';
    layer2_outputs(629) <= not(layer1_outputs(647));
    layer2_outputs(630) <= '0';
    layer2_outputs(631) <= not(layer1_outputs(4394));
    layer2_outputs(632) <= (layer1_outputs(980)) and (layer1_outputs(126));
    layer2_outputs(633) <= (layer1_outputs(91)) xor (layer1_outputs(4631));
    layer2_outputs(634) <= '0';
    layer2_outputs(635) <= layer1_outputs(405);
    layer2_outputs(636) <= not((layer1_outputs(134)) and (layer1_outputs(3739)));
    layer2_outputs(637) <= (layer1_outputs(4649)) or (layer1_outputs(4422));
    layer2_outputs(638) <= '1';
    layer2_outputs(639) <= layer1_outputs(1937);
    layer2_outputs(640) <= layer1_outputs(3884);
    layer2_outputs(641) <= (layer1_outputs(976)) and not (layer1_outputs(4842));
    layer2_outputs(642) <= not(layer1_outputs(5028));
    layer2_outputs(643) <= (layer1_outputs(3360)) and not (layer1_outputs(2902));
    layer2_outputs(644) <= not((layer1_outputs(2986)) or (layer1_outputs(620)));
    layer2_outputs(645) <= layer1_outputs(2544);
    layer2_outputs(646) <= layer1_outputs(4157);
    layer2_outputs(647) <= not(layer1_outputs(2221)) or (layer1_outputs(2416));
    layer2_outputs(648) <= not((layer1_outputs(1058)) or (layer1_outputs(254)));
    layer2_outputs(649) <= not((layer1_outputs(3370)) and (layer1_outputs(4181)));
    layer2_outputs(650) <= '0';
    layer2_outputs(651) <= layer1_outputs(1155);
    layer2_outputs(652) <= not(layer1_outputs(3230)) or (layer1_outputs(793));
    layer2_outputs(653) <= not((layer1_outputs(2820)) or (layer1_outputs(3085)));
    layer2_outputs(654) <= not(layer1_outputs(2493));
    layer2_outputs(655) <= not(layer1_outputs(2811)) or (layer1_outputs(1214));
    layer2_outputs(656) <= (layer1_outputs(4984)) and not (layer1_outputs(4250));
    layer2_outputs(657) <= not(layer1_outputs(2817));
    layer2_outputs(658) <= '1';
    layer2_outputs(659) <= layer1_outputs(3707);
    layer2_outputs(660) <= not(layer1_outputs(580));
    layer2_outputs(661) <= '1';
    layer2_outputs(662) <= not((layer1_outputs(1227)) and (layer1_outputs(4509)));
    layer2_outputs(663) <= (layer1_outputs(4148)) and not (layer1_outputs(3427));
    layer2_outputs(664) <= (layer1_outputs(1565)) and (layer1_outputs(3944));
    layer2_outputs(665) <= '1';
    layer2_outputs(666) <= '1';
    layer2_outputs(667) <= not(layer1_outputs(2191));
    layer2_outputs(668) <= layer1_outputs(3196);
    layer2_outputs(669) <= layer1_outputs(315);
    layer2_outputs(670) <= (layer1_outputs(2619)) xor (layer1_outputs(1534));
    layer2_outputs(671) <= (layer1_outputs(3725)) or (layer1_outputs(4211));
    layer2_outputs(672) <= (layer1_outputs(1444)) and (layer1_outputs(106));
    layer2_outputs(673) <= not(layer1_outputs(2671));
    layer2_outputs(674) <= layer1_outputs(3477);
    layer2_outputs(675) <= '1';
    layer2_outputs(676) <= not(layer1_outputs(3604)) or (layer1_outputs(609));
    layer2_outputs(677) <= layer1_outputs(2080);
    layer2_outputs(678) <= not(layer1_outputs(2161)) or (layer1_outputs(1532));
    layer2_outputs(679) <= not((layer1_outputs(559)) and (layer1_outputs(1112)));
    layer2_outputs(680) <= (layer1_outputs(1130)) and not (layer1_outputs(102));
    layer2_outputs(681) <= not(layer1_outputs(2743));
    layer2_outputs(682) <= not(layer1_outputs(3156));
    layer2_outputs(683) <= not(layer1_outputs(4514)) or (layer1_outputs(3799));
    layer2_outputs(684) <= (layer1_outputs(1677)) or (layer1_outputs(2167));
    layer2_outputs(685) <= not(layer1_outputs(25)) or (layer1_outputs(842));
    layer2_outputs(686) <= '1';
    layer2_outputs(687) <= not(layer1_outputs(1611));
    layer2_outputs(688) <= not(layer1_outputs(1989));
    layer2_outputs(689) <= not((layer1_outputs(2326)) or (layer1_outputs(674)));
    layer2_outputs(690) <= not(layer1_outputs(1161)) or (layer1_outputs(4423));
    layer2_outputs(691) <= not(layer1_outputs(3026));
    layer2_outputs(692) <= not((layer1_outputs(4945)) and (layer1_outputs(3535)));
    layer2_outputs(693) <= not(layer1_outputs(2561)) or (layer1_outputs(3720));
    layer2_outputs(694) <= layer1_outputs(4530);
    layer2_outputs(695) <= '0';
    layer2_outputs(696) <= not(layer1_outputs(136));
    layer2_outputs(697) <= (layer1_outputs(2606)) or (layer1_outputs(3612));
    layer2_outputs(698) <= not(layer1_outputs(3460)) or (layer1_outputs(696));
    layer2_outputs(699) <= (layer1_outputs(4231)) and not (layer1_outputs(1900));
    layer2_outputs(700) <= (layer1_outputs(3055)) and (layer1_outputs(586));
    layer2_outputs(701) <= not((layer1_outputs(3065)) or (layer1_outputs(1647)));
    layer2_outputs(702) <= (layer1_outputs(1690)) or (layer1_outputs(1077));
    layer2_outputs(703) <= (layer1_outputs(2527)) and not (layer1_outputs(1207));
    layer2_outputs(704) <= '0';
    layer2_outputs(705) <= not(layer1_outputs(1489));
    layer2_outputs(706) <= '1';
    layer2_outputs(707) <= layer1_outputs(767);
    layer2_outputs(708) <= not((layer1_outputs(2248)) or (layer1_outputs(3911)));
    layer2_outputs(709) <= (layer1_outputs(4471)) or (layer1_outputs(4881));
    layer2_outputs(710) <= '0';
    layer2_outputs(711) <= not((layer1_outputs(4035)) or (layer1_outputs(3231)));
    layer2_outputs(712) <= not(layer1_outputs(1127));
    layer2_outputs(713) <= not((layer1_outputs(450)) or (layer1_outputs(1267)));
    layer2_outputs(714) <= not(layer1_outputs(4215)) or (layer1_outputs(1411));
    layer2_outputs(715) <= '1';
    layer2_outputs(716) <= (layer1_outputs(3397)) or (layer1_outputs(1386));
    layer2_outputs(717) <= (layer1_outputs(4525)) or (layer1_outputs(5069));
    layer2_outputs(718) <= layer1_outputs(4262);
    layer2_outputs(719) <= not(layer1_outputs(618));
    layer2_outputs(720) <= (layer1_outputs(4036)) and (layer1_outputs(179));
    layer2_outputs(721) <= (layer1_outputs(3825)) and (layer1_outputs(1802));
    layer2_outputs(722) <= not(layer1_outputs(3653));
    layer2_outputs(723) <= not(layer1_outputs(4100));
    layer2_outputs(724) <= '1';
    layer2_outputs(725) <= '1';
    layer2_outputs(726) <= (layer1_outputs(259)) and (layer1_outputs(2729));
    layer2_outputs(727) <= not((layer1_outputs(442)) or (layer1_outputs(1050)));
    layer2_outputs(728) <= (layer1_outputs(3615)) and not (layer1_outputs(1949));
    layer2_outputs(729) <= layer1_outputs(4171);
    layer2_outputs(730) <= (layer1_outputs(3147)) and not (layer1_outputs(462));
    layer2_outputs(731) <= '0';
    layer2_outputs(732) <= (layer1_outputs(653)) or (layer1_outputs(354));
    layer2_outputs(733) <= '0';
    layer2_outputs(734) <= '0';
    layer2_outputs(735) <= not(layer1_outputs(531));
    layer2_outputs(736) <= layer1_outputs(4122);
    layer2_outputs(737) <= not(layer1_outputs(845));
    layer2_outputs(738) <= not(layer1_outputs(1256));
    layer2_outputs(739) <= '1';
    layer2_outputs(740) <= (layer1_outputs(2190)) and not (layer1_outputs(2041));
    layer2_outputs(741) <= '0';
    layer2_outputs(742) <= '0';
    layer2_outputs(743) <= not((layer1_outputs(3625)) or (layer1_outputs(582)));
    layer2_outputs(744) <= (layer1_outputs(824)) or (layer1_outputs(963));
    layer2_outputs(745) <= '1';
    layer2_outputs(746) <= layer1_outputs(3158);
    layer2_outputs(747) <= (layer1_outputs(906)) and not (layer1_outputs(4917));
    layer2_outputs(748) <= not(layer1_outputs(3987)) or (layer1_outputs(284));
    layer2_outputs(749) <= layer1_outputs(151);
    layer2_outputs(750) <= not(layer1_outputs(152)) or (layer1_outputs(2738));
    layer2_outputs(751) <= layer1_outputs(4858);
    layer2_outputs(752) <= layer1_outputs(3114);
    layer2_outputs(753) <= (layer1_outputs(4782)) or (layer1_outputs(4314));
    layer2_outputs(754) <= layer1_outputs(5103);
    layer2_outputs(755) <= (layer1_outputs(2529)) or (layer1_outputs(3063));
    layer2_outputs(756) <= not((layer1_outputs(4992)) and (layer1_outputs(4736)));
    layer2_outputs(757) <= (layer1_outputs(230)) xor (layer1_outputs(518));
    layer2_outputs(758) <= layer1_outputs(2461);
    layer2_outputs(759) <= (layer1_outputs(4175)) and (layer1_outputs(2085));
    layer2_outputs(760) <= (layer1_outputs(757)) and not (layer1_outputs(4868));
    layer2_outputs(761) <= not(layer1_outputs(1897)) or (layer1_outputs(4172));
    layer2_outputs(762) <= '1';
    layer2_outputs(763) <= (layer1_outputs(912)) or (layer1_outputs(2516));
    layer2_outputs(764) <= not((layer1_outputs(2230)) or (layer1_outputs(5072)));
    layer2_outputs(765) <= not((layer1_outputs(4370)) or (layer1_outputs(1808)));
    layer2_outputs(766) <= (layer1_outputs(2823)) and not (layer1_outputs(2399));
    layer2_outputs(767) <= not(layer1_outputs(553));
    layer2_outputs(768) <= (layer1_outputs(1763)) and not (layer1_outputs(3378));
    layer2_outputs(769) <= not(layer1_outputs(1059));
    layer2_outputs(770) <= not(layer1_outputs(313));
    layer2_outputs(771) <= layer1_outputs(2575);
    layer2_outputs(772) <= layer1_outputs(1658);
    layer2_outputs(773) <= (layer1_outputs(2615)) and not (layer1_outputs(2371));
    layer2_outputs(774) <= not(layer1_outputs(854));
    layer2_outputs(775) <= not(layer1_outputs(3744)) or (layer1_outputs(4826));
    layer2_outputs(776) <= (layer1_outputs(922)) and not (layer1_outputs(446));
    layer2_outputs(777) <= layer1_outputs(205);
    layer2_outputs(778) <= not((layer1_outputs(4867)) and (layer1_outputs(2761)));
    layer2_outputs(779) <= (layer1_outputs(44)) or (layer1_outputs(1773));
    layer2_outputs(780) <= not((layer1_outputs(1079)) or (layer1_outputs(4344)));
    layer2_outputs(781) <= (layer1_outputs(5012)) and not (layer1_outputs(4019));
    layer2_outputs(782) <= layer1_outputs(2420);
    layer2_outputs(783) <= not((layer1_outputs(3854)) or (layer1_outputs(4813)));
    layer2_outputs(784) <= layer1_outputs(207);
    layer2_outputs(785) <= not(layer1_outputs(3620));
    layer2_outputs(786) <= (layer1_outputs(4232)) or (layer1_outputs(2762));
    layer2_outputs(787) <= '1';
    layer2_outputs(788) <= not((layer1_outputs(2510)) and (layer1_outputs(3172)));
    layer2_outputs(789) <= not((layer1_outputs(2461)) or (layer1_outputs(3863)));
    layer2_outputs(790) <= (layer1_outputs(4021)) and not (layer1_outputs(4642));
    layer2_outputs(791) <= not(layer1_outputs(548)) or (layer1_outputs(3751));
    layer2_outputs(792) <= layer1_outputs(3359);
    layer2_outputs(793) <= not(layer1_outputs(4632));
    layer2_outputs(794) <= not(layer1_outputs(533)) or (layer1_outputs(685));
    layer2_outputs(795) <= (layer1_outputs(4331)) and (layer1_outputs(576));
    layer2_outputs(796) <= layer1_outputs(4841);
    layer2_outputs(797) <= '1';
    layer2_outputs(798) <= not(layer1_outputs(3300));
    layer2_outputs(799) <= not(layer1_outputs(2714));
    layer2_outputs(800) <= (layer1_outputs(2823)) and not (layer1_outputs(4086));
    layer2_outputs(801) <= not(layer1_outputs(1695));
    layer2_outputs(802) <= (layer1_outputs(3690)) and not (layer1_outputs(3552));
    layer2_outputs(803) <= layer1_outputs(946);
    layer2_outputs(804) <= '1';
    layer2_outputs(805) <= layer1_outputs(4908);
    layer2_outputs(806) <= '1';
    layer2_outputs(807) <= (layer1_outputs(4783)) and (layer1_outputs(3092));
    layer2_outputs(808) <= not((layer1_outputs(934)) xor (layer1_outputs(2827)));
    layer2_outputs(809) <= layer1_outputs(2642);
    layer2_outputs(810) <= not((layer1_outputs(604)) or (layer1_outputs(829)));
    layer2_outputs(811) <= (layer1_outputs(1904)) and (layer1_outputs(3991));
    layer2_outputs(812) <= (layer1_outputs(1760)) or (layer1_outputs(4188));
    layer2_outputs(813) <= not(layer1_outputs(116)) or (layer1_outputs(4694));
    layer2_outputs(814) <= not(layer1_outputs(4865));
    layer2_outputs(815) <= not((layer1_outputs(2351)) or (layer1_outputs(4407)));
    layer2_outputs(816) <= (layer1_outputs(4195)) and (layer1_outputs(4431));
    layer2_outputs(817) <= not(layer1_outputs(2021)) or (layer1_outputs(2529));
    layer2_outputs(818) <= not(layer1_outputs(4523));
    layer2_outputs(819) <= not(layer1_outputs(3309));
    layer2_outputs(820) <= layer1_outputs(2665);
    layer2_outputs(821) <= layer1_outputs(3718);
    layer2_outputs(822) <= (layer1_outputs(4631)) or (layer1_outputs(4075));
    layer2_outputs(823) <= not(layer1_outputs(2874)) or (layer1_outputs(60));
    layer2_outputs(824) <= (layer1_outputs(1060)) and not (layer1_outputs(810));
    layer2_outputs(825) <= layer1_outputs(2375);
    layer2_outputs(826) <= not(layer1_outputs(3430)) or (layer1_outputs(1066));
    layer2_outputs(827) <= not((layer1_outputs(4420)) or (layer1_outputs(2548)));
    layer2_outputs(828) <= not((layer1_outputs(1567)) or (layer1_outputs(1758)));
    layer2_outputs(829) <= not(layer1_outputs(4497));
    layer2_outputs(830) <= layer1_outputs(4069);
    layer2_outputs(831) <= not(layer1_outputs(3530));
    layer2_outputs(832) <= not((layer1_outputs(2121)) or (layer1_outputs(4446)));
    layer2_outputs(833) <= layer1_outputs(957);
    layer2_outputs(834) <= not(layer1_outputs(992));
    layer2_outputs(835) <= '1';
    layer2_outputs(836) <= (layer1_outputs(500)) and (layer1_outputs(4519));
    layer2_outputs(837) <= not(layer1_outputs(2264)) or (layer1_outputs(4176));
    layer2_outputs(838) <= not(layer1_outputs(461));
    layer2_outputs(839) <= (layer1_outputs(2226)) and not (layer1_outputs(1879));
    layer2_outputs(840) <= (layer1_outputs(2062)) and (layer1_outputs(1696));
    layer2_outputs(841) <= not(layer1_outputs(3865));
    layer2_outputs(842) <= '0';
    layer2_outputs(843) <= layer1_outputs(4249);
    layer2_outputs(844) <= '1';
    layer2_outputs(845) <= (layer1_outputs(278)) and (layer1_outputs(4879));
    layer2_outputs(846) <= not((layer1_outputs(299)) and (layer1_outputs(2842)));
    layer2_outputs(847) <= (layer1_outputs(512)) and not (layer1_outputs(718));
    layer2_outputs(848) <= layer1_outputs(1756);
    layer2_outputs(849) <= not(layer1_outputs(1116));
    layer2_outputs(850) <= (layer1_outputs(1223)) or (layer1_outputs(790));
    layer2_outputs(851) <= not(layer1_outputs(3242));
    layer2_outputs(852) <= (layer1_outputs(2208)) and (layer1_outputs(4418));
    layer2_outputs(853) <= '0';
    layer2_outputs(854) <= layer1_outputs(831);
    layer2_outputs(855) <= not(layer1_outputs(2003));
    layer2_outputs(856) <= (layer1_outputs(3901)) or (layer1_outputs(4008));
    layer2_outputs(857) <= layer1_outputs(2964);
    layer2_outputs(858) <= not(layer1_outputs(1830)) or (layer1_outputs(4425));
    layer2_outputs(859) <= (layer1_outputs(3263)) and (layer1_outputs(1437));
    layer2_outputs(860) <= not(layer1_outputs(3818));
    layer2_outputs(861) <= not((layer1_outputs(2795)) and (layer1_outputs(2989)));
    layer2_outputs(862) <= not(layer1_outputs(145));
    layer2_outputs(863) <= (layer1_outputs(2536)) and not (layer1_outputs(2082));
    layer2_outputs(864) <= (layer1_outputs(4712)) or (layer1_outputs(2768));
    layer2_outputs(865) <= not(layer1_outputs(3895)) or (layer1_outputs(2698));
    layer2_outputs(866) <= layer1_outputs(266);
    layer2_outputs(867) <= (layer1_outputs(4702)) or (layer1_outputs(2422));
    layer2_outputs(868) <= (layer1_outputs(2621)) and not (layer1_outputs(4029));
    layer2_outputs(869) <= layer1_outputs(4789);
    layer2_outputs(870) <= layer1_outputs(300);
    layer2_outputs(871) <= layer1_outputs(3478);
    layer2_outputs(872) <= '1';
    layer2_outputs(873) <= not((layer1_outputs(4833)) or (layer1_outputs(54)));
    layer2_outputs(874) <= not(layer1_outputs(1655));
    layer2_outputs(875) <= layer1_outputs(2550);
    layer2_outputs(876) <= not(layer1_outputs(1402));
    layer2_outputs(877) <= layer1_outputs(4763);
    layer2_outputs(878) <= not((layer1_outputs(746)) and (layer1_outputs(832)));
    layer2_outputs(879) <= '0';
    layer2_outputs(880) <= not(layer1_outputs(22));
    layer2_outputs(881) <= not(layer1_outputs(4291)) or (layer1_outputs(4752));
    layer2_outputs(882) <= '0';
    layer2_outputs(883) <= (layer1_outputs(1534)) and not (layer1_outputs(1663));
    layer2_outputs(884) <= '1';
    layer2_outputs(885) <= (layer1_outputs(1117)) or (layer1_outputs(3167));
    layer2_outputs(886) <= not((layer1_outputs(3749)) and (layer1_outputs(3361)));
    layer2_outputs(887) <= not(layer1_outputs(3376));
    layer2_outputs(888) <= (layer1_outputs(1305)) and not (layer1_outputs(4404));
    layer2_outputs(889) <= (layer1_outputs(2380)) and not (layer1_outputs(1889));
    layer2_outputs(890) <= not(layer1_outputs(695)) or (layer1_outputs(367));
    layer2_outputs(891) <= (layer1_outputs(3367)) and not (layer1_outputs(257));
    layer2_outputs(892) <= (layer1_outputs(3493)) and not (layer1_outputs(879));
    layer2_outputs(893) <= (layer1_outputs(305)) and not (layer1_outputs(2638));
    layer2_outputs(894) <= (layer1_outputs(2087)) or (layer1_outputs(1220));
    layer2_outputs(895) <= '0';
    layer2_outputs(896) <= not(layer1_outputs(1074));
    layer2_outputs(897) <= not((layer1_outputs(4910)) or (layer1_outputs(3571)));
    layer2_outputs(898) <= '1';
    layer2_outputs(899) <= '0';
    layer2_outputs(900) <= (layer1_outputs(1013)) xor (layer1_outputs(4458));
    layer2_outputs(901) <= layer1_outputs(4303);
    layer2_outputs(902) <= (layer1_outputs(4515)) and not (layer1_outputs(3355));
    layer2_outputs(903) <= not(layer1_outputs(3028)) or (layer1_outputs(4890));
    layer2_outputs(904) <= (layer1_outputs(2613)) or (layer1_outputs(3298));
    layer2_outputs(905) <= layer1_outputs(3329);
    layer2_outputs(906) <= not(layer1_outputs(2021));
    layer2_outputs(907) <= (layer1_outputs(1133)) and not (layer1_outputs(4022));
    layer2_outputs(908) <= (layer1_outputs(3180)) and not (layer1_outputs(4635));
    layer2_outputs(909) <= '0';
    layer2_outputs(910) <= not(layer1_outputs(40));
    layer2_outputs(911) <= '1';
    layer2_outputs(912) <= not(layer1_outputs(2376)) or (layer1_outputs(1595));
    layer2_outputs(913) <= (layer1_outputs(1967)) and not (layer1_outputs(3220));
    layer2_outputs(914) <= layer1_outputs(3682);
    layer2_outputs(915) <= '1';
    layer2_outputs(916) <= (layer1_outputs(1636)) or (layer1_outputs(1584));
    layer2_outputs(917) <= (layer1_outputs(4385)) and (layer1_outputs(2997));
    layer2_outputs(918) <= not(layer1_outputs(4166)) or (layer1_outputs(248));
    layer2_outputs(919) <= not(layer1_outputs(553));
    layer2_outputs(920) <= layer1_outputs(3701);
    layer2_outputs(921) <= '0';
    layer2_outputs(922) <= (layer1_outputs(4719)) xor (layer1_outputs(2377));
    layer2_outputs(923) <= '1';
    layer2_outputs(924) <= not(layer1_outputs(3798)) or (layer1_outputs(2727));
    layer2_outputs(925) <= not((layer1_outputs(229)) and (layer1_outputs(4926)));
    layer2_outputs(926) <= (layer1_outputs(2577)) and not (layer1_outputs(3194));
    layer2_outputs(927) <= layer1_outputs(1525);
    layer2_outputs(928) <= '1';
    layer2_outputs(929) <= not(layer1_outputs(4951));
    layer2_outputs(930) <= layer1_outputs(3013);
    layer2_outputs(931) <= not(layer1_outputs(2231)) or (layer1_outputs(3311));
    layer2_outputs(932) <= layer1_outputs(2382);
    layer2_outputs(933) <= not(layer1_outputs(999));
    layer2_outputs(934) <= not(layer1_outputs(2193));
    layer2_outputs(935) <= '1';
    layer2_outputs(936) <= not(layer1_outputs(844));
    layer2_outputs(937) <= not(layer1_outputs(1516)) or (layer1_outputs(1746));
    layer2_outputs(938) <= not((layer1_outputs(2708)) or (layer1_outputs(3118)));
    layer2_outputs(939) <= (layer1_outputs(3466)) and (layer1_outputs(5027));
    layer2_outputs(940) <= '0';
    layer2_outputs(941) <= layer1_outputs(1491);
    layer2_outputs(942) <= (layer1_outputs(2582)) and not (layer1_outputs(2406));
    layer2_outputs(943) <= '0';
    layer2_outputs(944) <= not((layer1_outputs(3886)) or (layer1_outputs(2066)));
    layer2_outputs(945) <= not((layer1_outputs(3783)) and (layer1_outputs(4384)));
    layer2_outputs(946) <= (layer1_outputs(2943)) or (layer1_outputs(4756));
    layer2_outputs(947) <= '1';
    layer2_outputs(948) <= '0';
    layer2_outputs(949) <= not(layer1_outputs(3238));
    layer2_outputs(950) <= layer1_outputs(417);
    layer2_outputs(951) <= (layer1_outputs(1304)) and (layer1_outputs(568));
    layer2_outputs(952) <= (layer1_outputs(393)) or (layer1_outputs(3939));
    layer2_outputs(953) <= not((layer1_outputs(2336)) and (layer1_outputs(2643)));
    layer2_outputs(954) <= '1';
    layer2_outputs(955) <= (layer1_outputs(2929)) and not (layer1_outputs(4383));
    layer2_outputs(956) <= (layer1_outputs(512)) or (layer1_outputs(1336));
    layer2_outputs(957) <= layer1_outputs(2492);
    layer2_outputs(958) <= not((layer1_outputs(3699)) or (layer1_outputs(1166)));
    layer2_outputs(959) <= (layer1_outputs(4490)) and not (layer1_outputs(370));
    layer2_outputs(960) <= not((layer1_outputs(4037)) and (layer1_outputs(4907)));
    layer2_outputs(961) <= not(layer1_outputs(978)) or (layer1_outputs(2406));
    layer2_outputs(962) <= layer1_outputs(547);
    layer2_outputs(963) <= (layer1_outputs(3188)) and not (layer1_outputs(3998));
    layer2_outputs(964) <= not(layer1_outputs(267)) or (layer1_outputs(4108));
    layer2_outputs(965) <= (layer1_outputs(2935)) or (layer1_outputs(4292));
    layer2_outputs(966) <= not((layer1_outputs(2123)) and (layer1_outputs(2784)));
    layer2_outputs(967) <= (layer1_outputs(4317)) and not (layer1_outputs(3377));
    layer2_outputs(968) <= not(layer1_outputs(2515));
    layer2_outputs(969) <= layer1_outputs(2339);
    layer2_outputs(970) <= not(layer1_outputs(4286)) or (layer1_outputs(3742));
    layer2_outputs(971) <= '0';
    layer2_outputs(972) <= not(layer1_outputs(260)) or (layer1_outputs(2354));
    layer2_outputs(973) <= (layer1_outputs(2342)) and not (layer1_outputs(1037));
    layer2_outputs(974) <= (layer1_outputs(3324)) and (layer1_outputs(1420));
    layer2_outputs(975) <= layer1_outputs(2796);
    layer2_outputs(976) <= not((layer1_outputs(3977)) and (layer1_outputs(1419)));
    layer2_outputs(977) <= not(layer1_outputs(4789)) or (layer1_outputs(1682));
    layer2_outputs(978) <= not(layer1_outputs(4698)) or (layer1_outputs(366));
    layer2_outputs(979) <= not(layer1_outputs(1451)) or (layer1_outputs(4712));
    layer2_outputs(980) <= (layer1_outputs(4764)) and not (layer1_outputs(2211));
    layer2_outputs(981) <= '1';
    layer2_outputs(982) <= not(layer1_outputs(2990));
    layer2_outputs(983) <= layer1_outputs(4274);
    layer2_outputs(984) <= (layer1_outputs(4048)) and not (layer1_outputs(4772));
    layer2_outputs(985) <= (layer1_outputs(2713)) or (layer1_outputs(3497));
    layer2_outputs(986) <= layer1_outputs(4077);
    layer2_outputs(987) <= not(layer1_outputs(2013)) or (layer1_outputs(2698));
    layer2_outputs(988) <= not((layer1_outputs(918)) and (layer1_outputs(239)));
    layer2_outputs(989) <= not(layer1_outputs(1086)) or (layer1_outputs(636));
    layer2_outputs(990) <= not((layer1_outputs(843)) and (layer1_outputs(4393)));
    layer2_outputs(991) <= not((layer1_outputs(1093)) and (layer1_outputs(713)));
    layer2_outputs(992) <= not(layer1_outputs(3876)) or (layer1_outputs(4196));
    layer2_outputs(993) <= (layer1_outputs(4793)) or (layer1_outputs(1550));
    layer2_outputs(994) <= not(layer1_outputs(980)) or (layer1_outputs(4247));
    layer2_outputs(995) <= not(layer1_outputs(4285));
    layer2_outputs(996) <= (layer1_outputs(706)) and not (layer1_outputs(2173));
    layer2_outputs(997) <= not(layer1_outputs(4298));
    layer2_outputs(998) <= (layer1_outputs(1850)) and not (layer1_outputs(3206));
    layer2_outputs(999) <= '0';
    layer2_outputs(1000) <= not(layer1_outputs(704));
    layer2_outputs(1001) <= not((layer1_outputs(1451)) and (layer1_outputs(3182)));
    layer2_outputs(1002) <= not(layer1_outputs(4718)) or (layer1_outputs(508));
    layer2_outputs(1003) <= not((layer1_outputs(4696)) and (layer1_outputs(3135)));
    layer2_outputs(1004) <= layer1_outputs(3817);
    layer2_outputs(1005) <= '1';
    layer2_outputs(1006) <= not((layer1_outputs(2956)) and (layer1_outputs(3899)));
    layer2_outputs(1007) <= not(layer1_outputs(2426));
    layer2_outputs(1008) <= not(layer1_outputs(569)) or (layer1_outputs(63));
    layer2_outputs(1009) <= not(layer1_outputs(427));
    layer2_outputs(1010) <= (layer1_outputs(2931)) and not (layer1_outputs(891));
    layer2_outputs(1011) <= '0';
    layer2_outputs(1012) <= not(layer1_outputs(1361));
    layer2_outputs(1013) <= (layer1_outputs(4874)) and not (layer1_outputs(788));
    layer2_outputs(1014) <= not(layer1_outputs(2824));
    layer2_outputs(1015) <= not((layer1_outputs(823)) xor (layer1_outputs(4847)));
    layer2_outputs(1016) <= not(layer1_outputs(791)) or (layer1_outputs(2773));
    layer2_outputs(1017) <= not((layer1_outputs(566)) xor (layer1_outputs(2460)));
    layer2_outputs(1018) <= layer1_outputs(3837);
    layer2_outputs(1019) <= layer1_outputs(1450);
    layer2_outputs(1020) <= not(layer1_outputs(2064));
    layer2_outputs(1021) <= not(layer1_outputs(2517)) or (layer1_outputs(1373));
    layer2_outputs(1022) <= '1';
    layer2_outputs(1023) <= not(layer1_outputs(966)) or (layer1_outputs(515));
    layer2_outputs(1024) <= (layer1_outputs(3601)) and not (layer1_outputs(3841));
    layer2_outputs(1025) <= (layer1_outputs(1219)) and not (layer1_outputs(2829));
    layer2_outputs(1026) <= not(layer1_outputs(4410)) or (layer1_outputs(5064));
    layer2_outputs(1027) <= (layer1_outputs(5051)) or (layer1_outputs(3674));
    layer2_outputs(1028) <= not(layer1_outputs(2611)) or (layer1_outputs(299));
    layer2_outputs(1029) <= not(layer1_outputs(974));
    layer2_outputs(1030) <= (layer1_outputs(1340)) and not (layer1_outputs(1884));
    layer2_outputs(1031) <= not(layer1_outputs(3068)) or (layer1_outputs(893));
    layer2_outputs(1032) <= not(layer1_outputs(1130));
    layer2_outputs(1033) <= not(layer1_outputs(5102));
    layer2_outputs(1034) <= not((layer1_outputs(4769)) and (layer1_outputs(842)));
    layer2_outputs(1035) <= '0';
    layer2_outputs(1036) <= layer1_outputs(782);
    layer2_outputs(1037) <= layer1_outputs(3752);
    layer2_outputs(1038) <= not(layer1_outputs(4029)) or (layer1_outputs(1314));
    layer2_outputs(1039) <= not(layer1_outputs(400));
    layer2_outputs(1040) <= (layer1_outputs(2225)) and (layer1_outputs(4936));
    layer2_outputs(1041) <= (layer1_outputs(3622)) and not (layer1_outputs(3988));
    layer2_outputs(1042) <= layer1_outputs(4733);
    layer2_outputs(1043) <= (layer1_outputs(4433)) and not (layer1_outputs(4998));
    layer2_outputs(1044) <= layer1_outputs(998);
    layer2_outputs(1045) <= not(layer1_outputs(1157));
    layer2_outputs(1046) <= layer1_outputs(2734);
    layer2_outputs(1047) <= not(layer1_outputs(841)) or (layer1_outputs(3661));
    layer2_outputs(1048) <= '0';
    layer2_outputs(1049) <= not(layer1_outputs(5014));
    layer2_outputs(1050) <= not(layer1_outputs(2890));
    layer2_outputs(1051) <= (layer1_outputs(2011)) or (layer1_outputs(4516));
    layer2_outputs(1052) <= (layer1_outputs(1119)) and (layer1_outputs(4434));
    layer2_outputs(1053) <= layer1_outputs(758);
    layer2_outputs(1054) <= (layer1_outputs(3816)) and not (layer1_outputs(5000));
    layer2_outputs(1055) <= (layer1_outputs(2462)) and not (layer1_outputs(2485));
    layer2_outputs(1056) <= '1';
    layer2_outputs(1057) <= not(layer1_outputs(4223));
    layer2_outputs(1058) <= not(layer1_outputs(4388)) or (layer1_outputs(3514));
    layer2_outputs(1059) <= (layer1_outputs(1030)) and not (layer1_outputs(2479));
    layer2_outputs(1060) <= (layer1_outputs(1842)) and not (layer1_outputs(5043));
    layer2_outputs(1061) <= not(layer1_outputs(4576));
    layer2_outputs(1062) <= (layer1_outputs(4617)) and not (layer1_outputs(3048));
    layer2_outputs(1063) <= '1';
    layer2_outputs(1064) <= layer1_outputs(2174);
    layer2_outputs(1065) <= '0';
    layer2_outputs(1066) <= layer1_outputs(3931);
    layer2_outputs(1067) <= '1';
    layer2_outputs(1068) <= '0';
    layer2_outputs(1069) <= not(layer1_outputs(2237)) or (layer1_outputs(689));
    layer2_outputs(1070) <= layer1_outputs(2721);
    layer2_outputs(1071) <= layer1_outputs(2262);
    layer2_outputs(1072) <= layer1_outputs(4768);
    layer2_outputs(1073) <= not(layer1_outputs(3998));
    layer2_outputs(1074) <= (layer1_outputs(3488)) and not (layer1_outputs(239));
    layer2_outputs(1075) <= not((layer1_outputs(1485)) and (layer1_outputs(1807)));
    layer2_outputs(1076) <= layer1_outputs(1170);
    layer2_outputs(1077) <= layer1_outputs(3081);
    layer2_outputs(1078) <= layer1_outputs(2835);
    layer2_outputs(1079) <= not(layer1_outputs(1741)) or (layer1_outputs(3178));
    layer2_outputs(1080) <= '1';
    layer2_outputs(1081) <= not(layer1_outputs(4965)) or (layer1_outputs(256));
    layer2_outputs(1082) <= (layer1_outputs(4386)) and (layer1_outputs(4774));
    layer2_outputs(1083) <= not(layer1_outputs(5016));
    layer2_outputs(1084) <= layer1_outputs(3905);
    layer2_outputs(1085) <= not(layer1_outputs(4284));
    layer2_outputs(1086) <= not(layer1_outputs(3044));
    layer2_outputs(1087) <= (layer1_outputs(2928)) and (layer1_outputs(1612));
    layer2_outputs(1088) <= layer1_outputs(2547);
    layer2_outputs(1089) <= '0';
    layer2_outputs(1090) <= (layer1_outputs(3599)) and (layer1_outputs(464));
    layer2_outputs(1091) <= layer1_outputs(2731);
    layer2_outputs(1092) <= '0';
    layer2_outputs(1093) <= (layer1_outputs(2458)) and not (layer1_outputs(154));
    layer2_outputs(1094) <= '1';
    layer2_outputs(1095) <= layer1_outputs(3973);
    layer2_outputs(1096) <= layer1_outputs(3828);
    layer2_outputs(1097) <= '1';
    layer2_outputs(1098) <= not(layer1_outputs(1387)) or (layer1_outputs(1222));
    layer2_outputs(1099) <= (layer1_outputs(4228)) and not (layer1_outputs(3642));
    layer2_outputs(1100) <= not(layer1_outputs(3417)) or (layer1_outputs(4461));
    layer2_outputs(1101) <= layer1_outputs(1010);
    layer2_outputs(1102) <= not(layer1_outputs(1793));
    layer2_outputs(1103) <= (layer1_outputs(672)) and not (layer1_outputs(4807));
    layer2_outputs(1104) <= '0';
    layer2_outputs(1105) <= not((layer1_outputs(4152)) or (layer1_outputs(1872)));
    layer2_outputs(1106) <= not((layer1_outputs(3908)) or (layer1_outputs(508)));
    layer2_outputs(1107) <= not(layer1_outputs(4158)) or (layer1_outputs(1267));
    layer2_outputs(1108) <= not((layer1_outputs(3322)) xor (layer1_outputs(1932)));
    layer2_outputs(1109) <= '1';
    layer2_outputs(1110) <= not(layer1_outputs(3352)) or (layer1_outputs(2414));
    layer2_outputs(1111) <= not(layer1_outputs(4593));
    layer2_outputs(1112) <= (layer1_outputs(2665)) and not (layer1_outputs(4289));
    layer2_outputs(1113) <= not(layer1_outputs(3858)) or (layer1_outputs(3864));
    layer2_outputs(1114) <= (layer1_outputs(4456)) and not (layer1_outputs(2821));
    layer2_outputs(1115) <= not(layer1_outputs(937)) or (layer1_outputs(4087));
    layer2_outputs(1116) <= not((layer1_outputs(3719)) or (layer1_outputs(268)));
    layer2_outputs(1117) <= (layer1_outputs(2410)) xor (layer1_outputs(4964));
    layer2_outputs(1118) <= '1';
    layer2_outputs(1119) <= layer1_outputs(1960);
    layer2_outputs(1120) <= layer1_outputs(2618);
    layer2_outputs(1121) <= '0';
    layer2_outputs(1122) <= (layer1_outputs(3415)) or (layer1_outputs(4134));
    layer2_outputs(1123) <= '1';
    layer2_outputs(1124) <= not(layer1_outputs(4502));
    layer2_outputs(1125) <= (layer1_outputs(2365)) and not (layer1_outputs(2255));
    layer2_outputs(1126) <= not(layer1_outputs(3826));
    layer2_outputs(1127) <= not(layer1_outputs(2495)) or (layer1_outputs(1482));
    layer2_outputs(1128) <= layer1_outputs(344);
    layer2_outputs(1129) <= layer1_outputs(2019);
    layer2_outputs(1130) <= '1';
    layer2_outputs(1131) <= layer1_outputs(737);
    layer2_outputs(1132) <= not(layer1_outputs(567));
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= not(layer1_outputs(754));
    layer2_outputs(1135) <= not(layer1_outputs(2588));
    layer2_outputs(1136) <= layer1_outputs(1348);
    layer2_outputs(1137) <= not(layer1_outputs(4287)) or (layer1_outputs(4112));
    layer2_outputs(1138) <= not(layer1_outputs(2046)) or (layer1_outputs(1857));
    layer2_outputs(1139) <= not(layer1_outputs(2747));
    layer2_outputs(1140) <= not(layer1_outputs(1022));
    layer2_outputs(1141) <= (layer1_outputs(1976)) xor (layer1_outputs(642));
    layer2_outputs(1142) <= not(layer1_outputs(4271));
    layer2_outputs(1143) <= not(layer1_outputs(1822));
    layer2_outputs(1144) <= (layer1_outputs(4641)) xor (layer1_outputs(4929));
    layer2_outputs(1145) <= '0';
    layer2_outputs(1146) <= not(layer1_outputs(3276));
    layer2_outputs(1147) <= not(layer1_outputs(748));
    layer2_outputs(1148) <= not(layer1_outputs(1903)) or (layer1_outputs(1009));
    layer2_outputs(1149) <= not((layer1_outputs(157)) and (layer1_outputs(1855)));
    layer2_outputs(1150) <= layer1_outputs(1172);
    layer2_outputs(1151) <= layer1_outputs(3873);
    layer2_outputs(1152) <= '0';
    layer2_outputs(1153) <= not(layer1_outputs(88));
    layer2_outputs(1154) <= layer1_outputs(4503);
    layer2_outputs(1155) <= (layer1_outputs(1345)) and not (layer1_outputs(4268));
    layer2_outputs(1156) <= (layer1_outputs(4539)) and (layer1_outputs(1367));
    layer2_outputs(1157) <= not(layer1_outputs(115)) or (layer1_outputs(872));
    layer2_outputs(1158) <= '0';
    layer2_outputs(1159) <= (layer1_outputs(1757)) and (layer1_outputs(4672));
    layer2_outputs(1160) <= (layer1_outputs(2312)) and (layer1_outputs(155));
    layer2_outputs(1161) <= (layer1_outputs(3098)) and not (layer1_outputs(4252));
    layer2_outputs(1162) <= (layer1_outputs(3470)) or (layer1_outputs(4791));
    layer2_outputs(1163) <= not(layer1_outputs(2803));
    layer2_outputs(1164) <= (layer1_outputs(3988)) or (layer1_outputs(3999));
    layer2_outputs(1165) <= layer1_outputs(398);
    layer2_outputs(1166) <= not((layer1_outputs(3954)) or (layer1_outputs(2251)));
    layer2_outputs(1167) <= not((layer1_outputs(1138)) or (layer1_outputs(351)));
    layer2_outputs(1168) <= not((layer1_outputs(1159)) and (layer1_outputs(3366)));
    layer2_outputs(1169) <= (layer1_outputs(5113)) and not (layer1_outputs(464));
    layer2_outputs(1170) <= layer1_outputs(2080);
    layer2_outputs(1171) <= layer1_outputs(2157);
    layer2_outputs(1172) <= not((layer1_outputs(703)) and (layer1_outputs(3910)));
    layer2_outputs(1173) <= (layer1_outputs(3766)) and not (layer1_outputs(3112));
    layer2_outputs(1174) <= not((layer1_outputs(1692)) and (layer1_outputs(1272)));
    layer2_outputs(1175) <= not(layer1_outputs(2104));
    layer2_outputs(1176) <= not(layer1_outputs(1755)) or (layer1_outputs(2039));
    layer2_outputs(1177) <= not(layer1_outputs(898)) or (layer1_outputs(3912));
    layer2_outputs(1178) <= not((layer1_outputs(386)) or (layer1_outputs(3913)));
    layer2_outputs(1179) <= (layer1_outputs(2789)) and not (layer1_outputs(2196));
    layer2_outputs(1180) <= (layer1_outputs(1995)) and not (layer1_outputs(4996));
    layer2_outputs(1181) <= not((layer1_outputs(2657)) or (layer1_outputs(4675)));
    layer2_outputs(1182) <= layer1_outputs(1087);
    layer2_outputs(1183) <= layer1_outputs(3468);
    layer2_outputs(1184) <= layer1_outputs(1817);
    layer2_outputs(1185) <= (layer1_outputs(2236)) and not (layer1_outputs(1744));
    layer2_outputs(1186) <= (layer1_outputs(3659)) or (layer1_outputs(207));
    layer2_outputs(1187) <= layer1_outputs(4044);
    layer2_outputs(1188) <= layer1_outputs(1175);
    layer2_outputs(1189) <= not(layer1_outputs(4308));
    layer2_outputs(1190) <= (layer1_outputs(4673)) and not (layer1_outputs(3057));
    layer2_outputs(1191) <= '0';
    layer2_outputs(1192) <= layer1_outputs(2856);
    layer2_outputs(1193) <= '1';
    layer2_outputs(1194) <= not(layer1_outputs(3013));
    layer2_outputs(1195) <= '0';
    layer2_outputs(1196) <= (layer1_outputs(3460)) and not (layer1_outputs(3575));
    layer2_outputs(1197) <= (layer1_outputs(2519)) or (layer1_outputs(2173));
    layer2_outputs(1198) <= (layer1_outputs(1426)) and (layer1_outputs(834));
    layer2_outputs(1199) <= (layer1_outputs(2639)) and not (layer1_outputs(2607));
    layer2_outputs(1200) <= not((layer1_outputs(881)) or (layer1_outputs(2486)));
    layer2_outputs(1201) <= not(layer1_outputs(1266));
    layer2_outputs(1202) <= (layer1_outputs(3871)) or (layer1_outputs(4684));
    layer2_outputs(1203) <= not(layer1_outputs(3386));
    layer2_outputs(1204) <= not(layer1_outputs(1581)) or (layer1_outputs(3554));
    layer2_outputs(1205) <= layer1_outputs(4492);
    layer2_outputs(1206) <= (layer1_outputs(4052)) and not (layer1_outputs(3212));
    layer2_outputs(1207) <= not(layer1_outputs(2367)) or (layer1_outputs(2693));
    layer2_outputs(1208) <= layer1_outputs(3023);
    layer2_outputs(1209) <= '1';
    layer2_outputs(1210) <= (layer1_outputs(510)) and not (layer1_outputs(209));
    layer2_outputs(1211) <= (layer1_outputs(668)) and not (layer1_outputs(1742));
    layer2_outputs(1212) <= '0';
    layer2_outputs(1213) <= not(layer1_outputs(1656)) or (layer1_outputs(1979));
    layer2_outputs(1214) <= not((layer1_outputs(3954)) and (layer1_outputs(3483)));
    layer2_outputs(1215) <= not((layer1_outputs(4336)) or (layer1_outputs(4047)));
    layer2_outputs(1216) <= not((layer1_outputs(4011)) and (layer1_outputs(4808)));
    layer2_outputs(1217) <= not((layer1_outputs(4909)) or (layer1_outputs(970)));
    layer2_outputs(1218) <= not(layer1_outputs(3801));
    layer2_outputs(1219) <= (layer1_outputs(5061)) and (layer1_outputs(1538));
    layer2_outputs(1220) <= not(layer1_outputs(2847)) or (layer1_outputs(611));
    layer2_outputs(1221) <= not(layer1_outputs(3945));
    layer2_outputs(1222) <= layer1_outputs(517);
    layer2_outputs(1223) <= layer1_outputs(1104);
    layer2_outputs(1224) <= (layer1_outputs(4587)) or (layer1_outputs(3346));
    layer2_outputs(1225) <= not((layer1_outputs(4561)) or (layer1_outputs(3521)));
    layer2_outputs(1226) <= not(layer1_outputs(4985)) or (layer1_outputs(4592));
    layer2_outputs(1227) <= not(layer1_outputs(1829));
    layer2_outputs(1228) <= not((layer1_outputs(2187)) or (layer1_outputs(2587)));
    layer2_outputs(1229) <= (layer1_outputs(2719)) and not (layer1_outputs(1528));
    layer2_outputs(1230) <= not((layer1_outputs(649)) or (layer1_outputs(3719)));
    layer2_outputs(1231) <= not(layer1_outputs(1781));
    layer2_outputs(1232) <= not(layer1_outputs(793)) or (layer1_outputs(1237));
    layer2_outputs(1233) <= '0';
    layer2_outputs(1234) <= layer1_outputs(4238);
    layer2_outputs(1235) <= (layer1_outputs(1973)) and (layer1_outputs(3862));
    layer2_outputs(1236) <= '1';
    layer2_outputs(1237) <= '0';
    layer2_outputs(1238) <= layer1_outputs(4889);
    layer2_outputs(1239) <= not(layer1_outputs(1583));
    layer2_outputs(1240) <= '0';
    layer2_outputs(1241) <= (layer1_outputs(817)) and not (layer1_outputs(3820));
    layer2_outputs(1242) <= (layer1_outputs(4800)) and (layer1_outputs(3974));
    layer2_outputs(1243) <= '1';
    layer2_outputs(1244) <= not(layer1_outputs(1659)) or (layer1_outputs(3848));
    layer2_outputs(1245) <= (layer1_outputs(4520)) and not (layer1_outputs(1126));
    layer2_outputs(1246) <= layer1_outputs(2587);
    layer2_outputs(1247) <= (layer1_outputs(3778)) and not (layer1_outputs(535));
    layer2_outputs(1248) <= (layer1_outputs(2081)) or (layer1_outputs(866));
    layer2_outputs(1249) <= '0';
    layer2_outputs(1250) <= not((layer1_outputs(3360)) or (layer1_outputs(4033)));
    layer2_outputs(1251) <= (layer1_outputs(4381)) and (layer1_outputs(388));
    layer2_outputs(1252) <= (layer1_outputs(4058)) and (layer1_outputs(2162));
    layer2_outputs(1253) <= (layer1_outputs(97)) and not (layer1_outputs(1005));
    layer2_outputs(1254) <= (layer1_outputs(1616)) and (layer1_outputs(4985));
    layer2_outputs(1255) <= not(layer1_outputs(876));
    layer2_outputs(1256) <= not(layer1_outputs(3));
    layer2_outputs(1257) <= layer1_outputs(483);
    layer2_outputs(1258) <= layer1_outputs(1706);
    layer2_outputs(1259) <= not(layer1_outputs(4148));
    layer2_outputs(1260) <= not(layer1_outputs(323));
    layer2_outputs(1261) <= not((layer1_outputs(1781)) xor (layer1_outputs(2506)));
    layer2_outputs(1262) <= not(layer1_outputs(2697));
    layer2_outputs(1263) <= (layer1_outputs(1838)) and not (layer1_outputs(2868));
    layer2_outputs(1264) <= '1';
    layer2_outputs(1265) <= (layer1_outputs(2275)) and not (layer1_outputs(3105));
    layer2_outputs(1266) <= (layer1_outputs(1211)) and (layer1_outputs(4610));
    layer2_outputs(1267) <= not(layer1_outputs(971)) or (layer1_outputs(744));
    layer2_outputs(1268) <= not(layer1_outputs(1562)) or (layer1_outputs(226));
    layer2_outputs(1269) <= not(layer1_outputs(199)) or (layer1_outputs(2932));
    layer2_outputs(1270) <= layer1_outputs(3128);
    layer2_outputs(1271) <= (layer1_outputs(3713)) and (layer1_outputs(3306));
    layer2_outputs(1272) <= not(layer1_outputs(2621)) or (layer1_outputs(679));
    layer2_outputs(1273) <= not(layer1_outputs(5109)) or (layer1_outputs(2484));
    layer2_outputs(1274) <= layer1_outputs(537);
    layer2_outputs(1275) <= not((layer1_outputs(714)) or (layer1_outputs(2301)));
    layer2_outputs(1276) <= (layer1_outputs(2390)) and not (layer1_outputs(2574));
    layer2_outputs(1277) <= not((layer1_outputs(4523)) and (layer1_outputs(4483)));
    layer2_outputs(1278) <= not(layer1_outputs(2031));
    layer2_outputs(1279) <= '1';
    layer2_outputs(1280) <= (layer1_outputs(3482)) or (layer1_outputs(4292));
    layer2_outputs(1281) <= (layer1_outputs(2095)) or (layer1_outputs(1325));
    layer2_outputs(1282) <= not(layer1_outputs(53)) or (layer1_outputs(2304));
    layer2_outputs(1283) <= not(layer1_outputs(4521)) or (layer1_outputs(1125));
    layer2_outputs(1284) <= '0';
    layer2_outputs(1285) <= not(layer1_outputs(1892));
    layer2_outputs(1286) <= (layer1_outputs(1720)) and (layer1_outputs(2169));
    layer2_outputs(1287) <= '1';
    layer2_outputs(1288) <= (layer1_outputs(3648)) and not (layer1_outputs(2521));
    layer2_outputs(1289) <= not(layer1_outputs(3509)) or (layer1_outputs(4727));
    layer2_outputs(1290) <= not((layer1_outputs(2843)) or (layer1_outputs(3811)));
    layer2_outputs(1291) <= not(layer1_outputs(2442));
    layer2_outputs(1292) <= not(layer1_outputs(1203)) or (layer1_outputs(334));
    layer2_outputs(1293) <= not(layer1_outputs(3806)) or (layer1_outputs(128));
    layer2_outputs(1294) <= not(layer1_outputs(4042));
    layer2_outputs(1295) <= layer1_outputs(2387);
    layer2_outputs(1296) <= layer1_outputs(3522);
    layer2_outputs(1297) <= (layer1_outputs(2235)) or (layer1_outputs(1122));
    layer2_outputs(1298) <= not((layer1_outputs(1376)) and (layer1_outputs(1784)));
    layer2_outputs(1299) <= not((layer1_outputs(1073)) and (layer1_outputs(2808)));
    layer2_outputs(1300) <= not((layer1_outputs(1041)) and (layer1_outputs(4044)));
    layer2_outputs(1301) <= layer1_outputs(2787);
    layer2_outputs(1302) <= (layer1_outputs(1935)) or (layer1_outputs(4580));
    layer2_outputs(1303) <= layer1_outputs(600);
    layer2_outputs(1304) <= '1';
    layer2_outputs(1305) <= (layer1_outputs(5047)) or (layer1_outputs(4656));
    layer2_outputs(1306) <= '0';
    layer2_outputs(1307) <= layer1_outputs(182);
    layer2_outputs(1308) <= (layer1_outputs(1533)) and not (layer1_outputs(2220));
    layer2_outputs(1309) <= (layer1_outputs(3379)) and (layer1_outputs(2005));
    layer2_outputs(1310) <= '0';
    layer2_outputs(1311) <= not((layer1_outputs(2782)) and (layer1_outputs(3510)));
    layer2_outputs(1312) <= '1';
    layer2_outputs(1313) <= '0';
    layer2_outputs(1314) <= layer1_outputs(621);
    layer2_outputs(1315) <= not(layer1_outputs(4895));
    layer2_outputs(1316) <= (layer1_outputs(3059)) xor (layer1_outputs(2054));
    layer2_outputs(1317) <= '0';
    layer2_outputs(1318) <= '0';
    layer2_outputs(1319) <= not((layer1_outputs(4521)) and (layer1_outputs(3257)));
    layer2_outputs(1320) <= (layer1_outputs(828)) or (layer1_outputs(319));
    layer2_outputs(1321) <= not(layer1_outputs(2043)) or (layer1_outputs(819));
    layer2_outputs(1322) <= not(layer1_outputs(4184)) or (layer1_outputs(2538));
    layer2_outputs(1323) <= '1';
    layer2_outputs(1324) <= layer1_outputs(5033);
    layer2_outputs(1325) <= layer1_outputs(4809);
    layer2_outputs(1326) <= layer1_outputs(3924);
    layer2_outputs(1327) <= (layer1_outputs(4880)) or (layer1_outputs(2838));
    layer2_outputs(1328) <= '0';
    layer2_outputs(1329) <= '1';
    layer2_outputs(1330) <= (layer1_outputs(1613)) and (layer1_outputs(1202));
    layer2_outputs(1331) <= layer1_outputs(721);
    layer2_outputs(1332) <= layer1_outputs(4012);
    layer2_outputs(1333) <= not(layer1_outputs(3547));
    layer2_outputs(1334) <= '1';
    layer2_outputs(1335) <= (layer1_outputs(2299)) and not (layer1_outputs(5100));
    layer2_outputs(1336) <= '1';
    layer2_outputs(1337) <= (layer1_outputs(734)) and not (layer1_outputs(2401));
    layer2_outputs(1338) <= '1';
    layer2_outputs(1339) <= '1';
    layer2_outputs(1340) <= not(layer1_outputs(541));
    layer2_outputs(1341) <= (layer1_outputs(4473)) and not (layer1_outputs(203));
    layer2_outputs(1342) <= not(layer1_outputs(3803)) or (layer1_outputs(1334));
    layer2_outputs(1343) <= not(layer1_outputs(4296)) or (layer1_outputs(3257));
    layer2_outputs(1344) <= (layer1_outputs(1621)) and not (layer1_outputs(1105));
    layer2_outputs(1345) <= '1';
    layer2_outputs(1346) <= not(layer1_outputs(2546));
    layer2_outputs(1347) <= (layer1_outputs(2320)) and not (layer1_outputs(155));
    layer2_outputs(1348) <= (layer1_outputs(4212)) and not (layer1_outputs(1620));
    layer2_outputs(1349) <= (layer1_outputs(4486)) and (layer1_outputs(1400));
    layer2_outputs(1350) <= (layer1_outputs(346)) and not (layer1_outputs(321));
    layer2_outputs(1351) <= '1';
    layer2_outputs(1352) <= '0';
    layer2_outputs(1353) <= layer1_outputs(2818);
    layer2_outputs(1354) <= not(layer1_outputs(2930));
    layer2_outputs(1355) <= layer1_outputs(4398);
    layer2_outputs(1356) <= not(layer1_outputs(425));
    layer2_outputs(1357) <= layer1_outputs(3709);
    layer2_outputs(1358) <= not(layer1_outputs(227)) or (layer1_outputs(3243));
    layer2_outputs(1359) <= not(layer1_outputs(2949));
    layer2_outputs(1360) <= not(layer1_outputs(698)) or (layer1_outputs(1119));
    layer2_outputs(1361) <= not((layer1_outputs(3868)) xor (layer1_outputs(4599)));
    layer2_outputs(1362) <= not(layer1_outputs(4360)) or (layer1_outputs(775));
    layer2_outputs(1363) <= (layer1_outputs(4321)) or (layer1_outputs(1953));
    layer2_outputs(1364) <= (layer1_outputs(3463)) and (layer1_outputs(383));
    layer2_outputs(1365) <= not(layer1_outputs(2865)) or (layer1_outputs(2888));
    layer2_outputs(1366) <= not(layer1_outputs(3655));
    layer2_outputs(1367) <= (layer1_outputs(275)) and not (layer1_outputs(4437));
    layer2_outputs(1368) <= not(layer1_outputs(3134)) or (layer1_outputs(2701));
    layer2_outputs(1369) <= not(layer1_outputs(389)) or (layer1_outputs(3426));
    layer2_outputs(1370) <= not(layer1_outputs(3399)) or (layer1_outputs(4205));
    layer2_outputs(1371) <= layer1_outputs(1631);
    layer2_outputs(1372) <= not((layer1_outputs(2375)) and (layer1_outputs(4973)));
    layer2_outputs(1373) <= (layer1_outputs(381)) and (layer1_outputs(2455));
    layer2_outputs(1374) <= not(layer1_outputs(1730));
    layer2_outputs(1375) <= layer1_outputs(4716);
    layer2_outputs(1376) <= not(layer1_outputs(908)) or (layer1_outputs(4777));
    layer2_outputs(1377) <= not((layer1_outputs(3923)) or (layer1_outputs(1799)));
    layer2_outputs(1378) <= (layer1_outputs(4277)) or (layer1_outputs(4611));
    layer2_outputs(1379) <= '1';
    layer2_outputs(1380) <= '0';
    layer2_outputs(1381) <= '1';
    layer2_outputs(1382) <= not(layer1_outputs(3582)) or (layer1_outputs(2508));
    layer2_outputs(1383) <= (layer1_outputs(4325)) or (layer1_outputs(4498));
    layer2_outputs(1384) <= '1';
    layer2_outputs(1385) <= (layer1_outputs(3121)) and not (layer1_outputs(225));
    layer2_outputs(1386) <= layer1_outputs(2494);
    layer2_outputs(1387) <= not(layer1_outputs(3501));
    layer2_outputs(1388) <= not(layer1_outputs(2777));
    layer2_outputs(1389) <= not(layer1_outputs(785));
    layer2_outputs(1390) <= (layer1_outputs(1894)) and not (layer1_outputs(2841));
    layer2_outputs(1391) <= '1';
    layer2_outputs(1392) <= not((layer1_outputs(5046)) and (layer1_outputs(3168)));
    layer2_outputs(1393) <= (layer1_outputs(2012)) and not (layer1_outputs(3128));
    layer2_outputs(1394) <= '0';
    layer2_outputs(1395) <= layer1_outputs(4536);
    layer2_outputs(1396) <= not(layer1_outputs(1977));
    layer2_outputs(1397) <= layer1_outputs(4927);
    layer2_outputs(1398) <= layer1_outputs(3750);
    layer2_outputs(1399) <= layer1_outputs(3557);
    layer2_outputs(1400) <= layer1_outputs(3209);
    layer2_outputs(1401) <= (layer1_outputs(4016)) or (layer1_outputs(4624));
    layer2_outputs(1402) <= not(layer1_outputs(3656));
    layer2_outputs(1403) <= not((layer1_outputs(4162)) and (layer1_outputs(2497)));
    layer2_outputs(1404) <= not(layer1_outputs(2066));
    layer2_outputs(1405) <= (layer1_outputs(3185)) or (layer1_outputs(68));
    layer2_outputs(1406) <= not((layer1_outputs(1253)) and (layer1_outputs(2617)));
    layer2_outputs(1407) <= '0';
    layer2_outputs(1408) <= not(layer1_outputs(3160));
    layer2_outputs(1409) <= not(layer1_outputs(2027));
    layer2_outputs(1410) <= not(layer1_outputs(2889));
    layer2_outputs(1411) <= not((layer1_outputs(3452)) and (layer1_outputs(3870)));
    layer2_outputs(1412) <= (layer1_outputs(2562)) and (layer1_outputs(3927));
    layer2_outputs(1413) <= (layer1_outputs(1161)) and not (layer1_outputs(3823));
    layer2_outputs(1414) <= not(layer1_outputs(2731)) or (layer1_outputs(1459));
    layer2_outputs(1415) <= not(layer1_outputs(2833)) or (layer1_outputs(678));
    layer2_outputs(1416) <= (layer1_outputs(3299)) or (layer1_outputs(5057));
    layer2_outputs(1417) <= (layer1_outputs(1893)) and not (layer1_outputs(2091));
    layer2_outputs(1418) <= not((layer1_outputs(2350)) or (layer1_outputs(3272)));
    layer2_outputs(1419) <= not(layer1_outputs(722));
    layer2_outputs(1420) <= layer1_outputs(3476);
    layer2_outputs(1421) <= '0';
    layer2_outputs(1422) <= not(layer1_outputs(2897));
    layer2_outputs(1423) <= not(layer1_outputs(2315));
    layer2_outputs(1424) <= '1';
    layer2_outputs(1425) <= layer1_outputs(4419);
    layer2_outputs(1426) <= not(layer1_outputs(4384)) or (layer1_outputs(1987));
    layer2_outputs(1427) <= layer1_outputs(3340);
    layer2_outputs(1428) <= not(layer1_outputs(3180)) or (layer1_outputs(4179));
    layer2_outputs(1429) <= not((layer1_outputs(4028)) or (layer1_outputs(2988)));
    layer2_outputs(1430) <= (layer1_outputs(2711)) and (layer1_outputs(2824));
    layer2_outputs(1431) <= layer1_outputs(117);
    layer2_outputs(1432) <= '0';
    layer2_outputs(1433) <= (layer1_outputs(2312)) and (layer1_outputs(1181));
    layer2_outputs(1434) <= (layer1_outputs(5040)) and not (layer1_outputs(992));
    layer2_outputs(1435) <= not(layer1_outputs(2370));
    layer2_outputs(1436) <= not((layer1_outputs(2717)) and (layer1_outputs(2877)));
    layer2_outputs(1437) <= layer1_outputs(2327);
    layer2_outputs(1438) <= layer1_outputs(1383);
    layer2_outputs(1439) <= not(layer1_outputs(2747));
    layer2_outputs(1440) <= '0';
    layer2_outputs(1441) <= (layer1_outputs(2757)) and not (layer1_outputs(930));
    layer2_outputs(1442) <= '0';
    layer2_outputs(1443) <= layer1_outputs(4914);
    layer2_outputs(1444) <= not(layer1_outputs(2222));
    layer2_outputs(1445) <= not(layer1_outputs(2910));
    layer2_outputs(1446) <= not(layer1_outputs(1582));
    layer2_outputs(1447) <= not(layer1_outputs(3384)) or (layer1_outputs(1346));
    layer2_outputs(1448) <= (layer1_outputs(2281)) and not (layer1_outputs(639));
    layer2_outputs(1449) <= '1';
    layer2_outputs(1450) <= (layer1_outputs(646)) and not (layer1_outputs(4901));
    layer2_outputs(1451) <= not((layer1_outputs(12)) and (layer1_outputs(434)));
    layer2_outputs(1452) <= '1';
    layer2_outputs(1453) <= '1';
    layer2_outputs(1454) <= not(layer1_outputs(773));
    layer2_outputs(1455) <= (layer1_outputs(346)) and (layer1_outputs(2802));
    layer2_outputs(1456) <= '1';
    layer2_outputs(1457) <= not((layer1_outputs(413)) or (layer1_outputs(117)));
    layer2_outputs(1458) <= (layer1_outputs(1038)) and not (layer1_outputs(2683));
    layer2_outputs(1459) <= not((layer1_outputs(2500)) and (layer1_outputs(638)));
    layer2_outputs(1460) <= (layer1_outputs(2954)) and not (layer1_outputs(402));
    layer2_outputs(1461) <= (layer1_outputs(3405)) or (layer1_outputs(4516));
    layer2_outputs(1462) <= not((layer1_outputs(4837)) and (layer1_outputs(1228)));
    layer2_outputs(1463) <= (layer1_outputs(4408)) or (layer1_outputs(4600));
    layer2_outputs(1464) <= not(layer1_outputs(649)) or (layer1_outputs(2146));
    layer2_outputs(1465) <= layer1_outputs(180);
    layer2_outputs(1466) <= (layer1_outputs(4942)) xor (layer1_outputs(2481));
    layer2_outputs(1467) <= not(layer1_outputs(2015)) or (layer1_outputs(2592));
    layer2_outputs(1468) <= not(layer1_outputs(3560)) or (layer1_outputs(4735));
    layer2_outputs(1469) <= not(layer1_outputs(2112));
    layer2_outputs(1470) <= not((layer1_outputs(2308)) and (layer1_outputs(3033)));
    layer2_outputs(1471) <= not((layer1_outputs(243)) and (layer1_outputs(3189)));
    layer2_outputs(1472) <= not((layer1_outputs(813)) and (layer1_outputs(1059)));
    layer2_outputs(1473) <= not(layer1_outputs(2825));
    layer2_outputs(1474) <= (layer1_outputs(1981)) or (layer1_outputs(1213));
    layer2_outputs(1475) <= not(layer1_outputs(2345));
    layer2_outputs(1476) <= layer1_outputs(1180);
    layer2_outputs(1477) <= not(layer1_outputs(4779));
    layer2_outputs(1478) <= (layer1_outputs(2477)) and not (layer1_outputs(2981));
    layer2_outputs(1479) <= not(layer1_outputs(2831)) or (layer1_outputs(1903));
    layer2_outputs(1480) <= (layer1_outputs(1003)) and (layer1_outputs(1381));
    layer2_outputs(1481) <= not(layer1_outputs(4838));
    layer2_outputs(1482) <= '1';
    layer2_outputs(1483) <= '0';
    layer2_outputs(1484) <= not(layer1_outputs(4167)) or (layer1_outputs(4984));
    layer2_outputs(1485) <= not(layer1_outputs(3630));
    layer2_outputs(1486) <= '1';
    layer2_outputs(1487) <= not((layer1_outputs(625)) or (layer1_outputs(511)));
    layer2_outputs(1488) <= (layer1_outputs(686)) and (layer1_outputs(121));
    layer2_outputs(1489) <= not(layer1_outputs(393)) or (layer1_outputs(2976));
    layer2_outputs(1490) <= '0';
    layer2_outputs(1491) <= not((layer1_outputs(311)) or (layer1_outputs(1369)));
    layer2_outputs(1492) <= not(layer1_outputs(1543));
    layer2_outputs(1493) <= '0';
    layer2_outputs(1494) <= '1';
    layer2_outputs(1495) <= not((layer1_outputs(2421)) or (layer1_outputs(1841)));
    layer2_outputs(1496) <= (layer1_outputs(4940)) or (layer1_outputs(1478));
    layer2_outputs(1497) <= (layer1_outputs(3205)) and not (layer1_outputs(1785));
    layer2_outputs(1498) <= not(layer1_outputs(1418)) or (layer1_outputs(3985));
    layer2_outputs(1499) <= (layer1_outputs(1282)) and not (layer1_outputs(1196));
    layer2_outputs(1500) <= layer1_outputs(3316);
    layer2_outputs(1501) <= not(layer1_outputs(2290)) or (layer1_outputs(2806));
    layer2_outputs(1502) <= not(layer1_outputs(3531));
    layer2_outputs(1503) <= not((layer1_outputs(1860)) and (layer1_outputs(2120)));
    layer2_outputs(1504) <= (layer1_outputs(4146)) and not (layer1_outputs(4218));
    layer2_outputs(1505) <= not(layer1_outputs(75)) or (layer1_outputs(3457));
    layer2_outputs(1506) <= not(layer1_outputs(1998)) or (layer1_outputs(4132));
    layer2_outputs(1507) <= not((layer1_outputs(2436)) or (layer1_outputs(1251)));
    layer2_outputs(1508) <= not(layer1_outputs(4706));
    layer2_outputs(1509) <= '1';
    layer2_outputs(1510) <= not(layer1_outputs(2985));
    layer2_outputs(1511) <= not((layer1_outputs(3410)) and (layer1_outputs(2913)));
    layer2_outputs(1512) <= not(layer1_outputs(2296));
    layer2_outputs(1513) <= not(layer1_outputs(3037)) or (layer1_outputs(4105));
    layer2_outputs(1514) <= layer1_outputs(3782);
    layer2_outputs(1515) <= not(layer1_outputs(290));
    layer2_outputs(1516) <= layer1_outputs(3269);
    layer2_outputs(1517) <= '1';
    layer2_outputs(1518) <= layer1_outputs(3169);
    layer2_outputs(1519) <= (layer1_outputs(1423)) and not (layer1_outputs(438));
    layer2_outputs(1520) <= not((layer1_outputs(3142)) and (layer1_outputs(4704)));
    layer2_outputs(1521) <= '1';
    layer2_outputs(1522) <= not((layer1_outputs(2955)) and (layer1_outputs(4424)));
    layer2_outputs(1523) <= not((layer1_outputs(2151)) and (layer1_outputs(490)));
    layer2_outputs(1524) <= not((layer1_outputs(1147)) and (layer1_outputs(1437)));
    layer2_outputs(1525) <= not(layer1_outputs(2976));
    layer2_outputs(1526) <= layer1_outputs(2065);
    layer2_outputs(1527) <= layer1_outputs(1455);
    layer2_outputs(1528) <= not(layer1_outputs(873));
    layer2_outputs(1529) <= layer1_outputs(697);
    layer2_outputs(1530) <= not((layer1_outputs(3109)) and (layer1_outputs(3483)));
    layer2_outputs(1531) <= not((layer1_outputs(4066)) or (layer1_outputs(807)));
    layer2_outputs(1532) <= not((layer1_outputs(1017)) or (layer1_outputs(3434)));
    layer2_outputs(1533) <= layer1_outputs(2283);
    layer2_outputs(1534) <= layer1_outputs(4616);
    layer2_outputs(1535) <= (layer1_outputs(204)) or (layer1_outputs(2108));
    layer2_outputs(1536) <= not(layer1_outputs(795)) or (layer1_outputs(2020));
    layer2_outputs(1537) <= layer1_outputs(4579);
    layer2_outputs(1538) <= not(layer1_outputs(2244));
    layer2_outputs(1539) <= '0';
    layer2_outputs(1540) <= not(layer1_outputs(1515)) or (layer1_outputs(2093));
    layer2_outputs(1541) <= not((layer1_outputs(2991)) and (layer1_outputs(2713)));
    layer2_outputs(1542) <= (layer1_outputs(4123)) and (layer1_outputs(3395));
    layer2_outputs(1543) <= not((layer1_outputs(3034)) or (layer1_outputs(3344)));
    layer2_outputs(1544) <= not((layer1_outputs(1368)) or (layer1_outputs(4548)));
    layer2_outputs(1545) <= not(layer1_outputs(3736));
    layer2_outputs(1546) <= layer1_outputs(4173);
    layer2_outputs(1547) <= not(layer1_outputs(1081)) or (layer1_outputs(3951));
    layer2_outputs(1548) <= '1';
    layer2_outputs(1549) <= not((layer1_outputs(2646)) and (layer1_outputs(4645)));
    layer2_outputs(1550) <= layer1_outputs(5091);
    layer2_outputs(1551) <= (layer1_outputs(2217)) xor (layer1_outputs(3453));
    layer2_outputs(1552) <= '0';
    layer2_outputs(1553) <= (layer1_outputs(2776)) and not (layer1_outputs(1796));
    layer2_outputs(1554) <= not(layer1_outputs(460));
    layer2_outputs(1555) <= layer1_outputs(4846);
    layer2_outputs(1556) <= not(layer1_outputs(2961));
    layer2_outputs(1557) <= '0';
    layer2_outputs(1558) <= not(layer1_outputs(60)) or (layer1_outputs(2175));
    layer2_outputs(1559) <= layer1_outputs(3141);
    layer2_outputs(1560) <= '1';
    layer2_outputs(1561) <= layer1_outputs(158);
    layer2_outputs(1562) <= (layer1_outputs(161)) and (layer1_outputs(2763));
    layer2_outputs(1563) <= not((layer1_outputs(784)) or (layer1_outputs(1506)));
    layer2_outputs(1564) <= not(layer1_outputs(4273));
    layer2_outputs(1565) <= not(layer1_outputs(3414));
    layer2_outputs(1566) <= not((layer1_outputs(4236)) and (layer1_outputs(3416)));
    layer2_outputs(1567) <= (layer1_outputs(1440)) and not (layer1_outputs(4820));
    layer2_outputs(1568) <= (layer1_outputs(4566)) and not (layer1_outputs(1222));
    layer2_outputs(1569) <= not(layer1_outputs(3870));
    layer2_outputs(1570) <= not((layer1_outputs(1057)) or (layer1_outputs(2921)));
    layer2_outputs(1571) <= not(layer1_outputs(3632));
    layer2_outputs(1572) <= layer1_outputs(4338);
    layer2_outputs(1573) <= (layer1_outputs(4113)) xor (layer1_outputs(2330));
    layer2_outputs(1574) <= not(layer1_outputs(1375));
    layer2_outputs(1575) <= not(layer1_outputs(3804)) or (layer1_outputs(1777));
    layer2_outputs(1576) <= not(layer1_outputs(1847)) or (layer1_outputs(2810));
    layer2_outputs(1577) <= not(layer1_outputs(4647));
    layer2_outputs(1578) <= not(layer1_outputs(1172));
    layer2_outputs(1579) <= '1';
    layer2_outputs(1580) <= layer1_outputs(84);
    layer2_outputs(1581) <= not(layer1_outputs(4759));
    layer2_outputs(1582) <= (layer1_outputs(1694)) or (layer1_outputs(254));
    layer2_outputs(1583) <= not(layer1_outputs(2682)) or (layer1_outputs(497));
    layer2_outputs(1584) <= layer1_outputs(3798);
    layer2_outputs(1585) <= not(layer1_outputs(1515)) or (layer1_outputs(2537));
    layer2_outputs(1586) <= not(layer1_outputs(2965));
    layer2_outputs(1587) <= not(layer1_outputs(2035));
    layer2_outputs(1588) <= not(layer1_outputs(4751));
    layer2_outputs(1589) <= '1';
    layer2_outputs(1590) <= not((layer1_outputs(4805)) and (layer1_outputs(5094)));
    layer2_outputs(1591) <= not((layer1_outputs(3802)) and (layer1_outputs(806)));
    layer2_outputs(1592) <= layer1_outputs(1629);
    layer2_outputs(1593) <= not(layer1_outputs(4606)) or (layer1_outputs(945));
    layer2_outputs(1594) <= (layer1_outputs(3550)) and (layer1_outputs(623));
    layer2_outputs(1595) <= not(layer1_outputs(3782)) or (layer1_outputs(46));
    layer2_outputs(1596) <= not(layer1_outputs(3035));
    layer2_outputs(1597) <= not(layer1_outputs(3082)) or (layer1_outputs(629));
    layer2_outputs(1598) <= (layer1_outputs(2653)) and not (layer1_outputs(3155));
    layer2_outputs(1599) <= (layer1_outputs(2585)) xor (layer1_outputs(1925));
    layer2_outputs(1600) <= '0';
    layer2_outputs(1601) <= not(layer1_outputs(1762)) or (layer1_outputs(2311));
    layer2_outputs(1602) <= layer1_outputs(3810);
    layer2_outputs(1603) <= not(layer1_outputs(896)) or (layer1_outputs(3545));
    layer2_outputs(1604) <= not(layer1_outputs(3423));
    layer2_outputs(1605) <= not(layer1_outputs(2463));
    layer2_outputs(1606) <= '1';
    layer2_outputs(1607) <= (layer1_outputs(1779)) and (layer1_outputs(3948));
    layer2_outputs(1608) <= layer1_outputs(3487);
    layer2_outputs(1609) <= '0';
    layer2_outputs(1610) <= not(layer1_outputs(941));
    layer2_outputs(1611) <= not(layer1_outputs(2603)) or (layer1_outputs(4162));
    layer2_outputs(1612) <= not((layer1_outputs(1239)) or (layer1_outputs(2440)));
    layer2_outputs(1613) <= '0';
    layer2_outputs(1614) <= layer1_outputs(813);
    layer2_outputs(1615) <= layer1_outputs(2114);
    layer2_outputs(1616) <= not(layer1_outputs(4414));
    layer2_outputs(1617) <= not(layer1_outputs(4954));
    layer2_outputs(1618) <= (layer1_outputs(3195)) or (layer1_outputs(3525));
    layer2_outputs(1619) <= not(layer1_outputs(337)) or (layer1_outputs(2586));
    layer2_outputs(1620) <= not(layer1_outputs(3304));
    layer2_outputs(1621) <= (layer1_outputs(3129)) and not (layer1_outputs(4266));
    layer2_outputs(1622) <= not(layer1_outputs(2705));
    layer2_outputs(1623) <= '1';
    layer2_outputs(1624) <= layer1_outputs(170);
    layer2_outputs(1625) <= layer1_outputs(1501);
    layer2_outputs(1626) <= not(layer1_outputs(2968));
    layer2_outputs(1627) <= '0';
    layer2_outputs(1628) <= not((layer1_outputs(1509)) or (layer1_outputs(1953)));
    layer2_outputs(1629) <= not(layer1_outputs(4003)) or (layer1_outputs(2470));
    layer2_outputs(1630) <= not(layer1_outputs(462));
    layer2_outputs(1631) <= '1';
    layer2_outputs(1632) <= not(layer1_outputs(2786)) or (layer1_outputs(33));
    layer2_outputs(1633) <= (layer1_outputs(1504)) and not (layer1_outputs(3787));
    layer2_outputs(1634) <= not((layer1_outputs(4129)) or (layer1_outputs(275)));
    layer2_outputs(1635) <= (layer1_outputs(1141)) and not (layer1_outputs(955));
    layer2_outputs(1636) <= not(layer1_outputs(163));
    layer2_outputs(1637) <= layer1_outputs(153);
    layer2_outputs(1638) <= '1';
    layer2_outputs(1639) <= layer1_outputs(215);
    layer2_outputs(1640) <= not((layer1_outputs(3102)) or (layer1_outputs(85)));
    layer2_outputs(1641) <= (layer1_outputs(4387)) and not (layer1_outputs(4801));
    layer2_outputs(1642) <= not(layer1_outputs(4319));
    layer2_outputs(1643) <= (layer1_outputs(1324)) or (layer1_outputs(2882));
    layer2_outputs(1644) <= not(layer1_outputs(4128));
    layer2_outputs(1645) <= (layer1_outputs(4368)) and not (layer1_outputs(409));
    layer2_outputs(1646) <= (layer1_outputs(4019)) xor (layer1_outputs(3593));
    layer2_outputs(1647) <= not((layer1_outputs(4673)) or (layer1_outputs(2662)));
    layer2_outputs(1648) <= layer1_outputs(29);
    layer2_outputs(1649) <= (layer1_outputs(2516)) and not (layer1_outputs(531));
    layer2_outputs(1650) <= not(layer1_outputs(1142)) or (layer1_outputs(641));
    layer2_outputs(1651) <= not((layer1_outputs(3014)) or (layer1_outputs(1703)));
    layer2_outputs(1652) <= not(layer1_outputs(1862));
    layer2_outputs(1653) <= not(layer1_outputs(3363));
    layer2_outputs(1654) <= not((layer1_outputs(863)) or (layer1_outputs(4004)));
    layer2_outputs(1655) <= not(layer1_outputs(2189));
    layer2_outputs(1656) <= not(layer1_outputs(1569)) or (layer1_outputs(3259));
    layer2_outputs(1657) <= not(layer1_outputs(3456)) or (layer1_outputs(4945));
    layer2_outputs(1658) <= not(layer1_outputs(3646));
    layer2_outputs(1659) <= not(layer1_outputs(3041)) or (layer1_outputs(5099));
    layer2_outputs(1660) <= '0';
    layer2_outputs(1661) <= not(layer1_outputs(4879));
    layer2_outputs(1662) <= (layer1_outputs(3174)) and (layer1_outputs(4372));
    layer2_outputs(1663) <= not(layer1_outputs(2669));
    layer2_outputs(1664) <= (layer1_outputs(4914)) or (layer1_outputs(4121));
    layer2_outputs(1665) <= '0';
    layer2_outputs(1666) <= (layer1_outputs(916)) and not (layer1_outputs(1191));
    layer2_outputs(1667) <= (layer1_outputs(4346)) xor (layer1_outputs(4461));
    layer2_outputs(1668) <= (layer1_outputs(4591)) or (layer1_outputs(1431));
    layer2_outputs(1669) <= layer1_outputs(2902);
    layer2_outputs(1670) <= '1';
    layer2_outputs(1671) <= (layer1_outputs(3610)) and not (layer1_outputs(3691));
    layer2_outputs(1672) <= not((layer1_outputs(2817)) and (layer1_outputs(2941)));
    layer2_outputs(1673) <= not(layer1_outputs(1505));
    layer2_outputs(1674) <= (layer1_outputs(1306)) or (layer1_outputs(2068));
    layer2_outputs(1675) <= not((layer1_outputs(2745)) and (layer1_outputs(2388)));
    layer2_outputs(1676) <= (layer1_outputs(1604)) and not (layer1_outputs(1167));
    layer2_outputs(1677) <= not((layer1_outputs(2198)) and (layer1_outputs(4891)));
    layer2_outputs(1678) <= (layer1_outputs(591)) and (layer1_outputs(2550));
    layer2_outputs(1679) <= not((layer1_outputs(3696)) and (layer1_outputs(906)));
    layer2_outputs(1680) <= not(layer1_outputs(1291));
    layer2_outputs(1681) <= not(layer1_outputs(2014));
    layer2_outputs(1682) <= not(layer1_outputs(4541));
    layer2_outputs(1683) <= (layer1_outputs(182)) and not (layer1_outputs(2523));
    layer2_outputs(1684) <= not((layer1_outputs(4147)) and (layer1_outputs(1313)));
    layer2_outputs(1685) <= not((layer1_outputs(1888)) or (layer1_outputs(4505)));
    layer2_outputs(1686) <= (layer1_outputs(2753)) and not (layer1_outputs(4227));
    layer2_outputs(1687) <= not(layer1_outputs(4508));
    layer2_outputs(1688) <= not(layer1_outputs(1576));
    layer2_outputs(1689) <= '0';
    layer2_outputs(1690) <= (layer1_outputs(1960)) and not (layer1_outputs(3253));
    layer2_outputs(1691) <= '0';
    layer2_outputs(1692) <= (layer1_outputs(3091)) and (layer1_outputs(4628));
    layer2_outputs(1693) <= layer1_outputs(1188);
    layer2_outputs(1694) <= not(layer1_outputs(457)) or (layer1_outputs(3240));
    layer2_outputs(1695) <= (layer1_outputs(3305)) and (layer1_outputs(4416));
    layer2_outputs(1696) <= layer1_outputs(1580);
    layer2_outputs(1697) <= not(layer1_outputs(2655));
    layer2_outputs(1698) <= not((layer1_outputs(4652)) and (layer1_outputs(3580)));
    layer2_outputs(1699) <= '0';
    layer2_outputs(1700) <= (layer1_outputs(4181)) and not (layer1_outputs(1552));
    layer2_outputs(1701) <= (layer1_outputs(3502)) and (layer1_outputs(4737));
    layer2_outputs(1702) <= not((layer1_outputs(1206)) and (layer1_outputs(3598)));
    layer2_outputs(1703) <= layer1_outputs(2206);
    layer2_outputs(1704) <= not(layer1_outputs(3943));
    layer2_outputs(1705) <= (layer1_outputs(1428)) or (layer1_outputs(3022));
    layer2_outputs(1706) <= not(layer1_outputs(4810)) or (layer1_outputs(577));
    layer2_outputs(1707) <= not(layer1_outputs(507));
    layer2_outputs(1708) <= (layer1_outputs(4622)) and not (layer1_outputs(3214));
    layer2_outputs(1709) <= layer1_outputs(4687);
    layer2_outputs(1710) <= (layer1_outputs(1814)) and not (layer1_outputs(4149));
    layer2_outputs(1711) <= '1';
    layer2_outputs(1712) <= (layer1_outputs(2998)) and not (layer1_outputs(4840));
    layer2_outputs(1713) <= '0';
    layer2_outputs(1714) <= not(layer1_outputs(517));
    layer2_outputs(1715) <= (layer1_outputs(4010)) and not (layer1_outputs(4112));
    layer2_outputs(1716) <= not(layer1_outputs(3249));
    layer2_outputs(1717) <= not(layer1_outputs(1148));
    layer2_outputs(1718) <= not(layer1_outputs(98)) or (layer1_outputs(1265));
    layer2_outputs(1719) <= layer1_outputs(4171);
    layer2_outputs(1720) <= not((layer1_outputs(2998)) and (layer1_outputs(5091)));
    layer2_outputs(1721) <= not(layer1_outputs(4440));
    layer2_outputs(1722) <= not(layer1_outputs(3274));
    layer2_outputs(1723) <= '1';
    layer2_outputs(1724) <= not((layer1_outputs(4263)) or (layer1_outputs(4320)));
    layer2_outputs(1725) <= '1';
    layer2_outputs(1726) <= (layer1_outputs(1856)) or (layer1_outputs(167));
    layer2_outputs(1727) <= '0';
    layer2_outputs(1728) <= not(layer1_outputs(4379)) or (layer1_outputs(4586));
    layer2_outputs(1729) <= not(layer1_outputs(3524)) or (layer1_outputs(489));
    layer2_outputs(1730) <= not((layer1_outputs(5001)) and (layer1_outputs(3481)));
    layer2_outputs(1731) <= (layer1_outputs(3722)) and not (layer1_outputs(3632));
    layer2_outputs(1732) <= not((layer1_outputs(3011)) or (layer1_outputs(1391)));
    layer2_outputs(1733) <= '0';
    layer2_outputs(1734) <= (layer1_outputs(1300)) and (layer1_outputs(3908));
    layer2_outputs(1735) <= not(layer1_outputs(8)) or (layer1_outputs(4910));
    layer2_outputs(1736) <= not((layer1_outputs(3509)) and (layer1_outputs(2985)));
    layer2_outputs(1737) <= (layer1_outputs(4324)) or (layer1_outputs(1495));
    layer2_outputs(1738) <= '0';
    layer2_outputs(1739) <= layer1_outputs(1577);
    layer2_outputs(1740) <= not((layer1_outputs(2832)) or (layer1_outputs(2366)));
    layer2_outputs(1741) <= not(layer1_outputs(1723));
    layer2_outputs(1742) <= not(layer1_outputs(1136));
    layer2_outputs(1743) <= not((layer1_outputs(4554)) or (layer1_outputs(3620)));
    layer2_outputs(1744) <= (layer1_outputs(2518)) and not (layer1_outputs(3708));
    layer2_outputs(1745) <= '0';
    layer2_outputs(1746) <= not(layer1_outputs(4705)) or (layer1_outputs(193));
    layer2_outputs(1747) <= (layer1_outputs(2365)) and (layer1_outputs(1343));
    layer2_outputs(1748) <= '0';
    layer2_outputs(1749) <= not(layer1_outputs(1818));
    layer2_outputs(1750) <= not(layer1_outputs(1556));
    layer2_outputs(1751) <= not(layer1_outputs(3390)) or (layer1_outputs(1831));
    layer2_outputs(1752) <= layer1_outputs(1862);
    layer2_outputs(1753) <= (layer1_outputs(3444)) and not (layer1_outputs(1890));
    layer2_outputs(1754) <= not(layer1_outputs(4761));
    layer2_outputs(1755) <= not(layer1_outputs(595));
    layer2_outputs(1756) <= layer1_outputs(2295);
    layer2_outputs(1757) <= not(layer1_outputs(1348));
    layer2_outputs(1758) <= layer1_outputs(765);
    layer2_outputs(1759) <= (layer1_outputs(1873)) or (layer1_outputs(2842));
    layer2_outputs(1760) <= not(layer1_outputs(616)) or (layer1_outputs(2651));
    layer2_outputs(1761) <= not(layer1_outputs(1143)) or (layer1_outputs(3978));
    layer2_outputs(1762) <= '1';
    layer2_outputs(1763) <= layer1_outputs(4854);
    layer2_outputs(1764) <= not(layer1_outputs(2160));
    layer2_outputs(1765) <= not(layer1_outputs(2057));
    layer2_outputs(1766) <= (layer1_outputs(1859)) xor (layer1_outputs(3218));
    layer2_outputs(1767) <= not((layer1_outputs(2307)) or (layer1_outputs(1067)));
    layer2_outputs(1768) <= not(layer1_outputs(4785));
    layer2_outputs(1769) <= not(layer1_outputs(3982));
    layer2_outputs(1770) <= '1';
    layer2_outputs(1771) <= '1';
    layer2_outputs(1772) <= '0';
    layer2_outputs(1773) <= layer1_outputs(4970);
    layer2_outputs(1774) <= not(layer1_outputs(3717));
    layer2_outputs(1775) <= (layer1_outputs(2788)) and not (layer1_outputs(3338));
    layer2_outputs(1776) <= not((layer1_outputs(55)) and (layer1_outputs(3096)));
    layer2_outputs(1777) <= layer1_outputs(96);
    layer2_outputs(1778) <= not(layer1_outputs(1896));
    layer2_outputs(1779) <= '1';
    layer2_outputs(1780) <= '1';
    layer2_outputs(1781) <= '1';
    layer2_outputs(1782) <= (layer1_outputs(1585)) and (layer1_outputs(3186));
    layer2_outputs(1783) <= not((layer1_outputs(571)) and (layer1_outputs(1691)));
    layer2_outputs(1784) <= (layer1_outputs(3157)) or (layer1_outputs(3256));
    layer2_outputs(1785) <= '0';
    layer2_outputs(1786) <= (layer1_outputs(1584)) and not (layer1_outputs(1008));
    layer2_outputs(1787) <= (layer1_outputs(639)) or (layer1_outputs(3608));
    layer2_outputs(1788) <= not(layer1_outputs(347));
    layer2_outputs(1789) <= layer1_outputs(4448);
    layer2_outputs(1790) <= '1';
    layer2_outputs(1791) <= layer1_outputs(1352);
    layer2_outputs(1792) <= not((layer1_outputs(3122)) and (layer1_outputs(627)));
    layer2_outputs(1793) <= not(layer1_outputs(1330));
    layer2_outputs(1794) <= (layer1_outputs(4350)) or (layer1_outputs(3695));
    layer2_outputs(1795) <= layer1_outputs(4222);
    layer2_outputs(1796) <= layer1_outputs(1292);
    layer2_outputs(1797) <= not((layer1_outputs(3123)) or (layer1_outputs(1020)));
    layer2_outputs(1798) <= not((layer1_outputs(2601)) and (layer1_outputs(40)));
    layer2_outputs(1799) <= not(layer1_outputs(2809)) or (layer1_outputs(894));
    layer2_outputs(1800) <= layer1_outputs(176);
    layer2_outputs(1801) <= not((layer1_outputs(3836)) and (layer1_outputs(4642)));
    layer2_outputs(1802) <= not(layer1_outputs(159));
    layer2_outputs(1803) <= '1';
    layer2_outputs(1804) <= '1';
    layer2_outputs(1805) <= not(layer1_outputs(4496));
    layer2_outputs(1806) <= '0';
    layer2_outputs(1807) <= not(layer1_outputs(1719)) or (layer1_outputs(4989));
    layer2_outputs(1808) <= (layer1_outputs(2475)) xor (layer1_outputs(2215));
    layer2_outputs(1809) <= not((layer1_outputs(2860)) and (layer1_outputs(4865)));
    layer2_outputs(1810) <= layer1_outputs(4587);
    layer2_outputs(1811) <= (layer1_outputs(2178)) xor (layer1_outputs(3371));
    layer2_outputs(1812) <= not(layer1_outputs(101));
    layer2_outputs(1813) <= not(layer1_outputs(3573));
    layer2_outputs(1814) <= not(layer1_outputs(4391)) or (layer1_outputs(3963));
    layer2_outputs(1815) <= layer1_outputs(5020);
    layer2_outputs(1816) <= layer1_outputs(3278);
    layer2_outputs(1817) <= '0';
    layer2_outputs(1818) <= not(layer1_outputs(4883));
    layer2_outputs(1819) <= not(layer1_outputs(1051));
    layer2_outputs(1820) <= (layer1_outputs(2555)) and not (layer1_outputs(3306));
    layer2_outputs(1821) <= not(layer1_outputs(325)) or (layer1_outputs(2786));
    layer2_outputs(1822) <= not((layer1_outputs(2863)) or (layer1_outputs(2211)));
    layer2_outputs(1823) <= '0';
    layer2_outputs(1824) <= '0';
    layer2_outputs(1825) <= not((layer1_outputs(861)) and (layer1_outputs(4170)));
    layer2_outputs(1826) <= '1';
    layer2_outputs(1827) <= '1';
    layer2_outputs(1828) <= not((layer1_outputs(385)) and (layer1_outputs(421)));
    layer2_outputs(1829) <= (layer1_outputs(1519)) or (layer1_outputs(2106));
    layer2_outputs(1830) <= layer1_outputs(4866);
    layer2_outputs(1831) <= layer1_outputs(1322);
    layer2_outputs(1832) <= not(layer1_outputs(4370)) or (layer1_outputs(1358));
    layer2_outputs(1833) <= not(layer1_outputs(1941));
    layer2_outputs(1834) <= not((layer1_outputs(825)) or (layer1_outputs(1068)));
    layer2_outputs(1835) <= layer1_outputs(2560);
    layer2_outputs(1836) <= not(layer1_outputs(3473));
    layer2_outputs(1837) <= layer1_outputs(1722);
    layer2_outputs(1838) <= (layer1_outputs(3361)) and (layer1_outputs(4269));
    layer2_outputs(1839) <= layer1_outputs(1615);
    layer2_outputs(1840) <= (layer1_outputs(3910)) and not (layer1_outputs(1609));
    layer2_outputs(1841) <= not((layer1_outputs(3984)) and (layer1_outputs(2686)));
    layer2_outputs(1842) <= not((layer1_outputs(437)) and (layer1_outputs(2505)));
    layer2_outputs(1843) <= layer1_outputs(143);
    layer2_outputs(1844) <= layer1_outputs(5);
    layer2_outputs(1845) <= not(layer1_outputs(1689));
    layer2_outputs(1846) <= layer1_outputs(236);
    layer2_outputs(1847) <= '1';
    layer2_outputs(1848) <= (layer1_outputs(3935)) and not (layer1_outputs(2115));
    layer2_outputs(1849) <= (layer1_outputs(274)) and not (layer1_outputs(2432));
    layer2_outputs(1850) <= layer1_outputs(2224);
    layer2_outputs(1851) <= layer1_outputs(4725);
    layer2_outputs(1852) <= '0';
    layer2_outputs(1853) <= (layer1_outputs(3154)) or (layer1_outputs(3851));
    layer2_outputs(1854) <= not((layer1_outputs(1521)) and (layer1_outputs(4435)));
    layer2_outputs(1855) <= (layer1_outputs(3469)) and (layer1_outputs(4260));
    layer2_outputs(1856) <= not((layer1_outputs(4049)) or (layer1_outputs(1412)));
    layer2_outputs(1857) <= (layer1_outputs(1219)) and (layer1_outputs(3101));
    layer2_outputs(1858) <= (layer1_outputs(2013)) and not (layer1_outputs(5094));
    layer2_outputs(1859) <= layer1_outputs(1442);
    layer2_outputs(1860) <= not(layer1_outputs(4032));
    layer2_outputs(1861) <= layer1_outputs(1380);
    layer2_outputs(1862) <= '0';
    layer2_outputs(1863) <= '0';
    layer2_outputs(1864) <= not(layer1_outputs(39));
    layer2_outputs(1865) <= (layer1_outputs(936)) or (layer1_outputs(2386));
    layer2_outputs(1866) <= not((layer1_outputs(1236)) and (layer1_outputs(2655)));
    layer2_outputs(1867) <= not(layer1_outputs(1431)) or (layer1_outputs(1164));
    layer2_outputs(1868) <= '1';
    layer2_outputs(1869) <= layer1_outputs(4953);
    layer2_outputs(1870) <= not(layer1_outputs(2272)) or (layer1_outputs(2203));
    layer2_outputs(1871) <= (layer1_outputs(3244)) and not (layer1_outputs(530));
    layer2_outputs(1872) <= not(layer1_outputs(2181));
    layer2_outputs(1873) <= layer1_outputs(2477);
    layer2_outputs(1874) <= '1';
    layer2_outputs(1875) <= not(layer1_outputs(902));
    layer2_outputs(1876) <= not((layer1_outputs(3589)) and (layer1_outputs(1127)));
    layer2_outputs(1877) <= (layer1_outputs(13)) and (layer1_outputs(2480));
    layer2_outputs(1878) <= (layer1_outputs(2873)) and not (layer1_outputs(4579));
    layer2_outputs(1879) <= layer1_outputs(242);
    layer2_outputs(1880) <= '1';
    layer2_outputs(1881) <= not((layer1_outputs(2355)) and (layer1_outputs(186)));
    layer2_outputs(1882) <= '1';
    layer2_outputs(1883) <= '0';
    layer2_outputs(1884) <= layer1_outputs(183);
    layer2_outputs(1885) <= '1';
    layer2_outputs(1886) <= layer1_outputs(242);
    layer2_outputs(1887) <= layer1_outputs(1939);
    layer2_outputs(1888) <= (layer1_outputs(1715)) and not (layer1_outputs(865));
    layer2_outputs(1889) <= not((layer1_outputs(2732)) or (layer1_outputs(1150)));
    layer2_outputs(1890) <= layer1_outputs(4200);
    layer2_outputs(1891) <= '0';
    layer2_outputs(1892) <= not(layer1_outputs(4944)) or (layer1_outputs(3261));
    layer2_outputs(1893) <= (layer1_outputs(664)) xor (layer1_outputs(1899));
    layer2_outputs(1894) <= '1';
    layer2_outputs(1895) <= '0';
    layer2_outputs(1896) <= not(layer1_outputs(3793)) or (layer1_outputs(2199));
    layer2_outputs(1897) <= (layer1_outputs(113)) and not (layer1_outputs(4919));
    layer2_outputs(1898) <= not(layer1_outputs(3996));
    layer2_outputs(1899) <= not(layer1_outputs(21)) or (layer1_outputs(630));
    layer2_outputs(1900) <= (layer1_outputs(4059)) or (layer1_outputs(251));
    layer2_outputs(1901) <= not(layer1_outputs(3831));
    layer2_outputs(1902) <= (layer1_outputs(414)) and not (layer1_outputs(4793));
    layer2_outputs(1903) <= '0';
    layer2_outputs(1904) <= layer1_outputs(811);
    layer2_outputs(1905) <= not(layer1_outputs(4974)) or (layer1_outputs(4043));
    layer2_outputs(1906) <= not(layer1_outputs(472)) or (layer1_outputs(2907));
    layer2_outputs(1907) <= (layer1_outputs(3881)) and not (layer1_outputs(1002));
    layer2_outputs(1908) <= '1';
    layer2_outputs(1909) <= '1';
    layer2_outputs(1910) <= not(layer1_outputs(968));
    layer2_outputs(1911) <= not(layer1_outputs(2450)) or (layer1_outputs(4537));
    layer2_outputs(1912) <= layer1_outputs(2554);
    layer2_outputs(1913) <= layer1_outputs(134);
    layer2_outputs(1914) <= (layer1_outputs(2400)) and not (layer1_outputs(4336));
    layer2_outputs(1915) <= not(layer1_outputs(2256));
    layer2_outputs(1916) <= '0';
    layer2_outputs(1917) <= not((layer1_outputs(3339)) and (layer1_outputs(2018)));
    layer2_outputs(1918) <= not((layer1_outputs(3333)) xor (layer1_outputs(770)));
    layer2_outputs(1919) <= not((layer1_outputs(1225)) and (layer1_outputs(3903)));
    layer2_outputs(1920) <= not(layer1_outputs(4257)) or (layer1_outputs(4466));
    layer2_outputs(1921) <= layer1_outputs(750);
    layer2_outputs(1922) <= (layer1_outputs(4313)) and not (layer1_outputs(2834));
    layer2_outputs(1923) <= layer1_outputs(4094);
    layer2_outputs(1924) <= layer1_outputs(4430);
    layer2_outputs(1925) <= not((layer1_outputs(352)) or (layer1_outputs(26)));
    layer2_outputs(1926) <= not(layer1_outputs(3149));
    layer2_outputs(1927) <= not((layer1_outputs(2332)) or (layer1_outputs(2328)));
    layer2_outputs(1928) <= not(layer1_outputs(3667));
    layer2_outputs(1929) <= not((layer1_outputs(1562)) and (layer1_outputs(1436)));
    layer2_outputs(1930) <= (layer1_outputs(4772)) and not (layer1_outputs(1687));
    layer2_outputs(1931) <= (layer1_outputs(3236)) xor (layer1_outputs(3289));
    layer2_outputs(1932) <= layer1_outputs(3894);
    layer2_outputs(1933) <= (layer1_outputs(4314)) or (layer1_outputs(3424));
    layer2_outputs(1934) <= '0';
    layer2_outputs(1935) <= not((layer1_outputs(1906)) and (layer1_outputs(1018)));
    layer2_outputs(1936) <= not(layer1_outputs(4411)) or (layer1_outputs(5075));
    layer2_outputs(1937) <= not(layer1_outputs(329));
    layer2_outputs(1938) <= not((layer1_outputs(4802)) or (layer1_outputs(3047)));
    layer2_outputs(1939) <= layer1_outputs(3698);
    layer2_outputs(1940) <= not(layer1_outputs(3901));
    layer2_outputs(1941) <= not(layer1_outputs(1720)) or (layer1_outputs(3705));
    layer2_outputs(1942) <= layer1_outputs(4293);
    layer2_outputs(1943) <= not(layer1_outputs(5059)) or (layer1_outputs(3472));
    layer2_outputs(1944) <= layer1_outputs(1902);
    layer2_outputs(1945) <= (layer1_outputs(1877)) and not (layer1_outputs(5090));
    layer2_outputs(1946) <= not((layer1_outputs(1714)) and (layer1_outputs(995)));
    layer2_outputs(1947) <= '0';
    layer2_outputs(1948) <= not(layer1_outputs(2548)) or (layer1_outputs(4761));
    layer2_outputs(1949) <= layer1_outputs(2958);
    layer2_outputs(1950) <= (layer1_outputs(3681)) and not (layer1_outputs(499));
    layer2_outputs(1951) <= layer1_outputs(2050);
    layer2_outputs(1952) <= not(layer1_outputs(124));
    layer2_outputs(1953) <= '0';
    layer2_outputs(1954) <= (layer1_outputs(1827)) and (layer1_outputs(1946));
    layer2_outputs(1955) <= not(layer1_outputs(318)) or (layer1_outputs(2110));
    layer2_outputs(1956) <= not(layer1_outputs(4815)) or (layer1_outputs(2348));
    layer2_outputs(1957) <= not(layer1_outputs(3223)) or (layer1_outputs(4282));
    layer2_outputs(1958) <= layer1_outputs(3431);
    layer2_outputs(1959) <= layer1_outputs(2837);
    layer2_outputs(1960) <= not(layer1_outputs(4006));
    layer2_outputs(1961) <= layer1_outputs(3755);
    layer2_outputs(1962) <= layer1_outputs(3576);
    layer2_outputs(1963) <= not(layer1_outputs(1938)) or (layer1_outputs(2203));
    layer2_outputs(1964) <= '1';
    layer2_outputs(1965) <= not(layer1_outputs(2858)) or (layer1_outputs(4770));
    layer2_outputs(1966) <= '0';
    layer2_outputs(1967) <= layer1_outputs(4947);
    layer2_outputs(1968) <= layer1_outputs(4046);
    layer2_outputs(1969) <= not((layer1_outputs(4406)) and (layer1_outputs(2294)));
    layer2_outputs(1970) <= layer1_outputs(1361);
    layer2_outputs(1971) <= not(layer1_outputs(370)) or (layer1_outputs(4621));
    layer2_outputs(1972) <= '0';
    layer2_outputs(1973) <= not(layer1_outputs(3315));
    layer2_outputs(1974) <= not(layer1_outputs(4006)) or (layer1_outputs(1538));
    layer2_outputs(1975) <= (layer1_outputs(4527)) and (layer1_outputs(3757));
    layer2_outputs(1976) <= layer1_outputs(2584);
    layer2_outputs(1977) <= (layer1_outputs(3513)) and not (layer1_outputs(1919));
    layer2_outputs(1978) <= (layer1_outputs(877)) and not (layer1_outputs(3002));
    layer2_outputs(1979) <= (layer1_outputs(1337)) and not (layer1_outputs(4287));
    layer2_outputs(1980) <= not(layer1_outputs(1975));
    layer2_outputs(1981) <= not(layer1_outputs(381));
    layer2_outputs(1982) <= (layer1_outputs(2861)) and (layer1_outputs(3060));
    layer2_outputs(1983) <= not((layer1_outputs(2182)) or (layer1_outputs(3209)));
    layer2_outputs(1984) <= (layer1_outputs(2182)) and not (layer1_outputs(4071));
    layer2_outputs(1985) <= '0';
    layer2_outputs(1986) <= layer1_outputs(3898);
    layer2_outputs(1987) <= not(layer1_outputs(3559)) or (layer1_outputs(1601));
    layer2_outputs(1988) <= '1';
    layer2_outputs(1989) <= not(layer1_outputs(1411));
    layer2_outputs(1990) <= (layer1_outputs(1630)) and (layer1_outputs(3466));
    layer2_outputs(1991) <= not((layer1_outputs(942)) or (layer1_outputs(4402)));
    layer2_outputs(1992) <= layer1_outputs(409);
    layer2_outputs(1993) <= (layer1_outputs(447)) and not (layer1_outputs(3428));
    layer2_outputs(1994) <= (layer1_outputs(371)) and not (layer1_outputs(885));
    layer2_outputs(1995) <= layer1_outputs(2535);
    layer2_outputs(1996) <= not(layer1_outputs(2933)) or (layer1_outputs(2635));
    layer2_outputs(1997) <= not(layer1_outputs(4486)) or (layer1_outputs(1927));
    layer2_outputs(1998) <= layer1_outputs(1427);
    layer2_outputs(1999) <= layer1_outputs(5085);
    layer2_outputs(2000) <= not(layer1_outputs(3246)) or (layer1_outputs(1712));
    layer2_outputs(2001) <= not(layer1_outputs(1487));
    layer2_outputs(2002) <= '1';
    layer2_outputs(2003) <= not(layer1_outputs(13));
    layer2_outputs(2004) <= (layer1_outputs(3672)) and not (layer1_outputs(2346));
    layer2_outputs(2005) <= layer1_outputs(2303);
    layer2_outputs(2006) <= not((layer1_outputs(1929)) and (layer1_outputs(1412)));
    layer2_outputs(2007) <= (layer1_outputs(1509)) and (layer1_outputs(468));
    layer2_outputs(2008) <= (layer1_outputs(4428)) and not (layer1_outputs(1175));
    layer2_outputs(2009) <= not(layer1_outputs(3061));
    layer2_outputs(2010) <= (layer1_outputs(1686)) and not (layer1_outputs(115));
    layer2_outputs(2011) <= layer1_outputs(727);
    layer2_outputs(2012) <= not(layer1_outputs(4406)) or (layer1_outputs(397));
    layer2_outputs(2013) <= not(layer1_outputs(224));
    layer2_outputs(2014) <= not(layer1_outputs(2740)) or (layer1_outputs(4416));
    layer2_outputs(2015) <= not((layer1_outputs(3475)) and (layer1_outputs(4969)));
    layer2_outputs(2016) <= '0';
    layer2_outputs(2017) <= not(layer1_outputs(1272)) or (layer1_outputs(4798));
    layer2_outputs(2018) <= layer1_outputs(1311);
    layer2_outputs(2019) <= not((layer1_outputs(3850)) or (layer1_outputs(3946)));
    layer2_outputs(2020) <= not(layer1_outputs(637));
    layer2_outputs(2021) <= (layer1_outputs(4446)) and not (layer1_outputs(5078));
    layer2_outputs(2022) <= not(layer1_outputs(468));
    layer2_outputs(2023) <= not(layer1_outputs(4110));
    layer2_outputs(2024) <= not(layer1_outputs(2598)) or (layer1_outputs(5080));
    layer2_outputs(2025) <= (layer1_outputs(633)) and not (layer1_outputs(2178));
    layer2_outputs(2026) <= not((layer1_outputs(2094)) or (layer1_outputs(3001)));
    layer2_outputs(2027) <= not(layer1_outputs(4366)) or (layer1_outputs(1871));
    layer2_outputs(2028) <= not(layer1_outputs(2077)) or (layer1_outputs(3769));
    layer2_outputs(2029) <= (layer1_outputs(3902)) xor (layer1_outputs(3161));
    layer2_outputs(2030) <= (layer1_outputs(3593)) and not (layer1_outputs(1103));
    layer2_outputs(2031) <= not(layer1_outputs(829));
    layer2_outputs(2032) <= layer1_outputs(653);
    layer2_outputs(2033) <= (layer1_outputs(3349)) and (layer1_outputs(3038));
    layer2_outputs(2034) <= not(layer1_outputs(378)) or (layer1_outputs(2513));
    layer2_outputs(2035) <= '1';
    layer2_outputs(2036) <= not((layer1_outputs(1844)) and (layer1_outputs(497)));
    layer2_outputs(2037) <= layer1_outputs(3465);
    layer2_outputs(2038) <= (layer1_outputs(1761)) or (layer1_outputs(193));
    layer2_outputs(2039) <= not(layer1_outputs(342));
    layer2_outputs(2040) <= not(layer1_outputs(3500));
    layer2_outputs(2041) <= not((layer1_outputs(179)) and (layer1_outputs(3190)));
    layer2_outputs(2042) <= (layer1_outputs(866)) and not (layer1_outputs(2806));
    layer2_outputs(2043) <= not((layer1_outputs(617)) and (layer1_outputs(646)));
    layer2_outputs(2044) <= not(layer1_outputs(228)) or (layer1_outputs(1821));
    layer2_outputs(2045) <= '1';
    layer2_outputs(2046) <= layer1_outputs(2467);
    layer2_outputs(2047) <= '0';
    layer2_outputs(2048) <= (layer1_outputs(334)) and not (layer1_outputs(4103));
    layer2_outputs(2049) <= not(layer1_outputs(3592));
    layer2_outputs(2050) <= '0';
    layer2_outputs(2051) <= '1';
    layer2_outputs(2052) <= '0';
    layer2_outputs(2053) <= layer1_outputs(222);
    layer2_outputs(2054) <= not((layer1_outputs(1283)) or (layer1_outputs(31)));
    layer2_outputs(2055) <= '1';
    layer2_outputs(2056) <= not(layer1_outputs(225)) or (layer1_outputs(2001));
    layer2_outputs(2057) <= '1';
    layer2_outputs(2058) <= not((layer1_outputs(4450)) and (layer1_outputs(305)));
    layer2_outputs(2059) <= not((layer1_outputs(5068)) or (layer1_outputs(1295)));
    layer2_outputs(2060) <= not((layer1_outputs(4144)) and (layer1_outputs(3039)));
    layer2_outputs(2061) <= '1';
    layer2_outputs(2062) <= layer1_outputs(1594);
    layer2_outputs(2063) <= not(layer1_outputs(4377));
    layer2_outputs(2064) <= (layer1_outputs(2643)) and not (layer1_outputs(79));
    layer2_outputs(2065) <= '1';
    layer2_outputs(2066) <= '0';
    layer2_outputs(2067) <= (layer1_outputs(3436)) and (layer1_outputs(2912));
    layer2_outputs(2068) <= layer1_outputs(5019);
    layer2_outputs(2069) <= layer1_outputs(224);
    layer2_outputs(2070) <= '1';
    layer2_outputs(2071) <= layer1_outputs(92);
    layer2_outputs(2072) <= (layer1_outputs(2901)) and not (layer1_outputs(3964));
    layer2_outputs(2073) <= layer1_outputs(3878);
    layer2_outputs(2074) <= not(layer1_outputs(3528));
    layer2_outputs(2075) <= not(layer1_outputs(3762)) or (layer1_outputs(4992));
    layer2_outputs(2076) <= not(layer1_outputs(3038)) or (layer1_outputs(421));
    layer2_outputs(2077) <= (layer1_outputs(3432)) and not (layer1_outputs(3980));
    layer2_outputs(2078) <= layer1_outputs(1162);
    layer2_outputs(2079) <= '1';
    layer2_outputs(2080) <= layer1_outputs(892);
    layer2_outputs(2081) <= '0';
    layer2_outputs(2082) <= not(layer1_outputs(3529)) or (layer1_outputs(3300));
    layer2_outputs(2083) <= not(layer1_outputs(156)) or (layer1_outputs(4711));
    layer2_outputs(2084) <= (layer1_outputs(3189)) or (layer1_outputs(291));
    layer2_outputs(2085) <= (layer1_outputs(5056)) or (layer1_outputs(4478));
    layer2_outputs(2086) <= not(layer1_outputs(2242));
    layer2_outputs(2087) <= layer1_outputs(4143);
    layer2_outputs(2088) <= (layer1_outputs(4168)) and (layer1_outputs(2045));
    layer2_outputs(2089) <= not((layer1_outputs(789)) or (layer1_outputs(2205)));
    layer2_outputs(2090) <= (layer1_outputs(595)) and (layer1_outputs(1837));
    layer2_outputs(2091) <= (layer1_outputs(3685)) and (layer1_outputs(3704));
    layer2_outputs(2092) <= not((layer1_outputs(2032)) or (layer1_outputs(3126)));
    layer2_outputs(2093) <= not((layer1_outputs(1807)) and (layer1_outputs(1392)));
    layer2_outputs(2094) <= not(layer1_outputs(1463));
    layer2_outputs(2095) <= not(layer1_outputs(3493)) or (layer1_outputs(976));
    layer2_outputs(2096) <= '0';
    layer2_outputs(2097) <= layer1_outputs(804);
    layer2_outputs(2098) <= (layer1_outputs(1864)) and not (layer1_outputs(569));
    layer2_outputs(2099) <= layer1_outputs(3132);
    layer2_outputs(2100) <= '1';
    layer2_outputs(2101) <= (layer1_outputs(4832)) and not (layer1_outputs(3605));
    layer2_outputs(2102) <= not(layer1_outputs(4949));
    layer2_outputs(2103) <= (layer1_outputs(3107)) or (layer1_outputs(2343));
    layer2_outputs(2104) <= not((layer1_outputs(4307)) or (layer1_outputs(897)));
    layer2_outputs(2105) <= (layer1_outputs(5053)) and not (layer1_outputs(3021));
    layer2_outputs(2106) <= '0';
    layer2_outputs(2107) <= (layer1_outputs(4476)) and (layer1_outputs(2233));
    layer2_outputs(2108) <= (layer1_outputs(1934)) and not (layer1_outputs(1617));
    layer2_outputs(2109) <= not(layer1_outputs(4884));
    layer2_outputs(2110) <= '1';
    layer2_outputs(2111) <= not(layer1_outputs(2780));
    layer2_outputs(2112) <= layer1_outputs(756);
    layer2_outputs(2113) <= not(layer1_outputs(2781));
    layer2_outputs(2114) <= (layer1_outputs(3588)) and (layer1_outputs(3453));
    layer2_outputs(2115) <= (layer1_outputs(873)) and (layer1_outputs(154));
    layer2_outputs(2116) <= not(layer1_outputs(3768)) or (layer1_outputs(2648));
    layer2_outputs(2117) <= (layer1_outputs(2402)) and not (layer1_outputs(2249));
    layer2_outputs(2118) <= layer1_outputs(717);
    layer2_outputs(2119) <= (layer1_outputs(1875)) or (layer1_outputs(1608));
    layer2_outputs(2120) <= not((layer1_outputs(3921)) or (layer1_outputs(925)));
    layer2_outputs(2121) <= (layer1_outputs(4823)) and (layer1_outputs(2487));
    layer2_outputs(2122) <= not(layer1_outputs(2901)) or (layer1_outputs(492));
    layer2_outputs(2123) <= (layer1_outputs(1739)) and not (layer1_outputs(3203));
    layer2_outputs(2124) <= not(layer1_outputs(2278)) or (layer1_outputs(892));
    layer2_outputs(2125) <= '1';
    layer2_outputs(2126) <= layer1_outputs(4297);
    layer2_outputs(2127) <= (layer1_outputs(5035)) or (layer1_outputs(2700));
    layer2_outputs(2128) <= '1';
    layer2_outputs(2129) <= not(layer1_outputs(705));
    layer2_outputs(2130) <= not(layer1_outputs(1954)) or (layer1_outputs(3391));
    layer2_outputs(2131) <= not((layer1_outputs(118)) or (layer1_outputs(482)));
    layer2_outputs(2132) <= not(layer1_outputs(3176));
    layer2_outputs(2133) <= not(layer1_outputs(353)) or (layer1_outputs(4002));
    layer2_outputs(2134) <= not(layer1_outputs(2574));
    layer2_outputs(2135) <= not((layer1_outputs(4958)) and (layer1_outputs(3814)));
    layer2_outputs(2136) <= (layer1_outputs(4721)) and not (layer1_outputs(2624));
    layer2_outputs(2137) <= not((layer1_outputs(374)) and (layer1_outputs(2722)));
    layer2_outputs(2138) <= not(layer1_outputs(2542));
    layer2_outputs(2139) <= not(layer1_outputs(404));
    layer2_outputs(2140) <= not(layer1_outputs(1417)) or (layer1_outputs(5000));
    layer2_outputs(2141) <= not(layer1_outputs(1894));
    layer2_outputs(2142) <= not(layer1_outputs(4542));
    layer2_outputs(2143) <= not(layer1_outputs(1156));
    layer2_outputs(2144) <= not(layer1_outputs(1038));
    layer2_outputs(2145) <= layer1_outputs(4130);
    layer2_outputs(2146) <= (layer1_outputs(2279)) or (layer1_outputs(2735));
    layer2_outputs(2147) <= not(layer1_outputs(4042)) or (layer1_outputs(3009));
    layer2_outputs(2148) <= not(layer1_outputs(4014)) or (layer1_outputs(461));
    layer2_outputs(2149) <= (layer1_outputs(2305)) or (layer1_outputs(165));
    layer2_outputs(2150) <= (layer1_outputs(652)) and not (layer1_outputs(406));
    layer2_outputs(2151) <= '0';
    layer2_outputs(2152) <= layer1_outputs(232);
    layer2_outputs(2153) <= not(layer1_outputs(423)) or (layer1_outputs(230));
    layer2_outputs(2154) <= not((layer1_outputs(145)) and (layer1_outputs(4518)));
    layer2_outputs(2155) <= layer1_outputs(3754);
    layer2_outputs(2156) <= '1';
    layer2_outputs(2157) <= layer1_outputs(1795);
    layer2_outputs(2158) <= '0';
    layer2_outputs(2159) <= (layer1_outputs(1323)) and not (layer1_outputs(3853));
    layer2_outputs(2160) <= not(layer1_outputs(4888)) or (layer1_outputs(495));
    layer2_outputs(2161) <= (layer1_outputs(671)) and (layer1_outputs(4460));
    layer2_outputs(2162) <= (layer1_outputs(1453)) and (layer1_outputs(2710));
    layer2_outputs(2163) <= not((layer1_outputs(3293)) and (layer1_outputs(749)));
    layer2_outputs(2164) <= (layer1_outputs(3971)) and not (layer1_outputs(4294));
    layer2_outputs(2165) <= layer1_outputs(94);
    layer2_outputs(2166) <= not((layer1_outputs(2051)) and (layer1_outputs(3073)));
    layer2_outputs(2167) <= not(layer1_outputs(3279));
    layer2_outputs(2168) <= not(layer1_outputs(1587));
    layer2_outputs(2169) <= not(layer1_outputs(944)) or (layer1_outputs(4166));
    layer2_outputs(2170) <= '0';
    layer2_outputs(2171) <= not(layer1_outputs(3780)) or (layer1_outputs(4666));
    layer2_outputs(2172) <= not(layer1_outputs(748));
    layer2_outputs(2173) <= layer1_outputs(4280);
    layer2_outputs(2174) <= not(layer1_outputs(2612)) or (layer1_outputs(2805));
    layer2_outputs(2175) <= (layer1_outputs(2569)) and (layer1_outputs(3262));
    layer2_outputs(2176) <= (layer1_outputs(3204)) or (layer1_outputs(4952));
    layer2_outputs(2177) <= layer1_outputs(2274);
    layer2_outputs(2178) <= (layer1_outputs(90)) or (layer1_outputs(2403));
    layer2_outputs(2179) <= layer1_outputs(3803);
    layer2_outputs(2180) <= not((layer1_outputs(4960)) xor (layer1_outputs(1427)));
    layer2_outputs(2181) <= '0';
    layer2_outputs(2182) <= '1';
    layer2_outputs(2183) <= '0';
    layer2_outputs(2184) <= not(layer1_outputs(4173));
    layer2_outputs(2185) <= '1';
    layer2_outputs(2186) <= not(layer1_outputs(3645));
    layer2_outputs(2187) <= (layer1_outputs(920)) and (layer1_outputs(3418));
    layer2_outputs(2188) <= (layer1_outputs(4494)) and not (layer1_outputs(4020));
    layer2_outputs(2189) <= (layer1_outputs(1282)) or (layer1_outputs(1403));
    layer2_outputs(2190) <= not(layer1_outputs(4809));
    layer2_outputs(2191) <= (layer1_outputs(2573)) and (layer1_outputs(180));
    layer2_outputs(2192) <= not((layer1_outputs(1558)) or (layer1_outputs(3082)));
    layer2_outputs(2193) <= layer1_outputs(3564);
    layer2_outputs(2194) <= not((layer1_outputs(4746)) and (layer1_outputs(1360)));
    layer2_outputs(2195) <= not((layer1_outputs(4335)) and (layer1_outputs(2155)));
    layer2_outputs(2196) <= not((layer1_outputs(406)) and (layer1_outputs(3409)));
    layer2_outputs(2197) <= (layer1_outputs(1794)) and not (layer1_outputs(360));
    layer2_outputs(2198) <= (layer1_outputs(2553)) or (layer1_outputs(188));
    layer2_outputs(2199) <= (layer1_outputs(2047)) xor (layer1_outputs(967));
    layer2_outputs(2200) <= '1';
    layer2_outputs(2201) <= layer1_outputs(4209);
    layer2_outputs(2202) <= not(layer1_outputs(4153));
    layer2_outputs(2203) <= layer1_outputs(875);
    layer2_outputs(2204) <= (layer1_outputs(4632)) and (layer1_outputs(2616));
    layer2_outputs(2205) <= not(layer1_outputs(4543));
    layer2_outputs(2206) <= not(layer1_outputs(1975));
    layer2_outputs(2207) <= (layer1_outputs(4819)) and (layer1_outputs(4509));
    layer2_outputs(2208) <= not(layer1_outputs(2878)) or (layer1_outputs(1721));
    layer2_outputs(2209) <= (layer1_outputs(2063)) xor (layer1_outputs(2836));
    layer2_outputs(2210) <= (layer1_outputs(3049)) or (layer1_outputs(4100));
    layer2_outputs(2211) <= not(layer1_outputs(2995));
    layer2_outputs(2212) <= not(layer1_outputs(1522)) or (layer1_outputs(2162));
    layer2_outputs(2213) <= not(layer1_outputs(5089));
    layer2_outputs(2214) <= (layer1_outputs(3296)) and not (layer1_outputs(4392));
    layer2_outputs(2215) <= (layer1_outputs(4604)) or (layer1_outputs(4470));
    layer2_outputs(2216) <= not(layer1_outputs(2851));
    layer2_outputs(2217) <= not(layer1_outputs(2606)) or (layer1_outputs(1144));
    layer2_outputs(2218) <= not(layer1_outputs(4001));
    layer2_outputs(2219) <= layer1_outputs(3565);
    layer2_outputs(2220) <= (layer1_outputs(2575)) or (layer1_outputs(4950));
    layer2_outputs(2221) <= '0';
    layer2_outputs(2222) <= '1';
    layer2_outputs(2223) <= not((layer1_outputs(310)) and (layer1_outputs(112)));
    layer2_outputs(2224) <= (layer1_outputs(833)) and not (layer1_outputs(4872));
    layer2_outputs(2225) <= not(layer1_outputs(4811));
    layer2_outputs(2226) <= '0';
    layer2_outputs(2227) <= not(layer1_outputs(4245));
    layer2_outputs(2228) <= (layer1_outputs(137)) or (layer1_outputs(3872));
    layer2_outputs(2229) <= (layer1_outputs(1653)) and not (layer1_outputs(856));
    layer2_outputs(2230) <= not((layer1_outputs(4494)) or (layer1_outputs(3371)));
    layer2_outputs(2231) <= (layer1_outputs(3000)) and not (layer1_outputs(4802));
    layer2_outputs(2232) <= (layer1_outputs(2204)) and not (layer1_outputs(804));
    layer2_outputs(2233) <= (layer1_outputs(3702)) or (layer1_outputs(719));
    layer2_outputs(2234) <= not(layer1_outputs(1053));
    layer2_outputs(2235) <= not(layer1_outputs(744));
    layer2_outputs(2236) <= not((layer1_outputs(993)) and (layer1_outputs(2419)));
    layer2_outputs(2237) <= not(layer1_outputs(650)) or (layer1_outputs(550));
    layer2_outputs(2238) <= layer1_outputs(4500);
    layer2_outputs(2239) <= (layer1_outputs(4340)) or (layer1_outputs(3398));
    layer2_outputs(2240) <= not((layer1_outputs(4754)) and (layer1_outputs(5041)));
    layer2_outputs(2241) <= layer1_outputs(58);
    layer2_outputs(2242) <= layer1_outputs(4868);
    layer2_outputs(2243) <= (layer1_outputs(1044)) and (layer1_outputs(4787));
    layer2_outputs(2244) <= not(layer1_outputs(3478)) or (layer1_outputs(2904));
    layer2_outputs(2245) <= (layer1_outputs(2888)) or (layer1_outputs(934));
    layer2_outputs(2246) <= not((layer1_outputs(5080)) or (layer1_outputs(3621)));
    layer2_outputs(2247) <= not(layer1_outputs(2869));
    layer2_outputs(2248) <= not(layer1_outputs(1882));
    layer2_outputs(2249) <= '0';
    layer2_outputs(2250) <= not(layer1_outputs(5001));
    layer2_outputs(2251) <= layer1_outputs(355);
    layer2_outputs(2252) <= '0';
    layer2_outputs(2253) <= '0';
    layer2_outputs(2254) <= (layer1_outputs(1555)) and not (layer1_outputs(4964));
    layer2_outputs(2255) <= not(layer1_outputs(4895));
    layer2_outputs(2256) <= (layer1_outputs(1493)) and not (layer1_outputs(2539));
    layer2_outputs(2257) <= layer1_outputs(4474);
    layer2_outputs(2258) <= not(layer1_outputs(3595));
    layer2_outputs(2259) <= not((layer1_outputs(1951)) or (layer1_outputs(1655)));
    layer2_outputs(2260) <= '0';
    layer2_outputs(2261) <= not(layer1_outputs(1149)) or (layer1_outputs(2072));
    layer2_outputs(2262) <= not(layer1_outputs(3084));
    layer2_outputs(2263) <= not(layer1_outputs(4708)) or (layer1_outputs(120));
    layer2_outputs(2264) <= layer1_outputs(2212);
    layer2_outputs(2265) <= not((layer1_outputs(898)) or (layer1_outputs(2191)));
    layer2_outputs(2266) <= not(layer1_outputs(4681));
    layer2_outputs(2267) <= layer1_outputs(3716);
    layer2_outputs(2268) <= layer1_outputs(395);
    layer2_outputs(2269) <= (layer1_outputs(425)) and not (layer1_outputs(4415));
    layer2_outputs(2270) <= not(layer1_outputs(1984));
    layer2_outputs(2271) <= (layer1_outputs(2594)) and not (layer1_outputs(589));
    layer2_outputs(2272) <= layer1_outputs(2137);
    layer2_outputs(2273) <= layer1_outputs(3712);
    layer2_outputs(2274) <= layer1_outputs(3036);
    layer2_outputs(2275) <= (layer1_outputs(3962)) or (layer1_outputs(3920));
    layer2_outputs(2276) <= layer1_outputs(1680);
    layer2_outputs(2277) <= (layer1_outputs(2785)) and not (layer1_outputs(1028));
    layer2_outputs(2278) <= not(layer1_outputs(1776));
    layer2_outputs(2279) <= not((layer1_outputs(3686)) and (layer1_outputs(1770)));
    layer2_outputs(2280) <= (layer1_outputs(816)) or (layer1_outputs(2609));
    layer2_outputs(2281) <= layer1_outputs(2576);
    layer2_outputs(2282) <= not((layer1_outputs(356)) or (layer1_outputs(4970)));
    layer2_outputs(2283) <= layer1_outputs(1304);
    layer2_outputs(2284) <= not(layer1_outputs(2057));
    layer2_outputs(2285) <= (layer1_outputs(4117)) and not (layer1_outputs(4261));
    layer2_outputs(2286) <= not(layer1_outputs(3230));
    layer2_outputs(2287) <= not((layer1_outputs(1045)) and (layer1_outputs(3016)));
    layer2_outputs(2288) <= (layer1_outputs(5112)) and not (layer1_outputs(1545));
    layer2_outputs(2289) <= '1';
    layer2_outputs(2290) <= layer1_outputs(1986);
    layer2_outputs(2291) <= (layer1_outputs(4978)) and (layer1_outputs(281));
    layer2_outputs(2292) <= not((layer1_outputs(2349)) and (layer1_outputs(3492)));
    layer2_outputs(2293) <= (layer1_outputs(1683)) and not (layer1_outputs(4182));
    layer2_outputs(2294) <= (layer1_outputs(975)) and not (layer1_outputs(2800));
    layer2_outputs(2295) <= not(layer1_outputs(3932)) or (layer1_outputs(160));
    layer2_outputs(2296) <= not(layer1_outputs(1218)) or (layer1_outputs(1813));
    layer2_outputs(2297) <= (layer1_outputs(2979)) and not (layer1_outputs(1553));
    layer2_outputs(2298) <= (layer1_outputs(3414)) and not (layer1_outputs(1839));
    layer2_outputs(2299) <= layer1_outputs(2501);
    layer2_outputs(2300) <= not((layer1_outputs(4164)) and (layer1_outputs(4692)));
    layer2_outputs(2301) <= not((layer1_outputs(2835)) or (layer1_outputs(3355)));
    layer2_outputs(2302) <= (layer1_outputs(2091)) and not (layer1_outputs(4694));
    layer2_outputs(2303) <= (layer1_outputs(2910)) and not (layer1_outputs(1586));
    layer2_outputs(2304) <= not(layer1_outputs(2659));
    layer2_outputs(2305) <= layer1_outputs(1878);
    layer2_outputs(2306) <= not(layer1_outputs(848));
    layer2_outputs(2307) <= not(layer1_outputs(2074));
    layer2_outputs(2308) <= '0';
    layer2_outputs(2309) <= '1';
    layer2_outputs(2310) <= not((layer1_outputs(231)) or (layer1_outputs(416)));
    layer2_outputs(2311) <= '1';
    layer2_outputs(2312) <= layer1_outputs(4752);
    layer2_outputs(2313) <= not(layer1_outputs(1228));
    layer2_outputs(2314) <= not((layer1_outputs(969)) and (layer1_outputs(1510)));
    layer2_outputs(2315) <= layer1_outputs(869);
    layer2_outputs(2316) <= not((layer1_outputs(883)) or (layer1_outputs(2508)));
    layer2_outputs(2317) <= not(layer1_outputs(513)) or (layer1_outputs(3207));
    layer2_outputs(2318) <= (layer1_outputs(3504)) and not (layer1_outputs(4787));
    layer2_outputs(2319) <= '0';
    layer2_outputs(2320) <= (layer1_outputs(3210)) and not (layer1_outputs(1397));
    layer2_outputs(2321) <= layer1_outputs(1229);
    layer2_outputs(2322) <= '1';
    layer2_outputs(2323) <= (layer1_outputs(4373)) or (layer1_outputs(981));
    layer2_outputs(2324) <= not(layer1_outputs(699)) or (layer1_outputs(4999));
    layer2_outputs(2325) <= (layer1_outputs(2960)) and not (layer1_outputs(2271));
    layer2_outputs(2326) <= layer1_outputs(1634);
    layer2_outputs(2327) <= not(layer1_outputs(4588));
    layer2_outputs(2328) <= '1';
    layer2_outputs(2329) <= (layer1_outputs(2209)) and not (layer1_outputs(4596));
    layer2_outputs(2330) <= (layer1_outputs(363)) and not (layer1_outputs(997));
    layer2_outputs(2331) <= not((layer1_outputs(2965)) and (layer1_outputs(2331)));
    layer2_outputs(2332) <= not(layer1_outputs(1612));
    layer2_outputs(2333) <= (layer1_outputs(377)) and not (layer1_outputs(2334));
    layer2_outputs(2334) <= not(layer1_outputs(2725));
    layer2_outputs(2335) <= not(layer1_outputs(4145));
    layer2_outputs(2336) <= not(layer1_outputs(3285));
    layer2_outputs(2337) <= layer1_outputs(4646);
    layer2_outputs(2338) <= not(layer1_outputs(606));
    layer2_outputs(2339) <= (layer1_outputs(1882)) or (layer1_outputs(4853));
    layer2_outputs(2340) <= (layer1_outputs(2695)) and not (layer1_outputs(2503));
    layer2_outputs(2341) <= not(layer1_outputs(1931));
    layer2_outputs(2342) <= not(layer1_outputs(2730));
    layer2_outputs(2343) <= not((layer1_outputs(4328)) and (layer1_outputs(34)));
    layer2_outputs(2344) <= not(layer1_outputs(4138)) or (layer1_outputs(871));
    layer2_outputs(2345) <= layer1_outputs(4727);
    layer2_outputs(2346) <= '0';
    layer2_outputs(2347) <= '1';
    layer2_outputs(2348) <= not(layer1_outputs(1299));
    layer2_outputs(2349) <= not(layer1_outputs(796));
    layer2_outputs(2350) <= not(layer1_outputs(3937));
    layer2_outputs(2351) <= not(layer1_outputs(2774)) or (layer1_outputs(1912));
    layer2_outputs(2352) <= not((layer1_outputs(4885)) and (layer1_outputs(2289)));
    layer2_outputs(2353) <= layer1_outputs(3893);
    layer2_outputs(2354) <= not(layer1_outputs(2334)) or (layer1_outputs(4080));
    layer2_outputs(2355) <= not(layer1_outputs(2577));
    layer2_outputs(2356) <= (layer1_outputs(4855)) and not (layer1_outputs(244));
    layer2_outputs(2357) <= (layer1_outputs(4791)) and (layer1_outputs(3734));
    layer2_outputs(2358) <= layer1_outputs(1752);
    layer2_outputs(2359) <= (layer1_outputs(70)) and not (layer1_outputs(2584));
    layer2_outputs(2360) <= '1';
    layer2_outputs(2361) <= not(layer1_outputs(968));
    layer2_outputs(2362) <= layer1_outputs(2026);
    layer2_outputs(2363) <= layer1_outputs(2881);
    layer2_outputs(2364) <= (layer1_outputs(440)) and not (layer1_outputs(2640));
    layer2_outputs(2365) <= not(layer1_outputs(2915));
    layer2_outputs(2366) <= '0';
    layer2_outputs(2367) <= not(layer1_outputs(3559));
    layer2_outputs(2368) <= '1';
    layer2_outputs(2369) <= not((layer1_outputs(3513)) or (layer1_outputs(4556)));
    layer2_outputs(2370) <= layer1_outputs(2181);
    layer2_outputs(2371) <= '1';
    layer2_outputs(2372) <= layer1_outputs(4942);
    layer2_outputs(2373) <= '1';
    layer2_outputs(2374) <= (layer1_outputs(3336)) and (layer1_outputs(4904));
    layer2_outputs(2375) <= not((layer1_outputs(2023)) or (layer1_outputs(1536)));
    layer2_outputs(2376) <= not(layer1_outputs(3201)) or (layer1_outputs(3937));
    layer2_outputs(2377) <= layer1_outputs(2594);
    layer2_outputs(2378) <= '0';
    layer2_outputs(2379) <= (layer1_outputs(1520)) and not (layer1_outputs(3480));
    layer2_outputs(2380) <= '1';
    layer2_outputs(2381) <= (layer1_outputs(4561)) and (layer1_outputs(1315));
    layer2_outputs(2382) <= not((layer1_outputs(1245)) and (layer1_outputs(2249)));
    layer2_outputs(2383) <= not(layer1_outputs(1390)) or (layer1_outputs(3037));
    layer2_outputs(2384) <= not((layer1_outputs(4066)) and (layer1_outputs(3110)));
    layer2_outputs(2385) <= (layer1_outputs(2612)) and not (layer1_outputs(940));
    layer2_outputs(2386) <= not(layer1_outputs(2928)) or (layer1_outputs(2269));
    layer2_outputs(2387) <= not(layer1_outputs(4605));
    layer2_outputs(2388) <= (layer1_outputs(3127)) or (layer1_outputs(2439));
    layer2_outputs(2389) <= not(layer1_outputs(267));
    layer2_outputs(2390) <= (layer1_outputs(4700)) or (layer1_outputs(2473));
    layer2_outputs(2391) <= not(layer1_outputs(2836));
    layer2_outputs(2392) <= not(layer1_outputs(2556));
    layer2_outputs(2393) <= not(layer1_outputs(4002));
    layer2_outputs(2394) <= (layer1_outputs(3095)) or (layer1_outputs(1898));
    layer2_outputs(2395) <= layer1_outputs(1393);
    layer2_outputs(2396) <= not(layer1_outputs(3083));
    layer2_outputs(2397) <= not((layer1_outputs(1710)) or (layer1_outputs(3214)));
    layer2_outputs(2398) <= layer1_outputs(1907);
    layer2_outputs(2399) <= (layer1_outputs(1467)) and not (layer1_outputs(57));
    layer2_outputs(2400) <= not(layer1_outputs(4726)) or (layer1_outputs(4583));
    layer2_outputs(2401) <= not((layer1_outputs(1328)) and (layer1_outputs(3061)));
    layer2_outputs(2402) <= not(layer1_outputs(3341));
    layer2_outputs(2403) <= not(layer1_outputs(1287)) or (layer1_outputs(2446));
    layer2_outputs(2404) <= layer1_outputs(1409);
    layer2_outputs(2405) <= not(layer1_outputs(20));
    layer2_outputs(2406) <= layer1_outputs(3647);
    layer2_outputs(2407) <= (layer1_outputs(2073)) and not (layer1_outputs(4902));
    layer2_outputs(2408) <= not(layer1_outputs(1967));
    layer2_outputs(2409) <= not(layer1_outputs(4118)) or (layer1_outputs(1338));
    layer2_outputs(2410) <= (layer1_outputs(3618)) and not (layer1_outputs(3441));
    layer2_outputs(2411) <= '1';
    layer2_outputs(2412) <= not(layer1_outputs(4451));
    layer2_outputs(2413) <= (layer1_outputs(5073)) and not (layer1_outputs(3976));
    layer2_outputs(2414) <= '0';
    layer2_outputs(2415) <= '1';
    layer2_outputs(2416) <= layer1_outputs(3115);
    layer2_outputs(2417) <= layer1_outputs(3395);
    layer2_outputs(2418) <= layer1_outputs(2895);
    layer2_outputs(2419) <= (layer1_outputs(3967)) and not (layer1_outputs(4718));
    layer2_outputs(2420) <= '1';
    layer2_outputs(2421) <= not(layer1_outputs(4524));
    layer2_outputs(2422) <= not(layer1_outputs(3949)) or (layer1_outputs(2669));
    layer2_outputs(2423) <= (layer1_outputs(524)) or (layer1_outputs(2828));
    layer2_outputs(2424) <= '1';
    layer2_outputs(2425) <= not(layer1_outputs(4819)) or (layer1_outputs(5084));
    layer2_outputs(2426) <= '0';
    layer2_outputs(2427) <= not(layer1_outputs(3710));
    layer2_outputs(2428) <= not(layer1_outputs(1530)) or (layer1_outputs(3124));
    layer2_outputs(2429) <= not(layer1_outputs(1787));
    layer2_outputs(2430) <= layer1_outputs(1963);
    layer2_outputs(2431) <= (layer1_outputs(3753)) xor (layer1_outputs(2660));
    layer2_outputs(2432) <= not(layer1_outputs(3935));
    layer2_outputs(2433) <= '0';
    layer2_outputs(2434) <= layer1_outputs(4948);
    layer2_outputs(2435) <= not((layer1_outputs(783)) or (layer1_outputs(3771)));
    layer2_outputs(2436) <= layer1_outputs(2792);
    layer2_outputs(2437) <= (layer1_outputs(3781)) or (layer1_outputs(2023));
    layer2_outputs(2438) <= not(layer1_outputs(4415)) or (layer1_outputs(2206));
    layer2_outputs(2439) <= (layer1_outputs(1401)) and not (layer1_outputs(998));
    layer2_outputs(2440) <= layer1_outputs(2896);
    layer2_outputs(2441) <= not((layer1_outputs(238)) and (layer1_outputs(85)));
    layer2_outputs(2442) <= '1';
    layer2_outputs(2443) <= layer1_outputs(3543);
    layer2_outputs(2444) <= '0';
    layer2_outputs(2445) <= not(layer1_outputs(490));
    layer2_outputs(2446) <= not((layer1_outputs(3163)) or (layer1_outputs(1483)));
    layer2_outputs(2447) <= not((layer1_outputs(3447)) or (layer1_outputs(4955)));
    layer2_outputs(2448) <= '1';
    layer2_outputs(2449) <= (layer1_outputs(5074)) or (layer1_outputs(2044));
    layer2_outputs(2450) <= not(layer1_outputs(4976)) or (layer1_outputs(3944));
    layer2_outputs(2451) <= not((layer1_outputs(1503)) or (layer1_outputs(4571)));
    layer2_outputs(2452) <= (layer1_outputs(2749)) and (layer1_outputs(1476));
    layer2_outputs(2453) <= not(layer1_outputs(2932));
    layer2_outputs(2454) <= not(layer1_outputs(4032));
    layer2_outputs(2455) <= layer1_outputs(2627);
    layer2_outputs(2456) <= (layer1_outputs(3198)) and not (layer1_outputs(1147));
    layer2_outputs(2457) <= not(layer1_outputs(4091));
    layer2_outputs(2458) <= layer1_outputs(4573);
    layer2_outputs(2459) <= (layer1_outputs(4959)) or (layer1_outputs(1046));
    layer2_outputs(2460) <= (layer1_outputs(218)) and (layer1_outputs(4578));
    layer2_outputs(2461) <= layer1_outputs(1218);
    layer2_outputs(2462) <= (layer1_outputs(487)) and (layer1_outputs(762));
    layer2_outputs(2463) <= not(layer1_outputs(3411)) or (layer1_outputs(4349));
    layer2_outputs(2464) <= not(layer1_outputs(493));
    layer2_outputs(2465) <= (layer1_outputs(1048)) and not (layer1_outputs(392));
    layer2_outputs(2466) <= (layer1_outputs(4595)) and not (layer1_outputs(197));
    layer2_outputs(2467) <= not((layer1_outputs(2927)) or (layer1_outputs(4137)));
    layer2_outputs(2468) <= not(layer1_outputs(4716));
    layer2_outputs(2469) <= layer1_outputs(5115);
    layer2_outputs(2470) <= not(layer1_outputs(1635));
    layer2_outputs(2471) <= not(layer1_outputs(2815)) or (layer1_outputs(1883));
    layer2_outputs(2472) <= not(layer1_outputs(1618)) or (layer1_outputs(1672));
    layer2_outputs(2473) <= not(layer1_outputs(723)) or (layer1_outputs(2022));
    layer2_outputs(2474) <= not((layer1_outputs(2704)) and (layer1_outputs(5008)));
    layer2_outputs(2475) <= not((layer1_outputs(2247)) or (layer1_outputs(1464)));
    layer2_outputs(2476) <= layer1_outputs(3977);
    layer2_outputs(2477) <= '0';
    layer2_outputs(2478) <= '0';
    layer2_outputs(2479) <= '0';
    layer2_outputs(2480) <= not((layer1_outputs(2413)) or (layer1_outputs(886)));
    layer2_outputs(2481) <= not((layer1_outputs(4651)) or (layer1_outputs(2632)));
    layer2_outputs(2482) <= not(layer1_outputs(3133));
    layer2_outputs(2483) <= layer1_outputs(2352);
    layer2_outputs(2484) <= '0';
    layer2_outputs(2485) <= not((layer1_outputs(4082)) and (layer1_outputs(3092)));
    layer2_outputs(2486) <= (layer1_outputs(3887)) and (layer1_outputs(4938));
    layer2_outputs(2487) <= not(layer1_outputs(4310));
    layer2_outputs(2488) <= not(layer1_outputs(2890));
    layer2_outputs(2489) <= (layer1_outputs(4363)) and (layer1_outputs(3776));
    layer2_outputs(2490) <= not(layer1_outputs(3515));
    layer2_outputs(2491) <= not(layer1_outputs(4591));
    layer2_outputs(2492) <= (layer1_outputs(1398)) and not (layer1_outputs(3704));
    layer2_outputs(2493) <= (layer1_outputs(1951)) and not (layer1_outputs(3756));
    layer2_outputs(2494) <= '0';
    layer2_outputs(2495) <= '1';
    layer2_outputs(2496) <= (layer1_outputs(770)) and not (layer1_outputs(3573));
    layer2_outputs(2497) <= not(layer1_outputs(4132));
    layer2_outputs(2498) <= not((layer1_outputs(2879)) or (layer1_outputs(2515)));
    layer2_outputs(2499) <= '0';
    layer2_outputs(2500) <= not(layer1_outputs(982));
    layer2_outputs(2501) <= '0';
    layer2_outputs(2502) <= not(layer1_outputs(962)) or (layer1_outputs(169));
    layer2_outputs(2503) <= layer1_outputs(3869);
    layer2_outputs(2504) <= (layer1_outputs(3874)) or (layer1_outputs(494));
    layer2_outputs(2505) <= (layer1_outputs(4104)) and not (layer1_outputs(4485));
    layer2_outputs(2506) <= layer1_outputs(1836);
    layer2_outputs(2507) <= layer1_outputs(549);
    layer2_outputs(2508) <= layer1_outputs(798);
    layer2_outputs(2509) <= not(layer1_outputs(4936)) or (layer1_outputs(3420));
    layer2_outputs(2510) <= not((layer1_outputs(2552)) or (layer1_outputs(3265)));
    layer2_outputs(2511) <= layer1_outputs(4187);
    layer2_outputs(2512) <= (layer1_outputs(597)) and not (layer1_outputs(528));
    layer2_outputs(2513) <= layer1_outputs(689);
    layer2_outputs(2514) <= '0';
    layer2_outputs(2515) <= not(layer1_outputs(4748));
    layer2_outputs(2516) <= '0';
    layer2_outputs(2517) <= not(layer1_outputs(3451)) or (layer1_outputs(519));
    layer2_outputs(2518) <= (layer1_outputs(683)) or (layer1_outputs(262));
    layer2_outputs(2519) <= not((layer1_outputs(240)) or (layer1_outputs(4084)));
    layer2_outputs(2520) <= not((layer1_outputs(2024)) and (layer1_outputs(1981)));
    layer2_outputs(2521) <= not(layer1_outputs(4528)) or (layer1_outputs(3131));
    layer2_outputs(2522) <= not(layer1_outputs(1480));
    layer2_outputs(2523) <= layer1_outputs(645);
    layer2_outputs(2524) <= '0';
    layer2_outputs(2525) <= not((layer1_outputs(948)) xor (layer1_outputs(1758)));
    layer2_outputs(2526) <= '0';
    layer2_outputs(2527) <= not(layer1_outputs(2210));
    layer2_outputs(2528) <= not(layer1_outputs(1289));
    layer2_outputs(2529) <= not(layer1_outputs(4580));
    layer2_outputs(2530) <= (layer1_outputs(2000)) and not (layer1_outputs(5015));
    layer2_outputs(2531) <= not(layer1_outputs(4281));
    layer2_outputs(2532) <= layer1_outputs(1496);
    layer2_outputs(2533) <= not((layer1_outputs(2556)) or (layer1_outputs(1075)));
    layer2_outputs(2534) <= layer1_outputs(61);
    layer2_outputs(2535) <= not(layer1_outputs(3358));
    layer2_outputs(2536) <= layer1_outputs(1052);
    layer2_outputs(2537) <= (layer1_outputs(1621)) or (layer1_outputs(4806));
    layer2_outputs(2538) <= layer1_outputs(2457);
    layer2_outputs(2539) <= layer1_outputs(2361);
    layer2_outputs(2540) <= (layer1_outputs(4893)) and not (layer1_outputs(1599));
    layer2_outputs(2541) <= '1';
    layer2_outputs(2542) <= (layer1_outputs(3741)) and not (layer1_outputs(2849));
    layer2_outputs(2543) <= '0';
    layer2_outputs(2544) <= (layer1_outputs(2775)) and not (layer1_outputs(4424));
    layer2_outputs(2545) <= '0';
    layer2_outputs(2546) <= '0';
    layer2_outputs(2547) <= (layer1_outputs(2435)) and not (layer1_outputs(3973));
    layer2_outputs(2548) <= '0';
    layer2_outputs(2549) <= not(layer1_outputs(2297)) or (layer1_outputs(2322));
    layer2_outputs(2550) <= (layer1_outputs(855)) xor (layer1_outputs(1577));
    layer2_outputs(2551) <= not((layer1_outputs(4176)) and (layer1_outputs(2706)));
    layer2_outputs(2552) <= '0';
    layer2_outputs(2553) <= not((layer1_outputs(4885)) and (layer1_outputs(3113)));
    layer2_outputs(2554) <= '1';
    layer2_outputs(2555) <= '0';
    layer2_outputs(2556) <= '0';
    layer2_outputs(2557) <= '1';
    layer2_outputs(2558) <= (layer1_outputs(3526)) and (layer1_outputs(263));
    layer2_outputs(2559) <= not(layer1_outputs(2994)) or (layer1_outputs(2489));
    layer2_outputs(2560) <= not(layer1_outputs(1527)) or (layer1_outputs(2709));
    layer2_outputs(2561) <= layer1_outputs(2336);
    layer2_outputs(2562) <= (layer1_outputs(2512)) and not (layer1_outputs(4612));
    layer2_outputs(2563) <= not((layer1_outputs(2002)) and (layer1_outputs(1809)));
    layer2_outputs(2564) <= '1';
    layer2_outputs(2565) <= (layer1_outputs(3245)) and (layer1_outputs(3530));
    layer2_outputs(2566) <= '0';
    layer2_outputs(2567) <= layer1_outputs(2622);
    layer2_outputs(2568) <= '1';
    layer2_outputs(2569) <= not((layer1_outputs(1362)) and (layer1_outputs(1628)));
    layer2_outputs(2570) <= (layer1_outputs(1980)) and (layer1_outputs(3990));
    layer2_outputs(2571) <= not((layer1_outputs(3467)) and (layer1_outputs(28)));
    layer2_outputs(2572) <= (layer1_outputs(4663)) and not (layer1_outputs(3635));
    layer2_outputs(2573) <= '0';
    layer2_outputs(2574) <= (layer1_outputs(301)) and not (layer1_outputs(1573));
    layer2_outputs(2575) <= not(layer1_outputs(1128));
    layer2_outputs(2576) <= layer1_outputs(4474);
    layer2_outputs(2577) <= layer1_outputs(3389);
    layer2_outputs(2578) <= (layer1_outputs(1271)) and not (layer1_outputs(2250));
    layer2_outputs(2579) <= not(layer1_outputs(4701)) or (layer1_outputs(4455));
    layer2_outputs(2580) <= (layer1_outputs(5108)) or (layer1_outputs(3714));
    layer2_outputs(2581) <= '1';
    layer2_outputs(2582) <= not(layer1_outputs(1820)) or (layer1_outputs(1011));
    layer2_outputs(2583) <= not((layer1_outputs(800)) and (layer1_outputs(614)));
    layer2_outputs(2584) <= (layer1_outputs(1069)) and not (layer1_outputs(321));
    layer2_outputs(2585) <= not(layer1_outputs(4365));
    layer2_outputs(2586) <= not(layer1_outputs(4072)) or (layer1_outputs(3125));
    layer2_outputs(2587) <= '0';
    layer2_outputs(2588) <= not(layer1_outputs(826));
    layer2_outputs(2589) <= '0';
    layer2_outputs(2590) <= layer1_outputs(1404);
    layer2_outputs(2591) <= not((layer1_outputs(752)) or (layer1_outputs(3224)));
    layer2_outputs(2592) <= (layer1_outputs(4339)) and (layer1_outputs(4990));
    layer2_outputs(2593) <= not((layer1_outputs(3255)) or (layer1_outputs(573)));
    layer2_outputs(2594) <= (layer1_outputs(2391)) and not (layer1_outputs(4662));
    layer2_outputs(2595) <= not((layer1_outputs(2185)) or (layer1_outputs(2766)));
    layer2_outputs(2596) <= not(layer1_outputs(2507)) or (layer1_outputs(2959));
    layer2_outputs(2597) <= layer1_outputs(3285);
    layer2_outputs(2598) <= not((layer1_outputs(3446)) and (layer1_outputs(2593)));
    layer2_outputs(2599) <= not((layer1_outputs(4781)) and (layer1_outputs(4583)));
    layer2_outputs(2600) <= not(layer1_outputs(2232)) or (layer1_outputs(575));
    layer2_outputs(2601) <= not(layer1_outputs(1323));
    layer2_outputs(2602) <= '0';
    layer2_outputs(2603) <= layer1_outputs(3959);
    layer2_outputs(2604) <= (layer1_outputs(4435)) and not (layer1_outputs(2101));
    layer2_outputs(2605) <= (layer1_outputs(763)) or (layer1_outputs(4274));
    layer2_outputs(2606) <= layer1_outputs(3763);
    layer2_outputs(2607) <= not(layer1_outputs(613)) or (layer1_outputs(3701));
    layer2_outputs(2608) <= not(layer1_outputs(110));
    layer2_outputs(2609) <= '1';
    layer2_outputs(2610) <= layer1_outputs(3151);
    layer2_outputs(2611) <= not((layer1_outputs(5007)) xor (layer1_outputs(64)));
    layer2_outputs(2612) <= not((layer1_outputs(4926)) or (layer1_outputs(4572)));
    layer2_outputs(2613) <= not((layer1_outputs(2739)) and (layer1_outputs(2019)));
    layer2_outputs(2614) <= not((layer1_outputs(3517)) and (layer1_outputs(2369)));
    layer2_outputs(2615) <= (layer1_outputs(1054)) or (layer1_outputs(3877));
    layer2_outputs(2616) <= not(layer1_outputs(710)) or (layer1_outputs(1991));
    layer2_outputs(2617) <= not(layer1_outputs(835));
    layer2_outputs(2618) <= not((layer1_outputs(1678)) or (layer1_outputs(4986)));
    layer2_outputs(2619) <= (layer1_outputs(2866)) xor (layer1_outputs(5024));
    layer2_outputs(2620) <= layer1_outputs(703);
    layer2_outputs(2621) <= not(layer1_outputs(1040)) or (layer1_outputs(3743));
    layer2_outputs(2622) <= layer1_outputs(788);
    layer2_outputs(2623) <= '1';
    layer2_outputs(2624) <= not((layer1_outputs(2951)) and (layer1_outputs(2681)));
    layer2_outputs(2625) <= '0';
    layer2_outputs(2626) <= layer1_outputs(732);
    layer2_outputs(2627) <= not(layer1_outputs(2670)) or (layer1_outputs(2536));
    layer2_outputs(2628) <= (layer1_outputs(127)) and not (layer1_outputs(2185));
    layer2_outputs(2629) <= layer1_outputs(539);
    layer2_outputs(2630) <= not((layer1_outputs(4476)) and (layer1_outputs(5093)));
    layer2_outputs(2631) <= (layer1_outputs(1212)) and (layer1_outputs(4267));
    layer2_outputs(2632) <= not(layer1_outputs(2220)) or (layer1_outputs(1737));
    layer2_outputs(2633) <= (layer1_outputs(1171)) and not (layer1_outputs(1426));
    layer2_outputs(2634) <= not(layer1_outputs(1072));
    layer2_outputs(2635) <= not(layer1_outputs(3436)) or (layer1_outputs(2338));
    layer2_outputs(2636) <= not(layer1_outputs(1955));
    layer2_outputs(2637) <= layer1_outputs(4126);
    layer2_outputs(2638) <= layer1_outputs(4144);
    layer2_outputs(2639) <= (layer1_outputs(4615)) and not (layer1_outputs(4671));
    layer2_outputs(2640) <= (layer1_outputs(662)) and not (layer1_outputs(2920));
    layer2_outputs(2641) <= '0';
    layer2_outputs(2642) <= '0';
    layer2_outputs(2643) <= (layer1_outputs(681)) or (layer1_outputs(3135));
    layer2_outputs(2644) <= '0';
    layer2_outputs(2645) <= not(layer1_outputs(2419)) or (layer1_outputs(1273));
    layer2_outputs(2646) <= not(layer1_outputs(3504)) or (layer1_outputs(2471));
    layer2_outputs(2647) <= layer1_outputs(105);
    layer2_outputs(2648) <= (layer1_outputs(577)) and (layer1_outputs(2293));
    layer2_outputs(2649) <= not(layer1_outputs(3072));
    layer2_outputs(2650) <= layer1_outputs(404);
    layer2_outputs(2651) <= (layer1_outputs(1357)) or (layer1_outputs(1785));
    layer2_outputs(2652) <= layer1_outputs(3652);
    layer2_outputs(2653) <= layer1_outputs(1004);
    layer2_outputs(2654) <= '1';
    layer2_outputs(2655) <= layer1_outputs(3439);
    layer2_outputs(2656) <= not(layer1_outputs(4894)) or (layer1_outputs(3847));
    layer2_outputs(2657) <= (layer1_outputs(2028)) and (layer1_outputs(2006));
    layer2_outputs(2658) <= not(layer1_outputs(819));
    layer2_outputs(2659) <= layer1_outputs(4313);
    layer2_outputs(2660) <= (layer1_outputs(2828)) and not (layer1_outputs(410));
    layer2_outputs(2661) <= '0';
    layer2_outputs(2662) <= '1';
    layer2_outputs(2663) <= (layer1_outputs(1465)) or (layer1_outputs(3647));
    layer2_outputs(2664) <= layer1_outputs(588);
    layer2_outputs(2665) <= not(layer1_outputs(4458));
    layer2_outputs(2666) <= not((layer1_outputs(5004)) xor (layer1_outputs(4738)));
    layer2_outputs(2667) <= (layer1_outputs(3431)) and (layer1_outputs(3176));
    layer2_outputs(2668) <= not((layer1_outputs(4076)) or (layer1_outputs(3883)));
    layer2_outputs(2669) <= (layer1_outputs(4199)) or (layer1_outputs(2103));
    layer2_outputs(2670) <= not(layer1_outputs(1833));
    layer2_outputs(2671) <= '1';
    layer2_outputs(2672) <= not((layer1_outputs(1045)) and (layer1_outputs(2451)));
    layer2_outputs(2673) <= (layer1_outputs(235)) and not (layer1_outputs(4552));
    layer2_outputs(2674) <= layer1_outputs(1895);
    layer2_outputs(2675) <= not(layer1_outputs(429)) or (layer1_outputs(465));
    layer2_outputs(2676) <= (layer1_outputs(4780)) and not (layer1_outputs(268));
    layer2_outputs(2677) <= layer1_outputs(1213);
    layer2_outputs(2678) <= '1';
    layer2_outputs(2679) <= not(layer1_outputs(868));
    layer2_outputs(2680) <= not(layer1_outputs(293));
    layer2_outputs(2681) <= not((layer1_outputs(3941)) or (layer1_outputs(2189)));
    layer2_outputs(2682) <= layer1_outputs(4876);
    layer2_outputs(2683) <= '1';
    layer2_outputs(2684) <= layer1_outputs(2790);
    layer2_outputs(2685) <= not(layer1_outputs(4060));
    layer2_outputs(2686) <= not((layer1_outputs(2916)) and (layer1_outputs(5004)));
    layer2_outputs(2687) <= '1';
    layer2_outputs(2688) <= not((layer1_outputs(1751)) xor (layer1_outputs(4369)));
    layer2_outputs(2689) <= not(layer1_outputs(2420));
    layer2_outputs(2690) <= not((layer1_outputs(1816)) or (layer1_outputs(814)));
    layer2_outputs(2691) <= not(layer1_outputs(4920));
    layer2_outputs(2692) <= (layer1_outputs(540)) xor (layer1_outputs(3152));
    layer2_outputs(2693) <= layer1_outputs(1748);
    layer2_outputs(2694) <= '0';
    layer2_outputs(2695) <= '1';
    layer2_outputs(2696) <= not((layer1_outputs(3651)) or (layer1_outputs(3638)));
    layer2_outputs(2697) <= (layer1_outputs(2926)) and not (layer1_outputs(4557));
    layer2_outputs(2698) <= not((layer1_outputs(2742)) or (layer1_outputs(5018)));
    layer2_outputs(2699) <= '1';
    layer2_outputs(2700) <= '1';
    layer2_outputs(2701) <= (layer1_outputs(4661)) and (layer1_outputs(4851));
    layer2_outputs(2702) <= (layer1_outputs(0)) and not (layer1_outputs(455));
    layer2_outputs(2703) <= not(layer1_outputs(4388));
    layer2_outputs(2704) <= '0';
    layer2_outputs(2705) <= (layer1_outputs(3819)) and (layer1_outputs(1210));
    layer2_outputs(2706) <= not(layer1_outputs(3669)) or (layer1_outputs(1110));
    layer2_outputs(2707) <= not(layer1_outputs(3725));
    layer2_outputs(2708) <= (layer1_outputs(2425)) and (layer1_outputs(1825));
    layer2_outputs(2709) <= '0';
    layer2_outputs(2710) <= (layer1_outputs(2639)) and not (layer1_outputs(3417));
    layer2_outputs(2711) <= layer1_outputs(1289);
    layer2_outputs(2712) <= not(layer1_outputs(1433)) or (layer1_outputs(4090));
    layer2_outputs(2713) <= not(layer1_outputs(4061));
    layer2_outputs(2714) <= (layer1_outputs(821)) and not (layer1_outputs(3684));
    layer2_outputs(2715) <= '1';
    layer2_outputs(2716) <= (layer1_outputs(2527)) and not (layer1_outputs(1335));
    layer2_outputs(2717) <= not((layer1_outputs(579)) or (layer1_outputs(1922)));
    layer2_outputs(2718) <= not(layer1_outputs(1669));
    layer2_outputs(2719) <= '1';
    layer2_outputs(2720) <= (layer1_outputs(4034)) and (layer1_outputs(3940));
    layer2_outputs(2721) <= (layer1_outputs(2978)) and (layer1_outputs(2952));
    layer2_outputs(2722) <= not(layer1_outputs(619));
    layer2_outputs(2723) <= '0';
    layer2_outputs(2724) <= layer1_outputs(329);
    layer2_outputs(2725) <= (layer1_outputs(4251)) and (layer1_outputs(2053));
    layer2_outputs(2726) <= not((layer1_outputs(4)) or (layer1_outputs(4484)));
    layer2_outputs(2727) <= layer1_outputs(3308);
    layer2_outputs(2728) <= '0';
    layer2_outputs(2729) <= not(layer1_outputs(1657)) or (layer1_outputs(3111));
    layer2_outputs(2730) <= (layer1_outputs(1166)) and not (layer1_outputs(812));
    layer2_outputs(2731) <= not((layer1_outputs(2)) and (layer1_outputs(3485)));
    layer2_outputs(2732) <= not(layer1_outputs(2208));
    layer2_outputs(2733) <= (layer1_outputs(378)) and not (layer1_outputs(4536));
    layer2_outputs(2734) <= (layer1_outputs(1163)) and not (layer1_outputs(1848));
    layer2_outputs(2735) <= (layer1_outputs(1308)) xor (layer1_outputs(424));
    layer2_outputs(2736) <= not(layer1_outputs(241));
    layer2_outputs(2737) <= not(layer1_outputs(2973));
    layer2_outputs(2738) <= '1';
    layer2_outputs(2739) <= not(layer1_outputs(4399));
    layer2_outputs(2740) <= not(layer1_outputs(2455)) or (layer1_outputs(4178));
    layer2_outputs(2741) <= not(layer1_outputs(234));
    layer2_outputs(2742) <= not(layer1_outputs(3648));
    layer2_outputs(2743) <= not(layer1_outputs(864)) or (layer1_outputs(4177));
    layer2_outputs(2744) <= not((layer1_outputs(66)) and (layer1_outputs(4283)));
    layer2_outputs(2745) <= (layer1_outputs(3644)) and (layer1_outputs(484));
    layer2_outputs(2746) <= layer1_outputs(249);
    layer2_outputs(2747) <= '0';
    layer2_outputs(2748) <= not(layer1_outputs(1522)) or (layer1_outputs(4154));
    layer2_outputs(2749) <= layer1_outputs(2001);
    layer2_outputs(2750) <= (layer1_outputs(3907)) and (layer1_outputs(506));
    layer2_outputs(2751) <= not(layer1_outputs(578)) or (layer1_outputs(269));
    layer2_outputs(2752) <= (layer1_outputs(1392)) and not (layer1_outputs(5031));
    layer2_outputs(2753) <= not((layer1_outputs(5116)) or (layer1_outputs(3104)));
    layer2_outputs(2754) <= (layer1_outputs(2680)) and not (layer1_outputs(3419));
    layer2_outputs(2755) <= layer1_outputs(499);
    layer2_outputs(2756) <= layer1_outputs(3890);
    layer2_outputs(2757) <= not((layer1_outputs(2846)) and (layer1_outputs(3966)));
    layer2_outputs(2758) <= '0';
    layer2_outputs(2759) <= layer1_outputs(1024);
    layer2_outputs(2760) <= (layer1_outputs(1183)) and (layer1_outputs(452));
    layer2_outputs(2761) <= (layer1_outputs(2315)) and (layer1_outputs(4469));
    layer2_outputs(2762) <= not(layer1_outputs(4894)) or (layer1_outputs(1801));
    layer2_outputs(2763) <= not(layer1_outputs(379)) or (layer1_outputs(2204));
    layer2_outputs(2764) <= layer1_outputs(3765);
    layer2_outputs(2765) <= not(layer1_outputs(2950)) or (layer1_outputs(938));
    layer2_outputs(2766) <= layer1_outputs(3518);
    layer2_outputs(2767) <= (layer1_outputs(1215)) and not (layer1_outputs(3187));
    layer2_outputs(2768) <= not(layer1_outputs(732));
    layer2_outputs(2769) <= layer1_outputs(3968);
    layer2_outputs(2770) <= (layer1_outputs(4310)) and (layer1_outputs(724));
    layer2_outputs(2771) <= not(layer1_outputs(4801)) or (layer1_outputs(2977));
    layer2_outputs(2772) <= layer1_outputs(143);
    layer2_outputs(2773) <= '1';
    layer2_outputs(2774) <= '0';
    layer2_outputs(2775) <= not(layer1_outputs(212)) or (layer1_outputs(3873));
    layer2_outputs(2776) <= layer1_outputs(2042);
    layer2_outputs(2777) <= layer1_outputs(3088);
    layer2_outputs(2778) <= not(layer1_outputs(854));
    layer2_outputs(2779) <= '1';
    layer2_outputs(2780) <= not(layer1_outputs(214)) or (layer1_outputs(1356));
    layer2_outputs(2781) <= layer1_outputs(3731);
    layer2_outputs(2782) <= not(layer1_outputs(1031)) or (layer1_outputs(3601));
    layer2_outputs(2783) <= not(layer1_outputs(2029)) or (layer1_outputs(159));
    layer2_outputs(2784) <= (layer1_outputs(146)) or (layer1_outputs(3675));
    layer2_outputs(2785) <= layer1_outputs(116);
    layer2_outputs(2786) <= layer1_outputs(2029);
    layer2_outputs(2787) <= layer1_outputs(1957);
    layer2_outputs(2788) <= not(layer1_outputs(1301));
    layer2_outputs(2789) <= not((layer1_outputs(1410)) or (layer1_outputs(1865)));
    layer2_outputs(2790) <= not((layer1_outputs(3017)) xor (layer1_outputs(2444)));
    layer2_outputs(2791) <= not(layer1_outputs(2472));
    layer2_outputs(2792) <= (layer1_outputs(667)) and (layer1_outputs(3676));
    layer2_outputs(2793) <= not(layer1_outputs(4246));
    layer2_outputs(2794) <= not(layer1_outputs(1992));
    layer2_outputs(2795) <= layer1_outputs(2252);
    layer2_outputs(2796) <= layer1_outputs(1316);
    layer2_outputs(2797) <= not((layer1_outputs(810)) or (layer1_outputs(1855)));
    layer2_outputs(2798) <= '1';
    layer2_outputs(2799) <= layer1_outputs(3148);
    layer2_outputs(2800) <= (layer1_outputs(3283)) and (layer1_outputs(823));
    layer2_outputs(2801) <= layer1_outputs(4492);
    layer2_outputs(2802) <= layer1_outputs(4328);
    layer2_outputs(2803) <= layer1_outputs(3861);
    layer2_outputs(2804) <= (layer1_outputs(220)) and (layer1_outputs(2764));
    layer2_outputs(2805) <= not(layer1_outputs(1835)) or (layer1_outputs(1499));
    layer2_outputs(2806) <= not(layer1_outputs(4858)) or (layer1_outputs(1247));
    layer2_outputs(2807) <= (layer1_outputs(2046)) and not (layer1_outputs(2335));
    layer2_outputs(2808) <= '0';
    layer2_outputs(2809) <= not(layer1_outputs(1277)) or (layer1_outputs(1502));
    layer2_outputs(2810) <= (layer1_outputs(1445)) xor (layer1_outputs(1071));
    layer2_outputs(2811) <= not(layer1_outputs(3780)) or (layer1_outputs(5083));
    layer2_outputs(2812) <= '0';
    layer2_outputs(2813) <= not((layer1_outputs(1943)) and (layer1_outputs(3824)));
    layer2_outputs(2814) <= (layer1_outputs(3235)) xor (layer1_outputs(132));
    layer2_outputs(2815) <= not(layer1_outputs(4684));
    layer2_outputs(2816) <= not(layer1_outputs(338)) or (layer1_outputs(250));
    layer2_outputs(2817) <= layer1_outputs(3677);
    layer2_outputs(2818) <= not((layer1_outputs(4264)) and (layer1_outputs(2351)));
    layer2_outputs(2819) <= not(layer1_outputs(2552));
    layer2_outputs(2820) <= not((layer1_outputs(3544)) or (layer1_outputs(4617)));
    layer2_outputs(2821) <= not((layer1_outputs(33)) or (layer1_outputs(135)));
    layer2_outputs(2822) <= (layer1_outputs(1360)) and not (layer1_outputs(2553));
    layer2_outputs(2823) <= not(layer1_outputs(4827)) or (layer1_outputs(4343));
    layer2_outputs(2824) <= not((layer1_outputs(4417)) or (layer1_outputs(3438)));
    layer2_outputs(2825) <= not(layer1_outputs(413));
    layer2_outputs(2826) <= '0';
    layer2_outputs(2827) <= '0';
    layer2_outputs(2828) <= layer1_outputs(244);
    layer2_outputs(2829) <= (layer1_outputs(1088)) and not (layer1_outputs(3896));
    layer2_outputs(2830) <= not(layer1_outputs(2590)) or (layer1_outputs(1132));
    layer2_outputs(2831) <= (layer1_outputs(2507)) and (layer1_outputs(4457));
    layer2_outputs(2832) <= not((layer1_outputs(5099)) or (layer1_outputs(4348)));
    layer2_outputs(2833) <= (layer1_outputs(4565)) and not (layer1_outputs(1269));
    layer2_outputs(2834) <= not(layer1_outputs(985)) or (layer1_outputs(4067));
    layer2_outputs(2835) <= not((layer1_outputs(4962)) and (layer1_outputs(3302)));
    layer2_outputs(2836) <= layer1_outputs(1716);
    layer2_outputs(2837) <= not(layer1_outputs(3649));
    layer2_outputs(2838) <= (layer1_outputs(3688)) or (layer1_outputs(4088));
    layer2_outputs(2839) <= not(layer1_outputs(3343));
    layer2_outputs(2840) <= not(layer1_outputs(3202));
    layer2_outputs(2841) <= not(layer1_outputs(657)) or (layer1_outputs(3315));
    layer2_outputs(2842) <= not(layer1_outputs(2531)) or (layer1_outputs(3282));
    layer2_outputs(2843) <= layer1_outputs(1458);
    layer2_outputs(2844) <= (layer1_outputs(3199)) or (layer1_outputs(1760));
    layer2_outputs(2845) <= (layer1_outputs(86)) and not (layer1_outputs(2582));
    layer2_outputs(2846) <= (layer1_outputs(1571)) or (layer1_outputs(1988));
    layer2_outputs(2847) <= not((layer1_outputs(4062)) and (layer1_outputs(368)));
    layer2_outputs(2848) <= (layer1_outputs(5039)) and (layer1_outputs(1909));
    layer2_outputs(2849) <= (layer1_outputs(4085)) and not (layer1_outputs(4434));
    layer2_outputs(2850) <= layer1_outputs(4443);
    layer2_outputs(2851) <= not(layer1_outputs(1936));
    layer2_outputs(2852) <= '1';
    layer2_outputs(2853) <= not((layer1_outputs(3507)) xor (layer1_outputs(2357)));
    layer2_outputs(2854) <= '0';
    layer2_outputs(2855) <= not(layer1_outputs(449));
    layer2_outputs(2856) <= (layer1_outputs(472)) and not (layer1_outputs(3458));
    layer2_outputs(2857) <= not(layer1_outputs(2244));
    layer2_outputs(2858) <= not(layer1_outputs(3217));
    layer2_outputs(2859) <= (layer1_outputs(3845)) and not (layer1_outputs(495));
    layer2_outputs(2860) <= '1';
    layer2_outputs(2861) <= (layer1_outputs(237)) and not (layer1_outputs(4275));
    layer2_outputs(2862) <= layer1_outputs(2361);
    layer2_outputs(2863) <= (layer1_outputs(5092)) and (layer1_outputs(2149));
    layer2_outputs(2864) <= not((layer1_outputs(1217)) or (layer1_outputs(2355)));
    layer2_outputs(2865) <= not((layer1_outputs(317)) or (layer1_outputs(2644)));
    layer2_outputs(2866) <= not(layer1_outputs(3807));
    layer2_outputs(2867) <= not(layer1_outputs(1660)) or (layer1_outputs(520));
    layer2_outputs(2868) <= not(layer1_outputs(475));
    layer2_outputs(2869) <= not(layer1_outputs(643));
    layer2_outputs(2870) <= '1';
    layer2_outputs(2871) <= layer1_outputs(1125);
    layer2_outputs(2872) <= not((layer1_outputs(1749)) or (layer1_outputs(2798)));
    layer2_outputs(2873) <= not((layer1_outputs(1468)) or (layer1_outputs(2170)));
    layer2_outputs(2874) <= not((layer1_outputs(2660)) and (layer1_outputs(2049)));
    layer2_outputs(2875) <= not(layer1_outputs(5074));
    layer2_outputs(2876) <= '0';
    layer2_outputs(2877) <= not(layer1_outputs(3314));
    layer2_outputs(2878) <= not(layer1_outputs(4660));
    layer2_outputs(2879) <= layer1_outputs(1670);
    layer2_outputs(2880) <= (layer1_outputs(2483)) and not (layer1_outputs(2879));
    layer2_outputs(2881) <= layer1_outputs(4265);
    layer2_outputs(2882) <= '0';
    layer2_outputs(2883) <= (layer1_outputs(387)) and (layer1_outputs(4395));
    layer2_outputs(2884) <= not(layer1_outputs(2466));
    layer2_outputs(2885) <= (layer1_outputs(3834)) and (layer1_outputs(4504));
    layer2_outputs(2886) <= (layer1_outputs(753)) and not (layer1_outputs(2135));
    layer2_outputs(2887) <= (layer1_outputs(4191)) or (layer1_outputs(1968));
    layer2_outputs(2888) <= (layer1_outputs(4142)) and not (layer1_outputs(4981));
    layer2_outputs(2889) <= '1';
    layer2_outputs(2890) <= '1';
    layer2_outputs(2891) <= not((layer1_outputs(4294)) and (layer1_outputs(2670)));
    layer2_outputs(2892) <= not(layer1_outputs(2109));
    layer2_outputs(2893) <= (layer1_outputs(2617)) and not (layer1_outputs(4594));
    layer2_outputs(2894) <= not(layer1_outputs(4669));
    layer2_outputs(2895) <= not(layer1_outputs(4164)) or (layer1_outputs(2166));
    layer2_outputs(2896) <= layer1_outputs(4821);
    layer2_outputs(2897) <= (layer1_outputs(897)) and (layer1_outputs(983));
    layer2_outputs(2898) <= not(layer1_outputs(2791)) or (layer1_outputs(138));
    layer2_outputs(2899) <= not(layer1_outputs(2234));
    layer2_outputs(2900) <= not(layer1_outputs(3629));
    layer2_outputs(2901) <= not(layer1_outputs(4825)) or (layer1_outputs(4183));
    layer2_outputs(2902) <= layer1_outputs(32);
    layer2_outputs(2903) <= not(layer1_outputs(4828));
    layer2_outputs(2904) <= '0';
    layer2_outputs(2905) <= layer1_outputs(1403);
    layer2_outputs(2906) <= not(layer1_outputs(2525)) or (layer1_outputs(4201));
    layer2_outputs(2907) <= (layer1_outputs(904)) and (layer1_outputs(1239));
    layer2_outputs(2908) <= '1';
    layer2_outputs(2909) <= '1';
    layer2_outputs(2910) <= not((layer1_outputs(3314)) xor (layer1_outputs(4699)));
    layer2_outputs(2911) <= (layer1_outputs(799)) and not (layer1_outputs(3735));
    layer2_outputs(2912) <= layer1_outputs(2358);
    layer2_outputs(2913) <= not(layer1_outputs(171)) or (layer1_outputs(1234));
    layer2_outputs(2914) <= not(layer1_outputs(4834));
    layer2_outputs(2915) <= (layer1_outputs(1863)) or (layer1_outputs(1824));
    layer2_outputs(2916) <= (layer1_outputs(3592)) and not (layer1_outputs(2924));
    layer2_outputs(2917) <= layer1_outputs(174);
    layer2_outputs(2918) <= not(layer1_outputs(424));
    layer2_outputs(2919) <= layer1_outputs(4344);
    layer2_outputs(2920) <= '0';
    layer2_outputs(2921) <= not(layer1_outputs(4156)) or (layer1_outputs(4054));
    layer2_outputs(2922) <= not(layer1_outputs(4875));
    layer2_outputs(2923) <= (layer1_outputs(955)) and not (layer1_outputs(5071));
    layer2_outputs(2924) <= not(layer1_outputs(4429));
    layer2_outputs(2925) <= layer1_outputs(3003);
    layer2_outputs(2926) <= '0';
    layer2_outputs(2927) <= (layer1_outputs(4574)) and not (layer1_outputs(3471));
    layer2_outputs(2928) <= (layer1_outputs(4967)) xor (layer1_outputs(2216));
    layer2_outputs(2929) <= not(layer1_outputs(1334));
    layer2_outputs(2930) <= '1';
    layer2_outputs(2931) <= (layer1_outputs(1971)) and not (layer1_outputs(144));
    layer2_outputs(2932) <= layer1_outputs(2378);
    layer2_outputs(2933) <= (layer1_outputs(3489)) and not (layer1_outputs(1108));
    layer2_outputs(2934) <= (layer1_outputs(2793)) and not (layer1_outputs(1389));
    layer2_outputs(2935) <= not(layer1_outputs(2304)) or (layer1_outputs(3035));
    layer2_outputs(2936) <= (layer1_outputs(3479)) and (layer1_outputs(3359));
    layer2_outputs(2937) <= not(layer1_outputs(1624));
    layer2_outputs(2938) <= (layer1_outputs(1909)) and not (layer1_outputs(769));
    layer2_outputs(2939) <= not(layer1_outputs(4667));
    layer2_outputs(2940) <= (layer1_outputs(3928)) and not (layer1_outputs(1215));
    layer2_outputs(2941) <= (layer1_outputs(2129)) and not (layer1_outputs(1575));
    layer2_outputs(2942) <= not((layer1_outputs(1740)) and (layer1_outputs(1799)));
    layer2_outputs(2943) <= not(layer1_outputs(52)) or (layer1_outputs(2948));
    layer2_outputs(2944) <= not(layer1_outputs(3012)) or (layer1_outputs(4041));
    layer2_outputs(2945) <= not(layer1_outputs(3060));
    layer2_outputs(2946) <= (layer1_outputs(4506)) and not (layer1_outputs(1413));
    layer2_outputs(2947) <= not(layer1_outputs(99));
    layer2_outputs(2948) <= (layer1_outputs(1190)) and (layer1_outputs(730));
    layer2_outputs(2949) <= (layer1_outputs(2591)) and not (layer1_outputs(3449));
    layer2_outputs(2950) <= (layer1_outputs(2615)) and (layer1_outputs(1438));
    layer2_outputs(2951) <= layer1_outputs(3330);
    layer2_outputs(2952) <= not((layer1_outputs(4612)) and (layer1_outputs(2636)));
    layer2_outputs(2953) <= '0';
    layer2_outputs(2954) <= not(layer1_outputs(2146));
    layer2_outputs(2955) <= not(layer1_outputs(5019)) or (layer1_outputs(1102));
    layer2_outputs(2956) <= layer1_outputs(4732);
    layer2_outputs(2957) <= not((layer1_outputs(3160)) and (layer1_outputs(4532)));
    layer2_outputs(2958) <= not(layer1_outputs(4359));
    layer2_outputs(2959) <= layer1_outputs(384);
    layer2_outputs(2960) <= '1';
    layer2_outputs(2961) <= layer1_outputs(2219);
    layer2_outputs(2962) <= '1';
    layer2_outputs(2963) <= not((layer1_outputs(2352)) and (layer1_outputs(3535)));
    layer2_outputs(2964) <= not(layer1_outputs(3936)) or (layer1_outputs(1843));
    layer2_outputs(2965) <= not(layer1_outputs(2407)) or (layer1_outputs(3907));
    layer2_outputs(2966) <= not(layer1_outputs(1320));
    layer2_outputs(2967) <= not((layer1_outputs(1945)) and (layer1_outputs(270)));
    layer2_outputs(2968) <= (layer1_outputs(5021)) and not (layer1_outputs(3266));
    layer2_outputs(2969) <= not(layer1_outputs(2428));
    layer2_outputs(2970) <= (layer1_outputs(3032)) xor (layer1_outputs(692));
    layer2_outputs(2971) <= layer1_outputs(5025);
    layer2_outputs(2972) <= layer1_outputs(1843);
    layer2_outputs(2973) <= not(layer1_outputs(2229));
    layer2_outputs(2974) <= (layer1_outputs(3071)) or (layer1_outputs(1117));
    layer2_outputs(2975) <= layer1_outputs(821);
    layer2_outputs(2976) <= layer1_outputs(880);
    layer2_outputs(2977) <= not(layer1_outputs(2325)) or (layer1_outputs(2121));
    layer2_outputs(2978) <= not(layer1_outputs(560)) or (layer1_outputs(709));
    layer2_outputs(2979) <= not((layer1_outputs(4475)) or (layer1_outputs(4968)));
    layer2_outputs(2980) <= not(layer1_outputs(4329));
    layer2_outputs(2981) <= not(layer1_outputs(3166)) or (layer1_outputs(2795));
    layer2_outputs(2982) <= (layer1_outputs(171)) and (layer1_outputs(3334));
    layer2_outputs(2983) <= (layer1_outputs(1805)) and not (layer1_outputs(5068));
    layer2_outputs(2984) <= (layer1_outputs(1990)) or (layer1_outputs(3845));
    layer2_outputs(2985) <= not((layer1_outputs(3574)) xor (layer1_outputs(4633)));
    layer2_outputs(2986) <= layer1_outputs(2382);
    layer2_outputs(2987) <= (layer1_outputs(2601)) and not (layer1_outputs(2749));
    layer2_outputs(2988) <= (layer1_outputs(2954)) and not (layer1_outputs(4453));
    layer2_outputs(2989) <= not(layer1_outputs(2980));
    layer2_outputs(2990) <= layer1_outputs(4861);
    layer2_outputs(2991) <= layer1_outputs(2983);
    layer2_outputs(2992) <= (layer1_outputs(2980)) and (layer1_outputs(674));
    layer2_outputs(2993) <= '0';
    layer2_outputs(2994) <= '1';
    layer2_outputs(2995) <= (layer1_outputs(2213)) and not (layer1_outputs(4715));
    layer2_outputs(2996) <= not((layer1_outputs(1148)) and (layer1_outputs(3192)));
    layer2_outputs(2997) <= not((layer1_outputs(2497)) or (layer1_outputs(3960)));
    layer2_outputs(2998) <= not(layer1_outputs(4397)) or (layer1_outputs(3312));
    layer2_outputs(2999) <= (layer1_outputs(3827)) and not (layer1_outputs(1494));
    layer2_outputs(3000) <= layer1_outputs(2027);
    layer2_outputs(3001) <= layer1_outputs(4770);
    layer2_outputs(3002) <= '1';
    layer2_outputs(3003) <= (layer1_outputs(3043)) and not (layer1_outputs(2035));
    layer2_outputs(3004) <= not(layer1_outputs(3490)) or (layer1_outputs(1288));
    layer2_outputs(3005) <= not(layer1_outputs(3373));
    layer2_outputs(3006) <= '1';
    layer2_outputs(3007) <= not((layer1_outputs(4998)) or (layer1_outputs(1874)));
    layer2_outputs(3008) <= not((layer1_outputs(3281)) or (layer1_outputs(4776)));
    layer2_outputs(3009) <= '1';
    layer2_outputs(3010) <= (layer1_outputs(1605)) or (layer1_outputs(3312));
    layer2_outputs(3011) <= not((layer1_outputs(3638)) or (layer1_outputs(1885)));
    layer2_outputs(3012) <= (layer1_outputs(4444)) or (layer1_outputs(1765));
    layer2_outputs(3013) <= '1';
    layer2_outputs(3014) <= (layer1_outputs(2470)) and (layer1_outputs(637));
    layer2_outputs(3015) <= not((layer1_outputs(2469)) and (layer1_outputs(3815)));
    layer2_outputs(3016) <= (layer1_outputs(3404)) or (layer1_outputs(4404));
    layer2_outputs(3017) <= not(layer1_outputs(4107));
    layer2_outputs(3018) <= '1';
    layer2_outputs(3019) <= not(layer1_outputs(308));
    layer2_outputs(3020) <= not(layer1_outputs(2018));
    layer2_outputs(3021) <= not(layer1_outputs(4782));
    layer2_outputs(3022) <= layer1_outputs(412);
    layer2_outputs(3023) <= (layer1_outputs(3972)) and (layer1_outputs(251));
    layer2_outputs(3024) <= not(layer1_outputs(4913));
    layer2_outputs(3025) <= (layer1_outputs(323)) or (layer1_outputs(1711));
    layer2_outputs(3026) <= '1';
    layer2_outputs(3027) <= layer1_outputs(886);
    layer2_outputs(3028) <= not((layer1_outputs(5087)) and (layer1_outputs(672)));
    layer2_outputs(3029) <= not((layer1_outputs(743)) and (layer1_outputs(80)));
    layer2_outputs(3030) <= '0';
    layer2_outputs(3031) <= not(layer1_outputs(1867)) or (layer1_outputs(961));
    layer2_outputs(3032) <= not((layer1_outputs(2706)) or (layer1_outputs(2025)));
    layer2_outputs(3033) <= (layer1_outputs(1911)) and not (layer1_outputs(1463));
    layer2_outputs(3034) <= layer1_outputs(3446);
    layer2_outputs(3035) <= layer1_outputs(3119);
    layer2_outputs(3036) <= layer1_outputs(3543);
    layer2_outputs(3037) <= not(layer1_outputs(2172));
    layer2_outputs(3038) <= layer1_outputs(4069);
    layer2_outputs(3039) <= (layer1_outputs(1012)) and (layer1_outputs(2573));
    layer2_outputs(3040) <= not(layer1_outputs(1540)) or (layer1_outputs(1024));
    layer2_outputs(3041) <= (layer1_outputs(341)) and (layer1_outputs(538));
    layer2_outputs(3042) <= (layer1_outputs(3524)) and (layer1_outputs(743));
    layer2_outputs(3043) <= (layer1_outputs(3237)) and not (layer1_outputs(3437));
    layer2_outputs(3044) <= (layer1_outputs(164)) and (layer1_outputs(2437));
    layer2_outputs(3045) <= not((layer1_outputs(1473)) or (layer1_outputs(2008)));
    layer2_outputs(3046) <= (layer1_outputs(471)) or (layer1_outputs(1331));
    layer2_outputs(3047) <= layer1_outputs(2679);
    layer2_outputs(3048) <= not((layer1_outputs(961)) and (layer1_outputs(2499)));
    layer2_outputs(3049) <= not((layer1_outputs(2649)) and (layer1_outputs(2919)));
    layer2_outputs(3050) <= layer1_outputs(768);
    layer2_outputs(3051) <= not((layer1_outputs(2397)) or (layer1_outputs(1106)));
    layer2_outputs(3052) <= (layer1_outputs(3009)) or (layer1_outputs(4915));
    layer2_outputs(3053) <= (layer1_outputs(2433)) and not (layer1_outputs(1011));
    layer2_outputs(3054) <= '1';
    layer2_outputs(3055) <= (layer1_outputs(3839)) or (layer1_outputs(120));
    layer2_outputs(3056) <= (layer1_outputs(3613)) and (layer1_outputs(2393));
    layer2_outputs(3057) <= not((layer1_outputs(456)) or (layer1_outputs(1455)));
    layer2_outputs(3058) <= (layer1_outputs(533)) or (layer1_outputs(3997));
    layer2_outputs(3059) <= not(layer1_outputs(3387)) or (layer1_outputs(982));
    layer2_outputs(3060) <= layer1_outputs(5083);
    layer2_outputs(3061) <= not((layer1_outputs(1851)) and (layer1_outputs(554)));
    layer2_outputs(3062) <= (layer1_outputs(286)) or (layer1_outputs(3208));
    layer2_outputs(3063) <= '1';
    layer2_outputs(3064) <= not(layer1_outputs(1985)) or (layer1_outputs(4529));
    layer2_outputs(3065) <= not(layer1_outputs(17));
    layer2_outputs(3066) <= not(layer1_outputs(836));
    layer2_outputs(3067) <= (layer1_outputs(163)) and (layer1_outputs(3287));
    layer2_outputs(3068) <= (layer1_outputs(1205)) and (layer1_outputs(103));
    layer2_outputs(3069) <= '0';
    layer2_outputs(3070) <= not(layer1_outputs(3334)) or (layer1_outputs(88));
    layer2_outputs(3071) <= (layer1_outputs(3735)) and not (layer1_outputs(236));
    layer2_outputs(3072) <= not(layer1_outputs(1818)) or (layer1_outputs(2568));
    layer2_outputs(3073) <= not(layer1_outputs(3076));
    layer2_outputs(3074) <= not(layer1_outputs(3385)) or (layer1_outputs(3606));
    layer2_outputs(3075) <= not(layer1_outputs(4115)) or (layer1_outputs(303));
    layer2_outputs(3076) <= (layer1_outputs(3623)) or (layer1_outputs(3077));
    layer2_outputs(3077) <= (layer1_outputs(178)) or (layer1_outputs(2258));
    layer2_outputs(3078) <= not(layer1_outputs(3181));
    layer2_outputs(3079) <= layer1_outputs(2492);
    layer2_outputs(3080) <= layer1_outputs(1185);
    layer2_outputs(3081) <= '0';
    layer2_outputs(3082) <= not((layer1_outputs(1588)) or (layer1_outputs(1031)));
    layer2_outputs(3083) <= not(layer1_outputs(931)) or (layer1_outputs(124));
    layer2_outputs(3084) <= '0';
    layer2_outputs(3085) <= (layer1_outputs(3765)) and (layer1_outputs(2176));
    layer2_outputs(3086) <= not(layer1_outputs(678)) or (layer1_outputs(1798));
    layer2_outputs(3087) <= not((layer1_outputs(1611)) xor (layer1_outputs(4543)));
    layer2_outputs(3088) <= (layer1_outputs(1098)) or (layer1_outputs(3867));
    layer2_outputs(3089) <= layer1_outputs(1557);
    layer2_outputs(3090) <= (layer1_outputs(3653)) and (layer1_outputs(565));
    layer2_outputs(3091) <= not(layer1_outputs(958));
    layer2_outputs(3092) <= not(layer1_outputs(433));
    layer2_outputs(3093) <= not(layer1_outputs(2241)) or (layer1_outputs(3737));
    layer2_outputs(3094) <= layer1_outputs(4207);
    layer2_outputs(3095) <= not(layer1_outputs(2693)) or (layer1_outputs(4447));
    layer2_outputs(3096) <= not(layer1_outputs(504));
    layer2_outputs(3097) <= '0';
    layer2_outputs(3098) <= (layer1_outputs(1249)) or (layer1_outputs(2863));
    layer2_outputs(3099) <= (layer1_outputs(4052)) and (layer1_outputs(391));
    layer2_outputs(3100) <= not(layer1_outputs(893)) or (layer1_outputs(1380));
    layer2_outputs(3101) <= '0';
    layer2_outputs(3102) <= '1';
    layer2_outputs(3103) <= not(layer1_outputs(565)) or (layer1_outputs(3113));
    layer2_outputs(3104) <= (layer1_outputs(532)) or (layer1_outputs(3030));
    layer2_outputs(3105) <= layer1_outputs(1923);
    layer2_outputs(3106) <= '1';
    layer2_outputs(3107) <= (layer1_outputs(3396)) or (layer1_outputs(4550));
    layer2_outputs(3108) <= not(layer1_outputs(3133)) or (layer1_outputs(1160));
    layer2_outputs(3109) <= (layer1_outputs(1040)) and not (layer1_outputs(4646));
    layer2_outputs(3110) <= layer1_outputs(1688);
    layer2_outputs(3111) <= not((layer1_outputs(4535)) and (layer1_outputs(1956)));
    layer2_outputs(3112) <= not(layer1_outputs(530));
    layer2_outputs(3113) <= '0';
    layer2_outputs(3114) <= not(layer1_outputs(2939));
    layer2_outputs(3115) <= (layer1_outputs(3635)) and not (layer1_outputs(2922));
    layer2_outputs(3116) <= layer1_outputs(3551);
    layer2_outputs(3117) <= not(layer1_outputs(1135)) or (layer1_outputs(2796));
    layer2_outputs(3118) <= '0';
    layer2_outputs(3119) <= not(layer1_outputs(3433)) or (layer1_outputs(4560));
    layer2_outputs(3120) <= layer1_outputs(295);
    layer2_outputs(3121) <= not((layer1_outputs(1394)) xor (layer1_outputs(3969)));
    layer2_outputs(3122) <= (layer1_outputs(2871)) and not (layer1_outputs(4598));
    layer2_outputs(3123) <= '0';
    layer2_outputs(3124) <= not((layer1_outputs(2476)) and (layer1_outputs(2229)));
    layer2_outputs(3125) <= not(layer1_outputs(3425));
    layer2_outputs(3126) <= not((layer1_outputs(4140)) and (layer1_outputs(4255)));
    layer2_outputs(3127) <= layer1_outputs(2372);
    layer2_outputs(3128) <= (layer1_outputs(1968)) and (layer1_outputs(4764));
    layer2_outputs(3129) <= not(layer1_outputs(1355));
    layer2_outputs(3130) <= layer1_outputs(2295);
    layer2_outputs(3131) <= layer1_outputs(505);
    layer2_outputs(3132) <= '0';
    layer2_outputs(3133) <= '0';
    layer2_outputs(3134) <= '0';
    layer2_outputs(3135) <= layer1_outputs(1775);
    layer2_outputs(3136) <= not(layer1_outputs(1554));
    layer2_outputs(3137) <= layer1_outputs(3353);
    layer2_outputs(3138) <= (layer1_outputs(4728)) or (layer1_outputs(1375));
    layer2_outputs(3139) <= layer1_outputs(538);
    layer2_outputs(3140) <= (layer1_outputs(1546)) and (layer1_outputs(3934));
    layer2_outputs(3141) <= not(layer1_outputs(4106)) or (layer1_outputs(1006));
    layer2_outputs(3142) <= not(layer1_outputs(2198));
    layer2_outputs(3143) <= (layer1_outputs(3942)) and (layer1_outputs(4558));
    layer2_outputs(3144) <= not(layer1_outputs(3866)) or (layer1_outputs(2725));
    layer2_outputs(3145) <= '1';
    layer2_outputs(3146) <= not(layer1_outputs(3564));
    layer2_outputs(3147) <= not(layer1_outputs(4677)) or (layer1_outputs(4615));
    layer2_outputs(3148) <= not((layer1_outputs(1541)) and (layer1_outputs(4330)));
    layer2_outputs(3149) <= not((layer1_outputs(1962)) or (layer1_outputs(1355)));
    layer2_outputs(3150) <= not(layer1_outputs(2541)) or (layer1_outputs(2779));
    layer2_outputs(3151) <= layer1_outputs(1178);
    layer2_outputs(3152) <= (layer1_outputs(4726)) and not (layer1_outputs(4921));
    layer2_outputs(3153) <= layer1_outputs(129);
    layer2_outputs(3154) <= (layer1_outputs(1255)) and not (layer1_outputs(1593));
    layer2_outputs(3155) <= not(layer1_outputs(320)) or (layer1_outputs(2604));
    layer2_outputs(3156) <= (layer1_outputs(1005)) and not (layer1_outputs(2531));
    layer2_outputs(3157) <= '1';
    layer2_outputs(3158) <= not(layer1_outputs(3663));
    layer2_outputs(3159) <= layer1_outputs(2107);
    layer2_outputs(3160) <= not((layer1_outputs(1698)) and (layer1_outputs(3841)));
    layer2_outputs(3161) <= not((layer1_outputs(2316)) xor (layer1_outputs(4471)));
    layer2_outputs(3162) <= not(layer1_outputs(3714)) or (layer1_outputs(1753));
    layer2_outputs(3163) <= not(layer1_outputs(715));
    layer2_outputs(3164) <= '1';
    layer2_outputs(3165) <= not(layer1_outputs(3844)) or (layer1_outputs(3367));
    layer2_outputs(3166) <= not(layer1_outputs(2281));
    layer2_outputs(3167) <= not(layer1_outputs(1819)) or (layer1_outputs(4456));
    layer2_outputs(3168) <= '0';
    layer2_outputs(3169) <= (layer1_outputs(4107)) xor (layer1_outputs(211));
    layer2_outputs(3170) <= (layer1_outputs(1114)) and not (layer1_outputs(4886));
    layer2_outputs(3171) <= not(layer1_outputs(2658));
    layer2_outputs(3172) <= not(layer1_outputs(2750)) or (layer1_outputs(3906));
    layer2_outputs(3173) <= layer1_outputs(419);
    layer2_outputs(3174) <= '1';
    layer2_outputs(3175) <= (layer1_outputs(2087)) and not (layer1_outputs(4776));
    layer2_outputs(3176) <= (layer1_outputs(4956)) or (layer1_outputs(4410));
    layer2_outputs(3177) <= (layer1_outputs(4506)) and (layer1_outputs(3609));
    layer2_outputs(3178) <= '1';
    layer2_outputs(3179) <= (layer1_outputs(1010)) and not (layer1_outputs(2443));
    layer2_outputs(3180) <= not((layer1_outputs(827)) or (layer1_outputs(3388)));
    layer2_outputs(3181) <= not(layer1_outputs(1132)) or (layer1_outputs(4794));
    layer2_outputs(3182) <= (layer1_outputs(2186)) and not (layer1_outputs(4312));
    layer2_outputs(3183) <= not(layer1_outputs(1258));
    layer2_outputs(3184) <= '0';
    layer2_outputs(3185) <= not(layer1_outputs(2853));
    layer2_outputs(3186) <= not(layer1_outputs(2761)) or (layer1_outputs(1668));
    layer2_outputs(3187) <= not((layer1_outputs(3866)) and (layer1_outputs(68)));
    layer2_outputs(3188) <= layer1_outputs(401);
    layer2_outputs(3189) <= (layer1_outputs(2618)) or (layer1_outputs(423));
    layer2_outputs(3190) <= not(layer1_outputs(2388));
    layer2_outputs(3191) <= (layer1_outputs(2369)) or (layer1_outputs(2992));
    layer2_outputs(3192) <= (layer1_outputs(3734)) and not (layer1_outputs(1786));
    layer2_outputs(3193) <= (layer1_outputs(1054)) and not (layer1_outputs(3664));
    layer2_outputs(3194) <= not((layer1_outputs(958)) xor (layer1_outputs(1051)));
    layer2_outputs(3195) <= layer1_outputs(3492);
    layer2_outputs(3196) <= '1';
    layer2_outputs(3197) <= not(layer1_outputs(3888)) or (layer1_outputs(661));
    layer2_outputs(3198) <= not(layer1_outputs(4627));
    layer2_outputs(3199) <= (layer1_outputs(4011)) xor (layer1_outputs(3264));
    layer2_outputs(3200) <= '1';
    layer2_outputs(3201) <= not(layer1_outputs(2354)) or (layer1_outputs(4312));
    layer2_outputs(3202) <= not((layer1_outputs(86)) or (layer1_outputs(3769)));
    layer2_outputs(3203) <= layer1_outputs(1663);
    layer2_outputs(3204) <= '1';
    layer2_outputs(3205) <= layer1_outputs(1261);
    layer2_outputs(3206) <= not(layer1_outputs(510)) or (layer1_outputs(1136));
    layer2_outputs(3207) <= not(layer1_outputs(4644));
    layer2_outputs(3208) <= not(layer1_outputs(4387));
    layer2_outputs(3209) <= '0';
    layer2_outputs(3210) <= '1';
    layer2_outputs(3211) <= not(layer1_outputs(4055));
    layer2_outputs(3212) <= (layer1_outputs(4114)) and not (layer1_outputs(1140));
    layer2_outputs(3213) <= (layer1_outputs(45)) and not (layer1_outputs(4692));
    layer2_outputs(3214) <= not(layer1_outputs(2380));
    layer2_outputs(3215) <= not(layer1_outputs(4279));
    layer2_outputs(3216) <= not(layer1_outputs(1661)) or (layer1_outputs(1389));
    layer2_outputs(3217) <= not(layer1_outputs(348));
    layer2_outputs(3218) <= (layer1_outputs(3858)) and not (layer1_outputs(1012));
    layer2_outputs(3219) <= (layer1_outputs(2716)) and not (layer1_outputs(1459));
    layer2_outputs(3220) <= not(layer1_outputs(2368));
    layer2_outputs(3221) <= not(layer1_outputs(3508)) or (layer1_outputs(2714));
    layer2_outputs(3222) <= layer1_outputs(4457);
    layer2_outputs(3223) <= layer1_outputs(2424);
    layer2_outputs(3224) <= (layer1_outputs(3165)) and not (layer1_outputs(760));
    layer2_outputs(3225) <= '0';
    layer2_outputs(3226) <= not((layer1_outputs(2869)) or (layer1_outputs(1357)));
    layer2_outputs(3227) <= not((layer1_outputs(4606)) and (layer1_outputs(3296)));
    layer2_outputs(3228) <= not(layer1_outputs(558)) or (layer1_outputs(1671));
    layer2_outputs(3229) <= not(layer1_outputs(3143));
    layer2_outputs(3230) <= (layer1_outputs(3925)) and not (layer1_outputs(1507));
    layer2_outputs(3231) <= '0';
    layer2_outputs(3232) <= not((layer1_outputs(4414)) and (layer1_outputs(1732)));
    layer2_outputs(3233) <= (layer1_outputs(1439)) and (layer1_outputs(1542));
    layer2_outputs(3234) <= not(layer1_outputs(1029)) or (layer1_outputs(3521));
    layer2_outputs(3235) <= not((layer1_outputs(3269)) and (layer1_outputs(3675)));
    layer2_outputs(3236) <= (layer1_outputs(1579)) and (layer1_outputs(3666));
    layer2_outputs(3237) <= not(layer1_outputs(4245)) or (layer1_outputs(1531));
    layer2_outputs(3238) <= layer1_outputs(3537);
    layer2_outputs(3239) <= not((layer1_outputs(2896)) and (layer1_outputs(4262)));
    layer2_outputs(3240) <= not(layer1_outputs(2715));
    layer2_outputs(3241) <= not(layer1_outputs(264)) or (layer1_outputs(4057));
    layer2_outputs(3242) <= not(layer1_outputs(4051)) or (layer1_outputs(1875));
    layer2_outputs(3243) <= layer1_outputs(1139);
    layer2_outputs(3244) <= not((layer1_outputs(292)) or (layer1_outputs(2424)));
    layer2_outputs(3245) <= '0';
    layer2_outputs(3246) <= (layer1_outputs(3073)) or (layer1_outputs(3356));
    layer2_outputs(3247) <= '0';
    layer2_outputs(3248) <= '1';
    layer2_outputs(3249) <= not(layer1_outputs(1340)) or (layer1_outputs(894));
    layer2_outputs(3250) <= layer1_outputs(1482);
    layer2_outputs(3251) <= (layer1_outputs(516)) or (layer1_outputs(4997));
    layer2_outputs(3252) <= (layer1_outputs(4830)) and not (layer1_outputs(1388));
    layer2_outputs(3253) <= (layer1_outputs(2927)) and (layer1_outputs(778));
    layer2_outputs(3254) <= not(layer1_outputs(199)) or (layer1_outputs(2174));
    layer2_outputs(3255) <= (layer1_outputs(1987)) and (layer1_outputs(3175));
    layer2_outputs(3256) <= layer1_outputs(95);
    layer2_outputs(3257) <= (layer1_outputs(2043)) xor (layer1_outputs(1111));
    layer2_outputs(3258) <= (layer1_outputs(3282)) and not (layer1_outputs(554));
    layer2_outputs(3259) <= not(layer1_outputs(1447)) or (layer1_outputs(3079));
    layer2_outputs(3260) <= not((layer1_outputs(1995)) and (layer1_outputs(2134)));
    layer2_outputs(3261) <= '0';
    layer2_outputs(3262) <= (layer1_outputs(2534)) and not (layer1_outputs(4493));
    layer2_outputs(3263) <= (layer1_outputs(546)) and (layer1_outputs(2082));
    layer2_outputs(3264) <= (layer1_outputs(2880)) or (layer1_outputs(486));
    layer2_outputs(3265) <= not(layer1_outputs(2886)) or (layer1_outputs(16));
    layer2_outputs(3266) <= (layer1_outputs(3321)) and not (layer1_outputs(1609));
    layer2_outputs(3267) <= (layer1_outputs(4250)) and not (layer1_outputs(3916));
    layer2_outputs(3268) <= (layer1_outputs(1950)) or (layer1_outputs(4840));
    layer2_outputs(3269) <= not((layer1_outputs(1666)) or (layer1_outputs(2855)));
    layer2_outputs(3270) <= not(layer1_outputs(2520));
    layer2_outputs(3271) <= (layer1_outputs(2126)) and (layer1_outputs(972));
    layer2_outputs(3272) <= (layer1_outputs(1592)) or (layer1_outputs(168));
    layer2_outputs(3273) <= layer1_outputs(2444);
    layer2_outputs(3274) <= not(layer1_outputs(3933)) or (layer1_outputs(879));
    layer2_outputs(3275) <= not(layer1_outputs(4229));
    layer2_outputs(3276) <= (layer1_outputs(2699)) and (layer1_outputs(3733));
    layer2_outputs(3277) <= not(layer1_outputs(2192));
    layer2_outputs(3278) <= not(layer1_outputs(2245));
    layer2_outputs(3279) <= '1';
    layer2_outputs(3280) <= not(layer1_outputs(3465));
    layer2_outputs(3281) <= '0';
    layer2_outputs(3282) <= not(layer1_outputs(2885)) or (layer1_outputs(1396));
    layer2_outputs(3283) <= (layer1_outputs(3849)) and not (layer1_outputs(3721));
    layer2_outputs(3284) <= not(layer1_outputs(2163));
    layer2_outputs(3285) <= '0';
    layer2_outputs(3286) <= layer1_outputs(2090);
    layer2_outputs(3287) <= '1';
    layer2_outputs(3288) <= not(layer1_outputs(4967));
    layer2_outputs(3289) <= not(layer1_outputs(4644)) or (layer1_outputs(951));
    layer2_outputs(3290) <= not(layer1_outputs(2533));
    layer2_outputs(3291) <= (layer1_outputs(4676)) and not (layer1_outputs(1576));
    layer2_outputs(3292) <= (layer1_outputs(3432)) xor (layer1_outputs(2408));
    layer2_outputs(3293) <= not(layer1_outputs(2283)) or (layer1_outputs(2909));
    layer2_outputs(3294) <= '1';
    layer2_outputs(3295) <= layer1_outputs(1759);
    layer2_outputs(3296) <= not(layer1_outputs(3617));
    layer2_outputs(3297) <= (layer1_outputs(844)) and (layer1_outputs(23));
    layer2_outputs(3298) <= layer1_outputs(959);
    layer2_outputs(3299) <= not((layer1_outputs(927)) or (layer1_outputs(2143)));
    layer2_outputs(3300) <= (layer1_outputs(22)) and not (layer1_outputs(3464));
    layer2_outputs(3301) <= not(layer1_outputs(4477));
    layer2_outputs(3302) <= not(layer1_outputs(3737));
    layer2_outputs(3303) <= (layer1_outputs(4847)) and not (layer1_outputs(4546));
    layer2_outputs(3304) <= layer1_outputs(518);
    layer2_outputs(3305) <= '1';
    layer2_outputs(3306) <= (layer1_outputs(4541)) and not (layer1_outputs(4993));
    layer2_outputs(3307) <= layer1_outputs(4625);
    layer2_outputs(3308) <= (layer1_outputs(4389)) and not (layer1_outputs(852));
    layer2_outputs(3309) <= not(layer1_outputs(1545)) or (layer1_outputs(4955));
    layer2_outputs(3310) <= (layer1_outputs(3636)) and (layer1_outputs(4550));
    layer2_outputs(3311) <= not(layer1_outputs(4149)) or (layer1_outputs(516));
    layer2_outputs(3312) <= not(layer1_outputs(2930));
    layer2_outputs(3313) <= not((layer1_outputs(4442)) or (layer1_outputs(2327)));
    layer2_outputs(3314) <= not(layer1_outputs(3830));
    layer2_outputs(3315) <= not(layer1_outputs(572)) or (layer1_outputs(4866));
    layer2_outputs(3316) <= not((layer1_outputs(2056)) and (layer1_outputs(1408)));
    layer2_outputs(3317) <= '0';
    layer2_outputs(3318) <= (layer1_outputs(2331)) or (layer1_outputs(4827));
    layer2_outputs(3319) <= (layer1_outputs(2340)) xor (layer1_outputs(1063));
    layer2_outputs(3320) <= not(layer1_outputs(1707));
    layer2_outputs(3321) <= not(layer1_outputs(4695)) or (layer1_outputs(4568));
    layer2_outputs(3322) <= layer1_outputs(3010);
    layer2_outputs(3323) <= '0';
    layer2_outputs(3324) <= not(layer1_outputs(3757));
    layer2_outputs(3325) <= '1';
    layer2_outputs(3326) <= layer1_outputs(688);
    layer2_outputs(3327) <= not(layer1_outputs(3442));
    layer2_outputs(3328) <= not((layer1_outputs(3400)) or (layer1_outputs(3434)));
    layer2_outputs(3329) <= not(layer1_outputs(1007));
    layer2_outputs(3330) <= not(layer1_outputs(1731));
    layer2_outputs(3331) <= (layer1_outputs(114)) or (layer1_outputs(4466));
    layer2_outputs(3332) <= (layer1_outputs(1118)) and (layer1_outputs(399));
    layer2_outputs(3333) <= '0';
    layer2_outputs(3334) <= not(layer1_outputs(1869)) or (layer1_outputs(2071));
    layer2_outputs(3335) <= not(layer1_outputs(2224)) or (layer1_outputs(59));
    layer2_outputs(3336) <= (layer1_outputs(1756)) and not (layer1_outputs(1646));
    layer2_outputs(3337) <= '1';
    layer2_outputs(3338) <= not(layer1_outputs(2626)) or (layer1_outputs(4745));
    layer2_outputs(3339) <= layer1_outputs(4932);
    layer2_outputs(3340) <= not((layer1_outputs(1303)) or (layer1_outputs(3506)));
    layer2_outputs(3341) <= '1';
    layer2_outputs(3342) <= (layer1_outputs(2999)) or (layer1_outputs(439));
    layer2_outputs(3343) <= '0';
    layer2_outputs(3344) <= (layer1_outputs(583)) and (layer1_outputs(2300));
    layer2_outputs(3345) <= (layer1_outputs(4897)) and (layer1_outputs(4754));
    layer2_outputs(3346) <= '0';
    layer2_outputs(3347) <= (layer1_outputs(984)) and not (layer1_outputs(4487));
    layer2_outputs(3348) <= not(layer1_outputs(4484)) or (layer1_outputs(4845));
    layer2_outputs(3349) <= layer1_outputs(2410);
    layer2_outputs(3350) <= '1';
    layer2_outputs(3351) <= not(layer1_outputs(3345)) or (layer1_outputs(3729));
    layer2_outputs(3352) <= (layer1_outputs(255)) and (layer1_outputs(3173));
    layer2_outputs(3353) <= not(layer1_outputs(4413));
    layer2_outputs(3354) <= layer1_outputs(5038);
    layer2_outputs(3355) <= (layer1_outputs(2373)) or (layer1_outputs(269));
    layer2_outputs(3356) <= not(layer1_outputs(2710));
    layer2_outputs(3357) <= layer1_outputs(2489);
    layer2_outputs(3358) <= not(layer1_outputs(4436));
    layer2_outputs(3359) <= (layer1_outputs(901)) and (layer1_outputs(3017));
    layer2_outputs(3360) <= layer1_outputs(935);
    layer2_outputs(3361) <= '0';
    layer2_outputs(3362) <= layer1_outputs(656);
    layer2_outputs(3363) <= layer1_outputs(2408);
    layer2_outputs(3364) <= (layer1_outputs(849)) and not (layer1_outputs(2688));
    layer2_outputs(3365) <= not(layer1_outputs(2961));
    layer2_outputs(3366) <= not((layer1_outputs(92)) or (layer1_outputs(1298)));
    layer2_outputs(3367) <= not(layer1_outputs(2445));
    layer2_outputs(3368) <= layer1_outputs(1563);
    layer2_outputs(3369) <= not((layer1_outputs(3025)) or (layer1_outputs(3393)));
    layer2_outputs(3370) <= not(layer1_outputs(4513));
    layer2_outputs(3371) <= '1';
    layer2_outputs(3372) <= (layer1_outputs(2487)) and not (layer1_outputs(2202));
    layer2_outputs(3373) <= '0';
    layer2_outputs(3374) <= not(layer1_outputs(587)) or (layer1_outputs(4756));
    layer2_outputs(3375) <= layer1_outputs(2769);
    layer2_outputs(3376) <= (layer1_outputs(2243)) and (layer1_outputs(2083));
    layer2_outputs(3377) <= not(layer1_outputs(296)) or (layer1_outputs(775));
    layer2_outputs(3378) <= (layer1_outputs(479)) and not (layer1_outputs(2974));
    layer2_outputs(3379) <= not(layer1_outputs(1076)) or (layer1_outputs(262));
    layer2_outputs(3380) <= not(layer1_outputs(1920));
    layer2_outputs(3381) <= layer1_outputs(4995);
    layer2_outputs(3382) <= (layer1_outputs(805)) and not (layer1_outputs(1530));
    layer2_outputs(3383) <= not(layer1_outputs(4741)) or (layer1_outputs(3050));
    layer2_outputs(3384) <= layer1_outputs(4165);
    layer2_outputs(3385) <= not((layer1_outputs(3233)) or (layer1_outputs(366)));
    layer2_outputs(3386) <= layer1_outputs(3663);
    layer2_outputs(3387) <= not(layer1_outputs(4073));
    layer2_outputs(3388) <= not((layer1_outputs(4781)) and (layer1_outputs(2033)));
    layer2_outputs(3389) <= '1';
    layer2_outputs(3390) <= not((layer1_outputs(2344)) or (layer1_outputs(4771)));
    layer2_outputs(3391) <= layer1_outputs(1573);
    layer2_outputs(3392) <= '1';
    layer2_outputs(3393) <= layer1_outputs(1571);
    layer2_outputs(3394) <= (layer1_outputs(2949)) and (layer1_outputs(673));
    layer2_outputs(3395) <= layer1_outputs(2971);
    layer2_outputs(3396) <= (layer1_outputs(365)) or (layer1_outputs(327));
    layer2_outputs(3397) <= not((layer1_outputs(4143)) and (layer1_outputs(731)));
    layer2_outputs(3398) <= not((layer1_outputs(2521)) and (layer1_outputs(1115)));
    layer2_outputs(3399) <= (layer1_outputs(2434)) and not (layer1_outputs(1284));
    layer2_outputs(3400) <= not(layer1_outputs(3266));
    layer2_outputs(3401) <= not(layer1_outputs(38)) or (layer1_outputs(2078));
    layer2_outputs(3402) <= not((layer1_outputs(3440)) and (layer1_outputs(41)));
    layer2_outputs(3403) <= not(layer1_outputs(4608));
    layer2_outputs(3404) <= (layer1_outputs(3713)) and (layer1_outputs(26));
    layer2_outputs(3405) <= layer1_outputs(3854);
    layer2_outputs(3406) <= '0';
    layer2_outputs(3407) <= not(layer1_outputs(1456)) or (layer1_outputs(1771));
    layer2_outputs(3408) <= not(layer1_outputs(564)) or (layer1_outputs(2308));
    layer2_outputs(3409) <= '0';
    layer2_outputs(3410) <= not(layer1_outputs(4353));
    layer2_outputs(3411) <= (layer1_outputs(5071)) or (layer1_outputs(2526));
    layer2_outputs(3412) <= (layer1_outputs(3068)) xor (layer1_outputs(3191));
    layer2_outputs(3413) <= (layer1_outputs(3673)) and not (layer1_outputs(1597));
    layer2_outputs(3414) <= not(layer1_outputs(4551));
    layer2_outputs(3415) <= (layer1_outputs(2258)) xor (layer1_outputs(4816));
    layer2_outputs(3416) <= not((layer1_outputs(4544)) or (layer1_outputs(5060)));
    layer2_outputs(3417) <= not(layer1_outputs(1681)) or (layer1_outputs(3640));
    layer2_outputs(3418) <= (layer1_outputs(200)) and not (layer1_outputs(2668));
    layer2_outputs(3419) <= layer1_outputs(2816);
    layer2_outputs(3420) <= (layer1_outputs(4678)) or (layer1_outputs(1285));
    layer2_outputs(3421) <= '0';
    layer2_outputs(3422) <= '0';
    layer2_outputs(3423) <= '0';
    layer2_outputs(3424) <= '1';
    layer2_outputs(3425) <= (layer1_outputs(3610)) and not (layer1_outputs(3572));
    layer2_outputs(3426) <= (layer1_outputs(293)) and not (layer1_outputs(41));
    layer2_outputs(3427) <= (layer1_outputs(449)) or (layer1_outputs(733));
    layer2_outputs(3428) <= layer1_outputs(4266);
    layer2_outputs(3429) <= '0';
    layer2_outputs(3430) <= not(layer1_outputs(190));
    layer2_outputs(3431) <= layer1_outputs(21);
    layer2_outputs(3432) <= not(layer1_outputs(362));
    layer2_outputs(3433) <= '1';
    layer2_outputs(3434) <= not(layer1_outputs(2880));
    layer2_outputs(3435) <= (layer1_outputs(4417)) or (layer1_outputs(3267));
    layer2_outputs(3436) <= not((layer1_outputs(1160)) and (layer1_outputs(4750)));
    layer2_outputs(3437) <= layer1_outputs(690);
    layer2_outputs(3438) <= (layer1_outputs(954)) and not (layer1_outputs(4348));
    layer2_outputs(3439) <= not((layer1_outputs(2452)) or (layer1_outputs(4053)));
    layer2_outputs(3440) <= layer1_outputs(923);
    layer2_outputs(3441) <= not(layer1_outputs(249));
    layer2_outputs(3442) <= (layer1_outputs(3979)) and not (layer1_outputs(411));
    layer2_outputs(3443) <= not(layer1_outputs(456)) or (layer1_outputs(1884));
    layer2_outputs(3444) <= not(layer1_outputs(2291));
    layer2_outputs(3445) <= not(layer1_outputs(969));
    layer2_outputs(3446) <= not((layer1_outputs(3023)) or (layer1_outputs(4037)));
    layer2_outputs(3447) <= '0';
    layer2_outputs(3448) <= '1';
    layer2_outputs(3449) <= (layer1_outputs(194)) and not (layer1_outputs(2630));
    layer2_outputs(3450) <= (layer1_outputs(3918)) and not (layer1_outputs(3634));
    layer2_outputs(3451) <= layer1_outputs(474);
    layer2_outputs(3452) <= layer1_outputs(2225);
    layer2_outputs(3453) <= layer1_outputs(4703);
    layer2_outputs(3454) <= layer1_outputs(2430);
    layer2_outputs(3455) <= not((layer1_outputs(3604)) and (layer1_outputs(1919)));
    layer2_outputs(3456) <= not(layer1_outputs(2758));
    layer2_outputs(3457) <= not((layer1_outputs(782)) or (layer1_outputs(3273)));
    layer2_outputs(3458) <= not(layer1_outputs(4669));
    layer2_outputs(3459) <= (layer1_outputs(3218)) and not (layer1_outputs(3680));
    layer2_outputs(3460) <= not(layer1_outputs(1419));
    layer2_outputs(3461) <= (layer1_outputs(1090)) and (layer1_outputs(1531));
    layer2_outputs(3462) <= not(layer1_outputs(4202)) or (layer1_outputs(1094));
    layer2_outputs(3463) <= '0';
    layer2_outputs(3464) <= '1';
    layer2_outputs(3465) <= not((layer1_outputs(1777)) or (layer1_outputs(71)));
    layer2_outputs(3466) <= layer1_outputs(122);
    layer2_outputs(3467) <= layer1_outputs(4742);
    layer2_outputs(3468) <= layer1_outputs(4798);
    layer2_outputs(3469) <= '0';
    layer2_outputs(3470) <= not(layer1_outputs(2104)) or (layer1_outputs(3332));
    layer2_outputs(3471) <= not(layer1_outputs(306)) or (layer1_outputs(2006));
    layer2_outputs(3472) <= not((layer1_outputs(2765)) xor (layer1_outputs(2599)));
    layer2_outputs(3473) <= (layer1_outputs(4409)) and (layer1_outputs(630));
    layer2_outputs(3474) <= (layer1_outputs(2047)) or (layer1_outputs(4396));
    layer2_outputs(3475) <= (layer1_outputs(4431)) or (layer1_outputs(2341));
    layer2_outputs(3476) <= '0';
    layer2_outputs(3477) <= not(layer1_outputs(2919)) or (layer1_outputs(1632));
    layer2_outputs(3478) <= not(layer1_outputs(4757));
    layer2_outputs(3479) <= (layer1_outputs(2837)) or (layer1_outputs(3542));
    layer2_outputs(3480) <= not((layer1_outputs(1217)) or (layer1_outputs(4608)));
    layer2_outputs(3481) <= (layer1_outputs(170)) or (layer1_outputs(4224));
    layer2_outputs(3482) <= not(layer1_outputs(2495)) or (layer1_outputs(3984));
    layer2_outputs(3483) <= (layer1_outputs(3196)) or (layer1_outputs(749));
    layer2_outputs(3484) <= '1';
    layer2_outputs(3485) <= layer1_outputs(1707);
    layer2_outputs(3486) <= (layer1_outputs(3900)) and not (layer1_outputs(521));
    layer2_outputs(3487) <= (layer1_outputs(2175)) and not (layer1_outputs(4293));
    layer2_outputs(3488) <= not((layer1_outputs(3216)) or (layer1_outputs(1550)));
    layer2_outputs(3489) <= layer1_outputs(3329);
    layer2_outputs(3490) <= layer1_outputs(1154);
    layer2_outputs(3491) <= not(layer1_outputs(1544));
    layer2_outputs(3492) <= '0';
    layer2_outputs(3493) <= (layer1_outputs(2052)) and not (layer1_outputs(1766));
    layer2_outputs(3494) <= not(layer1_outputs(4043)) or (layer1_outputs(4906));
    layer2_outputs(3495) <= not(layer1_outputs(1887));
    layer2_outputs(3496) <= layer1_outputs(210);
    layer2_outputs(3497) <= not((layer1_outputs(2282)) or (layer1_outputs(621)));
    layer2_outputs(3498) <= layer1_outputs(1871);
    layer2_outputs(3499) <= '0';
    layer2_outputs(3500) <= (layer1_outputs(853)) and not (layer1_outputs(3086));
    layer2_outputs(3501) <= not(layer1_outputs(1796));
    layer2_outputs(3502) <= layer1_outputs(680);
    layer2_outputs(3503) <= '1';
    layer2_outputs(3504) <= '1';
    layer2_outputs(3505) <= not((layer1_outputs(2671)) and (layer1_outputs(1709)));
    layer2_outputs(3506) <= '1';
    layer2_outputs(3507) <= (layer1_outputs(4833)) and not (layer1_outputs(4369));
    layer2_outputs(3508) <= (layer1_outputs(1933)) and not (layer1_outputs(3745));
    layer2_outputs(3509) <= not(layer1_outputs(4859));
    layer2_outputs(3510) <= not(layer1_outputs(908));
    layer2_outputs(3511) <= not((layer1_outputs(967)) xor (layer1_outputs(3764)));
    layer2_outputs(3512) <= (layer1_outputs(3703)) and not (layer1_outputs(4695));
    layer2_outputs(3513) <= (layer1_outputs(1535)) and (layer1_outputs(4342));
    layer2_outputs(3514) <= not((layer1_outputs(4137)) xor (layer1_outputs(4906)));
    layer2_outputs(3515) <= '0';
    layer2_outputs(3516) <= (layer1_outputs(509)) or (layer1_outputs(3455));
    layer2_outputs(3517) <= '0';
    layer2_outputs(3518) <= '1';
    layer2_outputs(3519) <= not((layer1_outputs(5088)) xor (layer1_outputs(4576)));
    layer2_outputs(3520) <= (layer1_outputs(4027)) and not (layer1_outputs(50));
    layer2_outputs(3521) <= (layer1_outputs(735)) and not (layer1_outputs(2040));
    layer2_outputs(3522) <= '1';
    layer2_outputs(3523) <= (layer1_outputs(557)) or (layer1_outputs(5118));
    layer2_outputs(3524) <= layer1_outputs(1671);
    layer2_outputs(3525) <= layer1_outputs(2784);
    layer2_outputs(3526) <= '0';
    layer2_outputs(3527) <= (layer1_outputs(3138)) and not (layer1_outputs(4977));
    layer2_outputs(3528) <= (layer1_outputs(2656)) and not (layer1_outputs(2874));
    layer2_outputs(3529) <= '0';
    layer2_outputs(3530) <= '1';
    layer2_outputs(3531) <= (layer1_outputs(1570)) and (layer1_outputs(4901));
    layer2_outputs(3532) <= (layer1_outputs(2567)) and not (layer1_outputs(279));
    layer2_outputs(3533) <= not(layer1_outputs(3888));
    layer2_outputs(3534) <= '0';
    layer2_outputs(3535) <= layer1_outputs(1008);
    layer2_outputs(3536) <= layer1_outputs(638);
    layer2_outputs(3537) <= not(layer1_outputs(335)) or (layer1_outputs(2798));
    layer2_outputs(3538) <= (layer1_outputs(49)) and not (layer1_outputs(118));
    layer2_outputs(3539) <= (layer1_outputs(4532)) or (layer1_outputs(3140));
    layer2_outputs(3540) <= not((layer1_outputs(1637)) and (layer1_outputs(371)));
    layer2_outputs(3541) <= not((layer1_outputs(4355)) or (layer1_outputs(2004)));
    layer2_outputs(3542) <= (layer1_outputs(271)) and not (layer1_outputs(380));
    layer2_outputs(3543) <= (layer1_outputs(3229)) or (layer1_outputs(2512));
    layer2_outputs(3544) <= (layer1_outputs(432)) and (layer1_outputs(99));
    layer2_outputs(3545) <= layer1_outputs(1687);
    layer2_outputs(3546) <= not(layer1_outputs(1804)) or (layer1_outputs(1752));
    layer2_outputs(3547) <= not((layer1_outputs(1174)) or (layer1_outputs(3795)));
    layer2_outputs(3548) <= not(layer1_outputs(1944));
    layer2_outputs(3549) <= (layer1_outputs(3244)) and (layer1_outputs(792));
    layer2_outputs(3550) <= layer1_outputs(4189);
    layer2_outputs(3551) <= not(layer1_outputs(459));
    layer2_outputs(3552) <= not(layer1_outputs(100));
    layer2_outputs(3553) <= layer1_outputs(2633);
    layer2_outputs(3554) <= not(layer1_outputs(4971));
    layer2_outputs(3555) <= not(layer1_outputs(1167)) or (layer1_outputs(1814));
    layer2_outputs(3556) <= '0';
    layer2_outputs(3557) <= '1';
    layer2_outputs(3558) <= '1';
    layer2_outputs(3559) <= not((layer1_outputs(4056)) and (layer1_outputs(551)));
    layer2_outputs(3560) <= '1';
    layer2_outputs(3561) <= '1';
    layer2_outputs(3562) <= not(layer1_outputs(4482));
    layer2_outputs(3563) <= not(layer1_outputs(2323));
    layer2_outputs(3564) <= not(layer1_outputs(165));
    layer2_outputs(3565) <= not(layer1_outputs(4449));
    layer2_outputs(3566) <= (layer1_outputs(2311)) and (layer1_outputs(4227));
    layer2_outputs(3567) <= not(layer1_outputs(4864)) or (layer1_outputs(2711));
    layer2_outputs(3568) <= not((layer1_outputs(5038)) or (layer1_outputs(815)));
    layer2_outputs(3569) <= (layer1_outputs(4007)) xor (layer1_outputs(3153));
    layer2_outputs(3570) <= not(layer1_outputs(4641)) or (layer1_outputs(708));
    layer2_outputs(3571) <= not(layer1_outputs(1642));
    layer2_outputs(3572) <= layer1_outputs(794);
    layer2_outputs(3573) <= layer1_outputs(4540);
    layer2_outputs(3574) <= not(layer1_outputs(1268));
    layer2_outputs(3575) <= (layer1_outputs(2073)) or (layer1_outputs(4896));
    layer2_outputs(3576) <= (layer1_outputs(485)) and not (layer1_outputs(4935));
    layer2_outputs(3577) <= layer1_outputs(4228);
    layer2_outputs(3578) <= (layer1_outputs(144)) and not (layer1_outputs(5115));
    layer2_outputs(3579) <= not((layer1_outputs(2218)) and (layer1_outputs(843)));
    layer2_outputs(3580) <= '0';
    layer2_outputs(3581) <= not(layer1_outputs(3489));
    layer2_outputs(3582) <= not((layer1_outputs(4610)) and (layer1_outputs(3430)));
    layer2_outputs(3583) <= '0';
    layer2_outputs(3584) <= not(layer1_outputs(1790));
    layer2_outputs(3585) <= layer1_outputs(1345);
    layer2_outputs(3586) <= layer1_outputs(847);
    layer2_outputs(3587) <= (layer1_outputs(1152)) and not (layer1_outputs(3730));
    layer2_outputs(3588) <= not((layer1_outputs(4980)) or (layer1_outputs(1959)));
    layer2_outputs(3589) <= layer1_outputs(2124);
    layer2_outputs(3590) <= '1';
    layer2_outputs(3591) <= (layer1_outputs(4377)) and (layer1_outputs(4530));
    layer2_outputs(3592) <= '1';
    layer2_outputs(3593) <= not(layer1_outputs(3303)) or (layer1_outputs(4254));
    layer2_outputs(3594) <= not(layer1_outputs(364)) or (layer1_outputs(301));
    layer2_outputs(3595) <= not(layer1_outputs(4514));
    layer2_outputs(3596) <= (layer1_outputs(519)) and not (layer1_outputs(4283));
    layer2_outputs(3597) <= (layer1_outputs(1315)) or (layer1_outputs(1636));
    layer2_outputs(3598) <= not(layer1_outputs(4047)) or (layer1_outputs(2520));
    layer2_outputs(3599) <= not(layer1_outputs(4784));
    layer2_outputs(3600) <= not(layer1_outputs(3894)) or (layer1_outputs(4098));
    layer2_outputs(3601) <= (layer1_outputs(1788)) or (layer1_outputs(1645));
    layer2_outputs(3602) <= not(layer1_outputs(259));
    layer2_outputs(3603) <= '0';
    layer2_outputs(3604) <= not(layer1_outputs(2179));
    layer2_outputs(3605) <= (layer1_outputs(1200)) and (layer1_outputs(2924));
    layer2_outputs(3606) <= not(layer1_outputs(1322)) or (layer1_outputs(3600));
    layer2_outputs(3607) <= '1';
    layer2_outputs(3608) <= not(layer1_outputs(4540)) or (layer1_outputs(3186));
    layer2_outputs(3609) <= '1';
    layer2_outputs(3610) <= (layer1_outputs(1572)) and not (layer1_outputs(3137));
    layer2_outputs(3611) <= not(layer1_outputs(4135)) or (layer1_outputs(809));
    layer2_outputs(3612) <= not((layer1_outputs(1359)) and (layer1_outputs(1533)));
    layer2_outputs(3613) <= layer1_outputs(3853);
    layer2_outputs(3614) <= '0';
    layer2_outputs(3615) <= '1';
    layer2_outputs(3616) <= (layer1_outputs(3046)) and not (layer1_outputs(2197));
    layer2_outputs(3617) <= not(layer1_outputs(671));
    layer2_outputs(3618) <= not((layer1_outputs(3551)) and (layer1_outputs(1114)));
    layer2_outputs(3619) <= (layer1_outputs(3724)) or (layer1_outputs(3210));
    layer2_outputs(3620) <= layer1_outputs(181);
    layer2_outputs(3621) <= '0';
    layer2_outputs(3622) <= '0';
    layer2_outputs(3623) <= (layer1_outputs(4860)) and (layer1_outputs(550));
    layer2_outputs(3624) <= '1';
    layer2_outputs(3625) <= '0';
    layer2_outputs(3626) <= '1';
    layer2_outputs(3627) <= (layer1_outputs(952)) and (layer1_outputs(4080));
    layer2_outputs(3628) <= (layer1_outputs(1857)) and (layer1_outputs(2572));
    layer2_outputs(3629) <= not(layer1_outputs(4577));
    layer2_outputs(3630) <= not((layer1_outputs(3930)) and (layer1_outputs(4508)));
    layer2_outputs(3631) <= not(layer1_outputs(3369));
    layer2_outputs(3632) <= not(layer1_outputs(4954));
    layer2_outputs(3633) <= not(layer1_outputs(2873)) or (layer1_outputs(2329));
    layer2_outputs(3634) <= (layer1_outputs(3882)) and not (layer1_outputs(3961));
    layer2_outputs(3635) <= not(layer1_outputs(1574));
    layer2_outputs(3636) <= not((layer1_outputs(2675)) or (layer1_outputs(1424)));
    layer2_outputs(3637) <= not(layer1_outputs(3862));
    layer2_outputs(3638) <= not((layer1_outputs(3904)) or (layer1_outputs(4163)));
    layer2_outputs(3639) <= not(layer1_outputs(3865));
    layer2_outputs(3640) <= '1';
    layer2_outputs(3641) <= (layer1_outputs(820)) and not (layer1_outputs(3602));
    layer2_outputs(3642) <= '0';
    layer2_outputs(3643) <= '0';
    layer2_outputs(3644) <= not(layer1_outputs(736));
    layer2_outputs(3645) <= layer1_outputs(1774);
    layer2_outputs(3646) <= not(layer1_outputs(2865)) or (layer1_outputs(3396));
    layer2_outputs(3647) <= not((layer1_outputs(3596)) or (layer1_outputs(3034)));
    layer2_outputs(3648) <= not((layer1_outputs(926)) or (layer1_outputs(3883)));
    layer2_outputs(3649) <= not(layer1_outputs(2005));
    layer2_outputs(3650) <= (layer1_outputs(2957)) and not (layer1_outputs(4815));
    layer2_outputs(3651) <= (layer1_outputs(1456)) and not (layer1_outputs(1065));
    layer2_outputs(3652) <= layer1_outputs(2392);
    layer2_outputs(3653) <= (layer1_outputs(4361)) and not (layer1_outputs(3662));
    layer2_outputs(3654) <= not(layer1_outputs(2482));
    layer2_outputs(3655) <= layer1_outputs(4169);
    layer2_outputs(3656) <= not(layer1_outputs(1580));
    layer2_outputs(3657) <= not((layer1_outputs(2201)) or (layer1_outputs(2518)));
    layer2_outputs(3658) <= not(layer1_outputs(3519));
    layer2_outputs(3659) <= '1';
    layer2_outputs(3660) <= '0';
    layer2_outputs(3661) <= '0';
    layer2_outputs(3662) <= (layer1_outputs(64)) or (layer1_outputs(373));
    layer2_outputs(3663) <= not(layer1_outputs(3240));
    layer2_outputs(3664) <= (layer1_outputs(245)) or (layer1_outputs(3895));
    layer2_outputs(3665) <= '1';
    layer2_outputs(3666) <= '1';
    layer2_outputs(3667) <= layer1_outputs(1398);
    layer2_outputs(3668) <= layer1_outputs(1333);
    layer2_outputs(3669) <= not(layer1_outputs(4267));
    layer2_outputs(3670) <= not(layer1_outputs(4887));
    layer2_outputs(3671) <= (layer1_outputs(722)) and not (layer1_outputs(3978));
    layer2_outputs(3672) <= layer1_outputs(4238);
    layer2_outputs(3673) <= not(layer1_outputs(1727));
    layer2_outputs(3674) <= not(layer1_outputs(3583)) or (layer1_outputs(4852));
    layer2_outputs(3675) <= not((layer1_outputs(3484)) or (layer1_outputs(2849)));
    layer2_outputs(3676) <= '1';
    layer2_outputs(3677) <= layer1_outputs(4941);
    layer2_outputs(3678) <= (layer1_outputs(2289)) and not (layer1_outputs(2534));
    layer2_outputs(3679) <= not(layer1_outputs(3251)) or (layer1_outputs(3722));
    layer2_outputs(3680) <= '1';
    layer2_outputs(3681) <= layer1_outputs(3353);
    layer2_outputs(3682) <= (layer1_outputs(3437)) and not (layer1_outputs(2030));
    layer2_outputs(3683) <= '0';
    layer2_outputs(3684) <= layer1_outputs(2360);
    layer2_outputs(3685) <= layer1_outputs(4731);
    layer2_outputs(3686) <= not(layer1_outputs(917));
    layer2_outputs(3687) <= '1';
    layer2_outputs(3688) <= not((layer1_outputs(1936)) or (layer1_outputs(2502)));
    layer2_outputs(3689) <= not(layer1_outputs(4330)) or (layer1_outputs(4300));
    layer2_outputs(3690) <= (layer1_outputs(433)) and (layer1_outputs(3433));
    layer2_outputs(3691) <= (layer1_outputs(4453)) and not (layer1_outputs(1296));
    layer2_outputs(3692) <= not(layer1_outputs(2449));
    layer2_outputs(3693) <= (layer1_outputs(4260)) and (layer1_outputs(1685));
    layer2_outputs(3694) <= (layer1_outputs(1462)) or (layer1_outputs(1839));
    layer2_outputs(3695) <= (layer1_outputs(4750)) and not (layer1_outputs(2458));
    layer2_outputs(3696) <= not(layer1_outputs(5034));
    layer2_outputs(3697) <= not((layer1_outputs(1309)) or (layer1_outputs(3413)));
    layer2_outputs(3698) <= '1';
    layer2_outputs(3699) <= not(layer1_outputs(3708)) or (layer1_outputs(172));
    layer2_outputs(3700) <= '1';
    layer2_outputs(3701) <= (layer1_outputs(2960)) and (layer1_outputs(2920));
    layer2_outputs(3702) <= (layer1_outputs(3298)) or (layer1_outputs(3761));
    layer2_outputs(3703) <= not(layer1_outputs(4931));
    layer2_outputs(3704) <= '0';
    layer2_outputs(3705) <= not(layer1_outputs(3712)) or (layer1_outputs(3239));
    layer2_outputs(3706) <= '1';
    layer2_outputs(3707) <= layer1_outputs(2732);
    layer2_outputs(3708) <= not((layer1_outputs(5104)) and (layer1_outputs(536)));
    layer2_outputs(3709) <= not(layer1_outputs(2310)) or (layer1_outputs(4316));
    layer2_outputs(3710) <= not(layer1_outputs(1347)) or (layer1_outputs(652));
    layer2_outputs(3711) <= (layer1_outputs(3339)) and not (layer1_outputs(1182));
    layer2_outputs(3712) <= not(layer1_outputs(2465));
    layer2_outputs(3713) <= layer1_outputs(643);
    layer2_outputs(3714) <= (layer1_outputs(2498)) and not (layer1_outputs(3419));
    layer2_outputs(3715) <= layer1_outputs(2171);
    layer2_outputs(3716) <= '1';
    layer2_outputs(3717) <= (layer1_outputs(5005)) and (layer1_outputs(3093));
    layer2_outputs(3718) <= not(layer1_outputs(2318));
    layer2_outputs(3719) <= '0';
    layer2_outputs(3720) <= not(layer1_outputs(3239));
    layer2_outputs(3721) <= layer1_outputs(3331);
    layer2_outputs(3722) <= not(layer1_outputs(4202));
    layer2_outputs(3723) <= (layer1_outputs(1519)) and not (layer1_outputs(4229));
    layer2_outputs(3724) <= (layer1_outputs(3345)) and (layer1_outputs(2385));
    layer2_outputs(3725) <= not(layer1_outputs(4463));
    layer2_outputs(3726) <= '0';
    layer2_outputs(3727) <= '1';
    layer2_outputs(3728) <= not(layer1_outputs(2083));
    layer2_outputs(3729) <= layer1_outputs(910);
    layer2_outputs(3730) <= '1';
    layer2_outputs(3731) <= '0';
    layer2_outputs(3732) <= not(layer1_outputs(2751));
    layer2_outputs(3733) <= not((layer1_outputs(4217)) and (layer1_outputs(3369)));
    layer2_outputs(3734) <= not((layer1_outputs(1542)) and (layer1_outputs(167)));
    layer2_outputs(3735) <= (layer1_outputs(1768)) and (layer1_outputs(4501));
    layer2_outputs(3736) <= not(layer1_outputs(4105));
    layer2_outputs(3737) <= '1';
    layer2_outputs(3738) <= '1';
    layer2_outputs(3739) <= '1';
    layer2_outputs(3740) <= (layer1_outputs(2453)) or (layer1_outputs(4290));
    layer2_outputs(3741) <= (layer1_outputs(4904)) and not (layer1_outputs(2377));
    layer2_outputs(3742) <= not(layer1_outputs(1371));
    layer2_outputs(3743) <= '1';
    layer2_outputs(3744) <= layer1_outputs(1644);
    layer2_outputs(3745) <= not(layer1_outputs(2812));
    layer2_outputs(3746) <= (layer1_outputs(745)) and not (layer1_outputs(4585));
    layer2_outputs(3747) <= not(layer1_outputs(3915));
    layer2_outputs(3748) <= (layer1_outputs(787)) or (layer1_outputs(4004));
    layer2_outputs(3749) <= '0';
    layer2_outputs(3750) <= (layer1_outputs(487)) and not (layer1_outputs(2868));
    layer2_outputs(3751) <= not(layer1_outputs(2666)) or (layer1_outputs(2851));
    layer2_outputs(3752) <= layer1_outputs(4846);
    layer2_outputs(3753) <= '1';
    layer2_outputs(3754) <= '0';
    layer2_outputs(3755) <= (layer1_outputs(543)) or (layer1_outputs(3633));
    layer2_outputs(3756) <= not(layer1_outputs(2898)) or (layer1_outputs(2975));
    layer2_outputs(3757) <= '1';
    layer2_outputs(3758) <= layer1_outputs(3885);
    layer2_outputs(3759) <= not((layer1_outputs(65)) xor (layer1_outputs(2095)));
    layer2_outputs(3760) <= not(layer1_outputs(4197));
    layer2_outputs(3761) <= layer1_outputs(1212);
    layer2_outputs(3762) <= layer1_outputs(315);
    layer2_outputs(3763) <= (layer1_outputs(80)) and (layer1_outputs(4598));
    layer2_outputs(3764) <= not((layer1_outputs(2684)) and (layer1_outputs(4480)));
    layer2_outputs(3765) <= layer1_outputs(3581);
    layer2_outputs(3766) <= not(layer1_outputs(1198)) or (layer1_outputs(3943));
    layer2_outputs(3767) <= not(layer1_outputs(3857)) or (layer1_outputs(2343));
    layer2_outputs(3768) <= '1';
    layer2_outputs(3769) <= layer1_outputs(3275);
    layer2_outputs(3770) <= (layer1_outputs(441)) or (layer1_outputs(3293));
    layer2_outputs(3771) <= not(layer1_outputs(527)) or (layer1_outputs(4296));
    layer2_outputs(3772) <= layer1_outputs(1050);
    layer2_outputs(3773) <= not((layer1_outputs(501)) or (layer1_outputs(4676)));
    layer2_outputs(3774) <= not((layer1_outputs(3228)) or (layer1_outputs(2016)));
    layer2_outputs(3775) <= not(layer1_outputs(4786)) or (layer1_outputs(1047));
    layer2_outputs(3776) <= '1';
    layer2_outputs(3777) <= (layer1_outputs(4505)) and not (layer1_outputs(1115));
    layer2_outputs(3778) <= (layer1_outputs(1970)) and not (layer1_outputs(3307));
    layer2_outputs(3779) <= not(layer1_outputs(2330));
    layer2_outputs(3780) <= not(layer1_outputs(2832)) or (layer1_outputs(2545));
    layer2_outputs(3781) <= layer1_outputs(1301);
    layer2_outputs(3782) <= (layer1_outputs(1061)) and not (layer1_outputs(2009));
    layer2_outputs(3783) <= not((layer1_outputs(3086)) and (layer1_outputs(161)));
    layer2_outputs(3784) <= '0';
    layer2_outputs(3785) <= not(layer1_outputs(3770)) or (layer1_outputs(298));
    layer2_outputs(3786) <= not(layer1_outputs(4835));
    layer2_outputs(3787) <= not(layer1_outputs(1770));
    layer2_outputs(3788) <= not((layer1_outputs(3294)) and (layer1_outputs(592)));
    layer2_outputs(3789) <= layer1_outputs(4856);
    layer2_outputs(3790) <= not((layer1_outputs(1662)) or (layer1_outputs(37)));
    layer2_outputs(3791) <= (layer1_outputs(4867)) or (layer1_outputs(4155));
    layer2_outputs(3792) <= not(layer1_outputs(4321)) or (layer1_outputs(1608));
    layer2_outputs(3793) <= (layer1_outputs(2844)) and not (layer1_outputs(3319));
    layer2_outputs(3794) <= not(layer1_outputs(1435)) or (layer1_outputs(1701));
    layer2_outputs(3795) <= layer1_outputs(2318);
    layer2_outputs(3796) <= layer1_outputs(1397);
    layer2_outputs(3797) <= layer1_outputs(2630);
    layer2_outputs(3798) <= not(layer1_outputs(2532)) or (layer1_outputs(560));
    layer2_outputs(3799) <= (layer1_outputs(5067)) and not (layer1_outputs(3947));
    layer2_outputs(3800) <= not(layer1_outputs(3790)) or (layer1_outputs(3788));
    layer2_outputs(3801) <= not((layer1_outputs(2876)) and (layer1_outputs(1196)));
    layer2_outputs(3802) <= (layer1_outputs(4723)) or (layer1_outputs(2292));
    layer2_outputs(3803) <= '0';
    layer2_outputs(3804) <= not(layer1_outputs(1590)) or (layer1_outputs(839));
    layer2_outputs(3805) <= '1';
    layer2_outputs(3806) <= (layer1_outputs(3946)) and not (layer1_outputs(1441));
    layer2_outputs(3807) <= not(layer1_outputs(1053));
    layer2_outputs(3808) <= (layer1_outputs(1260)) and not (layer1_outputs(2723));
    layer2_outputs(3809) <= not(layer1_outputs(42));
    layer2_outputs(3810) <= (layer1_outputs(475)) and not (layer1_outputs(3587));
    layer2_outputs(3811) <= not((layer1_outputs(160)) or (layer1_outputs(2862)));
    layer2_outputs(3812) <= (layer1_outputs(3541)) or (layer1_outputs(387));
    layer2_outputs(3813) <= '0';
    layer2_outputs(3814) <= (layer1_outputs(1941)) or (layer1_outputs(1626));
    layer2_outputs(3815) <= not(layer1_outputs(5081)) or (layer1_outputs(1595));
    layer2_outputs(3816) <= layer1_outputs(1263);
    layer2_outputs(3817) <= '0';
    layer2_outputs(3818) <= (layer1_outputs(4026)) and (layer1_outputs(4657));
    layer2_outputs(3819) <= (layer1_outputs(2207)) and not (layer1_outputs(4340));
    layer2_outputs(3820) <= layer1_outputs(4299);
    layer2_outputs(3821) <= (layer1_outputs(2754)) and not (layer1_outputs(601));
    layer2_outputs(3822) <= not((layer1_outputs(1444)) or (layer1_outputs(2503)));
    layer2_outputs(3823) <= '1';
    layer2_outputs(3824) <= '1';
    layer2_outputs(3825) <= '1';
    layer2_outputs(3826) <= layer1_outputs(3219);
    layer2_outputs(3827) <= not(layer1_outputs(4322)) or (layer1_outputs(3477));
    layer2_outputs(3828) <= not(layer1_outputs(3968));
    layer2_outputs(3829) <= layer1_outputs(4590);
    layer2_outputs(3830) <= not((layer1_outputs(4529)) and (layer1_outputs(1926)));
    layer2_outputs(3831) <= not(layer1_outputs(1149));
    layer2_outputs(3832) <= not((layer1_outputs(104)) xor (layer1_outputs(2273)));
    layer2_outputs(3833) <= '1';
    layer2_outputs(3834) <= '1';
    layer2_outputs(3835) <= (layer1_outputs(1244)) or (layer1_outputs(5117));
    layer2_outputs(3836) <= not(layer1_outputs(3101)) or (layer1_outputs(914));
    layer2_outputs(3837) <= not(layer1_outputs(4775)) or (layer1_outputs(1232));
    layer2_outputs(3838) <= not(layer1_outputs(1128));
    layer2_outputs(3839) <= (layer1_outputs(2314)) and (layer1_outputs(4519));
    layer2_outputs(3840) <= layer1_outputs(4748);
    layer2_outputs(3841) <= layer1_outputs(287);
    layer2_outputs(3842) <= not((layer1_outputs(3091)) or (layer1_outputs(4738)));
    layer2_outputs(3843) <= layer1_outputs(1999);
    layer2_outputs(3844) <= not(layer1_outputs(4200));
    layer2_outputs(3845) <= '0';
    layer2_outputs(3846) <= layer1_outputs(1745);
    layer2_outputs(3847) <= not(layer1_outputs(1238));
    layer2_outputs(3848) <= (layer1_outputs(3919)) and not (layer1_outputs(4357));
    layer2_outputs(3849) <= (layer1_outputs(2719)) and not (layer1_outputs(17));
    layer2_outputs(3850) <= layer1_outputs(1733);
    layer2_outputs(3851) <= (layer1_outputs(1816)) or (layer1_outputs(2187));
    layer2_outputs(3852) <= (layer1_outputs(4703)) and not (layer1_outputs(1216));
    layer2_outputs(3853) <= layer1_outputs(2270);
    layer2_outputs(3854) <= not(layer1_outputs(3100)) or (layer1_outputs(1377));
    layer2_outputs(3855) <= (layer1_outputs(1452)) and not (layer1_outputs(1466));
    layer2_outputs(3856) <= (layer1_outputs(2286)) xor (layer1_outputs(4436));
    layer2_outputs(3857) <= '1';
    layer2_outputs(3858) <= not((layer1_outputs(3116)) and (layer1_outputs(3950)));
    layer2_outputs(3859) <= not(layer1_outputs(3915));
    layer2_outputs(3860) <= not(layer1_outputs(69)) or (layer1_outputs(386));
    layer2_outputs(3861) <= not(layer1_outputs(2925)) or (layer1_outputs(598));
    layer2_outputs(3862) <= not(layer1_outputs(1302));
    layer2_outputs(3863) <= not(layer1_outputs(2313)) or (layer1_outputs(3445));
    layer2_outputs(3864) <= layer1_outputs(828);
    layer2_outputs(3865) <= (layer1_outputs(3594)) or (layer1_outputs(435));
    layer2_outputs(3866) <= (layer1_outputs(2061)) and (layer1_outputs(3381));
    layer2_outputs(3867) <= not(layer1_outputs(4648));
    layer2_outputs(3868) <= (layer1_outputs(3403)) and not (layer1_outputs(3732));
    layer2_outputs(3869) <= not(layer1_outputs(2589)) or (layer1_outputs(1047));
    layer2_outputs(3870) <= '0';
    layer2_outputs(3871) <= (layer1_outputs(697)) and not (layer1_outputs(3809));
    layer2_outputs(3872) <= (layer1_outputs(1048)) and (layer1_outputs(4596));
    layer2_outputs(3873) <= '1';
    layer2_outputs(3874) <= not(layer1_outputs(1));
    layer2_outputs(3875) <= not(layer1_outputs(445)) or (layer1_outputs(4358));
    layer2_outputs(3876) <= not(layer1_outputs(24));
    layer2_outputs(3877) <= layer1_outputs(2262);
    layer2_outputs(3878) <= (layer1_outputs(3678)) and (layer1_outputs(485));
    layer2_outputs(3879) <= (layer1_outputs(4113)) and (layer1_outputs(4765));
    layer2_outputs(3880) <= (layer1_outputs(1784)) and not (layer1_outputs(1254));
    layer2_outputs(3881) <= not((layer1_outputs(444)) and (layer1_outputs(3938)));
    layer2_outputs(3882) <= not(layer1_outputs(4813));
    layer2_outputs(3883) <= layer1_outputs(659);
    layer2_outputs(3884) <= (layer1_outputs(4251)) and (layer1_outputs(1295));
    layer2_outputs(3885) <= (layer1_outputs(2649)) or (layer1_outputs(1849));
    layer2_outputs(3886) <= (layer1_outputs(3723)) and not (layer1_outputs(2938));
    layer2_outputs(3887) <= '1';
    layer2_outputs(3888) <= not(layer1_outputs(4403));
    layer2_outputs(3889) <= '1';
    layer2_outputs(3890) <= not((layer1_outputs(4063)) and (layer1_outputs(2664)));
    layer2_outputs(3891) <= layer1_outputs(4775);
    layer2_outputs(3892) <= (layer1_outputs(307)) and not (layer1_outputs(2867));
    layer2_outputs(3893) <= (layer1_outputs(4220)) or (layer1_outputs(1247));
    layer2_outputs(3894) <= not(layer1_outputs(3380));
    layer2_outputs(3895) <= layer1_outputs(1082);
    layer2_outputs(3896) <= '0';
    layer2_outputs(3897) <= not(layer1_outputs(4544));
    layer2_outputs(3898) <= '1';
    layer2_outputs(3899) <= '1';
    layer2_outputs(3900) <= not(layer1_outputs(1992)) or (layer1_outputs(4395));
    layer2_outputs(3901) <= not((layer1_outputs(640)) and (layer1_outputs(4558)));
    layer2_outputs(3902) <= (layer1_outputs(2566)) or (layer1_outputs(2650));
    layer2_outputs(3903) <= not(layer1_outputs(3106));
    layer2_outputs(3904) <= layer1_outputs(5060);
    layer2_outputs(3905) <= not((layer1_outputs(4600)) or (layer1_outputs(839)));
    layer2_outputs(3906) <= layer1_outputs(2676);
    layer2_outputs(3907) <= (layer1_outputs(3981)) and not (layer1_outputs(71));
    layer2_outputs(3908) <= not(layer1_outputs(4822)) or (layer1_outputs(2894));
    layer2_outputs(3909) <= layer1_outputs(2391);
    layer2_outputs(3910) <= not(layer1_outputs(412)) or (layer1_outputs(3074));
    layer2_outputs(3911) <= not((layer1_outputs(2564)) and (layer1_outputs(692)));
    layer2_outputs(3912) <= not((layer1_outputs(3605)) and (layer1_outputs(4210)));
    layer2_outputs(3913) <= layer1_outputs(1270);
    layer2_outputs(3914) <= not(layer1_outputs(2395));
    layer2_outputs(3915) <= not(layer1_outputs(1959));
    layer2_outputs(3916) <= not(layer1_outputs(4459)) or (layer1_outputs(1689));
    layer2_outputs(3917) <= layer1_outputs(1860);
    layer2_outputs(3918) <= (layer1_outputs(4604)) and (layer1_outputs(1933));
    layer2_outputs(3919) <= (layer1_outputs(2131)) or (layer1_outputs(1517));
    layer2_outputs(3920) <= '0';
    layer2_outputs(3921) <= not((layer1_outputs(3177)) or (layer1_outputs(172)));
    layer2_outputs(3922) <= (layer1_outputs(1341)) and not (layer1_outputs(4763));
    layer2_outputs(3923) <= '1';
    layer2_outputs(3924) <= not(layer1_outputs(3947));
    layer2_outputs(3925) <= (layer1_outputs(4206)) or (layer1_outputs(1513));
    layer2_outputs(3926) <= layer1_outputs(561);
    layer2_outputs(3927) <= '1';
    layer2_outputs(3928) <= not((layer1_outputs(3807)) and (layer1_outputs(3036)));
    layer2_outputs(3929) <= not(layer1_outputs(2193)) or (layer1_outputs(2768));
    layer2_outputs(3930) <= (layer1_outputs(4563)) and not (layer1_outputs(1052));
    layer2_outputs(3931) <= '1';
    layer2_outputs(3932) <= (layer1_outputs(114)) and (layer1_outputs(2266));
    layer2_outputs(3933) <= '1';
    layer2_outputs(3934) <= '0';
    layer2_outputs(3935) <= not((layer1_outputs(4609)) and (layer1_outputs(4442)));
    layer2_outputs(3936) <= '1';
    layer2_outputs(3937) <= (layer1_outputs(483)) or (layer1_outputs(619));
    layer2_outputs(3938) <= not(layer1_outputs(1296)) or (layer1_outputs(3665));
    layer2_outputs(3939) <= not((layer1_outputs(382)) xor (layer1_outputs(2024)));
    layer2_outputs(3940) <= layer1_outputs(3426);
    layer2_outputs(3941) <= not(layer1_outputs(988)) or (layer1_outputs(933));
    layer2_outputs(3942) <= layer1_outputs(563);
    layer2_outputs(3943) <= not(layer1_outputs(887));
    layer2_outputs(3944) <= '0';
    layer2_outputs(3945) <= (layer1_outputs(2893)) and not (layer1_outputs(1713));
    layer2_outputs(3946) <= not((layer1_outputs(1354)) or (layer1_outputs(3799)));
    layer2_outputs(3947) <= '1';
    layer2_outputs(3948) <= layer1_outputs(1910);
    layer2_outputs(3949) <= '1';
    layer2_outputs(3950) <= (layer1_outputs(1619)) and not (layer1_outputs(3354));
    layer2_outputs(3951) <= (layer1_outputs(1592)) and not (layer1_outputs(1966));
    layer2_outputs(3952) <= '1';
    layer2_outputs(3953) <= not((layer1_outputs(1674)) and (layer1_outputs(5119)));
    layer2_outputs(3954) <= not((layer1_outputs(4350)) and (layer1_outputs(1331)));
    layer2_outputs(3955) <= layer1_outputs(2145);
    layer2_outputs(3956) <= '0';
    layer2_outputs(3957) <= not((layer1_outputs(4403)) or (layer1_outputs(4254)));
    layer2_outputs(3958) <= not(layer1_outputs(3472));
    layer2_outputs(3959) <= not((layer1_outputs(3172)) or (layer1_outputs(1523)));
    layer2_outputs(3960) <= layer1_outputs(1325);
    layer2_outputs(3961) <= (layer1_outputs(4629)) and (layer1_outputs(3886));
    layer2_outputs(3962) <= not((layer1_outputs(4893)) or (layer1_outputs(4729)));
    layer2_outputs(3963) <= '0';
    layer2_outputs(3964) <= '0';
    layer2_outputs(3965) <= '0';
    layer2_outputs(3966) <= not(layer1_outputs(183)) or (layer1_outputs(1418));
    layer2_outputs(3967) <= '0';
    layer2_outputs(3968) <= '0';
    layer2_outputs(3969) <= not(layer1_outputs(3221));
    layer2_outputs(3970) <= (layer1_outputs(1825)) and not (layer1_outputs(4647));
    layer2_outputs(3971) <= (layer1_outputs(3410)) and not (layer1_outputs(56));
    layer2_outputs(3972) <= not(layer1_outputs(436)) or (layer1_outputs(3286));
    layer2_outputs(3973) <= not((layer1_outputs(2632)) or (layer1_outputs(280)));
    layer2_outputs(3974) <= not((layer1_outputs(920)) and (layer1_outputs(2797)));
    layer2_outputs(3975) <= not(layer1_outputs(4038)) or (layer1_outputs(862));
    layer2_outputs(3976) <= not(layer1_outputs(4244)) or (layer1_outputs(4226));
    layer2_outputs(3977) <= (layer1_outputs(3495)) or (layer1_outputs(4445));
    layer2_outputs(3978) <= not(layer1_outputs(3544)) or (layer1_outputs(2132));
    layer2_outputs(3979) <= not((layer1_outputs(921)) and (layer1_outputs(2760)));
    layer2_outputs(3980) <= not(layer1_outputs(620)) or (layer1_outputs(1835));
    layer2_outputs(3981) <= (layer1_outputs(1248)) and not (layer1_outputs(1730));
    layer2_outputs(3982) <= (layer1_outputs(1372)) and (layer1_outputs(3443));
    layer2_outputs(3983) <= '1';
    layer2_outputs(3984) <= '0';
    layer2_outputs(3985) <= '0';
    layer2_outputs(3986) <= '1';
    layer2_outputs(3987) <= (layer1_outputs(427)) or (layer1_outputs(3671));
    layer2_outputs(3988) <= not(layer1_outputs(4915));
    layer2_outputs(3989) <= '0';
    layer2_outputs(3990) <= not(layer1_outputs(4586));
    layer2_outputs(3991) <= '1';
    layer2_outputs(3992) <= not(layer1_outputs(587));
    layer2_outputs(3993) <= not((layer1_outputs(4691)) or (layer1_outputs(2578)));
    layer2_outputs(3994) <= layer1_outputs(3595);
    layer2_outputs(3995) <= (layer1_outputs(1015)) and not (layer1_outputs(2782));
    layer2_outputs(3996) <= not(layer1_outputs(4831));
    layer2_outputs(3997) <= (layer1_outputs(3099)) and not (layer1_outputs(2572));
    layer2_outputs(3998) <= (layer1_outputs(3568)) or (layer1_outputs(96));
    layer2_outputs(3999) <= not(layer1_outputs(1229));
    layer2_outputs(4000) <= layer1_outputs(3224);
    layer2_outputs(4001) <= (layer1_outputs(4687)) and not (layer1_outputs(2109));
    layer2_outputs(4002) <= (layer1_outputs(4797)) and not (layer1_outputs(3502));
    layer2_outputs(4003) <= (layer1_outputs(2433)) and not (layer1_outputs(4537));
    layer2_outputs(4004) <= '0';
    layer2_outputs(4005) <= not(layer1_outputs(3848));
    layer2_outputs(4006) <= not((layer1_outputs(206)) and (layer1_outputs(816)));
    layer2_outputs(4007) <= (layer1_outputs(1764)) and not (layer1_outputs(3025));
    layer2_outputs(4008) <= layer1_outputs(3043);
    layer2_outputs(4009) <= '0';
    layer2_outputs(4010) <= not((layer1_outputs(667)) and (layer1_outputs(3039)));
    layer2_outputs(4011) <= not(layer1_outputs(1407)) or (layer1_outputs(5013));
    layer2_outputs(4012) <= '1';
    layer2_outputs(4013) <= not((layer1_outputs(2777)) or (layer1_outputs(4015)));
    layer2_outputs(4014) <= (layer1_outputs(4295)) and (layer1_outputs(209));
    layer2_outputs(4015) <= not(layer1_outputs(4059)) or (layer1_outputs(473));
    layer2_outputs(4016) <= '1';
    layer2_outputs(4017) <= '0';
    layer2_outputs(4018) <= not(layer1_outputs(192));
    layer2_outputs(4019) <= not((layer1_outputs(1294)) and (layer1_outputs(3394)));
    layer2_outputs(4020) <= layer1_outputs(2818);
    layer2_outputs(4021) <= not((layer1_outputs(3812)) and (layer1_outputs(2138)));
    layer2_outputs(4022) <= not(layer1_outputs(1382));
    layer2_outputs(4023) <= not(layer1_outputs(3983)) or (layer1_outputs(1432));
    layer2_outputs(4024) <= layer1_outputs(198);
    layer2_outputs(4025) <= not(layer1_outputs(2679));
    layer2_outputs(4026) <= not(layer1_outputs(4346)) or (layer1_outputs(3993));
    layer2_outputs(4027) <= layer1_outputs(3078);
    layer2_outputs(4028) <= (layer1_outputs(4562)) and not (layer1_outputs(87));
    layer2_outputs(4029) <= (layer1_outputs(3683)) or (layer1_outputs(3485));
    layer2_outputs(4030) <= layer1_outputs(166);
    layer2_outputs(4031) <= not(layer1_outputs(347));
    layer2_outputs(4032) <= layer1_outputs(3010);
    layer2_outputs(4033) <= not((layer1_outputs(3020)) and (layer1_outputs(1715)));
    layer2_outputs(4034) <= (layer1_outputs(4050)) and not (layer1_outputs(4804));
    layer2_outputs(4035) <= not(layer1_outputs(3019));
    layer2_outputs(4036) <= '1';
    layer2_outputs(4037) <= (layer1_outputs(1887)) and not (layer1_outputs(153));
    layer2_outputs(4038) <= (layer1_outputs(4248)) or (layer1_outputs(710));
    layer2_outputs(4039) <= not((layer1_outputs(3139)) or (layer1_outputs(2194)));
    layer2_outputs(4040) <= layer1_outputs(2814);
    layer2_outputs(4041) <= (layer1_outputs(2993)) or (layer1_outputs(3428));
    layer2_outputs(4042) <= not(layer1_outputs(2675));
    layer2_outputs(4043) <= not(layer1_outputs(2084));
    layer2_outputs(4044) <= layer1_outputs(2563);
    layer2_outputs(4045) <= not((layer1_outputs(3528)) and (layer1_outputs(3691)));
    layer2_outputs(4046) <= not(layer1_outputs(3669));
    layer2_outputs(4047) <= not(layer1_outputs(1187)) or (layer1_outputs(1001));
    layer2_outputs(4048) <= not((layer1_outputs(3925)) and (layer1_outputs(900)));
    layer2_outputs(4049) <= '0';
    layer2_outputs(4050) <= not(layer1_outputs(658)) or (layer1_outputs(3401));
    layer2_outputs(4051) <= (layer1_outputs(1370)) or (layer1_outputs(3992));
    layer2_outputs(4052) <= '1';
    layer2_outputs(4053) <= layer1_outputs(1761);
    layer2_outputs(4054) <= not((layer1_outputs(226)) or (layer1_outputs(3480)));
    layer2_outputs(4055) <= '1';
    layer2_outputs(4056) <= (layer1_outputs(3365)) or (layer1_outputs(4018));
    layer2_outputs(4057) <= not(layer1_outputs(4489)) or (layer1_outputs(4741));
    layer2_outputs(4058) <= not(layer1_outputs(3889));
    layer2_outputs(4059) <= not(layer1_outputs(786));
    layer2_outputs(4060) <= (layer1_outputs(4258)) or (layer1_outputs(4725));
    layer2_outputs(4061) <= layer1_outputs(558);
    layer2_outputs(4062) <= not(layer1_outputs(1560)) or (layer1_outputs(294));
    layer2_outputs(4063) <= '0';
    layer2_outputs(4064) <= layer1_outputs(2947);
    layer2_outputs(4065) <= (layer1_outputs(657)) and (layer1_outputs(4286));
    layer2_outputs(4066) <= not(layer1_outputs(3197)) or (layer1_outputs(428));
    layer2_outputs(4067) <= not((layer1_outputs(1489)) or (layer1_outputs(3772)));
    layer2_outputs(4068) <= layer1_outputs(2457);
    layer2_outputs(4069) <= not(layer1_outputs(4315));
    layer2_outputs(4070) <= (layer1_outputs(3241)) and not (layer1_outputs(3586));
    layer2_outputs(4071) <= not(layer1_outputs(1907)) or (layer1_outputs(627));
    layer2_outputs(4072) <= '0';
    layer2_outputs(4073) <= (layer1_outputs(2678)) and (layer1_outputs(3816));
    layer2_outputs(4074) <= not(layer1_outputs(1009));
    layer2_outputs(4075) <= not(layer1_outputs(3311));
    layer2_outputs(4076) <= layer1_outputs(3996);
    layer2_outputs(4077) <= '1';
    layer2_outputs(4078) <= layer1_outputs(1203);
    layer2_outputs(4079) <= '1';
    layer2_outputs(4080) <= not((layer1_outputs(684)) and (layer1_outputs(4575)));
    layer2_outputs(4081) <= not((layer1_outputs(3774)) and (layer1_outputs(4256)));
    layer2_outputs(4082) <= not(layer1_outputs(2072)) or (layer1_outputs(1121));
    layer2_outputs(4083) <= not(layer1_outputs(3479)) or (layer1_outputs(2379));
    layer2_outputs(4084) <= not(layer1_outputs(2972));
    layer2_outputs(4085) <= not(layer1_outputs(861)) or (layer1_outputs(1552));
    layer2_outputs(4086) <= (layer1_outputs(322)) and (layer1_outputs(4986));
    layer2_outputs(4087) <= not((layer1_outputs(3579)) and (layer1_outputs(467)));
    layer2_outputs(4088) <= not((layer1_outputs(5017)) or (layer1_outputs(2143)));
    layer2_outputs(4089) <= not((layer1_outputs(3760)) and (layer1_outputs(1652)));
    layer2_outputs(4090) <= not(layer1_outputs(4649)) or (layer1_outputs(4554));
    layer2_outputs(4091) <= '0';
    layer2_outputs(4092) <= '1';
    layer2_outputs(4093) <= (layer1_outputs(3606)) or (layer1_outputs(2659));
    layer2_outputs(4094) <= layer1_outputs(2728);
    layer2_outputs(4095) <= not(layer1_outputs(1089));
    layer2_outputs(4096) <= '0';
    layer2_outputs(4097) <= not((layer1_outputs(1466)) xor (layer1_outputs(2089)));
    layer2_outputs(4098) <= not((layer1_outputs(3896)) and (layer1_outputs(325)));
    layer2_outputs(4099) <= not(layer1_outputs(4862));
    layer2_outputs(4100) <= (layer1_outputs(1848)) and not (layer1_outputs(463));
    layer2_outputs(4101) <= (layer1_outputs(69)) and not (layer1_outputs(4734));
    layer2_outputs(4102) <= not(layer1_outputs(4730)) or (layer1_outputs(2664));
    layer2_outputs(4103) <= not(layer1_outputs(1994));
    layer2_outputs(4104) <= not(layer1_outputs(3760));
    layer2_outputs(4105) <= not(layer1_outputs(2197));
    layer2_outputs(4106) <= not(layer1_outputs(1168)) or (layer1_outputs(4075));
    layer2_outputs(4107) <= layer1_outputs(2499);
    layer2_outputs(4108) <= layer1_outputs(2744);
    layer2_outputs(4109) <= not(layer1_outputs(4301));
    layer2_outputs(4110) <= not(layer1_outputs(3484));
    layer2_outputs(4111) <= '1';
    layer2_outputs(4112) <= not((layer1_outputs(2723)) or (layer1_outputs(4863)));
    layer2_outputs(4113) <= not(layer1_outputs(1231));
    layer2_outputs(4114) <= not(layer1_outputs(3459)) or (layer1_outputs(4391));
    layer2_outputs(4115) <= (layer1_outputs(4183)) or (layer1_outputs(3934));
    layer2_outputs(4116) <= not(layer1_outputs(32));
    layer2_outputs(4117) <= not(layer1_outputs(4962)) or (layer1_outputs(2490));
    layer2_outputs(4118) <= layer1_outputs(1949);
    layer2_outputs(4119) <= layer1_outputs(1317);
    layer2_outputs(4120) <= not(layer1_outputs(1108));
    layer2_outputs(4121) <= '1';
    layer2_outputs(4122) <= (layer1_outputs(4619)) and not (layer1_outputs(5002));
    layer2_outputs(4123) <= not(layer1_outputs(2363)) or (layer1_outputs(4483));
    layer2_outputs(4124) <= (layer1_outputs(4083)) xor (layer1_outputs(2060));
    layer2_outputs(4125) <= not(layer1_outputs(3575));
    layer2_outputs(4126) <= not((layer1_outputs(2754)) and (layer1_outputs(4755)));
    layer2_outputs(4127) <= (layer1_outputs(149)) and not (layer1_outputs(407));
    layer2_outputs(4128) <= (layer1_outputs(2542)) or (layer1_outputs(709));
    layer2_outputs(4129) <= layer1_outputs(328);
    layer2_outputs(4130) <= not(layer1_outputs(5002));
    layer2_outputs(4131) <= not(layer1_outputs(2212)) or (layer1_outputs(1561));
    layer2_outputs(4132) <= layer1_outputs(4874);
    layer2_outputs(4133) <= (layer1_outputs(3840)) xor (layer1_outputs(359));
    layer2_outputs(4134) <= not(layer1_outputs(1911));
    layer2_outputs(4135) <= layer1_outputs(4130);
    layer2_outputs(4136) <= '1';
    layer2_outputs(4137) <= (layer1_outputs(398)) and not (layer1_outputs(4467));
    layer2_outputs(4138) <= not((layer1_outputs(952)) and (layer1_outputs(1097)));
    layer2_outputs(4139) <= not(layer1_outputs(2254));
    layer2_outputs(4140) <= layer1_outputs(878);
    layer2_outputs(4141) <= '1';
    layer2_outputs(4142) <= (layer1_outputs(5009)) and not (layer1_outputs(5008));
    layer2_outputs(4143) <= (layer1_outputs(4735)) or (layer1_outputs(4390));
    layer2_outputs(4144) <= (layer1_outputs(1181)) and not (layer1_outputs(4660));
    layer2_outputs(4145) <= '0';
    layer2_outputs(4146) <= layer1_outputs(4923);
    layer2_outputs(4147) <= not(layer1_outputs(913)) or (layer1_outputs(3088));
    layer2_outputs(4148) <= not(layer1_outputs(4650)) or (layer1_outputs(716));
    layer2_outputs(4149) <= '1';
    layer2_outputs(4150) <= (layer1_outputs(3533)) or (layer1_outputs(324));
    layer2_outputs(4151) <= layer1_outputs(3817);
    layer2_outputs(4152) <= (layer1_outputs(4654)) and not (layer1_outputs(2860));
    layer2_outputs(4153) <= '0';
    layer2_outputs(4154) <= not(layer1_outputs(2805)) or (layer1_outputs(415));
    layer2_outputs(4155) <= '1';
    layer2_outputs(4156) <= not(layer1_outputs(2579));
    layer2_outputs(4157) <= '0';
    layer2_outputs(4158) <= layer1_outputs(3116);
    layer2_outputs(4159) <= not(layer1_outputs(1157));
    layer2_outputs(4160) <= '0';
    layer2_outputs(4161) <= layer1_outputs(660);
    layer2_outputs(4162) <= not((layer1_outputs(1810)) xor (layer1_outputs(3578)));
    layer2_outputs(4163) <= (layer1_outputs(3246)) or (layer1_outputs(2848));
    layer2_outputs(4164) <= '0';
    layer2_outputs(4165) <= layer1_outputs(1725);
    layer2_outputs(4166) <= not((layer1_outputs(2982)) or (layer1_outputs(1622)));
    layer2_outputs(4167) <= not(layer1_outputs(1506)) or (layer1_outputs(1085));
    layer2_outputs(4168) <= (layer1_outputs(4889)) and (layer1_outputs(2372));
    layer2_outputs(4169) <= not((layer1_outputs(4518)) xor (layer1_outputs(5064)));
    layer2_outputs(4170) <= (layer1_outputs(1319)) or (layer1_outputs(4139));
    layer2_outputs(4171) <= '0';
    layer2_outputs(4172) <= not(layer1_outputs(3800));
    layer2_outputs(4173) <= not((layer1_outputs(4161)) or (layer1_outputs(2839)));
    layer2_outputs(4174) <= '0';
    layer2_outputs(4175) <= (layer1_outputs(3241)) xor (layer1_outputs(298));
    layer2_outputs(4176) <= '1';
    layer2_outputs(4177) <= not(layer1_outputs(4447)) or (layer1_outputs(4766));
    layer2_outputs(4178) <= not((layer1_outputs(3313)) xor (layer1_outputs(2576)));
    layer2_outputs(4179) <= not(layer1_outputs(81));
    layer2_outputs(4180) <= (layer1_outputs(615)) and not (layer1_outputs(4900));
    layer2_outputs(4181) <= not(layer1_outputs(476));
    layer2_outputs(4182) <= '1';
    layer2_outputs(4183) <= '1';
    layer2_outputs(4184) <= not(layer1_outputs(1570)) or (layer1_outputs(2537));
    layer2_outputs(4185) <= (layer1_outputs(2434)) and not (layer1_outputs(3989));
    layer2_outputs(4186) <= '0';
    layer2_outputs(4187) <= '0';
    layer2_outputs(4188) <= not(layer1_outputs(1556)) or (layer1_outputs(189));
    layer2_outputs(4189) <= (layer1_outputs(2464)) and (layer1_outputs(5030));
    layer2_outputs(4190) <= (layer1_outputs(2441)) and not (layer1_outputs(1347));
    layer2_outputs(4191) <= not(layer1_outputs(3667));
    layer2_outputs(4192) <= not(layer1_outputs(1409)) or (layer1_outputs(4295));
    layer2_outputs(4193) <= layer1_outputs(2077);
    layer2_outputs(4194) <= '0';
    layer2_outputs(4195) <= (layer1_outputs(3687)) xor (layer1_outputs(231));
    layer2_outputs(4196) <= layer1_outputs(215);
    layer2_outputs(4197) <= (layer1_outputs(3534)) and (layer1_outputs(489));
    layer2_outputs(4198) <= not(layer1_outputs(2530));
    layer2_outputs(4199) <= not(layer1_outputs(2983));
    layer2_outputs(4200) <= not(layer1_outputs(4356));
    layer2_outputs(4201) <= '1';
    layer2_outputs(4202) <= (layer1_outputs(3342)) and not (layer1_outputs(1847));
    layer2_outputs(4203) <= (layer1_outputs(1718)) or (layer1_outputs(1548));
    layer2_outputs(4204) <= '0';
    layer2_outputs(4205) <= '0';
    layer2_outputs(4206) <= not(layer1_outputs(4013));
    layer2_outputs(4207) <= not((layer1_outputs(505)) xor (layer1_outputs(1920)));
    layer2_outputs(4208) <= '0';
    layer2_outputs(4209) <= not(layer1_outputs(3999));
    layer2_outputs(4210) <= layer1_outputs(3813);
    layer2_outputs(4211) <= not((layer1_outputs(2319)) and (layer1_outputs(1414)));
    layer2_outputs(4212) <= (layer1_outputs(2349)) and not (layer1_outputs(2699));
    layer2_outputs(4213) <= layer1_outputs(4110);
    layer2_outputs(4214) <= not(layer1_outputs(1124)) or (layer1_outputs(1342));
    layer2_outputs(4215) <= (layer1_outputs(4597)) and not (layer1_outputs(761));
    layer2_outputs(4216) <= not(layer1_outputs(3590)) or (layer1_outputs(4734));
    layer2_outputs(4217) <= (layer1_outputs(4208)) and not (layer1_outputs(415));
    layer2_outputs(4218) <= not((layer1_outputs(4243)) and (layer1_outputs(3584)));
    layer2_outputs(4219) <= layer1_outputs(1371);
    layer2_outputs(4220) <= layer1_outputs(3455);
    layer2_outputs(4221) <= layer1_outputs(827);
    layer2_outputs(4222) <= not((layer1_outputs(641)) xor (layer1_outputs(1064)));
    layer2_outputs(4223) <= (layer1_outputs(699)) or (layer1_outputs(2025));
    layer2_outputs(4224) <= layer1_outputs(1044);
    layer2_outputs(4225) <= not(layer1_outputs(1921)) or (layer1_outputs(1511));
    layer2_outputs(4226) <= '0';
    layer2_outputs(4227) <= (layer1_outputs(2147)) or (layer1_outputs(2962));
    layer2_outputs(4228) <= not(layer1_outputs(4947)) or (layer1_outputs(1824));
    layer2_outputs(4229) <= not(layer1_outputs(1993)) or (layer1_outputs(5103));
    layer2_outputs(4230) <= '0';
    layer2_outputs(4231) <= '0';
    layer2_outputs(4232) <= layer1_outputs(2122);
    layer2_outputs(4233) <= (layer1_outputs(849)) or (layer1_outputs(4994));
    layer2_outputs(4234) <= '1';
    layer2_outputs(4235) <= not(layer1_outputs(4420)) or (layer1_outputs(4823));
    layer2_outputs(4236) <= not(layer1_outputs(930)) or (layer1_outputs(2068));
    layer2_outputs(4237) <= (layer1_outputs(4088)) and not (layer1_outputs(2688));
    layer2_outputs(4238) <= not(layer1_outputs(4689)) or (layer1_outputs(2701));
    layer2_outputs(4239) <= not(layer1_outputs(3228));
    layer2_outputs(4240) <= not(layer1_outputs(965));
    layer2_outputs(4241) <= not(layer1_outputs(824));
    layer2_outputs(4242) <= not(layer1_outputs(1461)) or (layer1_outputs(3029));
    layer2_outputs(4243) <= (layer1_outputs(4883)) or (layer1_outputs(4068));
    layer2_outputs(4244) <= not(layer1_outputs(4701)) or (layer1_outputs(2767));
    layer2_outputs(4245) <= (layer1_outputs(4747)) and (layer1_outputs(929));
    layer2_outputs(4246) <= not(layer1_outputs(1099));
    layer2_outputs(4247) <= (layer1_outputs(5112)) or (layer1_outputs(2718));
    layer2_outputs(4248) <= not(layer1_outputs(1789));
    layer2_outputs(4249) <= not(layer1_outputs(1022));
    layer2_outputs(4250) <= not(layer1_outputs(772)) or (layer1_outputs(1342));
    layer2_outputs(4251) <= (layer1_outputs(3689)) or (layer1_outputs(1231));
    layer2_outputs(4252) <= not(layer1_outputs(3607)) or (layer1_outputs(3219));
    layer2_outputs(4253) <= (layer1_outputs(4736)) xor (layer1_outputs(4682));
    layer2_outputs(4254) <= not((layer1_outputs(345)) or (layer1_outputs(3215)));
    layer2_outputs(4255) <= (layer1_outputs(3093)) or (layer1_outputs(3656));
    layer2_outputs(4256) <= (layer1_outputs(3272)) and (layer1_outputs(1079));
    layer2_outputs(4257) <= not(layer1_outputs(1726));
    layer2_outputs(4258) <= layer1_outputs(3042);
    layer2_outputs(4259) <= '0';
    layer2_outputs(4260) <= not(layer1_outputs(3917));
    layer2_outputs(4261) <= (layer1_outputs(4624)) and not (layer1_outputs(2689));
    layer2_outputs(4262) <= layer1_outputs(3516);
    layer2_outputs(4263) <= '1';
    layer2_outputs(4264) <= not(layer1_outputs(289));
    layer2_outputs(4265) <= '0';
    layer2_outputs(4266) <= not(layer1_outputs(2386));
    layer2_outputs(4267) <= not(layer1_outputs(2097));
    layer2_outputs(4268) <= not(layer1_outputs(2514)) or (layer1_outputs(4198));
    layer2_outputs(4269) <= not(layer1_outputs(5));
    layer2_outputs(4270) <= '0';
    layer2_outputs(4271) <= (layer1_outputs(4063)) and not (layer1_outputs(4273));
    layer2_outputs(4272) <= not((layer1_outputs(2296)) and (layer1_outputs(4257)));
    layer2_outputs(4273) <= layer1_outputs(4459);
    layer2_outputs(4274) <= (layer1_outputs(2494)) or (layer1_outputs(1256));
    layer2_outputs(4275) <= not(layer1_outputs(973)) or (layer1_outputs(3540));
    layer2_outputs(4276) <= not(layer1_outputs(3913)) or (layer1_outputs(3624));
    layer2_outputs(4277) <= not(layer1_outputs(3400)) or (layer1_outputs(4392));
    layer2_outputs(4278) <= layer1_outputs(3200);
    layer2_outputs(4279) <= (layer1_outputs(4072)) or (layer1_outputs(582));
    layer2_outputs(4280) <= (layer1_outputs(3383)) and (layer1_outputs(2826));
    layer2_outputs(4281) <= not((layer1_outputs(3767)) and (layer1_outputs(1261)));
    layer2_outputs(4282) <= '0';
    layer2_outputs(4283) <= '0';
    layer2_outputs(4284) <= layer1_outputs(4185);
    layer2_outputs(4285) <= not(layer1_outputs(2130));
    layer2_outputs(4286) <= (layer1_outputs(2917)) and not (layer1_outputs(4556));
    layer2_outputs(4287) <= (layer1_outputs(2128)) and not (layer1_outputs(1828));
    layer2_outputs(4288) <= not(layer1_outputs(2389));
    layer2_outputs(4289) <= not(layer1_outputs(999));
    layer2_outputs(4290) <= not(layer1_outputs(2381));
    layer2_outputs(4291) <= layer1_outputs(4853);
    layer2_outputs(4292) <= not((layer1_outputs(3594)) or (layer1_outputs(1640)));
    layer2_outputs(4293) <= (layer1_outputs(2686)) and not (layer1_outputs(4818));
    layer2_outputs(4294) <= (layer1_outputs(727)) and not (layer1_outputs(2783));
    layer2_outputs(4295) <= not(layer1_outputs(3893));
    layer2_outputs(4296) <= '0';
    layer2_outputs(4297) <= '1';
    layer2_outputs(4298) <= not(layer1_outputs(2780));
    layer2_outputs(4299) <= '1';
    layer2_outputs(4300) <= '0';
    layer2_outputs(4301) <= '0';
    layer2_outputs(4302) <= not(layer1_outputs(3045)) or (layer1_outputs(3486));
    layer2_outputs(4303) <= '0';
    layer2_outputs(4304) <= '1';
    layer2_outputs(4305) <= '0';
    layer2_outputs(4306) <= not((layer1_outputs(1076)) and (layer1_outputs(3011)));
    layer2_outputs(4307) <= (layer1_outputs(1568)) or (layer1_outputs(3258));
    layer2_outputs(4308) <= not(layer1_outputs(4464));
    layer2_outputs(4309) <= not((layer1_outputs(1164)) and (layer1_outputs(3619)));
    layer2_outputs(4310) <= not(layer1_outputs(3026)) or (layer1_outputs(3184));
    layer2_outputs(4311) <= not((layer1_outputs(993)) and (layer1_outputs(3767)));
    layer2_outputs(4312) <= '1';
    layer2_outputs(4313) <= layer1_outputs(889);
    layer2_outputs(4314) <= not(layer1_outputs(1163)) or (layer1_outputs(2443));
    layer2_outputs(4315) <= not(layer1_outputs(4309)) or (layer1_outputs(956));
    layer2_outputs(4316) <= not((layer1_outputs(2831)) or (layer1_outputs(23)));
    layer2_outputs(4317) <= layer1_outputs(966);
    layer2_outputs(4318) <= (layer1_outputs(3616)) and not (layer1_outputs(680));
    layer2_outputs(4319) <= (layer1_outputs(4831)) and not (layer1_outputs(1123));
    layer2_outputs(4320) <= layer1_outputs(454);
    layer2_outputs(4321) <= (layer1_outputs(936)) and (layer1_outputs(3402));
    layer2_outputs(4322) <= (layer1_outputs(1591)) and not (layer1_outputs(4507));
    layer2_outputs(4323) <= not((layer1_outputs(2371)) or (layer1_outputs(3630)));
    layer2_outputs(4324) <= layer1_outputs(1329);
    layer2_outputs(4325) <= (layer1_outputs(2268)) or (layer1_outputs(4230));
    layer2_outputs(4326) <= not(layer1_outputs(4400)) or (layer1_outputs(3193));
    layer2_outputs(4327) <= (layer1_outputs(302)) xor (layer1_outputs(2745));
    layer2_outputs(4328) <= not(layer1_outputs(3407));
    layer2_outputs(4329) <= not(layer1_outputs(850)) or (layer1_outputs(2460));
    layer2_outputs(4330) <= (layer1_outputs(2887)) and not (layer1_outputs(389));
    layer2_outputs(4331) <= (layer1_outputs(3139)) or (layer1_outputs(2712));
    layer2_outputs(4332) <= (layer1_outputs(3130)) or (layer1_outputs(3736));
    layer2_outputs(4333) <= not(layer1_outputs(4454));
    layer2_outputs(4334) <= '1';
    layer2_outputs(4335) <= layer1_outputs(807);
    layer2_outputs(4336) <= (layer1_outputs(4783)) and not (layer1_outputs(3706));
    layer2_outputs(4337) <= (layer1_outputs(1523)) and not (layer1_outputs(2359));
    layer2_outputs(4338) <= '0';
    layer2_outputs(4339) <= '0';
    layer2_outputs(4340) <= not(layer1_outputs(956)) or (layer1_outputs(2337));
    layer2_outputs(4341) <= not(layer1_outputs(960)) or (layer1_outputs(3389));
    layer2_outputs(4342) <= not(layer1_outputs(2486));
    layer2_outputs(4343) <= (layer1_outputs(2238)) and not (layer1_outputs(2812));
    layer2_outputs(4344) <= '1';
    layer2_outputs(4345) <= (layer1_outputs(3050)) xor (layer1_outputs(2180));
    layer2_outputs(4346) <= (layer1_outputs(705)) and not (layer1_outputs(2242));
    layer2_outputs(4347) <= not(layer1_outputs(4198));
    layer2_outputs(4348) <= layer1_outputs(5105);
    layer2_outputs(4349) <= '0';
    layer2_outputs(4350) <= layer1_outputs(2657);
    layer2_outputs(4351) <= layer1_outputs(3727);
    layer2_outputs(4352) <= not(layer1_outputs(2045));
    layer2_outputs(4353) <= '1';
    layer2_outputs(4354) <= (layer1_outputs(600)) and not (layer1_outputs(284));
    layer2_outputs(4355) <= layer1_outputs(2496);
    layer2_outputs(4356) <= '0';
    layer2_outputs(4357) <= '0';
    layer2_outputs(4358) <= (layer1_outputs(2438)) and not (layer1_outputs(2239));
    layer2_outputs(4359) <= '1';
    layer2_outputs(4360) <= layer1_outputs(4213);
    layer2_outputs(4361) <= layer1_outputs(77);
    layer2_outputs(4362) <= '0';
    layer2_outputs(4363) <= not(layer1_outputs(1929));
    layer2_outputs(4364) <= (layer1_outputs(513)) or (layer1_outputs(3555));
    layer2_outputs(4365) <= not(layer1_outputs(1452)) or (layer1_outputs(361));
    layer2_outputs(4366) <= layer1_outputs(287);
    layer2_outputs(4367) <= not((layer1_outputs(3538)) and (layer1_outputs(2000)));
    layer2_outputs(4368) <= not((layer1_outputs(3192)) or (layer1_outputs(4247)));
    layer2_outputs(4369) <= (layer1_outputs(1476)) and not (layer1_outputs(2207));
    layer2_outputs(4370) <= not(layer1_outputs(5085)) or (layer1_outputs(3539));
    layer2_outputs(4371) <= (layer1_outputs(1344)) and not (layer1_outputs(4533));
    layer2_outputs(4372) <= layer1_outputs(622);
    layer2_outputs(4373) <= not(layer1_outputs(2789));
    layer2_outputs(4374) <= layer1_outputs(4412);
    layer2_outputs(4375) <= not((layer1_outputs(593)) and (layer1_outputs(279)));
    layer2_outputs(4376) <= not(layer1_outputs(1600));
    layer2_outputs(4377) <= (layer1_outputs(2636)) and not (layer1_outputs(3271));
    layer2_outputs(4378) <= layer1_outputs(2972);
    layer2_outputs(4379) <= (layer1_outputs(1286)) and (layer1_outputs(2031));
    layer2_outputs(4380) <= '1';
    layer2_outputs(4381) <= not(layer1_outputs(1868)) or (layer1_outputs(29));
    layer2_outputs(4382) <= not(layer1_outputs(4361)) or (layer1_outputs(4796));
    layer2_outputs(4383) <= not((layer1_outputs(3000)) and (layer1_outputs(4216)));
    layer2_outputs(4384) <= not(layer1_outputs(3759));
    layer2_outputs(4385) <= not(layer1_outputs(4526)) or (layer1_outputs(2756));
    layer2_outputs(4386) <= layer1_outputs(235);
    layer2_outputs(4387) <= not(layer1_outputs(4828)) or (layer1_outputs(1292));
    layer2_outputs(4388) <= not(layer1_outputs(1698));
    layer2_outputs(4389) <= (layer1_outputs(1252)) and not (layer1_outputs(1062));
    layer2_outputs(4390) <= not(layer1_outputs(3173)) or (layer1_outputs(1539));
    layer2_outputs(4391) <= '1';
    layer2_outputs(4392) <= (layer1_outputs(4159)) and not (layer1_outputs(4232));
    layer2_outputs(4393) <= not(layer1_outputs(3784)) or (layer1_outputs(3499));
    layer2_outputs(4394) <= '1';
    layer2_outputs(4395) <= not(layer1_outputs(2117));
    layer2_outputs(4396) <= '0';
    layer2_outputs(4397) <= (layer1_outputs(1695)) and not (layer1_outputs(4688));
    layer2_outputs(4398) <= not((layer1_outputs(1639)) or (layer1_outputs(2148)));
    layer2_outputs(4399) <= '1';
    layer2_outputs(4400) <= (layer1_outputs(3959)) and not (layer1_outputs(339));
    layer2_outputs(4401) <= not((layer1_outputs(2119)) or (layer1_outputs(840)));
    layer2_outputs(4402) <= not(layer1_outputs(907)) or (layer1_outputs(474));
    layer2_outputs(4403) <= not((layer1_outputs(3831)) or (layer1_outputs(187)));
    layer2_outputs(4404) <= (layer1_outputs(4452)) or (layer1_outputs(45));
    layer2_outputs(4405) <= not(layer1_outputs(4811)) or (layer1_outputs(3852));
    layer2_outputs(4406) <= '1';
    layer2_outputs(4407) <= layer1_outputs(2599);
    layer2_outputs(4408) <= not(layer1_outputs(2554));
    layer2_outputs(4409) <= (layer1_outputs(5032)) and not (layer1_outputs(4091));
    layer2_outputs(4410) <= (layer1_outputs(4693)) and not (layer1_outputs(1661));
    layer2_outputs(4411) <= (layer1_outputs(683)) and not (layer1_outputs(4060));
    layer2_outputs(4412) <= (layer1_outputs(960)) and not (layer1_outputs(5113));
    layer2_outputs(4413) <= not(layer1_outputs(2674));
    layer2_outputs(4414) <= layer1_outputs(5010);
    layer2_outputs(4415) <= (layer1_outputs(4971)) or (layer1_outputs(2958));
    layer2_outputs(4416) <= (layer1_outputs(3926)) or (layer1_outputs(2610));
    layer2_outputs(4417) <= not(layer1_outputs(4040)) or (layer1_outputs(3981));
    layer2_outputs(4418) <= (layer1_outputs(1060)) or (layer1_outputs(2840));
    layer2_outputs(4419) <= (layer1_outputs(1041)) and not (layer1_outputs(1436));
    layer2_outputs(4420) <= '0';
    layer2_outputs(4421) <= not(layer1_outputs(4539));
    layer2_outputs(4422) <= '1';
    layer2_outputs(4423) <= '1';
    layer2_outputs(4424) <= layer1_outputs(1505);
    layer2_outputs(4425) <= not(layer1_outputs(1435)) or (layer1_outputs(3682));
    layer2_outputs(4426) <= (layer1_outputs(2771)) and not (layer1_outputs(4045));
    layer2_outputs(4427) <= '0';
    layer2_outputs(4428) <= not(layer1_outputs(326));
    layer2_outputs(4429) <= layer1_outputs(454);
    layer2_outputs(4430) <= not((layer1_outputs(5028)) or (layer1_outputs(685)));
    layer2_outputs(4431) <= not((layer1_outputs(5050)) and (layer1_outputs(4667)));
    layer2_outputs(4432) <= '0';
    layer2_outputs(4433) <= '0';
    layer2_outputs(4434) <= not((layer1_outputs(925)) or (layer1_outputs(3503)));
    layer2_outputs(4435) <= (layer1_outputs(3048)) and (layer1_outputs(4972));
    layer2_outputs(4436) <= (layer1_outputs(1686)) or (layer1_outputs(15));
    layer2_outputs(4437) <= not(layer1_outputs(651));
    layer2_outputs(4438) <= (layer1_outputs(4108)) and (layer1_outputs(1497));
    layer2_outputs(4439) <= not(layer1_outputs(3879)) or (layer1_outputs(822));
    layer2_outputs(4440) <= '0';
    layer2_outputs(4441) <= not(layer1_outputs(808)) or (layer1_outputs(53));
    layer2_outputs(4442) <= not((layer1_outputs(2673)) or (layer1_outputs(3332)));
    layer2_outputs(4443) <= layer1_outputs(1151);
    layer2_outputs(4444) <= (layer1_outputs(4621)) and not (layer1_outputs(2107));
    layer2_outputs(4445) <= '1';
    layer2_outputs(4446) <= layer1_outputs(4235);
    layer2_outputs(4447) <= layer1_outputs(629);
    layer2_outputs(4448) <= (layer1_outputs(277)) and (layer1_outputs(4152));
    layer2_outputs(4449) <= '1';
    layer2_outputs(4450) <= (layer1_outputs(3533)) and not (layer1_outputs(1036));
    layer2_outputs(4451) <= layer1_outputs(2580);
    layer2_outputs(4452) <= '0';
    layer2_outputs(4453) <= layer1_outputs(4691);
    layer2_outputs(4454) <= not((layer1_outputs(3746)) and (layer1_outputs(2938)));
    layer2_outputs(4455) <= (layer1_outputs(2387)) or (layer1_outputs(2347));
    layer2_outputs(4456) <= not(layer1_outputs(648));
    layer2_outputs(4457) <= (layer1_outputs(3362)) and not (layer1_outputs(690));
    layer2_outputs(4458) <= not(layer1_outputs(3562)) or (layer1_outputs(926));
    layer2_outputs(4459) <= not(layer1_outputs(83));
    layer2_outputs(4460) <= (layer1_outputs(1067)) and (layer1_outputs(4768));
    layer2_outputs(4461) <= not(layer1_outputs(593));
    layer2_outputs(4462) <= (layer1_outputs(3350)) and not (layer1_outputs(2970));
    layer2_outputs(4463) <= layer1_outputs(694);
    layer2_outputs(4464) <= '0';
    layer2_outputs(4465) <= (layer1_outputs(1963)) and not (layer1_outputs(2559));
    layer2_outputs(4466) <= layer1_outputs(664);
    layer2_outputs(4467) <= '0';
    layer2_outputs(4468) <= layer1_outputs(1628);
    layer2_outputs(4469) <= not(layer1_outputs(331)) or (layer1_outputs(635));
    layer2_outputs(4470) <= '0';
    layer2_outputs(4471) <= not(layer1_outputs(4222));
    layer2_outputs(4472) <= layer1_outputs(3307);
    layer2_outputs(4473) <= (layer1_outputs(5050)) and (layer1_outputs(496));
    layer2_outputs(4474) <= '1';
    layer2_outputs(4475) <= '0';
    layer2_outputs(4476) <= '0';
    layer2_outputs(4477) <= '1';
    layer2_outputs(4478) <= (layer1_outputs(4025)) or (layer1_outputs(3494));
    layer2_outputs(4479) <= layer1_outputs(3109);
    layer2_outputs(4480) <= not(layer1_outputs(3014)) or (layer1_outputs(552));
    layer2_outputs(4481) <= not(layer1_outputs(2050));
    layer2_outputs(4482) <= not(layer1_outputs(4635)) or (layer1_outputs(4668));
    layer2_outputs(4483) <= not(layer1_outputs(3183));
    layer2_outputs(4484) <= (layer1_outputs(1070)) and (layer1_outputs(4934));
    layer2_outputs(4485) <= not(layer1_outputs(1589));
    layer2_outputs(4486) <= not(layer1_outputs(4745));
    layer2_outputs(4487) <= layer1_outputs(4699);
    layer2_outputs(4488) <= '0';
    layer2_outputs(4489) <= (layer1_outputs(4899)) and (layer1_outputs(3070));
    layer2_outputs(4490) <= (layer1_outputs(4740)) and not (layer1_outputs(1209));
    layer2_outputs(4491) <= (layer1_outputs(1927)) and (layer1_outputs(3838));
    layer2_outputs(4492) <= layer1_outputs(2906);
    layer2_outputs(4493) <= not((layer1_outputs(903)) or (layer1_outputs(4952)));
    layer2_outputs(4494) <= not((layer1_outputs(2708)) or (layer1_outputs(2947)));
    layer2_outputs(4495) <= (layer1_outputs(336)) or (layer1_outputs(1246));
    layer2_outputs(4496) <= not(layer1_outputs(668));
    layer2_outputs(4497) <= (layer1_outputs(238)) or (layer1_outputs(3263));
    layer2_outputs(4498) <= not(layer1_outputs(2694));
    layer2_outputs(4499) <= not(layer1_outputs(3880));
    layer2_outputs(4500) <= not(layer1_outputs(3797));
    layer2_outputs(4501) <= (layer1_outputs(2989)) and not (layer1_outputs(2415));
    layer2_outputs(4502) <= layer1_outputs(5097);
    layer2_outputs(4503) <= layer1_outputs(1610);
    layer2_outputs(4504) <= (layer1_outputs(2403)) and not (layer1_outputs(1511));
    layer2_outputs(4505) <= not(layer1_outputs(2456)) or (layer1_outputs(247));
    layer2_outputs(4506) <= (layer1_outputs(1454)) and (layer1_outputs(4961));
    layer2_outputs(4507) <= not(layer1_outputs(731)) or (layer1_outputs(2977));
    layer2_outputs(4508) <= not((layer1_outputs(752)) or (layer1_outputs(4697)));
    layer2_outputs(4509) <= '1';
    layer2_outputs(4510) <= not(layer1_outputs(1724)) or (layer1_outputs(4609));
    layer2_outputs(4511) <= layer1_outputs(1015);
    layer2_outputs(4512) <= not(layer1_outputs(5029)) or (layer1_outputs(175));
    layer2_outputs(4513) <= '0';
    layer2_outputs(4514) <= not(layer1_outputs(2347)) or (layer1_outputs(2840));
    layer2_outputs(4515) <= layer1_outputs(2692);
    layer2_outputs(4516) <= not(layer1_outputs(2478));
    layer2_outputs(4517) <= not(layer1_outputs(348));
    layer2_outputs(4518) <= (layer1_outputs(4869)) or (layer1_outputs(3539));
    layer2_outputs(4519) <= (layer1_outputs(4488)) and not (layer1_outputs(3584));
    layer2_outputs(4520) <= not(layer1_outputs(768)) or (layer1_outputs(754));
    layer2_outputs(4521) <= not(layer1_outputs(401)) or (layer1_outputs(1637));
    layer2_outputs(4522) <= '0';
    layer2_outputs(4523) <= (layer1_outputs(3374)) and (layer1_outputs(2167));
    layer2_outputs(4524) <= layer1_outputs(4707);
    layer2_outputs(4525) <= (layer1_outputs(728)) and not (layer1_outputs(3280));
    layer2_outputs(4526) <= (layer1_outputs(407)) and (layer1_outputs(3103));
    layer2_outputs(4527) <= (layer1_outputs(2994)) and not (layer1_outputs(3007));
    layer2_outputs(4528) <= '1';
    layer2_outputs(4529) <= not(layer1_outputs(282));
    layer2_outputs(4530) <= not(layer1_outputs(837));
    layer2_outputs(4531) <= layer1_outputs(1197);
    layer2_outputs(4532) <= not(layer1_outputs(4433)) or (layer1_outputs(1947));
    layer2_outputs(4533) <= layer1_outputs(1794);
    layer2_outputs(4534) <= not(layer1_outputs(3177)) or (layer1_outputs(1827));
    layer2_outputs(4535) <= layer1_outputs(4119);
    layer2_outputs(4536) <= '1';
    layer2_outputs(4537) <= '1';
    layer2_outputs(4538) <= (layer1_outputs(2300)) and not (layer1_outputs(3804));
    layer2_outputs(4539) <= layer1_outputs(3614);
    layer2_outputs(4540) <= not((layer1_outputs(4585)) and (layer1_outputs(1447)));
    layer2_outputs(4541) <= '1';
    layer2_outputs(4542) <= layer1_outputs(4463);
    layer2_outputs(4543) <= not(layer1_outputs(4773));
    layer2_outputs(4544) <= '1';
    layer2_outputs(4545) <= (layer1_outputs(1544)) or (layer1_outputs(610));
    layer2_outputs(4546) <= not(layer1_outputs(5061));
    layer2_outputs(4547) <= not(layer1_outputs(3864));
    layer2_outputs(4548) <= (layer1_outputs(157)) and not (layer1_outputs(2885));
    layer2_outputs(4549) <= not(layer1_outputs(1385));
    layer2_outputs(4550) <= '1';
    layer2_outputs(4551) <= (layer1_outputs(5062)) and (layer1_outputs(4700));
    layer2_outputs(4552) <= layer1_outputs(363);
    layer2_outputs(4553) <= not(layer1_outputs(1280));
    layer2_outputs(4554) <= (layer1_outputs(1945)) xor (layer1_outputs(747));
    layer2_outputs(4555) <= (layer1_outputs(5032)) and (layer1_outputs(2184));
    layer2_outputs(4556) <= '0';
    layer2_outputs(4557) <= not(layer1_outputs(2580)) or (layer1_outputs(927));
    layer2_outputs(4558) <= '0';
    layer2_outputs(4559) <= '1';
    layer2_outputs(4560) <= not((layer1_outputs(2214)) or (layer1_outputs(2903)));
    layer2_outputs(4561) <= (layer1_outputs(2123)) and not (layer1_outputs(1500));
    layer2_outputs(4562) <= (layer1_outputs(150)) or (layer1_outputs(2111));
    layer2_outputs(4563) <= (layer1_outputs(1561)) and not (layer1_outputs(1896));
    layer2_outputs(4564) <= not((layer1_outputs(2411)) and (layer1_outputs(3537)));
    layer2_outputs(4565) <= layer1_outputs(1122);
    layer2_outputs(4566) <= layer1_outputs(5095);
    layer2_outputs(4567) <= layer1_outputs(2522);
    layer2_outputs(4568) <= (layer1_outputs(2854)) and not (layer1_outputs(3474));
    layer2_outputs(4569) <= (layer1_outputs(4282)) or (layer1_outputs(273));
    layer2_outputs(4570) <= layer1_outputs(2597);
    layer2_outputs(4571) <= (layer1_outputs(2692)) and (layer1_outputs(559));
    layer2_outputs(4572) <= (layer1_outputs(3276)) and not (layer1_outputs(527));
    layer2_outputs(4573) <= not((layer1_outputs(2532)) and (layer1_outputs(3957)));
    layer2_outputs(4574) <= layer1_outputs(3680);
    layer2_outputs(4575) <= '1';
    layer2_outputs(4576) <= '1';
    layer2_outputs(4577) <= not((layer1_outputs(716)) or (layer1_outputs(4481)));
    layer2_outputs(4578) <= layer1_outputs(679);
    layer2_outputs(4579) <= layer1_outputs(5024);
    layer2_outputs(4580) <= not(layer1_outputs(4785));
    layer2_outputs(4581) <= (layer1_outputs(5025)) and not (layer1_outputs(1178));
    layer2_outputs(4582) <= layer1_outputs(2472);
    layer2_outputs(4583) <= '0';
    layer2_outputs(4584) <= '0';
    layer2_outputs(4585) <= not(layer1_outputs(1484)) or (layer1_outputs(2763));
    layer2_outputs(4586) <= (layer1_outputs(375)) and (layer1_outputs(1762));
    layer2_outputs(4587) <= not(layer1_outputs(391));
    layer2_outputs(4588) <= (layer1_outputs(458)) and (layer1_outputs(792));
    layer2_outputs(4589) <= not((layer1_outputs(3268)) or (layer1_outputs(1767)));
    layer2_outputs(4590) <= not((layer1_outputs(4951)) and (layer1_outputs(3628)));
    layer2_outputs(4591) <= not(layer1_outputs(1106));
    layer2_outputs(4592) <= '1';
    layer2_outputs(4593) <= (layer1_outputs(5013)) and (layer1_outputs(4663));
    layer2_outputs(4594) <= layer1_outputs(3546);
    layer2_outputs(4595) <= (layer1_outputs(2321)) and (layer1_outputs(3274));
    layer2_outputs(4596) <= (layer1_outputs(2004)) or (layer1_outputs(605));
    layer2_outputs(4597) <= (layer1_outputs(2581)) and not (layer1_outputs(395));
    layer2_outputs(4598) <= (layer1_outputs(4443)) and not (layer1_outputs(2418));
    layer2_outputs(4599) <= (layer1_outputs(4490)) and not (layer1_outputs(3670));
    layer2_outputs(4600) <= layer1_outputs(3385);
    layer2_outputs(4601) <= (layer1_outputs(3488)) and not (layer1_outputs(350));
    layer2_outputs(4602) <= not(layer1_outputs(2858)) or (layer1_outputs(5040));
    layer2_outputs(4603) <= (layer1_outputs(1393)) and not (layer1_outputs(3007));
    layer2_outputs(4604) <= '1';
    layer2_outputs(4605) <= '1';
    layer2_outputs(4606) <= '1';
    layer2_outputs(4607) <= '0';
    layer2_outputs(4608) <= not(layer1_outputs(4570)) or (layer1_outputs(584));
    layer2_outputs(4609) <= not(layer1_outputs(4495));
    layer2_outputs(4610) <= not(layer1_outputs(3569));
    layer2_outputs(4611) <= '1';
    layer2_outputs(4612) <= not((layer1_outputs(2468)) and (layer1_outputs(221)));
    layer2_outputs(4613) <= not((layer1_outputs(4322)) and (layer1_outputs(1025)));
    layer2_outputs(4614) <= (layer1_outputs(3482)) and not (layer1_outputs(917));
    layer2_outputs(4615) <= '1';
    layer2_outputs(4616) <= not(layer1_outputs(28));
    layer2_outputs(4617) <= '1';
    layer2_outputs(4618) <= not(layer1_outputs(4625));
    layer2_outputs(4619) <= layer1_outputs(2628);
    layer2_outputs(4620) <= layer1_outputs(4603);
    layer2_outputs(4621) <= '1';
    layer2_outputs(4622) <= not(layer1_outputs(2654));
    layer2_outputs(4623) <= not(layer1_outputs(2528));
    layer2_outputs(4624) <= not(layer1_outputs(1173)) or (layer1_outputs(1230));
    layer2_outputs(4625) <= not((layer1_outputs(4325)) and (layer1_outputs(493)));
    layer2_outputs(4626) <= '1';
    layer2_outputs(4627) <= not((layer1_outputs(1055)) or (layer1_outputs(2116)));
    layer2_outputs(4628) <= not((layer1_outputs(4510)) or (layer1_outputs(3548)));
    layer2_outputs(4629) <= '1';
    layer2_outputs(4630) <= not(layer1_outputs(4333));
    layer2_outputs(4631) <= (layer1_outputs(3692)) and not (layer1_outputs(4065));
    layer2_outputs(4632) <= '0';
    layer2_outputs(4633) <= (layer1_outputs(5087)) and not (layer1_outputs(1241));
    layer2_outputs(4634) <= not(layer1_outputs(4399)) or (layer1_outputs(3184));
    layer2_outputs(4635) <= not((layer1_outputs(2152)) and (layer1_outputs(1733)));
    layer2_outputs(4636) <= not((layer1_outputs(93)) and (layer1_outputs(2459)));
    layer2_outputs(4637) <= (layer1_outputs(3563)) and not (layer1_outputs(4896));
    layer2_outputs(4638) <= not((layer1_outputs(2878)) and (layer1_outputs(2450)));
    layer2_outputs(4639) <= not((layer1_outputs(1139)) or (layer1_outputs(1078)));
    layer2_outputs(4640) <= not((layer1_outputs(4626)) or (layer1_outputs(2103)));
    layer2_outputs(4641) <= layer1_outputs(3805);
    layer2_outputs(4642) <= (layer1_outputs(3762)) or (layer1_outputs(4922));
    layer2_outputs(4643) <= not(layer1_outputs(3566)) or (layer1_outputs(675));
    layer2_outputs(4644) <= not(layer1_outputs(2752));
    layer2_outputs(4645) <= layer1_outputs(1886);
    layer2_outputs(4646) <= '1';
    layer2_outputs(4647) <= '0';
    layer2_outputs(4648) <= (layer1_outputs(1723)) and (layer1_outputs(3698));
    layer2_outputs(4649) <= '1';
    layer2_outputs(4650) <= '1';
    layer2_outputs(4651) <= layer1_outputs(2801);
    layer2_outputs(4652) <= not(layer1_outputs(1030));
    layer2_outputs(4653) <= not(layer1_outputs(1811));
    layer2_outputs(4654) <= not(layer1_outputs(2647)) or (layer1_outputs(335));
    layer2_outputs(4655) <= not(layer1_outputs(1300));
    layer2_outputs(4656) <= '0';
    layer2_outputs(4657) <= not((layer1_outputs(5069)) and (layer1_outputs(3435)));
    layer2_outputs(4658) <= not(layer1_outputs(599)) or (layer1_outputs(983));
    layer2_outputs(4659) <= '1';
    layer2_outputs(4660) <= not(layer1_outputs(1193)) or (layer1_outputs(3671));
    layer2_outputs(4661) <= (layer1_outputs(592)) and not (layer1_outputs(3855));
    layer2_outputs(4662) <= not(layer1_outputs(1077));
    layer2_outputs(4663) <= not(layer1_outputs(2125)) or (layer1_outputs(198));
    layer2_outputs(4664) <= not((layer1_outputs(1623)) xor (layer1_outputs(1182)));
    layer2_outputs(4665) <= not(layer1_outputs(2)) or (layer1_outputs(4318));
    layer2_outputs(4666) <= '0';
    layer2_outputs(4667) <= not(layer1_outputs(1806));
    layer2_outputs(4668) <= (layer1_outputs(1471)) and not (layer1_outputs(3105));
    layer2_outputs(4669) <= '1';
    layer2_outputs(4670) <= not(layer1_outputs(4169));
    layer2_outputs(4671) <= not(layer1_outputs(4479));
    layer2_outputs(4672) <= '1';
    layer2_outputs(4673) <= (layer1_outputs(1641)) and not (layer1_outputs(745));
    layer2_outputs(4674) <= layer1_outputs(2100);
    layer2_outputs(4675) <= (layer1_outputs(2678)) or (layer1_outputs(2605));
    layer2_outputs(4676) <= not((layer1_outputs(4623)) or (layer1_outputs(4236)));
    layer2_outputs(4677) <= (layer1_outputs(1619)) and not (layer1_outputs(3833));
    layer2_outputs(4678) <= not(layer1_outputs(4916));
    layer2_outputs(4679) <= '1';
    layer2_outputs(4680) <= not(layer1_outputs(4437));
    layer2_outputs(4681) <= (layer1_outputs(2156)) and (layer1_outputs(1262));
    layer2_outputs(4682) <= not((layer1_outputs(3673)) and (layer1_outputs(3019)));
    layer2_outputs(4683) <= (layer1_outputs(3253)) or (layer1_outputs(137));
    layer2_outputs(4684) <= '0';
    layer2_outputs(4685) <= (layer1_outputs(891)) and not (layer1_outputs(102));
    layer2_outputs(4686) <= layer1_outputs(3640);
    layer2_outputs(4687) <= (layer1_outputs(3791)) and not (layer1_outputs(3320));
    layer2_outputs(4688) <= (layer1_outputs(3791)) and (layer1_outputs(3324));
    layer2_outputs(4689) <= not(layer1_outputs(1606));
    layer2_outputs(4690) <= not(layer1_outputs(3195));
    layer2_outputs(4691) <= (layer1_outputs(3850)) and not (layer1_outputs(3654));
    layer2_outputs(4692) <= not((layer1_outputs(3553)) and (layer1_outputs(1264)));
    layer2_outputs(4693) <= not(layer1_outputs(1113));
    layer2_outputs(4694) <= layer1_outputs(3909);
    layer2_outputs(4695) <= not(layer1_outputs(5049));
    layer2_outputs(4696) <= not((layer1_outputs(2993)) or (layer1_outputs(1823)));
    layer2_outputs(4697) <= (layer1_outputs(740)) or (layer1_outputs(2341));
    layer2_outputs(4698) <= (layer1_outputs(4634)) and (layer1_outputs(164));
    layer2_outputs(4699) <= layer1_outputs(147);
    layer2_outputs(4700) <= not(layer1_outputs(3137));
    layer2_outputs(4701) <= not((layer1_outputs(2528)) or (layer1_outputs(3454)));
    layer2_outputs(4702) <= '0';
    layer2_outputs(4703) <= (layer1_outputs(1660)) and not (layer1_outputs(43));
    layer2_outputs(4704) <= (layer1_outputs(634)) and not (layer1_outputs(1013));
    layer2_outputs(4705) <= (layer1_outputs(1854)) and (layer1_outputs(1744));
    layer2_outputs(4706) <= not((layer1_outputs(3852)) or (layer1_outputs(2759)));
    layer2_outputs(4707) <= not((layer1_outputs(3490)) and (layer1_outputs(1615)));
    layer2_outputs(4708) <= (layer1_outputs(3225)) and not (layer1_outputs(4017));
    layer2_outputs(4709) <= (layer1_outputs(2478)) and not (layer1_outputs(140));
    layer2_outputs(4710) <= (layer1_outputs(3110)) or (layer1_outputs(2447));
    layer2_outputs(4711) <= not((layer1_outputs(4593)) and (layer1_outputs(4983)));
    layer2_outputs(4712) <= (layer1_outputs(3018)) and not (layer1_outputs(3842));
    layer2_outputs(4713) <= (layer1_outputs(4318)) and not (layer1_outputs(557));
    layer2_outputs(4714) <= (layer1_outputs(4109)) and not (layer1_outputs(1627));
    layer2_outputs(4715) <= '0';
    layer2_outputs(4716) <= (layer1_outputs(9)) and not (layer1_outputs(4284));
    layer2_outputs(4717) <= '0';
    layer2_outputs(4718) <= not((layer1_outputs(4636)) and (layer1_outputs(4389)));
    layer2_outputs(4719) <= not(layer1_outputs(5096)) or (layer1_outputs(1020));
    layer2_outputs(4720) <= (layer1_outputs(4499)) and not (layer1_outputs(4103));
    layer2_outputs(4721) <= not((layer1_outputs(881)) xor (layer1_outputs(2485)));
    layer2_outputs(4722) <= not(layer1_outputs(2830));
    layer2_outputs(4723) <= '1';
    layer2_outputs(4724) <= layer1_outputs(3252);
    layer2_outputs(4725) <= not((layer1_outputs(903)) or (layer1_outputs(4241)));
    layer2_outputs(4726) <= not(layer1_outputs(3707));
    layer2_outputs(4727) <= '1';
    layer2_outputs(4728) <= not((layer1_outputs(35)) or (layer1_outputs(4843)));
    layer2_outputs(4729) <= '0';
    layer2_outputs(4730) <= (layer1_outputs(1074)) and (layer1_outputs(1625));
    layer2_outputs(4731) <= '1';
    layer2_outputs(4732) <= not((layer1_outputs(1224)) or (layer1_outputs(3627)));
    layer2_outputs(4733) <= not(layer1_outputs(4213)) or (layer1_outputs(1536));
    layer2_outputs(4734) <= not(layer1_outputs(2600)) or (layer1_outputs(1280));
    layer2_outputs(4735) <= not(layer1_outputs(798));
    layer2_outputs(4736) <= not(layer1_outputs(742)) or (layer1_outputs(959));
    layer2_outputs(4737) <= '1';
    layer2_outputs(4738) <= not((layer1_outputs(4574)) and (layer1_outputs(2094)));
    layer2_outputs(4739) <= (layer1_outputs(1121)) or (layer1_outputs(4401));
    layer2_outputs(4740) <= (layer1_outputs(2129)) and (layer1_outputs(3412));
    layer2_outputs(4741) <= layer1_outputs(4278);
    layer2_outputs(4742) <= '1';
    layer2_outputs(4743) <= not((layer1_outputs(1035)) or (layer1_outputs(2076)));
    layer2_outputs(4744) <= '1';
    layer2_outputs(4745) <= not(layer1_outputs(573));
    layer2_outputs(4746) <= not((layer1_outputs(15)) and (layer1_outputs(4913)));
    layer2_outputs(4747) <= layer1_outputs(4766);
    layer2_outputs(4748) <= (layer1_outputs(1939)) and (layer1_outputs(3694));
    layer2_outputs(4749) <= (layer1_outputs(780)) and (layer1_outputs(1143));
    layer2_outputs(4750) <= '0';
    layer2_outputs(4751) <= not(layer1_outputs(832));
    layer2_outputs(4752) <= layer1_outputs(442);
    layer2_outputs(4753) <= '1';
    layer2_outputs(4754) <= not(layer1_outputs(846));
    layer2_outputs(4755) <= not(layer1_outputs(1018)) or (layer1_outputs(3247));
    layer2_outputs(4756) <= not((layer1_outputs(76)) and (layer1_outputs(3811)));
    layer2_outputs(4757) <= layer1_outputs(4020);
    layer2_outputs(4758) <= layer1_outputs(5078);
    layer2_outputs(4759) <= (layer1_outputs(4054)) xor (layer1_outputs(1838));
    layer2_outputs(4760) <= layer1_outputs(2070);
    layer2_outputs(4761) <= not(layer1_outputs(59));
    layer2_outputs(4762) <= not(layer1_outputs(3094));
    layer2_outputs(4763) <= (layer1_outputs(4129)) and not (layer1_outputs(48));
    layer2_outputs(4764) <= (layer1_outputs(3938)) and not (layer1_outputs(78));
    layer2_outputs(4765) <= (layer1_outputs(1653)) and not (layer1_outputs(1650));
    layer2_outputs(4766) <= not(layer1_outputs(356));
    layer2_outputs(4767) <= layer1_outputs(2605);
    layer2_outputs(4768) <= '0';
    layer2_outputs(4769) <= not(layer1_outputs(2288)) or (layer1_outputs(2939));
    layer2_outputs(4770) <= (layer1_outputs(2482)) and not (layer1_outputs(4217));
    layer2_outputs(4771) <= (layer1_outputs(2953)) and (layer1_outputs(1443));
    layer2_outputs(4772) <= not(layer1_outputs(1634)) or (layer1_outputs(694));
    layer2_outputs(4773) <= not((layer1_outputs(5006)) or (layer1_outputs(3005)));
    layer2_outputs(4774) <= (layer1_outputs(3227)) and not (layer1_outputs(426));
    layer2_outputs(4775) <= not((layer1_outputs(3190)) and (layer1_outputs(2644)));
    layer2_outputs(4776) <= not(layer1_outputs(2463)) or (layer1_outputs(2217));
    layer2_outputs(4777) <= not(layer1_outputs(4359));
    layer2_outputs(4778) <= '1';
    layer2_outputs(4779) <= '1';
    layer2_outputs(4780) <= not(layer1_outputs(3486));
    layer2_outputs(4781) <= not(layer1_outputs(2979));
    layer2_outputs(4782) <= not(layer1_outputs(1472)) or (layer1_outputs(4345));
    layer2_outputs(4783) <= not(layer1_outputs(2933)) or (layer1_outputs(929));
    layer2_outputs(4784) <= layer1_outputs(2596);
    layer2_outputs(4785) <= (layer1_outputs(4820)) and (layer1_outputs(1815));
    layer2_outputs(4786) <= (layer1_outputs(3194)) and not (layer1_outputs(1656));
    layer2_outputs(4787) <= not((layer1_outputs(2041)) and (layer1_outputs(1782)));
    layer2_outputs(4788) <= layer1_outputs(1007);
    layer2_outputs(4789) <= not((layer1_outputs(1878)) and (layer1_outputs(4850)));
    layer2_outputs(4790) <= '0';
    layer2_outputs(4791) <= (layer1_outputs(2474)) or (layer1_outputs(1598));
    layer2_outputs(4792) <= not(layer1_outputs(1023));
    layer2_outputs(4793) <= not(layer1_outputs(4116));
    layer2_outputs(4794) <= '0';
    layer2_outputs(4795) <= (layer1_outputs(1243)) or (layer1_outputs(4836));
    layer2_outputs(4796) <= (layer1_outputs(3597)) and (layer1_outputs(1366));
    layer2_outputs(4797) <= '0';
    layer2_outputs(4798) <= layer1_outputs(431);
    layer2_outputs(4799) <= not(layer1_outputs(3740));
    layer2_outputs(4800) <= (layer1_outputs(4991)) and (layer1_outputs(1722));
    layer2_outputs(4801) <= '0';
    layer2_outputs(4802) <= '1';
    layer2_outputs(4803) <= layer1_outputs(4737);
    layer2_outputs(4804) <= not(layer1_outputs(39)) or (layer1_outputs(3945));
    layer2_outputs(4805) <= '1';
    layer2_outputs(4806) <= not(layer1_outputs(4562)) or (layer1_outputs(711));
    layer2_outputs(4807) <= not(layer1_outputs(4569));
    layer2_outputs(4808) <= (layer1_outputs(54)) and not (layer1_outputs(4226));
    layer2_outputs(4809) <= (layer1_outputs(3205)) and not (layer1_outputs(591));
    layer2_outputs(4810) <= (layer1_outputs(1126)) and not (layer1_outputs(973));
    layer2_outputs(4811) <= (layer1_outputs(4744)) and not (layer1_outputs(2696));
    layer2_outputs(4812) <= layer1_outputs(3275);
    layer2_outputs(4813) <= not(layer1_outputs(1350));
    layer2_outputs(4814) <= not(layer1_outputs(440)) or (layer1_outputs(1351));
    layer2_outputs(4815) <= not(layer1_outputs(108));
    layer2_outputs(4816) <= not(layer1_outputs(1832)) or (layer1_outputs(3822));
    layer2_outputs(4817) <= (layer1_outputs(4814)) and not (layer1_outputs(3202));
    layer2_outputs(4818) <= (layer1_outputs(1778)) or (layer1_outputs(2937));
    layer2_outputs(4819) <= '0';
    layer2_outputs(4820) <= '0';
    layer2_outputs(4821) <= not((layer1_outputs(1908)) and (layer1_outputs(1783)));
    layer2_outputs(4822) <= '1';
    layer2_outputs(4823) <= not(layer1_outputs(3451));
    layer2_outputs(4824) <= layer1_outputs(1787);
    layer2_outputs(4825) <= '1';
    layer2_outputs(4826) <= (layer1_outputs(1095)) and not (layer1_outputs(3795));
    layer2_outputs(4827) <= not(layer1_outputs(2007));
    layer2_outputs(4828) <= layer1_outputs(2773);
    layer2_outputs(4829) <= not(layer1_outputs(4000));
    layer2_outputs(4830) <= (layer1_outputs(4341)) and (layer1_outputs(3323));
    layer2_outputs(4831) <= not((layer1_outputs(3459)) or (layer1_outputs(4010)));
    layer2_outputs(4832) <= not((layer1_outputs(4261)) or (layer1_outputs(146)));
    layer2_outputs(4833) <= '1';
    layer2_outputs(4834) <= (layer1_outputs(2238)) and (layer1_outputs(761));
    layer2_outputs(4835) <= not(layer1_outputs(2667));
    layer2_outputs(4836) <= not(layer1_outputs(4040)) or (layer1_outputs(2767));
    layer2_outputs(4837) <= layer1_outputs(3169);
    layer2_outputs(4838) <= '1';
    layer2_outputs(4839) <= '0';
    layer2_outputs(4840) <= (layer1_outputs(2971)) or (layer1_outputs(317));
    layer2_outputs(4841) <= (layer1_outputs(856)) or (layer1_outputs(3321));
    layer2_outputs(4842) <= '1';
    layer2_outputs(4843) <= not((layer1_outputs(1735)) or (layer1_outputs(3552)));
    layer2_outputs(4844) <= not(layer1_outputs(5101)) or (layer1_outputs(3291));
    layer2_outputs(4845) <= layer1_outputs(4899);
    layer2_outputs(4846) <= not(layer1_outputs(1033));
    layer2_outputs(4847) <= not(layer1_outputs(14));
    layer2_outputs(4848) <= not(layer1_outputs(2273));
    layer2_outputs(4849) <= not(layer1_outputs(1084));
    layer2_outputs(4850) <= layer1_outputs(4666);
    layer2_outputs(4851) <= layer1_outputs(4030);
    layer2_outputs(4852) <= '0';
    layer2_outputs(4853) <= not((layer1_outputs(1977)) and (layer1_outputs(1235)));
    layer2_outputs(4854) <= '1';
    layer2_outputs(4855) <= not((layer1_outputs(488)) and (layer1_outputs(2056)));
    layer2_outputs(4856) <= '0';
    layer2_outputs(4857) <= '0';
    layer2_outputs(4858) <= not(layer1_outputs(3008)) or (layer1_outputs(3364));
    layer2_outputs(4859) <= (layer1_outputs(5100)) and not (layer1_outputs(4127));
    layer2_outputs(4860) <= (layer1_outputs(4438)) and (layer1_outputs(1904));
    layer2_outputs(4861) <= not(layer1_outputs(3505));
    layer2_outputs(4862) <= not((layer1_outputs(3994)) and (layer1_outputs(1585)));
    layer2_outputs(4863) <= not((layer1_outputs(4855)) and (layer1_outputs(4898)));
    layer2_outputs(4864) <= not(layer1_outputs(3066));
    layer2_outputs(4865) <= layer1_outputs(2456);
    layer2_outputs(4866) <= (layer1_outputs(884)) xor (layer1_outputs(4845));
    layer2_outputs(4867) <= not(layer1_outputs(3982)) or (layer1_outputs(3226));
    layer2_outputs(4868) <= (layer1_outputs(2266)) or (layer1_outputs(4812));
    layer2_outputs(4869) <= layer1_outputs(2353);
    layer2_outputs(4870) <= layer1_outputs(4767);
    layer2_outputs(4871) <= '1';
    layer2_outputs(4872) <= not(layer1_outputs(1643));
    layer2_outputs(4873) <= not(layer1_outputs(3217));
    layer2_outputs(4874) <= not((layer1_outputs(3077)) or (layer1_outputs(1027)));
    layer2_outputs(4875) <= not((layer1_outputs(4589)) and (layer1_outputs(4146)));
    layer2_outputs(4876) <= layer1_outputs(618);
    layer2_outputs(4877) <= not(layer1_outputs(62));
    layer2_outputs(4878) <= layer1_outputs(1697);
    layer2_outputs(4879) <= not(layer1_outputs(2593)) or (layer1_outputs(477));
    layer2_outputs(4880) <= not(layer1_outputs(1978)) or (layer1_outputs(1297));
    layer2_outputs(4881) <= '0';
    layer2_outputs(4882) <= not(layer1_outputs(4441));
    layer2_outputs(4883) <= not((layer1_outputs(2783)) and (layer1_outputs(3352)));
    layer2_outputs(4884) <= '0';
    layer2_outputs(4885) <= (layer1_outputs(2423)) and not (layer1_outputs(970));
    layer2_outputs(4886) <= not(layer1_outputs(1363));
    layer2_outputs(4887) <= not(layer1_outputs(1415)) or (layer1_outputs(3745));
    layer2_outputs(4888) <= not((layer1_outputs(1938)) or (layer1_outputs(452)));
    layer2_outputs(4889) <= layer1_outputs(4356);
    layer2_outputs(4890) <= not(layer1_outputs(4023));
    layer2_outputs(4891) <= layer1_outputs(3508);
    layer2_outputs(4892) <= not(layer1_outputs(3703));
    layer2_outputs(4893) <= not(layer1_outputs(2401)) or (layer1_outputs(217));
    layer2_outputs(4894) <= not((layer1_outputs(2415)) xor (layer1_outputs(3526)));
    layer2_outputs(4895) <= not(layer1_outputs(390));
    layer2_outputs(4896) <= not(layer1_outputs(1462)) or (layer1_outputs(3955));
    layer2_outputs(4897) <= not(layer1_outputs(3622));
    layer2_outputs(4898) <= not((layer1_outputs(4343)) or (layer1_outputs(3723)));
    layer2_outputs(4899) <= (layer1_outputs(4800)) and not (layer1_outputs(4578));
    layer2_outputs(4900) <= not(layer1_outputs(3236)) or (layer1_outputs(3941));
    layer2_outputs(4901) <= not(layer1_outputs(1997));
    layer2_outputs(4902) <= '0';
    layer2_outputs(4903) <= layer1_outputs(1528);
    layer2_outputs(4904) <= (layer1_outputs(1234)) or (layer1_outputs(1613));
    layer2_outputs(4905) <= (layer1_outputs(847)) and (layer1_outputs(1658));
    layer2_outputs(4906) <= layer1_outputs(4124);
    layer2_outputs(4907) <= (layer1_outputs(884)) and (layer1_outputs(2875));
    layer2_outputs(4908) <= layer1_outputs(2051);
    layer2_outputs(4909) <= layer1_outputs(2172);
    layer2_outputs(4910) <= not(layer1_outputs(2558));
    layer2_outputs(4911) <= not(layer1_outputs(4924));
    layer2_outputs(4912) <= layer1_outputs(3652);
    layer2_outputs(4913) <= layer1_outputs(1180);
    layer2_outputs(4914) <= (layer1_outputs(686)) and not (layer1_outputs(1439));
    layer2_outputs(4915) <= not(layer1_outputs(1640)) or (layer1_outputs(2755));
    layer2_outputs(4916) <= '1';
    layer2_outputs(4917) <= layer1_outputs(3784);
    layer2_outputs(4918) <= layer1_outputs(4363);
    layer2_outputs(4919) <= not(layer1_outputs(4097));
    layer2_outputs(4920) <= not((layer1_outputs(3684)) or (layer1_outputs(3625)));
    layer2_outputs(4921) <= not(layer1_outputs(1488));
    layer2_outputs(4922) <= (layer1_outputs(1191)) and (layer1_outputs(3003));
    layer2_outputs(4923) <= (layer1_outputs(3366)) or (layer1_outputs(1999));
    layer2_outputs(4924) <= '1';
    layer2_outputs(4925) <= not(layer1_outputs(2691)) or (layer1_outputs(73));
    layer2_outputs(4926) <= (layer1_outputs(2042)) and not (layer1_outputs(1725));
    layer2_outputs(4927) <= not(layer1_outputs(1681)) or (layer1_outputs(2815));
    layer2_outputs(4928) <= not(layer1_outputs(2681));
    layer2_outputs(4929) <= not(layer1_outputs(2240));
    layer2_outputs(4930) <= layer1_outputs(1202);
    layer2_outputs(4931) <= (layer1_outputs(1120)) and not (layer1_outputs(3475));
    layer2_outputs(4932) <= (layer1_outputs(94)) or (layer1_outputs(3102));
    layer2_outputs(4933) <= layer1_outputs(4009);
    layer2_outputs(4934) <= (layer1_outputs(1177)) and (layer1_outputs(4920));
    layer2_outputs(4935) <= layer1_outputs(3768);
    layer2_outputs(4936) <= '1';
    layer2_outputs(4937) <= not(layer1_outputs(3344));
    layer2_outputs(4938) <= not(layer1_outputs(2568));
    layer2_outputs(4939) <= not(layer1_outputs(4720)) or (layer1_outputs(2440));
    layer2_outputs(4940) <= not((layer1_outputs(1682)) and (layer1_outputs(1386)));
    layer2_outputs(4941) <= '0';
    layer2_outputs(4942) <= (layer1_outputs(328)) or (layer1_outputs(394));
    layer2_outputs(4943) <= '0';
    layer2_outputs(4944) <= layer1_outputs(5031);
    layer2_outputs(4945) <= '0';
    layer2_outputs(4946) <= (layer1_outputs(2735)) and (layer1_outputs(3129));
    layer2_outputs(4947) <= (layer1_outputs(4428)) and not (layer1_outputs(1273));
    layer2_outputs(4948) <= '0';
    layer2_outputs(4949) <= not(layer1_outputs(1624));
    layer2_outputs(4950) <= layer1_outputs(1549);
    layer2_outputs(4951) <= not(layer1_outputs(3305));
    layer2_outputs(4952) <= '0';
    layer2_outputs(4953) <= layer1_outputs(2344);
    layer2_outputs(4954) <= not((layer1_outputs(2984)) and (layer1_outputs(4999)));
    layer2_outputs(4955) <= not(layer1_outputs(3912)) or (layer1_outputs(4255));
    layer2_outputs(4956) <= not(layer1_outputs(1632));
    layer2_outputs(4957) <= '0';
    layer2_outputs(4958) <= layer1_outputs(4611);
    layer2_outputs(4959) <= not(layer1_outputs(258));
    layer2_outputs(4960) <= (layer1_outputs(1442)) and not (layer1_outputs(3792));
    layer2_outputs(4961) <= layer1_outputs(3516);
    layer2_outputs(4962) <= (layer1_outputs(4618)) and not (layer1_outputs(1006));
    layer2_outputs(4963) <= layer1_outputs(5046);
    layer2_outputs(4964) <= not((layer1_outputs(979)) and (layer1_outputs(106)));
    layer2_outputs(4965) <= not(layer1_outputs(875)) or (layer1_outputs(4246));
    layer2_outputs(4966) <= '0';
    layer2_outputs(4967) <= (layer1_outputs(1495)) and not (layer1_outputs(2269));
    layer2_outputs(4968) <= not(layer1_outputs(4094));
    layer2_outputs(4969) <= '0';
    layer2_outputs(4970) <= '1';
    layer2_outputs(4971) <= not(layer1_outputs(532)) or (layer1_outputs(3560));
    layer2_outputs(4972) <= layer1_outputs(1759);
    layer2_outputs(4973) <= not(layer1_outputs(2396));
    layer2_outputs(4974) <= '0';
    layer2_outputs(4975) <= '1';
    layer2_outputs(4976) <= not((layer1_outputs(1065)) or (layer1_outputs(1091)));
    layer2_outputs(4977) <= not(layer1_outputs(30)) or (layer1_outputs(4444));
    layer2_outputs(4978) <= (layer1_outputs(2746)) and not (layer1_outputs(3342));
    layer2_outputs(4979) <= not(layer1_outputs(324)) or (layer1_outputs(2748));
    layer2_outputs(4980) <= layer1_outputs(4111);
    layer2_outputs(4981) <= not((layer1_outputs(3692)) and (layer1_outputs(443)));
    layer2_outputs(4982) <= not(layer1_outputs(4765)) or (layer1_outputs(1265));
    layer2_outputs(4983) <= not(layer1_outputs(3520)) or (layer1_outputs(1986));
    layer2_outputs(4984) <= not((layer1_outputs(4352)) and (layer1_outputs(1924)));
    layer2_outputs(4985) <= layer1_outputs(2059);
    layer2_outputs(4986) <= (layer1_outputs(3619)) and (layer1_outputs(2122));
    layer2_outputs(4987) <= not((layer1_outputs(1985)) and (layer1_outputs(631)));
    layer2_outputs(4988) <= not((layer1_outputs(4680)) or (layer1_outputs(3842)));
    layer2_outputs(4989) <= (layer1_outputs(174)) and (layer1_outputs(3860));
    layer2_outputs(4990) <= not((layer1_outputs(7)) xor (layer1_outputs(4645)));
    layer2_outputs(4991) <= not((layer1_outputs(3441)) and (layer1_outputs(4064)));
    layer2_outputs(4992) <= not(layer1_outputs(2114)) or (layer1_outputs(147));
    layer2_outputs(4993) <= layer1_outputs(2845);
    layer2_outputs(4994) <= (layer1_outputs(1958)) and not (layer1_outputs(1405));
    layer2_outputs(4995) <= not(layer1_outputs(1153));
    layer2_outputs(4996) <= not((layer1_outputs(4290)) and (layer1_outputs(3983)));
    layer2_outputs(4997) <= not(layer1_outputs(2870)) or (layer1_outputs(4566));
    layer2_outputs(4998) <= (layer1_outputs(3271)) and not (layer1_outputs(3570));
    layer2_outputs(4999) <= not(layer1_outputs(2325)) or (layer1_outputs(2322));
    layer2_outputs(5000) <= not(layer1_outputs(4230));
    layer2_outputs(5001) <= layer1_outputs(2413);
    layer2_outputs(5002) <= not((layer1_outputs(403)) and (layer1_outputs(594)));
    layer2_outputs(5003) <= (layer1_outputs(1537)) and not (layer1_outputs(4013));
    layer2_outputs(5004) <= (layer1_outputs(2205)) and not (layer1_outputs(3056));
    layer2_outputs(5005) <= '0';
    layer2_outputs(5006) <= (layer1_outputs(4022)) and not (layer1_outputs(2127));
    layer2_outputs(5007) <= not(layer1_outputs(1271));
    layer2_outputs(5008) <= (layer1_outputs(4510)) or (layer1_outputs(1874));
    layer2_outputs(5009) <= (layer1_outputs(4935)) and not (layer1_outputs(14));
    layer2_outputs(5010) <= not(layer1_outputs(3792));
    layer2_outputs(5011) <= not((layer1_outputs(4974)) xor (layer1_outputs(1705)));
    layer2_outputs(5012) <= not((layer1_outputs(4997)) xor (layer1_outputs(4996)));
    layer2_outputs(5013) <= '1';
    layer2_outputs(5014) <= (layer1_outputs(25)) or (layer1_outputs(392));
    layer2_outputs(5015) <= '1';
    layer2_outputs(5016) <= (layer1_outputs(4603)) and not (layer1_outputs(4382));
    layer2_outputs(5017) <= (layer1_outputs(589)) and not (layer1_outputs(1479));
    layer2_outputs(5018) <= layer1_outputs(2111);
    layer2_outputs(5019) <= (layer1_outputs(874)) or (layer1_outputs(2481));
    layer2_outputs(5020) <= (layer1_outputs(3200)) and (layer1_outputs(610));
    layer2_outputs(5021) <= (layer1_outputs(3378)) and (layer1_outputs(724));
    layer2_outputs(5022) <= '0';
    layer2_outputs(5023) <= '0';
    layer2_outputs(5024) <= '0';
    layer2_outputs(5025) <= not(layer1_outputs(655));
    layer2_outputs(5026) <= (layer1_outputs(717)) and not (layer1_outputs(5102));
    layer2_outputs(5027) <= layer1_outputs(4465);
    layer2_outputs(5028) <= layer1_outputs(4637);
    layer2_outputs(5029) <= not(layer1_outputs(1324));
    layer2_outputs(5030) <= not(layer1_outputs(4192));
    layer2_outputs(5031) <= not(layer1_outputs(1344));
    layer2_outputs(5032) <= (layer1_outputs(4511)) and (layer1_outputs(2656));
    layer2_outputs(5033) <= (layer1_outputs(1287)) and (layer1_outputs(984));
    layer2_outputs(5034) <= '1';
    layer2_outputs(5035) <= (layer1_outputs(544)) and not (layer1_outputs(2390));
    layer2_outputs(5036) <= '0';
    layer2_outputs(5037) <= not(layer1_outputs(1564)) or (layer1_outputs(2183));
    layer2_outputs(5038) <= not((layer1_outputs(34)) xor (layer1_outputs(3006)));
    layer2_outputs(5039) <= (layer1_outputs(3182)) and (layer1_outputs(3063));
    layer2_outputs(5040) <= (layer1_outputs(4386)) and not (layer1_outputs(867));
    layer2_outputs(5041) <= not((layer1_outputs(3420)) or (layer1_outputs(469)));
    layer2_outputs(5042) <= layer1_outputs(3030);
    layer2_outputs(5043) <= '0';
    layer2_outputs(5044) <= (layer1_outputs(1085)) and not (layer1_outputs(2756));
    layer2_outputs(5045) <= (layer1_outputs(3726)) and not (layer1_outputs(3496));
    layer2_outputs(5046) <= not(layer1_outputs(201)) or (layer1_outputs(1200));
    layer2_outputs(5047) <= not((layer1_outputs(1221)) or (layer1_outputs(278)));
    layer2_outputs(5048) <= layer1_outputs(2911);
    layer2_outputs(5049) <= not(layer1_outputs(2285)) or (layer1_outputs(2165));
    layer2_outputs(5050) <= not((layer1_outputs(3612)) and (layer1_outputs(2213)));
    layer2_outputs(5051) <= not((layer1_outputs(1819)) and (layer1_outputs(3089)));
    layer2_outputs(5052) <= '0';
    layer2_outputs(5053) <= not(layer1_outputs(122));
    layer2_outputs(5054) <= layer1_outputs(3955);
    layer2_outputs(5055) <= layer1_outputs(2852);
    layer2_outputs(5056) <= (layer1_outputs(4976)) or (layer1_outputs(4125));
    layer2_outputs(5057) <= layer1_outputs(2429);
    layer2_outputs(5058) <= not(layer1_outputs(2179));
    layer2_outputs(5059) <= not((layer1_outputs(2028)) or (layer1_outputs(757)));
    layer2_outputs(5060) <= '1';
    layer2_outputs(5061) <= (layer1_outputs(1753)) and (layer1_outputs(2256));
    layer2_outputs(5062) <= layer1_outputs(36);
    layer2_outputs(5063) <= (layer1_outputs(3049)) and (layer1_outputs(3476));
    layer2_outputs(5064) <= not(layer1_outputs(422)) or (layer1_outputs(3499));
    layer2_outputs(5065) <= '0';
    layer2_outputs(5066) <= (layer1_outputs(1259)) and not (layer1_outputs(5063));
    layer2_outputs(5067) <= (layer1_outputs(1691)) and not (layer1_outputs(4136));
    layer2_outputs(5068) <= not(layer1_outputs(3522)) or (layer1_outputs(2070));
    layer2_outputs(5069) <= not(layer1_outputs(3065)) or (layer1_outputs(181));
    layer2_outputs(5070) <= (layer1_outputs(2892)) and not (layer1_outputs(3024));
    layer2_outputs(5071) <= (layer1_outputs(2645)) and not (layer1_outputs(2975));
    layer2_outputs(5072) <= '1';
    layer2_outputs(5073) <= layer1_outputs(1782);
    layer2_outputs(5074) <= not((layer1_outputs(2150)) or (layer1_outputs(2428)));
    layer2_outputs(5075) <= not(layer1_outputs(4426));
    layer2_outputs(5076) <= not((layer1_outputs(3284)) xor (layer1_outputs(4661)));
    layer2_outputs(5077) <= not((layer1_outputs(4714)) or (layer1_outputs(12)));
    layer2_outputs(5078) <= not(layer1_outputs(4886));
    layer2_outputs(5079) <= layer1_outputs(4731);
    layer2_outputs(5080) <= layer1_outputs(2176);
    layer2_outputs(5081) <= not(layer1_outputs(2493));
    layer2_outputs(5082) <= layer1_outputs(4111);
    layer2_outputs(5083) <= (layer1_outputs(2881)) and not (layer1_outputs(2194));
    layer2_outputs(5084) <= layer1_outputs(4903);
    layer2_outputs(5085) <= '0';
    layer2_outputs(5086) <= layer1_outputs(1279);
    layer2_outputs(5087) <= (layer1_outputs(2150)) and not (layer1_outputs(3743));
    layer2_outputs(5088) <= not(layer1_outputs(4445));
    layer2_outputs(5089) <= '0';
    layer2_outputs(5090) <= (layer1_outputs(1712)) and not (layer1_outputs(3047));
    layer2_outputs(5091) <= not((layer1_outputs(991)) and (layer1_outputs(2118)));
    layer2_outputs(5092) <= (layer1_outputs(1477)) and not (layer1_outputs(2259));
    layer2_outputs(5093) <= not((layer1_outputs(1320)) or (layer1_outputs(2504)));
    layer2_outputs(5094) <= (layer1_outputs(1867)) xor (layer1_outputs(1591));
    layer2_outputs(5095) <= '0';
    layer2_outputs(5096) <= not((layer1_outputs(3677)) or (layer1_outputs(871)));
    layer2_outputs(5097) <= layer1_outputs(24);
    layer2_outputs(5098) <= not(layer1_outputs(3407)) or (layer1_outputs(2969));
    layer2_outputs(5099) <= (layer1_outputs(2195)) and not (layer1_outputs(4560));
    layer2_outputs(5100) <= layer1_outputs(3744);
    layer2_outputs(5101) <= not(layer1_outputs(2491)) or (layer1_outputs(555));
    layer2_outputs(5102) <= not((layer1_outputs(360)) and (layer1_outputs(50)));
    layer2_outputs(5103) <= not(layer1_outputs(4719));
    layer2_outputs(5104) <= not(layer1_outputs(3740));
    layer2_outputs(5105) <= (layer1_outputs(2834)) and (layer1_outputs(3170));
    layer2_outputs(5106) <= not((layer1_outputs(1083)) xor (layer1_outputs(196)));
    layer2_outputs(5107) <= not(layer1_outputs(3880));
    layer2_outputs(5108) <= '0';
    layer2_outputs(5109) <= layer1_outputs(848);
    layer2_outputs(5110) <= layer1_outputs(1275);
    layer2_outputs(5111) <= not((layer1_outputs(2171)) and (layer1_outputs(2411)));
    layer2_outputs(5112) <= not(layer1_outputs(394)) or (layer1_outputs(4922));
    layer2_outputs(5113) <= not(layer1_outputs(2471));
    layer2_outputs(5114) <= '1';
    layer2_outputs(5115) <= layer1_outputs(3081);
    layer2_outputs(5116) <= not(layer1_outputs(384));
    layer2_outputs(5117) <= not((layer1_outputs(1235)) and (layer1_outputs(602)));
    layer2_outputs(5118) <= not(layer1_outputs(3917));
    layer2_outputs(5119) <= layer1_outputs(4376);
    layer3_outputs(0) <= (layer2_outputs(975)) and not (layer2_outputs(1965));
    layer3_outputs(1) <= not(layer2_outputs(2853));
    layer3_outputs(2) <= (layer2_outputs(4198)) and not (layer2_outputs(349));
    layer3_outputs(3) <= '1';
    layer3_outputs(4) <= (layer2_outputs(3546)) or (layer2_outputs(35));
    layer3_outputs(5) <= layer2_outputs(2921);
    layer3_outputs(6) <= (layer2_outputs(2884)) and not (layer2_outputs(4042));
    layer3_outputs(7) <= layer2_outputs(2532);
    layer3_outputs(8) <= '1';
    layer3_outputs(9) <= not(layer2_outputs(2201));
    layer3_outputs(10) <= not(layer2_outputs(1513));
    layer3_outputs(11) <= '0';
    layer3_outputs(12) <= (layer2_outputs(2567)) and not (layer2_outputs(3392));
    layer3_outputs(13) <= not((layer2_outputs(1404)) or (layer2_outputs(1129)));
    layer3_outputs(14) <= not(layer2_outputs(1860)) or (layer2_outputs(3452));
    layer3_outputs(15) <= not(layer2_outputs(4482));
    layer3_outputs(16) <= (layer2_outputs(3925)) or (layer2_outputs(4610));
    layer3_outputs(17) <= not((layer2_outputs(600)) and (layer2_outputs(3332)));
    layer3_outputs(18) <= not(layer2_outputs(112));
    layer3_outputs(19) <= not(layer2_outputs(207));
    layer3_outputs(20) <= not(layer2_outputs(3613));
    layer3_outputs(21) <= '1';
    layer3_outputs(22) <= not(layer2_outputs(2957));
    layer3_outputs(23) <= not(layer2_outputs(4792));
    layer3_outputs(24) <= not(layer2_outputs(4622));
    layer3_outputs(25) <= layer2_outputs(2018);
    layer3_outputs(26) <= '1';
    layer3_outputs(27) <= not((layer2_outputs(2281)) or (layer2_outputs(3420)));
    layer3_outputs(28) <= layer2_outputs(4972);
    layer3_outputs(29) <= not(layer2_outputs(1414)) or (layer2_outputs(2286));
    layer3_outputs(30) <= layer2_outputs(4046);
    layer3_outputs(31) <= (layer2_outputs(1743)) and not (layer2_outputs(463));
    layer3_outputs(32) <= not(layer2_outputs(3938)) or (layer2_outputs(3748));
    layer3_outputs(33) <= not((layer2_outputs(3583)) and (layer2_outputs(999)));
    layer3_outputs(34) <= not(layer2_outputs(1845)) or (layer2_outputs(2150));
    layer3_outputs(35) <= '1';
    layer3_outputs(36) <= (layer2_outputs(1188)) and not (layer2_outputs(4804));
    layer3_outputs(37) <= (layer2_outputs(2528)) or (layer2_outputs(4710));
    layer3_outputs(38) <= layer2_outputs(3052);
    layer3_outputs(39) <= not(layer2_outputs(3903));
    layer3_outputs(40) <= not(layer2_outputs(2867));
    layer3_outputs(41) <= layer2_outputs(1976);
    layer3_outputs(42) <= not((layer2_outputs(1699)) and (layer2_outputs(2638)));
    layer3_outputs(43) <= layer2_outputs(4039);
    layer3_outputs(44) <= not(layer2_outputs(3729));
    layer3_outputs(45) <= (layer2_outputs(2464)) xor (layer2_outputs(3369));
    layer3_outputs(46) <= (layer2_outputs(4122)) and (layer2_outputs(4566));
    layer3_outputs(47) <= not(layer2_outputs(5078)) or (layer2_outputs(3778));
    layer3_outputs(48) <= not(layer2_outputs(14));
    layer3_outputs(49) <= '0';
    layer3_outputs(50) <= '1';
    layer3_outputs(51) <= not((layer2_outputs(1909)) and (layer2_outputs(3199)));
    layer3_outputs(52) <= not(layer2_outputs(2390));
    layer3_outputs(53) <= layer2_outputs(3513);
    layer3_outputs(54) <= layer2_outputs(3251);
    layer3_outputs(55) <= not(layer2_outputs(3252)) or (layer2_outputs(116));
    layer3_outputs(56) <= not((layer2_outputs(3683)) or (layer2_outputs(2174)));
    layer3_outputs(57) <= layer2_outputs(1);
    layer3_outputs(58) <= '1';
    layer3_outputs(59) <= not(layer2_outputs(593));
    layer3_outputs(60) <= '0';
    layer3_outputs(61) <= '1';
    layer3_outputs(62) <= '1';
    layer3_outputs(63) <= not(layer2_outputs(3994));
    layer3_outputs(64) <= layer2_outputs(3966);
    layer3_outputs(65) <= layer2_outputs(4663);
    layer3_outputs(66) <= (layer2_outputs(4766)) and not (layer2_outputs(2998));
    layer3_outputs(67) <= not(layer2_outputs(2652));
    layer3_outputs(68) <= (layer2_outputs(3179)) and (layer2_outputs(3007));
    layer3_outputs(69) <= layer2_outputs(1559);
    layer3_outputs(70) <= layer2_outputs(2152);
    layer3_outputs(71) <= layer2_outputs(4119);
    layer3_outputs(72) <= (layer2_outputs(2501)) and not (layer2_outputs(274));
    layer3_outputs(73) <= not(layer2_outputs(3668));
    layer3_outputs(74) <= not(layer2_outputs(4683));
    layer3_outputs(75) <= not(layer2_outputs(1391)) or (layer2_outputs(2380));
    layer3_outputs(76) <= not((layer2_outputs(687)) and (layer2_outputs(157)));
    layer3_outputs(77) <= not(layer2_outputs(3951));
    layer3_outputs(78) <= not(layer2_outputs(802)) or (layer2_outputs(3644));
    layer3_outputs(79) <= (layer2_outputs(4424)) and not (layer2_outputs(4123));
    layer3_outputs(80) <= layer2_outputs(3722);
    layer3_outputs(81) <= layer2_outputs(1737);
    layer3_outputs(82) <= not(layer2_outputs(1968));
    layer3_outputs(83) <= not((layer2_outputs(3299)) or (layer2_outputs(2164)));
    layer3_outputs(84) <= (layer2_outputs(4777)) and not (layer2_outputs(4355));
    layer3_outputs(85) <= not(layer2_outputs(460));
    layer3_outputs(86) <= layer2_outputs(185);
    layer3_outputs(87) <= not(layer2_outputs(2199));
    layer3_outputs(88) <= layer2_outputs(350);
    layer3_outputs(89) <= layer2_outputs(3554);
    layer3_outputs(90) <= (layer2_outputs(2224)) or (layer2_outputs(2453));
    layer3_outputs(91) <= not(layer2_outputs(421)) or (layer2_outputs(3547));
    layer3_outputs(92) <= not(layer2_outputs(2384)) or (layer2_outputs(4377));
    layer3_outputs(93) <= (layer2_outputs(4846)) and (layer2_outputs(1361));
    layer3_outputs(94) <= (layer2_outputs(2513)) and not (layer2_outputs(3065));
    layer3_outputs(95) <= not(layer2_outputs(796)) or (layer2_outputs(2806));
    layer3_outputs(96) <= '0';
    layer3_outputs(97) <= (layer2_outputs(1745)) and not (layer2_outputs(2079));
    layer3_outputs(98) <= not((layer2_outputs(4586)) and (layer2_outputs(2178)));
    layer3_outputs(99) <= not(layer2_outputs(2473));
    layer3_outputs(100) <= (layer2_outputs(4455)) and not (layer2_outputs(2280));
    layer3_outputs(101) <= not(layer2_outputs(4500));
    layer3_outputs(102) <= not((layer2_outputs(1081)) or (layer2_outputs(3208)));
    layer3_outputs(103) <= '1';
    layer3_outputs(104) <= not(layer2_outputs(1197));
    layer3_outputs(105) <= not(layer2_outputs(5014));
    layer3_outputs(106) <= layer2_outputs(1462);
    layer3_outputs(107) <= not(layer2_outputs(1159)) or (layer2_outputs(1563));
    layer3_outputs(108) <= '1';
    layer3_outputs(109) <= '1';
    layer3_outputs(110) <= not((layer2_outputs(4657)) xor (layer2_outputs(493)));
    layer3_outputs(111) <= not((layer2_outputs(3765)) and (layer2_outputs(3051)));
    layer3_outputs(112) <= not(layer2_outputs(230));
    layer3_outputs(113) <= layer2_outputs(1956);
    layer3_outputs(114) <= layer2_outputs(4193);
    layer3_outputs(115) <= '1';
    layer3_outputs(116) <= (layer2_outputs(4282)) and (layer2_outputs(4617));
    layer3_outputs(117) <= not((layer2_outputs(124)) or (layer2_outputs(1273)));
    layer3_outputs(118) <= layer2_outputs(3975);
    layer3_outputs(119) <= (layer2_outputs(4139)) or (layer2_outputs(3734));
    layer3_outputs(120) <= not((layer2_outputs(3191)) xor (layer2_outputs(4128)));
    layer3_outputs(121) <= '1';
    layer3_outputs(122) <= (layer2_outputs(1758)) or (layer2_outputs(2303));
    layer3_outputs(123) <= not(layer2_outputs(560));
    layer3_outputs(124) <= '0';
    layer3_outputs(125) <= not(layer2_outputs(697));
    layer3_outputs(126) <= (layer2_outputs(74)) and not (layer2_outputs(3853));
    layer3_outputs(127) <= not((layer2_outputs(3539)) and (layer2_outputs(2848)));
    layer3_outputs(128) <= layer2_outputs(2230);
    layer3_outputs(129) <= not(layer2_outputs(3996));
    layer3_outputs(130) <= '0';
    layer3_outputs(131) <= (layer2_outputs(351)) and not (layer2_outputs(611));
    layer3_outputs(132) <= not(layer2_outputs(571));
    layer3_outputs(133) <= (layer2_outputs(1124)) and not (layer2_outputs(3163));
    layer3_outputs(134) <= layer2_outputs(1071);
    layer3_outputs(135) <= not(layer2_outputs(3154)) or (layer2_outputs(2846));
    layer3_outputs(136) <= not((layer2_outputs(4491)) xor (layer2_outputs(877)));
    layer3_outputs(137) <= layer2_outputs(57);
    layer3_outputs(138) <= (layer2_outputs(3102)) or (layer2_outputs(4038));
    layer3_outputs(139) <= not(layer2_outputs(4514)) or (layer2_outputs(541));
    layer3_outputs(140) <= '0';
    layer3_outputs(141) <= layer2_outputs(2802);
    layer3_outputs(142) <= (layer2_outputs(4906)) and not (layer2_outputs(626));
    layer3_outputs(143) <= not((layer2_outputs(3601)) and (layer2_outputs(4444)));
    layer3_outputs(144) <= not((layer2_outputs(3539)) or (layer2_outputs(911)));
    layer3_outputs(145) <= not((layer2_outputs(4844)) or (layer2_outputs(2020)));
    layer3_outputs(146) <= not((layer2_outputs(2866)) and (layer2_outputs(3711)));
    layer3_outputs(147) <= (layer2_outputs(1429)) and not (layer2_outputs(3383));
    layer3_outputs(148) <= not((layer2_outputs(4338)) and (layer2_outputs(672)));
    layer3_outputs(149) <= not((layer2_outputs(3742)) or (layer2_outputs(4505)));
    layer3_outputs(150) <= not(layer2_outputs(4879));
    layer3_outputs(151) <= not((layer2_outputs(4056)) and (layer2_outputs(712)));
    layer3_outputs(152) <= not(layer2_outputs(3046));
    layer3_outputs(153) <= not((layer2_outputs(1614)) xor (layer2_outputs(877)));
    layer3_outputs(154) <= not((layer2_outputs(1232)) or (layer2_outputs(1275)));
    layer3_outputs(155) <= not(layer2_outputs(2575)) or (layer2_outputs(133));
    layer3_outputs(156) <= not(layer2_outputs(2891)) or (layer2_outputs(2408));
    layer3_outputs(157) <= layer2_outputs(3576);
    layer3_outputs(158) <= (layer2_outputs(436)) and not (layer2_outputs(1516));
    layer3_outputs(159) <= layer2_outputs(4695);
    layer3_outputs(160) <= '0';
    layer3_outputs(161) <= not((layer2_outputs(3766)) or (layer2_outputs(3472)));
    layer3_outputs(162) <= not((layer2_outputs(1988)) or (layer2_outputs(3608)));
    layer3_outputs(163) <= (layer2_outputs(4927)) or (layer2_outputs(2138));
    layer3_outputs(164) <= not(layer2_outputs(570)) or (layer2_outputs(2816));
    layer3_outputs(165) <= (layer2_outputs(742)) or (layer2_outputs(1989));
    layer3_outputs(166) <= not(layer2_outputs(3153)) or (layer2_outputs(2160));
    layer3_outputs(167) <= not(layer2_outputs(3867));
    layer3_outputs(168) <= not(layer2_outputs(5045)) or (layer2_outputs(671));
    layer3_outputs(169) <= '0';
    layer3_outputs(170) <= (layer2_outputs(1398)) or (layer2_outputs(1524));
    layer3_outputs(171) <= (layer2_outputs(4091)) and (layer2_outputs(4595));
    layer3_outputs(172) <= layer2_outputs(3353);
    layer3_outputs(173) <= (layer2_outputs(4412)) and not (layer2_outputs(4751));
    layer3_outputs(174) <= (layer2_outputs(656)) and (layer2_outputs(2681));
    layer3_outputs(175) <= (layer2_outputs(4041)) or (layer2_outputs(4342));
    layer3_outputs(176) <= not(layer2_outputs(3243));
    layer3_outputs(177) <= '0';
    layer3_outputs(178) <= (layer2_outputs(2958)) and (layer2_outputs(3271));
    layer3_outputs(179) <= (layer2_outputs(3817)) and (layer2_outputs(648));
    layer3_outputs(180) <= (layer2_outputs(866)) or (layer2_outputs(905));
    layer3_outputs(181) <= (layer2_outputs(1302)) or (layer2_outputs(2352));
    layer3_outputs(182) <= layer2_outputs(3196);
    layer3_outputs(183) <= (layer2_outputs(182)) and not (layer2_outputs(231));
    layer3_outputs(184) <= layer2_outputs(3936);
    layer3_outputs(185) <= not(layer2_outputs(1614)) or (layer2_outputs(4286));
    layer3_outputs(186) <= not(layer2_outputs(2015));
    layer3_outputs(187) <= not(layer2_outputs(475));
    layer3_outputs(188) <= layer2_outputs(2306);
    layer3_outputs(189) <= (layer2_outputs(3146)) or (layer2_outputs(3072));
    layer3_outputs(190) <= not(layer2_outputs(2591)) or (layer2_outputs(4085));
    layer3_outputs(191) <= (layer2_outputs(3124)) or (layer2_outputs(2915));
    layer3_outputs(192) <= not(layer2_outputs(4978));
    layer3_outputs(193) <= layer2_outputs(4973);
    layer3_outputs(194) <= layer2_outputs(1076);
    layer3_outputs(195) <= layer2_outputs(791);
    layer3_outputs(196) <= not(layer2_outputs(4302)) or (layer2_outputs(129));
    layer3_outputs(197) <= (layer2_outputs(3995)) or (layer2_outputs(4446));
    layer3_outputs(198) <= (layer2_outputs(4006)) and not (layer2_outputs(3923));
    layer3_outputs(199) <= not(layer2_outputs(859));
    layer3_outputs(200) <= not((layer2_outputs(1192)) or (layer2_outputs(1798)));
    layer3_outputs(201) <= not(layer2_outputs(1984));
    layer3_outputs(202) <= (layer2_outputs(3879)) and not (layer2_outputs(4559));
    layer3_outputs(203) <= layer2_outputs(2866);
    layer3_outputs(204) <= layer2_outputs(949);
    layer3_outputs(205) <= (layer2_outputs(4623)) and not (layer2_outputs(1578));
    layer3_outputs(206) <= (layer2_outputs(302)) and not (layer2_outputs(3664));
    layer3_outputs(207) <= not((layer2_outputs(4904)) or (layer2_outputs(2187)));
    layer3_outputs(208) <= not(layer2_outputs(3365));
    layer3_outputs(209) <= (layer2_outputs(4237)) and not (layer2_outputs(2002));
    layer3_outputs(210) <= (layer2_outputs(2220)) or (layer2_outputs(5003));
    layer3_outputs(211) <= (layer2_outputs(3672)) and not (layer2_outputs(971));
    layer3_outputs(212) <= not(layer2_outputs(2303));
    layer3_outputs(213) <= '1';
    layer3_outputs(214) <= layer2_outputs(3848);
    layer3_outputs(215) <= not((layer2_outputs(1388)) and (layer2_outputs(672)));
    layer3_outputs(216) <= layer2_outputs(1666);
    layer3_outputs(217) <= not(layer2_outputs(235)) or (layer2_outputs(2629));
    layer3_outputs(218) <= not((layer2_outputs(1520)) or (layer2_outputs(1604)));
    layer3_outputs(219) <= layer2_outputs(2538);
    layer3_outputs(220) <= not(layer2_outputs(4827)) or (layer2_outputs(4975));
    layer3_outputs(221) <= not((layer2_outputs(986)) and (layer2_outputs(3984)));
    layer3_outputs(222) <= not((layer2_outputs(2273)) and (layer2_outputs(2549)));
    layer3_outputs(223) <= not(layer2_outputs(629));
    layer3_outputs(224) <= not(layer2_outputs(1601));
    layer3_outputs(225) <= not((layer2_outputs(3626)) or (layer2_outputs(3674)));
    layer3_outputs(226) <= (layer2_outputs(1702)) or (layer2_outputs(4083));
    layer3_outputs(227) <= (layer2_outputs(4530)) xor (layer2_outputs(2759));
    layer3_outputs(228) <= layer2_outputs(4847);
    layer3_outputs(229) <= layer2_outputs(4192);
    layer3_outputs(230) <= not(layer2_outputs(597));
    layer3_outputs(231) <= not(layer2_outputs(1719));
    layer3_outputs(232) <= not(layer2_outputs(2941));
    layer3_outputs(233) <= layer2_outputs(4788);
    layer3_outputs(234) <= (layer2_outputs(4405)) or (layer2_outputs(2399));
    layer3_outputs(235) <= layer2_outputs(973);
    layer3_outputs(236) <= '1';
    layer3_outputs(237) <= not((layer2_outputs(3174)) or (layer2_outputs(3045)));
    layer3_outputs(238) <= not((layer2_outputs(511)) or (layer2_outputs(1492)));
    layer3_outputs(239) <= '0';
    layer3_outputs(240) <= layer2_outputs(3041);
    layer3_outputs(241) <= (layer2_outputs(636)) or (layer2_outputs(4732));
    layer3_outputs(242) <= layer2_outputs(1101);
    layer3_outputs(243) <= not(layer2_outputs(790));
    layer3_outputs(244) <= not(layer2_outputs(4492));
    layer3_outputs(245) <= layer2_outputs(2525);
    layer3_outputs(246) <= not((layer2_outputs(1516)) or (layer2_outputs(4704)));
    layer3_outputs(247) <= (layer2_outputs(2987)) and not (layer2_outputs(627));
    layer3_outputs(248) <= '0';
    layer3_outputs(249) <= not((layer2_outputs(4072)) and (layer2_outputs(2652)));
    layer3_outputs(250) <= (layer2_outputs(3465)) and not (layer2_outputs(4493));
    layer3_outputs(251) <= layer2_outputs(2405);
    layer3_outputs(252) <= not(layer2_outputs(171)) or (layer2_outputs(3791));
    layer3_outputs(253) <= layer2_outputs(1553);
    layer3_outputs(254) <= (layer2_outputs(3991)) or (layer2_outputs(1971));
    layer3_outputs(255) <= layer2_outputs(2918);
    layer3_outputs(256) <= not(layer2_outputs(550));
    layer3_outputs(257) <= not(layer2_outputs(3291));
    layer3_outputs(258) <= not(layer2_outputs(5083));
    layer3_outputs(259) <= layer2_outputs(3368);
    layer3_outputs(260) <= '1';
    layer3_outputs(261) <= not(layer2_outputs(2421)) or (layer2_outputs(33));
    layer3_outputs(262) <= not(layer2_outputs(2740));
    layer3_outputs(263) <= not(layer2_outputs(3023));
    layer3_outputs(264) <= '0';
    layer3_outputs(265) <= (layer2_outputs(4773)) and (layer2_outputs(3000));
    layer3_outputs(266) <= (layer2_outputs(4129)) or (layer2_outputs(1870));
    layer3_outputs(267) <= '1';
    layer3_outputs(268) <= layer2_outputs(732);
    layer3_outputs(269) <= not(layer2_outputs(373));
    layer3_outputs(270) <= not((layer2_outputs(2727)) or (layer2_outputs(1378)));
    layer3_outputs(271) <= not(layer2_outputs(3203));
    layer3_outputs(272) <= (layer2_outputs(2155)) or (layer2_outputs(247));
    layer3_outputs(273) <= '1';
    layer3_outputs(274) <= layer2_outputs(2007);
    layer3_outputs(275) <= layer2_outputs(2238);
    layer3_outputs(276) <= '1';
    layer3_outputs(277) <= not(layer2_outputs(3151)) or (layer2_outputs(1140));
    layer3_outputs(278) <= layer2_outputs(2527);
    layer3_outputs(279) <= layer2_outputs(2076);
    layer3_outputs(280) <= (layer2_outputs(1571)) and not (layer2_outputs(3753));
    layer3_outputs(281) <= (layer2_outputs(2420)) and not (layer2_outputs(472));
    layer3_outputs(282) <= not(layer2_outputs(3090));
    layer3_outputs(283) <= (layer2_outputs(2577)) or (layer2_outputs(987));
    layer3_outputs(284) <= (layer2_outputs(5054)) or (layer2_outputs(1041));
    layer3_outputs(285) <= not((layer2_outputs(2025)) and (layer2_outputs(71)));
    layer3_outputs(286) <= not((layer2_outputs(1268)) and (layer2_outputs(175)));
    layer3_outputs(287) <= layer2_outputs(812);
    layer3_outputs(288) <= (layer2_outputs(470)) or (layer2_outputs(3750));
    layer3_outputs(289) <= (layer2_outputs(4921)) and not (layer2_outputs(3106));
    layer3_outputs(290) <= not(layer2_outputs(3596)) or (layer2_outputs(870));
    layer3_outputs(291) <= '0';
    layer3_outputs(292) <= not((layer2_outputs(267)) or (layer2_outputs(3092)));
    layer3_outputs(293) <= (layer2_outputs(921)) and not (layer2_outputs(1731));
    layer3_outputs(294) <= (layer2_outputs(3782)) and (layer2_outputs(4852));
    layer3_outputs(295) <= not(layer2_outputs(2593));
    layer3_outputs(296) <= not((layer2_outputs(3518)) or (layer2_outputs(2220)));
    layer3_outputs(297) <= not(layer2_outputs(3119));
    layer3_outputs(298) <= not((layer2_outputs(4834)) or (layer2_outputs(1254)));
    layer3_outputs(299) <= '0';
    layer3_outputs(300) <= layer2_outputs(3782);
    layer3_outputs(301) <= not((layer2_outputs(4772)) and (layer2_outputs(808)));
    layer3_outputs(302) <= '0';
    layer3_outputs(303) <= (layer2_outputs(3977)) and not (layer2_outputs(1459));
    layer3_outputs(304) <= not(layer2_outputs(2257));
    layer3_outputs(305) <= not(layer2_outputs(4762)) or (layer2_outputs(1762));
    layer3_outputs(306) <= '1';
    layer3_outputs(307) <= (layer2_outputs(2222)) or (layer2_outputs(3235));
    layer3_outputs(308) <= (layer2_outputs(1149)) and not (layer2_outputs(4864));
    layer3_outputs(309) <= not(layer2_outputs(2893)) or (layer2_outputs(3278));
    layer3_outputs(310) <= layer2_outputs(1101);
    layer3_outputs(311) <= (layer2_outputs(1693)) and not (layer2_outputs(4719));
    layer3_outputs(312) <= layer2_outputs(629);
    layer3_outputs(313) <= (layer2_outputs(1653)) and (layer2_outputs(2484));
    layer3_outputs(314) <= not(layer2_outputs(4946));
    layer3_outputs(315) <= (layer2_outputs(996)) and (layer2_outputs(648));
    layer3_outputs(316) <= layer2_outputs(3736);
    layer3_outputs(317) <= not(layer2_outputs(1083)) or (layer2_outputs(75));
    layer3_outputs(318) <= layer2_outputs(1262);
    layer3_outputs(319) <= not((layer2_outputs(4604)) and (layer2_outputs(4360)));
    layer3_outputs(320) <= '0';
    layer3_outputs(321) <= layer2_outputs(2200);
    layer3_outputs(322) <= not((layer2_outputs(79)) and (layer2_outputs(108)));
    layer3_outputs(323) <= (layer2_outputs(2714)) and (layer2_outputs(3087));
    layer3_outputs(324) <= not((layer2_outputs(4798)) and (layer2_outputs(4612)));
    layer3_outputs(325) <= (layer2_outputs(517)) and (layer2_outputs(3864));
    layer3_outputs(326) <= layer2_outputs(3617);
    layer3_outputs(327) <= not(layer2_outputs(2130)) or (layer2_outputs(3598));
    layer3_outputs(328) <= not((layer2_outputs(2939)) and (layer2_outputs(1647)));
    layer3_outputs(329) <= not((layer2_outputs(195)) and (layer2_outputs(2043)));
    layer3_outputs(330) <= not(layer2_outputs(2252)) or (layer2_outputs(3245));
    layer3_outputs(331) <= layer2_outputs(5039);
    layer3_outputs(332) <= (layer2_outputs(4991)) and not (layer2_outputs(73));
    layer3_outputs(333) <= layer2_outputs(4793);
    layer3_outputs(334) <= (layer2_outputs(3433)) and not (layer2_outputs(960));
    layer3_outputs(335) <= (layer2_outputs(3359)) and not (layer2_outputs(4997));
    layer3_outputs(336) <= (layer2_outputs(911)) or (layer2_outputs(2005));
    layer3_outputs(337) <= not(layer2_outputs(2));
    layer3_outputs(338) <= (layer2_outputs(4112)) or (layer2_outputs(1118));
    layer3_outputs(339) <= not(layer2_outputs(2114));
    layer3_outputs(340) <= (layer2_outputs(4307)) or (layer2_outputs(2624));
    layer3_outputs(341) <= (layer2_outputs(137)) and (layer2_outputs(5033));
    layer3_outputs(342) <= '0';
    layer3_outputs(343) <= not(layer2_outputs(1729)) or (layer2_outputs(1259));
    layer3_outputs(344) <= not((layer2_outputs(3138)) or (layer2_outputs(3964)));
    layer3_outputs(345) <= (layer2_outputs(156)) and not (layer2_outputs(1803));
    layer3_outputs(346) <= (layer2_outputs(2118)) and not (layer2_outputs(1890));
    layer3_outputs(347) <= layer2_outputs(1866);
    layer3_outputs(348) <= not(layer2_outputs(1957));
    layer3_outputs(349) <= (layer2_outputs(4968)) and (layer2_outputs(938));
    layer3_outputs(350) <= not(layer2_outputs(3416));
    layer3_outputs(351) <= (layer2_outputs(405)) or (layer2_outputs(3612));
    layer3_outputs(352) <= (layer2_outputs(2142)) and (layer2_outputs(4697));
    layer3_outputs(353) <= '1';
    layer3_outputs(354) <= not((layer2_outputs(1479)) or (layer2_outputs(1326)));
    layer3_outputs(355) <= '1';
    layer3_outputs(356) <= layer2_outputs(2179);
    layer3_outputs(357) <= (layer2_outputs(2103)) xor (layer2_outputs(4905));
    layer3_outputs(358) <= (layer2_outputs(3431)) and not (layer2_outputs(3250));
    layer3_outputs(359) <= not(layer2_outputs(2835));
    layer3_outputs(360) <= (layer2_outputs(997)) xor (layer2_outputs(4556));
    layer3_outputs(361) <= not((layer2_outputs(126)) or (layer2_outputs(2115)));
    layer3_outputs(362) <= not(layer2_outputs(3677)) or (layer2_outputs(4550));
    layer3_outputs(363) <= not((layer2_outputs(3474)) and (layer2_outputs(4705)));
    layer3_outputs(364) <= not(layer2_outputs(1921));
    layer3_outputs(365) <= '0';
    layer3_outputs(366) <= not((layer2_outputs(351)) and (layer2_outputs(4479)));
    layer3_outputs(367) <= not(layer2_outputs(1301));
    layer3_outputs(368) <= (layer2_outputs(4811)) and not (layer2_outputs(902));
    layer3_outputs(369) <= not((layer2_outputs(1343)) and (layer2_outputs(2714)));
    layer3_outputs(370) <= (layer2_outputs(2208)) or (layer2_outputs(731));
    layer3_outputs(371) <= (layer2_outputs(3584)) and not (layer2_outputs(1772));
    layer3_outputs(372) <= not((layer2_outputs(3176)) or (layer2_outputs(271)));
    layer3_outputs(373) <= not(layer2_outputs(4147)) or (layer2_outputs(2316));
    layer3_outputs(374) <= not(layer2_outputs(1374));
    layer3_outputs(375) <= layer2_outputs(1247);
    layer3_outputs(376) <= not((layer2_outputs(2237)) and (layer2_outputs(5037)));
    layer3_outputs(377) <= (layer2_outputs(4599)) and (layer2_outputs(3170));
    layer3_outputs(378) <= not(layer2_outputs(4956));
    layer3_outputs(379) <= (layer2_outputs(3880)) and not (layer2_outputs(660));
    layer3_outputs(380) <= not((layer2_outputs(2628)) and (layer2_outputs(3657)));
    layer3_outputs(381) <= (layer2_outputs(3950)) and not (layer2_outputs(4606));
    layer3_outputs(382) <= (layer2_outputs(3865)) and not (layer2_outputs(4023));
    layer3_outputs(383) <= (layer2_outputs(1706)) or (layer2_outputs(3688));
    layer3_outputs(384) <= (layer2_outputs(326)) and not (layer2_outputs(2683));
    layer3_outputs(385) <= not(layer2_outputs(2109));
    layer3_outputs(386) <= layer2_outputs(2163);
    layer3_outputs(387) <= '0';
    layer3_outputs(388) <= (layer2_outputs(1808)) and not (layer2_outputs(3978));
    layer3_outputs(389) <= not((layer2_outputs(3838)) and (layer2_outputs(4716)));
    layer3_outputs(390) <= not(layer2_outputs(3895));
    layer3_outputs(391) <= (layer2_outputs(1203)) and (layer2_outputs(184));
    layer3_outputs(392) <= not(layer2_outputs(2682));
    layer3_outputs(393) <= not(layer2_outputs(4714));
    layer3_outputs(394) <= layer2_outputs(785);
    layer3_outputs(395) <= not(layer2_outputs(3312));
    layer3_outputs(396) <= '0';
    layer3_outputs(397) <= '1';
    layer3_outputs(398) <= not(layer2_outputs(876));
    layer3_outputs(399) <= not(layer2_outputs(315));
    layer3_outputs(400) <= not((layer2_outputs(3019)) or (layer2_outputs(3847)));
    layer3_outputs(401) <= layer2_outputs(4836);
    layer3_outputs(402) <= layer2_outputs(5032);
    layer3_outputs(403) <= not(layer2_outputs(3081));
    layer3_outputs(404) <= layer2_outputs(2506);
    layer3_outputs(405) <= not(layer2_outputs(264));
    layer3_outputs(406) <= layer2_outputs(2381);
    layer3_outputs(407) <= layer2_outputs(3829);
    layer3_outputs(408) <= not(layer2_outputs(4564)) or (layer2_outputs(1580));
    layer3_outputs(409) <= '1';
    layer3_outputs(410) <= '1';
    layer3_outputs(411) <= '0';
    layer3_outputs(412) <= (layer2_outputs(2777)) or (layer2_outputs(443));
    layer3_outputs(413) <= '0';
    layer3_outputs(414) <= not(layer2_outputs(3720)) or (layer2_outputs(3768));
    layer3_outputs(415) <= not(layer2_outputs(3384));
    layer3_outputs(416) <= not(layer2_outputs(2315));
    layer3_outputs(417) <= layer2_outputs(4837);
    layer3_outputs(418) <= not(layer2_outputs(2278));
    layer3_outputs(419) <= not((layer2_outputs(4738)) or (layer2_outputs(4900)));
    layer3_outputs(420) <= not((layer2_outputs(1643)) xor (layer2_outputs(621)));
    layer3_outputs(421) <= not(layer2_outputs(1069));
    layer3_outputs(422) <= (layer2_outputs(478)) and not (layer2_outputs(809));
    layer3_outputs(423) <= not(layer2_outputs(153));
    layer3_outputs(424) <= layer2_outputs(3600);
    layer3_outputs(425) <= (layer2_outputs(3707)) and not (layer2_outputs(754));
    layer3_outputs(426) <= not((layer2_outputs(2051)) xor (layer2_outputs(811)));
    layer3_outputs(427) <= not((layer2_outputs(655)) or (layer2_outputs(2923)));
    layer3_outputs(428) <= not(layer2_outputs(1535));
    layer3_outputs(429) <= not(layer2_outputs(5015));
    layer3_outputs(430) <= not(layer2_outputs(4960));
    layer3_outputs(431) <= '1';
    layer3_outputs(432) <= '1';
    layer3_outputs(433) <= layer2_outputs(2855);
    layer3_outputs(434) <= layer2_outputs(3086);
    layer3_outputs(435) <= layer2_outputs(1630);
    layer3_outputs(436) <= not((layer2_outputs(116)) and (layer2_outputs(2460)));
    layer3_outputs(437) <= (layer2_outputs(4086)) or (layer2_outputs(172));
    layer3_outputs(438) <= not(layer2_outputs(4737)) or (layer2_outputs(1703));
    layer3_outputs(439) <= (layer2_outputs(3027)) and not (layer2_outputs(3229));
    layer3_outputs(440) <= not((layer2_outputs(941)) and (layer2_outputs(1313)));
    layer3_outputs(441) <= not(layer2_outputs(423));
    layer3_outputs(442) <= (layer2_outputs(3446)) and (layer2_outputs(83));
    layer3_outputs(443) <= not(layer2_outputs(2438));
    layer3_outputs(444) <= '1';
    layer3_outputs(445) <= '0';
    layer3_outputs(446) <= (layer2_outputs(2717)) and not (layer2_outputs(1878));
    layer3_outputs(447) <= layer2_outputs(3314);
    layer3_outputs(448) <= layer2_outputs(1155);
    layer3_outputs(449) <= (layer2_outputs(4000)) or (layer2_outputs(356));
    layer3_outputs(450) <= layer2_outputs(1288);
    layer3_outputs(451) <= not(layer2_outputs(4580));
    layer3_outputs(452) <= (layer2_outputs(1162)) and (layer2_outputs(4400));
    layer3_outputs(453) <= not(layer2_outputs(3387)) or (layer2_outputs(265));
    layer3_outputs(454) <= (layer2_outputs(1891)) and (layer2_outputs(543));
    layer3_outputs(455) <= not(layer2_outputs(1375));
    layer3_outputs(456) <= (layer2_outputs(4452)) and not (layer2_outputs(3632));
    layer3_outputs(457) <= layer2_outputs(4148);
    layer3_outputs(458) <= '0';
    layer3_outputs(459) <= layer2_outputs(1940);
    layer3_outputs(460) <= (layer2_outputs(3820)) xor (layer2_outputs(3377));
    layer3_outputs(461) <= layer2_outputs(4949);
    layer3_outputs(462) <= (layer2_outputs(3751)) and (layer2_outputs(2727));
    layer3_outputs(463) <= '0';
    layer3_outputs(464) <= not(layer2_outputs(1191)) or (layer2_outputs(2344));
    layer3_outputs(465) <= layer2_outputs(2056);
    layer3_outputs(466) <= layer2_outputs(298);
    layer3_outputs(467) <= (layer2_outputs(861)) and (layer2_outputs(5097));
    layer3_outputs(468) <= layer2_outputs(3692);
    layer3_outputs(469) <= not((layer2_outputs(3303)) and (layer2_outputs(2356)));
    layer3_outputs(470) <= not((layer2_outputs(1840)) xor (layer2_outputs(1613)));
    layer3_outputs(471) <= not(layer2_outputs(5013));
    layer3_outputs(472) <= '1';
    layer3_outputs(473) <= (layer2_outputs(1621)) and not (layer2_outputs(4111));
    layer3_outputs(474) <= '0';
    layer3_outputs(475) <= not(layer2_outputs(3826));
    layer3_outputs(476) <= (layer2_outputs(4860)) and not (layer2_outputs(127));
    layer3_outputs(477) <= not(layer2_outputs(1263)) or (layer2_outputs(2989));
    layer3_outputs(478) <= not(layer2_outputs(512)) or (layer2_outputs(1016));
    layer3_outputs(479) <= not(layer2_outputs(4140));
    layer3_outputs(480) <= '0';
    layer3_outputs(481) <= '0';
    layer3_outputs(482) <= not(layer2_outputs(4037));
    layer3_outputs(483) <= not(layer2_outputs(352));
    layer3_outputs(484) <= '0';
    layer3_outputs(485) <= not((layer2_outputs(2973)) or (layer2_outputs(3106)));
    layer3_outputs(486) <= layer2_outputs(1471);
    layer3_outputs(487) <= '0';
    layer3_outputs(488) <= '1';
    layer3_outputs(489) <= layer2_outputs(146);
    layer3_outputs(490) <= (layer2_outputs(2634)) and not (layer2_outputs(1746));
    layer3_outputs(491) <= layer2_outputs(4317);
    layer3_outputs(492) <= layer2_outputs(4276);
    layer3_outputs(493) <= layer2_outputs(1625);
    layer3_outputs(494) <= layer2_outputs(94);
    layer3_outputs(495) <= not((layer2_outputs(3684)) xor (layer2_outputs(2871)));
    layer3_outputs(496) <= not(layer2_outputs(1827));
    layer3_outputs(497) <= not(layer2_outputs(4866));
    layer3_outputs(498) <= layer2_outputs(617);
    layer3_outputs(499) <= (layer2_outputs(4597)) and not (layer2_outputs(945));
    layer3_outputs(500) <= '1';
    layer3_outputs(501) <= '0';
    layer3_outputs(502) <= not(layer2_outputs(4809));
    layer3_outputs(503) <= not(layer2_outputs(983));
    layer3_outputs(504) <= not(layer2_outputs(2292));
    layer3_outputs(505) <= not(layer2_outputs(415)) or (layer2_outputs(3084));
    layer3_outputs(506) <= layer2_outputs(1395);
    layer3_outputs(507) <= '0';
    layer3_outputs(508) <= not((layer2_outputs(545)) and (layer2_outputs(3750)));
    layer3_outputs(509) <= not(layer2_outputs(4777)) or (layer2_outputs(3430));
    layer3_outputs(510) <= not(layer2_outputs(1172));
    layer3_outputs(511) <= not((layer2_outputs(1449)) or (layer2_outputs(761)));
    layer3_outputs(512) <= '0';
    layer3_outputs(513) <= not(layer2_outputs(455)) or (layer2_outputs(1133));
    layer3_outputs(514) <= layer2_outputs(2739);
    layer3_outputs(515) <= (layer2_outputs(3566)) and (layer2_outputs(1815));
    layer3_outputs(516) <= not(layer2_outputs(3902));
    layer3_outputs(517) <= not(layer2_outputs(777)) or (layer2_outputs(2660));
    layer3_outputs(518) <= layer2_outputs(1295);
    layer3_outputs(519) <= layer2_outputs(2722);
    layer3_outputs(520) <= layer2_outputs(4901);
    layer3_outputs(521) <= (layer2_outputs(2967)) and not (layer2_outputs(1460));
    layer3_outputs(522) <= (layer2_outputs(1766)) and not (layer2_outputs(4621));
    layer3_outputs(523) <= not((layer2_outputs(118)) or (layer2_outputs(2028)));
    layer3_outputs(524) <= '0';
    layer3_outputs(525) <= '0';
    layer3_outputs(526) <= not(layer2_outputs(2266)) or (layer2_outputs(2230));
    layer3_outputs(527) <= (layer2_outputs(1126)) and not (layer2_outputs(1891));
    layer3_outputs(528) <= not(layer2_outputs(1032)) or (layer2_outputs(3468));
    layer3_outputs(529) <= not((layer2_outputs(273)) xor (layer2_outputs(3932)));
    layer3_outputs(530) <= layer2_outputs(3188);
    layer3_outputs(531) <= not(layer2_outputs(1903)) or (layer2_outputs(894));
    layer3_outputs(532) <= '1';
    layer3_outputs(533) <= layer2_outputs(4948);
    layer3_outputs(534) <= (layer2_outputs(1230)) and (layer2_outputs(887));
    layer3_outputs(535) <= (layer2_outputs(995)) and (layer2_outputs(3512));
    layer3_outputs(536) <= (layer2_outputs(1038)) and (layer2_outputs(1769));
    layer3_outputs(537) <= (layer2_outputs(2892)) and not (layer2_outputs(4337));
    layer3_outputs(538) <= not((layer2_outputs(3676)) and (layer2_outputs(1954)));
    layer3_outputs(539) <= not(layer2_outputs(2707)) or (layer2_outputs(3108));
    layer3_outputs(540) <= not(layer2_outputs(4066)) or (layer2_outputs(568));
    layer3_outputs(541) <= not((layer2_outputs(4230)) and (layer2_outputs(4301)));
    layer3_outputs(542) <= layer2_outputs(1569);
    layer3_outputs(543) <= layer2_outputs(4861);
    layer3_outputs(544) <= layer2_outputs(3846);
    layer3_outputs(545) <= '1';
    layer3_outputs(546) <= (layer2_outputs(4734)) or (layer2_outputs(275));
    layer3_outputs(547) <= not(layer2_outputs(1837));
    layer3_outputs(548) <= layer2_outputs(1729);
    layer3_outputs(549) <= not(layer2_outputs(1090));
    layer3_outputs(550) <= layer2_outputs(659);
    layer3_outputs(551) <= not((layer2_outputs(211)) xor (layer2_outputs(3923)));
    layer3_outputs(552) <= (layer2_outputs(1881)) xor (layer2_outputs(3158));
    layer3_outputs(553) <= '0';
    layer3_outputs(554) <= (layer2_outputs(5005)) and not (layer2_outputs(1909));
    layer3_outputs(555) <= not(layer2_outputs(305));
    layer3_outputs(556) <= (layer2_outputs(3603)) and not (layer2_outputs(2357));
    layer3_outputs(557) <= not(layer2_outputs(1251)) or (layer2_outputs(4108));
    layer3_outputs(558) <= not((layer2_outputs(3110)) or (layer2_outputs(3238)));
    layer3_outputs(559) <= not(layer2_outputs(4209));
    layer3_outputs(560) <= (layer2_outputs(3264)) or (layer2_outputs(3481));
    layer3_outputs(561) <= '1';
    layer3_outputs(562) <= not(layer2_outputs(1611));
    layer3_outputs(563) <= layer2_outputs(920);
    layer3_outputs(564) <= layer2_outputs(3313);
    layer3_outputs(565) <= layer2_outputs(3160);
    layer3_outputs(566) <= '0';
    layer3_outputs(567) <= not(layer2_outputs(836));
    layer3_outputs(568) <= layer2_outputs(1004);
    layer3_outputs(569) <= '1';
    layer3_outputs(570) <= (layer2_outputs(4365)) or (layer2_outputs(4474));
    layer3_outputs(571) <= layer2_outputs(1058);
    layer3_outputs(572) <= (layer2_outputs(669)) and not (layer2_outputs(840));
    layer3_outputs(573) <= not(layer2_outputs(1831)) or (layer2_outputs(518));
    layer3_outputs(574) <= '1';
    layer3_outputs(575) <= not(layer2_outputs(985));
    layer3_outputs(576) <= '1';
    layer3_outputs(577) <= not(layer2_outputs(4308)) or (layer2_outputs(4983));
    layer3_outputs(578) <= not((layer2_outputs(1911)) or (layer2_outputs(993)));
    layer3_outputs(579) <= (layer2_outputs(5020)) and not (layer2_outputs(4835));
    layer3_outputs(580) <= (layer2_outputs(3922)) and not (layer2_outputs(4214));
    layer3_outputs(581) <= layer2_outputs(2042);
    layer3_outputs(582) <= not((layer2_outputs(3265)) or (layer2_outputs(3900)));
    layer3_outputs(583) <= (layer2_outputs(3550)) xor (layer2_outputs(4628));
    layer3_outputs(584) <= not(layer2_outputs(5119)) or (layer2_outputs(4568));
    layer3_outputs(585) <= (layer2_outputs(111)) or (layer2_outputs(5078));
    layer3_outputs(586) <= (layer2_outputs(2774)) and not (layer2_outputs(1306));
    layer3_outputs(587) <= not((layer2_outputs(1180)) and (layer2_outputs(3098)));
    layer3_outputs(588) <= not(layer2_outputs(25)) or (layer2_outputs(4971));
    layer3_outputs(589) <= (layer2_outputs(2212)) xor (layer2_outputs(780));
    layer3_outputs(590) <= not(layer2_outputs(1775));
    layer3_outputs(591) <= not((layer2_outputs(4587)) or (layer2_outputs(649)));
    layer3_outputs(592) <= not(layer2_outputs(566));
    layer3_outputs(593) <= not(layer2_outputs(855));
    layer3_outputs(594) <= '0';
    layer3_outputs(595) <= '1';
    layer3_outputs(596) <= (layer2_outputs(3939)) and not (layer2_outputs(2086));
    layer3_outputs(597) <= layer2_outputs(2993);
    layer3_outputs(598) <= (layer2_outputs(399)) or (layer2_outputs(3455));
    layer3_outputs(599) <= not(layer2_outputs(5090)) or (layer2_outputs(3963));
    layer3_outputs(600) <= (layer2_outputs(3748)) or (layer2_outputs(3536));
    layer3_outputs(601) <= (layer2_outputs(931)) or (layer2_outputs(1442));
    layer3_outputs(602) <= not(layer2_outputs(3403));
    layer3_outputs(603) <= layer2_outputs(4542);
    layer3_outputs(604) <= (layer2_outputs(505)) or (layer2_outputs(3986));
    layer3_outputs(605) <= '0';
    layer3_outputs(606) <= '1';
    layer3_outputs(607) <= '0';
    layer3_outputs(608) <= (layer2_outputs(1280)) and (layer2_outputs(3798));
    layer3_outputs(609) <= layer2_outputs(1825);
    layer3_outputs(610) <= not(layer2_outputs(441));
    layer3_outputs(611) <= not(layer2_outputs(4438)) or (layer2_outputs(522));
    layer3_outputs(612) <= not(layer2_outputs(2965)) or (layer2_outputs(2333));
    layer3_outputs(613) <= (layer2_outputs(3060)) and not (layer2_outputs(868));
    layer3_outputs(614) <= not(layer2_outputs(5002)) or (layer2_outputs(2067));
    layer3_outputs(615) <= (layer2_outputs(288)) and not (layer2_outputs(355));
    layer3_outputs(616) <= not(layer2_outputs(4009));
    layer3_outputs(617) <= not((layer2_outputs(2910)) or (layer2_outputs(3978)));
    layer3_outputs(618) <= layer2_outputs(1973);
    layer3_outputs(619) <= (layer2_outputs(2928)) and not (layer2_outputs(781));
    layer3_outputs(620) <= not((layer2_outputs(4120)) and (layer2_outputs(2698)));
    layer3_outputs(621) <= not(layer2_outputs(2515));
    layer3_outputs(622) <= not(layer2_outputs(3123)) or (layer2_outputs(4686));
    layer3_outputs(623) <= (layer2_outputs(3042)) or (layer2_outputs(171));
    layer3_outputs(624) <= not(layer2_outputs(3818));
    layer3_outputs(625) <= layer2_outputs(3537);
    layer3_outputs(626) <= not(layer2_outputs(4277));
    layer3_outputs(627) <= not(layer2_outputs(1045));
    layer3_outputs(628) <= not(layer2_outputs(1010)) or (layer2_outputs(3058));
    layer3_outputs(629) <= (layer2_outputs(1901)) and not (layer2_outputs(2694));
    layer3_outputs(630) <= not(layer2_outputs(2896)) or (layer2_outputs(2024));
    layer3_outputs(631) <= '0';
    layer3_outputs(632) <= not((layer2_outputs(450)) or (layer2_outputs(278)));
    layer3_outputs(633) <= (layer2_outputs(3169)) and not (layer2_outputs(2361));
    layer3_outputs(634) <= not((layer2_outputs(3916)) and (layer2_outputs(213)));
    layer3_outputs(635) <= (layer2_outputs(3825)) and not (layer2_outputs(2513));
    layer3_outputs(636) <= (layer2_outputs(726)) or (layer2_outputs(3303));
    layer3_outputs(637) <= not(layer2_outputs(2091)) or (layer2_outputs(2761));
    layer3_outputs(638) <= '0';
    layer3_outputs(639) <= not(layer2_outputs(4426)) or (layer2_outputs(4149));
    layer3_outputs(640) <= not(layer2_outputs(2145)) or (layer2_outputs(704));
    layer3_outputs(641) <= not(layer2_outputs(348)) or (layer2_outputs(840));
    layer3_outputs(642) <= not(layer2_outputs(80)) or (layer2_outputs(3013));
    layer3_outputs(643) <= (layer2_outputs(4326)) and not (layer2_outputs(3172));
    layer3_outputs(644) <= '0';
    layer3_outputs(645) <= not(layer2_outputs(3816));
    layer3_outputs(646) <= not(layer2_outputs(4692));
    layer3_outputs(647) <= '1';
    layer3_outputs(648) <= not(layer2_outputs(1187)) or (layer2_outputs(3528));
    layer3_outputs(649) <= (layer2_outputs(852)) and not (layer2_outputs(535));
    layer3_outputs(650) <= (layer2_outputs(1210)) and (layer2_outputs(3450));
    layer3_outputs(651) <= not((layer2_outputs(4136)) xor (layer2_outputs(4152)));
    layer3_outputs(652) <= (layer2_outputs(46)) and (layer2_outputs(3737));
    layer3_outputs(653) <= layer2_outputs(3457);
    layer3_outputs(654) <= (layer2_outputs(542)) and not (layer2_outputs(3020));
    layer3_outputs(655) <= (layer2_outputs(1638)) and not (layer2_outputs(2806));
    layer3_outputs(656) <= not(layer2_outputs(1700)) or (layer2_outputs(2437));
    layer3_outputs(657) <= not((layer2_outputs(4590)) and (layer2_outputs(3101)));
    layer3_outputs(658) <= (layer2_outputs(4907)) and (layer2_outputs(2329));
    layer3_outputs(659) <= '1';
    layer3_outputs(660) <= not(layer2_outputs(3681)) or (layer2_outputs(1785));
    layer3_outputs(661) <= not(layer2_outputs(1339));
    layer3_outputs(662) <= not(layer2_outputs(1247));
    layer3_outputs(663) <= '0';
    layer3_outputs(664) <= not(layer2_outputs(4489)) or (layer2_outputs(416));
    layer3_outputs(665) <= '1';
    layer3_outputs(666) <= (layer2_outputs(1113)) and (layer2_outputs(2532));
    layer3_outputs(667) <= layer2_outputs(4692);
    layer3_outputs(668) <= not(layer2_outputs(5084)) or (layer2_outputs(1774));
    layer3_outputs(669) <= (layer2_outputs(3456)) and not (layer2_outputs(4467));
    layer3_outputs(670) <= not(layer2_outputs(3114));
    layer3_outputs(671) <= '1';
    layer3_outputs(672) <= not(layer2_outputs(3731)) or (layer2_outputs(559));
    layer3_outputs(673) <= '1';
    layer3_outputs(674) <= not(layer2_outputs(2396));
    layer3_outputs(675) <= not(layer2_outputs(3579));
    layer3_outputs(676) <= not((layer2_outputs(4029)) or (layer2_outputs(3520)));
    layer3_outputs(677) <= (layer2_outputs(1697)) or (layer2_outputs(1141));
    layer3_outputs(678) <= (layer2_outputs(1704)) and (layer2_outputs(2423));
    layer3_outputs(679) <= '1';
    layer3_outputs(680) <= layer2_outputs(2023);
    layer3_outputs(681) <= not(layer2_outputs(1346));
    layer3_outputs(682) <= layer2_outputs(2210);
    layer3_outputs(683) <= layer2_outputs(953);
    layer3_outputs(684) <= not(layer2_outputs(1346)) or (layer2_outputs(141));
    layer3_outputs(685) <= layer2_outputs(3128);
    layer3_outputs(686) <= not(layer2_outputs(2159));
    layer3_outputs(687) <= (layer2_outputs(3060)) and not (layer2_outputs(3362));
    layer3_outputs(688) <= (layer2_outputs(1811)) and not (layer2_outputs(2796));
    layer3_outputs(689) <= not(layer2_outputs(2946));
    layer3_outputs(690) <= '1';
    layer3_outputs(691) <= (layer2_outputs(613)) and not (layer2_outputs(1316));
    layer3_outputs(692) <= not(layer2_outputs(8));
    layer3_outputs(693) <= not(layer2_outputs(110));
    layer3_outputs(694) <= '0';
    layer3_outputs(695) <= (layer2_outputs(2094)) and not (layer2_outputs(2275));
    layer3_outputs(696) <= (layer2_outputs(2472)) and not (layer2_outputs(1153));
    layer3_outputs(697) <= not(layer2_outputs(4540)) or (layer2_outputs(4704));
    layer3_outputs(698) <= not(layer2_outputs(834));
    layer3_outputs(699) <= layer2_outputs(2324);
    layer3_outputs(700) <= (layer2_outputs(1126)) and not (layer2_outputs(3984));
    layer3_outputs(701) <= not(layer2_outputs(4005)) or (layer2_outputs(853));
    layer3_outputs(702) <= not(layer2_outputs(2232));
    layer3_outputs(703) <= layer2_outputs(1556);
    layer3_outputs(704) <= not((layer2_outputs(4094)) and (layer2_outputs(2551)));
    layer3_outputs(705) <= not((layer2_outputs(4511)) and (layer2_outputs(270)));
    layer3_outputs(706) <= '1';
    layer3_outputs(707) <= layer2_outputs(2157);
    layer3_outputs(708) <= not((layer2_outputs(1420)) and (layer2_outputs(776)));
    layer3_outputs(709) <= not(layer2_outputs(3111));
    layer3_outputs(710) <= not(layer2_outputs(3958));
    layer3_outputs(711) <= layer2_outputs(3839);
    layer3_outputs(712) <= layer2_outputs(4862);
    layer3_outputs(713) <= layer2_outputs(4213);
    layer3_outputs(714) <= (layer2_outputs(695)) or (layer2_outputs(2377));
    layer3_outputs(715) <= not((layer2_outputs(1594)) xor (layer2_outputs(1767)));
    layer3_outputs(716) <= layer2_outputs(3701);
    layer3_outputs(717) <= not((layer2_outputs(5101)) or (layer2_outputs(1469)));
    layer3_outputs(718) <= (layer2_outputs(2618)) or (layer2_outputs(1648));
    layer3_outputs(719) <= (layer2_outputs(2440)) and not (layer2_outputs(4178));
    layer3_outputs(720) <= not((layer2_outputs(3615)) and (layer2_outputs(4330)));
    layer3_outputs(721) <= layer2_outputs(3352);
    layer3_outputs(722) <= layer2_outputs(866);
    layer3_outputs(723) <= not((layer2_outputs(1039)) and (layer2_outputs(2248)));
    layer3_outputs(724) <= not(layer2_outputs(2587)) or (layer2_outputs(882));
    layer3_outputs(725) <= not(layer2_outputs(1966)) or (layer2_outputs(4915));
    layer3_outputs(726) <= not(layer2_outputs(2592));
    layer3_outputs(727) <= not(layer2_outputs(3681)) or (layer2_outputs(1865));
    layer3_outputs(728) <= layer2_outputs(1044);
    layer3_outputs(729) <= '1';
    layer3_outputs(730) <= '0';
    layer3_outputs(731) <= layer2_outputs(3779);
    layer3_outputs(732) <= '0';
    layer3_outputs(733) <= (layer2_outputs(3382)) and not (layer2_outputs(4758));
    layer3_outputs(734) <= not((layer2_outputs(156)) and (layer2_outputs(4918)));
    layer3_outputs(735) <= not((layer2_outputs(1054)) and (layer2_outputs(670)));
    layer3_outputs(736) <= not(layer2_outputs(2012));
    layer3_outputs(737) <= not(layer2_outputs(3381));
    layer3_outputs(738) <= not((layer2_outputs(3379)) or (layer2_outputs(3029)));
    layer3_outputs(739) <= not(layer2_outputs(4053)) or (layer2_outputs(1086));
    layer3_outputs(740) <= '1';
    layer3_outputs(741) <= layer2_outputs(4238);
    layer3_outputs(742) <= not(layer2_outputs(2167));
    layer3_outputs(743) <= not(layer2_outputs(1123)) or (layer2_outputs(3351));
    layer3_outputs(744) <= '1';
    layer3_outputs(745) <= '1';
    layer3_outputs(746) <= not(layer2_outputs(3859));
    layer3_outputs(747) <= (layer2_outputs(602)) and not (layer2_outputs(604));
    layer3_outputs(748) <= not(layer2_outputs(3988));
    layer3_outputs(749) <= layer2_outputs(3192);
    layer3_outputs(750) <= layer2_outputs(906);
    layer3_outputs(751) <= layer2_outputs(4022);
    layer3_outputs(752) <= (layer2_outputs(16)) or (layer2_outputs(428));
    layer3_outputs(753) <= not(layer2_outputs(2357)) or (layer2_outputs(3771));
    layer3_outputs(754) <= (layer2_outputs(3970)) and not (layer2_outputs(2195));
    layer3_outputs(755) <= (layer2_outputs(893)) and not (layer2_outputs(1579));
    layer3_outputs(756) <= not(layer2_outputs(519));
    layer3_outputs(757) <= (layer2_outputs(2458)) and not (layer2_outputs(3157));
    layer3_outputs(758) <= layer2_outputs(4887);
    layer3_outputs(759) <= not(layer2_outputs(358));
    layer3_outputs(760) <= not(layer2_outputs(959));
    layer3_outputs(761) <= not(layer2_outputs(753));
    layer3_outputs(762) <= (layer2_outputs(2253)) and not (layer2_outputs(4019));
    layer3_outputs(763) <= (layer2_outputs(3840)) and not (layer2_outputs(507));
    layer3_outputs(764) <= (layer2_outputs(242)) and not (layer2_outputs(915));
    layer3_outputs(765) <= (layer2_outputs(1762)) and not (layer2_outputs(2849));
    layer3_outputs(766) <= not(layer2_outputs(4900));
    layer3_outputs(767) <= layer2_outputs(3708);
    layer3_outputs(768) <= layer2_outputs(3883);
    layer3_outputs(769) <= '1';
    layer3_outputs(770) <= '0';
    layer3_outputs(771) <= layer2_outputs(4346);
    layer3_outputs(772) <= not(layer2_outputs(2940)) or (layer2_outputs(5064));
    layer3_outputs(773) <= layer2_outputs(2876);
    layer3_outputs(774) <= (layer2_outputs(2767)) and (layer2_outputs(3944));
    layer3_outputs(775) <= layer2_outputs(2679);
    layer3_outputs(776) <= (layer2_outputs(3349)) and (layer2_outputs(315));
    layer3_outputs(777) <= '0';
    layer3_outputs(778) <= not(layer2_outputs(3497)) or (layer2_outputs(2279));
    layer3_outputs(779) <= (layer2_outputs(4410)) or (layer2_outputs(1565));
    layer3_outputs(780) <= not(layer2_outputs(2533)) or (layer2_outputs(1298));
    layer3_outputs(781) <= not((layer2_outputs(268)) and (layer2_outputs(4430)));
    layer3_outputs(782) <= not(layer2_outputs(190)) or (layer2_outputs(3199));
    layer3_outputs(783) <= not(layer2_outputs(2377));
    layer3_outputs(784) <= (layer2_outputs(2583)) and not (layer2_outputs(3457));
    layer3_outputs(785) <= not((layer2_outputs(2506)) xor (layer2_outputs(5087)));
    layer3_outputs(786) <= not(layer2_outputs(2579)) or (layer2_outputs(3448));
    layer3_outputs(787) <= '1';
    layer3_outputs(788) <= not(layer2_outputs(2982));
    layer3_outputs(789) <= layer2_outputs(639);
    layer3_outputs(790) <= not(layer2_outputs(2576)) or (layer2_outputs(3740));
    layer3_outputs(791) <= not(layer2_outputs(4037));
    layer3_outputs(792) <= not((layer2_outputs(4532)) and (layer2_outputs(699)));
    layer3_outputs(793) <= not(layer2_outputs(641));
    layer3_outputs(794) <= '0';
    layer3_outputs(795) <= not(layer2_outputs(3807));
    layer3_outputs(796) <= not((layer2_outputs(125)) and (layer2_outputs(4634)));
    layer3_outputs(797) <= '0';
    layer3_outputs(798) <= layer2_outputs(2630);
    layer3_outputs(799) <= not(layer2_outputs(1669));
    layer3_outputs(800) <= '0';
    layer3_outputs(801) <= not((layer2_outputs(4647)) or (layer2_outputs(4210)));
    layer3_outputs(802) <= not((layer2_outputs(2928)) and (layer2_outputs(3963)));
    layer3_outputs(803) <= not(layer2_outputs(5102)) or (layer2_outputs(3066));
    layer3_outputs(804) <= layer2_outputs(2132);
    layer3_outputs(805) <= not(layer2_outputs(3601));
    layer3_outputs(806) <= (layer2_outputs(3419)) or (layer2_outputs(4624));
    layer3_outputs(807) <= not((layer2_outputs(347)) and (layer2_outputs(92)));
    layer3_outputs(808) <= not((layer2_outputs(2934)) or (layer2_outputs(2454)));
    layer3_outputs(809) <= layer2_outputs(74);
    layer3_outputs(810) <= layer2_outputs(2940);
    layer3_outputs(811) <= layer2_outputs(2778);
    layer3_outputs(812) <= (layer2_outputs(3766)) and not (layer2_outputs(91));
    layer3_outputs(813) <= not(layer2_outputs(4996));
    layer3_outputs(814) <= layer2_outputs(17);
    layer3_outputs(815) <= (layer2_outputs(4494)) and not (layer2_outputs(5065));
    layer3_outputs(816) <= (layer2_outputs(4868)) and not (layer2_outputs(303));
    layer3_outputs(817) <= not((layer2_outputs(4908)) or (layer2_outputs(2561)));
    layer3_outputs(818) <= layer2_outputs(3535);
    layer3_outputs(819) <= '1';
    layer3_outputs(820) <= layer2_outputs(2143);
    layer3_outputs(821) <= not(layer2_outputs(1001));
    layer3_outputs(822) <= not(layer2_outputs(3298));
    layer3_outputs(823) <= layer2_outputs(4840);
    layer3_outputs(824) <= not(layer2_outputs(2849)) or (layer2_outputs(3899));
    layer3_outputs(825) <= layer2_outputs(1714);
    layer3_outputs(826) <= not((layer2_outputs(2990)) or (layer2_outputs(1602)));
    layer3_outputs(827) <= '0';
    layer3_outputs(828) <= layer2_outputs(2583);
    layer3_outputs(829) <= not((layer2_outputs(1948)) or (layer2_outputs(1278)));
    layer3_outputs(830) <= not(layer2_outputs(2554));
    layer3_outputs(831) <= not(layer2_outputs(2980));
    layer3_outputs(832) <= not((layer2_outputs(3342)) or (layer2_outputs(3202)));
    layer3_outputs(833) <= not(layer2_outputs(3573));
    layer3_outputs(834) <= not(layer2_outputs(5030));
    layer3_outputs(835) <= (layer2_outputs(4964)) or (layer2_outputs(1933));
    layer3_outputs(836) <= not((layer2_outputs(4658)) or (layer2_outputs(3592)));
    layer3_outputs(837) <= layer2_outputs(4867);
    layer3_outputs(838) <= not(layer2_outputs(1274));
    layer3_outputs(839) <= layer2_outputs(1897);
    layer3_outputs(840) <= not(layer2_outputs(2159));
    layer3_outputs(841) <= not(layer2_outputs(4003)) or (layer2_outputs(3606));
    layer3_outputs(842) <= layer2_outputs(2179);
    layer3_outputs(843) <= '0';
    layer3_outputs(844) <= (layer2_outputs(772)) and not (layer2_outputs(952));
    layer3_outputs(845) <= not((layer2_outputs(4421)) or (layer2_outputs(683)));
    layer3_outputs(846) <= layer2_outputs(2416);
    layer3_outputs(847) <= not((layer2_outputs(3640)) and (layer2_outputs(4984)));
    layer3_outputs(848) <= not(layer2_outputs(10));
    layer3_outputs(849) <= layer2_outputs(2401);
    layer3_outputs(850) <= (layer2_outputs(510)) and not (layer2_outputs(276));
    layer3_outputs(851) <= '0';
    layer3_outputs(852) <= not(layer2_outputs(4731));
    layer3_outputs(853) <= not(layer2_outputs(2023));
    layer3_outputs(854) <= layer2_outputs(3800);
    layer3_outputs(855) <= not((layer2_outputs(3351)) xor (layer2_outputs(1801)));
    layer3_outputs(856) <= not(layer2_outputs(572));
    layer3_outputs(857) <= not(layer2_outputs(719));
    layer3_outputs(858) <= layer2_outputs(1203);
    layer3_outputs(859) <= layer2_outputs(2010);
    layer3_outputs(860) <= (layer2_outputs(4398)) xor (layer2_outputs(4364));
    layer3_outputs(861) <= layer2_outputs(2349);
    layer3_outputs(862) <= (layer2_outputs(4264)) and (layer2_outputs(4298));
    layer3_outputs(863) <= '1';
    layer3_outputs(864) <= layer2_outputs(4921);
    layer3_outputs(865) <= not((layer2_outputs(534)) and (layer2_outputs(1011)));
    layer3_outputs(866) <= (layer2_outputs(4528)) xor (layer2_outputs(4929));
    layer3_outputs(867) <= layer2_outputs(3166);
    layer3_outputs(868) <= layer2_outputs(2078);
    layer3_outputs(869) <= (layer2_outputs(2855)) and not (layer2_outputs(95));
    layer3_outputs(870) <= layer2_outputs(4324);
    layer3_outputs(871) <= (layer2_outputs(2165)) or (layer2_outputs(2027));
    layer3_outputs(872) <= (layer2_outputs(395)) and not (layer2_outputs(3565));
    layer3_outputs(873) <= (layer2_outputs(2338)) and (layer2_outputs(824));
    layer3_outputs(874) <= not(layer2_outputs(3589));
    layer3_outputs(875) <= not(layer2_outputs(5102)) or (layer2_outputs(3214));
    layer3_outputs(876) <= layer2_outputs(105);
    layer3_outputs(877) <= layer2_outputs(898);
    layer3_outputs(878) <= not(layer2_outputs(4535)) or (layer2_outputs(2966));
    layer3_outputs(879) <= (layer2_outputs(4688)) and (layer2_outputs(2004));
    layer3_outputs(880) <= (layer2_outputs(2710)) or (layer2_outputs(4022));
    layer3_outputs(881) <= (layer2_outputs(3294)) or (layer2_outputs(3902));
    layer3_outputs(882) <= (layer2_outputs(1308)) and not (layer2_outputs(4971));
    layer3_outputs(883) <= not(layer2_outputs(3652));
    layer3_outputs(884) <= '0';
    layer3_outputs(885) <= (layer2_outputs(3852)) and (layer2_outputs(2800));
    layer3_outputs(886) <= layer2_outputs(1281);
    layer3_outputs(887) <= '1';
    layer3_outputs(888) <= layer2_outputs(1454);
    layer3_outputs(889) <= not((layer2_outputs(310)) or (layer2_outputs(1374)));
    layer3_outputs(890) <= not(layer2_outputs(1427));
    layer3_outputs(891) <= not(layer2_outputs(1027)) or (layer2_outputs(403));
    layer3_outputs(892) <= not((layer2_outputs(1006)) xor (layer2_outputs(2493)));
    layer3_outputs(893) <= (layer2_outputs(657)) or (layer2_outputs(200));
    layer3_outputs(894) <= '0';
    layer3_outputs(895) <= (layer2_outputs(1862)) or (layer2_outputs(1939));
    layer3_outputs(896) <= not(layer2_outputs(1808));
    layer3_outputs(897) <= '0';
    layer3_outputs(898) <= not(layer2_outputs(2841)) or (layer2_outputs(3335));
    layer3_outputs(899) <= layer2_outputs(4620);
    layer3_outputs(900) <= (layer2_outputs(96)) and not (layer2_outputs(784));
    layer3_outputs(901) <= '1';
    layer3_outputs(902) <= '0';
    layer3_outputs(903) <= not((layer2_outputs(2332)) or (layer2_outputs(3102)));
    layer3_outputs(904) <= layer2_outputs(4105);
    layer3_outputs(905) <= not(layer2_outputs(3458));
    layer3_outputs(906) <= not(layer2_outputs(2283));
    layer3_outputs(907) <= layer2_outputs(1996);
    layer3_outputs(908) <= not(layer2_outputs(3050)) or (layer2_outputs(2895));
    layer3_outputs(909) <= (layer2_outputs(1151)) and not (layer2_outputs(4589));
    layer3_outputs(910) <= layer2_outputs(2571);
    layer3_outputs(911) <= layer2_outputs(585);
    layer3_outputs(912) <= not(layer2_outputs(1610));
    layer3_outputs(913) <= layer2_outputs(299);
    layer3_outputs(914) <= not(layer2_outputs(3073));
    layer3_outputs(915) <= (layer2_outputs(4519)) and not (layer2_outputs(1125));
    layer3_outputs(916) <= (layer2_outputs(1051)) and not (layer2_outputs(1245));
    layer3_outputs(917) <= (layer2_outputs(4645)) and not (layer2_outputs(3503));
    layer3_outputs(918) <= (layer2_outputs(2266)) and (layer2_outputs(4354));
    layer3_outputs(919) <= (layer2_outputs(2214)) and (layer2_outputs(3168));
    layer3_outputs(920) <= not(layer2_outputs(2790)) or (layer2_outputs(3253));
    layer3_outputs(921) <= not((layer2_outputs(2843)) or (layer2_outputs(3697)));
    layer3_outputs(922) <= not(layer2_outputs(1960));
    layer3_outputs(923) <= not(layer2_outputs(4947)) or (layer2_outputs(2432));
    layer3_outputs(924) <= not(layer2_outputs(569)) or (layer2_outputs(2113));
    layer3_outputs(925) <= (layer2_outputs(424)) and (layer2_outputs(5107));
    layer3_outputs(926) <= (layer2_outputs(3942)) or (layer2_outputs(665));
    layer3_outputs(927) <= (layer2_outputs(4065)) and not (layer2_outputs(2452));
    layer3_outputs(928) <= (layer2_outputs(2181)) xor (layer2_outputs(1997));
    layer3_outputs(929) <= not(layer2_outputs(4399));
    layer3_outputs(930) <= (layer2_outputs(2061)) and not (layer2_outputs(833));
    layer3_outputs(931) <= not((layer2_outputs(201)) or (layer2_outputs(2479)));
    layer3_outputs(932) <= not(layer2_outputs(110));
    layer3_outputs(933) <= (layer2_outputs(3001)) and (layer2_outputs(3552));
    layer3_outputs(934) <= not(layer2_outputs(673));
    layer3_outputs(935) <= not(layer2_outputs(234)) or (layer2_outputs(2688));
    layer3_outputs(936) <= (layer2_outputs(4195)) and (layer2_outputs(3974));
    layer3_outputs(937) <= layer2_outputs(2905);
    layer3_outputs(938) <= (layer2_outputs(1393)) and not (layer2_outputs(413));
    layer3_outputs(939) <= not(layer2_outputs(4055));
    layer3_outputs(940) <= '0';
    layer3_outputs(941) <= layer2_outputs(4320);
    layer3_outputs(942) <= layer2_outputs(1673);
    layer3_outputs(943) <= not(layer2_outputs(2793));
    layer3_outputs(944) <= not(layer2_outputs(1260));
    layer3_outputs(945) <= '0';
    layer3_outputs(946) <= not((layer2_outputs(4647)) xor (layer2_outputs(914)));
    layer3_outputs(947) <= layer2_outputs(2421);
    layer3_outputs(948) <= not(layer2_outputs(4241)) or (layer2_outputs(4698));
    layer3_outputs(949) <= (layer2_outputs(4569)) or (layer2_outputs(18));
    layer3_outputs(950) <= layer2_outputs(4453);
    layer3_outputs(951) <= not(layer2_outputs(2523)) or (layer2_outputs(2544));
    layer3_outputs(952) <= not(layer2_outputs(2649));
    layer3_outputs(953) <= not(layer2_outputs(1548)) or (layer2_outputs(3560));
    layer3_outputs(954) <= (layer2_outputs(850)) or (layer2_outputs(1079));
    layer3_outputs(955) <= not(layer2_outputs(1728));
    layer3_outputs(956) <= layer2_outputs(1629);
    layer3_outputs(957) <= layer2_outputs(512);
    layer3_outputs(958) <= (layer2_outputs(2469)) and not (layer2_outputs(4036));
    layer3_outputs(959) <= not((layer2_outputs(2935)) or (layer2_outputs(2705)));
    layer3_outputs(960) <= (layer2_outputs(1626)) and not (layer2_outputs(4303));
    layer3_outputs(961) <= not(layer2_outputs(584));
    layer3_outputs(962) <= '1';
    layer3_outputs(963) <= not(layer2_outputs(4134));
    layer3_outputs(964) <= not(layer2_outputs(485));
    layer3_outputs(965) <= not(layer2_outputs(2492));
    layer3_outputs(966) <= '1';
    layer3_outputs(967) <= not((layer2_outputs(1593)) or (layer2_outputs(3181)));
    layer3_outputs(968) <= (layer2_outputs(1064)) and not (layer2_outputs(343));
    layer3_outputs(969) <= not(layer2_outputs(1034)) or (layer2_outputs(3814));
    layer3_outputs(970) <= (layer2_outputs(2582)) and (layer2_outputs(1036));
    layer3_outputs(971) <= not(layer2_outputs(2556));
    layer3_outputs(972) <= not(layer2_outputs(2746));
    layer3_outputs(973) <= not(layer2_outputs(2258));
    layer3_outputs(974) <= layer2_outputs(4421);
    layer3_outputs(975) <= not(layer2_outputs(4157));
    layer3_outputs(976) <= not((layer2_outputs(3882)) xor (layer2_outputs(734)));
    layer3_outputs(977) <= not(layer2_outputs(3116));
    layer3_outputs(978) <= '0';
    layer3_outputs(979) <= layer2_outputs(1421);
    layer3_outputs(980) <= layer2_outputs(4268);
    layer3_outputs(981) <= not(layer2_outputs(3418)) or (layer2_outputs(4472));
    layer3_outputs(982) <= '0';
    layer3_outputs(983) <= '0';
    layer3_outputs(984) <= (layer2_outputs(1352)) and not (layer2_outputs(3414));
    layer3_outputs(985) <= (layer2_outputs(3568)) and not (layer2_outputs(2892));
    layer3_outputs(986) <= not(layer2_outputs(3725));
    layer3_outputs(987) <= '1';
    layer3_outputs(988) <= layer2_outputs(3008);
    layer3_outputs(989) <= not(layer2_outputs(4865));
    layer3_outputs(990) <= (layer2_outputs(3523)) and not (layer2_outputs(4572));
    layer3_outputs(991) <= '1';
    layer3_outputs(992) <= not((layer2_outputs(2157)) or (layer2_outputs(310)));
    layer3_outputs(993) <= layer2_outputs(1294);
    layer3_outputs(994) <= not((layer2_outputs(4209)) or (layer2_outputs(5119)));
    layer3_outputs(995) <= not(layer2_outputs(5001));
    layer3_outputs(996) <= not(layer2_outputs(3234)) or (layer2_outputs(4082));
    layer3_outputs(997) <= '0';
    layer3_outputs(998) <= '1';
    layer3_outputs(999) <= not(layer2_outputs(3247)) or (layer2_outputs(2347));
    layer3_outputs(1000) <= (layer2_outputs(4011)) and not (layer2_outputs(3656));
    layer3_outputs(1001) <= '0';
    layer3_outputs(1002) <= not(layer2_outputs(3935)) or (layer2_outputs(631));
    layer3_outputs(1003) <= (layer2_outputs(1368)) xor (layer2_outputs(848));
    layer3_outputs(1004) <= '0';
    layer3_outputs(1005) <= not(layer2_outputs(4427));
    layer3_outputs(1006) <= not((layer2_outputs(4636)) or (layer2_outputs(4633)));
    layer3_outputs(1007) <= (layer2_outputs(3364)) and not (layer2_outputs(1073));
    layer3_outputs(1008) <= (layer2_outputs(2417)) or (layer2_outputs(335));
    layer3_outputs(1009) <= (layer2_outputs(3258)) and not (layer2_outputs(3220));
    layer3_outputs(1010) <= not((layer2_outputs(1951)) or (layer2_outputs(1080)));
    layer3_outputs(1011) <= not(layer2_outputs(4441));
    layer3_outputs(1012) <= (layer2_outputs(4182)) and not (layer2_outputs(2013));
    layer3_outputs(1013) <= (layer2_outputs(3767)) and not (layer2_outputs(4120));
    layer3_outputs(1014) <= not(layer2_outputs(2206)) or (layer2_outputs(3248));
    layer3_outputs(1015) <= layer2_outputs(1696);
    layer3_outputs(1016) <= not((layer2_outputs(1970)) or (layer2_outputs(803)));
    layer3_outputs(1017) <= not(layer2_outputs(4024));
    layer3_outputs(1018) <= (layer2_outputs(2489)) and not (layer2_outputs(2085));
    layer3_outputs(1019) <= layer2_outputs(3894);
    layer3_outputs(1020) <= layer2_outputs(970);
    layer3_outputs(1021) <= not(layer2_outputs(2359)) or (layer2_outputs(1712));
    layer3_outputs(1022) <= not(layer2_outputs(1742)) or (layer2_outputs(2289));
    layer3_outputs(1023) <= not(layer2_outputs(2112));
    layer3_outputs(1024) <= (layer2_outputs(2621)) or (layer2_outputs(1691));
    layer3_outputs(1025) <= '0';
    layer3_outputs(1026) <= not(layer2_outputs(4651));
    layer3_outputs(1027) <= (layer2_outputs(4184)) or (layer2_outputs(4281));
    layer3_outputs(1028) <= not(layer2_outputs(1194));
    layer3_outputs(1029) <= not(layer2_outputs(4572));
    layer3_outputs(1030) <= layer2_outputs(396);
    layer3_outputs(1031) <= layer2_outputs(2135);
    layer3_outputs(1032) <= not(layer2_outputs(2817));
    layer3_outputs(1033) <= not(layer2_outputs(2259));
    layer3_outputs(1034) <= not(layer2_outputs(4749));
    layer3_outputs(1035) <= not(layer2_outputs(2487));
    layer3_outputs(1036) <= not(layer2_outputs(3773));
    layer3_outputs(1037) <= not(layer2_outputs(4760));
    layer3_outputs(1038) <= '0';
    layer3_outputs(1039) <= not(layer2_outputs(781)) or (layer2_outputs(961));
    layer3_outputs(1040) <= layer2_outputs(4015);
    layer3_outputs(1041) <= '0';
    layer3_outputs(1042) <= not((layer2_outputs(1184)) and (layer2_outputs(1911)));
    layer3_outputs(1043) <= layer2_outputs(3148);
    layer3_outputs(1044) <= not(layer2_outputs(229)) or (layer2_outputs(3215));
    layer3_outputs(1045) <= '0';
    layer3_outputs(1046) <= layer2_outputs(723);
    layer3_outputs(1047) <= (layer2_outputs(1874)) and (layer2_outputs(357));
    layer3_outputs(1048) <= not(layer2_outputs(616));
    layer3_outputs(1049) <= not(layer2_outputs(3815));
    layer3_outputs(1050) <= (layer2_outputs(2563)) and (layer2_outputs(1694));
    layer3_outputs(1051) <= (layer2_outputs(1939)) or (layer2_outputs(4773));
    layer3_outputs(1052) <= '0';
    layer3_outputs(1053) <= not(layer2_outputs(4166)) or (layer2_outputs(353));
    layer3_outputs(1054) <= not((layer2_outputs(97)) or (layer2_outputs(1278)));
    layer3_outputs(1055) <= (layer2_outputs(1828)) or (layer2_outputs(3201));
    layer3_outputs(1056) <= (layer2_outputs(2217)) and not (layer2_outputs(3487));
    layer3_outputs(1057) <= not(layer2_outputs(363)) or (layer2_outputs(3659));
    layer3_outputs(1058) <= not(layer2_outputs(2792));
    layer3_outputs(1059) <= not(layer2_outputs(483));
    layer3_outputs(1060) <= not((layer2_outputs(1110)) xor (layer2_outputs(4837)));
    layer3_outputs(1061) <= not(layer2_outputs(3525)) or (layer2_outputs(3832));
    layer3_outputs(1062) <= not(layer2_outputs(596)) or (layer2_outputs(196));
    layer3_outputs(1063) <= not(layer2_outputs(3581));
    layer3_outputs(1064) <= layer2_outputs(2451);
    layer3_outputs(1065) <= layer2_outputs(3774);
    layer3_outputs(1066) <= '1';
    layer3_outputs(1067) <= (layer2_outputs(4992)) and not (layer2_outputs(857));
    layer3_outputs(1068) <= not(layer2_outputs(3508));
    layer3_outputs(1069) <= not((layer2_outputs(4124)) and (layer2_outputs(1311)));
    layer3_outputs(1070) <= not((layer2_outputs(2908)) or (layer2_outputs(2870)));
    layer3_outputs(1071) <= layer2_outputs(4693);
    layer3_outputs(1072) <= not(layer2_outputs(773)) or (layer2_outputs(994));
    layer3_outputs(1073) <= layer2_outputs(465);
    layer3_outputs(1074) <= not(layer2_outputs(1915)) or (layer2_outputs(851));
    layer3_outputs(1075) <= not((layer2_outputs(5109)) or (layer2_outputs(701)));
    layer3_outputs(1076) <= not(layer2_outputs(4913));
    layer3_outputs(1077) <= not(layer2_outputs(258)) or (layer2_outputs(646));
    layer3_outputs(1078) <= not((layer2_outputs(2150)) or (layer2_outputs(3809)));
    layer3_outputs(1079) <= '0';
    layer3_outputs(1080) <= (layer2_outputs(4700)) or (layer2_outputs(2374));
    layer3_outputs(1081) <= (layer2_outputs(498)) and not (layer2_outputs(2669));
    layer3_outputs(1082) <= not(layer2_outputs(883)) or (layer2_outputs(4851));
    layer3_outputs(1083) <= layer2_outputs(127);
    layer3_outputs(1084) <= '1';
    layer3_outputs(1085) <= not(layer2_outputs(4795));
    layer3_outputs(1086) <= not(layer2_outputs(4680)) or (layer2_outputs(1959));
    layer3_outputs(1087) <= (layer2_outputs(260)) and (layer2_outputs(4496));
    layer3_outputs(1088) <= not(layer2_outputs(686)) or (layer2_outputs(763));
    layer3_outputs(1089) <= layer2_outputs(1098);
    layer3_outputs(1090) <= (layer2_outputs(4211)) or (layer2_outputs(638));
    layer3_outputs(1091) <= layer2_outputs(701);
    layer3_outputs(1092) <= layer2_outputs(4278);
    layer3_outputs(1093) <= (layer2_outputs(2264)) and not (layer2_outputs(1885));
    layer3_outputs(1094) <= layer2_outputs(4694);
    layer3_outputs(1095) <= not((layer2_outputs(762)) or (layer2_outputs(1392)));
    layer3_outputs(1096) <= not((layer2_outputs(1461)) or (layer2_outputs(3389)));
    layer3_outputs(1097) <= (layer2_outputs(4775)) or (layer2_outputs(2936));
    layer3_outputs(1098) <= not(layer2_outputs(119)) or (layer2_outputs(4216));
    layer3_outputs(1099) <= not(layer2_outputs(578)) or (layer2_outputs(4747));
    layer3_outputs(1100) <= (layer2_outputs(1279)) and not (layer2_outputs(3743));
    layer3_outputs(1101) <= not((layer2_outputs(1685)) or (layer2_outputs(5023)));
    layer3_outputs(1102) <= layer2_outputs(4877);
    layer3_outputs(1103) <= layer2_outputs(3791);
    layer3_outputs(1104) <= layer2_outputs(1472);
    layer3_outputs(1105) <= not((layer2_outputs(2630)) and (layer2_outputs(526)));
    layer3_outputs(1106) <= layer2_outputs(1859);
    layer3_outputs(1107) <= not(layer2_outputs(401));
    layer3_outputs(1108) <= not((layer2_outputs(3005)) or (layer2_outputs(1598)));
    layer3_outputs(1109) <= not(layer2_outputs(1389));
    layer3_outputs(1110) <= layer2_outputs(2968);
    layer3_outputs(1111) <= not(layer2_outputs(4730));
    layer3_outputs(1112) <= (layer2_outputs(4562)) and (layer2_outputs(2045));
    layer3_outputs(1113) <= not((layer2_outputs(5033)) and (layer2_outputs(703)));
    layer3_outputs(1114) <= '1';
    layer3_outputs(1115) <= '1';
    layer3_outputs(1116) <= (layer2_outputs(4850)) and not (layer2_outputs(4935));
    layer3_outputs(1117) <= not(layer2_outputs(1676));
    layer3_outputs(1118) <= not(layer2_outputs(1616));
    layer3_outputs(1119) <= not(layer2_outputs(809));
    layer3_outputs(1120) <= not(layer2_outputs(161));
    layer3_outputs(1121) <= not((layer2_outputs(3586)) and (layer2_outputs(4942)));
    layer3_outputs(1122) <= not(layer2_outputs(4615));
    layer3_outputs(1123) <= not((layer2_outputs(3070)) and (layer2_outputs(1868)));
    layer3_outputs(1124) <= '1';
    layer3_outputs(1125) <= not((layer2_outputs(4523)) or (layer2_outputs(3604)));
    layer3_outputs(1126) <= not(layer2_outputs(285));
    layer3_outputs(1127) <= not(layer2_outputs(4454));
    layer3_outputs(1128) <= not(layer2_outputs(2809)) or (layer2_outputs(367));
    layer3_outputs(1129) <= (layer2_outputs(3355)) or (layer2_outputs(4048));
    layer3_outputs(1130) <= not(layer2_outputs(1454)) or (layer2_outputs(3590));
    layer3_outputs(1131) <= '1';
    layer3_outputs(1132) <= '1';
    layer3_outputs(1133) <= layer2_outputs(2077);
    layer3_outputs(1134) <= '0';
    layer3_outputs(1135) <= not(layer2_outputs(1469));
    layer3_outputs(1136) <= '1';
    layer3_outputs(1137) <= not((layer2_outputs(1782)) or (layer2_outputs(4637)));
    layer3_outputs(1138) <= layer2_outputs(3836);
    layer3_outputs(1139) <= not(layer2_outputs(1465));
    layer3_outputs(1140) <= layer2_outputs(2914);
    layer3_outputs(1141) <= not(layer2_outputs(3047));
    layer3_outputs(1142) <= not((layer2_outputs(2954)) and (layer2_outputs(1181)));
    layer3_outputs(1143) <= not(layer2_outputs(1788));
    layer3_outputs(1144) <= '0';
    layer3_outputs(1145) <= not(layer2_outputs(4896)) or (layer2_outputs(2375));
    layer3_outputs(1146) <= layer2_outputs(1701);
    layer3_outputs(1147) <= not(layer2_outputs(3405));
    layer3_outputs(1148) <= not(layer2_outputs(4238));
    layer3_outputs(1149) <= not(layer2_outputs(1197));
    layer3_outputs(1150) <= layer2_outputs(3273);
    layer3_outputs(1151) <= (layer2_outputs(4440)) and not (layer2_outputs(338));
    layer3_outputs(1152) <= (layer2_outputs(3084)) and not (layer2_outputs(2499));
    layer3_outputs(1153) <= (layer2_outputs(4650)) and (layer2_outputs(2664));
    layer3_outputs(1154) <= not(layer2_outputs(1814)) or (layer2_outputs(3273));
    layer3_outputs(1155) <= (layer2_outputs(1714)) and (layer2_outputs(3744));
    layer3_outputs(1156) <= not((layer2_outputs(982)) or (layer2_outputs(1143)));
    layer3_outputs(1157) <= (layer2_outputs(1823)) and not (layer2_outputs(2580));
    layer3_outputs(1158) <= not((layer2_outputs(3370)) xor (layer2_outputs(4611)));
    layer3_outputs(1159) <= not(layer2_outputs(3899));
    layer3_outputs(1160) <= not(layer2_outputs(467)) or (layer2_outputs(4114));
    layer3_outputs(1161) <= (layer2_outputs(3440)) and (layer2_outputs(2228));
    layer3_outputs(1162) <= not(layer2_outputs(1208));
    layer3_outputs(1163) <= not(layer2_outputs(2627)) or (layer2_outputs(1740));
    layer3_outputs(1164) <= (layer2_outputs(3878)) and (layer2_outputs(4982));
    layer3_outputs(1165) <= not(layer2_outputs(2695));
    layer3_outputs(1166) <= not(layer2_outputs(1634)) or (layer2_outputs(1342));
    layer3_outputs(1167) <= not(layer2_outputs(430));
    layer3_outputs(1168) <= (layer2_outputs(1565)) or (layer2_outputs(1091));
    layer3_outputs(1169) <= (layer2_outputs(2151)) and not (layer2_outputs(3054));
    layer3_outputs(1170) <= '1';
    layer3_outputs(1171) <= not((layer2_outputs(5115)) and (layer2_outputs(2945)));
    layer3_outputs(1172) <= '1';
    layer3_outputs(1173) <= '0';
    layer3_outputs(1174) <= layer2_outputs(491);
    layer3_outputs(1175) <= not(layer2_outputs(4411));
    layer3_outputs(1176) <= not(layer2_outputs(2778));
    layer3_outputs(1177) <= layer2_outputs(5081);
    layer3_outputs(1178) <= (layer2_outputs(2111)) and not (layer2_outputs(3627));
    layer3_outputs(1179) <= layer2_outputs(3998);
    layer3_outputs(1180) <= not((layer2_outputs(4442)) and (layer2_outputs(4097)));
    layer3_outputs(1181) <= layer2_outputs(4419);
    layer3_outputs(1182) <= layer2_outputs(841);
    layer3_outputs(1183) <= (layer2_outputs(2880)) and not (layer2_outputs(1107));
    layer3_outputs(1184) <= '1';
    layer3_outputs(1185) <= not(layer2_outputs(144)) or (layer2_outputs(4759));
    layer3_outputs(1186) <= not(layer2_outputs(907)) or (layer2_outputs(961));
    layer3_outputs(1187) <= not(layer2_outputs(1340));
    layer3_outputs(1188) <= not(layer2_outputs(3580)) or (layer2_outputs(3986));
    layer3_outputs(1189) <= (layer2_outputs(1259)) or (layer2_outputs(3879));
    layer3_outputs(1190) <= not(layer2_outputs(618));
    layer3_outputs(1191) <= layer2_outputs(2268);
    layer3_outputs(1192) <= not((layer2_outputs(2648)) and (layer2_outputs(184)));
    layer3_outputs(1193) <= not(layer2_outputs(2255));
    layer3_outputs(1194) <= (layer2_outputs(2540)) or (layer2_outputs(4970));
    layer3_outputs(1195) <= not(layer2_outputs(637));
    layer3_outputs(1196) <= '1';
    layer3_outputs(1197) <= not(layer2_outputs(4124)) or (layer2_outputs(943));
    layer3_outputs(1198) <= layer2_outputs(2189);
    layer3_outputs(1199) <= not(layer2_outputs(3371));
    layer3_outputs(1200) <= not(layer2_outputs(1998));
    layer3_outputs(1201) <= not(layer2_outputs(5027));
    layer3_outputs(1202) <= not((layer2_outputs(3014)) or (layer2_outputs(3021)));
    layer3_outputs(1203) <= (layer2_outputs(998)) xor (layer2_outputs(3628));
    layer3_outputs(1204) <= (layer2_outputs(2732)) or (layer2_outputs(4147));
    layer3_outputs(1205) <= (layer2_outputs(2361)) or (layer2_outputs(4357));
    layer3_outputs(1206) <= (layer2_outputs(1922)) and not (layer2_outputs(4545));
    layer3_outputs(1207) <= layer2_outputs(496);
    layer3_outputs(1208) <= '1';
    layer3_outputs(1209) <= not(layer2_outputs(4711)) or (layer2_outputs(4881));
    layer3_outputs(1210) <= layer2_outputs(4057);
    layer3_outputs(1211) <= layer2_outputs(2134);
    layer3_outputs(1212) <= layer2_outputs(3777);
    layer3_outputs(1213) <= (layer2_outputs(445)) and not (layer2_outputs(340));
    layer3_outputs(1214) <= not(layer2_outputs(1805));
    layer3_outputs(1215) <= not((layer2_outputs(242)) or (layer2_outputs(155)));
    layer3_outputs(1216) <= '0';
    layer3_outputs(1217) <= not(layer2_outputs(4747));
    layer3_outputs(1218) <= '1';
    layer3_outputs(1219) <= not(layer2_outputs(3599));
    layer3_outputs(1220) <= not(layer2_outputs(2251));
    layer3_outputs(1221) <= '0';
    layer3_outputs(1222) <= '0';
    layer3_outputs(1223) <= layer2_outputs(2750);
    layer3_outputs(1224) <= '1';
    layer3_outputs(1225) <= '1';
    layer3_outputs(1226) <= not(layer2_outputs(1645)) or (layer2_outputs(4356));
    layer3_outputs(1227) <= not(layer2_outputs(718));
    layer3_outputs(1228) <= (layer2_outputs(2871)) and not (layer2_outputs(4681));
    layer3_outputs(1229) <= '1';
    layer3_outputs(1230) <= (layer2_outputs(2492)) and not (layer2_outputs(2144));
    layer3_outputs(1231) <= '1';
    layer3_outputs(1232) <= '1';
    layer3_outputs(1233) <= not(layer2_outputs(1694)) or (layer2_outputs(3322));
    layer3_outputs(1234) <= not(layer2_outputs(4549));
    layer3_outputs(1235) <= not(layer2_outputs(3152));
    layer3_outputs(1236) <= layer2_outputs(1385);
    layer3_outputs(1237) <= not(layer2_outputs(3256));
    layer3_outputs(1238) <= layer2_outputs(2001);
    layer3_outputs(1239) <= layer2_outputs(2677);
    layer3_outputs(1240) <= '0';
    layer3_outputs(1241) <= not(layer2_outputs(3170));
    layer3_outputs(1242) <= (layer2_outputs(1364)) and not (layer2_outputs(154));
    layer3_outputs(1243) <= layer2_outputs(43);
    layer3_outputs(1244) <= '0';
    layer3_outputs(1245) <= not(layer2_outputs(542)) or (layer2_outputs(177));
    layer3_outputs(1246) <= not(layer2_outputs(797)) or (layer2_outputs(4600));
    layer3_outputs(1247) <= '1';
    layer3_outputs(1248) <= not((layer2_outputs(3694)) or (layer2_outputs(1202)));
    layer3_outputs(1249) <= (layer2_outputs(2810)) and not (layer2_outputs(4726));
    layer3_outputs(1250) <= (layer2_outputs(3998)) and not (layer2_outputs(3282));
    layer3_outputs(1251) <= not(layer2_outputs(4537));
    layer3_outputs(1252) <= (layer2_outputs(346)) and (layer2_outputs(2821));
    layer3_outputs(1253) <= not(layer2_outputs(5117)) or (layer2_outputs(4525));
    layer3_outputs(1254) <= '1';
    layer3_outputs(1255) <= not(layer2_outputs(671));
    layer3_outputs(1256) <= not(layer2_outputs(1298));
    layer3_outputs(1257) <= not(layer2_outputs(1102)) or (layer2_outputs(2887));
    layer3_outputs(1258) <= not((layer2_outputs(4882)) or (layer2_outputs(1280)));
    layer3_outputs(1259) <= layer2_outputs(845);
    layer3_outputs(1260) <= '0';
    layer3_outputs(1261) <= '0';
    layer3_outputs(1262) <= layer2_outputs(1005);
    layer3_outputs(1263) <= not(layer2_outputs(4102));
    layer3_outputs(1264) <= not(layer2_outputs(2881));
    layer3_outputs(1265) <= not(layer2_outputs(4220));
    layer3_outputs(1266) <= layer2_outputs(496);
    layer3_outputs(1267) <= not((layer2_outputs(2272)) or (layer2_outputs(3970)));
    layer3_outputs(1268) <= not(layer2_outputs(1838)) or (layer2_outputs(513));
    layer3_outputs(1269) <= not((layer2_outputs(2485)) or (layer2_outputs(1299)));
    layer3_outputs(1270) <= layer2_outputs(2815);
    layer3_outputs(1271) <= (layer2_outputs(1300)) and (layer2_outputs(3067));
    layer3_outputs(1272) <= not(layer2_outputs(3919));
    layer3_outputs(1273) <= not(layer2_outputs(1282));
    layer3_outputs(1274) <= not(layer2_outputs(4735)) or (layer2_outputs(1189));
    layer3_outputs(1275) <= '1';
    layer3_outputs(1276) <= (layer2_outputs(1117)) and not (layer2_outputs(1680));
    layer3_outputs(1277) <= (layer2_outputs(4193)) and (layer2_outputs(3930));
    layer3_outputs(1278) <= not((layer2_outputs(486)) and (layer2_outputs(1017)));
    layer3_outputs(1279) <= '1';
    layer3_outputs(1280) <= layer2_outputs(3581);
    layer3_outputs(1281) <= layer2_outputs(3822);
    layer3_outputs(1282) <= not(layer2_outputs(1560)) or (layer2_outputs(884));
    layer3_outputs(1283) <= layer2_outputs(557);
    layer3_outputs(1284) <= '1';
    layer3_outputs(1285) <= not(layer2_outputs(3297)) or (layer2_outputs(4783));
    layer3_outputs(1286) <= not(layer2_outputs(1290));
    layer3_outputs(1287) <= (layer2_outputs(32)) or (layer2_outputs(1279));
    layer3_outputs(1288) <= '1';
    layer3_outputs(1289) <= not((layer2_outputs(1026)) or (layer2_outputs(1153)));
    layer3_outputs(1290) <= not(layer2_outputs(5004));
    layer3_outputs(1291) <= layer2_outputs(509);
    layer3_outputs(1292) <= not(layer2_outputs(1640));
    layer3_outputs(1293) <= not(layer2_outputs(4264)) or (layer2_outputs(894));
    layer3_outputs(1294) <= '0';
    layer3_outputs(1295) <= not((layer2_outputs(3767)) and (layer2_outputs(4989)));
    layer3_outputs(1296) <= not(layer2_outputs(2395));
    layer3_outputs(1297) <= '0';
    layer3_outputs(1298) <= not(layer2_outputs(2553));
    layer3_outputs(1299) <= (layer2_outputs(4188)) or (layer2_outputs(2185));
    layer3_outputs(1300) <= (layer2_outputs(3718)) and not (layer2_outputs(3219));
    layer3_outputs(1301) <= (layer2_outputs(1359)) xor (layer2_outputs(2701));
    layer3_outputs(1302) <= layer2_outputs(2887);
    layer3_outputs(1303) <= '0';
    layer3_outputs(1304) <= not(layer2_outputs(2608));
    layer3_outputs(1305) <= (layer2_outputs(3685)) and (layer2_outputs(2424));
    layer3_outputs(1306) <= not(layer2_outputs(1673)) or (layer2_outputs(4490));
    layer3_outputs(1307) <= not(layer2_outputs(1886));
    layer3_outputs(1308) <= layer2_outputs(3198);
    layer3_outputs(1309) <= not(layer2_outputs(2851));
    layer3_outputs(1310) <= not(layer2_outputs(2694)) or (layer2_outputs(2731));
    layer3_outputs(1311) <= (layer2_outputs(209)) and (layer2_outputs(2218));
    layer3_outputs(1312) <= not(layer2_outputs(1922));
    layer3_outputs(1313) <= (layer2_outputs(1681)) and (layer2_outputs(69));
    layer3_outputs(1314) <= layer2_outputs(2001);
    layer3_outputs(1315) <= not((layer2_outputs(4162)) or (layer2_outputs(2687)));
    layer3_outputs(1316) <= (layer2_outputs(2659)) xor (layer2_outputs(2800));
    layer3_outputs(1317) <= (layer2_outputs(1246)) and not (layer2_outputs(3468));
    layer3_outputs(1318) <= not(layer2_outputs(14));
    layer3_outputs(1319) <= layer2_outputs(1752);
    layer3_outputs(1320) <= not(layer2_outputs(2563)) or (layer2_outputs(3856));
    layer3_outputs(1321) <= not(layer2_outputs(4340)) or (layer2_outputs(2401));
    layer3_outputs(1322) <= not(layer2_outputs(364));
    layer3_outputs(1323) <= (layer2_outputs(625)) xor (layer2_outputs(4963));
    layer3_outputs(1324) <= not(layer2_outputs(3095));
    layer3_outputs(1325) <= layer2_outputs(3525);
    layer3_outputs(1326) <= (layer2_outputs(3551)) or (layer2_outputs(1001));
    layer3_outputs(1327) <= not(layer2_outputs(950));
    layer3_outputs(1328) <= not(layer2_outputs(4262));
    layer3_outputs(1329) <= (layer2_outputs(3850)) and not (layer2_outputs(4598));
    layer3_outputs(1330) <= not(layer2_outputs(4842));
    layer3_outputs(1331) <= (layer2_outputs(1552)) and not (layer2_outputs(3420));
    layer3_outputs(1332) <= not(layer2_outputs(1999));
    layer3_outputs(1333) <= (layer2_outputs(2602)) and not (layer2_outputs(3574));
    layer3_outputs(1334) <= layer2_outputs(3618);
    layer3_outputs(1335) <= layer2_outputs(3569);
    layer3_outputs(1336) <= not(layer2_outputs(3454)) or (layer2_outputs(1970));
    layer3_outputs(1337) <= (layer2_outputs(2701)) and not (layer2_outputs(850));
    layer3_outputs(1338) <= layer2_outputs(4071);
    layer3_outputs(1339) <= (layer2_outputs(2529)) xor (layer2_outputs(3189));
    layer3_outputs(1340) <= not(layer2_outputs(4919));
    layer3_outputs(1341) <= not(layer2_outputs(2815));
    layer3_outputs(1342) <= layer2_outputs(2335);
    layer3_outputs(1343) <= '1';
    layer3_outputs(1344) <= layer2_outputs(3283);
    layer3_outputs(1345) <= (layer2_outputs(263)) and not (layer2_outputs(1646));
    layer3_outputs(1346) <= not((layer2_outputs(884)) or (layer2_outputs(3451)));
    layer3_outputs(1347) <= not((layer2_outputs(142)) or (layer2_outputs(3795)));
    layer3_outputs(1348) <= (layer2_outputs(3474)) and not (layer2_outputs(4249));
    layer3_outputs(1349) <= (layer2_outputs(4353)) and not (layer2_outputs(2576));
    layer3_outputs(1350) <= not(layer2_outputs(951)) or (layer2_outputs(3775));
    layer3_outputs(1351) <= (layer2_outputs(2238)) and not (layer2_outputs(1705));
    layer3_outputs(1352) <= (layer2_outputs(4267)) xor (layer2_outputs(4830));
    layer3_outputs(1353) <= '1';
    layer3_outputs(1354) <= not(layer2_outputs(4691));
    layer3_outputs(1355) <= (layer2_outputs(53)) or (layer2_outputs(2009));
    layer3_outputs(1356) <= not(layer2_outputs(2345));
    layer3_outputs(1357) <= '0';
    layer3_outputs(1358) <= layer2_outputs(2184);
    layer3_outputs(1359) <= not(layer2_outputs(4670));
    layer3_outputs(1360) <= not(layer2_outputs(2667)) or (layer2_outputs(936));
    layer3_outputs(1361) <= (layer2_outputs(1707)) and not (layer2_outputs(2733));
    layer3_outputs(1362) <= not(layer2_outputs(3122)) or (layer2_outputs(1343));
    layer3_outputs(1363) <= (layer2_outputs(1849)) xor (layer2_outputs(4383));
    layer3_outputs(1364) <= layer2_outputs(1918);
    layer3_outputs(1365) <= not(layer2_outputs(3917));
    layer3_outputs(1366) <= '0';
    layer3_outputs(1367) <= '0';
    layer3_outputs(1368) <= not(layer2_outputs(4480));
    layer3_outputs(1369) <= not(layer2_outputs(130));
    layer3_outputs(1370) <= (layer2_outputs(4654)) and not (layer2_outputs(3329));
    layer3_outputs(1371) <= not(layer2_outputs(1102));
    layer3_outputs(1372) <= layer2_outputs(3542);
    layer3_outputs(1373) <= not(layer2_outputs(3254));
    layer3_outputs(1374) <= not(layer2_outputs(5086));
    layer3_outputs(1375) <= (layer2_outputs(1100)) and (layer2_outputs(4090));
    layer3_outputs(1376) <= (layer2_outputs(1949)) and not (layer2_outputs(4206));
    layer3_outputs(1377) <= (layer2_outputs(2555)) and not (layer2_outputs(823));
    layer3_outputs(1378) <= (layer2_outputs(992)) and not (layer2_outputs(3221));
    layer3_outputs(1379) <= '1';
    layer3_outputs(1380) <= (layer2_outputs(2883)) and not (layer2_outputs(2356));
    layer3_outputs(1381) <= '0';
    layer3_outputs(1382) <= not(layer2_outputs(839)) or (layer2_outputs(4132));
    layer3_outputs(1383) <= layer2_outputs(845);
    layer3_outputs(1384) <= layer2_outputs(3612);
    layer3_outputs(1385) <= not(layer2_outputs(2558));
    layer3_outputs(1386) <= '1';
    layer3_outputs(1387) <= (layer2_outputs(1004)) and not (layer2_outputs(3852));
    layer3_outputs(1388) <= not((layer2_outputs(410)) and (layer2_outputs(4162)));
    layer3_outputs(1389) <= not(layer2_outputs(1684)) or (layer2_outputs(4319));
    layer3_outputs(1390) <= not(layer2_outputs(488)) or (layer2_outputs(445));
    layer3_outputs(1391) <= not(layer2_outputs(1505)) or (layer2_outputs(5057));
    layer3_outputs(1392) <= (layer2_outputs(978)) xor (layer2_outputs(3570));
    layer3_outputs(1393) <= (layer2_outputs(381)) or (layer2_outputs(4106));
    layer3_outputs(1394) <= (layer2_outputs(2560)) or (layer2_outputs(559));
    layer3_outputs(1395) <= not(layer2_outputs(3853));
    layer3_outputs(1396) <= (layer2_outputs(5117)) or (layer2_outputs(361));
    layer3_outputs(1397) <= not((layer2_outputs(3226)) or (layer2_outputs(1092)));
    layer3_outputs(1398) <= layer2_outputs(1039);
    layer3_outputs(1399) <= not(layer2_outputs(344)) or (layer2_outputs(3469));
    layer3_outputs(1400) <= (layer2_outputs(4140)) and not (layer2_outputs(3284));
    layer3_outputs(1401) <= layer2_outputs(2872);
    layer3_outputs(1402) <= layer2_outputs(3535);
    layer3_outputs(1403) <= not(layer2_outputs(2864)) or (layer2_outputs(3011));
    layer3_outputs(1404) <= layer2_outputs(1566);
    layer3_outputs(1405) <= (layer2_outputs(357)) and not (layer2_outputs(3215));
    layer3_outputs(1406) <= layer2_outputs(358);
    layer3_outputs(1407) <= (layer2_outputs(2785)) or (layer2_outputs(658));
    layer3_outputs(1408) <= not(layer2_outputs(2629));
    layer3_outputs(1409) <= not(layer2_outputs(766));
    layer3_outputs(1410) <= not((layer2_outputs(1534)) or (layer2_outputs(1875)));
    layer3_outputs(1411) <= (layer2_outputs(1406)) or (layer2_outputs(378));
    layer3_outputs(1412) <= (layer2_outputs(1711)) and (layer2_outputs(4651));
    layer3_outputs(1413) <= not(layer2_outputs(885)) or (layer2_outputs(4326));
    layer3_outputs(1414) <= '0';
    layer3_outputs(1415) <= layer2_outputs(3047);
    layer3_outputs(1416) <= not(layer2_outputs(286));
    layer3_outputs(1417) <= (layer2_outputs(28)) and (layer2_outputs(3494));
    layer3_outputs(1418) <= '1';
    layer3_outputs(1419) <= (layer2_outputs(2538)) and not (layer2_outputs(3268));
    layer3_outputs(1420) <= '1';
    layer3_outputs(1421) <= (layer2_outputs(1984)) and (layer2_outputs(3475));
    layer3_outputs(1422) <= '0';
    layer3_outputs(1423) <= layer2_outputs(3643);
    layer3_outputs(1424) <= not(layer2_outputs(1671)) or (layer2_outputs(139));
    layer3_outputs(1425) <= layer2_outputs(4159);
    layer3_outputs(1426) <= not(layer2_outputs(3086));
    layer3_outputs(1427) <= layer2_outputs(3135);
    layer3_outputs(1428) <= layer2_outputs(1365);
    layer3_outputs(1429) <= '0';
    layer3_outputs(1430) <= not(layer2_outputs(4001)) or (layer2_outputs(3553));
    layer3_outputs(1431) <= '0';
    layer3_outputs(1432) <= (layer2_outputs(2030)) and not (layer2_outputs(4678));
    layer3_outputs(1433) <= '1';
    layer3_outputs(1434) <= layer2_outputs(1121);
    layer3_outputs(1435) <= not((layer2_outputs(3333)) or (layer2_outputs(2236)));
    layer3_outputs(1436) <= not(layer2_outputs(622));
    layer3_outputs(1437) <= not(layer2_outputs(1742));
    layer3_outputs(1438) <= layer2_outputs(3146);
    layer3_outputs(1439) <= (layer2_outputs(1962)) and not (layer2_outputs(1894));
    layer3_outputs(1440) <= not(layer2_outputs(2097));
    layer3_outputs(1441) <= not((layer2_outputs(1883)) xor (layer2_outputs(3884)));
    layer3_outputs(1442) <= not(layer2_outputs(1607)) or (layer2_outputs(2573));
    layer3_outputs(1443) <= '1';
    layer3_outputs(1444) <= not(layer2_outputs(4253));
    layer3_outputs(1445) <= not(layer2_outputs(2014));
    layer3_outputs(1446) <= not(layer2_outputs(1500));
    layer3_outputs(1447) <= (layer2_outputs(3720)) or (layer2_outputs(112));
    layer3_outputs(1448) <= (layer2_outputs(1719)) and (layer2_outputs(1753));
    layer3_outputs(1449) <= not((layer2_outputs(5090)) or (layer2_outputs(4853)));
    layer3_outputs(1450) <= layer2_outputs(1015);
    layer3_outputs(1451) <= (layer2_outputs(1443)) or (layer2_outputs(2593));
    layer3_outputs(1452) <= not((layer2_outputs(3628)) and (layer2_outputs(1986)));
    layer3_outputs(1453) <= (layer2_outputs(2263)) or (layer2_outputs(1523));
    layer3_outputs(1454) <= not((layer2_outputs(2797)) or (layer2_outputs(452)));
    layer3_outputs(1455) <= not((layer2_outputs(5082)) or (layer2_outputs(4253)));
    layer3_outputs(1456) <= not(layer2_outputs(1040)) or (layer2_outputs(2267));
    layer3_outputs(1457) <= not(layer2_outputs(2032));
    layer3_outputs(1458) <= not((layer2_outputs(1438)) and (layer2_outputs(4554)));
    layer3_outputs(1459) <= (layer2_outputs(4708)) or (layer2_outputs(400));
    layer3_outputs(1460) <= '0';
    layer3_outputs(1461) <= (layer2_outputs(1179)) and not (layer2_outputs(2062));
    layer3_outputs(1462) <= not((layer2_outputs(2040)) and (layer2_outputs(4143)));
    layer3_outputs(1463) <= (layer2_outputs(1030)) and (layer2_outputs(710));
    layer3_outputs(1464) <= not(layer2_outputs(4464)) or (layer2_outputs(4351));
    layer3_outputs(1465) <= (layer2_outputs(3327)) and (layer2_outputs(5094));
    layer3_outputs(1466) <= not(layer2_outputs(1205));
    layer3_outputs(1467) <= (layer2_outputs(2216)) and not (layer2_outputs(4917));
    layer3_outputs(1468) <= '1';
    layer3_outputs(1469) <= not(layer2_outputs(3613));
    layer3_outputs(1470) <= '0';
    layer3_outputs(1471) <= (layer2_outputs(1996)) and (layer2_outputs(2102));
    layer3_outputs(1472) <= (layer2_outputs(1148)) and not (layer2_outputs(458));
    layer3_outputs(1473) <= not(layer2_outputs(4059));
    layer3_outputs(1474) <= layer2_outputs(1315);
    layer3_outputs(1475) <= layer2_outputs(2343);
    layer3_outputs(1476) <= not(layer2_outputs(432)) or (layer2_outputs(4877));
    layer3_outputs(1477) <= layer2_outputs(56);
    layer3_outputs(1478) <= layer2_outputs(4020);
    layer3_outputs(1479) <= layer2_outputs(1532);
    layer3_outputs(1480) <= '1';
    layer3_outputs(1481) <= not((layer2_outputs(3906)) or (layer2_outputs(4128)));
    layer3_outputs(1482) <= not(layer2_outputs(2147));
    layer3_outputs(1483) <= not(layer2_outputs(3622)) or (layer2_outputs(210));
    layer3_outputs(1484) <= (layer2_outputs(4856)) and (layer2_outputs(4695));
    layer3_outputs(1485) <= (layer2_outputs(3395)) xor (layer2_outputs(5079));
    layer3_outputs(1486) <= (layer2_outputs(4721)) and (layer2_outputs(3886));
    layer3_outputs(1487) <= not((layer2_outputs(2611)) and (layer2_outputs(1752)));
    layer3_outputs(1488) <= layer2_outputs(4258);
    layer3_outputs(1489) <= not(layer2_outputs(1332));
    layer3_outputs(1490) <= (layer2_outputs(4097)) or (layer2_outputs(5051));
    layer3_outputs(1491) <= '0';
    layer3_outputs(1492) <= (layer2_outputs(1009)) and not (layer2_outputs(3812));
    layer3_outputs(1493) <= '1';
    layer3_outputs(1494) <= not(layer2_outputs(60));
    layer3_outputs(1495) <= not(layer2_outputs(4743));
    layer3_outputs(1496) <= layer2_outputs(3218);
    layer3_outputs(1497) <= '0';
    layer3_outputs(1498) <= '1';
    layer3_outputs(1499) <= not(layer2_outputs(1342)) or (layer2_outputs(2262));
    layer3_outputs(1500) <= (layer2_outputs(2141)) and not (layer2_outputs(4061));
    layer3_outputs(1501) <= (layer2_outputs(3220)) and (layer2_outputs(370));
    layer3_outputs(1502) <= not((layer2_outputs(4723)) and (layer2_outputs(926)));
    layer3_outputs(1503) <= not((layer2_outputs(2832)) and (layer2_outputs(4788)));
    layer3_outputs(1504) <= not((layer2_outputs(1468)) and (layer2_outputs(1672)));
    layer3_outputs(1505) <= layer2_outputs(2386);
    layer3_outputs(1506) <= (layer2_outputs(1791)) and (layer2_outputs(1040));
    layer3_outputs(1507) <= layer2_outputs(626);
    layer3_outputs(1508) <= layer2_outputs(3669);
    layer3_outputs(1509) <= '1';
    layer3_outputs(1510) <= (layer2_outputs(909)) and (layer2_outputs(4661));
    layer3_outputs(1511) <= layer2_outputs(394);
    layer3_outputs(1512) <= layer2_outputs(3844);
    layer3_outputs(1513) <= not((layer2_outputs(3723)) or (layer2_outputs(4924)));
    layer3_outputs(1514) <= '1';
    layer3_outputs(1515) <= (layer2_outputs(3390)) and not (layer2_outputs(2482));
    layer3_outputs(1516) <= (layer2_outputs(1946)) and not (layer2_outputs(3441));
    layer3_outputs(1517) <= layer2_outputs(584);
    layer3_outputs(1518) <= not(layer2_outputs(5031));
    layer3_outputs(1519) <= layer2_outputs(2894);
    layer3_outputs(1520) <= '0';
    layer3_outputs(1521) <= layer2_outputs(3480);
    layer3_outputs(1522) <= layer2_outputs(1046);
    layer3_outputs(1523) <= (layer2_outputs(617)) or (layer2_outputs(2033));
    layer3_outputs(1524) <= (layer2_outputs(1431)) and not (layer2_outputs(476));
    layer3_outputs(1525) <= not((layer2_outputs(3787)) or (layer2_outputs(632)));
    layer3_outputs(1526) <= (layer2_outputs(925)) and not (layer2_outputs(3348));
    layer3_outputs(1527) <= (layer2_outputs(414)) and not (layer2_outputs(4441));
    layer3_outputs(1528) <= (layer2_outputs(4703)) and (layer2_outputs(1919));
    layer3_outputs(1529) <= not(layer2_outputs(4408));
    layer3_outputs(1530) <= (layer2_outputs(2995)) and (layer2_outputs(2325));
    layer3_outputs(1531) <= not(layer2_outputs(4959));
    layer3_outputs(1532) <= (layer2_outputs(1419)) and (layer2_outputs(1711));
    layer3_outputs(1533) <= (layer2_outputs(685)) or (layer2_outputs(6));
    layer3_outputs(1534) <= not(layer2_outputs(4008));
    layer3_outputs(1535) <= not(layer2_outputs(2280));
    layer3_outputs(1536) <= (layer2_outputs(2705)) or (layer2_outputs(858));
    layer3_outputs(1537) <= (layer2_outputs(251)) and not (layer2_outputs(2411));
    layer3_outputs(1538) <= not(layer2_outputs(1955)) or (layer2_outputs(145));
    layer3_outputs(1539) <= (layer2_outputs(454)) and (layer2_outputs(3207));
    layer3_outputs(1540) <= (layer2_outputs(661)) and not (layer2_outputs(3979));
    layer3_outputs(1541) <= (layer2_outputs(2000)) and not (layer2_outputs(4742));
    layer3_outputs(1542) <= not(layer2_outputs(2205));
    layer3_outputs(1543) <= '0';
    layer3_outputs(1544) <= (layer2_outputs(719)) or (layer2_outputs(2544));
    layer3_outputs(1545) <= not(layer2_outputs(544));
    layer3_outputs(1546) <= not((layer2_outputs(262)) or (layer2_outputs(3031)));
    layer3_outputs(1547) <= '1';
    layer3_outputs(1548) <= layer2_outputs(2168);
    layer3_outputs(1549) <= not(layer2_outputs(583));
    layer3_outputs(1550) <= layer2_outputs(4714);
    layer3_outputs(1551) <= not(layer2_outputs(2391)) or (layer2_outputs(5100));
    layer3_outputs(1552) <= not(layer2_outputs(3131)) or (layer2_outputs(4225));
    layer3_outputs(1553) <= (layer2_outputs(159)) and not (layer2_outputs(3946));
    layer3_outputs(1554) <= (layer2_outputs(4565)) or (layer2_outputs(1076));
    layer3_outputs(1555) <= not(layer2_outputs(2384));
    layer3_outputs(1556) <= not(layer2_outputs(3033));
    layer3_outputs(1557) <= not(layer2_outputs(4381));
    layer3_outputs(1558) <= not(layer2_outputs(4746));
    layer3_outputs(1559) <= '0';
    layer3_outputs(1560) <= layer2_outputs(2456);
    layer3_outputs(1561) <= layer2_outputs(468);
    layer3_outputs(1562) <= not((layer2_outputs(1529)) and (layer2_outputs(3712)));
    layer3_outputs(1563) <= '1';
    layer3_outputs(1564) <= (layer2_outputs(4017)) and not (layer2_outputs(1416));
    layer3_outputs(1565) <= (layer2_outputs(4740)) and (layer2_outputs(2943));
    layer3_outputs(1566) <= layer2_outputs(1649);
    layer3_outputs(1567) <= (layer2_outputs(3387)) and not (layer2_outputs(3478));
    layer3_outputs(1568) <= not(layer2_outputs(2068));
    layer3_outputs(1569) <= (layer2_outputs(3833)) xor (layer2_outputs(4816));
    layer3_outputs(1570) <= not(layer2_outputs(8));
    layer3_outputs(1571) <= '1';
    layer3_outputs(1572) <= not((layer2_outputs(4853)) and (layer2_outputs(1077)));
    layer3_outputs(1573) <= not(layer2_outputs(3055)) or (layer2_outputs(772));
    layer3_outputs(1574) <= layer2_outputs(1658);
    layer3_outputs(1575) <= not(layer2_outputs(4194)) or (layer2_outputs(1864));
    layer3_outputs(1576) <= (layer2_outputs(2657)) and not (layer2_outputs(3400));
    layer3_outputs(1577) <= not(layer2_outputs(456)) or (layer2_outputs(3793));
    layer3_outputs(1578) <= (layer2_outputs(747)) and (layer2_outputs(2254));
    layer3_outputs(1579) <= not((layer2_outputs(90)) or (layer2_outputs(506)));
    layer3_outputs(1580) <= not((layer2_outputs(4677)) or (layer2_outputs(3129)));
    layer3_outputs(1581) <= '0';
    layer3_outputs(1582) <= not(layer2_outputs(846)) or (layer2_outputs(2445));
    layer3_outputs(1583) <= layer2_outputs(4095);
    layer3_outputs(1584) <= not(layer2_outputs(1175));
    layer3_outputs(1585) <= (layer2_outputs(4585)) or (layer2_outputs(1779));
    layer3_outputs(1586) <= not(layer2_outputs(1886));
    layer3_outputs(1587) <= not(layer2_outputs(4233));
    layer3_outputs(1588) <= not(layer2_outputs(4725)) or (layer2_outputs(1816));
    layer3_outputs(1589) <= (layer2_outputs(2953)) and not (layer2_outputs(4275));
    layer3_outputs(1590) <= (layer2_outputs(3482)) or (layer2_outputs(2314));
    layer3_outputs(1591) <= '0';
    layer3_outputs(1592) <= (layer2_outputs(2438)) and (layer2_outputs(785));
    layer3_outputs(1593) <= '1';
    layer3_outputs(1594) <= not(layer2_outputs(758)) or (layer2_outputs(2241));
    layer3_outputs(1595) <= not(layer2_outputs(3301));
    layer3_outputs(1596) <= '1';
    layer3_outputs(1597) <= not(layer2_outputs(203));
    layer3_outputs(1598) <= layer2_outputs(2658);
    layer3_outputs(1599) <= not(layer2_outputs(4222)) or (layer2_outputs(4344));
    layer3_outputs(1600) <= layer2_outputs(220);
    layer3_outputs(1601) <= not(layer2_outputs(4208)) or (layer2_outputs(1336));
    layer3_outputs(1602) <= not(layer2_outputs(1492)) or (layer2_outputs(2541));
    layer3_outputs(1603) <= not(layer2_outputs(2404));
    layer3_outputs(1604) <= layer2_outputs(2961);
    layer3_outputs(1605) <= (layer2_outputs(1016)) and not (layer2_outputs(3562));
    layer3_outputs(1606) <= (layer2_outputs(2805)) and not (layer2_outputs(2957));
    layer3_outputs(1607) <= layer2_outputs(3545);
    layer3_outputs(1608) <= not(layer2_outputs(5057)) or (layer2_outputs(1175));
    layer3_outputs(1609) <= (layer2_outputs(691)) or (layer2_outputs(4259));
    layer3_outputs(1610) <= not(layer2_outputs(4329));
    layer3_outputs(1611) <= not(layer2_outputs(55)) or (layer2_outputs(275));
    layer3_outputs(1612) <= not(layer2_outputs(717)) or (layer2_outputs(2466));
    layer3_outputs(1613) <= (layer2_outputs(729)) and not (layer2_outputs(3897));
    layer3_outputs(1614) <= layer2_outputs(1572);
    layer3_outputs(1615) <= (layer2_outputs(4588)) and not (layer2_outputs(4070));
    layer3_outputs(1616) <= layer2_outputs(2051);
    layer3_outputs(1617) <= layer2_outputs(3917);
    layer3_outputs(1618) <= (layer2_outputs(3421)) and not (layer2_outputs(9));
    layer3_outputs(1619) <= not(layer2_outputs(1892));
    layer3_outputs(1620) <= (layer2_outputs(3396)) and (layer2_outputs(1044));
    layer3_outputs(1621) <= (layer2_outputs(2845)) and not (layer2_outputs(2500));
    layer3_outputs(1622) <= not((layer2_outputs(4610)) or (layer2_outputs(1561)));
    layer3_outputs(1623) <= not(layer2_outputs(4171)) or (layer2_outputs(131));
    layer3_outputs(1624) <= layer2_outputs(3258);
    layer3_outputs(1625) <= not((layer2_outputs(2909)) and (layer2_outputs(303)));
    layer3_outputs(1626) <= not(layer2_outputs(3490));
    layer3_outputs(1627) <= not((layer2_outputs(1402)) and (layer2_outputs(691)));
    layer3_outputs(1628) <= (layer2_outputs(2049)) or (layer2_outputs(4168));
    layer3_outputs(1629) <= not(layer2_outputs(3940)) or (layer2_outputs(2649));
    layer3_outputs(1630) <= not(layer2_outputs(535));
    layer3_outputs(1631) <= (layer2_outputs(2399)) xor (layer2_outputs(3260));
    layer3_outputs(1632) <= (layer2_outputs(2383)) or (layer2_outputs(4592));
    layer3_outputs(1633) <= not(layer2_outputs(4694)) or (layer2_outputs(4868));
    layer3_outputs(1634) <= not((layer2_outputs(1643)) or (layer2_outputs(292)));
    layer3_outputs(1635) <= layer2_outputs(1273);
    layer3_outputs(1636) <= layer2_outputs(336);
    layer3_outputs(1637) <= (layer2_outputs(3610)) and not (layer2_outputs(2095));
    layer3_outputs(1638) <= layer2_outputs(3263);
    layer3_outputs(1639) <= not(layer2_outputs(1786)) or (layer2_outputs(4676));
    layer3_outputs(1640) <= (layer2_outputs(4030)) xor (layer2_outputs(4077));
    layer3_outputs(1641) <= layer2_outputs(2535);
    layer3_outputs(1642) <= not(layer2_outputs(916));
    layer3_outputs(1643) <= not((layer2_outputs(497)) and (layer2_outputs(4729)));
    layer3_outputs(1644) <= not((layer2_outputs(3624)) and (layer2_outputs(2433)));
    layer3_outputs(1645) <= not(layer2_outputs(480));
    layer3_outputs(1646) <= '1';
    layer3_outputs(1647) <= not(layer2_outputs(4655));
    layer3_outputs(1648) <= not(layer2_outputs(3079));
    layer3_outputs(1649) <= not(layer2_outputs(1555));
    layer3_outputs(1650) <= layer2_outputs(436);
    layer3_outputs(1651) <= '0';
    layer3_outputs(1652) <= (layer2_outputs(5039)) and (layer2_outputs(318));
    layer3_outputs(1653) <= not((layer2_outputs(516)) and (layer2_outputs(3695)));
    layer3_outputs(1654) <= not((layer2_outputs(4888)) and (layer2_outputs(4436)));
    layer3_outputs(1655) <= not((layer2_outputs(493)) and (layer2_outputs(4937)));
    layer3_outputs(1656) <= not(layer2_outputs(4498));
    layer3_outputs(1657) <= (layer2_outputs(2703)) or (layer2_outputs(3187));
    layer3_outputs(1658) <= not((layer2_outputs(791)) or (layer2_outputs(5105)));
    layer3_outputs(1659) <= not((layer2_outputs(3898)) or (layer2_outputs(1730)));
    layer3_outputs(1660) <= layer2_outputs(4912);
    layer3_outputs(1661) <= (layer2_outputs(5006)) and (layer2_outputs(2745));
    layer3_outputs(1662) <= not(layer2_outputs(714));
    layer3_outputs(1663) <= not(layer2_outputs(4270));
    layer3_outputs(1664) <= (layer2_outputs(3390)) and not (layer2_outputs(3506));
    layer3_outputs(1665) <= '0';
    layer3_outputs(1666) <= not((layer2_outputs(3270)) or (layer2_outputs(807)));
    layer3_outputs(1667) <= not((layer2_outputs(269)) or (layer2_outputs(1917)));
    layer3_outputs(1668) <= not(layer2_outputs(1439));
    layer3_outputs(1669) <= not((layer2_outputs(606)) and (layer2_outputs(3173)));
    layer3_outputs(1670) <= not(layer2_outputs(3785)) or (layer2_outputs(3559));
    layer3_outputs(1671) <= (layer2_outputs(4783)) or (layer2_outputs(163));
    layer3_outputs(1672) <= layer2_outputs(871);
    layer3_outputs(1673) <= not(layer2_outputs(1135));
    layer3_outputs(1674) <= '0';
    layer3_outputs(1675) <= not((layer2_outputs(457)) and (layer2_outputs(4968)));
    layer3_outputs(1676) <= '0';
    layer3_outputs(1677) <= (layer2_outputs(3644)) and not (layer2_outputs(4926));
    layer3_outputs(1678) <= '1';
    layer3_outputs(1679) <= (layer2_outputs(380)) xor (layer2_outputs(2480));
    layer3_outputs(1680) <= layer2_outputs(4180);
    layer3_outputs(1681) <= (layer2_outputs(752)) and not (layer2_outputs(4308));
    layer3_outputs(1682) <= layer2_outputs(314);
    layer3_outputs(1683) <= '1';
    layer3_outputs(1684) <= not(layer2_outputs(2364));
    layer3_outputs(1685) <= not(layer2_outputs(667)) or (layer2_outputs(4718));
    layer3_outputs(1686) <= '1';
    layer3_outputs(1687) <= '0';
    layer3_outputs(1688) <= layer2_outputs(3012);
    layer3_outputs(1689) <= layer2_outputs(2393);
    layer3_outputs(1690) <= not(layer2_outputs(5013));
    layer3_outputs(1691) <= (layer2_outputs(1027)) and not (layer2_outputs(1114));
    layer3_outputs(1692) <= not((layer2_outputs(4995)) and (layer2_outputs(272)));
    layer3_outputs(1693) <= not(layer2_outputs(362));
    layer3_outputs(1694) <= layer2_outputs(2897);
    layer3_outputs(1695) <= (layer2_outputs(4574)) and not (layer2_outputs(2972));
    layer3_outputs(1696) <= (layer2_outputs(4439)) and not (layer2_outputs(1805));
    layer3_outputs(1697) <= not(layer2_outputs(3729));
    layer3_outputs(1698) <= (layer2_outputs(3109)) and not (layer2_outputs(2689));
    layer3_outputs(1699) <= '1';
    layer3_outputs(1700) <= (layer2_outputs(2858)) xor (layer2_outputs(2889));
    layer3_outputs(1701) <= (layer2_outputs(1961)) and (layer2_outputs(4686));
    layer3_outputs(1702) <= '0';
    layer3_outputs(1703) <= layer2_outputs(2810);
    layer3_outputs(1704) <= (layer2_outputs(929)) and not (layer2_outputs(86));
    layer3_outputs(1705) <= not(layer2_outputs(982));
    layer3_outputs(1706) <= (layer2_outputs(619)) or (layer2_outputs(3096));
    layer3_outputs(1707) <= not(layer2_outputs(269));
    layer3_outputs(1708) <= (layer2_outputs(1331)) or (layer2_outputs(1304));
    layer3_outputs(1709) <= '1';
    layer3_outputs(1710) <= not(layer2_outputs(4305)) or (layer2_outputs(4987));
    layer3_outputs(1711) <= layer2_outputs(2102);
    layer3_outputs(1712) <= (layer2_outputs(1853)) or (layer2_outputs(483));
    layer3_outputs(1713) <= not(layer2_outputs(4103));
    layer3_outputs(1714) <= (layer2_outputs(3835)) or (layer2_outputs(366));
    layer3_outputs(1715) <= not((layer2_outputs(1060)) or (layer2_outputs(3253)));
    layer3_outputs(1716) <= not(layer2_outputs(1912));
    layer3_outputs(1717) <= not(layer2_outputs(3616)) or (layer2_outputs(3046));
    layer3_outputs(1718) <= (layer2_outputs(4934)) and not (layer2_outputs(4870));
    layer3_outputs(1719) <= (layer2_outputs(4428)) xor (layer2_outputs(3756));
    layer3_outputs(1720) <= layer2_outputs(1851);
    layer3_outputs(1721) <= (layer2_outputs(5105)) and not (layer2_outputs(1739));
    layer3_outputs(1722) <= (layer2_outputs(1266)) and not (layer2_outputs(2169));
    layer3_outputs(1723) <= not((layer2_outputs(265)) or (layer2_outputs(3063)));
    layer3_outputs(1724) <= not(layer2_outputs(3618));
    layer3_outputs(1725) <= (layer2_outputs(3393)) and not (layer2_outputs(391));
    layer3_outputs(1726) <= layer2_outputs(4332);
    layer3_outputs(1727) <= (layer2_outputs(892)) and (layer2_outputs(4292));
    layer3_outputs(1728) <= not(layer2_outputs(777));
    layer3_outputs(1729) <= not(layer2_outputs(2639));
    layer3_outputs(1730) <= layer2_outputs(1692);
    layer3_outputs(1731) <= not(layer2_outputs(3135)) or (layer2_outputs(2172));
    layer3_outputs(1732) <= layer2_outputs(4177);
    layer3_outputs(1733) <= not(layer2_outputs(4798)) or (layer2_outputs(2388));
    layer3_outputs(1734) <= (layer2_outputs(3558)) or (layer2_outputs(362));
    layer3_outputs(1735) <= not((layer2_outputs(370)) xor (layer2_outputs(1060)));
    layer3_outputs(1736) <= not(layer2_outputs(2947));
    layer3_outputs(1737) <= '0';
    layer3_outputs(1738) <= (layer2_outputs(1221)) and not (layer2_outputs(213));
    layer3_outputs(1739) <= not(layer2_outputs(787));
    layer3_outputs(1740) <= layer2_outputs(3311);
    layer3_outputs(1741) <= layer2_outputs(2779);
    layer3_outputs(1742) <= not(layer2_outputs(4342)) or (layer2_outputs(5026));
    layer3_outputs(1743) <= not(layer2_outputs(186)) or (layer2_outputs(3496));
    layer3_outputs(1744) <= not(layer2_outputs(3595));
    layer3_outputs(1745) <= not(layer2_outputs(736));
    layer3_outputs(1746) <= not(layer2_outputs(2798));
    layer3_outputs(1747) <= (layer2_outputs(1005)) and not (layer2_outputs(1119));
    layer3_outputs(1748) <= (layer2_outputs(39)) and (layer2_outputs(3055));
    layer3_outputs(1749) <= not(layer2_outputs(2416));
    layer3_outputs(1750) <= (layer2_outputs(816)) and not (layer2_outputs(1913));
    layer3_outputs(1751) <= not(layer2_outputs(2115)) or (layer2_outputs(4279));
    layer3_outputs(1752) <= not((layer2_outputs(1708)) and (layer2_outputs(1236)));
    layer3_outputs(1753) <= layer2_outputs(3596);
    layer3_outputs(1754) <= not(layer2_outputs(5091));
    layer3_outputs(1755) <= layer2_outputs(5020);
    layer3_outputs(1756) <= not(layer2_outputs(1794)) or (layer2_outputs(279));
    layer3_outputs(1757) <= layer2_outputs(4721);
    layer3_outputs(1758) <= (layer2_outputs(2870)) or (layer2_outputs(460));
    layer3_outputs(1759) <= layer2_outputs(220);
    layer3_outputs(1760) <= not(layer2_outputs(3537));
    layer3_outputs(1761) <= layer2_outputs(3269);
    layer3_outputs(1762) <= '1';
    layer3_outputs(1763) <= '1';
    layer3_outputs(1764) <= '0';
    layer3_outputs(1765) <= layer2_outputs(317);
    layer3_outputs(1766) <= not(layer2_outputs(4631));
    layer3_outputs(1767) <= not((layer2_outputs(2461)) xor (layer2_outputs(797)));
    layer3_outputs(1768) <= not((layer2_outputs(4457)) or (layer2_outputs(2006)));
    layer3_outputs(1769) <= not((layer2_outputs(2651)) and (layer2_outputs(509)));
    layer3_outputs(1770) <= (layer2_outputs(2106)) or (layer2_outputs(6));
    layer3_outputs(1771) <= '1';
    layer3_outputs(1772) <= not(layer2_outputs(647));
    layer3_outputs(1773) <= not((layer2_outputs(2949)) or (layer2_outputs(1510)));
    layer3_outputs(1774) <= '1';
    layer3_outputs(1775) <= (layer2_outputs(2524)) and not (layer2_outputs(2390));
    layer3_outputs(1776) <= not(layer2_outputs(2711)) or (layer2_outputs(1138));
    layer3_outputs(1777) <= not(layer2_outputs(3470)) or (layer2_outputs(86));
    layer3_outputs(1778) <= (layer2_outputs(788)) and not (layer2_outputs(5065));
    layer3_outputs(1779) <= not(layer2_outputs(2478)) or (layer2_outputs(1399));
    layer3_outputs(1780) <= not(layer2_outputs(4928));
    layer3_outputs(1781) <= layer2_outputs(2405);
    layer3_outputs(1782) <= (layer2_outputs(4444)) and not (layer2_outputs(4746));
    layer3_outputs(1783) <= (layer2_outputs(741)) and (layer2_outputs(1716));
    layer3_outputs(1784) <= '1';
    layer3_outputs(1785) <= not(layer2_outputs(3180));
    layer3_outputs(1786) <= not(layer2_outputs(82));
    layer3_outputs(1787) <= layer2_outputs(522);
    layer3_outputs(1788) <= (layer2_outputs(2044)) and not (layer2_outputs(3533));
    layer3_outputs(1789) <= (layer2_outputs(4517)) xor (layer2_outputs(2785));
    layer3_outputs(1790) <= layer2_outputs(2670);
    layer3_outputs(1791) <= '1';
    layer3_outputs(1792) <= (layer2_outputs(3213)) and not (layer2_outputs(1425));
    layer3_outputs(1793) <= not((layer2_outputs(62)) or (layer2_outputs(4078)));
    layer3_outputs(1794) <= not(layer2_outputs(1077));
    layer3_outputs(1795) <= layer2_outputs(1928);
    layer3_outputs(1796) <= (layer2_outputs(2433)) or (layer2_outputs(932));
    layer3_outputs(1797) <= (layer2_outputs(2005)) and not (layer2_outputs(928));
    layer3_outputs(1798) <= not((layer2_outputs(2305)) and (layer2_outputs(4014)));
    layer3_outputs(1799) <= '1';
    layer3_outputs(1800) <= layer2_outputs(1491);
    layer3_outputs(1801) <= not(layer2_outputs(1319));
    layer3_outputs(1802) <= not(layer2_outputs(1002)) or (layer2_outputs(1356));
    layer3_outputs(1803) <= layer2_outputs(2069);
    layer3_outputs(1804) <= not((layer2_outputs(4045)) xor (layer2_outputs(1818)));
    layer3_outputs(1805) <= layer2_outputs(3841);
    layer3_outputs(1806) <= not(layer2_outputs(3049));
    layer3_outputs(1807) <= not((layer2_outputs(1736)) and (layer2_outputs(4869)));
    layer3_outputs(1808) <= not(layer2_outputs(2817));
    layer3_outputs(1809) <= not((layer2_outputs(3857)) or (layer2_outputs(4891)));
    layer3_outputs(1810) <= (layer2_outputs(324)) and (layer2_outputs(3281));
    layer3_outputs(1811) <= (layer2_outputs(3007)) and not (layer2_outputs(658));
    layer3_outputs(1812) <= (layer2_outputs(4336)) or (layer2_outputs(4391));
    layer3_outputs(1813) <= (layer2_outputs(2896)) and not (layer2_outputs(4581));
    layer3_outputs(1814) <= not((layer2_outputs(4208)) xor (layer2_outputs(369)));
    layer3_outputs(1815) <= not(layer2_outputs(2956));
    layer3_outputs(1816) <= not(layer2_outputs(3255));
    layer3_outputs(1817) <= not(layer2_outputs(4861));
    layer3_outputs(1818) <= (layer2_outputs(461)) and (layer2_outputs(4466));
    layer3_outputs(1819) <= not(layer2_outputs(4261)) or (layer2_outputs(1057));
    layer3_outputs(1820) <= not(layer2_outputs(589));
    layer3_outputs(1821) <= layer2_outputs(4956);
    layer3_outputs(1822) <= not(layer2_outputs(2950)) or (layer2_outputs(3398));
    layer3_outputs(1823) <= not(layer2_outputs(4027));
    layer3_outputs(1824) <= (layer2_outputs(4515)) and not (layer2_outputs(3925));
    layer3_outputs(1825) <= not((layer2_outputs(2314)) or (layer2_outputs(708)));
    layer3_outputs(1826) <= not(layer2_outputs(3787)) or (layer2_outputs(4170));
    layer3_outputs(1827) <= (layer2_outputs(37)) xor (layer2_outputs(1768));
    layer3_outputs(1828) <= not((layer2_outputs(3200)) or (layer2_outputs(3279)));
    layer3_outputs(1829) <= (layer2_outputs(4974)) xor (layer2_outputs(3466));
    layer3_outputs(1830) <= layer2_outputs(4273);
    layer3_outputs(1831) <= layer2_outputs(3510);
    layer3_outputs(1832) <= layer2_outputs(4494);
    layer3_outputs(1833) <= (layer2_outputs(2752)) and (layer2_outputs(2907));
    layer3_outputs(1834) <= '1';
    layer3_outputs(1835) <= not(layer2_outputs(3881)) or (layer2_outputs(4107));
    layer3_outputs(1836) <= (layer2_outputs(3411)) and not (layer2_outputs(2792));
    layer3_outputs(1837) <= layer2_outputs(2929);
    layer3_outputs(1838) <= not((layer2_outputs(4666)) and (layer2_outputs(3563)));
    layer3_outputs(1839) <= '1';
    layer3_outputs(1840) <= layer2_outputs(896);
    layer3_outputs(1841) <= layer2_outputs(933);
    layer3_outputs(1842) <= not((layer2_outputs(1689)) xor (layer2_outputs(2828)));
    layer3_outputs(1843) <= not((layer2_outputs(2244)) or (layer2_outputs(4048)));
    layer3_outputs(1844) <= '0';
    layer3_outputs(1845) <= layer2_outputs(4104);
    layer3_outputs(1846) <= (layer2_outputs(3625)) or (layer2_outputs(3715));
    layer3_outputs(1847) <= not(layer2_outputs(2836));
    layer3_outputs(1848) <= not(layer2_outputs(2436));
    layer3_outputs(1849) <= not(layer2_outputs(676));
    layer3_outputs(1850) <= '0';
    layer3_outputs(1851) <= (layer2_outputs(4944)) or (layer2_outputs(1390));
    layer3_outputs(1852) <= not(layer2_outputs(3250));
    layer3_outputs(1853) <= not(layer2_outputs(1436));
    layer3_outputs(1854) <= not(layer2_outputs(4873));
    layer3_outputs(1855) <= not(layer2_outputs(2435));
    layer3_outputs(1856) <= not(layer2_outputs(3761));
    layer3_outputs(1857) <= not(layer2_outputs(4291));
    layer3_outputs(1858) <= (layer2_outputs(1474)) and not (layer2_outputs(2296));
    layer3_outputs(1859) <= not((layer2_outputs(2050)) and (layer2_outputs(4004)));
    layer3_outputs(1860) <= layer2_outputs(3838);
    layer3_outputs(1861) <= (layer2_outputs(4672)) and not (layer2_outputs(2167));
    layer3_outputs(1862) <= (layer2_outputs(1990)) and (layer2_outputs(3801));
    layer3_outputs(1863) <= (layer2_outputs(4317)) or (layer2_outputs(398));
    layer3_outputs(1864) <= not(layer2_outputs(1219)) or (layer2_outputs(3776));
    layer3_outputs(1865) <= not(layer2_outputs(236)) or (layer2_outputs(1807));
    layer3_outputs(1866) <= (layer2_outputs(595)) and not (layer2_outputs(4473));
    layer3_outputs(1867) <= (layer2_outputs(3092)) or (layer2_outputs(936));
    layer3_outputs(1868) <= layer2_outputs(4483);
    layer3_outputs(1869) <= (layer2_outputs(2944)) xor (layer2_outputs(3247));
    layer3_outputs(1870) <= not(layer2_outputs(2248));
    layer3_outputs(1871) <= (layer2_outputs(3602)) or (layer2_outputs(4881));
    layer3_outputs(1872) <= not(layer2_outputs(4237)) or (layer2_outputs(1093));
    layer3_outputs(1873) <= not(layer2_outputs(3605)) or (layer2_outputs(1198));
    layer3_outputs(1874) <= not((layer2_outputs(2651)) or (layer2_outputs(126)));
    layer3_outputs(1875) <= not(layer2_outputs(4420)) or (layer2_outputs(3689));
    layer3_outputs(1876) <= not(layer2_outputs(693));
    layer3_outputs(1877) <= not(layer2_outputs(2223)) or (layer2_outputs(3257));
    layer3_outputs(1878) <= (layer2_outputs(2845)) and not (layer2_outputs(3716));
    layer3_outputs(1879) <= layer2_outputs(3264);
    layer3_outputs(1880) <= (layer2_outputs(4393)) or (layer2_outputs(2536));
    layer3_outputs(1881) <= layer2_outputs(2355);
    layer3_outputs(1882) <= (layer2_outputs(3428)) or (layer2_outputs(2344));
    layer3_outputs(1883) <= layer2_outputs(456);
    layer3_outputs(1884) <= (layer2_outputs(2709)) and (layer2_outputs(4467));
    layer3_outputs(1885) <= not(layer2_outputs(835));
    layer3_outputs(1886) <= not(layer2_outputs(2696));
    layer3_outputs(1887) <= layer2_outputs(4486);
    layer3_outputs(1888) <= not(layer2_outputs(331)) or (layer2_outputs(3924));
    layer3_outputs(1889) <= '1';
    layer3_outputs(1890) <= not(layer2_outputs(650)) or (layer2_outputs(3849));
    layer3_outputs(1891) <= '0';
    layer3_outputs(1892) <= layer2_outputs(2577);
    layer3_outputs(1893) <= '0';
    layer3_outputs(1894) <= '1';
    layer3_outputs(1895) <= not((layer2_outputs(4456)) and (layer2_outputs(425)));
    layer3_outputs(1896) <= not(layer2_outputs(2822)) or (layer2_outputs(1033));
    layer3_outputs(1897) <= not((layer2_outputs(3506)) or (layer2_outputs(1814)));
    layer3_outputs(1898) <= '1';
    layer3_outputs(1899) <= not(layer2_outputs(3817)) or (layer2_outputs(3743));
    layer3_outputs(1900) <= (layer2_outputs(1054)) and not (layer2_outputs(4397));
    layer3_outputs(1901) <= not(layer2_outputs(748)) or (layer2_outputs(1567));
    layer3_outputs(1902) <= not(layer2_outputs(3509));
    layer3_outputs(1903) <= '0';
    layer3_outputs(1904) <= '1';
    layer3_outputs(1905) <= layer2_outputs(917);
    layer3_outputs(1906) <= not(layer2_outputs(4855)) or (layer2_outputs(898));
    layer3_outputs(1907) <= (layer2_outputs(2613)) and (layer2_outputs(3643));
    layer3_outputs(1908) <= (layer2_outputs(1163)) and not (layer2_outputs(899));
    layer3_outputs(1909) <= (layer2_outputs(4977)) and (layer2_outputs(3679));
    layer3_outputs(1910) <= (layer2_outputs(2813)) or (layer2_outputs(3599));
    layer3_outputs(1911) <= (layer2_outputs(1796)) and not (layer2_outputs(3930));
    layer3_outputs(1912) <= '1';
    layer3_outputs(1913) <= (layer2_outputs(157)) and not (layer2_outputs(4555));
    layer3_outputs(1914) <= '1';
    layer3_outputs(1915) <= layer2_outputs(3635);
    layer3_outputs(1916) <= not(layer2_outputs(3401));
    layer3_outputs(1917) <= layer2_outputs(4590);
    layer3_outputs(1918) <= not(layer2_outputs(4657));
    layer3_outputs(1919) <= (layer2_outputs(3692)) and (layer2_outputs(3211));
    layer3_outputs(1920) <= (layer2_outputs(2061)) or (layer2_outputs(1809));
    layer3_outputs(1921) <= (layer2_outputs(4073)) and (layer2_outputs(3467));
    layer3_outputs(1922) <= not(layer2_outputs(2676)) or (layer2_outputs(3759));
    layer3_outputs(1923) <= layer2_outputs(4950);
    layer3_outputs(1924) <= not(layer2_outputs(632)) or (layer2_outputs(2811));
    layer3_outputs(1925) <= not(layer2_outputs(1328));
    layer3_outputs(1926) <= not(layer2_outputs(4150)) or (layer2_outputs(4985));
    layer3_outputs(1927) <= layer2_outputs(411);
    layer3_outputs(1928) <= layer2_outputs(114);
    layer3_outputs(1929) <= not(layer2_outputs(2556)) or (layer2_outputs(2035));
    layer3_outputs(1930) <= (layer2_outputs(5107)) and not (layer2_outputs(4609));
    layer3_outputs(1931) <= not(layer2_outputs(4715)) or (layer2_outputs(818));
    layer3_outputs(1932) <= layer2_outputs(683);
    layer3_outputs(1933) <= (layer2_outputs(1136)) and not (layer2_outputs(3670));
    layer3_outputs(1934) <= not((layer2_outputs(4542)) or (layer2_outputs(1444)));
    layer3_outputs(1935) <= not(layer2_outputs(1674));
    layer3_outputs(1936) <= not(layer2_outputs(4676)) or (layer2_outputs(2773));
    layer3_outputs(1937) <= not(layer2_outputs(2922));
    layer3_outputs(1938) <= not((layer2_outputs(2573)) or (layer2_outputs(1382)));
    layer3_outputs(1939) <= (layer2_outputs(1887)) and not (layer2_outputs(4668));
    layer3_outputs(1940) <= layer2_outputs(4333);
    layer3_outputs(1941) <= not(layer2_outputs(4856)) or (layer2_outputs(1082));
    layer3_outputs(1942) <= (layer2_outputs(2802)) and (layer2_outputs(1061));
    layer3_outputs(1943) <= not((layer2_outputs(2121)) and (layer2_outputs(4607)));
    layer3_outputs(1944) <= '0';
    layer3_outputs(1945) <= (layer2_outputs(3097)) xor (layer2_outputs(2481));
    layer3_outputs(1946) <= (layer2_outputs(2884)) and not (layer2_outputs(61));
    layer3_outputs(1947) <= '1';
    layer3_outputs(1948) <= '0';
    layer3_outputs(1949) <= layer2_outputs(2850);
    layer3_outputs(1950) <= not(layer2_outputs(3495));
    layer3_outputs(1951) <= not((layer2_outputs(4057)) or (layer2_outputs(2243)));
    layer3_outputs(1952) <= not(layer2_outputs(2819)) or (layer2_outputs(5081));
    layer3_outputs(1953) <= not(layer2_outputs(856));
    layer3_outputs(1954) <= layer2_outputs(423);
    layer3_outputs(1955) <= layer2_outputs(3855);
    layer3_outputs(1956) <= not((layer2_outputs(4387)) or (layer2_outputs(4577)));
    layer3_outputs(1957) <= not(layer2_outputs(970)) or (layer2_outputs(2744));
    layer3_outputs(1958) <= '1';
    layer3_outputs(1959) <= not((layer2_outputs(4250)) and (layer2_outputs(3467)));
    layer3_outputs(1960) <= layer2_outputs(440);
    layer3_outputs(1961) <= not((layer2_outputs(4502)) xor (layer2_outputs(3018)));
    layer3_outputs(1962) <= not(layer2_outputs(3749)) or (layer2_outputs(2653));
    layer3_outputs(1963) <= not(layer2_outputs(295));
    layer3_outputs(1964) <= '0';
    layer3_outputs(1965) <= not(layer2_outputs(4506));
    layer3_outputs(1966) <= not(layer2_outputs(1433));
    layer3_outputs(1967) <= (layer2_outputs(4370)) or (layer2_outputs(3562));
    layer3_outputs(1968) <= '1';
    layer3_outputs(1969) <= (layer2_outputs(4614)) and not (layer2_outputs(4752));
    layer3_outputs(1970) <= not(layer2_outputs(2455));
    layer3_outputs(1971) <= not(layer2_outputs(1765)) or (layer2_outputs(4845));
    layer3_outputs(1972) <= '0';
    layer3_outputs(1973) <= layer2_outputs(746);
    layer3_outputs(1974) <= layer2_outputs(2638);
    layer3_outputs(1975) <= '1';
    layer3_outputs(1976) <= '0';
    layer3_outputs(1977) <= not(layer2_outputs(3846)) or (layer2_outputs(1757));
    layer3_outputs(1978) <= not(layer2_outputs(1998));
    layer3_outputs(1979) <= (layer2_outputs(3650)) or (layer2_outputs(687));
    layer3_outputs(1980) <= not((layer2_outputs(2868)) or (layer2_outputs(1083)));
    layer3_outputs(1981) <= not((layer2_outputs(4394)) or (layer2_outputs(4279)));
    layer3_outputs(1982) <= not((layer2_outputs(1257)) and (layer2_outputs(3171)));
    layer3_outputs(1983) <= not(layer2_outputs(612)) or (layer2_outputs(4175));
    layer3_outputs(1984) <= (layer2_outputs(3367)) and not (layer2_outputs(4838));
    layer3_outputs(1985) <= not((layer2_outputs(3085)) or (layer2_outputs(1290)));
    layer3_outputs(1986) <= layer2_outputs(1448);
    layer3_outputs(1987) <= not(layer2_outputs(2654)) or (layer2_outputs(434));
    layer3_outputs(1988) <= not((layer2_outputs(4779)) or (layer2_outputs(2328)));
    layer3_outputs(1989) <= not((layer2_outputs(3483)) or (layer2_outputs(1202)));
    layer3_outputs(1990) <= layer2_outputs(1910);
    layer3_outputs(1991) <= layer2_outputs(2618);
    layer3_outputs(1992) <= layer2_outputs(4032);
    layer3_outputs(1993) <= (layer2_outputs(2964)) or (layer2_outputs(2351));
    layer3_outputs(1994) <= not(layer2_outputs(799));
    layer3_outputs(1995) <= (layer2_outputs(3491)) and not (layer2_outputs(1585));
    layer3_outputs(1996) <= not(layer2_outputs(2054));
    layer3_outputs(1997) <= layer2_outputs(4886);
    layer3_outputs(1998) <= not(layer2_outputs(3144));
    layer3_outputs(1999) <= not((layer2_outputs(2279)) and (layer2_outputs(3212)));
    layer3_outputs(2000) <= (layer2_outputs(3799)) and not (layer2_outputs(1592));
    layer3_outputs(2001) <= layer2_outputs(4715);
    layer3_outputs(2002) <= (layer2_outputs(3843)) and not (layer2_outputs(4501));
    layer3_outputs(2003) <= not(layer2_outputs(2757));
    layer3_outputs(2004) <= '0';
    layer3_outputs(2005) <= '1';
    layer3_outputs(2006) <= not((layer2_outputs(4337)) or (layer2_outputs(1623)));
    layer3_outputs(2007) <= not((layer2_outputs(1350)) and (layer2_outputs(4230)));
    layer3_outputs(2008) <= not((layer2_outputs(1015)) or (layer2_outputs(666)));
    layer3_outputs(2009) <= layer2_outputs(3806);
    layer3_outputs(2010) <= not(layer2_outputs(3227));
    layer3_outputs(2011) <= not(layer2_outputs(3721));
    layer3_outputs(2012) <= layer2_outputs(2041);
    layer3_outputs(2013) <= not(layer2_outputs(1532));
    layer3_outputs(2014) <= not(layer2_outputs(408)) or (layer2_outputs(1242));
    layer3_outputs(2015) <= not(layer2_outputs(2337)) or (layer2_outputs(2962));
    layer3_outputs(2016) <= not(layer2_outputs(3044)) or (layer2_outputs(345));
    layer3_outputs(2017) <= not(layer2_outputs(412)) or (layer2_outputs(68));
    layer3_outputs(2018) <= not(layer2_outputs(4181));
    layer3_outputs(2019) <= (layer2_outputs(3735)) and not (layer2_outputs(404));
    layer3_outputs(2020) <= layer2_outputs(4736);
    layer3_outputs(2021) <= layer2_outputs(974);
    layer3_outputs(2022) <= '1';
    layer3_outputs(2023) <= '0';
    layer3_outputs(2024) <= not(layer2_outputs(3136));
    layer3_outputs(2025) <= (layer2_outputs(3105)) and not (layer2_outputs(4643));
    layer3_outputs(2026) <= not(layer2_outputs(4205)) or (layer2_outputs(410));
    layer3_outputs(2027) <= not(layer2_outputs(2032));
    layer3_outputs(2028) <= '0';
    layer3_outputs(2029) <= not((layer2_outputs(4348)) and (layer2_outputs(607)));
    layer3_outputs(2030) <= not(layer2_outputs(1796)) or (layer2_outputs(2953));
    layer3_outputs(2031) <= '0';
    layer3_outputs(2032) <= '0';
    layer3_outputs(2033) <= (layer2_outputs(1019)) or (layer2_outputs(4319));
    layer3_outputs(2034) <= layer2_outputs(2083);
    layer3_outputs(2035) <= not(layer2_outputs(576));
    layer3_outputs(2036) <= not(layer2_outputs(4336));
    layer3_outputs(2037) <= not(layer2_outputs(1856));
    layer3_outputs(2038) <= layer2_outputs(2960);
    layer3_outputs(2039) <= not(layer2_outputs(99));
    layer3_outputs(2040) <= layer2_outputs(2527);
    layer3_outputs(2041) <= not((layer2_outputs(495)) and (layer2_outputs(363)));
    layer3_outputs(2042) <= not(layer2_outputs(4324));
    layer3_outputs(2043) <= layer2_outputs(654);
    layer3_outputs(2044) <= layer2_outputs(2686);
    layer3_outputs(2045) <= not((layer2_outputs(1777)) or (layer2_outputs(2726)));
    layer3_outputs(2046) <= layer2_outputs(2334);
    layer3_outputs(2047) <= not(layer2_outputs(1424));
    layer3_outputs(2048) <= (layer2_outputs(3120)) and not (layer2_outputs(1857));
    layer3_outputs(2049) <= not(layer2_outputs(1667));
    layer3_outputs(2050) <= not(layer2_outputs(5089)) or (layer2_outputs(1190));
    layer3_outputs(2051) <= (layer2_outputs(1218)) and not (layer2_outputs(1082));
    layer3_outputs(2052) <= not((layer2_outputs(2362)) or (layer2_outputs(4876)));
    layer3_outputs(2053) <= (layer2_outputs(2862)) and not (layer2_outputs(3260));
    layer3_outputs(2054) <= (layer2_outputs(3077)) and not (layer2_outputs(1734));
    layer3_outputs(2055) <= not(layer2_outputs(3277));
    layer3_outputs(2056) <= not(layer2_outputs(4966)) or (layer2_outputs(4999));
    layer3_outputs(2057) <= (layer2_outputs(3499)) and not (layer2_outputs(1149));
    layer3_outputs(2058) <= '0';
    layer3_outputs(2059) <= not((layer2_outputs(1644)) and (layer2_outputs(5115)));
    layer3_outputs(2060) <= not(layer2_outputs(1168)) or (layer2_outputs(793));
    layer3_outputs(2061) <= '1';
    layer3_outputs(2062) <= layer2_outputs(4561);
    layer3_outputs(2063) <= not(layer2_outputs(4185));
    layer3_outputs(2064) <= not((layer2_outputs(4461)) and (layer2_outputs(2874)));
    layer3_outputs(2065) <= not(layer2_outputs(4103));
    layer3_outputs(2066) <= not((layer2_outputs(2084)) or (layer2_outputs(4889)));
    layer3_outputs(2067) <= not((layer2_outputs(2331)) or (layer2_outputs(500)));
    layer3_outputs(2068) <= (layer2_outputs(1375)) and (layer2_outputs(309));
    layer3_outputs(2069) <= not(layer2_outputs(3548)) or (layer2_outputs(1824));
    layer3_outputs(2070) <= (layer2_outputs(3492)) and not (layer2_outputs(4771));
    layer3_outputs(2071) <= (layer2_outputs(1704)) and (layer2_outputs(4726));
    layer3_outputs(2072) <= not(layer2_outputs(1546)) or (layer2_outputs(3526));
    layer3_outputs(2073) <= (layer2_outputs(802)) and (layer2_outputs(721));
    layer3_outputs(2074) <= not(layer2_outputs(2565)) or (layer2_outputs(3561));
    layer3_outputs(2075) <= layer2_outputs(3402);
    layer3_outputs(2076) <= not((layer2_outputs(1094)) xor (layer2_outputs(2434)));
    layer3_outputs(2077) <= layer2_outputs(3306);
    layer3_outputs(2078) <= not(layer2_outputs(2086)) or (layer2_outputs(4569));
    layer3_outputs(2079) <= '0';
    layer3_outputs(2080) <= '0';
    layer3_outputs(2081) <= '0';
    layer3_outputs(2082) <= not(layer2_outputs(3877)) or (layer2_outputs(4538));
    layer3_outputs(2083) <= (layer2_outputs(831)) and not (layer2_outputs(4637));
    layer3_outputs(2084) <= not(layer2_outputs(5021)) or (layer2_outputs(730));
    layer3_outputs(2085) <= layer2_outputs(2938);
    layer3_outputs(2086) <= not((layer2_outputs(823)) or (layer2_outputs(628)));
    layer3_outputs(2087) <= not((layer2_outputs(1134)) or (layer2_outputs(312)));
    layer3_outputs(2088) <= not((layer2_outputs(608)) and (layer2_outputs(3491)));
    layer3_outputs(2089) <= (layer2_outputs(4200)) or (layer2_outputs(1556));
    layer3_outputs(2090) <= not(layer2_outputs(4952)) or (layer2_outputs(1837));
    layer3_outputs(2091) <= (layer2_outputs(812)) and (layer2_outputs(3266));
    layer3_outputs(2092) <= not((layer2_outputs(188)) or (layer2_outputs(2211)));
    layer3_outputs(2093) <= layer2_outputs(466);
    layer3_outputs(2094) <= not(layer2_outputs(2974));
    layer3_outputs(2095) <= not((layer2_outputs(554)) or (layer2_outputs(670)));
    layer3_outputs(2096) <= not(layer2_outputs(397)) or (layer2_outputs(2486));
    layer3_outputs(2097) <= (layer2_outputs(345)) and not (layer2_outputs(4151));
    layer3_outputs(2098) <= (layer2_outputs(1089)) and not (layer2_outputs(1607));
    layer3_outputs(2099) <= (layer2_outputs(2750)) and not (layer2_outputs(3242));
    layer3_outputs(2100) <= (layer2_outputs(2642)) and not (layer2_outputs(430));
    layer3_outputs(2101) <= (layer2_outputs(1962)) and not (layer2_outputs(1446));
    layer3_outputs(2102) <= layer2_outputs(1249);
    layer3_outputs(2103) <= not((layer2_outputs(2794)) and (layer2_outputs(0)));
    layer3_outputs(2104) <= (layer2_outputs(3019)) and not (layer2_outputs(738));
    layer3_outputs(2105) <= not((layer2_outputs(4191)) and (layer2_outputs(3799)));
    layer3_outputs(2106) <= (layer2_outputs(2636)) and not (layer2_outputs(1843));
    layer3_outputs(2107) <= (layer2_outputs(4703)) and not (layer2_outputs(170));
    layer3_outputs(2108) <= layer2_outputs(1586);
    layer3_outputs(2109) <= layer2_outputs(4245);
    layer3_outputs(2110) <= layer2_outputs(4806);
    layer3_outputs(2111) <= layer2_outputs(1418);
    layer3_outputs(2112) <= (layer2_outputs(2137)) and (layer2_outputs(3246));
    layer3_outputs(2113) <= not(layer2_outputs(2874));
    layer3_outputs(2114) <= (layer2_outputs(4132)) and not (layer2_outputs(4328));
    layer3_outputs(2115) <= not(layer2_outputs(1269)) or (layer2_outputs(1967));
    layer3_outputs(2116) <= not(layer2_outputs(1759)) or (layer2_outputs(4962));
    layer3_outputs(2117) <= (layer2_outputs(4179)) and not (layer2_outputs(577));
    layer3_outputs(2118) <= '0';
    layer3_outputs(2119) <= not((layer2_outputs(1882)) or (layer2_outputs(724)));
    layer3_outputs(2120) <= (layer2_outputs(5062)) and not (layer2_outputs(3546));
    layer3_outputs(2121) <= '1';
    layer3_outputs(2122) <= '0';
    layer3_outputs(2123) <= not(layer2_outputs(4567)) or (layer2_outputs(3526));
    layer3_outputs(2124) <= not(layer2_outputs(1875));
    layer3_outputs(2125) <= (layer2_outputs(3770)) and not (layer2_outputs(2393));
    layer3_outputs(2126) <= not(layer2_outputs(879)) or (layer2_outputs(3153));
    layer3_outputs(2127) <= layer2_outputs(916);
    layer3_outputs(2128) <= not(layer2_outputs(1400));
    layer3_outputs(2129) <= layer2_outputs(3834);
    layer3_outputs(2130) <= layer2_outputs(2083);
    layer3_outputs(2131) <= layer2_outputs(2621);
    layer3_outputs(2132) <= (layer2_outputs(1708)) and (layer2_outputs(3803));
    layer3_outputs(2133) <= not(layer2_outputs(2814));
    layer3_outputs(2134) <= not((layer2_outputs(957)) xor (layer2_outputs(4558)));
    layer3_outputs(2135) <= '0';
    layer3_outputs(2136) <= '0';
    layer3_outputs(2137) <= layer2_outputs(2348);
    layer3_outputs(2138) <= not(layer2_outputs(4210)) or (layer2_outputs(2087));
    layer3_outputs(2139) <= layer2_outputs(5032);
    layer3_outputs(2140) <= not((layer2_outputs(2978)) xor (layer2_outputs(2435)));
    layer3_outputs(2141) <= '0';
    layer3_outputs(2142) <= (layer2_outputs(1722)) and not (layer2_outputs(435));
    layer3_outputs(2143) <= not(layer2_outputs(4616));
    layer3_outputs(2144) <= '0';
    layer3_outputs(2145) <= not((layer2_outputs(2336)) xor (layer2_outputs(1938)));
    layer3_outputs(2146) <= layer2_outputs(5007);
    layer3_outputs(2147) <= (layer2_outputs(1613)) and (layer2_outputs(1749));
    layer3_outputs(2148) <= not(layer2_outputs(1087));
    layer3_outputs(2149) <= not(layer2_outputs(1654));
    layer3_outputs(2150) <= not(layer2_outputs(3469)) or (layer2_outputs(3873));
    layer3_outputs(2151) <= (layer2_outputs(3564)) or (layer2_outputs(695));
    layer3_outputs(2152) <= (layer2_outputs(1307)) and (layer2_outputs(515));
    layer3_outputs(2153) <= not((layer2_outputs(2055)) and (layer2_outputs(4859)));
    layer3_outputs(2154) <= not((layer2_outputs(1820)) or (layer2_outputs(4942)));
    layer3_outputs(2155) <= '1';
    layer3_outputs(2156) <= not((layer2_outputs(3169)) xor (layer2_outputs(1687)));
    layer3_outputs(2157) <= not(layer2_outputs(1503));
    layer3_outputs(2158) <= (layer2_outputs(1214)) and (layer2_outputs(3487));
    layer3_outputs(2159) <= not((layer2_outputs(525)) and (layer2_outputs(3636)));
    layer3_outputs(2160) <= layer2_outputs(5106);
    layer3_outputs(2161) <= '0';
    layer3_outputs(2162) <= (layer2_outputs(2304)) and not (layer2_outputs(1606));
    layer3_outputs(2163) <= layer2_outputs(136);
    layer3_outputs(2164) <= layer2_outputs(107);
    layer3_outputs(2165) <= not((layer2_outputs(1849)) and (layer2_outputs(2489)));
    layer3_outputs(2166) <= not((layer2_outputs(1224)) or (layer2_outputs(3843)));
    layer3_outputs(2167) <= (layer2_outputs(3655)) and not (layer2_outputs(786));
    layer3_outputs(2168) <= not(layer2_outputs(147));
    layer3_outputs(2169) <= '1';
    layer3_outputs(2170) <= (layer2_outputs(3645)) or (layer2_outputs(1584));
    layer3_outputs(2171) <= not(layer2_outputs(4589)) or (layer2_outputs(3987));
    layer3_outputs(2172) <= (layer2_outputs(1330)) and not (layer2_outputs(1502));
    layer3_outputs(2173) <= layer2_outputs(3802);
    layer3_outputs(2174) <= not((layer2_outputs(386)) or (layer2_outputs(3029)));
    layer3_outputs(2175) <= '0';
    layer3_outputs(2176) <= (layer2_outputs(4660)) and (layer2_outputs(3069));
    layer3_outputs(2177) <= '0';
    layer3_outputs(2178) <= layer2_outputs(4760);
    layer3_outputs(2179) <= layer2_outputs(2202);
    layer3_outputs(2180) <= not(layer2_outputs(4142));
    layer3_outputs(2181) <= not(layer2_outputs(246)) or (layer2_outputs(1186));
    layer3_outputs(2182) <= not(layer2_outputs(710)) or (layer2_outputs(185));
    layer3_outputs(2183) <= layer2_outputs(2740);
    layer3_outputs(2184) <= (layer2_outputs(2414)) and not (layer2_outputs(2675));
    layer3_outputs(2185) <= (layer2_outputs(3797)) and not (layer2_outputs(2608));
    layer3_outputs(2186) <= not(layer2_outputs(4187)) or (layer2_outputs(4021));
    layer3_outputs(2187) <= layer2_outputs(3427);
    layer3_outputs(2188) <= layer2_outputs(2378);
    layer3_outputs(2189) <= (layer2_outputs(3904)) and not (layer2_outputs(2586));
    layer3_outputs(2190) <= not((layer2_outputs(4673)) xor (layer2_outputs(2330)));
    layer3_outputs(2191) <= (layer2_outputs(4702)) and not (layer2_outputs(3026));
    layer3_outputs(2192) <= not((layer2_outputs(250)) xor (layer2_outputs(196)));
    layer3_outputs(2193) <= layer2_outputs(3790);
    layer3_outputs(2194) <= not((layer2_outputs(4636)) and (layer2_outputs(2600)));
    layer3_outputs(2195) <= (layer2_outputs(4335)) or (layer2_outputs(3072));
    layer3_outputs(2196) <= (layer2_outputs(1171)) xor (layer2_outputs(3401));
    layer3_outputs(2197) <= layer2_outputs(4447);
    layer3_outputs(2198) <= (layer2_outputs(2808)) and not (layer2_outputs(3422));
    layer3_outputs(2199) <= not(layer2_outputs(500));
    layer3_outputs(2200) <= (layer2_outputs(3348)) xor (layer2_outputs(1503));
    layer3_outputs(2201) <= not((layer2_outputs(4960)) or (layer2_outputs(2190)));
    layer3_outputs(2202) <= not(layer2_outputs(2716));
    layer3_outputs(2203) <= '1';
    layer3_outputs(2204) <= (layer2_outputs(301)) xor (layer2_outputs(4304));
    layer3_outputs(2205) <= (layer2_outputs(3574)) xor (layer2_outputs(2153));
    layer3_outputs(2206) <= (layer2_outputs(2176)) and not (layer2_outputs(2276));
    layer3_outputs(2207) <= not((layer2_outputs(4775)) or (layer2_outputs(1484)));
    layer3_outputs(2208) <= '0';
    layer3_outputs(2209) <= layer2_outputs(3436);
    layer3_outputs(2210) <= '0';
    layer3_outputs(2211) <= not(layer2_outputs(2088));
    layer3_outputs(2212) <= not(layer2_outputs(4841));
    layer3_outputs(2213) <= not((layer2_outputs(3848)) and (layer2_outputs(504)));
    layer3_outputs(2214) <= not(layer2_outputs(258));
    layer3_outputs(2215) <= (layer2_outputs(3249)) and not (layer2_outputs(2493));
    layer3_outputs(2216) <= '1';
    layer3_outputs(2217) <= not((layer2_outputs(5018)) and (layer2_outputs(694)));
    layer3_outputs(2218) <= not(layer2_outputs(3553));
    layer3_outputs(2219) <= (layer2_outputs(4615)) or (layer2_outputs(551));
    layer3_outputs(2220) <= not((layer2_outputs(1201)) or (layer2_outputs(144)));
    layer3_outputs(2221) <= not(layer2_outputs(3797));
    layer3_outputs(2222) <= not((layer2_outputs(397)) and (layer2_outputs(717)));
    layer3_outputs(2223) <= layer2_outputs(891);
    layer3_outputs(2224) <= (layer2_outputs(5095)) and not (layer2_outputs(4922));
    layer3_outputs(2225) <= not((layer2_outputs(2431)) and (layer2_outputs(1789)));
    layer3_outputs(2226) <= (layer2_outputs(1246)) or (layer2_outputs(3908));
    layer3_outputs(2227) <= not((layer2_outputs(2468)) and (layer2_outputs(575)));
    layer3_outputs(2228) <= not((layer2_outputs(4247)) and (layer2_outputs(4963)));
    layer3_outputs(2229) <= not((layer2_outputs(865)) and (layer2_outputs(2033)));
    layer3_outputs(2230) <= layer2_outputs(1778);
    layer3_outputs(2231) <= layer2_outputs(567);
    layer3_outputs(2232) <= '1';
    layer3_outputs(2233) <= layer2_outputs(1792);
    layer3_outputs(2234) <= layer2_outputs(966);
    layer3_outputs(2235) <= not(layer2_outputs(1801));
    layer3_outputs(2236) <= not(layer2_outputs(1041));
    layer3_outputs(2237) <= (layer2_outputs(4887)) and not (layer2_outputs(2811));
    layer3_outputs(2238) <= layer2_outputs(4836);
    layer3_outputs(2239) <= not(layer2_outputs(3882)) or (layer2_outputs(2784));
    layer3_outputs(2240) <= not(layer2_outputs(3654));
    layer3_outputs(2241) <= not((layer2_outputs(1432)) and (layer2_outputs(1557)));
    layer3_outputs(2242) <= (layer2_outputs(2272)) and not (layer2_outputs(1747));
    layer3_outputs(2243) <= (layer2_outputs(4243)) or (layer2_outputs(4002));
    layer3_outputs(2244) <= (layer2_outputs(1618)) or (layer2_outputs(2775));
    layer3_outputs(2245) <= (layer2_outputs(693)) and not (layer2_outputs(141));
    layer3_outputs(2246) <= layer2_outputs(2764);
    layer3_outputs(2247) <= (layer2_outputs(923)) and (layer2_outputs(84));
    layer3_outputs(2248) <= not(layer2_outputs(3604)) or (layer2_outputs(2643));
    layer3_outputs(2249) <= (layer2_outputs(2330)) and not (layer2_outputs(3938));
    layer3_outputs(2250) <= (layer2_outputs(3933)) or (layer2_outputs(4244));
    layer3_outputs(2251) <= layer2_outputs(3035);
    layer3_outputs(2252) <= not(layer2_outputs(3005));
    layer3_outputs(2253) <= not(layer2_outputs(4065)) or (layer2_outputs(2780));
    layer3_outputs(2254) <= (layer2_outputs(87)) and (layer2_outputs(4226));
    layer3_outputs(2255) <= (layer2_outputs(236)) and not (layer2_outputs(2354));
    layer3_outputs(2256) <= not(layer2_outputs(4889)) or (layer2_outputs(2229));
    layer3_outputs(2257) <= (layer2_outputs(903)) or (layer2_outputs(319));
    layer3_outputs(2258) <= not((layer2_outputs(238)) or (layer2_outputs(2768)));
    layer3_outputs(2259) <= not((layer2_outputs(3784)) and (layer2_outputs(3845)));
    layer3_outputs(2260) <= not(layer2_outputs(1488)) or (layer2_outputs(872));
    layer3_outputs(2261) <= '1';
    layer3_outputs(2262) <= not(layer2_outputs(608));
    layer3_outputs(2263) <= not(layer2_outputs(3577));
    layer3_outputs(2264) <= not(layer2_outputs(1458));
    layer3_outputs(2265) <= not((layer2_outputs(1806)) and (layer2_outputs(975)));
    layer3_outputs(2266) <= (layer2_outputs(967)) and (layer2_outputs(4999));
    layer3_outputs(2267) <= not(layer2_outputs(696)) or (layer2_outputs(2643));
    layer3_outputs(2268) <= not(layer2_outputs(502));
    layer3_outputs(2269) <= '0';
    layer3_outputs(2270) <= (layer2_outputs(3571)) or (layer2_outputs(4565));
    layer3_outputs(2271) <= (layer2_outputs(3818)) or (layer2_outputs(3459));
    layer3_outputs(2272) <= layer2_outputs(2925);
    layer3_outputs(2273) <= layer2_outputs(3345);
    layer3_outputs(2274) <= not(layer2_outputs(1905)) or (layer2_outputs(1591));
    layer3_outputs(2275) <= (layer2_outputs(4941)) xor (layer2_outputs(3758));
    layer3_outputs(2276) <= layer2_outputs(4291);
    layer3_outputs(2277) <= not((layer2_outputs(2790)) or (layer2_outputs(2604)));
    layer3_outputs(2278) <= (layer2_outputs(3432)) and not (layer2_outputs(2747));
    layer3_outputs(2279) <= layer2_outputs(1830);
    layer3_outputs(2280) <= layer2_outputs(2645);
    layer3_outputs(2281) <= not(layer2_outputs(854));
    layer3_outputs(2282) <= not((layer2_outputs(1291)) and (layer2_outputs(1749)));
    layer3_outputs(2283) <= '1';
    layer3_outputs(2284) <= not((layer2_outputs(2986)) or (layer2_outputs(1293)));
    layer3_outputs(2285) <= (layer2_outputs(2198)) and (layer2_outputs(1319));
    layer3_outputs(2286) <= (layer2_outputs(707)) and not (layer2_outputs(735));
    layer3_outputs(2287) <= not(layer2_outputs(2728));
    layer3_outputs(2288) <= layer2_outputs(3532);
    layer3_outputs(2289) <= (layer2_outputs(2419)) and not (layer2_outputs(2566));
    layer3_outputs(2290) <= (layer2_outputs(4911)) or (layer2_outputs(4972));
    layer3_outputs(2291) <= not((layer2_outputs(3999)) or (layer2_outputs(5056)));
    layer3_outputs(2292) <= (layer2_outputs(1264)) or (layer2_outputs(4298));
    layer3_outputs(2293) <= '1';
    layer3_outputs(2294) <= not(layer2_outputs(254));
    layer3_outputs(2295) <= layer2_outputs(4408);
    layer3_outputs(2296) <= not(layer2_outputs(2519)) or (layer2_outputs(1322));
    layer3_outputs(2297) <= layer2_outputs(792);
    layer3_outputs(2298) <= layer2_outputs(4561);
    layer3_outputs(2299) <= not((layer2_outputs(3705)) or (layer2_outputs(4518)));
    layer3_outputs(2300) <= not((layer2_outputs(2911)) or (layer2_outputs(1124)));
    layer3_outputs(2301) <= (layer2_outputs(2415)) and (layer2_outputs(1642));
    layer3_outputs(2302) <= (layer2_outputs(409)) and not (layer2_outputs(4592));
    layer3_outputs(2303) <= '1';
    layer3_outputs(2304) <= layer2_outputs(4909);
    layer3_outputs(2305) <= layer2_outputs(1791);
    layer3_outputs(2306) <= not(layer2_outputs(2378)) or (layer2_outputs(3018));
    layer3_outputs(2307) <= not((layer2_outputs(151)) or (layer2_outputs(3648)));
    layer3_outputs(2308) <= '1';
    layer3_outputs(2309) <= not(layer2_outputs(3641)) or (layer2_outputs(206));
    layer3_outputs(2310) <= not(layer2_outputs(1352)) or (layer2_outputs(4875));
    layer3_outputs(2311) <= (layer2_outputs(2420)) or (layer2_outputs(2309));
    layer3_outputs(2312) <= layer2_outputs(3521);
    layer3_outputs(2313) <= layer2_outputs(1914);
    layer3_outputs(2314) <= (layer2_outputs(2326)) or (layer2_outputs(1223));
    layer3_outputs(2315) <= not(layer2_outputs(4546));
    layer3_outputs(2316) <= (layer2_outputs(3261)) and (layer2_outputs(1043));
    layer3_outputs(2317) <= not((layer2_outputs(1429)) and (layer2_outputs(3914)));
    layer3_outputs(2318) <= (layer2_outputs(1386)) and not (layer2_outputs(2451));
    layer3_outputs(2319) <= (layer2_outputs(3327)) or (layer2_outputs(4727));
    layer3_outputs(2320) <= (layer2_outputs(4928)) and not (layer2_outputs(1398));
    layer3_outputs(2321) <= not(layer2_outputs(1721));
    layer3_outputs(2322) <= not(layer2_outputs(4784));
    layer3_outputs(2323) <= (layer2_outputs(2741)) xor (layer2_outputs(1724));
    layer3_outputs(2324) <= not((layer2_outputs(2296)) xor (layer2_outputs(825)));
    layer3_outputs(2325) <= not(layer2_outputs(2600));
    layer3_outputs(2326) <= layer2_outputs(1844);
    layer3_outputs(2327) <= not((layer2_outputs(3184)) or (layer2_outputs(2194)));
    layer3_outputs(2328) <= not(layer2_outputs(4613));
    layer3_outputs(2329) <= (layer2_outputs(2276)) and not (layer2_outputs(57));
    layer3_outputs(2330) <= layer2_outputs(464);
    layer3_outputs(2331) <= '0';
    layer3_outputs(2332) <= layer2_outputs(2722);
    layer3_outputs(2333) <= '0';
    layer3_outputs(2334) <= (layer2_outputs(19)) and not (layer2_outputs(1723));
    layer3_outputs(2335) <= (layer2_outputs(2256)) and not (layer2_outputs(2763));
    layer3_outputs(2336) <= (layer2_outputs(2702)) or (layer2_outputs(2931));
    layer3_outputs(2337) <= (layer2_outputs(1829)) and (layer2_outputs(2777));
    layer3_outputs(2338) <= '0';
    layer3_outputs(2339) <= (layer2_outputs(4980)) and not (layer2_outputs(4620));
    layer3_outputs(2340) <= (layer2_outputs(2614)) or (layer2_outputs(3407));
    layer3_outputs(2341) <= layer2_outputs(17);
    layer3_outputs(2342) <= not(layer2_outputs(3473));
    layer3_outputs(2343) <= (layer2_outputs(876)) and not (layer2_outputs(3347));
    layer3_outputs(2344) <= (layer2_outputs(277)) or (layer2_outputs(814));
    layer3_outputs(2345) <= (layer2_outputs(4581)) and not (layer2_outputs(4509));
    layer3_outputs(2346) <= (layer2_outputs(1148)) or (layer2_outputs(3700));
    layer3_outputs(2347) <= not(layer2_outputs(2035)) or (layer2_outputs(197));
    layer3_outputs(2348) <= not(layer2_outputs(4385));
    layer3_outputs(2349) <= '1';
    layer3_outputs(2350) <= not((layer2_outputs(3557)) or (layer2_outputs(1541)));
    layer3_outputs(2351) <= layer2_outputs(1912);
    layer3_outputs(2352) <= (layer2_outputs(1990)) and (layer2_outputs(2515));
    layer3_outputs(2353) <= not(layer2_outputs(2194)) or (layer2_outputs(789));
    layer3_outputs(2354) <= not(layer2_outputs(2667));
    layer3_outputs(2355) <= '0';
    layer3_outputs(2356) <= layer2_outputs(4910);
    layer3_outputs(2357) <= layer2_outputs(830);
    layer3_outputs(2358) <= (layer2_outputs(1059)) and not (layer2_outputs(2696));
    layer3_outputs(2359) <= not(layer2_outputs(3300));
    layer3_outputs(2360) <= not(layer2_outputs(4353));
    layer3_outputs(2361) <= not(layer2_outputs(4926));
    layer3_outputs(2362) <= '1';
    layer3_outputs(2363) <= '0';
    layer3_outputs(2364) <= layer2_outputs(2650);
    layer3_outputs(2365) <= layer2_outputs(2372);
    layer3_outputs(2366) <= layer2_outputs(2099);
    layer3_outputs(2367) <= (layer2_outputs(1160)) and (layer2_outputs(1690));
    layer3_outputs(2368) <= not(layer2_outputs(3343));
    layer3_outputs(2369) <= '1';
    layer3_outputs(2370) <= not((layer2_outputs(3835)) or (layer2_outputs(960)));
    layer3_outputs(2371) <= not((layer2_outputs(4961)) or (layer2_outputs(4608)));
    layer3_outputs(2372) <= (layer2_outputs(36)) and not (layer2_outputs(3949));
    layer3_outputs(2373) <= (layer2_outputs(4687)) and not (layer2_outputs(3511));
    layer3_outputs(2374) <= '1';
    layer3_outputs(2375) <= (layer2_outputs(2599)) and not (layer2_outputs(2622));
    layer3_outputs(2376) <= not(layer2_outputs(4511));
    layer3_outputs(2377) <= not(layer2_outputs(3376));
    layer3_outputs(2378) <= layer2_outputs(4864);
    layer3_outputs(2379) <= not(layer2_outputs(3674));
    layer3_outputs(2380) <= '1';
    layer3_outputs(2381) <= not(layer2_outputs(4468));
    layer3_outputs(2382) <= not(layer2_outputs(1784)) or (layer2_outputs(685));
    layer3_outputs(2383) <= not((layer2_outputs(1324)) and (layer2_outputs(1435)));
    layer3_outputs(2384) <= '1';
    layer3_outputs(2385) <= '1';
    layer3_outputs(2386) <= not(layer2_outputs(4834)) or (layer2_outputs(479));
    layer3_outputs(2387) <= not((layer2_outputs(4108)) or (layer2_outputs(1473)));
    layer3_outputs(2388) <= (layer2_outputs(5045)) and (layer2_outputs(1655));
    layer3_outputs(2389) <= layer2_outputs(1942);
    layer3_outputs(2390) <= not(layer2_outputs(4063)) or (layer2_outputs(1924));
    layer3_outputs(2391) <= not(layer2_outputs(4395));
    layer3_outputs(2392) <= (layer2_outputs(1559)) and not (layer2_outputs(4380));
    layer3_outputs(2393) <= not(layer2_outputs(789)) or (layer2_outputs(3316));
    layer3_outputs(2394) <= (layer2_outputs(209)) and not (layer2_outputs(1438));
    layer3_outputs(2395) <= (layer2_outputs(4176)) or (layer2_outputs(2731));
    layer3_outputs(2396) <= not((layer2_outputs(3196)) or (layer2_outputs(3885)));
    layer3_outputs(2397) <= '1';
    layer3_outputs(2398) <= not(layer2_outputs(2567));
    layer3_outputs(2399) <= not((layer2_outputs(3519)) or (layer2_outputs(1187)));
    layer3_outputs(2400) <= (layer2_outputs(803)) and not (layer2_outputs(1002));
    layer3_outputs(2401) <= not(layer2_outputs(2814)) or (layer2_outputs(1950));
    layer3_outputs(2402) <= (layer2_outputs(2277)) xor (layer2_outputs(1871));
    layer3_outputs(2403) <= not(layer2_outputs(334)) or (layer2_outputs(2302));
    layer3_outputs(2404) <= (layer2_outputs(2548)) and not (layer2_outputs(41));
    layer3_outputs(2405) <= not((layer2_outputs(167)) and (layer2_outputs(115)));
    layer3_outputs(2406) <= not(layer2_outputs(2450));
    layer3_outputs(2407) <= '1';
    layer3_outputs(2408) <= (layer2_outputs(2011)) and (layer2_outputs(3271));
    layer3_outputs(2409) <= layer2_outputs(4594);
    layer3_outputs(2410) <= layer2_outputs(4502);
    layer3_outputs(2411) <= (layer2_outputs(1930)) or (layer2_outputs(2039));
    layer3_outputs(2412) <= not(layer2_outputs(935));
    layer3_outputs(2413) <= '0';
    layer3_outputs(2414) <= (layer2_outputs(3224)) and (layer2_outputs(1157));
    layer3_outputs(2415) <= layer2_outputs(1497);
    layer3_outputs(2416) <= not((layer2_outputs(2048)) or (layer2_outputs(1568)));
    layer3_outputs(2417) <= '1';
    layer3_outputs(2418) <= (layer2_outputs(1020)) and not (layer2_outputs(4504));
    layer3_outputs(2419) <= layer2_outputs(3760);
    layer3_outputs(2420) <= (layer2_outputs(2122)) and not (layer2_outputs(1271));
    layer3_outputs(2421) <= layer2_outputs(214);
    layer3_outputs(2422) <= (layer2_outputs(5063)) and not (layer2_outputs(4501));
    layer3_outputs(2423) <= (layer2_outputs(3950)) and not (layer2_outputs(2865));
    layer3_outputs(2424) <= (layer2_outputs(928)) and (layer2_outputs(5112));
    layer3_outputs(2425) <= (layer2_outputs(3386)) or (layer2_outputs(1920));
    layer3_outputs(2426) <= not(layer2_outputs(4114));
    layer3_outputs(2427) <= (layer2_outputs(4706)) and not (layer2_outputs(1276));
    layer3_outputs(2428) <= not((layer2_outputs(4981)) and (layer2_outputs(1501)));
    layer3_outputs(2429) <= not(layer2_outputs(134)) or (layer2_outputs(5114));
    layer3_outputs(2430) <= layer2_outputs(293);
    layer3_outputs(2431) <= '1';
    layer3_outputs(2432) <= not(layer2_outputs(586)) or (layer2_outputs(2901));
    layer3_outputs(2433) <= (layer2_outputs(4584)) and not (layer2_outputs(969));
    layer3_outputs(2434) <= '0';
    layer3_outputs(2435) <= not(layer2_outputs(3498));
    layer3_outputs(2436) <= not((layer2_outputs(2585)) or (layer2_outputs(1118)));
    layer3_outputs(2437) <= not(layer2_outputs(3464)) or (layer2_outputs(65));
    layer3_outputs(2438) <= layer2_outputs(5041);
    layer3_outputs(2439) <= not(layer2_outputs(1651)) or (layer2_outputs(323));
    layer3_outputs(2440) <= not(layer2_outputs(2840));
    layer3_outputs(2441) <= not(layer2_outputs(2139)) or (layer2_outputs(4893));
    layer3_outputs(2442) <= not(layer2_outputs(2258)) or (layer2_outputs(2826));
    layer3_outputs(2443) <= '0';
    layer3_outputs(2444) <= (layer2_outputs(3572)) and not (layer2_outputs(4555));
    layer3_outputs(2445) <= (layer2_outputs(2301)) or (layer2_outputs(738));
    layer3_outputs(2446) <= not((layer2_outputs(2034)) and (layer2_outputs(1327)));
    layer3_outputs(2447) <= not((layer2_outputs(1479)) and (layer2_outputs(290)));
    layer3_outputs(2448) <= not(layer2_outputs(2829)) or (layer2_outputs(1025));
    layer3_outputs(2449) <= not((layer2_outputs(3972)) or (layer2_outputs(3676)));
    layer3_outputs(2450) <= not(layer2_outputs(1775)) or (layer2_outputs(1790));
    layer3_outputs(2451) <= '1';
    layer3_outputs(2452) <= (layer2_outputs(3257)) and not (layer2_outputs(192));
    layer3_outputs(2453) <= not((layer2_outputs(3114)) and (layer2_outputs(2772)));
    layer3_outputs(2454) <= (layer2_outputs(2900)) or (layer2_outputs(1860));
    layer3_outputs(2455) <= (layer2_outputs(4095)) or (layer2_outputs(4008));
    layer3_outputs(2456) <= '1';
    layer3_outputs(2457) <= (layer2_outputs(1256)) and not (layer2_outputs(180));
    layer3_outputs(2458) <= not(layer2_outputs(2394));
    layer3_outputs(2459) <= layer2_outputs(399);
    layer3_outputs(2460) <= layer2_outputs(1981);
    layer3_outputs(2461) <= layer2_outputs(548);
    layer3_outputs(2462) <= layer2_outputs(3076);
    layer3_outputs(2463) <= layer2_outputs(1315);
    layer3_outputs(2464) <= not(layer2_outputs(1502)) or (layer2_outputs(2906));
    layer3_outputs(2465) <= (layer2_outputs(2654)) and not (layer2_outputs(3505));
    layer3_outputs(2466) <= layer2_outputs(4172);
    layer3_outputs(2467) <= layer2_outputs(1396);
    layer3_outputs(2468) <= not(layer2_outputs(2109));
    layer3_outputs(2469) <= (layer2_outputs(1562)) and not (layer2_outputs(2656));
    layer3_outputs(2470) <= layer2_outputs(4546);
    layer3_outputs(2471) <= not(layer2_outputs(650)) or (layer2_outputs(1351));
    layer3_outputs(2472) <= (layer2_outputs(4472)) and not (layer2_outputs(2981));
    layer3_outputs(2473) <= '0';
    layer3_outputs(2474) <= (layer2_outputs(4493)) and not (layer2_outputs(2057));
    layer3_outputs(2475) <= not((layer2_outputs(1132)) and (layer2_outputs(1977)));
    layer3_outputs(2476) <= (layer2_outputs(3698)) and not (layer2_outputs(4863));
    layer3_outputs(2477) <= not(layer2_outputs(1554));
    layer3_outputs(2478) <= not((layer2_outputs(3009)) or (layer2_outputs(4799)));
    layer3_outputs(2479) <= '1';
    layer3_outputs(2480) <= (layer2_outputs(2130)) and not (layer2_outputs(3139));
    layer3_outputs(2481) <= layer2_outputs(3035);
    layer3_outputs(2482) <= not(layer2_outputs(4158));
    layer3_outputs(2483) <= not(layer2_outputs(2488)) or (layer2_outputs(920));
    layer3_outputs(2484) <= not((layer2_outputs(1112)) and (layer2_outputs(3549)));
    layer3_outputs(2485) <= not((layer2_outputs(822)) and (layer2_outputs(223)));
    layer3_outputs(2486) <= not(layer2_outputs(2503));
    layer3_outputs(2487) <= (layer2_outputs(1119)) or (layer2_outputs(2246));
    layer3_outputs(2488) <= not((layer2_outputs(4544)) or (layer2_outputs(48)));
    layer3_outputs(2489) <= not(layer2_outputs(3129));
    layer3_outputs(2490) <= (layer2_outputs(1115)) and not (layer2_outputs(561));
    layer3_outputs(2491) <= not((layer2_outputs(3955)) or (layer2_outputs(2300)));
    layer3_outputs(2492) <= layer2_outputs(1688);
    layer3_outputs(2493) <= layer2_outputs(4745);
    layer3_outputs(2494) <= not(layer2_outputs(2073));
    layer3_outputs(2495) <= (layer2_outputs(1948)) or (layer2_outputs(3210));
    layer3_outputs(2496) <= not(layer2_outputs(5022)) or (layer2_outputs(696));
    layer3_outputs(2497) <= not((layer2_outputs(2733)) or (layer2_outputs(880)));
    layer3_outputs(2498) <= not(layer2_outputs(1682)) or (layer2_outputs(1657));
    layer3_outputs(2499) <= (layer2_outputs(1021)) xor (layer2_outputs(1527));
    layer3_outputs(2500) <= (layer2_outputs(4809)) or (layer2_outputs(2666));
    layer3_outputs(2501) <= not((layer2_outputs(3947)) xor (layer2_outputs(4872)));
    layer3_outputs(2502) <= not((layer2_outputs(3913)) and (layer2_outputs(1545)));
    layer3_outputs(2503) <= not(layer2_outputs(2976));
    layer3_outputs(2504) <= not((layer2_outputs(578)) and (layer2_outputs(3021)));
    layer3_outputs(2505) <= (layer2_outputs(2632)) and not (layer2_outputs(1969));
    layer3_outputs(2506) <= not(layer2_outputs(241));
    layer3_outputs(2507) <= (layer2_outputs(3538)) and not (layer2_outputs(1097));
    layer3_outputs(2508) <= not((layer2_outputs(1162)) and (layer2_outputs(368)));
    layer3_outputs(2509) <= not(layer2_outputs(3772));
    layer3_outputs(2510) <= not(layer2_outputs(3184));
    layer3_outputs(2511) <= not((layer2_outputs(2776)) xor (layer2_outputs(2886)));
    layer3_outputs(2512) <= not(layer2_outputs(4514)) or (layer2_outputs(438));
    layer3_outputs(2513) <= '0';
    layer3_outputs(2514) <= not(layer2_outputs(1663));
    layer3_outputs(2515) <= (layer2_outputs(2104)) and not (layer2_outputs(2991));
    layer3_outputs(2516) <= not(layer2_outputs(3981));
    layer3_outputs(2517) <= (layer2_outputs(1806)) and (layer2_outputs(5058));
    layer3_outputs(2518) <= not(layer2_outputs(2954)) or (layer2_outputs(1557));
    layer3_outputs(2519) <= not(layer2_outputs(229));
    layer3_outputs(2520) <= layer2_outputs(2240);
    layer3_outputs(2521) <= layer2_outputs(2026);
    layer3_outputs(2522) <= layer2_outputs(4186);
    layer3_outputs(2523) <= not(layer2_outputs(3371));
    layer3_outputs(2524) <= not((layer2_outputs(4069)) and (layer2_outputs(2426)));
    layer3_outputs(2525) <= not(layer2_outputs(3754)) or (layer2_outputs(1456));
    layer3_outputs(2526) <= '0';
    layer3_outputs(2527) <= '1';
    layer3_outputs(2528) <= (layer2_outputs(1800)) or (layer2_outputs(3235));
    layer3_outputs(2529) <= (layer2_outputs(3942)) or (layer2_outputs(3269));
    layer3_outputs(2530) <= (layer2_outputs(4084)) and (layer2_outputs(4366));
    layer3_outputs(2531) <= not(layer2_outputs(1354));
    layer3_outputs(2532) <= not(layer2_outputs(1324));
    layer3_outputs(2533) <= not(layer2_outputs(3391));
    layer3_outputs(2534) <= not((layer2_outputs(1718)) or (layer2_outputs(4586)));
    layer3_outputs(2535) <= (layer2_outputs(1636)) or (layer2_outputs(4251));
    layer3_outputs(2536) <= not(layer2_outputs(4711));
    layer3_outputs(2537) <= not((layer2_outputs(1241)) and (layer2_outputs(4113)));
    layer3_outputs(2538) <= not(layer2_outputs(2456));
    layer3_outputs(2539) <= '1';
    layer3_outputs(2540) <= layer2_outputs(2952);
    layer3_outputs(2541) <= (layer2_outputs(3607)) and not (layer2_outputs(3740));
    layer3_outputs(2542) <= layer2_outputs(939);
    layer3_outputs(2543) <= '0';
    layer3_outputs(2544) <= (layer2_outputs(2569)) and not (layer2_outputs(111));
    layer3_outputs(2545) <= layer2_outputs(3430);
    layer3_outputs(2546) <= layer2_outputs(774);
    layer3_outputs(2547) <= layer2_outputs(2434);
    layer3_outputs(2548) <= layer2_outputs(2096);
    layer3_outputs(2549) <= (layer2_outputs(614)) and not (layer2_outputs(4707));
    layer3_outputs(2550) <= not((layer2_outputs(343)) or (layer2_outputs(3412)));
    layer3_outputs(2551) <= not(layer2_outputs(119));
    layer3_outputs(2552) <= not((layer2_outputs(2430)) or (layer2_outputs(912)));
    layer3_outputs(2553) <= not((layer2_outputs(4262)) or (layer2_outputs(1696)));
    layer3_outputs(2554) <= (layer2_outputs(3236)) and (layer2_outputs(1686));
    layer3_outputs(2555) <= not(layer2_outputs(4178));
    layer3_outputs(2556) <= not(layer2_outputs(3001));
    layer3_outputs(2557) <= not(layer2_outputs(3913)) or (layer2_outputs(4903));
    layer3_outputs(2558) <= (layer2_outputs(5116)) or (layer2_outputs(3133));
    layer3_outputs(2559) <= (layer2_outputs(4519)) and not (layer2_outputs(1987));
    layer3_outputs(2560) <= not((layer2_outputs(2897)) or (layer2_outputs(1953)));
    layer3_outputs(2561) <= (layer2_outputs(214)) and not (layer2_outputs(2997));
    layer3_outputs(2562) <= not((layer2_outputs(432)) or (layer2_outputs(1942)));
    layer3_outputs(2563) <= '1';
    layer3_outputs(2564) <= (layer2_outputs(633)) or (layer2_outputs(4358));
    layer3_outputs(2565) <= not(layer2_outputs(2241)) or (layer2_outputs(568));
    layer3_outputs(2566) <= not(layer2_outputs(3711)) or (layer2_outputs(2239));
    layer3_outputs(2567) <= layer2_outputs(487);
    layer3_outputs(2568) <= (layer2_outputs(2366)) and (layer2_outputs(3034));
    layer3_outputs(2569) <= (layer2_outputs(1524)) or (layer2_outputs(2205));
    layer3_outputs(2570) <= layer2_outputs(3717);
    layer3_outputs(2571) <= '0';
    layer3_outputs(2572) <= not(layer2_outputs(4771)) or (layer2_outputs(4842));
    layer3_outputs(2573) <= (layer2_outputs(2841)) or (layer2_outputs(3771));
    layer3_outputs(2574) <= not((layer2_outputs(2596)) and (layer2_outputs(4662)));
    layer3_outputs(2575) <= not(layer2_outputs(4761)) or (layer2_outputs(447));
    layer3_outputs(2576) <= not(layer2_outputs(3726)) or (layer2_outputs(4482));
    layer3_outputs(2577) <= not((layer2_outputs(3594)) and (layer2_outputs(2268)));
    layer3_outputs(2578) <= '0';
    layer3_outputs(2579) <= '1';
    layer3_outputs(2580) <= not(layer2_outputs(3579)) or (layer2_outputs(4624));
    layer3_outputs(2581) <= not(layer2_outputs(2213));
    layer3_outputs(2582) <= not((layer2_outputs(3502)) or (layer2_outputs(4056)));
    layer3_outputs(2583) <= not(layer2_outputs(3310));
    layer3_outputs(2584) <= layer2_outputs(3009);
    layer3_outputs(2585) <= '1';
    layer3_outputs(2586) <= not((layer2_outputs(760)) or (layer2_outputs(857)));
    layer3_outputs(2587) <= not(layer2_outputs(281)) or (layer2_outputs(652));
    layer3_outputs(2588) <= not(layer2_outputs(1635)) or (layer2_outputs(523));
    layer3_outputs(2589) <= not(layer2_outputs(790));
    layer3_outputs(2590) <= '1';
    layer3_outputs(2591) <= '1';
    layer3_outputs(2592) <= (layer2_outputs(203)) or (layer2_outputs(4040));
    layer3_outputs(2593) <= (layer2_outputs(2228)) and not (layer2_outputs(2677));
    layer3_outputs(2594) <= '1';
    layer3_outputs(2595) <= (layer2_outputs(4437)) and (layer2_outputs(3370));
    layer3_outputs(2596) <= '1';
    layer3_outputs(2597) <= (layer2_outputs(2987)) and not (layer2_outputs(3013));
    layer3_outputs(2598) <= not(layer2_outputs(4644)) or (layer2_outputs(1681));
    layer3_outputs(2599) <= not(layer2_outputs(4551));
    layer3_outputs(2600) <= not(layer2_outputs(1023));
    layer3_outputs(2601) <= (layer2_outputs(2507)) or (layer2_outputs(1166));
    layer3_outputs(2602) <= (layer2_outputs(3586)) and (layer2_outputs(12));
    layer3_outputs(2603) <= not(layer2_outputs(2648));
    layer3_outputs(2604) <= layer2_outputs(123);
    layer3_outputs(2605) <= (layer2_outputs(4027)) and not (layer2_outputs(1623));
    layer3_outputs(2606) <= (layer2_outputs(1839)) and not (layer2_outputs(4744));
    layer3_outputs(2607) <= (layer2_outputs(4026)) and not (layer2_outputs(191));
    layer3_outputs(2608) <= not(layer2_outputs(676));
    layer3_outputs(2609) <= '0';
    layer3_outputs(2610) <= not((layer2_outputs(4556)) xor (layer2_outputs(4533)));
    layer3_outputs(2611) <= not(layer2_outputs(204));
    layer3_outputs(2612) <= (layer2_outputs(956)) and not (layer2_outputs(1369));
    layer3_outputs(2613) <= not(layer2_outputs(5026));
    layer3_outputs(2614) <= (layer2_outputs(3048)) or (layer2_outputs(4949));
    layer3_outputs(2615) <= (layer2_outputs(1458)) and not (layer2_outputs(3516));
    layer3_outputs(2616) <= not(layer2_outputs(1511));
    layer3_outputs(2617) <= layer2_outputs(2795);
    layer3_outputs(2618) <= layer2_outputs(3746);
    layer3_outputs(2619) <= layer2_outputs(806);
    layer3_outputs(2620) <= (layer2_outputs(759)) and not (layer2_outputs(3706));
    layer3_outputs(2621) <= not(layer2_outputs(473)) or (layer2_outputs(228));
    layer3_outputs(2622) <= '1';
    layer3_outputs(2623) <= not(layer2_outputs(4576)) or (layer2_outputs(3362));
    layer3_outputs(2624) <= not(layer2_outputs(2917)) or (layer2_outputs(4168));
    layer3_outputs(2625) <= layer2_outputs(2071);
    layer3_outputs(2626) <= layer2_outputs(3704);
    layer3_outputs(2627) <= not((layer2_outputs(1074)) or (layer2_outputs(1174)));
    layer3_outputs(2628) <= (layer2_outputs(2858)) and not (layer2_outputs(2232));
    layer3_outputs(2629) <= (layer2_outputs(468)) or (layer2_outputs(4696));
    layer3_outputs(2630) <= (layer2_outputs(3544)) or (layer2_outputs(3866));
    layer3_outputs(2631) <= layer2_outputs(1930);
    layer3_outputs(2632) <= not(layer2_outputs(863)) or (layer2_outputs(605));
    layer3_outputs(2633) <= '1';
    layer3_outputs(2634) <= not(layer2_outputs(3205));
    layer3_outputs(2635) <= layer2_outputs(4151);
    layer3_outputs(2636) <= not(layer2_outputs(3831));
    layer3_outputs(2637) <= not(layer2_outputs(3017));
    layer3_outputs(2638) <= not(layer2_outputs(1705));
    layer3_outputs(2639) <= '0';
    layer3_outputs(2640) <= not((layer2_outputs(1038)) or (layer2_outputs(5080)));
    layer3_outputs(2641) <= layer2_outputs(4697);
    layer3_outputs(2642) <= not(layer2_outputs(2754));
    layer3_outputs(2643) <= layer2_outputs(3380);
    layer3_outputs(2644) <= layer2_outputs(1057);
    layer3_outputs(2645) <= (layer2_outputs(1138)) and (layer2_outputs(3398));
    layer3_outputs(2646) <= layer2_outputs(4937);
    layer3_outputs(2647) <= '1';
    layer3_outputs(2648) <= (layer2_outputs(2304)) and (layer2_outputs(3810));
    layer3_outputs(2649) <= not(layer2_outputs(1629)) or (layer2_outputs(4918));
    layer3_outputs(2650) <= (layer2_outputs(1303)) and not (layer2_outputs(4641));
    layer3_outputs(2651) <= not(layer2_outputs(443));
    layer3_outputs(2652) <= '0';
    layer3_outputs(2653) <= (layer2_outputs(2052)) and not (layer2_outputs(3160));
    layer3_outputs(2654) <= not((layer2_outputs(4632)) and (layer2_outputs(4794)));
    layer3_outputs(2655) <= layer2_outputs(4355);
    layer3_outputs(2656) <= not(layer2_outputs(1507));
    layer3_outputs(2657) <= not(layer2_outputs(2812));
    layer3_outputs(2658) <= layer2_outputs(3997);
    layer3_outputs(2659) <= not(layer2_outputs(2294)) or (layer2_outputs(3580));
    layer3_outputs(2660) <= '1';
    layer3_outputs(2661) <= not(layer2_outputs(3736));
    layer3_outputs(2662) <= '0';
    layer3_outputs(2663) <= layer2_outputs(3888);
    layer3_outputs(2664) <= not(layer2_outputs(2148));
    layer3_outputs(2665) <= not((layer2_outputs(2225)) and (layer2_outputs(4218)));
    layer3_outputs(2666) <= layer2_outputs(1161);
    layer3_outputs(2667) <= '0';
    layer3_outputs(2668) <= not(layer2_outputs(1032)) or (layer2_outputs(3775));
    layer3_outputs(2669) <= not(layer2_outputs(4925));
    layer3_outputs(2670) <= not(layer2_outputs(2685));
    layer3_outputs(2671) <= (layer2_outputs(2095)) and not (layer2_outputs(4806));
    layer3_outputs(2672) <= layer2_outputs(4557);
    layer3_outputs(2673) <= layer2_outputs(198);
    layer3_outputs(2674) <= (layer2_outputs(1475)) and (layer2_outputs(4360));
    layer3_outputs(2675) <= layer2_outputs(2883);
    layer3_outputs(2676) <= not(layer2_outputs(985));
    layer3_outputs(2677) <= not((layer2_outputs(5075)) or (layer2_outputs(1457)));
    layer3_outputs(2678) <= (layer2_outputs(4040)) and (layer2_outputs(4938));
    layer3_outputs(2679) <= layer2_outputs(225);
    layer3_outputs(2680) <= not(layer2_outputs(3849));
    layer3_outputs(2681) <= layer2_outputs(3297);
    layer3_outputs(2682) <= not(layer2_outputs(3344));
    layer3_outputs(2683) <= not((layer2_outputs(5101)) and (layer2_outputs(1936)));
    layer3_outputs(2684) <= not(layer2_outputs(292));
    layer3_outputs(2685) <= not((layer2_outputs(1770)) or (layer2_outputs(4390)));
    layer3_outputs(2686) <= not(layer2_outputs(3713));
    layer3_outputs(2687) <= not(layer2_outputs(4729)) or (layer2_outputs(128));
    layer3_outputs(2688) <= (layer2_outputs(3744)) or (layer2_outputs(3875));
    layer3_outputs(2689) <= '1';
    layer3_outputs(2690) <= not(layer2_outputs(5096)) or (layer2_outputs(24));
    layer3_outputs(2691) <= not((layer2_outputs(4268)) or (layer2_outputs(2508)));
    layer3_outputs(2692) <= (layer2_outputs(3862)) and not (layer2_outputs(4379));
    layer3_outputs(2693) <= (layer2_outputs(941)) or (layer2_outputs(4720));
    layer3_outputs(2694) <= '0';
    layer3_outputs(2695) <= not((layer2_outputs(2691)) and (layer2_outputs(4170)));
    layer3_outputs(2696) <= (layer2_outputs(4278)) or (layer2_outputs(664));
    layer3_outputs(2697) <= '1';
    layer3_outputs(2698) <= '1';
    layer3_outputs(2699) <= layer2_outputs(1061);
    layer3_outputs(2700) <= layer2_outputs(250);
    layer3_outputs(2701) <= layer2_outputs(259);
    layer3_outputs(2702) <= layer2_outputs(3312);
    layer3_outputs(2703) <= not(layer2_outputs(1709)) or (layer2_outputs(3059));
    layer3_outputs(2704) <= not((layer2_outputs(4242)) and (layer2_outputs(4265)));
    layer3_outputs(2705) <= layer2_outputs(4304);
    layer3_outputs(2706) <= not(layer2_outputs(2718)) or (layer2_outputs(4405));
    layer3_outputs(2707) <= layer2_outputs(2878);
    layer3_outputs(2708) <= layer2_outputs(2770);
    layer3_outputs(2709) <= layer2_outputs(640);
    layer3_outputs(2710) <= (layer2_outputs(3451)) and not (layer2_outputs(3));
    layer3_outputs(2711) <= layer2_outputs(4269);
    layer3_outputs(2712) <= '1';
    layer3_outputs(2713) <= (layer2_outputs(600)) or (layer2_outputs(3422));
    layer3_outputs(2714) <= not(layer2_outputs(3022));
    layer3_outputs(2715) <= layer2_outputs(1926);
    layer3_outputs(2716) <= layer2_outputs(4171);
    layer3_outputs(2717) <= (layer2_outputs(651)) xor (layer2_outputs(3971));
    layer3_outputs(2718) <= not(layer2_outputs(4848)) or (layer2_outputs(3334));
    layer3_outputs(2719) <= not((layer2_outputs(4294)) xor (layer2_outputs(2599)));
    layer3_outputs(2720) <= (layer2_outputs(3149)) or (layer2_outputs(4419));
    layer3_outputs(2721) <= layer2_outputs(4909);
    layer3_outputs(2722) <= (layer2_outputs(1355)) and not (layer2_outputs(1754));
    layer3_outputs(2723) <= not(layer2_outputs(1733)) or (layer2_outputs(508));
    layer3_outputs(2724) <= (layer2_outputs(1436)) and (layer2_outputs(3874));
    layer3_outputs(2725) <= layer2_outputs(1053);
    layer3_outputs(2726) <= not((layer2_outputs(4674)) or (layer2_outputs(2762)));
    layer3_outputs(2727) <= layer2_outputs(2875);
    layer3_outputs(2728) <= (layer2_outputs(378)) and not (layer2_outputs(3300));
    layer3_outputs(2729) <= (layer2_outputs(3638)) or (layer2_outputs(4791));
    layer3_outputs(2730) <= '0';
    layer3_outputs(2731) <= not(layer2_outputs(2809)) or (layer2_outputs(749));
    layer3_outputs(2732) <= (layer2_outputs(3862)) or (layer2_outputs(1904));
    layer3_outputs(2733) <= not(layer2_outputs(1554));
    layer3_outputs(2734) <= '0';
    layer3_outputs(2735) <= not(layer2_outputs(581));
    layer3_outputs(2736) <= '0';
    layer3_outputs(2737) <= layer2_outputs(978);
    layer3_outputs(2738) <= '1';
    layer3_outputs(2739) <= (layer2_outputs(2791)) or (layer2_outputs(1222));
    layer3_outputs(2740) <= not(layer2_outputs(4605));
    layer3_outputs(2741) <= not(layer2_outputs(2900));
    layer3_outputs(2742) <= layer2_outputs(3372);
    layer3_outputs(2743) <= '0';
    layer3_outputs(2744) <= not(layer2_outputs(955)) or (layer2_outputs(1735));
    layer3_outputs(2745) <= layer2_outputs(846);
    layer3_outputs(2746) <= not((layer2_outputs(2683)) or (layer2_outputs(5029)));
    layer3_outputs(2747) <= not(layer2_outputs(1254));
    layer3_outputs(2748) <= not(layer2_outputs(1355));
    layer3_outputs(2749) <= not((layer2_outputs(1043)) and (layer2_outputs(3067)));
    layer3_outputs(2750) <= '1';
    layer3_outputs(2751) <= layer2_outputs(4980);
    layer3_outputs(2752) <= '0';
    layer3_outputs(2753) <= not(layer2_outputs(3025)) or (layer2_outputs(4224));
    layer3_outputs(2754) <= not(layer2_outputs(3049));
    layer3_outputs(2755) <= not((layer2_outputs(822)) or (layer2_outputs(4741)));
    layer3_outputs(2756) <= layer2_outputs(808);
    layer3_outputs(2757) <= (layer2_outputs(329)) and (layer2_outputs(4510));
    layer3_outputs(2758) <= not((layer2_outputs(1744)) and (layer2_outputs(2064)));
    layer3_outputs(2759) <= layer2_outputs(5114);
    layer3_outputs(2760) <= '0';
    layer3_outputs(2761) <= not(layer2_outputs(4236));
    layer3_outputs(2762) <= (layer2_outputs(4203)) and not (layer2_outputs(1495));
    layer3_outputs(2763) <= not(layer2_outputs(289)) or (layer2_outputs(887));
    layer3_outputs(2764) <= '0';
    layer3_outputs(2765) <= not(layer2_outputs(565)) or (layer2_outputs(3881));
    layer3_outputs(2766) <= layer2_outputs(3466);
    layer3_outputs(2767) <= not(layer2_outputs(4477));
    layer3_outputs(2768) <= (layer2_outputs(2468)) and (layer2_outputs(591));
    layer3_outputs(2769) <= (layer2_outputs(547)) and (layer2_outputs(3319));
    layer3_outputs(2770) <= '1';
    layer3_outputs(2771) <= not(layer2_outputs(4394)) or (layer2_outputs(998));
    layer3_outputs(2772) <= '1';
    layer3_outputs(2773) <= (layer2_outputs(4682)) xor (layer2_outputs(4035));
    layer3_outputs(2774) <= '0';
    layer3_outputs(2775) <= not(layer2_outputs(3937)) or (layer2_outputs(3267));
    layer3_outputs(2776) <= not(layer2_outputs(4954));
    layer3_outputs(2777) <= not(layer2_outputs(4476));
    layer3_outputs(2778) <= not(layer2_outputs(487));
    layer3_outputs(2779) <= not(layer2_outputs(2018));
    layer3_outputs(2780) <= '1';
    layer3_outputs(2781) <= (layer2_outputs(1489)) xor (layer2_outputs(918));
    layer3_outputs(2782) <= layer2_outputs(189);
    layer3_outputs(2783) <= (layer2_outputs(3195)) and not (layer2_outputs(4149));
    layer3_outputs(2784) <= (layer2_outputs(299)) or (layer2_outputs(2404));
    layer3_outputs(2785) <= not(layer2_outputs(2490));
    layer3_outputs(2786) <= not(layer2_outputs(88));
    layer3_outputs(2787) <= (layer2_outputs(2295)) and not (layer2_outputs(3510));
    layer3_outputs(2788) <= not(layer2_outputs(173));
    layer3_outputs(2789) <= (layer2_outputs(930)) and (layer2_outputs(1604));
    layer3_outputs(2790) <= not(layer2_outputs(3295));
    layer3_outputs(2791) <= not((layer2_outputs(4096)) and (layer2_outputs(4156)));
    layer3_outputs(2792) <= not(layer2_outputs(4616));
    layer3_outputs(2793) <= layer2_outputs(895);
    layer3_outputs(2794) <= not(layer2_outputs(4374));
    layer3_outputs(2795) <= '0';
    layer3_outputs(2796) <= not((layer2_outputs(3385)) and (layer2_outputs(4)));
    layer3_outputs(2797) <= '0';
    layer3_outputs(2798) <= (layer2_outputs(1610)) and not (layer2_outputs(140));
    layer3_outputs(2799) <= not(layer2_outputs(5113));
    layer3_outputs(2800) <= (layer2_outputs(2341)) or (layer2_outputs(2550));
    layer3_outputs(2801) <= not(layer2_outputs(194)) or (layer2_outputs(3919));
    layer3_outputs(2802) <= not((layer2_outputs(3463)) xor (layer2_outputs(3880)));
    layer3_outputs(2803) <= (layer2_outputs(965)) or (layer2_outputs(4932));
    layer3_outputs(2804) <= (layer2_outputs(4831)) and (layer2_outputs(1907));
    layer3_outputs(2805) <= '1';
    layer3_outputs(2806) <= not(layer2_outputs(1831));
    layer3_outputs(2807) <= (layer2_outputs(4944)) or (layer2_outputs(596));
    layer3_outputs(2808) <= not((layer2_outputs(66)) and (layer2_outputs(595)));
    layer3_outputs(2809) <= not((layer2_outputs(3288)) and (layer2_outputs(120)));
    layer3_outputs(2810) <= not(layer2_outputs(2918));
    layer3_outputs(2811) <= layer2_outputs(4600);
    layer3_outputs(2812) <= layer2_outputs(85);
    layer3_outputs(2813) <= layer2_outputs(1958);
    layer3_outputs(2814) <= (layer2_outputs(1267)) or (layer2_outputs(3107));
    layer3_outputs(2815) <= '1';
    layer3_outputs(2816) <= '1';
    layer3_outputs(2817) <= (layer2_outputs(1037)) and (layer2_outputs(1131));
    layer3_outputs(2818) <= (layer2_outputs(504)) and not (layer2_outputs(2443));
    layer3_outputs(2819) <= (layer2_outputs(799)) or (layer2_outputs(1024));
    layer3_outputs(2820) <= not(layer2_outputs(3338)) or (layer2_outputs(2002));
    layer3_outputs(2821) <= layer2_outputs(4553);
    layer3_outputs(2822) <= layer2_outputs(773);
    layer3_outputs(2823) <= layer2_outputs(519);
    layer3_outputs(2824) <= layer2_outputs(4061);
    layer3_outputs(2825) <= (layer2_outputs(5075)) or (layer2_outputs(1852));
    layer3_outputs(2826) <= not((layer2_outputs(756)) or (layer2_outputs(497)));
    layer3_outputs(2827) <= not(layer2_outputs(708)) or (layer2_outputs(3940));
    layer3_outputs(2828) <= not(layer2_outputs(3471));
    layer3_outputs(2829) <= (layer2_outputs(1360)) and (layer2_outputs(3319));
    layer3_outputs(2830) <= layer2_outputs(2546);
    layer3_outputs(2831) <= not(layer2_outputs(3841));
    layer3_outputs(2832) <= '1';
    layer3_outputs(2833) <= layer2_outputs(4287);
    layer3_outputs(2834) <= not(layer2_outputs(919)) or (layer2_outputs(1847));
    layer3_outputs(2835) <= not(layer2_outputs(1267));
    layer3_outputs(2836) <= not(layer2_outputs(1963)) or (layer2_outputs(3686));
    layer3_outputs(2837) <= not((layer2_outputs(3796)) or (layer2_outputs(1592)));
    layer3_outputs(2838) <= not((layer2_outputs(1821)) or (layer2_outputs(1609)));
    layer3_outputs(2839) <= not(layer2_outputs(4361));
    layer3_outputs(2840) <= '0';
    layer3_outputs(2841) <= not(layer2_outputs(996));
    layer3_outputs(2842) <= '0';
    layer3_outputs(2843) <= not(layer2_outputs(2519));
    layer3_outputs(2844) <= layer2_outputs(4407);
    layer3_outputs(2845) <= not(layer2_outputs(3828));
    layer3_outputs(2846) <= not(layer2_outputs(4153)) or (layer2_outputs(847));
    layer3_outputs(2847) <= not((layer2_outputs(3589)) or (layer2_outputs(1022)));
    layer3_outputs(2848) <= '0';
    layer3_outputs(2849) <= '0';
    layer3_outputs(2850) <= (layer2_outputs(643)) or (layer2_outputs(104));
    layer3_outputs(2851) <= layer2_outputs(4845);
    layer3_outputs(2852) <= not((layer2_outputs(442)) xor (layer2_outputs(165)));
    layer3_outputs(2853) <= not(layer2_outputs(3011));
    layer3_outputs(2854) <= not(layer2_outputs(5021));
    layer3_outputs(2855) <= layer2_outputs(3088);
    layer3_outputs(2856) <= not(layer2_outputs(2998));
    layer3_outputs(2857) <= not(layer2_outputs(2590));
    layer3_outputs(2858) <= '1';
    layer3_outputs(2859) <= not((layer2_outputs(700)) and (layer2_outputs(3768)));
    layer3_outputs(2860) <= '0';
    layer3_outputs(2861) <= '0';
    layer3_outputs(2862) <= not(layer2_outputs(2483)) or (layer2_outputs(1403));
    layer3_outputs(2863) <= '0';
    layer3_outputs(2864) <= not((layer2_outputs(5038)) or (layer2_outputs(2899)));
    layer3_outputs(2865) <= '0';
    layer3_outputs(2866) <= not((layer2_outputs(2465)) or (layer2_outputs(1480)));
    layer3_outputs(2867) <= not(layer2_outputs(3179));
    layer3_outputs(2868) <= not(layer2_outputs(2641));
    layer3_outputs(2869) <= not(layer2_outputs(2730)) or (layer2_outputs(932));
    layer3_outputs(2870) <= not((layer2_outputs(2394)) or (layer2_outputs(3936)));
    layer3_outputs(2871) <= layer2_outputs(3861);
    layer3_outputs(2872) <= '1';
    layer3_outputs(2873) <= (layer2_outputs(3533)) or (layer2_outputs(923));
    layer3_outputs(2874) <= layer2_outputs(2027);
    layer3_outputs(2875) <= '0';
    layer3_outputs(2876) <= (layer2_outputs(798)) and (layer2_outputs(4653));
    layer3_outputs(2877) <= layer2_outputs(382);
    layer3_outputs(2878) <= (layer2_outputs(1538)) and not (layer2_outputs(1994));
    layer3_outputs(2879) <= not(layer2_outputs(3854));
    layer3_outputs(2880) <= (layer2_outputs(4251)) and not (layer2_outputs(4032));
    layer3_outputs(2881) <= not((layer2_outputs(1646)) and (layer2_outputs(1915)));
    layer3_outputs(2882) <= layer2_outputs(4813);
    layer3_outputs(2883) <= (layer2_outputs(3476)) and not (layer2_outputs(1842));
    layer3_outputs(2884) <= not((layer2_outputs(1821)) and (layer2_outputs(1478)));
    layer3_outputs(2885) <= not((layer2_outputs(1413)) and (layer2_outputs(3241)));
    layer3_outputs(2886) <= layer2_outputs(4406);
    layer3_outputs(2887) <= not(layer2_outputs(2072));
    layer3_outputs(2888) <= not(layer2_outputs(4035));
    layer3_outputs(2889) <= layer2_outputs(2242);
    layer3_outputs(2890) <= not((layer2_outputs(2512)) and (layer2_outputs(1653)));
    layer3_outputs(2891) <= (layer2_outputs(4201)) and (layer2_outputs(167));
    layer3_outputs(2892) <= '1';
    layer3_outputs(2893) <= layer2_outputs(4883);
    layer3_outputs(2894) <= not(layer2_outputs(1065)) or (layer2_outputs(4012));
    layer3_outputs(2895) <= not(layer2_outputs(5009));
    layer3_outputs(2896) <= '1';
    layer3_outputs(2897) <= not((layer2_outputs(1418)) and (layer2_outputs(3340)));
    layer3_outputs(2898) <= not(layer2_outputs(1698));
    layer3_outputs(2899) <= not(layer2_outputs(4736));
    layer3_outputs(2900) <= layer2_outputs(1310);
    layer3_outputs(2901) <= layer2_outputs(2562);
    layer3_outputs(2902) <= not(layer2_outputs(4335));
    layer3_outputs(2903) <= (layer2_outputs(2060)) or (layer2_outputs(243));
    layer3_outputs(2904) <= not(layer2_outputs(2758));
    layer3_outputs(2905) <= (layer2_outputs(5064)) and (layer2_outputs(4387));
    layer3_outputs(2906) <= layer2_outputs(3754);
    layer3_outputs(2907) <= not((layer2_outputs(3157)) and (layer2_outputs(1104)));
    layer3_outputs(2908) <= (layer2_outputs(847)) or (layer2_outputs(3147));
    layer3_outputs(2909) <= not(layer2_outputs(1257));
    layer3_outputs(2910) <= layer2_outputs(4139);
    layer3_outputs(2911) <= layer2_outputs(431);
    layer3_outputs(2912) <= (layer2_outputs(3954)) or (layer2_outputs(3376));
    layer3_outputs(2913) <= (layer2_outputs(2721)) and not (layer2_outputs(3739));
    layer3_outputs(2914) <= (layer2_outputs(1943)) and (layer2_outputs(19));
    layer3_outputs(2915) <= (layer2_outputs(1092)) and (layer2_outputs(2161));
    layer3_outputs(2916) <= not(layer2_outputs(96)) or (layer2_outputs(3150));
    layer3_outputs(2917) <= not((layer2_outputs(3851)) or (layer2_outputs(5082)));
    layer3_outputs(2918) <= layer2_outputs(195);
    layer3_outputs(2919) <= not(layer2_outputs(3696));
    layer3_outputs(2920) <= not(layer2_outputs(1335)) or (layer2_outputs(2117));
    layer3_outputs(2921) <= layer2_outputs(2688);
    layer3_outputs(2922) <= layer2_outputs(979);
    layer3_outputs(2923) <= (layer2_outputs(4780)) and (layer2_outputs(2056));
    layer3_outputs(2924) <= '0';
    layer3_outputs(2925) <= layer2_outputs(2067);
    layer3_outputs(2926) <= (layer2_outputs(1868)) xor (layer2_outputs(4554));
    layer3_outputs(2927) <= not(layer2_outputs(831));
    layer3_outputs(2928) <= layer2_outputs(472);
    layer3_outputs(2929) <= not(layer2_outputs(1018));
    layer3_outputs(2930) <= not(layer2_outputs(3465));
    layer3_outputs(2931) <= '0';
    layer3_outputs(2932) <= '0';
    layer3_outputs(2933) <= layer2_outputs(359);
    layer3_outputs(2934) <= layer2_outputs(4733);
    layer3_outputs(2935) <= (layer2_outputs(2787)) or (layer2_outputs(3082));
    layer3_outputs(2936) <= (layer2_outputs(352)) and not (layer2_outputs(508));
    layer3_outputs(2937) <= layer2_outputs(4803);
    layer3_outputs(2938) <= not(layer2_outputs(3218));
    layer3_outputs(2939) <= layer2_outputs(4912);
    layer3_outputs(2940) <= not(layer2_outputs(72));
    layer3_outputs(2941) <= layer2_outputs(646);
    layer3_outputs(2942) <= not(layer2_outputs(2497)) or (layer2_outputs(2502));
    layer3_outputs(2943) <= '1';
    layer3_outputs(2944) <= not(layer2_outputs(1106)) or (layer2_outputs(440));
    layer3_outputs(2945) <= (layer2_outputs(3784)) xor (layer2_outputs(5029));
    layer3_outputs(2946) <= (layer2_outputs(4660)) and not (layer2_outputs(2311));
    layer3_outputs(2947) <= (layer2_outputs(1971)) or (layer2_outputs(3965));
    layer3_outputs(2948) <= (layer2_outputs(4443)) or (layer2_outputs(3219));
    layer3_outputs(2949) <= (layer2_outputs(2307)) and not (layer2_outputs(2988));
    layer3_outputs(2950) <= layer2_outputs(2819);
    layer3_outputs(2951) <= layer2_outputs(374);
    layer3_outputs(2952) <= (layer2_outputs(2175)) and not (layer2_outputs(2418));
    layer3_outputs(2953) <= layer2_outputs(4812);
    layer3_outputs(2954) <= layer2_outputs(3439);
    layer3_outputs(2955) <= not(layer2_outputs(2460));
    layer3_outputs(2956) <= '1';
    layer3_outputs(2957) <= (layer2_outputs(3186)) and not (layer2_outputs(1720));
    layer3_outputs(2958) <= not(layer2_outputs(3037));
    layer3_outputs(2959) <= not(layer2_outputs(843));
    layer3_outputs(2960) <= not((layer2_outputs(769)) or (layer2_outputs(4846)));
    layer3_outputs(2961) <= layer2_outputs(2162);
    layer3_outputs(2962) <= (layer2_outputs(3226)) and (layer2_outputs(1992));
    layer3_outputs(2963) <= '1';
    layer3_outputs(2964) <= (layer2_outputs(20)) or (layer2_outputs(4810));
    layer3_outputs(2965) <= '0';
    layer3_outputs(2966) <= layer2_outputs(2428);
    layer3_outputs(2967) <= not(layer2_outputs(1183));
    layer3_outputs(2968) <= (layer2_outputs(1272)) and (layer2_outputs(1864));
    layer3_outputs(2969) <= not((layer2_outputs(4299)) and (layer2_outputs(4199)));
    layer3_outputs(2970) <= (layer2_outputs(4221)) and not (layer2_outputs(645));
    layer3_outputs(2971) <= (layer2_outputs(833)) or (layer2_outputs(2092));
    layer3_outputs(2972) <= not((layer2_outputs(730)) and (layer2_outputs(895)));
    layer3_outputs(2973) <= '0';
    layer3_outputs(2974) <= (layer2_outputs(2713)) and not (layer2_outputs(2839));
    layer3_outputs(2975) <= not((layer2_outputs(2403)) or (layer2_outputs(555)));
    layer3_outputs(2976) <= layer2_outputs(4154);
    layer3_outputs(2977) <= '1';
    layer3_outputs(2978) <= not(layer2_outputs(3036));
    layer3_outputs(2979) <= layer2_outputs(1220);
    layer3_outputs(2980) <= '1';
    layer3_outputs(2981) <= (layer2_outputs(3317)) and not (layer2_outputs(3920));
    layer3_outputs(2982) <= not(layer2_outputs(4188));
    layer3_outputs(2983) <= not(layer2_outputs(4720));
    layer3_outputs(2984) <= not(layer2_outputs(4362)) or (layer2_outputs(4352));
    layer3_outputs(2985) <= (layer2_outputs(2782)) and not (layer2_outputs(2753));
    layer3_outputs(2986) <= (layer2_outputs(1285)) and not (layer2_outputs(3232));
    layer3_outputs(2987) <= not(layer2_outputs(2074));
    layer3_outputs(2988) <= layer2_outputs(3825);
    layer3_outputs(2989) <= not((layer2_outputs(4099)) and (layer2_outputs(1960)));
    layer3_outputs(2990) <= '1';
    layer3_outputs(2991) <= not((layer2_outputs(4558)) and (layer2_outputs(1261)));
    layer3_outputs(2992) <= (layer2_outputs(893)) and not (layer2_outputs(2140));
    layer3_outputs(2993) <= not((layer2_outputs(4583)) or (layer2_outputs(2125)));
    layer3_outputs(2994) <= layer2_outputs(2003);
    layer3_outputs(2995) <= '1';
    layer3_outputs(2996) <= not(layer2_outputs(4371));
    layer3_outputs(2997) <= (layer2_outputs(190)) xor (layer2_outputs(1876));
    layer3_outputs(2998) <= layer2_outputs(914);
    layer3_outputs(2999) <= '1';
    layer3_outputs(3000) <= not(layer2_outputs(2209));
    layer3_outputs(3001) <= not(layer2_outputs(2197)) or (layer2_outputs(1334));
    layer3_outputs(3002) <= (layer2_outputs(237)) and (layer2_outputs(1730));
    layer3_outputs(3003) <= (layer2_outputs(4996)) and not (layer2_outputs(4859));
    layer3_outputs(3004) <= (layer2_outputs(4527)) or (layer2_outputs(967));
    layer3_outputs(3005) <= not((layer2_outputs(1137)) or (layer2_outputs(4115)));
    layer3_outputs(3006) <= '0';
    layer3_outputs(3007) <= layer2_outputs(117);
    layer3_outputs(3008) <= not(layer2_outputs(2419));
    layer3_outputs(3009) <= not((layer2_outputs(4982)) xor (layer2_outputs(4626)));
    layer3_outputs(3010) <= (layer2_outputs(1747)) and not (layer2_outputs(98));
    layer3_outputs(3011) <= (layer2_outputs(3656)) and not (layer2_outputs(5048));
    layer3_outputs(3012) <= (layer2_outputs(4769)) or (layer2_outputs(302));
    layer3_outputs(3013) <= not((layer2_outputs(2048)) or (layer2_outputs(4571)));
    layer3_outputs(3014) <= (layer2_outputs(4823)) and not (layer2_outputs(3878));
    layer3_outputs(3015) <= not(layer2_outputs(2512)) or (layer2_outputs(4414));
    layer3_outputs(3016) <= not(layer2_outputs(2606));
    layer3_outputs(3017) <= layer2_outputs(3594);
    layer3_outputs(3018) <= not((layer2_outputs(4562)) and (layer2_outputs(1281)));
    layer3_outputs(3019) <= layer2_outputs(4769);
    layer3_outputs(3020) <= not(layer2_outputs(5011));
    layer3_outputs(3021) <= not(layer2_outputs(2473));
    layer3_outputs(3022) <= not(layer2_outputs(4890)) or (layer2_outputs(3800));
    layer3_outputs(3023) <= not((layer2_outputs(4260)) and (layer2_outputs(152)));
    layer3_outputs(3024) <= not(layer2_outputs(4054));
    layer3_outputs(3025) <= (layer2_outputs(1533)) or (layer2_outputs(2547));
    layer3_outputs(3026) <= '0';
    layer3_outputs(3027) <= (layer2_outputs(1921)) and (layer2_outputs(1379));
    layer3_outputs(3028) <= layer2_outputs(1176);
    layer3_outputs(3029) <= layer2_outputs(3691);
    layer3_outputs(3030) <= '1';
    layer3_outputs(3031) <= layer2_outputs(2821);
    layer3_outputs(3032) <= (layer2_outputs(15)) xor (layer2_outputs(161));
    layer3_outputs(3033) <= (layer2_outputs(1978)) and not (layer2_outputs(3210));
    layer3_outputs(3034) <= not(layer2_outputs(2937));
    layer3_outputs(3035) <= (layer2_outputs(104)) and not (layer2_outputs(3056));
    layer3_outputs(3036) <= not(layer2_outputs(4129));
    layer3_outputs(3037) <= layer2_outputs(54);
    layer3_outputs(3038) <= '1';
    layer3_outputs(3039) <= (layer2_outputs(2805)) and (layer2_outputs(4525));
    layer3_outputs(3040) <= (layer2_outputs(4992)) and not (layer2_outputs(4156));
    layer3_outputs(3041) <= not(layer2_outputs(2291)) or (layer2_outputs(417));
    layer3_outputs(3042) <= not((layer2_outputs(2975)) or (layer2_outputs(4978)));
    layer3_outputs(3043) <= (layer2_outputs(3911)) or (layer2_outputs(1670));
    layer3_outputs(3044) <= layer2_outputs(2818);
    layer3_outputs(3045) <= not(layer2_outputs(1351)) or (layer2_outputs(3463));
    layer3_outputs(3046) <= not(layer2_outputs(1925));
    layer3_outputs(3047) <= not((layer2_outputs(459)) and (layer2_outputs(2723)));
    layer3_outputs(3048) <= not((layer2_outputs(2233)) or (layer2_outputs(1059)));
    layer3_outputs(3049) <= '1';
    layer3_outputs(3050) <= '1';
    layer3_outputs(3051) <= layer2_outputs(4154);
    layer3_outputs(3052) <= (layer2_outputs(322)) and not (layer2_outputs(3732));
    layer3_outputs(3053) <= layer2_outputs(1238);
    layer3_outputs(3054) <= not(layer2_outputs(247));
    layer3_outputs(3055) <= '0';
    layer3_outputs(3056) <= not(layer2_outputs(2313));
    layer3_outputs(3057) <= '0';
    layer3_outputs(3058) <= layer2_outputs(1146);
    layer3_outputs(3059) <= layer2_outputs(3854);
    layer3_outputs(3060) <= not(layer2_outputs(2628)) or (layer2_outputs(320));
    layer3_outputs(3061) <= not((layer2_outputs(1401)) and (layer2_outputs(1402)));
    layer3_outputs(3062) <= not(layer2_outputs(4630));
    layer3_outputs(3063) <= layer2_outputs(747);
    layer3_outputs(3064) <= not(layer2_outputs(3961));
    layer3_outputs(3065) <= not((layer2_outputs(4687)) or (layer2_outputs(4754)));
    layer3_outputs(3066) <= not(layer2_outputs(3545));
    layer3_outputs(3067) <= (layer2_outputs(934)) and not (layer2_outputs(810));
    layer3_outputs(3068) <= (layer2_outputs(3638)) and not (layer2_outputs(3415));
    layer3_outputs(3069) <= layer2_outputs(1327);
    layer3_outputs(3070) <= layer2_outputs(1802);
    layer3_outputs(3071) <= not(layer2_outputs(1542)) or (layer2_outputs(4875));
    layer3_outputs(3072) <= (layer2_outputs(1021)) xor (layer2_outputs(2285));
    layer3_outputs(3073) <= not((layer2_outputs(4212)) or (layer2_outputs(3893)));
    layer3_outputs(3074) <= layer2_outputs(2191);
    layer3_outputs(3075) <= not(layer2_outputs(22)) or (layer2_outputs(5035));
    layer3_outputs(3076) <= layer2_outputs(762);
    layer3_outputs(3077) <= not(layer2_outputs(560));
    layer3_outputs(3078) <= not((layer2_outputs(293)) or (layer2_outputs(1529)));
    layer3_outputs(3079) <= (layer2_outputs(150)) or (layer2_outputs(341));
    layer3_outputs(3080) <= not(layer2_outputs(3142));
    layer3_outputs(3081) <= not(layer2_outputs(5055));
    layer3_outputs(3082) <= (layer2_outputs(289)) and not (layer2_outputs(222));
    layer3_outputs(3083) <= layer2_outputs(4363);
    layer3_outputs(3084) <= not(layer2_outputs(4051));
    layer3_outputs(3085) <= not(layer2_outputs(2931));
    layer3_outputs(3086) <= not(layer2_outputs(682)) or (layer2_outputs(4235));
    layer3_outputs(3087) <= '1';
    layer3_outputs(3088) <= not(layer2_outputs(139));
    layer3_outputs(3089) <= (layer2_outputs(1036)) and (layer2_outputs(2771));
    layer3_outputs(3090) <= not(layer2_outputs(3414)) or (layer2_outputs(165));
    layer3_outputs(3091) <= layer2_outputs(3156);
    layer3_outputs(3092) <= layer2_outputs(4429);
    layer3_outputs(3093) <= (layer2_outputs(4585)) or (layer2_outputs(239));
    layer3_outputs(3094) <= (layer2_outputs(2963)) and not (layer2_outputs(782));
    layer3_outputs(3095) <= '1';
    layer3_outputs(3096) <= not((layer2_outputs(513)) or (layer2_outputs(1744)));
    layer3_outputs(3097) <= not((layer2_outputs(609)) and (layer2_outputs(3081)));
    layer3_outputs(3098) <= not((layer2_outputs(3336)) and (layer2_outputs(1252)));
    layer3_outputs(3099) <= '1';
    layer3_outputs(3100) <= not(layer2_outputs(1200));
    layer3_outputs(3101) <= not((layer2_outputs(2120)) and (layer2_outputs(3222)));
    layer3_outputs(3102) <= not(layer2_outputs(3958)) or (layer2_outputs(2449));
    layer3_outputs(3103) <= not(layer2_outputs(1577));
    layer3_outputs(3104) <= not(layer2_outputs(4709));
    layer3_outputs(3105) <= layer2_outputs(3034);
    layer3_outputs(3106) <= '1';
    layer3_outputs(3107) <= not((layer2_outputs(5050)) or (layer2_outputs(1051)));
    layer3_outputs(3108) <= '0';
    layer3_outputs(3109) <= (layer2_outputs(3071)) and not (layer2_outputs(3719));
    layer3_outputs(3110) <= layer2_outputs(3322);
    layer3_outputs(3111) <= (layer2_outputs(3452)) and not (layer2_outputs(4583));
    layer3_outputs(3112) <= not(layer2_outputs(2559));
    layer3_outputs(3113) <= not(layer2_outputs(3040));
    layer3_outputs(3114) <= (layer2_outputs(1003)) and not (layer2_outputs(4495));
    layer3_outputs(3115) <= (layer2_outputs(3290)) and not (layer2_outputs(4644));
    layer3_outputs(3116) <= not(layer2_outputs(1594));
    layer3_outputs(3117) <= not(layer2_outputs(662)) or (layer2_outputs(221));
    layer3_outputs(3118) <= not(layer2_outputs(2488)) or (layer2_outputs(1725));
    layer3_outputs(3119) <= (layer2_outputs(989)) and (layer2_outputs(3449));
    layer3_outputs(3120) <= not(layer2_outputs(5070));
    layer3_outputs(3121) <= (layer2_outputs(4993)) and (layer2_outputs(1622));
    layer3_outputs(3122) <= layer2_outputs(2229);
    layer3_outputs(3123) <= (layer2_outputs(609)) and (layer2_outputs(1979));
    layer3_outputs(3124) <= '1';
    layer3_outputs(3125) <= not((layer2_outputs(1193)) or (layer2_outputs(482)));
    layer3_outputs(3126) <= not(layer2_outputs(744));
    layer3_outputs(3127) <= '1';
    layer3_outputs(3128) <= layer2_outputs(2440);
    layer3_outputs(3129) <= not(layer2_outputs(1553)) or (layer2_outputs(4936));
    layer3_outputs(3130) <= (layer2_outputs(1621)) and not (layer2_outputs(3073));
    layer3_outputs(3131) <= '1';
    layer3_outputs(3132) <= (layer2_outputs(123)) and not (layer2_outputs(3424));
    layer3_outputs(3133) <= (layer2_outputs(4826)) and not (layer2_outputs(2783));
    layer3_outputs(3134) <= not(layer2_outputs(4539)) or (layer2_outputs(4635));
    layer3_outputs(3135) <= layer2_outputs(2454);
    layer3_outputs(3136) <= (layer2_outputs(3142)) or (layer2_outputs(4410));
    layer3_outputs(3137) <= layer2_outputs(1470);
    layer3_outputs(3138) <= layer2_outputs(1217);
    layer3_outputs(3139) <= not(layer2_outputs(2471)) or (layer2_outputs(3591));
    layer3_outputs(3140) <= (layer2_outputs(77)) or (layer2_outputs(1142));
    layer3_outputs(3141) <= not(layer2_outputs(3356));
    layer3_outputs(3142) <= '1';
    layer3_outputs(3143) <= not((layer2_outputs(837)) and (layer2_outputs(4437)));
    layer3_outputs(3144) <= layer2_outputs(740);
    layer3_outputs(3145) <= (layer2_outputs(4855)) and not (layer2_outputs(3988));
    layer3_outputs(3146) <= not((layer2_outputs(1858)) and (layer2_outputs(3037)));
    layer3_outputs(3147) <= (layer2_outputs(3010)) and not (layer2_outputs(3435));
    layer3_outputs(3148) <= (layer2_outputs(3738)) or (layer2_outputs(4955));
    layer3_outputs(3149) <= (layer2_outputs(454)) and not (layer2_outputs(1500));
    layer3_outputs(3150) <= layer2_outputs(3330);
    layer3_outputs(3151) <= (layer2_outputs(3982)) and not (layer2_outputs(2365));
    layer3_outputs(3152) <= '0';
    layer3_outputs(3153) <= '0';
    layer3_outputs(3154) <= not((layer2_outputs(5003)) or (layer2_outputs(2744)));
    layer3_outputs(3155) <= not((layer2_outputs(2919)) or (layer2_outputs(51)));
    layer3_outputs(3156) <= layer2_outputs(3660);
    layer3_outputs(3157) <= (layer2_outputs(2379)) and not (layer2_outputs(2623));
    layer3_outputs(3158) <= layer2_outputs(2053);
    layer3_outputs(3159) <= not(layer2_outputs(439));
    layer3_outputs(3160) <= (layer2_outputs(3962)) and (layer2_outputs(2959));
    layer3_outputs(3161) <= '1';
    layer3_outputs(3162) <= layer2_outputs(1964);
    layer3_outputs(3163) <= layer2_outputs(1258);
    layer3_outputs(3164) <= not((layer2_outputs(3564)) or (layer2_outputs(529)));
    layer3_outputs(3165) <= not(layer2_outputs(3357));
    layer3_outputs(3166) <= layer2_outputs(2446);
    layer3_outputs(3167) <= not(layer2_outputs(3648)) or (layer2_outputs(1616));
    layer3_outputs(3168) <= not(layer2_outputs(147));
    layer3_outputs(3169) <= layer2_outputs(494);
    layer3_outputs(3170) <= (layer2_outputs(713)) and not (layer2_outputs(1034));
    layer3_outputs(3171) <= '0';
    layer3_outputs(3172) <= not((layer2_outputs(106)) and (layer2_outputs(2647)));
    layer3_outputs(3173) <= not((layer2_outputs(3993)) or (layer2_outputs(4350)));
    layer3_outputs(3174) <= (layer2_outputs(1515)) and not (layer2_outputs(1825));
    layer3_outputs(3175) <= (layer2_outputs(3671)) and not (layer2_outputs(1908));
    layer3_outputs(3176) <= (layer2_outputs(918)) and not (layer2_outputs(3714));
    layer3_outputs(3177) <= (layer2_outputs(1328)) and not (layer2_outputs(2659));
    layer3_outputs(3178) <= not((layer2_outputs(3339)) or (layer2_outputs(1488)));
    layer3_outputs(3179) <= not((layer2_outputs(4215)) and (layer2_outputs(4211)));
    layer3_outputs(3180) <= not(layer2_outputs(484));
    layer3_outputs(3181) <= not(layer2_outputs(4886));
    layer3_outputs(3182) <= not(layer2_outputs(4758));
    layer3_outputs(3183) <= not(layer2_outputs(1823)) or (layer2_outputs(3732));
    layer3_outputs(3184) <= not(layer2_outputs(1844)) or (layer2_outputs(4774));
    layer3_outputs(3185) <= not(layer2_outputs(1991));
    layer3_outputs(3186) <= not(layer2_outputs(3288));
    layer3_outputs(3187) <= not(layer2_outputs(4351));
    layer3_outputs(3188) <= layer2_outputs(253);
    layer3_outputs(3189) <= not(layer2_outputs(3364));
    layer3_outputs(3190) <= not(layer2_outputs(3721));
    layer3_outputs(3191) <= not((layer2_outputs(2154)) or (layer2_outputs(1064)));
    layer3_outputs(3192) <= not(layer2_outputs(4135));
    layer3_outputs(3193) <= '0';
    layer3_outputs(3194) <= (layer2_outputs(2966)) and not (layer2_outputs(2144));
    layer3_outputs(3195) <= not(layer2_outputs(1789)) or (layer2_outputs(1549));
    layer3_outputs(3196) <= not((layer2_outputs(528)) or (layer2_outputs(968)));
    layer3_outputs(3197) <= layer2_outputs(4404);
    layer3_outputs(3198) <= not(layer2_outputs(2912));
    layer3_outputs(3199) <= not((layer2_outputs(2017)) or (layer2_outputs(2613)));
    layer3_outputs(3200) <= not(layer2_outputs(3512));
    layer3_outputs(3201) <= layer2_outputs(2180);
    layer3_outputs(3202) <= not(layer2_outputs(1069));
    layer3_outputs(3203) <= not(layer2_outputs(4231));
    layer3_outputs(3204) <= not((layer2_outputs(3890)) or (layer2_outputs(3048)));
    layer3_outputs(3205) <= '1';
    layer3_outputs(3206) <= not(layer2_outputs(2392));
    layer3_outputs(3207) <= not((layer2_outputs(1678)) and (layer2_outputs(3255)));
    layer3_outputs(3208) <= not((layer2_outputs(2318)) and (layer2_outputs(958)));
    layer3_outputs(3209) <= '0';
    layer3_outputs(3210) <= not((layer2_outputs(2082)) or (layer2_outputs(1668)));
    layer3_outputs(3211) <= not(layer2_outputs(3735));
    layer3_outputs(3212) <= (layer2_outputs(925)) and not (layer2_outputs(3053));
    layer3_outputs(3213) <= not(layer2_outputs(5069));
    layer3_outputs(3214) <= (layer2_outputs(4776)) or (layer2_outputs(2591));
    layer3_outputs(3215) <= layer2_outputs(2905);
    layer3_outputs(3216) <= not(layer2_outputs(1096));
    layer3_outputs(3217) <= not(layer2_outputs(1235));
    layer3_outputs(3218) <= '1';
    layer3_outputs(3219) <= layer2_outputs(1239);
    layer3_outputs(3220) <= (layer2_outputs(4824)) and not (layer2_outputs(3423));
    layer3_outputs(3221) <= not(layer2_outputs(3829));
    layer3_outputs(3222) <= not(layer2_outputs(4910));
    layer3_outputs(3223) <= (layer2_outputs(4412)) and not (layer2_outputs(3558));
    layer3_outputs(3224) <= not(layer2_outputs(3481));
    layer3_outputs(3225) <= '0';
    layer3_outputs(3226) <= not((layer2_outputs(4093)) and (layer2_outputs(427)));
    layer3_outputs(3227) <= layer2_outputs(4080);
    layer3_outputs(3228) <= not(layer2_outputs(4258));
    layer3_outputs(3229) <= not(layer2_outputs(4219)) or (layer2_outputs(1297));
    layer3_outputs(3230) <= layer2_outputs(3216);
    layer3_outputs(3231) <= not((layer2_outputs(2977)) or (layer2_outputs(2783)));
    layer3_outputs(3232) <= not(layer2_outputs(3686));
    layer3_outputs(3233) <= not((layer2_outputs(1972)) and (layer2_outputs(625)));
    layer3_outputs(3234) <= (layer2_outputs(1103)) xor (layer2_outputs(149));
    layer3_outputs(3235) <= (layer2_outputs(3921)) and not (layer2_outputs(5110));
    layer3_outputs(3236) <= not((layer2_outputs(3380)) xor (layer2_outputs(4367)));
    layer3_outputs(3237) <= layer2_outputs(4332);
    layer3_outputs(3238) <= (layer2_outputs(2520)) or (layer2_outputs(29));
    layer3_outputs(3239) <= not(layer2_outputs(3960));
    layer3_outputs(3240) <= (layer2_outputs(724)) or (layer2_outputs(3089));
    layer3_outputs(3241) <= not((layer2_outputs(1735)) xor (layer2_outputs(2171)));
    layer3_outputs(3242) <= (layer2_outputs(1447)) and not (layer2_outputs(2945));
    layer3_outputs(3243) <= not(layer2_outputs(5079)) or (layer2_outputs(3332));
    layer3_outputs(3244) <= '1';
    layer3_outputs(3245) <= '0';
    layer3_outputs(3246) <= not(layer2_outputs(3496));
    layer3_outputs(3247) <= not((layer2_outputs(4520)) and (layer2_outputs(757)));
    layer3_outputs(3248) <= not(layer2_outputs(4914));
    layer3_outputs(3249) <= '1';
    layer3_outputs(3250) <= not(layer2_outputs(4347));
    layer3_outputs(3251) <= (layer2_outputs(3731)) or (layer2_outputs(2331));
    layer3_outputs(3252) <= '1';
    layer3_outputs(3253) <= layer2_outputs(283);
    layer3_outputs(3254) <= not(layer2_outputs(3052));
    layer3_outputs(3255) <= not(layer2_outputs(3209));
    layer3_outputs(3256) <= not((layer2_outputs(1354)) and (layer2_outputs(3204)));
    layer3_outputs(3257) <= not((layer2_outputs(1047)) and (layer2_outputs(3645)));
    layer3_outputs(3258) <= not((layer2_outputs(407)) or (layer2_outputs(2775)));
    layer3_outputs(3259) <= not(layer2_outputs(3117)) or (layer2_outputs(1445));
    layer3_outputs(3260) <= '0';
    layer3_outputs(3261) <= (layer2_outputs(1689)) and not (layer2_outputs(4778));
    layer3_outputs(3262) <= '1';
    layer3_outputs(3263) <= (layer2_outputs(1097)) and not (layer2_outputs(4377));
    layer3_outputs(3264) <= '1';
    layer3_outputs(3265) <= '1';
    layer3_outputs(3266) <= not(layer2_outputs(5093));
    layer3_outputs(3267) <= not(layer2_outputs(4722));
    layer3_outputs(3268) <= not(layer2_outputs(4935));
    layer3_outputs(3269) <= not(layer2_outputs(2549)) or (layer2_outputs(5025));
    layer3_outputs(3270) <= not(layer2_outputs(4607));
    layer3_outputs(3271) <= not(layer2_outputs(1073)) or (layer2_outputs(3246));
    layer3_outputs(3272) <= '0';
    layer3_outputs(3273) <= layer2_outputs(1392);
    layer3_outputs(3274) <= not((layer2_outputs(674)) and (layer2_outputs(4391)));
    layer3_outputs(3275) <= (layer2_outputs(4217)) and not (layer2_outputs(4940));
    layer3_outputs(3276) <= layer2_outputs(2407);
    layer3_outputs(3277) <= not(layer2_outputs(5061)) or (layer2_outputs(3657));
    layer3_outputs(3278) <= not(layer2_outputs(1120));
    layer3_outputs(3279) <= not(layer2_outputs(3242));
    layer3_outputs(3280) <= not(layer2_outputs(2543)) or (layer2_outputs(1070));
    layer3_outputs(3281) <= not((layer2_outputs(643)) or (layer2_outputs(4843)));
    layer3_outputs(3282) <= not(layer2_outputs(976));
    layer3_outputs(3283) <= (layer2_outputs(2345)) and not (layer2_outputs(2219));
    layer3_outputs(3284) <= not(layer2_outputs(3275));
    layer3_outputs(3285) <= layer2_outputs(2184);
    layer3_outputs(3286) <= (layer2_outputs(102)) and not (layer2_outputs(4490));
    layer3_outputs(3287) <= (layer2_outputs(3713)) and (layer2_outputs(657));
    layer3_outputs(3288) <= not(layer2_outputs(4277));
    layer3_outputs(3289) <= '0';
    layer3_outputs(3290) <= layer2_outputs(4179);
    layer3_outputs(3291) <= layer2_outputs(1841);
    layer3_outputs(3292) <= not(layer2_outputs(4507)) or (layer2_outputs(4573));
    layer3_outputs(3293) <= (layer2_outputs(1368)) and (layer2_outputs(838));
    layer3_outputs(3294) <= not(layer2_outputs(3112)) or (layer2_outputs(4270));
    layer3_outputs(3295) <= not((layer2_outputs(1396)) or (layer2_outputs(896)));
    layer3_outputs(3296) <= (layer2_outputs(2913)) or (layer2_outputs(58));
    layer3_outputs(3297) <= not(layer2_outputs(2049));
    layer3_outputs(3298) <= not(layer2_outputs(2031));
    layer3_outputs(3299) <= layer2_outputs(2363);
    layer3_outputs(3300) <= layer2_outputs(461);
    layer3_outputs(3301) <= not(layer2_outputs(5001));
    layer3_outputs(3302) <= layer2_outputs(3);
    layer3_outputs(3303) <= not(layer2_outputs(782));
    layer3_outputs(3304) <= '1';
    layer3_outputs(3305) <= not(layer2_outputs(883)) or (layer2_outputs(3115));
    layer3_outputs(3306) <= layer2_outputs(4283);
    layer3_outputs(3307) <= layer2_outputs(4602);
    layer3_outputs(3308) <= not(layer2_outputs(1408)) or (layer2_outputs(2322));
    layer3_outputs(3309) <= (layer2_outputs(1072)) and (layer2_outputs(122));
    layer3_outputs(3310) <= not((layer2_outputs(1741)) or (layer2_outputs(4228)));
    layer3_outputs(3311) <= not(layer2_outputs(2147));
    layer3_outputs(3312) <= not(layer2_outputs(651));
    layer3_outputs(3313) <= layer2_outputs(4401);
    layer3_outputs(3314) <= not(layer2_outputs(1000));
    layer3_outputs(3315) <= layer2_outputs(2242);
    layer3_outputs(3316) <= (layer2_outputs(4957)) and not (layer2_outputs(1952));
    layer3_outputs(3317) <= (layer2_outputs(3111)) and not (layer2_outputs(4503));
    layer3_outputs(3318) <= (layer2_outputs(4138)) or (layer2_outputs(70));
    layer3_outputs(3319) <= (layer2_outputs(934)) and (layer2_outputs(3292));
    layer3_outputs(3320) <= (layer2_outputs(4690)) and not (layer2_outputs(4885));
    layer3_outputs(3321) <= not(layer2_outputs(2085));
    layer3_outputs(3322) <= '1';
    layer3_outputs(3323) <= not(layer2_outputs(211));
    layer3_outputs(3324) <= (layer2_outputs(2664)) or (layer2_outputs(2135));
    layer3_outputs(3325) <= layer2_outputs(849);
    layer3_outputs(3326) <= not(layer2_outputs(1544)) or (layer2_outputs(3062));
    layer3_outputs(3327) <= layer2_outputs(689);
    layer3_outputs(3328) <= layer2_outputs(1473);
    layer3_outputs(3329) <= (layer2_outputs(2831)) and (layer2_outputs(4440));
    layer3_outputs(3330) <= not(layer2_outputs(4487)) or (layer2_outputs(3907));
    layer3_outputs(3331) <= (layer2_outputs(748)) and not (layer2_outputs(2748));
    layer3_outputs(3332) <= not(layer2_outputs(3636));
    layer3_outputs(3333) <= not(layer2_outputs(1485));
    layer3_outputs(3334) <= not(layer2_outputs(2077));
    layer3_outputs(3335) <= layer2_outputs(5004);
    layer3_outputs(3336) <= not((layer2_outputs(4521)) or (layer2_outputs(1505)));
    layer3_outputs(3337) <= (layer2_outputs(180)) and not (layer2_outputs(3567));
    layer3_outputs(3338) <= not((layer2_outputs(3066)) and (layer2_outputs(1717)));
    layer3_outputs(3339) <= not(layer2_outputs(3442)) or (layer2_outputs(4818));
    layer3_outputs(3340) <= not(layer2_outputs(1672));
    layer3_outputs(3341) <= (layer2_outputs(1572)) and not (layer2_outputs(4051));
    layer3_outputs(3342) <= not(layer2_outputs(5110)) or (layer2_outputs(3093));
    layer3_outputs(3343) <= not(layer2_outputs(983));
    layer3_outputs(3344) <= layer2_outputs(1071);
    layer3_outputs(3345) <= '1';
    layer3_outputs(3346) <= layer2_outputs(4516);
    layer3_outputs(3347) <= layer2_outputs(2317);
    layer3_outputs(3348) <= '1';
    layer3_outputs(3349) <= (layer2_outputs(3682)) xor (layer2_outputs(3957));
    layer3_outputs(3350) <= not(layer2_outputs(4814));
    layer3_outputs(3351) <= not(layer2_outputs(3339));
    layer3_outputs(3352) <= not(layer2_outputs(1085)) or (layer2_outputs(311));
    layer3_outputs(3353) <= not(layer2_outputs(2656));
    layer3_outputs(3354) <= not(layer2_outputs(980));
    layer3_outputs(3355) <= '1';
    layer3_outputs(3356) <= (layer2_outputs(3552)) and not (layer2_outputs(4325));
    layer3_outputs(3357) <= layer2_outputs(4058);
    layer3_outputs(3358) <= (layer2_outputs(2235)) or (layer2_outputs(471));
    layer3_outputs(3359) <= (layer2_outputs(4618)) and not (layer2_outputs(4677));
    layer3_outputs(3360) <= not(layer2_outputs(3795));
    layer3_outputs(3361) <= '0';
    layer3_outputs(3362) <= '0';
    layer3_outputs(3363) <= not((layer2_outputs(2716)) and (layer2_outputs(1164)));
    layer3_outputs(3364) <= not(layer2_outputs(1501)) or (layer2_outputs(769));
    layer3_outputs(3365) <= not(layer2_outputs(1228));
    layer3_outputs(3366) <= not(layer2_outputs(2635)) or (layer2_outputs(4068));
    layer3_outputs(3367) <= layer2_outputs(677);
    layer3_outputs(3368) <= not(layer2_outputs(746)) or (layer2_outputs(2503));
    layer3_outputs(3369) <= not(layer2_outputs(1240)) or (layer2_outputs(5111));
    layer3_outputs(3370) <= '0';
    layer3_outputs(3371) <= (layer2_outputs(2616)) or (layer2_outputs(3869));
    layer3_outputs(3372) <= '1';
    layer3_outputs(3373) <= '1';
    layer3_outputs(3374) <= (layer2_outputs(4630)) and not (layer2_outputs(4531));
    layer3_outputs(3375) <= not((layer2_outputs(4907)) and (layer2_outputs(2068)));
    layer3_outputs(3376) <= (layer2_outputs(742)) and not (layer2_outputs(321));
    layer3_outputs(3377) <= (layer2_outputs(4488)) xor (layer2_outputs(2327));
    layer3_outputs(3378) <= not(layer2_outputs(2992));
    layer3_outputs(3379) <= not((layer2_outputs(4110)) or (layer2_outputs(532)));
    layer3_outputs(3380) <= not(layer2_outputs(4082)) or (layer2_outputs(2177));
    layer3_outputs(3381) <= not(layer2_outputs(4435));
    layer3_outputs(3382) <= layer2_outputs(3139);
    layer3_outputs(3383) <= (layer2_outputs(2921)) and not (layer2_outputs(4373));
    layer3_outputs(3384) <= (layer2_outputs(3633)) and not (layer2_outputs(2386));
    layer3_outputs(3385) <= not(layer2_outputs(4020));
    layer3_outputs(3386) <= not(layer2_outputs(2693)) or (layer2_outputs(3080));
    layer3_outputs(3387) <= '0';
    layer3_outputs(3388) <= '0';
    layer3_outputs(3389) <= (layer2_outputs(1697)) and (layer2_outputs(1380));
    layer3_outputs(3390) <= not((layer2_outputs(4552)) and (layer2_outputs(219)));
    layer3_outputs(3391) <= layer2_outputs(4227);
    layer3_outputs(3392) <= not(layer2_outputs(2226));
    layer3_outputs(3393) <= layer2_outputs(5071);
    layer3_outputs(3394) <= not((layer2_outputs(2411)) or (layer2_outputs(4393)));
    layer3_outputs(3395) <= layer2_outputs(2588);
    layer3_outputs(3396) <= '1';
    layer3_outputs(3397) <= not(layer2_outputs(3003));
    layer3_outputs(3398) <= layer2_outputs(586);
    layer3_outputs(3399) <= not(layer2_outputs(3948));
    layer3_outputs(3400) <= not(layer2_outputs(4233));
    layer3_outputs(3401) <= not((layer2_outputs(3197)) and (layer2_outputs(4130)));
    layer3_outputs(3402) <= not(layer2_outputs(2038));
    layer3_outputs(3403) <= '0';
    layer3_outputs(3404) <= '0';
    layer3_outputs(3405) <= not((layer2_outputs(1174)) or (layer2_outputs(474)));
    layer3_outputs(3406) <= not(layer2_outputs(4099)) or (layer2_outputs(2028));
    layer3_outputs(3407) <= layer2_outputs(2793);
    layer3_outputs(3408) <= layer2_outputs(3400);
    layer3_outputs(3409) <= '0';
    layer3_outputs(3410) <= layer2_outputs(3098);
    layer3_outputs(3411) <= not((layer2_outputs(2882)) xor (layer2_outputs(3187)));
    layer3_outputs(3412) <= (layer2_outputs(4774)) and not (layer2_outputs(3582));
    layer3_outputs(3413) <= not(layer2_outputs(4084)) or (layer2_outputs(1764));
    layer3_outputs(3414) <= not(layer2_outputs(2724));
    layer3_outputs(3415) <= layer2_outputs(516);
    layer3_outputs(3416) <= (layer2_outputs(4548)) and (layer2_outputs(821));
    layer3_outputs(3417) <= (layer2_outputs(1949)) and not (layer2_outputs(2661));
    layer3_outputs(3418) <= (layer2_outputs(1292)) xor (layer2_outputs(452));
    layer3_outputs(3419) <= '1';
    layer3_outputs(3420) <= layer2_outputs(2060);
    layer3_outputs(3421) <= not(layer2_outputs(4776));
    layer3_outputs(3422) <= '0';
    layer3_outputs(3423) <= (layer2_outputs(379)) or (layer2_outputs(3812));
    layer3_outputs(3424) <= layer2_outputs(20);
    layer3_outputs(3425) <= not(layer2_outputs(1048)) or (layer2_outputs(3872));
    layer3_outputs(3426) <= not((layer2_outputs(3550)) and (layer2_outputs(1008)));
    layer3_outputs(3427) <= (layer2_outputs(1495)) and (layer2_outputs(70));
    layer3_outputs(3428) <= '0';
    layer3_outputs(3429) <= (layer2_outputs(1382)) or (layer2_outputs(1170));
    layer3_outputs(3430) <= (layer2_outputs(2409)) xor (layer2_outputs(1216));
    layer3_outputs(3431) <= (layer2_outputs(2719)) or (layer2_outputs(3905));
    layer3_outputs(3432) <= not((layer2_outputs(4118)) and (layer2_outputs(1829)));
    layer3_outputs(3433) <= '1';
    layer3_outputs(3434) <= (layer2_outputs(3324)) and not (layer2_outputs(1286));
    layer3_outputs(3435) <= not(layer2_outputs(183));
    layer3_outputs(3436) <= not((layer2_outputs(3949)) xor (layer2_outputs(995)));
    layer3_outputs(3437) <= (layer2_outputs(520)) and (layer2_outputs(577));
    layer3_outputs(3438) <= (layer2_outputs(1851)) and (layer2_outputs(1923));
    layer3_outputs(3439) <= not(layer2_outputs(3089));
    layer3_outputs(3440) <= (layer2_outputs(4507)) and not (layer2_outputs(4235));
    layer3_outputs(3441) <= not(layer2_outputs(2850));
    layer3_outputs(3442) <= layer2_outputs(1383);
    layer3_outputs(3443) <= not((layer2_outputs(3328)) and (layer2_outputs(3673)));
    layer3_outputs(3444) <= not((layer2_outputs(3461)) and (layer2_outputs(1943)));
    layer3_outputs(3445) <= not(layer2_outputs(1810));
    layer3_outputs(3446) <= not(layer2_outputs(3785));
    layer3_outputs(3447) <= not((layer2_outputs(3642)) and (layer2_outputs(3529)));
    layer3_outputs(3448) <= not(layer2_outputs(1410));
    layer3_outputs(3449) <= (layer2_outputs(453)) and (layer2_outputs(3582));
    layer3_outputs(3450) <= (layer2_outputs(4009)) and (layer2_outputs(940));
    layer3_outputs(3451) <= (layer2_outputs(3760)) xor (layer2_outputs(1068));
    layer3_outputs(3452) <= (layer2_outputs(418)) and not (layer2_outputs(2687));
    layer3_outputs(3453) <= not(layer2_outputs(4488)) or (layer2_outputs(1411));
    layer3_outputs(3454) <= (layer2_outputs(3945)) xor (layer2_outputs(2774));
    layer3_outputs(3455) <= not(layer2_outputs(2751));
    layer3_outputs(3456) <= layer2_outputs(3318);
    layer3_outputs(3457) <= (layer2_outputs(3383)) and (layer2_outputs(1887));
    layer3_outputs(3458) <= '1';
    layer3_outputs(3459) <= not(layer2_outputs(2903));
    layer3_outputs(3460) <= '1';
    layer3_outputs(3461) <= layer2_outputs(39);
    layer3_outputs(3462) <= not(layer2_outputs(956));
    layer3_outputs(3463) <= (layer2_outputs(1393)) and (layer2_outputs(2183));
    layer3_outputs(3464) <= not((layer2_outputs(1544)) xor (layer2_outputs(3472)));
    layer3_outputs(3465) <= '1';
    layer3_outputs(3466) <= (layer2_outputs(1596)) and not (layer2_outputs(1677));
    layer3_outputs(3467) <= not((layer2_outputs(2448)) and (layer2_outputs(4024)));
    layer3_outputs(3468) <= not(layer2_outputs(3914));
    layer3_outputs(3469) <= layer2_outputs(1417);
    layer3_outputs(3470) <= not((layer2_outputs(4665)) or (layer2_outputs(3125)));
    layer3_outputs(3471) <= not(layer2_outputs(4354));
    layer3_outputs(3472) <= not(layer2_outputs(4069)) or (layer2_outputs(2110));
    layer3_outputs(3473) <= not(layer2_outputs(3663));
    layer3_outputs(3474) <= (layer2_outputs(44)) xor (layer2_outputs(280));
    layer3_outputs(3475) <= (layer2_outputs(1834)) and (layer2_outputs(2202));
    layer3_outputs(3476) <= not(layer2_outputs(3284));
    layer3_outputs(3477) <= not((layer2_outputs(3809)) or (layer2_outputs(3191)));
    layer3_outputs(3478) <= '1';
    layer3_outputs(3479) <= not(layer2_outputs(5010));
    layer3_outputs(3480) <= not(layer2_outputs(2531));
    layer3_outputs(3481) <= (layer2_outputs(1048)) and not (layer2_outputs(64));
    layer3_outputs(3482) <= layer2_outputs(2127);
    layer3_outputs(3483) <= (layer2_outputs(1109)) and not (layer2_outputs(4839));
    layer3_outputs(3484) <= not(layer2_outputs(4165)) or (layer2_outputs(3690));
    layer3_outputs(3485) <= not(layer2_outputs(2039));
    layer3_outputs(3486) <= (layer2_outputs(212)) and not (layer2_outputs(3519));
    layer3_outputs(3487) <= not(layer2_outputs(5025));
    layer3_outputs(3488) <= (layer2_outputs(145)) and not (layer2_outputs(2269));
    layer3_outputs(3489) <= not(layer2_outputs(1843));
    layer3_outputs(3490) <= (layer2_outputs(2784)) and (layer2_outputs(2326));
    layer3_outputs(3491) <= (layer2_outputs(492)) or (layer2_outputs(2203));
    layer3_outputs(3492) <= not(layer2_outputs(4902));
    layer3_outputs(3493) <= not(layer2_outputs(4016)) or (layer2_outputs(4025));
    layer3_outputs(3494) <= '0';
    layer3_outputs(3495) <= (layer2_outputs(4196)) and not (layer2_outputs(4847));
    layer3_outputs(3496) <= layer2_outputs(1731);
    layer3_outputs(3497) <= not(layer2_outputs(385));
    layer3_outputs(3498) <= (layer2_outputs(4369)) and not (layer2_outputs(3896));
    layer3_outputs(3499) <= not(layer2_outputs(2661)) or (layer2_outputs(1028));
    layer3_outputs(3500) <= '0';
    layer3_outputs(3501) <= not(layer2_outputs(1314)) or (layer2_outputs(305));
    layer3_outputs(3502) <= layer2_outputs(3148);
    layer3_outputs(3503) <= layer2_outputs(2227);
    layer3_outputs(3504) <= not(layer2_outputs(3842));
    layer3_outputs(3505) <= layer2_outputs(1816);
    layer3_outputs(3506) <= (layer2_outputs(3912)) xor (layer2_outputs(3315));
    layer3_outputs(3507) <= not((layer2_outputs(3845)) and (layer2_outputs(1185)));
    layer3_outputs(3508) <= not(layer2_outputs(2019)) or (layer2_outputs(4256));
    layer3_outputs(3509) <= layer2_outputs(4173);
    layer3_outputs(3510) <= not((layer2_outputs(3206)) and (layer2_outputs(4618)));
    layer3_outputs(3511) <= not(layer2_outputs(2211));
    layer3_outputs(3512) <= (layer2_outputs(661)) or (layer2_outputs(806));
    layer3_outputs(3513) <= not(layer2_outputs(3366)) or (layer2_outputs(2213));
    layer3_outputs(3514) <= not((layer2_outputs(164)) and (layer2_outputs(4945)));
    layer3_outputs(3515) <= not((layer2_outputs(4605)) or (layer2_outputs(2006)));
    layer3_outputs(3516) <= not(layer2_outputs(551)) or (layer2_outputs(964));
    layer3_outputs(3517) <= not((layer2_outputs(444)) and (layer2_outputs(3113)));
    layer3_outputs(3518) <= '0';
    layer3_outputs(3519) <= layer2_outputs(4034);
    layer3_outputs(3520) <= '1';
    layer3_outputs(3521) <= '1';
    layer3_outputs(3522) <= not(layer2_outputs(3872));
    layer3_outputs(3523) <= (layer2_outputs(1661)) or (layer2_outputs(1595));
    layer3_outputs(3524) <= (layer2_outputs(4664)) xor (layer2_outputs(4380));
    layer3_outputs(3525) <= (layer2_outputs(2642)) and (layer2_outputs(5071));
    layer3_outputs(3526) <= not((layer2_outputs(3173)) or (layer2_outputs(3221)));
    layer3_outputs(3527) <= not(layer2_outputs(3296)) or (layer2_outputs(1362));
    layer3_outputs(3528) <= '0';
    layer3_outputs(3529) <= not(layer2_outputs(1422));
    layer3_outputs(3530) <= not((layer2_outputs(4534)) or (layer2_outputs(455)));
    layer3_outputs(3531) <= layer2_outputs(2343);
    layer3_outputs(3532) <= not((layer2_outputs(4895)) or (layer2_outputs(4905)));
    layer3_outputs(3533) <= not(layer2_outputs(266));
    layer3_outputs(3534) <= (layer2_outputs(207)) or (layer2_outputs(1183));
    layer3_outputs(3535) <= not((layer2_outputs(2929)) and (layer2_outputs(3103)));
    layer3_outputs(3536) <= not((layer2_outputs(1865)) xor (layer2_outputs(3230)));
    layer3_outputs(3537) <= not(layer2_outputs(248)) or (layer2_outputs(1568));
    layer3_outputs(3538) <= layer2_outputs(3627);
    layer3_outputs(3539) <= not((layer2_outputs(3509)) or (layer2_outputs(1530)));
    layer3_outputs(3540) <= layer2_outputs(4664);
    layer3_outputs(3541) <= (layer2_outputs(3847)) and (layer2_outputs(2851));
    layer3_outputs(3542) <= '0';
    layer3_outputs(3543) <= not(layer2_outputs(4433));
    layer3_outputs(3544) <= (layer2_outputs(598)) and not (layer2_outputs(3325));
    layer3_outputs(3545) <= not(layer2_outputs(2312));
    layer3_outputs(3546) <= not(layer2_outputs(2787));
    layer3_outputs(3547) <= not((layer2_outputs(1164)) xor (layer2_outputs(3770)));
    layer3_outputs(3548) <= (layer2_outputs(704)) and not (layer2_outputs(4505));
    layer3_outputs(3549) <= layer2_outputs(4954);
    layer3_outputs(3550) <= '1';
    layer3_outputs(3551) <= '1';
    layer3_outputs(3552) <= (layer2_outputs(1628)) and (layer2_outputs(864));
    layer3_outputs(3553) <= layer2_outputs(3650);
    layer3_outputs(3554) <= layer2_outputs(4415);
    layer3_outputs(3555) <= (layer2_outputs(1322)) or (layer2_outputs(2700));
    layer3_outputs(3556) <= not(layer2_outputs(622)) or (layer2_outputs(1899));
    layer3_outputs(3557) <= not(layer2_outputs(536));
    layer3_outputs(3558) <= (layer2_outputs(4652)) or (layer2_outputs(2261));
    layer3_outputs(3559) <= '1';
    layer3_outputs(3560) <= not(layer2_outputs(1754));
    layer3_outputs(3561) <= not(layer2_outputs(501)) or (layer2_outputs(1243));
    layer3_outputs(3562) <= not(layer2_outputs(3130));
    layer3_outputs(3563) <= not((layer2_outputs(2665)) or (layer2_outputs(3871)));
    layer3_outputs(3564) <= not((layer2_outputs(4093)) or (layer2_outputs(1817)));
    layer3_outputs(3565) <= layer2_outputs(2516);
    layer3_outputs(3566) <= layer2_outputs(1007);
    layer3_outputs(3567) <= '1';
    layer3_outputs(3568) <= not(layer2_outputs(834));
    layer3_outputs(3569) <= not((layer2_outputs(284)) or (layer2_outputs(4531)));
    layer3_outputs(3570) <= (layer2_outputs(3793)) or (layer2_outputs(4443));
    layer3_outputs(3571) <= not(layer2_outputs(2462));
    layer3_outputs(3572) <= not(layer2_outputs(249));
    layer3_outputs(3573) <= (layer2_outputs(3959)) and (layer2_outputs(1620));
    layer3_outputs(3574) <= not(layer2_outputs(1160));
    layer3_outputs(3575) <= not(layer2_outputs(2320));
    layer3_outputs(3576) <= not(layer2_outputs(921));
    layer3_outputs(3577) <= layer2_outputs(1171);
    layer3_outputs(3578) <= (layer2_outputs(2009)) xor (layer2_outputs(3039));
    layer3_outputs(3579) <= not(layer2_outputs(61));
    layer3_outputs(3580) <= layer2_outputs(4675);
    layer3_outputs(3581) <= not((layer2_outputs(4330)) or (layer2_outputs(2568)));
    layer3_outputs(3582) <= (layer2_outputs(406)) and (layer2_outputs(4984));
    layer3_outputs(3583) <= not(layer2_outputs(132)) or (layer2_outputs(1255));
    layer3_outputs(3584) <= (layer2_outputs(122)) and not (layer2_outputs(3426));
    layer3_outputs(3585) <= '1';
    layer3_outputs(3586) <= not(layer2_outputs(4892));
    layer3_outputs(3587) <= not(layer2_outputs(3905)) or (layer2_outputs(3118));
    layer3_outputs(3588) <= (layer2_outputs(3515)) and (layer2_outputs(3634));
    layer3_outputs(3589) <= layer2_outputs(488);
    layer3_outputs(3590) <= layer2_outputs(880);
    layer3_outputs(3591) <= '1';
    layer3_outputs(3592) <= (layer2_outputs(574)) and not (layer2_outputs(2986));
    layer3_outputs(3593) <= not((layer2_outputs(1661)) and (layer2_outputs(2758)));
    layer3_outputs(3594) <= layer2_outputs(1800);
    layer3_outputs(3595) <= not((layer2_outputs(4700)) or (layer2_outputs(5053)));
    layer3_outputs(3596) <= not((layer2_outputs(2429)) or (layer2_outputs(325)));
    layer3_outputs(3597) <= layer2_outputs(3329);
    layer3_outputs(3598) <= not(layer2_outputs(5093));
    layer3_outputs(3599) <= layer2_outputs(1765);
    layer3_outputs(3600) <= (layer2_outputs(2977)) and not (layer2_outputs(3183));
    layer3_outputs(3601) <= not(layer2_outputs(743)) or (layer2_outputs(121));
    layer3_outputs(3602) <= not(layer2_outputs(4010));
    layer3_outputs(3603) <= '0';
    layer3_outputs(3604) <= not(layer2_outputs(1633));
    layer3_outputs(3605) <= layer2_outputs(795);
    layer3_outputs(3606) <= not(layer2_outputs(1869));
    layer3_outputs(3607) <= not((layer2_outputs(4300)) or (layer2_outputs(3703)));
    layer3_outputs(3608) <= '0';
    layer3_outputs(3609) <= (layer2_outputs(3112)) and not (layer2_outputs(1950));
    layer3_outputs(3610) <= (layer2_outputs(2912)) and (layer2_outputs(3755));
    layer3_outputs(3611) <= '0';
    layer3_outputs(3612) <= (layer2_outputs(2116)) and not (layer2_outputs(1655));
    layer3_outputs(3613) <= '0';
    layer3_outputs(3614) <= not(layer2_outputs(285)) or (layer2_outputs(3522));
    layer3_outputs(3615) <= layer2_outputs(570);
    layer3_outputs(3616) <= '1';
    layer3_outputs(3617) <= not((layer2_outputs(3742)) xor (layer2_outputs(539)));
    layer3_outputs(3618) <= layer2_outputs(3078);
    layer3_outputs(3619) <= '1';
    layer3_outputs(3620) <= (layer2_outputs(466)) xor (layer2_outputs(4011));
    layer3_outputs(3621) <= layer2_outputs(2672);
    layer3_outputs(3622) <= not((layer2_outputs(2612)) and (layer2_outputs(4648)));
    layer3_outputs(3623) <= not(layer2_outputs(4361));
    layer3_outputs(3624) <= not(layer2_outputs(1522));
    layer3_outputs(3625) <= not(layer2_outputs(1783));
    layer3_outputs(3626) <= layer2_outputs(4110);
    layer3_outputs(3627) <= not(layer2_outputs(1937)) or (layer2_outputs(1799));
    layer3_outputs(3628) <= not(layer2_outputs(2321));
    layer3_outputs(3629) <= not(layer2_outputs(3036));
    layer3_outputs(3630) <= not(layer2_outputs(5037));
    layer3_outputs(3631) <= layer2_outputs(2072);
    layer3_outputs(3632) <= layer2_outputs(4372);
    layer3_outputs(3633) <= not(layer2_outputs(1531)) or (layer2_outputs(1867));
    layer3_outputs(3634) <= not(layer2_outputs(3163));
    layer3_outputs(3635) <= '0';
    layer3_outputs(3636) <= '0';
    layer3_outputs(3637) <= (layer2_outputs(2008)) or (layer2_outputs(4212));
    layer3_outputs(3638) <= layer2_outputs(4198);
    layer3_outputs(3639) <= not(layer2_outputs(638));
    layer3_outputs(3640) <= not(layer2_outputs(3708));
    layer3_outputs(3641) <= (layer2_outputs(2984)) or (layer2_outputs(2364));
    layer3_outputs(3642) <= '0';
    layer3_outputs(3643) <= layer2_outputs(3038);
    layer3_outputs(3644) <= layer2_outputs(1361);
    layer3_outputs(3645) <= not(layer2_outputs(3185)) or (layer2_outputs(1647));
    layer3_outputs(3646) <= not((layer2_outputs(4044)) and (layer2_outputs(4543)));
    layer3_outputs(3647) <= not(layer2_outputs(4318)) or (layer2_outputs(635));
    layer3_outputs(3648) <= (layer2_outputs(1947)) and not (layer2_outputs(2058));
    layer3_outputs(3649) <= layer2_outputs(4392);
    layer3_outputs(3650) <= '1';
    layer3_outputs(3651) <= not(layer2_outputs(4090)) or (layer2_outputs(4995));
    layer3_outputs(3652) <= not(layer2_outputs(545)) or (layer2_outputs(3211));
    layer3_outputs(3653) <= not((layer2_outputs(261)) and (layer2_outputs(1129)));
    layer3_outputs(3654) <= not((layer2_outputs(2882)) and (layer2_outputs(2526)));
    layer3_outputs(3655) <= not(layer2_outputs(1045));
    layer3_outputs(3656) <= layer2_outputs(765);
    layer3_outputs(3657) <= not(layer2_outputs(1602)) or (layer2_outputs(819));
    layer3_outputs(3658) <= layer2_outputs(4409);
    layer3_outputs(3659) <= (layer2_outputs(4104)) and (layer2_outputs(4257));
    layer3_outputs(3660) <= (layer2_outputs(4770)) and not (layer2_outputs(1384));
    layer3_outputs(3661) <= layer2_outputs(2942);
    layer3_outputs(3662) <= not(layer2_outputs(1079));
    layer3_outputs(3663) <= not((layer2_outputs(4359)) and (layer2_outputs(5073)));
    layer3_outputs(3664) <= not(layer2_outputs(3293));
    layer3_outputs(3665) <= not(layer2_outputs(5));
    layer3_outputs(3666) <= not(layer2_outputs(3006));
    layer3_outputs(3667) <= layer2_outputs(4295);
    layer3_outputs(3668) <= layer2_outputs(3652);
    layer3_outputs(3669) <= not(layer2_outputs(2766));
    layer3_outputs(3670) <= layer2_outputs(4655);
    layer3_outputs(3671) <= layer2_outputs(4101);
    layer3_outputs(3672) <= (layer2_outputs(422)) and not (layer2_outputs(2215));
    layer3_outputs(3673) <= not(layer2_outputs(2385));
    layer3_outputs(3674) <= not(layer2_outputs(1487)) or (layer2_outputs(1900));
    layer3_outputs(3675) <= layer2_outputs(2059);
    layer3_outputs(3676) <= not(layer2_outputs(2742));
    layer3_outputs(3677) <= '0';
    layer3_outputs(3678) <= '0';
    layer3_outputs(3679) <= (layer2_outputs(428)) or (layer2_outputs(4285));
    layer3_outputs(3680) <= not((layer2_outputs(45)) and (layer2_outputs(1695)));
    layer3_outputs(3681) <= (layer2_outputs(2178)) and (layer2_outputs(4028));
    layer3_outputs(3682) <= layer2_outputs(3649);
    layer3_outputs(3683) <= not(layer2_outputs(1611));
    layer3_outputs(3684) <= '0';
    layer3_outputs(3685) <= not((layer2_outputs(5118)) and (layer2_outputs(3166)));
    layer3_outputs(3686) <= not((layer2_outputs(828)) and (layer2_outputs(1446)));
    layer3_outputs(3687) <= not(layer2_outputs(121));
    layer3_outputs(3688) <= (layer2_outputs(3541)) or (layer2_outputs(5018));
    layer3_outputs(3689) <= (layer2_outputs(3724)) and (layer2_outputs(4403));
    layer3_outputs(3690) <= (layer2_outputs(4379)) and (layer2_outputs(4696));
    layer3_outputs(3691) <= not(layer2_outputs(4499));
    layer3_outputs(3692) <= not((layer2_outputs(716)) and (layer2_outputs(4315)));
    layer3_outputs(3693) <= (layer2_outputs(2637)) or (layer2_outputs(341));
    layer3_outputs(3694) <= (layer2_outputs(3094)) and not (layer2_outputs(3399));
    layer3_outputs(3695) <= '0';
    layer3_outputs(3696) <= layer2_outputs(1389);
    layer3_outputs(3697) <= not(layer2_outputs(2561));
    layer3_outputs(3698) <= (layer2_outputs(4967)) and (layer2_outputs(4829));
    layer3_outputs(3699) <= (layer2_outputs(728)) and (layer2_outputs(778));
    layer3_outputs(3700) <= layer2_outputs(3373);
    layer3_outputs(3701) <= not(layer2_outputs(3321));
    layer3_outputs(3702) <= (layer2_outputs(3429)) and not (layer2_outputs(3064));
    layer3_outputs(3703) <= (layer2_outputs(4791)) and (layer2_outputs(479));
    layer3_outputs(3704) <= (layer2_outputs(1935)) or (layer2_outputs(3002));
    layer3_outputs(3705) <= (layer2_outputs(1596)) and not (layer2_outputs(1855));
    layer3_outputs(3706) <= layer2_outputs(48);
    layer3_outputs(3707) <= (layer2_outputs(771)) and (layer2_outputs(4296));
    layer3_outputs(3708) <= layer2_outputs(262);
    layer3_outputs(3709) <= '1';
    layer3_outputs(3710) <= not(layer2_outputs(2090)) or (layer2_outputs(291));
    layer3_outputs(3711) <= '1';
    layer3_outputs(3712) <= not(layer2_outputs(2487)) or (layer2_outputs(1014));
    layer3_outputs(3713) <= (layer2_outputs(38)) and not (layer2_outputs(2516));
    layer3_outputs(3714) <= '1';
    layer3_outputs(3715) <= (layer2_outputs(2772)) or (layer2_outputs(5007));
    layer3_outputs(3716) <= not((layer2_outputs(1062)) and (layer2_outputs(4392)));
    layer3_outputs(3717) <= (layer2_outputs(85)) or (layer2_outputs(4422));
    layer3_outputs(3718) <= not(layer2_outputs(2400));
    layer3_outputs(3719) <= not(layer2_outputs(4122)) or (layer2_outputs(2375));
    layer3_outputs(3720) <= '1';
    layer3_outputs(3721) <= (layer2_outputs(2224)) and not (layer2_outputs(3753));
    layer3_outputs(3722) <= not(layer2_outputs(1268));
    layer3_outputs(3723) <= not(layer2_outputs(3798));
    layer3_outputs(3724) <= '1';
    layer3_outputs(3725) <= (layer2_outputs(4874)) and not (layer2_outputs(4625));
    layer3_outputs(3726) <= not(layer2_outputs(4893)) or (layer2_outputs(1802));
    layer3_outputs(3727) <= not(layer2_outputs(1690)) or (layer2_outputs(270));
    layer3_outputs(3728) <= layer2_outputs(3588);
    layer3_outputs(3729) <= not(layer2_outputs(4239)) or (layer2_outputs(4520));
    layer3_outputs(3730) <= not((layer2_outputs(2755)) xor (layer2_outputs(457)));
    layer3_outputs(3731) <= layer2_outputs(4255);
    layer3_outputs(3732) <= not(layer2_outputs(599)) or (layer2_outputs(2839));
    layer3_outputs(3733) <= (layer2_outputs(1121)) and not (layer2_outputs(1482));
    layer3_outputs(3734) <= not(layer2_outputs(2334));
    layer3_outputs(3735) <= layer2_outputs(3927);
    layer3_outputs(3736) <= (layer2_outputs(4087)) and not (layer2_outputs(3781));
    layer3_outputs(3737) <= '0';
    layer3_outputs(3738) <= '1';
    layer3_outputs(3739) <= layer2_outputs(729);
    layer3_outputs(3740) <= not(layer2_outputs(1981)) or (layer2_outputs(2908));
    layer3_outputs(3741) <= (layer2_outputs(191)) or (layer2_outputs(2834));
    layer3_outputs(3742) <= not((layer2_outputs(784)) or (layer2_outputs(1232)));
    layer3_outputs(3743) <= not((layer2_outputs(2720)) xor (layer2_outputs(4019)));
    layer3_outputs(3744) <= not(layer2_outputs(1675));
    layer3_outputs(3745) <= not(layer2_outputs(768));
    layer3_outputs(3746) <= layer2_outputs(4160);
    layer3_outputs(3747) <= not(layer2_outputs(1234)) or (layer2_outputs(2367));
    layer3_outputs(3748) <= '1';
    layer3_outputs(3749) <= '1';
    layer3_outputs(3750) <= layer2_outputs(4349);
    layer3_outputs(3751) <= layer2_outputs(576);
    layer3_outputs(3752) <= '1';
    layer3_outputs(3753) <= not(layer2_outputs(4454));
    layer3_outputs(3754) <= not(layer2_outputs(1134)) or (layer2_outputs(3889));
    layer3_outputs(3755) <= not(layer2_outputs(874));
    layer3_outputs(3756) <= layer2_outputs(438);
    layer3_outputs(3757) <= not(layer2_outputs(2161)) or (layer2_outputs(1384));
    layer3_outputs(3758) <= not(layer2_outputs(1205));
    layer3_outputs(3759) <= layer2_outputs(420);
    layer3_outputs(3760) <= (layer2_outputs(4816)) or (layer2_outputs(3983));
    layer3_outputs(3761) <= (layer2_outputs(3244)) xor (layer2_outputs(2166));
    layer3_outputs(3762) <= (layer2_outputs(2323)) or (layer2_outputs(4568));
    layer3_outputs(3763) <= (layer2_outputs(3870)) and not (layer2_outputs(763));
    layer3_outputs(3764) <= layer2_outputs(2181);
    layer3_outputs(3765) <= (layer2_outputs(3256)) xor (layer2_outputs(1817));
    layer3_outputs(3766) <= not(layer2_outputs(3819));
    layer3_outputs(3767) <= (layer2_outputs(1269)) and not (layer2_outputs(3038));
    layer3_outputs(3768) <= not(layer2_outputs(1348)) or (layer2_outputs(4838));
    layer3_outputs(3769) <= not(layer2_outputs(1555));
    layer3_outputs(3770) <= (layer2_outputs(3244)) and (layer2_outputs(938));
    layer3_outputs(3771) <= '0';
    layer3_outputs(3772) <= not((layer2_outputs(948)) xor (layer2_outputs(3611)));
    layer3_outputs(3773) <= (layer2_outputs(4283)) and not (layer2_outputs(1066));
    layer3_outputs(3774) <= (layer2_outputs(1550)) and not (layer2_outputs(4159));
    layer3_outputs(3775) <= not(layer2_outputs(2210)) or (layer2_outputs(4825));
    layer3_outputs(3776) <= not((layer2_outputs(2726)) and (layer2_outputs(1499)));
    layer3_outputs(3777) <= not((layer2_outputs(3361)) xor (layer2_outputs(2626)));
    layer3_outputs(3778) <= '0';
    layer3_outputs(3779) <= layer2_outputs(4681);
    layer3_outputs(3780) <= not((layer2_outputs(1833)) and (layer2_outputs(2655)));
    layer3_outputs(3781) <= not(layer2_outputs(727)) or (layer2_outputs(3243));
    layer3_outputs(3782) <= layer2_outputs(67);
    layer3_outputs(3783) <= (layer2_outputs(1035)) and not (layer2_outputs(1733));
    layer3_outputs(3784) <= (layer2_outputs(3308)) and not (layer2_outputs(1804));
    layer3_outputs(3785) <= not(layer2_outputs(4628)) or (layer2_outputs(256));
    layer3_outputs(3786) <= (layer2_outputs(4049)) xor (layer2_outputs(3555));
    layer3_outputs(3787) <= not((layer2_outputs(68)) and (layer2_outputs(668)));
    layer3_outputs(3788) <= not((layer2_outputs(2590)) or (layer2_outputs(968)));
    layer3_outputs(3789) <= layer2_outputs(1514);
    layer3_outputs(3790) <= (layer2_outputs(4638)) and not (layer2_outputs(861));
    layer3_outputs(3791) <= layer2_outputs(1405);
    layer3_outputs(3792) <= not(layer2_outputs(160));
    layer3_outputs(3793) <= (layer2_outputs(4802)) xor (layer2_outputs(2898));
    layer3_outputs(3794) <= not(layer2_outputs(4510));
    layer3_outputs(3795) <= '1';
    layer3_outputs(3796) <= '1';
    layer3_outputs(3797) <= not(layer2_outputs(1049));
    layer3_outputs(3798) <= '1';
    layer3_outputs(3799) <= not(layer2_outputs(92)) or (layer2_outputs(1657));
    layer3_outputs(3800) <= not((layer2_outputs(4016)) xor (layer2_outputs(4951)));
    layer3_outputs(3801) <= not(layer2_outputs(3901)) or (layer2_outputs(4309));
    layer3_outputs(3802) <= not((layer2_outputs(3291)) xor (layer2_outputs(2843)));
    layer3_outputs(3803) <= not((layer2_outputs(3959)) and (layer2_outputs(4547)));
    layer3_outputs(3804) <= not((layer2_outputs(3272)) or (layer2_outputs(1595)));
    layer3_outputs(3805) <= (layer2_outputs(2107)) and not (layer2_outputs(3789));
    layer3_outputs(3806) <= (layer2_outputs(4920)) and not (layer2_outputs(1345));
    layer3_outputs(3807) <= not(layer2_outputs(3378));
    layer3_outputs(3808) <= '1';
    layer3_outputs(3809) <= not((layer2_outputs(4461)) or (layer2_outputs(1514)));
    layer3_outputs(3810) <= not((layer2_outputs(2645)) or (layer2_outputs(3151)));
    layer3_outputs(3811) <= layer2_outputs(3082);
    layer3_outputs(3812) <= layer2_outputs(459);
    layer3_outputs(3813) <= (layer2_outputs(2631)) and not (layer2_outputs(1879));
    layer3_outputs(3814) <= not((layer2_outputs(2408)) or (layer2_outputs(1959)));
    layer3_outputs(3815) <= layer2_outputs(3432);
    layer3_outputs(3816) <= not(layer2_outputs(380)) or (layer2_outputs(3436));
    layer3_outputs(3817) <= layer2_outputs(1958);
    layer3_outputs(3818) <= not((layer2_outputs(2414)) and (layer2_outputs(4884)));
    layer3_outputs(3819) <= layer2_outputs(2692);
    layer3_outputs(3820) <= (layer2_outputs(3615)) and not (layer2_outputs(2459));
    layer3_outputs(3821) <= not(layer2_outputs(2412));
    layer3_outputs(3822) <= not(layer2_outputs(4023));
    layer3_outputs(3823) <= not(layer2_outputs(227));
    layer3_outputs(3824) <= (layer2_outputs(4214)) or (layer2_outputs(1830));
    layer3_outputs(3825) <= not((layer2_outputs(3216)) or (layer2_outputs(4557)));
    layer3_outputs(3826) <= layer2_outputs(1669);
    layer3_outputs(3827) <= (layer2_outputs(1228)) and not (layer2_outputs(349));
    layer3_outputs(3828) <= (layer2_outputs(1451)) and not (layer2_outputs(1847));
    layer3_outputs(3829) <= not((layer2_outputs(2735)) and (layer2_outputs(5067)));
    layer3_outputs(3830) <= (layer2_outputs(962)) and not (layer2_outputs(1902));
    layer3_outputs(3831) <= (layer2_outputs(4445)) or (layer2_outputs(3399));
    layer3_outputs(3832) <= not(layer2_outputs(2301)) or (layer2_outputs(2234));
    layer3_outputs(3833) <= not(layer2_outputs(4815));
    layer3_outputs(3834) <= layer2_outputs(4965);
    layer3_outputs(3835) <= (layer2_outputs(2474)) or (layer2_outputs(2398));
    layer3_outputs(3836) <= not(layer2_outputs(4078));
    layer3_outputs(3837) <= (layer2_outputs(711)) and not (layer2_outputs(3762));
    layer3_outputs(3838) <= not(layer2_outputs(499));
    layer3_outputs(3839) <= layer2_outputs(4043);
    layer3_outputs(3840) <= layer2_outputs(2761);
    layer3_outputs(3841) <= not(layer2_outputs(1461)) or (layer2_outputs(1154));
    layer3_outputs(3842) <= not(layer2_outputs(4725)) or (layer2_outputs(1520));
    layer3_outputs(3843) <= not(layer2_outputs(3405));
    layer3_outputs(3844) <= (layer2_outputs(841)) or (layer2_outputs(1423));
    layer3_outputs(3845) <= '1';
    layer3_outputs(3846) <= not((layer2_outputs(2820)) or (layer2_outputs(3178)));
    layer3_outputs(3847) <= not(layer2_outputs(2902));
    layer3_outputs(3848) <= not(layer2_outputs(2592)) or (layer2_outputs(3449));
    layer3_outputs(3849) <= layer2_outputs(3639);
    layer3_outputs(3850) <= layer2_outputs(420);
    layer3_outputs(3851) <= not(layer2_outputs(2937));
    layer3_outputs(3852) <= not(layer2_outputs(1985)) or (layer2_outputs(1334));
    layer3_outputs(3853) <= '0';
    layer3_outputs(3854) <= not(layer2_outputs(1726));
    layer3_outputs(3855) <= (layer2_outputs(2899)) and not (layer2_outputs(4939));
    layer3_outputs(3856) <= not(layer2_outputs(373));
    layer3_outputs(3857) <= (layer2_outputs(2182)) or (layer2_outputs(3096));
    layer3_outputs(3858) <= not(layer2_outputs(1353));
    layer3_outputs(3859) <= '1';
    layer3_outputs(3860) <= (layer2_outputs(1679)) and (layer2_outputs(1167));
    layer3_outputs(3861) <= not(layer2_outputs(4551));
    layer3_outputs(3862) <= not((layer2_outputs(3575)) or (layer2_outputs(3585)));
    layer3_outputs(3863) <= not((layer2_outputs(2111)) and (layer2_outputs(22)));
    layer3_outputs(3864) <= not(layer2_outputs(1112)) or (layer2_outputs(2222));
    layer3_outputs(3865) <= layer2_outputs(4534);
    layer3_outputs(3866) <= not(layer2_outputs(678));
    layer3_outputs(3867) <= not((layer2_outputs(644)) and (layer2_outputs(2872)));
    layer3_outputs(3868) <= '0';
    layer3_outputs(3869) <= not(layer2_outputs(1331));
    layer3_outputs(3870) <= not(layer2_outputs(2251));
    layer3_outputs(3871) <= not(layer2_outputs(538));
    layer3_outputs(3872) <= layer2_outputs(2894);
    layer3_outputs(3873) <= (layer2_outputs(949)) and not (layer2_outputs(2594));
    layer3_outputs(3874) <= not(layer2_outputs(2193)) or (layer2_outputs(663));
    layer3_outputs(3875) <= not((layer2_outputs(3915)) and (layer2_outputs(514)));
    layer3_outputs(3876) <= not((layer2_outputs(4612)) and (layer2_outputs(3338)));
    layer3_outputs(3877) <= not((layer2_outputs(4743)) xor (layer2_outputs(13)));
    layer3_outputs(3878) <= not(layer2_outputs(1542));
    layer3_outputs(3879) <= (layer2_outputs(2852)) and not (layer2_outputs(1026));
    layer3_outputs(3880) <= layer2_outputs(3305);
    layer3_outputs(3881) <= not((layer2_outputs(1931)) and (layer2_outputs(1146)));
    layer3_outputs(3882) <= not(layer2_outputs(2757));
    layer3_outputs(3883) <= not(layer2_outputs(4289));
    layer3_outputs(3884) <= layer2_outputs(1262);
    layer3_outputs(3885) <= not(layer2_outputs(372)) or (layer2_outputs(4821));
    layer3_outputs(3886) <= (layer2_outputs(1177)) and not (layer2_outputs(1050));
    layer3_outputs(3887) <= not(layer2_outputs(5016));
    layer3_outputs(3888) <= layer2_outputs(3699);
    layer3_outputs(3889) <= not(layer2_outputs(2076));
    layer3_outputs(3890) <= not(layer2_outputs(34));
    layer3_outputs(3891) <= layer2_outputs(2718);
    layer3_outputs(3892) <= (layer2_outputs(4286)) and not (layer2_outputs(3783));
    layer3_outputs(3893) <= layer2_outputs(3974);
    layer3_outputs(3894) <= layer2_outputs(4100);
    layer3_outputs(3895) <= not(layer2_outputs(1632));
    layer3_outputs(3896) <= '1';
    layer3_outputs(3897) <= layer2_outputs(3115);
    layer3_outputs(3898) <= (layer2_outputs(757)) and (layer2_outputs(4661));
    layer3_outputs(3899) <= not(layer2_outputs(2353));
    layer3_outputs(3900) <= layer2_outputs(2825);
    layer3_outputs(3901) <= layer2_outputs(4994);
    layer3_outputs(3902) <= not((layer2_outputs(4373)) and (layer2_outputs(4471)));
    layer3_outputs(3903) <= layer2_outputs(709);
    layer3_outputs(3904) <= '0';
    layer3_outputs(3905) <= layer2_outputs(1717);
    layer3_outputs(3906) <= not((layer2_outputs(3080)) and (layer2_outputs(562)));
    layer3_outputs(3907) <= (layer2_outputs(681)) and not (layer2_outputs(4346));
    layer3_outputs(3908) <= (layer2_outputs(1238)) and not (layer2_outputs(23));
    layer3_outputs(3909) <= (layer2_outputs(253)) and not (layer2_outputs(11));
    layer3_outputs(3910) <= layer2_outputs(1974);
    layer3_outputs(3911) <= '0';
    layer3_outputs(3912) <= (layer2_outputs(588)) and not (layer2_outputs(3353));
    layer3_outputs(3913) <= (layer2_outputs(3649)) or (layer2_outputs(3821));
    layer3_outputs(3914) <= (layer2_outputs(3658)) and not (layer2_outputs(1260));
    layer3_outputs(3915) <= not(layer2_outputs(4316)) or (layer2_outputs(4690));
    layer3_outputs(3916) <= layer2_outputs(446);
    layer3_outputs(3917) <= (layer2_outputs(1182)) and (layer2_outputs(3769));
    layer3_outputs(3918) <= layer2_outputs(4574);
    layer3_outputs(3919) <= (layer2_outputs(2923)) and not (layer2_outputs(2398));
    layer3_outputs(3920) <= (layer2_outputs(4522)) and (layer2_outputs(805));
    layer3_outputs(3921) <= not(layer2_outputs(2828));
    layer3_outputs(3922) <= (layer2_outputs(1388)) and not (layer2_outputs(2837));
    layer3_outputs(3923) <= layer2_outputs(3099);
    layer3_outputs(3924) <= not(layer2_outputs(1640)) or (layer2_outputs(1114));
    layer3_outputs(3925) <= not(layer2_outputs(624));
    layer3_outputs(3926) <= (layer2_outputs(2050)) or (layer2_outputs(1743));
    layer3_outputs(3927) <= not(layer2_outputs(1042)) or (layer2_outputs(4601));
    layer3_outputs(3928) <= (layer2_outputs(4699)) and not (layer2_outputs(4873));
    layer3_outputs(3929) <= '0';
    layer3_outputs(3930) <= not(layer2_outputs(93));
    layer3_outputs(3931) <= (layer2_outputs(4799)) and not (layer2_outputs(1932));
    layer3_outputs(3932) <= not(layer2_outputs(1337)) or (layer2_outputs(148));
    layer3_outputs(3933) <= not(layer2_outputs(3065));
    layer3_outputs(3934) <= layer2_outputs(2274);
    layer3_outputs(3935) <= not(layer2_outputs(620));
    layer3_outputs(3936) <= not(layer2_outputs(65)) or (layer2_outputs(553));
    layer3_outputs(3937) <= '1';
    layer3_outputs(3938) <= (layer2_outputs(3417)) and not (layer2_outputs(2388));
    layer3_outputs(3939) <= not((layer2_outputs(2195)) xor (layer2_outputs(1256)));
    layer3_outputs(3940) <= not(layer2_outputs(3180));
    layer3_outputs(3941) <= '0';
    layer3_outputs(3942) <= not(layer2_outputs(1748)) or (layer2_outputs(3159));
    layer3_outputs(3943) <= not((layer2_outputs(1323)) or (layer2_outputs(4682)));
    layer3_outputs(3944) <= not(layer2_outputs(2133));
    layer3_outputs(3945) <= not(layer2_outputs(5000));
    layer3_outputs(3946) <= not(layer2_outputs(1972));
    layer3_outputs(3947) <= layer2_outputs(1211);
    layer3_outputs(3948) <= not(layer2_outputs(3386));
    layer3_outputs(3949) <= not(layer2_outputs(606)) or (layer2_outputs(2100));
    layer3_outputs(3950) <= (layer2_outputs(1099)) or (layer2_outputs(3010));
    layer3_outputs(3951) <= '0';
    layer3_outputs(3952) <= layer2_outputs(1819);
    layer3_outputs(3953) <= layer2_outputs(580);
    layer3_outputs(3954) <= layer2_outputs(950);
    layer3_outputs(3955) <= (layer2_outputs(2991)) or (layer2_outputs(1302));
    layer3_outputs(3956) <= (layer2_outputs(993)) and not (layer2_outputs(2713));
    layer3_outputs(3957) <= not((layer2_outputs(392)) and (layer2_outputs(2284)));
    layer3_outputs(3958) <= not(layer2_outputs(3477));
    layer3_outputs(3959) <= '1';
    layer3_outputs(3960) <= not(layer2_outputs(3360));
    layer3_outputs(3961) <= not(layer2_outputs(554));
    layer3_outputs(3962) <= layer2_outputs(4497);
    layer3_outputs(3963) <= not(layer2_outputs(564));
    layer3_outputs(3964) <= not(layer2_outputs(391));
    layer3_outputs(3965) <= '1';
    layer3_outputs(3966) <= not((layer2_outputs(2978)) and (layer2_outputs(3321)));
    layer3_outputs(3967) <= not(layer2_outputs(4870));
    layer3_outputs(3968) <= (layer2_outputs(4652)) and not (layer2_outputs(294));
    layer3_outputs(3969) <= not((layer2_outputs(2764)) and (layer2_outputs(2471)));
    layer3_outputs(3970) <= not(layer2_outputs(3208)) or (layer2_outputs(1139));
    layer3_outputs(3971) <= (layer2_outputs(2101)) and not (layer2_outputs(4000));
    layer3_outputs(3972) <= '1';
    layer3_outputs(3973) <= not((layer2_outputs(3987)) or (layer2_outputs(4274)));
    layer3_outputs(3974) <= (layer2_outputs(2046)) and (layer2_outputs(4584));
    layer3_outputs(3975) <= (layer2_outputs(5052)) and (layer2_outputs(3438));
    layer3_outputs(3976) <= not(layer2_outputs(1732));
    layer3_outputs(3977) <= not((layer2_outputs(3716)) or (layer2_outputs(183)));
    layer3_outputs(3978) <= layer2_outputs(873);
    layer3_outputs(3979) <= '1';
    layer3_outputs(3980) <= not((layer2_outputs(1888)) and (layer2_outputs(783)));
    layer3_outputs(3981) <= (layer2_outputs(4549)) and not (layer2_outputs(4404));
    layer3_outputs(3982) <= not((layer2_outputs(2214)) and (layer2_outputs(2644)));
    layer3_outputs(3983) <= not(layer2_outputs(1774));
    layer3_outputs(3984) <= (layer2_outputs(1347)) and not (layer2_outputs(2358));
    layer3_outputs(3985) <= layer2_outputs(1850);
    layer3_outputs(3986) <= not(layer2_outputs(694)) or (layer2_outputs(3898));
    layer3_outputs(3987) <= (layer2_outputs(1067)) and not (layer2_outputs(3441));
    layer3_outputs(3988) <= (layer2_outputs(4643)) and (layer2_outputs(3263));
    layer3_outputs(3989) <= '0';
    layer3_outputs(3990) <= not((layer2_outputs(4485)) xor (layer2_outputs(4481)));
    layer3_outputs(3991) <= layer2_outputs(1732);
    layer3_outputs(3992) <= not((layer2_outputs(4649)) or (layer2_outputs(260)));
    layer3_outputs(3993) <= not(layer2_outputs(333)) or (layer2_outputs(1787));
    layer3_outputs(3994) <= layer2_outputs(3954);
    layer3_outputs(3995) <= not(layer2_outputs(634)) or (layer2_outputs(2909));
    layer3_outputs(3996) <= not((layer2_outputs(1836)) or (layer2_outputs(1286)));
    layer3_outputs(3997) <= not(layer2_outputs(4897));
    layer3_outputs(3998) <= '0';
    layer3_outputs(3999) <= not(layer2_outputs(3358)) or (layer2_outputs(980));
    layer3_outputs(4000) <= (layer2_outputs(955)) and not (layer2_outputs(1329));
    layer3_outputs(4001) <= not(layer2_outputs(1601));
    layer3_outputs(4002) <= not(layer2_outputs(2042));
    layer3_outputs(4003) <= not(layer2_outputs(4321)) or (layer2_outputs(2658));
    layer3_outputs(4004) <= not((layer2_outputs(25)) or (layer2_outputs(3442)));
    layer3_outputs(4005) <= (layer2_outputs(4888)) and not (layer2_outputs(3237));
    layer3_outputs(4006) <= not(layer2_outputs(899));
    layer3_outputs(4007) <= (layer2_outputs(1781)) or (layer2_outputs(3164));
    layer3_outputs(4008) <= '0';
    layer3_outputs(4009) <= not(layer2_outputs(2562)) or (layer2_outputs(450));
    layer3_outputs(4010) <= layer2_outputs(4570);
    layer3_outputs(4011) <= (layer2_outputs(3932)) and (layer2_outputs(1639));
    layer3_outputs(4012) <= '1';
    layer3_outputs(4013) <= not(layer2_outputs(1084)) or (layer2_outputs(3734));
    layer3_outputs(4014) <= not(layer2_outputs(26)) or (layer2_outputs(1409));
    layer3_outputs(4015) <= (layer2_outputs(4762)) and not (layer2_outputs(1961));
    layer3_outputs(4016) <= (layer2_outputs(3804)) or (layer2_outputs(4112));
    layer3_outputs(4017) <= not((layer2_outputs(1892)) and (layer2_outputs(2370)));
    layer3_outputs(4018) <= not((layer2_outputs(12)) or (layer2_outputs(304)));
    layer3_outputs(4019) <= (layer2_outputs(2578)) and not (layer2_outputs(2497));
    layer3_outputs(4020) <= not((layer2_outputs(313)) or (layer2_outputs(4066)));
    layer3_outputs(4021) <= '1';
    layer3_outputs(4022) <= (layer2_outputs(4427)) and not (layer2_outputs(3239));
    layer3_outputs(4023) <= (layer2_outputs(610)) and not (layer2_outputs(3228));
    layer3_outputs(4024) <= (layer2_outputs(2582)) or (layer2_outputs(163));
    layer3_outputs(4025) <= layer2_outputs(1599);
    layer3_outputs(4026) <= '0';
    layer3_outputs(4027) <= '0';
    layer3_outputs(4028) <= not((layer2_outputs(2058)) or (layer2_outputs(2070)));
    layer3_outputs(4029) <= '1';
    layer3_outputs(4030) <= not((layer2_outputs(3152)) and (layer2_outputs(2878)));
    layer3_outputs(4031) <= not(layer2_outputs(5099)) or (layer2_outputs(2149));
    layer3_outputs(4032) <= not(layer2_outputs(4403)) or (layer2_outputs(1547));
    layer3_outputs(4033) <= not((layer2_outputs(891)) and (layer2_outputs(328)));
    layer3_outputs(4034) <= layer2_outputs(4232);
    layer3_outputs(4035) <= (layer2_outputs(1812)) or (layer2_outputs(2380));
    layer3_outputs(4036) <= not((layer2_outputs(3324)) or (layer2_outputs(3240)));
    layer3_outputs(4037) <= layer2_outputs(4839);
    layer3_outputs(4038) <= (layer2_outputs(4306)) and not (layer2_outputs(2403));
    layer3_outputs(4039) <= not(layer2_outputs(3099));
    layer3_outputs(4040) <= not(layer2_outputs(3024)) or (layer2_outputs(470));
    layer3_outputs(4041) <= not(layer2_outputs(2803));
    layer3_outputs(4042) <= layer2_outputs(3937);
    layer3_outputs(4043) <= not((layer2_outputs(89)) or (layer2_outputs(30)));
    layer3_outputs(4044) <= (layer2_outputs(2927)) and (layer2_outputs(1181));
    layer3_outputs(4045) <= '0';
    layer3_outputs(4046) <= not(layer2_outputs(490)) or (layer2_outputs(4146));
    layer3_outputs(4047) <= layer2_outputs(1637);
    layer3_outputs(4048) <= '0';
    layer3_outputs(4049) <= (layer2_outputs(1999)) or (layer2_outputs(2469));
    layer3_outputs(4050) <= not(layer2_outputs(4295)) or (layer2_outputs(1219));
    layer3_outputs(4051) <= not((layer2_outputs(4820)) and (layer2_outputs(2753)));
    layer3_outputs(4052) <= not(layer2_outputs(1287)) or (layer2_outputs(2387));
    layer3_outputs(4053) <= not(layer2_outputs(4341)) or (layer2_outputs(2166));
    layer3_outputs(4054) <= '1';
    layer3_outputs(4055) <= '1';
    layer3_outputs(4056) <= layer2_outputs(760);
    layer3_outputs(4057) <= layer2_outputs(5104);
    layer3_outputs(4058) <= not((layer2_outputs(2104)) and (layer2_outputs(2397)));
    layer3_outputs(4059) <= layer2_outputs(217);
    layer3_outputs(4060) <= (layer2_outputs(1439)) and (layer2_outputs(1095));
    layer3_outputs(4061) <= '1';
    layer3_outputs(4062) <= (layer2_outputs(2078)) and (layer2_outputs(2339));
    layer3_outputs(4063) <= '0';
    layer3_outputs(4064) <= not(layer2_outputs(2287)) or (layer2_outputs(3924));
    layer3_outputs(4065) <= '0';
    layer3_outputs(4066) <= layer2_outputs(4734);
    layer3_outputs(4067) <= not(layer2_outputs(95));
    layer3_outputs(4068) <= layer2_outputs(3689);
    layer3_outputs(4069) <= not((layer2_outputs(4445)) or (layer2_outputs(3193)));
    layer3_outputs(4070) <= not(layer2_outputs(527));
    layer3_outputs(4071) <= not((layer2_outputs(618)) or (layer2_outputs(4985)));
    layer3_outputs(4072) <= not(layer2_outputs(3967)) or (layer2_outputs(4608));
    layer3_outputs(4073) <= '1';
    layer3_outputs(4074) <= not((layer2_outputs(2428)) or (layer2_outputs(2298)));
    layer3_outputs(4075) <= (layer2_outputs(4650)) or (layer2_outputs(2518));
    layer3_outputs(4076) <= layer2_outputs(4401);
    layer3_outputs(4077) <= layer2_outputs(1188);
    layer3_outputs(4078) <= (layer2_outputs(530)) and not (layer2_outputs(768));
    layer3_outputs(4079) <= '0';
    layer3_outputs(4080) <= not((layer2_outputs(1376)) or (layer2_outputs(2865)));
    layer3_outputs(4081) <= not(layer2_outputs(1605)) or (layer2_outputs(4724));
    layer3_outputs(4082) <= (layer2_outputs(3556)) or (layer2_outputs(524));
    layer3_outputs(4083) <= not(layer2_outputs(3331));
    layer3_outputs(4084) <= '0';
    layer3_outputs(4085) <= '1';
    layer3_outputs(4086) <= (layer2_outputs(721)) and (layer2_outputs(541));
    layer3_outputs(4087) <= (layer2_outputs(1521)) xor (layer2_outputs(1358));
    layer3_outputs(4088) <= layer2_outputs(2327);
    layer3_outputs(4089) <= '1';
    layer3_outputs(4090) <= not(layer2_outputs(3808));
    layer3_outputs(4091) <= layer2_outputs(2231);
    layer3_outputs(4092) <= '1';
    layer3_outputs(4093) <= '1';
    layer3_outputs(4094) <= not(layer2_outputs(4451));
    layer3_outputs(4095) <= (layer2_outputs(1562)) and not (layer2_outputs(1305));
    layer3_outputs(4096) <= layer2_outputs(2188);
    layer3_outputs(4097) <= layer2_outputs(533);
    layer3_outputs(4098) <= not((layer2_outputs(1634)) or (layer2_outputs(2765)));
    layer3_outputs(4099) <= (layer2_outputs(4402)) and (layer2_outputs(2975));
    layer3_outputs(4100) <= '1';
    layer3_outputs(4101) <= '1';
    layer3_outputs(4102) <= layer2_outputs(1768);
    layer3_outputs(4103) <= not(layer2_outputs(1357));
    layer3_outputs(4104) <= not(layer2_outputs(3983));
    layer3_outputs(4105) <= not(layer2_outputs(669));
    layer3_outputs(4106) <= layer2_outputs(2462);
    layer3_outputs(4107) <= not((layer2_outputs(3023)) and (layer2_outputs(2942)));
    layer3_outputs(4108) <= (layer2_outputs(243)) and not (layer2_outputs(573));
    layer3_outputs(4109) <= '1';
    layer3_outputs(4110) <= not(layer2_outputs(957)) or (layer2_outputs(507));
    layer3_outputs(4111) <= (layer2_outputs(2924)) and not (layer2_outputs(1009));
    layer3_outputs(4112) <= (layer2_outputs(2542)) and not (layer2_outputs(3397));
    layer3_outputs(4113) <= not(layer2_outputs(227)) or (layer2_outputs(628));
    layer3_outputs(4114) <= not(layer2_outputs(3665));
    layer3_outputs(4115) <= '0';
    layer3_outputs(4116) <= (layer2_outputs(518)) and not (layer2_outputs(5028));
    layer3_outputs(4117) <= layer2_outputs(5031);
    layer3_outputs(4118) <= (layer2_outputs(4244)) xor (layer2_outputs(1471));
    layer3_outputs(4119) <= not((layer2_outputs(3222)) and (layer2_outputs(4964)));
    layer3_outputs(4120) <= layer2_outputs(4671);
    layer3_outputs(4121) <= not(layer2_outputs(536));
    layer3_outputs(4122) <= (layer2_outputs(494)) xor (layer2_outputs(1266));
    layer3_outputs(4123) <= (layer2_outputs(556)) and not (layer2_outputs(4068));
    layer3_outputs(4124) <= layer2_outputs(1587);
    layer3_outputs(4125) <= not((layer2_outputs(2756)) xor (layer2_outputs(4256)));
    layer3_outputs(4126) <= layer2_outputs(2830);
    layer3_outputs(4127) <= '0';
    layer3_outputs(4128) <= not((layer2_outputs(172)) or (layer2_outputs(3138)));
    layer3_outputs(4129) <= not(layer2_outputs(257)) or (layer2_outputs(5012));
    layer3_outputs(4130) <= not((layer2_outputs(1301)) or (layer2_outputs(192)));
    layer3_outputs(4131) <= (layer2_outputs(3124)) and not (layer2_outputs(2193));
    layer3_outputs(4132) <= '1';
    layer3_outputs(4133) <= (layer2_outputs(3074)) and not (layer2_outputs(383));
    layer3_outputs(4134) <= (layer2_outputs(4229)) xor (layer2_outputs(1377));
    layer3_outputs(4135) <= not(layer2_outputs(722));
    layer3_outputs(4136) <= layer2_outputs(2478);
    layer3_outputs(4137) <= not(layer2_outputs(446));
    layer3_outputs(4138) <= (layer2_outputs(1879)) and not (layer2_outputs(1371));
    layer3_outputs(4139) <= not(layer2_outputs(3501));
    layer3_outputs(4140) <= (layer2_outputs(605)) or (layer2_outputs(1506));
    layer3_outputs(4141) <= (layer2_outputs(1234)) and not (layer2_outputs(2968));
    layer3_outputs(4142) <= '0';
    layer3_outputs(4143) <= layer2_outputs(3320);
    layer3_outputs(4144) <= (layer2_outputs(4026)) and not (layer2_outputs(1037));
    layer3_outputs(4145) <= layer2_outputs(346);
    layer3_outputs(4146) <= (layer2_outputs(4146)) and not (layer2_outputs(3831));
    layer3_outputs(4147) <= layer2_outputs(181);
    layer3_outputs(4148) <= layer2_outputs(4745);
    layer3_outputs(4149) <= '1';
    layer3_outputs(4150) <= layer2_outputs(4666);
    layer3_outputs(4151) <= (layer2_outputs(3972)) or (layer2_outputs(1803));
    layer3_outputs(4152) <= not(layer2_outputs(684)) or (layer2_outputs(4932));
    layer3_outputs(4153) <= not(layer2_outputs(3195)) or (layer2_outputs(849));
    layer3_outputs(4154) <= layer2_outputs(3214);
    layer3_outputs(4155) <= not(layer2_outputs(1973));
    layer3_outputs(4156) <= (layer2_outputs(1019)) and (layer2_outputs(1193));
    layer3_outputs(4157) <= not(layer2_outputs(1588));
    layer3_outputs(4158) <= (layer2_outputs(2376)) or (layer2_outputs(1212));
    layer3_outputs(4159) <= not(layer2_outputs(2768));
    layer3_outputs(4160) <= not((layer2_outputs(2158)) and (layer2_outputs(2788)));
    layer3_outputs(4161) <= '1';
    layer3_outputs(4162) <= '0';
    layer3_outputs(4163) <= not(layer2_outputs(1013));
    layer3_outputs(4164) <= (layer2_outputs(3056)) and (layer2_outputs(531));
    layer3_outputs(4165) <= not(layer2_outputs(1282));
    layer3_outputs(4166) <= layer2_outputs(4242);
    layer3_outputs(4167) <= not((layer2_outputs(58)) or (layer2_outputs(2149)));
    layer3_outputs(4168) <= layer2_outputs(221);
    layer3_outputs(4169) <= (layer2_outputs(2389)) and not (layer2_outputs(1226));
    layer3_outputs(4170) <= not((layer2_outputs(1477)) and (layer2_outputs(3132)));
    layer3_outputs(4171) <= not((layer2_outputs(862)) and (layer2_outputs(4272)));
    layer3_outputs(4172) <= layer2_outputs(2939);
    layer3_outputs(4173) <= not(layer2_outputs(2776)) or (layer2_outputs(2738));
    layer3_outputs(4174) <= not(layer2_outputs(3413)) or (layer2_outputs(1271));
    layer3_outputs(4175) <= (layer2_outputs(4395)) and (layer2_outputs(3306));
    layer3_outputs(4176) <= (layer2_outputs(1103)) and (layer2_outputs(4796));
    layer3_outputs(4177) <= (layer2_outputs(3981)) and not (layer2_outputs(2368));
    layer3_outputs(4178) <= '1';
    layer3_outputs(4179) <= '1';
    layer3_outputs(4180) <= (layer2_outputs(2961)) and not (layer2_outputs(700));
    layer3_outputs(4181) <= '0';
    layer3_outputs(4182) <= not(layer2_outputs(767));
    layer3_outputs(4183) <= '1';
    layer3_outputs(4184) <= layer2_outputs(2284);
    layer3_outputs(4185) <= layer2_outputs(1687);
    layer3_outputs(4186) <= layer2_outputs(4223);
    layer3_outputs(4187) <= not(layer2_outputs(4042));
    layer3_outputs(4188) <= layer2_outputs(4548);
    layer3_outputs(4189) <= not((layer2_outputs(4349)) and (layer2_outputs(603)));
    layer3_outputs(4190) <= (layer2_outputs(1848)) and (layer2_outputs(3773));
    layer3_outputs(4191) <= layer2_outputs(2697);
    layer3_outputs(4192) <= layer2_outputs(475);
    layer3_outputs(4193) <= (layer2_outputs(2585)) or (layer2_outputs(1578));
    layer3_outputs(4194) <= (layer2_outputs(5063)) xor (layer2_outputs(2674));
    layer3_outputs(4195) <= not(layer2_outputs(1317));
    layer3_outputs(4196) <= layer2_outputs(2550);
    layer3_outputs(4197) <= (layer2_outputs(4409)) and not (layer2_outputs(3764));
    layer3_outputs(4198) <= (layer2_outputs(2749)) and not (layer2_outputs(3820));
    layer3_outputs(4199) <= (layer2_outputs(4290)) and not (layer2_outputs(155));
    layer3_outputs(4200) <= not(layer2_outputs(2720));
    layer3_outputs(4201) <= layer2_outputs(3042);
    layer3_outputs(4202) <= (layer2_outputs(1499)) and not (layer2_outputs(300));
    layer3_outputs(4203) <= not(layer2_outputs(3295));
    layer3_outputs(4204) <= layer2_outputs(2432);
    layer3_outputs(4205) <= '0';
    layer3_outputs(4206) <= (layer2_outputs(4145)) and not (layer2_outputs(3557));
    layer3_outputs(4207) <= (layer2_outputs(1356)) and not (layer2_outputs(4288));
    layer3_outputs(4208) <= '1';
    layer3_outputs(4209) <= not(layer2_outputs(4728)) or (layer2_outputs(1227));
    layer3_outputs(4210) <= (layer2_outputs(740)) and not (layer2_outputs(3943));
    layer3_outputs(4211) <= layer2_outputs(4958);
    layer3_outputs(4212) <= (layer2_outputs(2379)) and not (layer2_outputs(4167));
    layer3_outputs(4213) <= not(layer2_outputs(3607));
    layer3_outputs(4214) <= not((layer2_outputs(2376)) and (layer2_outputs(3177)));
    layer3_outputs(4215) <= not((layer2_outputs(682)) or (layer2_outputs(451)));
    layer3_outputs(4216) <= not((layer2_outputs(4215)) and (layer2_outputs(4579)));
    layer3_outputs(4217) <= not(layer2_outputs(2297));
    layer3_outputs(4218) <= not((layer2_outputs(4448)) and (layer2_outputs(4904)));
    layer3_outputs(4219) <= layer2_outputs(323);
    layer3_outputs(4220) <= '0';
    layer3_outputs(4221) <= (layer2_outputs(388)) and not (layer2_outputs(1508));
    layer3_outputs(4222) <= not(layer2_outputs(4469));
    layer3_outputs(4223) <= not(layer2_outputs(3181));
    layer3_outputs(4224) <= not((layer2_outputs(627)) or (layer2_outputs(1678)));
    layer3_outputs(4225) <= (layer2_outputs(109)) xor (layer2_outputs(3521));
    layer3_outputs(4226) <= not((layer2_outputs(3745)) and (layer2_outputs(828)));
    layer3_outputs(4227) <= '0';
    layer3_outputs(4228) <= layer2_outputs(1476);
    layer3_outputs(4229) <= not(layer2_outputs(587)) or (layer2_outputs(4503));
    layer3_outputs(4230) <= not(layer2_outputs(792)) or (layer2_outputs(675));
    layer3_outputs(4231) <= '1';
    layer3_outputs(4232) <= not(layer2_outputs(4701)) or (layer2_outputs(681));
    layer3_outputs(4233) <= '1';
    layer3_outputs(4234) <= layer2_outputs(348);
    layer3_outputs(4235) <= (layer2_outputs(1951)) and not (layer2_outputs(3309));
    layer3_outputs(4236) <= layer2_outputs(3855);
    layer3_outputs(4237) <= not((layer2_outputs(741)) and (layer2_outputs(360)));
    layer3_outputs(4238) <= not((layer2_outputs(1929)) xor (layer2_outputs(4536)));
    layer3_outputs(4239) <= not(layer2_outputs(2490));
    layer3_outputs(4240) <= '0';
    layer3_outputs(4241) <= not(layer2_outputs(1545));
    layer3_outputs(4242) <= layer2_outputs(4352);
    layer3_outputs(4243) <= not(layer2_outputs(801));
    layer3_outputs(4244) <= not((layer2_outputs(3702)) and (layer2_outputs(2350)));
    layer3_outputs(4245) <= layer2_outputs(3402);
    layer3_outputs(4246) <= layer2_outputs(3460);
    layer3_outputs(4247) <= (layer2_outputs(3190)) xor (layer2_outputs(1029));
    layer3_outputs(4248) <= layer2_outputs(1624);
    layer3_outputs(4249) <= (layer2_outputs(897)) xor (layer2_outputs(1522));
    layer3_outputs(4250) <= not(layer2_outputs(2439));
    layer3_outputs(4251) <= layer2_outputs(1675);
    layer3_outputs(4252) <= (layer2_outputs(2595)) and not (layer2_outputs(1866));
    layer3_outputs(4253) <= (layer2_outputs(2889)) and not (layer2_outputs(2804));
    layer3_outputs(4254) <= layer2_outputs(4152);
    layer3_outputs(4255) <= not((layer2_outputs(2335)) and (layer2_outputs(1853)));
    layer3_outputs(4256) <= (layer2_outputs(1207)) and not (layer2_outputs(3357));
    layer3_outputs(4257) <= '0';
    layer3_outputs(4258) <= (layer2_outputs(795)) and not (layer2_outputs(2862));
    layer3_outputs(4259) <= '0';
    layer3_outputs(4260) <= (layer2_outputs(3788)) and not (layer2_outputs(1511));
    layer3_outputs(4261) <= (layer2_outputs(2676)) and not (layer2_outputs(1883));
    layer3_outputs(4262) <= not((layer2_outputs(151)) or (layer2_outputs(5011)));
    layer3_outputs(4263) <= (layer2_outputs(654)) or (layer2_outputs(2704));
    layer3_outputs(4264) <= not(layer2_outputs(3443));
    layer3_outputs(4265) <= (layer2_outputs(3143)) and not (layer2_outputs(449));
    layer3_outputs(4266) <= (layer2_outputs(1662)) and (layer2_outputs(1332));
    layer3_outputs(4267) <= not((layer2_outputs(2441)) or (layer2_outputs(2589)));
    layer3_outputs(4268) <= (layer2_outputs(3885)) or (layer2_outputs(2543));
    layer3_outputs(4269) <= not(layer2_outputs(129));
    layer3_outputs(4270) <= '1';
    layer3_outputs(4271) <= not((layer2_outputs(143)) and (layer2_outputs(1110)));
    layer3_outputs(4272) <= (layer2_outputs(1416)) or (layer2_outputs(1401));
    layer3_outputs(4273) <= not(layer2_outputs(2103)) or (layer2_outputs(2734));
    layer3_outputs(4274) <= (layer2_outputs(1173)) and (layer2_outputs(3952));
    layer3_outputs(4275) <= not((layer2_outputs(4111)) or (layer2_outputs(1540)));
    layer3_outputs(4276) <= '0';
    layer3_outputs(4277) <= (layer2_outputs(4064)) or (layer2_outputs(46));
    layer3_outputs(4278) <= not((layer2_outputs(751)) and (layer2_outputs(1906)));
    layer3_outputs(4279) <= not(layer2_outputs(3540));
    layer3_outputs(4280) <= '1';
    layer3_outputs(4281) <= not((layer2_outputs(1658)) or (layer2_outputs(4005)));
    layer3_outputs(4282) <= not((layer2_outputs(3020)) and (layer2_outputs(800)));
    layer3_outputs(4283) <= (layer2_outputs(1116)) xor (layer2_outputs(4407));
    layer3_outputs(4284) <= (layer2_outputs(1130)) or (layer2_outputs(3952));
    layer3_outputs(4285) <= not((layer2_outputs(1100)) and (layer2_outputs(2223)));
    layer3_outputs(4286) <= (layer2_outputs(4993)) xor (layer2_outputs(2756));
    layer3_outputs(4287) <= not(layer2_outputs(852)) or (layer2_outputs(826));
    layer3_outputs(4288) <= (layer2_outputs(4313)) xor (layer2_outputs(3592));
    layer3_outputs(4289) <= layer2_outputs(2869);
    layer3_outputs(4290) <= not(layer2_outputs(3359));
    layer3_outputs(4291) <= layer2_outputs(1630);
    layer3_outputs(4292) <= (layer2_outputs(3083)) xor (layer2_outputs(2529));
    layer3_outputs(4293) <= layer2_outputs(1165);
    layer3_outputs(4294) <= (layer2_outputs(1481)) or (layer2_outputs(264));
    layer3_outputs(4295) <= (layer2_outputs(1739)) or (layer2_outputs(3254));
    layer3_outputs(4296) <= '0';
    layer3_outputs(4297) <= layer2_outputs(4906);
    layer3_outputs(4298) <= layer2_outputs(1585);
    layer3_outputs(4299) <= not((layer2_outputs(1993)) or (layer2_outputs(2153)));
    layer3_outputs(4300) <= not(layer2_outputs(3372));
    layer3_outputs(4301) <= not(layer2_outputs(705)) or (layer2_outputs(2029));
    layer3_outputs(4302) <= layer2_outputs(1325);
    layer3_outputs(4303) <= '1';
    layer3_outputs(4304) <= (layer2_outputs(4087)) or (layer2_outputs(1443));
    layer3_outputs(4305) <= not(layer2_outputs(4018));
    layer3_outputs(4306) <= not(layer2_outputs(864)) or (layer2_outputs(3726));
    layer3_outputs(4307) <= (layer2_outputs(2093)) or (layer2_outputs(3756));
    layer3_outputs(4308) <= not((layer2_outputs(4133)) or (layer2_outputs(1390)));
    layer3_outputs(4309) <= not(layer2_outputs(4418));
    layer3_outputs(4310) <= not((layer2_outputs(3233)) xor (layer2_outputs(2856)));
    layer3_outputs(4311) <= not((layer2_outputs(3394)) or (layer2_outputs(3895)));
    layer3_outputs(4312) <= not(layer2_outputs(4263)) or (layer2_outputs(2014));
    layer3_outputs(4313) <= not((layer2_outputs(677)) or (layer2_outputs(4767)));
    layer3_outputs(4314) <= not(layer2_outputs(4792));
    layer3_outputs(4315) <= not(layer2_outputs(2252));
    layer3_outputs(4316) <= layer2_outputs(540);
    layer3_outputs(4317) <= not(layer2_outputs(286)) or (layer2_outputs(804));
    layer3_outputs(4318) <= not(layer2_outputs(2668)) or (layer2_outputs(2508));
    layer3_outputs(4319) <= not((layer2_outputs(2217)) xor (layer2_outputs(3471)));
    layer3_outputs(4320) <= layer2_outputs(1811);
    layer3_outputs(4321) <= not(layer2_outputs(592));
    layer3_outputs(4322) <= '1';
    layer3_outputs(4323) <= not((layer2_outputs(3614)) and (layer2_outputs(601)));
    layer3_outputs(4324) <= (layer2_outputs(467)) xor (layer2_outputs(1155));
    layer3_outputs(4325) <= (layer2_outputs(4357)) or (layer2_outputs(4382));
    layer3_outputs(4326) <= layer2_outputs(3808);
    layer3_outputs(4327) <= not(layer2_outputs(807));
    layer3_outputs(4328) <= not(layer2_outputs(2218));
    layer3_outputs(4329) <= not(layer2_outputs(1645)) or (layer2_outputs(3695));
    layer3_outputs(4330) <= (layer2_outputs(1683)) and not (layer2_outputs(3004));
    layer3_outputs(4331) <= layer2_outputs(4622);
    layer3_outputs(4332) <= (layer2_outputs(4254)) and not (layer2_outputs(1236));
    layer3_outputs(4333) <= layer2_outputs(2691);
    layer3_outputs(4334) <= not(layer2_outputs(3165));
    layer3_outputs(4335) <= not(layer2_outputs(1275)) or (layer2_outputs(2863));
    layer3_outputs(4336) <= not((layer2_outputs(1489)) and (layer2_outputs(4563)));
    layer3_outputs(4337) <= '1';
    layer3_outputs(4338) <= not(layer2_outputs(2260));
    layer3_outputs(4339) <= not((layer2_outputs(1159)) and (layer2_outputs(2747)));
    layer3_outputs(4340) <= (layer2_outputs(4967)) and (layer2_outputs(3068));
    layer3_outputs(4341) <= '0';
    layer3_outputs(4342) <= (layer2_outputs(1111)) and (layer2_outputs(4190));
    layer3_outputs(4343) <= not((layer2_outputs(7)) and (layer2_outputs(3666)));
    layer3_outputs(4344) <= (layer2_outputs(4333)) and not (layer2_outputs(1650));
    layer3_outputs(4345) <= layer2_outputs(4424);
    layer3_outputs(4346) <= not((layer2_outputs(935)) and (layer2_outputs(4453)));
    layer3_outputs(4347) <= layer2_outputs(1599);
    layer3_outputs(4348) <= (layer2_outputs(4818)) xor (layer2_outputs(3434));
    layer3_outputs(4349) <= not(layer2_outputs(2770)) or (layer2_outputs(2065));
    layer3_outputs(4350) <= layer2_outputs(4028);
    layer3_outputs(4351) <= (layer2_outputs(3016)) and not (layer2_outputs(2372));
    layer3_outputs(4352) <= '1';
    layer3_outputs(4353) <= layer2_outputs(566);
    layer3_outputs(4354) <= '1';
    layer3_outputs(4355) <= not(layer2_outputs(2760));
    layer3_outputs(4356) <= '1';
    layer3_outputs(4357) <= (layer2_outputs(1476)) and not (layer2_outputs(4808));
    layer3_outputs(4358) <= '1';
    layer3_outputs(4359) <= layer2_outputs(3282);
    layer3_outputs(4360) <= not((layer2_outputs(4560)) or (layer2_outputs(62)));
    layer3_outputs(4361) <= (layer2_outputs(4901)) and not (layer2_outputs(1383));
    layer3_outputs(4362) <= layer2_outputs(755);
    layer3_outputs(4363) <= layer2_outputs(2580);
    layer3_outputs(4364) <= layer2_outputs(2514);
    layer3_outputs(4365) <= (layer2_outputs(1980)) and not (layer2_outputs(1052));
    layer3_outputs(4366) <= (layer2_outputs(1593)) and not (layer2_outputs(245));
    layer3_outputs(4367) <= (layer2_outputs(2916)) and not (layer2_outputs(837));
    layer3_outputs(4368) <= '0';
    layer3_outputs(4369) <= not((layer2_outputs(3563)) xor (layer2_outputs(2967)));
    layer3_outputs(4370) <= '0';
    layer3_outputs(4371) <= layer2_outputs(4603);
    layer3_outputs(4372) <= not(layer2_outputs(775));
    layer3_outputs(4373) <= not(layer2_outputs(4243)) or (layer2_outputs(656));
    layer3_outputs(4374) <= layer2_outputs(4897);
    layer3_outputs(4375) <= '0';
    layer3_outputs(4376) <= '0';
    layer3_outputs(4377) <= (layer2_outputs(1815)) and (layer2_outputs(3900));
    layer3_outputs(4378) <= not(layer2_outputs(1716));
    layer3_outputs(4379) <= layer2_outputs(4484);
    layer3_outputs(4380) <= not((layer2_outputs(2690)) and (layer2_outputs(1855)));
    layer3_outputs(4381) <= '1';
    layer3_outputs(4382) <= not(layer2_outputs(2725)) or (layer2_outputs(4047));
    layer3_outputs(4383) <= not((layer2_outputs(3262)) and (layer2_outputs(4763)));
    layer3_outputs(4384) <= '1';
    layer3_outputs(4385) <= (layer2_outputs(1846)) and (layer2_outputs(3345));
    layer3_outputs(4386) <= (layer2_outputs(2108)) xor (layer2_outputs(1348));
    layer3_outputs(4387) <= (layer2_outputs(1143)) and not (layer2_outputs(2476));
    layer3_outputs(4388) <= not(layer2_outputs(2737));
    layer3_outputs(4389) <= not(layer2_outputs(3217)) or (layer2_outputs(1147));
    layer3_outputs(4390) <= not(layer2_outputs(1105)) or (layer2_outputs(977));
    layer3_outputs(4391) <= '1';
    layer3_outputs(4392) <= (layer2_outputs(3223)) or (layer2_outputs(1684));
    layer3_outputs(4393) <= (layer2_outputs(1888)) and not (layer2_outputs(3520));
    layer3_outputs(4394) <= (layer2_outputs(3373)) and not (layer2_outputs(2981));
    layer3_outputs(4395) <= (layer2_outputs(5055)) and (layer2_outputs(3190));
    layer3_outputs(4396) <= not(layer2_outputs(2353));
    layer3_outputs(4397) <= '1';
    layer3_outputs(4398) <= not(layer2_outputs(4137));
    layer3_outputs(4399) <= '0';
    layer3_outputs(4400) <= not((layer2_outputs(3445)) and (layer2_outputs(1983)));
    layer3_outputs(4401) <= not((layer2_outputs(3856)) and (layer2_outputs(1820)));
    layer3_outputs(4402) <= not(layer2_outputs(3945));
    layer3_outputs(4403) <= layer2_outputs(1898);
    layer3_outputs(4404) <= (layer2_outputs(3502)) or (layer2_outputs(579));
    layer3_outputs(4405) <= not((layer2_outputs(3075)) and (layer2_outputs(4827)));
    layer3_outputs(4406) <= not((layer2_outputs(4883)) and (layer2_outputs(2173)));
    layer3_outputs(4407) <= '1';
    layer3_outputs(4408) <= '0';
    layer3_outputs(4409) <= not(layer2_outputs(4597));
    layer3_outputs(4410) <= not(layer2_outputs(3631));
    layer3_outputs(4411) <= not(layer2_outputs(4952)) or (layer2_outputs(1189));
    layer3_outputs(4412) <= layer2_outputs(4821);
    layer3_outputs(4413) <= not(layer2_outputs(4121)) or (layer2_outputs(890));
    layer3_outputs(4414) <= (layer2_outputs(1347)) and not (layer2_outputs(1790));
    layer3_outputs(4415) <= layer2_outputs(1799);
    layer3_outputs(4416) <= (layer2_outputs(2992)) and (layer2_outputs(1150));
    layer3_outputs(4417) <= not(layer2_outputs(2457));
    layer3_outputs(4418) <= not((layer2_outputs(655)) and (layer2_outputs(2623)));
    layer3_outputs(4419) <= not(layer2_outputs(3358));
    layer3_outputs(4420) <= '1';
    layer3_outputs(4421) <= (layer2_outputs(4192)) and not (layer2_outputs(4619));
    layer3_outputs(4422) <= not((layer2_outputs(2017)) xor (layer2_outputs(2717)));
    layer3_outputs(4423) <= layer2_outputs(1795);
    layer3_outputs(4424) <= not(layer2_outputs(1467)) or (layer2_outputs(766));
    layer3_outputs(4425) <= not(layer2_outputs(1227));
    layer3_outputs(4426) <= (layer2_outputs(355)) and (layer2_outputs(3850));
    layer3_outputs(4427) <= (layer2_outputs(2698)) and not (layer2_outputs(794));
    layer3_outputs(4428) <= (layer2_outputs(5092)) xor (layer2_outputs(118));
    layer3_outputs(4429) <= layer2_outputs(5038);
    layer3_outputs(4430) <= (layer2_outputs(5027)) and (layer2_outputs(153));
    layer3_outputs(4431) <= not(layer2_outputs(1590)) or (layer2_outputs(1424));
    layer3_outputs(4432) <= (layer2_outputs(389)) xor (layer2_outputs(3992));
    layer3_outputs(4433) <= '1';
    layer3_outputs(4434) <= not((layer2_outputs(53)) or (layer2_outputs(1321)));
    layer3_outputs(4435) <= layer2_outputs(1870);
    layer3_outputs(4436) <= not(layer2_outputs(4134)) or (layer2_outputs(4802));
    layer3_outputs(4437) <= (layer2_outputs(4582)) and not (layer2_outputs(2572));
    layer3_outputs(4438) <= layer2_outputs(649);
    layer3_outputs(4439) <= not((layer2_outputs(4423)) and (layer2_outputs(667)));
    layer3_outputs(4440) <= '1';
    layer3_outputs(4441) <= not(layer2_outputs(3485));
    layer3_outputs(4442) <= not((layer2_outputs(3765)) or (layer2_outputs(865)));
    layer3_outputs(4443) <= (layer2_outputs(2511)) and not (layer2_outputs(4591));
    layer3_outputs(4444) <= (layer2_outputs(552)) or (layer2_outputs(4931));
    layer3_outputs(4445) <= '1';
    layer3_outputs(4446) <= not(layer2_outputs(311)) or (layer2_outputs(344));
    layer3_outputs(4447) <= not(layer2_outputs(82));
    layer3_outputs(4448) <= not(layer2_outputs(997));
    layer3_outputs(4449) <= '0';
    layer3_outputs(4450) <= '1';
    layer3_outputs(4451) <= '1';
    layer3_outputs(4452) <= not(layer2_outputs(1753));
    layer3_outputs(4453) <= not((layer2_outputs(2054)) and (layer2_outputs(333)));
    layer3_outputs(4454) <= not(layer2_outputs(1546));
    layer3_outputs(4455) <= not((layer2_outputs(4376)) or (layer2_outputs(108)));
    layer3_outputs(4456) <= (layer2_outputs(1323)) or (layer2_outputs(3448));
    layer3_outputs(4457) <= '1';
    layer3_outputs(4458) <= (layer2_outputs(786)) and not (layer2_outputs(2407));
    layer3_outputs(4459) <= not((layer2_outputs(2603)) or (layer2_outputs(1150)));
    layer3_outputs(4460) <= (layer2_outputs(1618)) xor (layer2_outputs(5095));
    layer3_outputs(4461) <= not((layer2_outputs(4770)) and (layer2_outputs(2170)));
    layer3_outputs(4462) <= layer2_outputs(734);
    layer3_outputs(4463) <= '1';
    layer3_outputs(4464) <= (layer2_outputs(1641)) or (layer2_outputs(2396));
    layer3_outputs(4465) <= (layer2_outputs(3777)) xor (layer2_outputs(2486));
    layer3_outputs(4466) <= not((layer2_outputs(1047)) and (layer2_outputs(3859)));
    layer3_outputs(4467) <= (layer2_outputs(3440)) and not (layer2_outputs(771));
    layer3_outputs(4468) <= not(layer2_outputs(4780));
    layer3_outputs(4469) <= not(layer2_outputs(3761)) or (layer2_outputs(2129));
    layer3_outputs(4470) <= not((layer2_outputs(2037)) and (layer2_outputs(1380)));
    layer3_outputs(4471) <= '1';
    layer3_outputs(4472) <= layer2_outputs(1564);
    layer3_outputs(4473) <= layer2_outputs(2342);
    layer3_outputs(4474) <= '0';
    layer3_outputs(4475) <= (layer2_outputs(3116)) or (layer2_outputs(130));
    layer3_outputs(4476) <= not(layer2_outputs(1312)) or (layer2_outputs(2767));
    layer3_outputs(4477) <= not((layer2_outputs(3892)) or (layer2_outputs(241)));
    layer3_outputs(4478) <= layer2_outputs(1240);
    layer3_outputs(4479) <= not(layer2_outputs(2154));
    layer3_outputs(4480) <= not(layer2_outputs(2969)) or (layer2_outputs(1022));
    layer3_outputs(4481) <= not((layer2_outputs(3137)) and (layer2_outputs(1141)));
    layer3_outputs(4482) <= layer2_outputs(5016);
    layer3_outputs(4483) <= (layer2_outputs(4740)) and not (layer2_outputs(2911));
    layer3_outputs(4484) <= not(layer2_outputs(499));
    layer3_outputs(4485) <= not((layer2_outputs(1861)) or (layer2_outputs(5100)));
    layer3_outputs(4486) <= '1';
    layer3_outputs(4487) <= not(layer2_outputs(2443)) or (layer2_outputs(4876));
    layer3_outputs(4488) <= not(layer2_outputs(3973));
    layer3_outputs(4489) <= not((layer2_outputs(5094)) and (layer2_outputs(4529)));
    layer3_outputs(4490) <= layer2_outputs(557);
    layer3_outputs(4491) <= not(layer2_outputs(5118));
    layer3_outputs(4492) <= (layer2_outputs(3815)) and (layer2_outputs(3418));
    layer3_outputs(4493) <= not(layer2_outputs(3032)) or (layer2_outputs(168));
    layer3_outputs(4494) <= not(layer2_outputs(1371)) or (layer2_outputs(1778));
    layer3_outputs(4495) <= (layer2_outputs(4311)) or (layer2_outputs(27));
    layer3_outputs(4496) <= not((layer2_outputs(412)) and (layer2_outputs(3690)));
    layer3_outputs(4497) <= not(layer2_outputs(4800));
    layer3_outputs(4498) <= not((layer2_outputs(2198)) or (layer2_outputs(3261)));
    layer3_outputs(4499) <= (layer2_outputs(832)) and not (layer2_outputs(2715));
    layer3_outputs(4500) <= not(layer2_outputs(1444)) or (layer2_outputs(3141));
    layer3_outputs(4501) <= not(layer2_outputs(2801));
    layer3_outputs(4502) <= not(layer2_outputs(2097));
    layer3_outputs(4503) <= (layer2_outputs(33)) and not (layer2_outputs(1296));
    layer3_outputs(4504) <= not((layer2_outputs(2958)) and (layer2_outputs(1519)));
    layer3_outputs(4505) <= not(layer2_outputs(427));
    layer3_outputs(4506) <= (layer2_outputs(5009)) or (layer2_outputs(3769));
    layer3_outputs(4507) <= not(layer2_outputs(3159)) or (layer2_outputs(2847));
    layer3_outputs(4508) <= (layer2_outputs(2552)) and not (layer2_outputs(4062));
    layer3_outputs(4509) <= not(layer2_outputs(4371)) or (layer2_outputs(4310));
    layer3_outputs(4510) <= not((layer2_outputs(2724)) and (layer2_outputs(2825)));
    layer3_outputs(4511) <= (layer2_outputs(3985)) and not (layer2_outputs(3814));
    layer3_outputs(4512) <= not(layer2_outputs(2132));
    layer3_outputs(4513) <= not(layer2_outputs(2837)) or (layer2_outputs(1412));
    layer3_outputs(4514) <= not((layer2_outputs(300)) or (layer2_outputs(2852)));
    layer3_outputs(4515) <= layer2_outputs(1698);
    layer3_outputs(4516) <= not(layer2_outputs(1169));
    layer3_outputs(4517) <= '0';
    layer3_outputs(4518) <= layer2_outputs(3906);
    layer3_outputs(4519) <= layer2_outputs(2288);
    layer3_outputs(4520) <= layer2_outputs(3639);
    layer3_outputs(4521) <= (layer2_outputs(2429)) or (layer2_outputs(2675));
    layer3_outputs(4522) <= not((layer2_outputs(3378)) and (layer2_outputs(2122)));
    layer3_outputs(4523) <= layer2_outputs(890);
    layer3_outputs(4524) <= (layer2_outputs(2807)) and not (layer2_outputs(4641));
    layer3_outputs(4525) <= (layer2_outputs(4161)) and not (layer2_outputs(1023));
    layer3_outputs(4526) <= (layer2_outputs(2318)) and not (layer2_outputs(3860));
    layer3_outputs(4527) <= not(layer2_outputs(2537));
    layer3_outputs(4528) <= not(layer2_outputs(1664));
    layer3_outputs(4529) <= '0';
    layer3_outputs(4530) <= not(layer2_outputs(1512)) or (layer2_outputs(633));
    layer3_outputs(4531) <= (layer2_outputs(4923)) and (layer2_outputs(255));
    layer3_outputs(4532) <= not((layer2_outputs(4669)) or (layer2_outputs(5049)));
    layer3_outputs(4533) <= (layer2_outputs(3781)) and not (layer2_outputs(4049));
    layer3_outputs(4534) <= (layer2_outputs(563)) and (layer2_outputs(2751));
    layer3_outputs(4535) <= not(layer2_outputs(3573)) or (layer2_outputs(1216));
    layer3_outputs(4536) <= not(layer2_outputs(239)) or (layer2_outputs(3728));
    layer3_outputs(4537) <= layer2_outputs(3480);
    layer3_outputs(4538) <= '0';
    layer3_outputs(4539) <= '1';
    layer3_outputs(4540) <= (layer2_outputs(2415)) and not (layer2_outputs(3087));
    layer3_outputs(4541) <= layer2_outputs(3723);
    layer3_outputs(4542) <= not((layer2_outputs(3240)) and (layer2_outputs(1309)));
    layer3_outputs(4543) <= (layer2_outputs(3294)) or (layer2_outputs(4055));
    layer3_outputs(4544) <= not(layer2_outputs(3127));
    layer3_outputs(4545) <= layer2_outputs(306);
    layer3_outputs(4546) <= not(layer2_outputs(143)) or (layer2_outputs(1090));
    layer3_outputs(4547) <= (layer2_outputs(3385)) xor (layer2_outputs(1518));
    layer3_outputs(4548) <= not((layer2_outputs(1606)) or (layer2_outputs(1316)));
    layer3_outputs(4549) <= (layer2_outputs(3802)) or (layer2_outputs(1583));
    layer3_outputs(4550) <= (layer2_outputs(1760)) or (layer2_outputs(976));
    layer3_outputs(4551) <= '0';
    layer3_outputs(4552) <= (layer2_outputs(892)) and not (layer2_outputs(308));
    layer3_outputs(4553) <= layer2_outputs(4119);
    layer3_outputs(4554) <= not((layer2_outputs(4430)) xor (layer2_outputs(4161)));
    layer3_outputs(4555) <= (layer2_outputs(591)) or (layer2_outputs(3366));
    layer3_outputs(4556) <= layer2_outputs(4917);
    layer3_outputs(4557) <= not((layer2_outputs(2539)) xor (layer2_outputs(755)));
    layer3_outputs(4558) <= '0';
    layer3_outputs(4559) <= not((layer2_outputs(224)) and (layer2_outputs(5041)));
    layer3_outputs(4560) <= not(layer2_outputs(409));
    layer3_outputs(4561) <= layer2_outputs(1577);
    layer3_outputs(4562) <= layer2_outputs(548);
    layer3_outputs(4563) <= not((layer2_outputs(492)) or (layer2_outputs(1786)));
    layer3_outputs(4564) <= '1';
    layer3_outputs(4565) <= '1';
    layer3_outputs(4566) <= layer2_outputs(4940);
    layer3_outputs(4567) <= layer2_outputs(1787);
    layer3_outputs(4568) <= layer2_outputs(4127);
    layer3_outputs(4569) <= layer2_outputs(2910);
    layer3_outputs(4570) <= (layer2_outputs(4828)) and (layer2_outputs(3043));
    layer3_outputs(4571) <= (layer2_outputs(4801)) or (layer2_outputs(4021));
    layer3_outputs(4572) <= not((layer2_outputs(4075)) and (layer2_outputs(1095)));
    layer3_outputs(4573) <= not(layer2_outputs(764));
    layer3_outputs(4574) <= '0';
    layer3_outputs(4575) <= layer2_outputs(2879);
    layer3_outputs(4576) <= not((layer2_outputs(3912)) or (layer2_outputs(403)));
    layer3_outputs(4577) <= (layer2_outputs(1206)) and not (layer2_outputs(3653));
    layer3_outputs(4578) <= layer2_outputs(825);
    layer3_outputs(4579) <= layer2_outputs(2310);
    layer3_outputs(4580) <= (layer2_outputs(325)) and (layer2_outputs(453));
    layer3_outputs(4581) <= (layer2_outputs(851)) and not (layer2_outputs(1154));
    layer3_outputs(4582) <= '1';
    layer3_outputs(4583) <= (layer2_outputs(962)) and not (layer2_outputs(1220));
    layer3_outputs(4584) <= not(layer2_outputs(1893));
    layer3_outputs(4585) <= not(layer2_outputs(1590));
    layer3_outputs(4586) <= (layer2_outputs(4663)) and not (layer2_outputs(2312));
    layer3_outputs(4587) <= '1';
    layer3_outputs(4588) <= (layer2_outputs(1483)) and not (layer2_outputs(4234));
    layer3_outputs(4589) <= (layer2_outputs(1635)) and not (layer2_outputs(2635));
    layer3_outputs(4590) <= '0';
    layer3_outputs(4591) <= (layer2_outputs(587)) or (layer2_outputs(3083));
    layer3_outputs(4592) <= not(layer2_outputs(1072));
    layer3_outputs(4593) <= not(layer2_outputs(712));
    layer3_outputs(4594) <= (layer2_outputs(737)) and not (layer2_outputs(901));
    layer3_outputs(4595) <= not(layer2_outputs(5040));
    layer3_outputs(4596) <= (layer2_outputs(2594)) and not (layer2_outputs(3337));
    layer3_outputs(4597) <= not(layer2_outputs(2827)) or (layer2_outputs(974));
    layer3_outputs(4598) <= not(layer2_outputs(2535));
    layer3_outputs(4599) <= not(layer2_outputs(4965));
    layer3_outputs(4600) <= (layer2_outputs(1065)) and not (layer2_outputs(3609));
    layer3_outputs(4601) <= '1';
    layer3_outputs(4602) <= layer2_outputs(1793);
    layer3_outputs(4603) <= layer2_outputs(642);
    layer3_outputs(4604) <= '0';
    layer3_outputs(4605) <= (layer2_outputs(2650)) and not (layer2_outputs(3947));
    layer3_outputs(4606) <= (layer2_outputs(3806)) and not (layer2_outputs(4033));
    layer3_outputs(4607) <= (layer2_outputs(5042)) and not (layer2_outputs(4232));
    layer3_outputs(4608) <= not((layer2_outputs(4406)) and (layer2_outputs(3454)));
    layer3_outputs(4609) <= not(layer2_outputs(173)) or (layer2_outputs(4691));
    layer3_outputs(4610) <= (layer2_outputs(4911)) or (layer2_outputs(3492));
    layer3_outputs(4611) <= layer2_outputs(371);
    layer3_outputs(4612) <= (layer2_outputs(4220)) or (layer2_outputs(1904));
    layer3_outputs(4613) <= (layer2_outputs(607)) and not (layer2_outputs(4205));
    layer3_outputs(4614) <= (layer2_outputs(4417)) or (layer2_outputs(4523));
    layer3_outputs(4615) <= not((layer2_outputs(2269)) xor (layer2_outputs(3662)));
    layer3_outputs(4616) <= (layer2_outputs(3870)) and not (layer2_outputs(517));
    layer3_outputs(4617) <= (layer2_outputs(4067)) and not (layer2_outputs(1403));
    layer3_outputs(4618) <= not(layer2_outputs(4219));
    layer3_outputs(4619) <= (layer2_outputs(3014)) and (layer2_outputs(4305));
    layer3_outputs(4620) <= not(layer2_outputs(27));
    layer3_outputs(4621) <= '0';
    layer3_outputs(4622) <= '0';
    layer3_outputs(4623) <= (layer2_outputs(779)) and (layer2_outputs(4288));
    layer3_outputs(4624) <= not(layer2_outputs(2685));
    layer3_outputs(4625) <= not((layer2_outputs(1450)) and (layer2_outputs(4038)));
    layer3_outputs(4626) <= not(layer2_outputs(1497));
    layer3_outputs(4627) <= (layer2_outputs(2616)) and not (layer2_outputs(2152));
    layer3_outputs(4628) <= not(layer2_outputs(5096)) or (layer2_outputs(3570));
    layer3_outputs(4629) <= not(layer2_outputs(109)) or (layer2_outputs(1377));
    layer3_outputs(4630) <= not(layer2_outputs(2307));
    layer3_outputs(4631) <= layer2_outputs(281);
    layer3_outputs(4632) <= not(layer2_outputs(801));
    layer3_outputs(4633) <= not((layer2_outputs(2557)) xor (layer2_outputs(330)));
    layer3_outputs(4634) <= (layer2_outputs(1660)) or (layer2_outputs(4058));
    layer3_outputs(4635) <= layer2_outputs(5074);
    layer3_outputs(4636) <= not(layer2_outputs(736));
    layer3_outputs(4637) <= '1';
    layer3_outputs(4638) <= '1';
    layer3_outputs(4639) <= (layer2_outputs(4384)) or (layer2_outputs(1957));
    layer3_outputs(4640) <= layer2_outputs(2245);
    layer3_outputs(4641) <= layer2_outputs(3365);
    layer3_outputs(4642) <= '1';
    layer3_outputs(4643) <= '0';
    layer3_outputs(4644) <= layer2_outputs(2782);
    layer3_outputs(4645) <= (layer2_outputs(1179)) and (layer2_outputs(2285));
    layer3_outputs(4646) <= layer2_outputs(3012);
    layer3_outputs(4647) <= not(layer2_outputs(3876)) or (layer2_outputs(3680));
    layer3_outputs(4648) <= not((layer2_outputs(3572)) and (layer2_outputs(5022)));
    layer3_outputs(4649) <= (layer2_outputs(2466)) and not (layer2_outputs(3070));
    layer3_outputs(4650) <= not((layer2_outputs(441)) xor (layer2_outputs(3990)));
    layer3_outputs(4651) <= not(layer2_outputs(2427)) or (layer2_outputs(1483));
    layer3_outputs(4652) <= not((layer2_outputs(2971)) or (layer2_outputs(3149)));
    layer3_outputs(4653) <= layer2_outputs(15);
    layer3_outputs(4654) <= not((layer2_outputs(1255)) or (layer2_outputs(393)));
    layer3_outputs(4655) <= (layer2_outputs(4994)) and not (layer2_outputs(1496));
    layer3_outputs(4656) <= '1';
    layer3_outputs(4657) <= (layer2_outputs(4781)) and not (layer2_outputs(3063));
    layer3_outputs(4658) <= layer2_outputs(4223);
    layer3_outputs(4659) <= (layer2_outputs(176)) or (layer2_outputs(973));
    layer3_outputs(4660) <= not((layer2_outputs(2755)) and (layer2_outputs(2521)));
    layer3_outputs(4661) <= not(layer2_outputs(2168));
    layer3_outputs(4662) <= layer2_outputs(2305);
    layer3_outputs(4663) <= not((layer2_outputs(3704)) or (layer2_outputs(1459)));
    layer3_outputs(4664) <= (layer2_outputs(2708)) and not (layer2_outputs(917));
    layer3_outputs(4665) <= layer2_outputs(637);
    layer3_outputs(4666) <= '0';
    layer3_outputs(4667) <= (layer2_outputs(3495)) xor (layer2_outputs(621));
    layer3_outputs(4668) <= (layer2_outputs(2075)) and not (layer2_outputs(4739));
    layer3_outputs(4669) <= '0';
    layer3_outputs(4670) <= (layer2_outputs(1509)) or (layer2_outputs(1509));
    layer3_outputs(4671) <= not(layer2_outputs(3262));
    layer3_outputs(4672) <= '0';
    layer3_outputs(4673) <= not(layer2_outputs(2904)) or (layer2_outputs(3444));
    layer3_outputs(4674) <= (layer2_outputs(912)) and not (layer2_outputs(4671));
    layer3_outputs(4675) <= not((layer2_outputs(393)) or (layer2_outputs(3611)));
    layer3_outputs(4676) <= '0';
    layer3_outputs(4677) <= not((layer2_outputs(31)) or (layer2_outputs(3494)));
    layer3_outputs(4678) <= not((layer2_outputs(4241)) and (layer2_outputs(394)));
    layer3_outputs(4679) <= '0';
    layer3_outputs(4680) <= not(layer2_outputs(5109)) or (layer2_outputs(4174));
    layer3_outputs(4681) <= layer2_outputs(4448);
    layer3_outputs(4682) <= not(layer2_outputs(644)) or (layer2_outputs(177));
    layer3_outputs(4683) <= '0';
    layer3_outputs(4684) <= not(layer2_outputs(902)) or (layer2_outputs(4896));
    layer3_outputs(4685) <= '0';
    layer3_outputs(4686) <= not(layer2_outputs(2257));
    layer3_outputs(4687) <= not(layer2_outputs(5068)) or (layer2_outputs(652));
    layer3_outputs(4688) <= layer2_outputs(3381);
    layer3_outputs(4689) <= '1';
    layer3_outputs(4690) <= not(layer2_outputs(4073));
    layer3_outputs(4691) <= not((layer2_outputs(1474)) and (layer2_outputs(3623)));
    layer3_outputs(4692) <= layer2_outputs(377);
    layer3_outputs(4693) <= (layer2_outputs(2831)) and not (layer2_outputs(1573));
    layer3_outputs(4694) <= layer2_outputs(1818);
    layer3_outputs(4695) <= layer2_outputs(3774);
    layer3_outputs(4696) <= (layer2_outputs(4571)) and (layer2_outputs(113));
    layer3_outputs(4697) <= not(layer2_outputs(4227));
    layer3_outputs(4698) <= layer2_outputs(2417);
    layer3_outputs(4699) <= (layer2_outputs(2521)) and not (layer2_outputs(947));
    layer3_outputs(4700) <= (layer2_outputs(2526)) and not (layer2_outputs(3719));
    layer3_outputs(4701) <= not(layer2_outputs(4803));
    layer3_outputs(4702) <= layer2_outputs(3679);
    layer3_outputs(4703) <= (layer2_outputs(2491)) and not (layer2_outputs(4389));
    layer3_outputs(4704) <= layer2_outputs(1);
    layer3_outputs(4705) <= layer2_outputs(3997);
    layer3_outputs(4706) <= (layer2_outputs(1995)) or (layer2_outputs(2924));
    layer3_outputs(4707) <= '1';
    layer3_outputs(4708) <= '0';
    layer3_outputs(4709) <= (layer2_outputs(282)) and not (layer2_outputs(3325));
    layer3_outputs(4710) <= (layer2_outputs(4790)) or (layer2_outputs(2674));
    layer3_outputs(4711) <= (layer2_outputs(2933)) and not (layer2_outputs(3667));
    layer3_outputs(4712) <= not(layer2_outputs(986));
    layer3_outputs(4713) <= not(layer2_outputs(4701)) or (layer2_outputs(1190));
    layer3_outputs(4714) <= layer2_outputs(814);
    layer3_outputs(4715) <= layer2_outputs(540);
    layer3_outputs(4716) <= not((layer2_outputs(3290)) xor (layer2_outputs(2525)));
    layer3_outputs(4717) <= not(layer2_outputs(2622));
    layer3_outputs(4718) <= not(layer2_outputs(1551));
    layer3_outputs(4719) <= not(layer2_outputs(3194));
    layer3_outputs(4720) <= not((layer2_outputs(4064)) and (layer2_outputs(2137)));
    layer3_outputs(4721) <= not(layer2_outputs(2245));
    layer3_outputs(4722) <= not((layer2_outputs(3696)) and (layer2_outputs(927)));
    layer3_outputs(4723) <= not(layer2_outputs(1841)) or (layer2_outputs(3675));
    layer3_outputs(4724) <= (layer2_outputs(2129)) and not (layer2_outputs(3176));
    layer3_outputs(4725) <= layer2_outputs(288);
    layer3_outputs(4726) <= (layer2_outputs(4598)) and (layer2_outputs(1624));
    layer3_outputs(4727) <= '0';
    layer3_outputs(4728) <= (layer2_outputs(261)) and not (layer2_outputs(2262));
    layer3_outputs(4729) <= layer2_outputs(4550);
    layer3_outputs(4730) <= '0';
    layer3_outputs(4731) <= '1';
    layer3_outputs(4732) <= (layer2_outputs(4930)) and not (layer2_outputs(820));
    layer3_outputs(4733) <= (layer2_outputs(4225)) or (layer2_outputs(4331));
    layer3_outputs(4734) <= not((layer2_outputs(2271)) and (layer2_outputs(2959)));
    layer3_outputs(4735) <= not((layer2_outputs(901)) or (layer2_outputs(4869)));
    layer3_outputs(4736) <= layer2_outputs(175);
    layer3_outputs(4737) <= (layer2_outputs(3995)) or (layer2_outputs(2382));
    layer3_outputs(4738) <= '1';
    layer3_outputs(4739) <= not(layer2_outputs(3439));
    layer3_outputs(4740) <= (layer2_outputs(2522)) and not (layer2_outputs(1880));
    layer3_outputs(4741) <= not(layer2_outputs(3578));
    layer3_outputs(4742) <= not(layer2_outputs(2636)) or (layer2_outputs(217));
    layer3_outputs(4743) <= (layer2_outputs(5112)) and not (layer2_outputs(1773));
    layer3_outputs(4744) <= layer2_outputs(26);
    layer3_outputs(4745) <= (layer2_outputs(1648)) or (layer2_outputs(592));
    layer3_outputs(4746) <= (layer2_outputs(2352)) and (layer2_outputs(1639));
    layer3_outputs(4747) <= '0';
    layer3_outputs(4748) <= '1';
    layer3_outputs(4749) <= not(layer2_outputs(4246));
    layer3_outputs(4750) <= not((layer2_outputs(100)) xor (layer2_outputs(2552)));
    layer3_outputs(4751) <= (layer2_outputs(2795)) and not (layer2_outputs(1782));
    layer3_outputs(4752) <= (layer2_outputs(1426)) or (layer2_outputs(2598));
    layer3_outputs(4753) <= not(layer2_outputs(3515));
    layer3_outputs(4754) <= not(layer2_outputs(3431)) or (layer2_outputs(274));
    layer3_outputs(4755) <= not(layer2_outputs(1372));
    layer3_outputs(4756) <= not((layer2_outputs(3482)) or (layer2_outputs(1780)));
    layer3_outputs(4757) <= layer2_outputs(1210);
    layer3_outputs(4758) <= '1';
    layer3_outputs(4759) <= (layer2_outputs(2728)) and (layer2_outputs(67));
    layer3_outputs(4760) <= not(layer2_outputs(4450)) or (layer2_outputs(4077));
    layer3_outputs(4761) <= not((layer2_outputs(5044)) xor (layer2_outputs(3897)));
    layer3_outputs(4762) <= '0';
    layer3_outputs(4763) <= not(layer2_outputs(3667));
    layer3_outputs(4764) <= layer2_outputs(3280);
    layer3_outputs(4765) <= not((layer2_outputs(102)) xor (layer2_outputs(4267)));
    layer3_outputs(4766) <= not(layer2_outputs(2973));
    layer3_outputs(4767) <= (layer2_outputs(788)) or (layer2_outputs(4757));
    layer3_outputs(4768) <= not((layer2_outputs(1472)) or (layer2_outputs(1902)));
    layer3_outputs(4769) <= layer2_outputs(4309);
    layer3_outputs(4770) <= layer2_outputs(1168);
    layer3_outputs(4771) <= not(layer2_outputs(4874)) or (layer2_outputs(3141));
    layer3_outputs(4772) <= not(layer2_outputs(3125));
    layer3_outputs(4773) <= layer2_outputs(1755);
    layer3_outputs(4774) <= not(layer2_outputs(1863));
    layer3_outputs(4775) <= not(layer2_outputs(2308)) or (layer2_outputs(2930));
    layer3_outputs(4776) <= '1';
    layer3_outputs(4777) <= not(layer2_outputs(5052));
    layer3_outputs(4778) <= not(layer2_outputs(495)) or (layer2_outputs(989));
    layer3_outputs(4779) <= layer2_outputs(2337);
    layer3_outputs(4780) <= (layer2_outputs(1637)) and not (layer2_outputs(3884));
    layer3_outputs(4781) <= '0';
    layer3_outputs(4782) <= layer2_outputs(1676);
    layer3_outputs(4783) <= not((layer2_outputs(971)) or (layer2_outputs(4854)));
    layer3_outputs(4784) <= (layer2_outputs(3490)) and not (layer2_outputs(2036));
    layer3_outputs(4785) <= not(layer2_outputs(40));
    layer3_outputs(4786) <= layer2_outputs(2840);
    layer3_outputs(4787) <= '1';
    layer3_outputs(4788) <= (layer2_outputs(4508)) and not (layer2_outputs(843));
    layer3_outputs(4789) <= not(layer2_outputs(2707));
    layer3_outputs(4790) <= not(layer2_outputs(2873));
    layer3_outputs(4791) <= not(layer2_outputs(2823));
    layer3_outputs(4792) <= (layer2_outputs(3617)) or (layer2_outputs(3738));
    layer3_outputs(4793) <= (layer2_outputs(3966)) and not (layer2_outputs(4416));
    layer3_outputs(4794) <= layer2_outputs(3314);
    layer3_outputs(4795) <= layer2_outputs(3710);
    layer3_outputs(4796) <= not(layer2_outputs(332)) or (layer2_outputs(906));
    layer3_outputs(4797) <= not(layer2_outputs(2328));
    layer3_outputs(4798) <= layer2_outputs(1576);
    layer3_outputs(4799) <= '1';
    layer3_outputs(4800) <= not(layer2_outputs(4386)) or (layer2_outputs(2639));
    layer3_outputs(4801) <= layer2_outputs(356);
    layer3_outputs(4802) <= '1';
    layer3_outputs(4803) <= (layer2_outputs(2281)) or (layer2_outputs(2703));
    layer3_outputs(4804) <= not(layer2_outputs(1581)) or (layer2_outputs(3858));
    layer3_outputs(4805) <= (layer2_outputs(3071)) and not (layer2_outputs(805));
    layer3_outputs(4806) <= not(layer2_outputs(4860)) or (layer2_outputs(4767));
    layer3_outputs(4807) <= (layer2_outputs(2916)) and (layer2_outputs(881));
    layer3_outputs(4808) <= '0';
    layer3_outputs(4809) <= not(layer2_outputs(2943));
    layer3_outputs(4810) <= not(layer2_outputs(4133));
    layer3_outputs(4811) <= (layer2_outputs(4832)) and not (layer2_outputs(1558));
    layer3_outputs(4812) <= not(layer2_outputs(2477));
    layer3_outputs(4813) <= layer2_outputs(856);
    layer3_outputs(4814) <= (layer2_outputs(2895)) and not (layer2_outputs(2926));
    layer3_outputs(4815) <= (layer2_outputs(3145)) xor (layer2_outputs(2476));
    layer3_outputs(4816) <= (layer2_outputs(1784)) and not (layer2_outputs(4413));
    layer3_outputs(4817) <= not(layer2_outputs(4378)) or (layer2_outputs(2989));
    layer3_outputs(4818) <= (layer2_outputs(2267)) and not (layer2_outputs(879));
    layer3_outputs(4819) <= not(layer2_outputs(4089)) or (layer2_outputs(804));
    layer3_outputs(4820) <= '0';
    layer3_outputs(4821) <= not(layer2_outputs(3527));
    layer3_outputs(4822) <= layer2_outputs(1321);
    layer3_outputs(4823) <= '0';
    layer3_outputs(4824) <= not(layer2_outputs(1840));
    layer3_outputs(4825) <= not(layer2_outputs(3340));
    layer3_outputs(4826) <= not((layer2_outputs(2934)) and (layer2_outputs(1128)));
    layer3_outputs(4827) <= (layer2_outputs(4915)) or (layer2_outputs(611));
    layer3_outputs(4828) <= '1';
    layer3_outputs(4829) <= (layer2_outputs(761)) or (layer2_outputs(2680));
    layer3_outputs(4830) <= layer2_outputs(1451);
    layer3_outputs(4831) <= layer2_outputs(4814);
    layer3_outputs(4832) <= (layer2_outputs(4397)) and not (layer2_outputs(2999));
    layer3_outputs(4833) <= (layer2_outputs(47)) and not (layer2_outputs(1133));
    layer3_outputs(4834) <= not(layer2_outputs(1838)) or (layer2_outputs(3225));
    layer3_outputs(4835) <= not(layer2_outputs(1178));
    layer3_outputs(4836) <= layer2_outputs(1756);
    layer3_outputs(4837) <= not((layer2_outputs(3990)) and (layer2_outputs(966)));
    layer3_outputs(4838) <= layer2_outputs(490);
    layer3_outputs(4839) <= '1';
    layer3_outputs(4840) <= (layer2_outputs(2663)) and (layer2_outputs(4007));
    layer3_outputs(4841) <= (layer2_outputs(4030)) and not (layer2_outputs(4248));
    layer3_outputs(4842) <= layer2_outputs(1385);
    layer3_outputs(4843) <= not(layer2_outputs(4533)) or (layer2_outputs(2110));
    layer3_outputs(4844) <= (layer2_outputs(1945)) and not (layer2_outputs(4955));
    layer3_outputs(4845) <= (layer2_outputs(3409)) xor (layer2_outputs(418));
    layer3_outputs(4846) <= not(layer2_outputs(287)) or (layer2_outputs(2105));
    layer3_outputs(4847) <= not((layer2_outputs(1408)) or (layer2_outputs(4498)));
    layer3_outputs(4848) <= (layer2_outputs(1058)) and (layer2_outputs(4463));
    layer3_outputs(4849) <= layer2_outputs(3342);
    layer3_outputs(4850) <= not((layer2_outputs(1020)) xor (layer2_outputs(4524)));
    layer3_outputs(4851) <= layer2_outputs(4070);
    layer3_outputs(4852) <= not(layer2_outputs(3456)) or (layer2_outputs(1000));
    layer3_outputs(4853) <= (layer2_outputs(744)) xor (layer2_outputs(4329));
    layer3_outputs(4854) <= not(layer2_outputs(5008));
    layer3_outputs(4855) <= not(layer2_outputs(2706));
    layer3_outputs(4856) <= not(layer2_outputs(951));
    layer3_outputs(4857) <= (layer2_outputs(2657)) and not (layer2_outputs(2485));
    layer3_outputs(4858) <= not(layer2_outputs(4596)) or (layer2_outputs(4631));
    layer3_outputs(4859) <= layer2_outputs(1632);
    layer3_outputs(4860) <= (layer2_outputs(2207)) and not (layer2_outputs(3445));
    layer3_outputs(4861) <= layer2_outputs(1448);
    layer3_outputs(4862) <= not(layer2_outputs(4079));
    layer3_outputs(4863) <= (layer2_outputs(4858)) and not (layer2_outputs(3960));
    layer3_outputs(4864) <= '1';
    layer3_outputs(4865) <= not(layer2_outputs(1809));
    layer3_outputs(4866) <= (layer2_outputs(4508)) and (layer2_outputs(308));
    layer3_outputs(4867) <= layer2_outputs(3703);
    layer3_outputs(4868) <= not(layer2_outputs(2640));
    layer3_outputs(4869) <= (layer2_outputs(106)) and (layer2_outputs(1263));
    layer3_outputs(4870) <= not(layer2_outputs(579)) or (layer2_outputs(2444));
    layer3_outputs(4871) <= not((layer2_outputs(4255)) xor (layer2_outputs(752)));
    layer3_outputs(4872) <= (layer2_outputs(1364)) and not (layer2_outputs(991));
    layer3_outputs(4873) <= (layer2_outputs(1457)) and not (layer2_outputs(5054));
    layer3_outputs(4874) <= (layer2_outputs(179)) or (layer2_outputs(2699));
    layer3_outputs(4875) <= '1';
    layer3_outputs(4876) <= (layer2_outputs(3747)) or (layer2_outputs(1641));
    layer3_outputs(4877) <= (layer2_outputs(1580)) or (layer2_outputs(1222));
    layer3_outputs(4878) <= layer2_outputs(2736);
    layer3_outputs(4879) <= layer2_outputs(2043);
    layer3_outputs(4880) <= not(layer2_outputs(164)) or (layer2_outputs(908));
    layer3_outputs(4881) <= not(layer2_outputs(2026));
    layer3_outputs(4882) <= '0';
    layer3_outputs(4883) <= layer2_outputs(3395);
    layer3_outputs(4884) <= '1';
    layer3_outputs(4885) <= (layer2_outputs(3746)) and (layer2_outputs(2293));
    layer3_outputs(4886) <= '0';
    layer3_outputs(4887) <= layer2_outputs(528);
    layer3_outputs(4888) <= not(layer2_outputs(3162));
    layer3_outputs(4889) <= (layer2_outputs(42)) and (layer2_outputs(1477));
    layer3_outputs(4890) <= (layer2_outputs(1003)) and (layer2_outputs(848));
    layer3_outputs(4891) <= not(layer2_outputs(462));
    layer3_outputs(4892) <= layer2_outputs(4229);
    layer3_outputs(4893) <= (layer2_outputs(4953)) and not (layer2_outputs(5062));
    layer3_outputs(4894) <= '1';
    layer3_outputs(4895) <= (layer2_outputs(4594)) and (layer2_outputs(2824));
    layer3_outputs(4896) <= layer2_outputs(4411);
    layer3_outputs(4897) <= (layer2_outputs(3194)) and not (layer2_outputs(2653));
    layer3_outputs(4898) <= not(layer2_outputs(4898));
    layer3_outputs(4899) <= '1';
    layer3_outputs(4900) <= '0';
    layer3_outputs(4901) <= layer2_outputs(2071);
    layer3_outputs(4902) <= not(layer2_outputs(5091)) or (layer2_outputs(2084));
    layer3_outputs(4903) <= layer2_outputs(4137);
    layer3_outputs(4904) <= '1';
    layer3_outputs(4905) <= '0';
    layer3_outputs(4906) <= not(layer2_outputs(1013)) or (layer2_outputs(842));
    layer3_outputs(4907) <= (layer2_outputs(1517)) and not (layer2_outputs(735));
    layer3_outputs(4908) <= (layer2_outputs(1231)) and not (layer2_outputs(977));
    layer3_outputs(4909) <= (layer2_outputs(4515)) or (layer2_outputs(1080));
    layer3_outputs(4910) <= (layer2_outputs(1415)) and not (layer2_outputs(2788));
    layer3_outputs(4911) <= not((layer2_outputs(1906)) and (layer2_outputs(1056)));
    layer3_outputs(4912) <= layer2_outputs(1218);
    layer3_outputs(4913) <= not(layer2_outputs(2292));
    layer3_outputs(4914) <= not((layer2_outputs(3928)) or (layer2_outputs(984)));
    layer3_outputs(4915) <= '1';
    layer3_outputs(4916) <= (layer2_outputs(4462)) and (layer2_outputs(631));
    layer3_outputs(4917) <= '1';
    layer3_outputs(4918) <= (layer2_outputs(1139)) and not (layer2_outputs(3091));
    layer3_outputs(4919) <= layer2_outputs(4645);
    layer3_outputs(4920) <= (layer2_outputs(4858)) and (layer2_outputs(1157));
    layer3_outputs(4921) <= (layer2_outputs(4203)) and (layer2_outputs(4898));
    layer3_outputs(4922) <= '0';
    layer3_outputs(4923) <= '0';
    layer3_outputs(4924) <= (layer2_outputs(1225)) and not (layer2_outputs(1720));
    layer3_outputs(4925) <= not(layer2_outputs(3602));
    layer3_outputs(4926) <= not(layer2_outputs(829));
    layer3_outputs(4927) <= (layer2_outputs(3323)) and not (layer2_outputs(202));
    layer3_outputs(4928) <= not(layer2_outputs(4857));
    layer3_outputs(4929) <= not(layer2_outputs(1372)) or (layer2_outputs(63));
    layer3_outputs(4930) <= not(layer2_outputs(1163));
    layer3_outputs(4931) <= (layer2_outputs(1852)) and not (layer2_outputs(337));
    layer3_outputs(4932) <= (layer2_outputs(3961)) and not (layer2_outputs(2118));
    layer3_outputs(4933) <= (layer2_outputs(1755)) or (layer2_outputs(1724));
    layer3_outputs(4934) <= not(layer2_outputs(690)) or (layer2_outputs(2315));
    layer3_outputs(4935) <= not((layer2_outputs(5005)) and (layer2_outputs(97)));
    layer3_outputs(4936) <= layer2_outputs(3522);
    layer3_outputs(4937) <= not(layer2_outputs(3033));
    layer3_outputs(4938) <= not((layer2_outputs(4044)) and (layer2_outputs(2237)));
    layer3_outputs(4939) <= not(layer2_outputs(3634)) or (layer2_outputs(1581));
    layer3_outputs(4940) <= '1';
    layer3_outputs(4941) <= (layer2_outputs(889)) and not (layer2_outputs(2974));
    layer3_outputs(4942) <= not(layer2_outputs(3691)) or (layer2_outputs(1833));
    layer3_outputs(4943) <= not(layer2_outputs(749));
    layer3_outputs(4944) <= (layer2_outputs(2475)) or (layer2_outputs(988));
    layer3_outputs(4945) <= '1';
    layer3_outputs(4946) <= (layer2_outputs(4086)) and not (layer2_outputs(4824));
    layer3_outputs(4947) <= layer2_outputs(216);
    layer3_outputs(4948) <= layer2_outputs(3326);
    layer3_outputs(4949) <= layer2_outputs(1900);
    layer3_outputs(4950) <= '1';
    layer3_outputs(4951) <= not(layer2_outputs(3786));
    layer3_outputs(4952) <= layer2_outputs(4535);
    layer3_outputs(4953) <= (layer2_outputs(4423)) xor (layer2_outputs(1759));
    layer3_outputs(4954) <= '0';
    layer3_outputs(4955) <= '0';
    layer3_outputs(4956) <= layer2_outputs(368);
    layer3_outputs(4957) <= layer2_outputs(3203);
    layer3_outputs(4958) <= (layer2_outputs(1692)) and (layer2_outputs(5066));
    layer3_outputs(4959) <= not(layer2_outputs(1099));
    layer3_outputs(4960) <= layer2_outputs(3391);
    layer3_outputs(4961) <= (layer2_outputs(4398)) and (layer2_outputs(3968));
    layer3_outputs(4962) <= '0';
    layer3_outputs(4963) <= not(layer2_outputs(146));
    layer3_outputs(4964) <= (layer2_outputs(1608)) and not (layer2_outputs(2881));
    layer3_outputs(4965) <= (layer2_outputs(688)) xor (layer2_outputs(1615));
    layer3_outputs(4966) <= (layer2_outputs(565)) and not (layer2_outputs(88));
    layer3_outputs(4967) <= (layer2_outputs(2617)) and not (layer2_outputs(4998));
    layer3_outputs(4968) <= not((layer2_outputs(4629)) or (layer2_outputs(4646)));
    layer3_outputs(4969) <= '0';
    layer3_outputs(4970) <= '0';
    layer3_outputs(4971) <= (layer2_outputs(1659)) and not (layer2_outputs(1575));
    layer3_outputs(4972) <= layer2_outputs(4180);
    layer3_outputs(4973) <= not(layer2_outputs(4109));
    layer3_outputs(4974) <= not(layer2_outputs(1201));
    layer3_outputs(4975) <= layer2_outputs(1846);
    layer3_outputs(4976) <= not(layer2_outputs(4050));
    layer3_outputs(4977) <= (layer2_outputs(2877)) and (layer2_outputs(2022));
    layer3_outputs(4978) <= layer2_outputs(2574);
    layer3_outputs(4979) <= layer2_outputs(642);
    layer3_outputs(4980) <= not(layer2_outputs(1504));
    layer3_outputs(4981) <= not(layer2_outputs(4290)) or (layer2_outputs(3865));
    layer3_outputs(4982) <= not(layer2_outputs(4485));
    layer3_outputs(4983) <= not(layer2_outputs(2886));
    layer3_outputs(4984) <= not((layer2_outputs(1270)) xor (layer2_outputs(2270)));
    layer3_outputs(4985) <= '1';
    layer3_outputs(4986) <= not(layer2_outputs(4422)) or (layer2_outputs(1726));
    layer3_outputs(4987) <= not(layer2_outputs(2088)) or (layer2_outputs(4500));
    layer3_outputs(4988) <= '0';
    layer3_outputs(4989) <= layer2_outputs(2041);
    layer3_outputs(4990) <= (layer2_outputs(3606)) and not (layer2_outputs(5014));
    layer3_outputs(4991) <= not(layer2_outputs(2936)) or (layer2_outputs(1144));
    layer3_outputs(4992) <= not((layer2_outputs(839)) and (layer2_outputs(374)));
    layer3_outputs(4993) <= (layer2_outputs(1974)) or (layer2_outputs(1127));
    layer3_outputs(4994) <= '0';
    layer3_outputs(4995) <= '0';
    layer3_outputs(4996) <= not((layer2_outputs(2313)) and (layer2_outputs(2834)));
    layer3_outputs(4997) <= (layer2_outputs(2965)) and not (layer2_outputs(3991));
    layer3_outputs(4998) <= not(layer2_outputs(1165));
    layer3_outputs(4999) <= not(layer2_outputs(1835)) or (layer2_outputs(263));
    layer3_outputs(5000) <= not(layer2_outputs(1510)) or (layer2_outputs(5083));
    layer3_outputs(5001) <= '1';
    layer3_outputs(5002) <= not(layer2_outputs(5085)) or (layer2_outputs(4596));
    layer3_outputs(5003) <= not(layer2_outputs(384));
    layer3_outputs(5004) <= (layer2_outputs(4325)) and not (layer2_outputs(1421));
    layer3_outputs(5005) <= not(layer2_outputs(3293)) or (layer2_outputs(1437));
    layer3_outputs(5006) <= not(layer2_outputs(1046));
    layer3_outputs(5007) <= '1';
    layer3_outputs(5008) <= not(layer2_outputs(1250)) or (layer2_outputs(1434));
    layer3_outputs(5009) <= (layer2_outputs(3836)) and not (layer2_outputs(3304));
    layer3_outputs(5010) <= (layer2_outputs(1252)) and not (layer2_outputs(4148));
    layer3_outputs(5011) <= layer2_outputs(3088);
    layer3_outputs(5012) <= not(layer2_outputs(4130));
    layer3_outputs(5013) <= layer2_outputs(4105);
    layer3_outputs(5014) <= layer2_outputs(1136);
    layer3_outputs(5015) <= (layer2_outputs(5040)) and not (layer2_outputs(3833));
    layer3_outputs(5016) <= not((layer2_outputs(307)) and (layer2_outputs(1475)));
    layer3_outputs(5017) <= layer2_outputs(1695);
    layer3_outputs(5018) <= layer2_outputs(783);
    layer3_outputs(5019) <= not(layer2_outputs(3576)) or (layer2_outputs(1172));
    layer3_outputs(5020) <= '1';
    layer3_outputs(5021) <= (layer2_outputs(1312)) xor (layer2_outputs(4867));
    layer3_outputs(5022) <= not((layer2_outputs(2226)) or (layer2_outputs(3780)));
    layer3_outputs(5023) <= '1';
    layer3_outputs(5024) <= (layer2_outputs(4973)) or (layer2_outputs(4248));
    layer3_outputs(5025) <= layer2_outputs(675);
    layer3_outputs(5026) <= layer2_outputs(3675);
    layer3_outputs(5027) <= not(layer2_outputs(1764));
    layer3_outputs(5028) <= not(layer2_outputs(711));
    layer3_outputs(5029) <= (layer2_outputs(3752)) and not (layer2_outputs(199));
    layer3_outputs(5030) <= not(layer2_outputs(2020));
    layer3_outputs(5031) <= not(layer2_outputs(4266)) or (layer2_outputs(780));
    layer3_outputs(5032) <= not((layer2_outputs(1582)) xor (layer2_outputs(4010)));
    layer3_outputs(5033) <= (layer2_outputs(2617)) and not (layer2_outputs(3901));
    layer3_outputs(5034) <= not(layer2_outputs(5086));
    layer3_outputs(5035) <= not(layer2_outputs(4314)) or (layer2_outputs(2620));
    layer3_outputs(5036) <= '1';
    layer3_outputs(5037) <= '1';
    layer3_outputs(5038) <= layer2_outputs(1987);
    layer3_outputs(5039) <= not((layer2_outputs(2589)) and (layer2_outputs(1237)));
    layer3_outputs(5040) <= (layer2_outputs(1363)) and not (layer2_outputs(2291));
    layer3_outputs(5041) <= not((layer2_outputs(1105)) or (layer2_outputs(4840)));
    layer3_outputs(5042) <= '0';
    layer3_outputs(5043) <= not(layer2_outputs(2395));
    layer3_outputs(5044) <= (layer2_outputs(4843)) and not (layer2_outputs(4529));
    layer3_outputs(5045) <= (layer2_outputs(4761)) and not (layer2_outputs(1526));
    layer3_outputs(5046) <= layer2_outputs(924);
    layer3_outputs(5047) <= not(layer2_outputs(1196));
    layer3_outputs(5048) <= not(layer2_outputs(817));
    layer3_outputs(5049) <= not(layer2_outputs(2710));
    layer3_outputs(5050) <= (layer2_outputs(1528)) and not (layer2_outputs(636));
    layer3_outputs(5051) <= '1';
    layer3_outputs(5052) <= '1';
    layer3_outputs(5053) <= layer2_outputs(4489);
    layer3_outputs(5054) <= not(layer2_outputs(3678)) or (layer2_outputs(3479));
    layer3_outputs(5055) <= '1';
    layer3_outputs(5056) <= (layer2_outputs(1884)) and not (layer2_outputs(1245));
    layer3_outputs(5057) <= not(layer2_outputs(503)) or (layer2_outputs(2316));
    layer3_outputs(5058) <= not(layer2_outputs(4245));
    layer3_outputs(5059) <= '1';
    layer3_outputs(5060) <= (layer2_outputs(404)) and (layer2_outputs(1794));
    layer3_outputs(5061) <= layer2_outputs(2976);
    layer3_outputs(5062) <= not(layer2_outputs(3100));
    layer3_outputs(5063) <= '0';
    layer3_outputs(5064) <= '0';
    layer3_outputs(5065) <= not(layer2_outputs(4684)) or (layer2_outputs(4879));
    layer3_outputs(5066) <= (layer2_outputs(320)) and not (layer2_outputs(2861));
    layer3_outputs(5067) <= '0';
    layer3_outputs(5068) <= '0';
    layer3_outputs(5069) <= not((layer2_outputs(1523)) xor (layer2_outputs(4451)));
    layer3_outputs(5070) <= layer2_outputs(1583);
    layer3_outputs(5071) <= not((layer2_outputs(4280)) and (layer2_outputs(1797)));
    layer3_outputs(5072) <= layer2_outputs(3499);
    layer3_outputs(5073) <= not(layer2_outputs(3091)) or (layer2_outputs(4181));
    layer3_outputs(5074) <= layer2_outputs(278);
    layer3_outputs(5075) <= not(layer2_outputs(1226)) or (layer2_outputs(1750));
    layer3_outputs(5076) <= (layer2_outputs(1130)) and (layer2_outputs(4475));
    layer3_outputs(5077) <= not(layer2_outputs(697));
    layer3_outputs(5078) <= '1';
    layer3_outputs(5079) <= (layer2_outputs(4107)) and not (layer2_outputs(1463));
    layer3_outputs(5080) <= layer2_outputs(4045);
    layer3_outputs(5081) <= not(layer2_outputs(2079)) or (layer2_outputs(2632));
    layer3_outputs(5082) <= (layer2_outputs(1464)) and not (layer2_outputs(1761));
    layer3_outputs(5083) <= layer2_outputs(162);
    layer3_outputs(5084) <= not(layer2_outputs(2738)) or (layer2_outputs(4457));
    layer3_outputs(5085) <= (layer2_outputs(2930)) or (layer2_outputs(5106));
    layer3_outputs(5086) <= (layer2_outputs(1842)) xor (layer2_outputs(1440));
    layer3_outputs(5087) <= '1';
    layer3_outputs(5088) <= (layer2_outputs(2320)) and (layer2_outputs(3828));
    layer3_outputs(5089) <= '1';
    layer3_outputs(5090) <= not(layer2_outputs(813));
    layer3_outputs(5091) <= layer2_outputs(3377);
    layer3_outputs(5092) <= '1';
    layer3_outputs(5093) <= not(layer2_outputs(870)) or (layer2_outputs(4293));
    layer3_outputs(5094) <= layer2_outputs(1910);
    layer3_outputs(5095) <= (layer2_outputs(4202)) or (layer2_outputs(4094));
    layer3_outputs(5096) <= not(layer2_outputs(922)) or (layer2_outputs(1571));
    layer3_outputs(5097) <= '1';
    layer3_outputs(5098) <= layer2_outputs(1620);
    layer3_outputs(5099) <= not((layer2_outputs(2003)) and (layer2_outputs(4832)));
    layer3_outputs(5100) <= not(layer2_outputs(1007)) or (layer2_outputs(4218));
    layer3_outputs(5101) <= not(layer2_outputs(684));
    layer3_outputs(5102) <= (layer2_outputs(1370)) or (layer2_outputs(1147));
    layer3_outputs(5103) <= not(layer2_outputs(1025));
    layer3_outputs(5104) <= not((layer2_outputs(2298)) and (layer2_outputs(4131)));
    layer3_outputs(5105) <= '1';
    layer3_outputs(5106) <= layer2_outputs(4249);
    layer3_outputs(5107) <= not(layer2_outputs(963));
    layer3_outputs(5108) <= not(layer2_outputs(1584));
    layer3_outputs(5109) <= not(layer2_outputs(2873)) or (layer2_outputs(1603));
    layer3_outputs(5110) <= not(layer2_outputs(385));
    layer3_outputs(5111) <= (layer2_outputs(539)) and not (layer2_outputs(3161));
    layer3_outputs(5112) <= (layer2_outputs(4076)) and not (layer2_outputs(3933));
    layer3_outputs(5113) <= layer2_outputs(1294);
    layer3_outputs(5114) <= not(layer2_outputs(1485));
    layer3_outputs(5115) <= '0';
    layer3_outputs(5116) <= (layer2_outputs(3286)) and not (layer2_outputs(337));
    layer3_outputs(5117) <= layer2_outputs(1506);
    layer3_outputs(5118) <= not(layer2_outputs(1012));
    layer3_outputs(5119) <= '1';
    layer4_outputs(0) <= not(layer3_outputs(1488));
    layer4_outputs(1) <= (layer3_outputs(4369)) or (layer3_outputs(2901));
    layer4_outputs(2) <= layer3_outputs(2557);
    layer4_outputs(3) <= (layer3_outputs(2486)) and (layer3_outputs(5042));
    layer4_outputs(4) <= (layer3_outputs(3775)) or (layer3_outputs(621));
    layer4_outputs(5) <= (layer3_outputs(139)) and not (layer3_outputs(722));
    layer4_outputs(6) <= not(layer3_outputs(1837)) or (layer3_outputs(2015));
    layer4_outputs(7) <= not((layer3_outputs(301)) and (layer3_outputs(1153)));
    layer4_outputs(8) <= (layer3_outputs(3546)) and (layer3_outputs(326));
    layer4_outputs(9) <= (layer3_outputs(3465)) and not (layer3_outputs(340));
    layer4_outputs(10) <= not(layer3_outputs(967));
    layer4_outputs(11) <= not(layer3_outputs(4064));
    layer4_outputs(12) <= not(layer3_outputs(4366));
    layer4_outputs(13) <= '1';
    layer4_outputs(14) <= not((layer3_outputs(11)) and (layer3_outputs(403)));
    layer4_outputs(15) <= not(layer3_outputs(255));
    layer4_outputs(16) <= layer3_outputs(3482);
    layer4_outputs(17) <= layer3_outputs(958);
    layer4_outputs(18) <= not(layer3_outputs(4004));
    layer4_outputs(19) <= not(layer3_outputs(1217));
    layer4_outputs(20) <= layer3_outputs(3660);
    layer4_outputs(21) <= layer3_outputs(731);
    layer4_outputs(22) <= layer3_outputs(3284);
    layer4_outputs(23) <= not(layer3_outputs(2430)) or (layer3_outputs(2195));
    layer4_outputs(24) <= not(layer3_outputs(2924));
    layer4_outputs(25) <= (layer3_outputs(916)) and (layer3_outputs(855));
    layer4_outputs(26) <= not(layer3_outputs(2959));
    layer4_outputs(27) <= not(layer3_outputs(1713)) or (layer3_outputs(1081));
    layer4_outputs(28) <= layer3_outputs(1077);
    layer4_outputs(29) <= not(layer3_outputs(4123));
    layer4_outputs(30) <= not(layer3_outputs(1788)) or (layer3_outputs(3551));
    layer4_outputs(31) <= layer3_outputs(4250);
    layer4_outputs(32) <= not((layer3_outputs(4373)) xor (layer3_outputs(599)));
    layer4_outputs(33) <= '0';
    layer4_outputs(34) <= not(layer3_outputs(4840)) or (layer3_outputs(1736));
    layer4_outputs(35) <= (layer3_outputs(1554)) and not (layer3_outputs(4953));
    layer4_outputs(36) <= (layer3_outputs(913)) and (layer3_outputs(5088));
    layer4_outputs(37) <= '1';
    layer4_outputs(38) <= not(layer3_outputs(1854));
    layer4_outputs(39) <= (layer3_outputs(3439)) and not (layer3_outputs(4104));
    layer4_outputs(40) <= not((layer3_outputs(4209)) or (layer3_outputs(548)));
    layer4_outputs(41) <= not(layer3_outputs(5105));
    layer4_outputs(42) <= (layer3_outputs(2646)) xor (layer3_outputs(1380));
    layer4_outputs(43) <= not(layer3_outputs(642)) or (layer3_outputs(148));
    layer4_outputs(44) <= not((layer3_outputs(1794)) and (layer3_outputs(4903)));
    layer4_outputs(45) <= '0';
    layer4_outputs(46) <= not((layer3_outputs(1870)) or (layer3_outputs(216)));
    layer4_outputs(47) <= not(layer3_outputs(2228)) or (layer3_outputs(481));
    layer4_outputs(48) <= not(layer3_outputs(2836));
    layer4_outputs(49) <= not((layer3_outputs(4887)) xor (layer3_outputs(1442)));
    layer4_outputs(50) <= layer3_outputs(3136);
    layer4_outputs(51) <= layer3_outputs(2958);
    layer4_outputs(52) <= '0';
    layer4_outputs(53) <= '0';
    layer4_outputs(54) <= (layer3_outputs(3128)) xor (layer3_outputs(4602));
    layer4_outputs(55) <= (layer3_outputs(3984)) and not (layer3_outputs(934));
    layer4_outputs(56) <= not(layer3_outputs(2045));
    layer4_outputs(57) <= not(layer3_outputs(1032));
    layer4_outputs(58) <= layer3_outputs(208);
    layer4_outputs(59) <= not(layer3_outputs(555));
    layer4_outputs(60) <= not(layer3_outputs(3988));
    layer4_outputs(61) <= not(layer3_outputs(4819));
    layer4_outputs(62) <= (layer3_outputs(758)) and not (layer3_outputs(3043));
    layer4_outputs(63) <= layer3_outputs(66);
    layer4_outputs(64) <= layer3_outputs(3587);
    layer4_outputs(65) <= (layer3_outputs(1532)) or (layer3_outputs(415));
    layer4_outputs(66) <= not(layer3_outputs(4915));
    layer4_outputs(67) <= not(layer3_outputs(4528)) or (layer3_outputs(3481));
    layer4_outputs(68) <= (layer3_outputs(1521)) and (layer3_outputs(5060));
    layer4_outputs(69) <= not(layer3_outputs(2992));
    layer4_outputs(70) <= (layer3_outputs(4297)) and (layer3_outputs(4833));
    layer4_outputs(71) <= not(layer3_outputs(3393)) or (layer3_outputs(2447));
    layer4_outputs(72) <= not(layer3_outputs(2610)) or (layer3_outputs(3325));
    layer4_outputs(73) <= '1';
    layer4_outputs(74) <= '1';
    layer4_outputs(75) <= not((layer3_outputs(1319)) or (layer3_outputs(3330)));
    layer4_outputs(76) <= (layer3_outputs(1190)) and not (layer3_outputs(2727));
    layer4_outputs(77) <= layer3_outputs(4308);
    layer4_outputs(78) <= '1';
    layer4_outputs(79) <= not(layer3_outputs(2508)) or (layer3_outputs(3237));
    layer4_outputs(80) <= layer3_outputs(3350);
    layer4_outputs(81) <= (layer3_outputs(2951)) and (layer3_outputs(4323));
    layer4_outputs(82) <= not(layer3_outputs(3580));
    layer4_outputs(83) <= layer3_outputs(3628);
    layer4_outputs(84) <= (layer3_outputs(705)) and not (layer3_outputs(2757));
    layer4_outputs(85) <= layer3_outputs(91);
    layer4_outputs(86) <= (layer3_outputs(4989)) and not (layer3_outputs(1475));
    layer4_outputs(87) <= not((layer3_outputs(1451)) or (layer3_outputs(3555)));
    layer4_outputs(88) <= not(layer3_outputs(1574));
    layer4_outputs(89) <= '1';
    layer4_outputs(90) <= not((layer3_outputs(4341)) xor (layer3_outputs(3511)));
    layer4_outputs(91) <= not((layer3_outputs(2569)) and (layer3_outputs(404)));
    layer4_outputs(92) <= not(layer3_outputs(4087)) or (layer3_outputs(4825));
    layer4_outputs(93) <= layer3_outputs(1281);
    layer4_outputs(94) <= layer3_outputs(937);
    layer4_outputs(95) <= '1';
    layer4_outputs(96) <= not(layer3_outputs(603));
    layer4_outputs(97) <= layer3_outputs(3646);
    layer4_outputs(98) <= not(layer3_outputs(4911)) or (layer3_outputs(834));
    layer4_outputs(99) <= layer3_outputs(2728);
    layer4_outputs(100) <= not(layer3_outputs(5059));
    layer4_outputs(101) <= (layer3_outputs(3149)) or (layer3_outputs(4728));
    layer4_outputs(102) <= not(layer3_outputs(4878));
    layer4_outputs(103) <= layer3_outputs(388);
    layer4_outputs(104) <= not((layer3_outputs(2952)) and (layer3_outputs(1146)));
    layer4_outputs(105) <= not(layer3_outputs(2600));
    layer4_outputs(106) <= not(layer3_outputs(156)) or (layer3_outputs(2944));
    layer4_outputs(107) <= (layer3_outputs(4236)) and not (layer3_outputs(67));
    layer4_outputs(108) <= not(layer3_outputs(1865)) or (layer3_outputs(1246));
    layer4_outputs(109) <= layer3_outputs(127);
    layer4_outputs(110) <= (layer3_outputs(2101)) and not (layer3_outputs(4774));
    layer4_outputs(111) <= layer3_outputs(4509);
    layer4_outputs(112) <= not((layer3_outputs(61)) or (layer3_outputs(3434)));
    layer4_outputs(113) <= not((layer3_outputs(1053)) and (layer3_outputs(4346)));
    layer4_outputs(114) <= layer3_outputs(2637);
    layer4_outputs(115) <= not((layer3_outputs(1153)) or (layer3_outputs(3698)));
    layer4_outputs(116) <= (layer3_outputs(857)) or (layer3_outputs(150));
    layer4_outputs(117) <= not((layer3_outputs(4327)) xor (layer3_outputs(654)));
    layer4_outputs(118) <= not(layer3_outputs(4662));
    layer4_outputs(119) <= not(layer3_outputs(643));
    layer4_outputs(120) <= not(layer3_outputs(128));
    layer4_outputs(121) <= not((layer3_outputs(3429)) and (layer3_outputs(4415)));
    layer4_outputs(122) <= '0';
    layer4_outputs(123) <= not(layer3_outputs(2716));
    layer4_outputs(124) <= not((layer3_outputs(1564)) and (layer3_outputs(459)));
    layer4_outputs(125) <= not((layer3_outputs(4627)) and (layer3_outputs(1630)));
    layer4_outputs(126) <= layer3_outputs(4592);
    layer4_outputs(127) <= layer3_outputs(1055);
    layer4_outputs(128) <= (layer3_outputs(4705)) and not (layer3_outputs(808));
    layer4_outputs(129) <= (layer3_outputs(4814)) xor (layer3_outputs(913));
    layer4_outputs(130) <= (layer3_outputs(1494)) or (layer3_outputs(2412));
    layer4_outputs(131) <= not(layer3_outputs(73)) or (layer3_outputs(2782));
    layer4_outputs(132) <= not((layer3_outputs(2580)) or (layer3_outputs(2910)));
    layer4_outputs(133) <= not((layer3_outputs(678)) and (layer3_outputs(2141)));
    layer4_outputs(134) <= layer3_outputs(3503);
    layer4_outputs(135) <= not((layer3_outputs(3447)) and (layer3_outputs(110)));
    layer4_outputs(136) <= layer3_outputs(122);
    layer4_outputs(137) <= '0';
    layer4_outputs(138) <= '0';
    layer4_outputs(139) <= not(layer3_outputs(3402));
    layer4_outputs(140) <= (layer3_outputs(158)) and not (layer3_outputs(4675));
    layer4_outputs(141) <= layer3_outputs(96);
    layer4_outputs(142) <= not((layer3_outputs(4813)) and (layer3_outputs(3587)));
    layer4_outputs(143) <= layer3_outputs(4203);
    layer4_outputs(144) <= layer3_outputs(2792);
    layer4_outputs(145) <= not((layer3_outputs(4063)) and (layer3_outputs(116)));
    layer4_outputs(146) <= not(layer3_outputs(3949)) or (layer3_outputs(4798));
    layer4_outputs(147) <= layer3_outputs(5022);
    layer4_outputs(148) <= (layer3_outputs(1738)) and not (layer3_outputs(4559));
    layer4_outputs(149) <= (layer3_outputs(3452)) and (layer3_outputs(2685));
    layer4_outputs(150) <= (layer3_outputs(344)) and not (layer3_outputs(3376));
    layer4_outputs(151) <= '1';
    layer4_outputs(152) <= '0';
    layer4_outputs(153) <= not((layer3_outputs(3063)) and (layer3_outputs(3367)));
    layer4_outputs(154) <= layer3_outputs(3924);
    layer4_outputs(155) <= '0';
    layer4_outputs(156) <= (layer3_outputs(4854)) and not (layer3_outputs(3550));
    layer4_outputs(157) <= '1';
    layer4_outputs(158) <= layer3_outputs(4025);
    layer4_outputs(159) <= not(layer3_outputs(2146));
    layer4_outputs(160) <= '0';
    layer4_outputs(161) <= not((layer3_outputs(408)) xor (layer3_outputs(226)));
    layer4_outputs(162) <= (layer3_outputs(2879)) and not (layer3_outputs(2654));
    layer4_outputs(163) <= (layer3_outputs(4379)) or (layer3_outputs(3408));
    layer4_outputs(164) <= layer3_outputs(4875);
    layer4_outputs(165) <= not(layer3_outputs(4599));
    layer4_outputs(166) <= not((layer3_outputs(1326)) and (layer3_outputs(2592)));
    layer4_outputs(167) <= layer3_outputs(2382);
    layer4_outputs(168) <= not(layer3_outputs(666));
    layer4_outputs(169) <= layer3_outputs(2);
    layer4_outputs(170) <= not(layer3_outputs(777));
    layer4_outputs(171) <= '0';
    layer4_outputs(172) <= (layer3_outputs(3213)) and not (layer3_outputs(2961));
    layer4_outputs(173) <= layer3_outputs(3444);
    layer4_outputs(174) <= not(layer3_outputs(28));
    layer4_outputs(175) <= (layer3_outputs(4309)) and not (layer3_outputs(2904));
    layer4_outputs(176) <= layer3_outputs(3674);
    layer4_outputs(177) <= layer3_outputs(1239);
    layer4_outputs(178) <= not(layer3_outputs(4282)) or (layer3_outputs(703));
    layer4_outputs(179) <= not((layer3_outputs(2255)) xor (layer3_outputs(1625)));
    layer4_outputs(180) <= not((layer3_outputs(112)) and (layer3_outputs(279)));
    layer4_outputs(181) <= layer3_outputs(3732);
    layer4_outputs(182) <= layer3_outputs(763);
    layer4_outputs(183) <= (layer3_outputs(1324)) and (layer3_outputs(834));
    layer4_outputs(184) <= not((layer3_outputs(1662)) and (layer3_outputs(2636)));
    layer4_outputs(185) <= layer3_outputs(2438);
    layer4_outputs(186) <= not((layer3_outputs(4310)) or (layer3_outputs(953)));
    layer4_outputs(187) <= not(layer3_outputs(2629));
    layer4_outputs(188) <= not(layer3_outputs(791));
    layer4_outputs(189) <= layer3_outputs(2568);
    layer4_outputs(190) <= (layer3_outputs(2967)) or (layer3_outputs(963));
    layer4_outputs(191) <= not(layer3_outputs(380));
    layer4_outputs(192) <= layer3_outputs(1943);
    layer4_outputs(193) <= '1';
    layer4_outputs(194) <= (layer3_outputs(266)) and not (layer3_outputs(1681));
    layer4_outputs(195) <= (layer3_outputs(3044)) and not (layer3_outputs(2776));
    layer4_outputs(196) <= (layer3_outputs(1942)) and not (layer3_outputs(465));
    layer4_outputs(197) <= '1';
    layer4_outputs(198) <= not(layer3_outputs(3610));
    layer4_outputs(199) <= not(layer3_outputs(2343));
    layer4_outputs(200) <= '0';
    layer4_outputs(201) <= (layer3_outputs(2701)) or (layer3_outputs(1661));
    layer4_outputs(202) <= '1';
    layer4_outputs(203) <= layer3_outputs(2799);
    layer4_outputs(204) <= not(layer3_outputs(3814));
    layer4_outputs(205) <= not((layer3_outputs(3161)) or (layer3_outputs(1121)));
    layer4_outputs(206) <= not(layer3_outputs(2399));
    layer4_outputs(207) <= not(layer3_outputs(2378));
    layer4_outputs(208) <= not(layer3_outputs(1871)) or (layer3_outputs(4029));
    layer4_outputs(209) <= (layer3_outputs(203)) and not (layer3_outputs(94));
    layer4_outputs(210) <= (layer3_outputs(5012)) xor (layer3_outputs(1895));
    layer4_outputs(211) <= not(layer3_outputs(1619)) or (layer3_outputs(2886));
    layer4_outputs(212) <= not(layer3_outputs(3519)) or (layer3_outputs(1382));
    layer4_outputs(213) <= layer3_outputs(3442);
    layer4_outputs(214) <= (layer3_outputs(3542)) and (layer3_outputs(3415));
    layer4_outputs(215) <= not(layer3_outputs(1857));
    layer4_outputs(216) <= (layer3_outputs(4574)) xor (layer3_outputs(3476));
    layer4_outputs(217) <= '1';
    layer4_outputs(218) <= layer3_outputs(3827);
    layer4_outputs(219) <= (layer3_outputs(556)) or (layer3_outputs(1440));
    layer4_outputs(220) <= not((layer3_outputs(1953)) xor (layer3_outputs(207)));
    layer4_outputs(221) <= not(layer3_outputs(1448));
    layer4_outputs(222) <= not((layer3_outputs(1068)) or (layer3_outputs(2059)));
    layer4_outputs(223) <= '1';
    layer4_outputs(224) <= not(layer3_outputs(4633));
    layer4_outputs(225) <= '0';
    layer4_outputs(226) <= (layer3_outputs(3839)) and not (layer3_outputs(1051));
    layer4_outputs(227) <= not((layer3_outputs(3020)) and (layer3_outputs(4606)));
    layer4_outputs(228) <= not(layer3_outputs(3734));
    layer4_outputs(229) <= not(layer3_outputs(3044));
    layer4_outputs(230) <= (layer3_outputs(4001)) and not (layer3_outputs(3466));
    layer4_outputs(231) <= layer3_outputs(648);
    layer4_outputs(232) <= layer3_outputs(1028);
    layer4_outputs(233) <= not(layer3_outputs(3042)) or (layer3_outputs(3567));
    layer4_outputs(234) <= not(layer3_outputs(3931)) or (layer3_outputs(4017));
    layer4_outputs(235) <= not(layer3_outputs(3112));
    layer4_outputs(236) <= '1';
    layer4_outputs(237) <= not((layer3_outputs(2254)) and (layer3_outputs(3299)));
    layer4_outputs(238) <= not((layer3_outputs(2097)) and (layer3_outputs(1103)));
    layer4_outputs(239) <= (layer3_outputs(1666)) and not (layer3_outputs(3199));
    layer4_outputs(240) <= not(layer3_outputs(1524));
    layer4_outputs(241) <= (layer3_outputs(1589)) or (layer3_outputs(4331));
    layer4_outputs(242) <= not((layer3_outputs(4015)) and (layer3_outputs(3258)));
    layer4_outputs(243) <= not((layer3_outputs(1702)) or (layer3_outputs(872)));
    layer4_outputs(244) <= (layer3_outputs(1148)) and not (layer3_outputs(1990));
    layer4_outputs(245) <= (layer3_outputs(925)) and not (layer3_outputs(33));
    layer4_outputs(246) <= (layer3_outputs(253)) and not (layer3_outputs(322));
    layer4_outputs(247) <= not(layer3_outputs(3197));
    layer4_outputs(248) <= not(layer3_outputs(1156));
    layer4_outputs(249) <= layer3_outputs(1925);
    layer4_outputs(250) <= not((layer3_outputs(2992)) and (layer3_outputs(2288)));
    layer4_outputs(251) <= layer3_outputs(3167);
    layer4_outputs(252) <= layer3_outputs(2168);
    layer4_outputs(253) <= layer3_outputs(5032);
    layer4_outputs(254) <= (layer3_outputs(1377)) and (layer3_outputs(3984));
    layer4_outputs(255) <= not(layer3_outputs(3757));
    layer4_outputs(256) <= (layer3_outputs(4836)) and (layer3_outputs(4886));
    layer4_outputs(257) <= not(layer3_outputs(1149)) or (layer3_outputs(1742));
    layer4_outputs(258) <= not(layer3_outputs(1206)) or (layer3_outputs(4163));
    layer4_outputs(259) <= layer3_outputs(2196);
    layer4_outputs(260) <= not(layer3_outputs(1732));
    layer4_outputs(261) <= (layer3_outputs(3550)) and not (layer3_outputs(4582));
    layer4_outputs(262) <= (layer3_outputs(1279)) and (layer3_outputs(3045));
    layer4_outputs(263) <= layer3_outputs(2463);
    layer4_outputs(264) <= not(layer3_outputs(2142));
    layer4_outputs(265) <= layer3_outputs(2200);
    layer4_outputs(266) <= '1';
    layer4_outputs(267) <= (layer3_outputs(232)) xor (layer3_outputs(4548));
    layer4_outputs(268) <= not(layer3_outputs(1486));
    layer4_outputs(269) <= not((layer3_outputs(3986)) or (layer3_outputs(4893)));
    layer4_outputs(270) <= not((layer3_outputs(2196)) or (layer3_outputs(1185)));
    layer4_outputs(271) <= not(layer3_outputs(499)) or (layer3_outputs(4647));
    layer4_outputs(272) <= '1';
    layer4_outputs(273) <= '1';
    layer4_outputs(274) <= layer3_outputs(790);
    layer4_outputs(275) <= layer3_outputs(3684);
    layer4_outputs(276) <= not((layer3_outputs(3515)) xor (layer3_outputs(1574)));
    layer4_outputs(277) <= (layer3_outputs(3355)) and (layer3_outputs(356));
    layer4_outputs(278) <= (layer3_outputs(4053)) and not (layer3_outputs(1671));
    layer4_outputs(279) <= layer3_outputs(947);
    layer4_outputs(280) <= not(layer3_outputs(4665)) or (layer3_outputs(4189));
    layer4_outputs(281) <= not(layer3_outputs(707));
    layer4_outputs(282) <= layer3_outputs(4969);
    layer4_outputs(283) <= (layer3_outputs(2878)) xor (layer3_outputs(3167));
    layer4_outputs(284) <= (layer3_outputs(1786)) and not (layer3_outputs(2781));
    layer4_outputs(285) <= (layer3_outputs(2367)) and (layer3_outputs(3234));
    layer4_outputs(286) <= not(layer3_outputs(4448));
    layer4_outputs(287) <= not(layer3_outputs(4505));
    layer4_outputs(288) <= layer3_outputs(3646);
    layer4_outputs(289) <= not(layer3_outputs(2785)) or (layer3_outputs(46));
    layer4_outputs(290) <= not(layer3_outputs(1245));
    layer4_outputs(291) <= not((layer3_outputs(4734)) or (layer3_outputs(4770)));
    layer4_outputs(292) <= layer3_outputs(2059);
    layer4_outputs(293) <= '0';
    layer4_outputs(294) <= (layer3_outputs(915)) xor (layer3_outputs(770));
    layer4_outputs(295) <= not((layer3_outputs(1706)) or (layer3_outputs(1721)));
    layer4_outputs(296) <= not((layer3_outputs(823)) and (layer3_outputs(333)));
    layer4_outputs(297) <= layer3_outputs(500);
    layer4_outputs(298) <= not(layer3_outputs(1487)) or (layer3_outputs(1021));
    layer4_outputs(299) <= layer3_outputs(3860);
    layer4_outputs(300) <= layer3_outputs(1145);
    layer4_outputs(301) <= not(layer3_outputs(2838)) or (layer3_outputs(1416));
    layer4_outputs(302) <= not((layer3_outputs(2620)) and (layer3_outputs(218)));
    layer4_outputs(303) <= layer3_outputs(1111);
    layer4_outputs(304) <= (layer3_outputs(1513)) and not (layer3_outputs(3007));
    layer4_outputs(305) <= not(layer3_outputs(1534)) or (layer3_outputs(3354));
    layer4_outputs(306) <= not(layer3_outputs(2235)) or (layer3_outputs(3951));
    layer4_outputs(307) <= '0';
    layer4_outputs(308) <= (layer3_outputs(893)) xor (layer3_outputs(2317));
    layer4_outputs(309) <= (layer3_outputs(786)) or (layer3_outputs(3709));
    layer4_outputs(310) <= not((layer3_outputs(577)) or (layer3_outputs(217)));
    layer4_outputs(311) <= not(layer3_outputs(1363)) or (layer3_outputs(1067));
    layer4_outputs(312) <= not(layer3_outputs(573));
    layer4_outputs(313) <= '0';
    layer4_outputs(314) <= layer3_outputs(3445);
    layer4_outputs(315) <= not(layer3_outputs(933));
    layer4_outputs(316) <= not(layer3_outputs(4949));
    layer4_outputs(317) <= not(layer3_outputs(4262));
    layer4_outputs(318) <= not(layer3_outputs(1542));
    layer4_outputs(319) <= layer3_outputs(4201);
    layer4_outputs(320) <= not((layer3_outputs(1078)) or (layer3_outputs(3391)));
    layer4_outputs(321) <= not(layer3_outputs(3137)) or (layer3_outputs(1370));
    layer4_outputs(322) <= not(layer3_outputs(1543));
    layer4_outputs(323) <= layer3_outputs(93);
    layer4_outputs(324) <= (layer3_outputs(1538)) and (layer3_outputs(3799));
    layer4_outputs(325) <= (layer3_outputs(2274)) and (layer3_outputs(2091));
    layer4_outputs(326) <= (layer3_outputs(1)) or (layer3_outputs(3647));
    layer4_outputs(327) <= layer3_outputs(1806);
    layer4_outputs(328) <= (layer3_outputs(4952)) and (layer3_outputs(3108));
    layer4_outputs(329) <= (layer3_outputs(1323)) or (layer3_outputs(977));
    layer4_outputs(330) <= (layer3_outputs(2103)) or (layer3_outputs(4597));
    layer4_outputs(331) <= not(layer3_outputs(4586));
    layer4_outputs(332) <= not((layer3_outputs(2684)) and (layer3_outputs(4527)));
    layer4_outputs(333) <= '1';
    layer4_outputs(334) <= (layer3_outputs(3990)) or (layer3_outputs(4009));
    layer4_outputs(335) <= layer3_outputs(2178);
    layer4_outputs(336) <= layer3_outputs(2275);
    layer4_outputs(337) <= not(layer3_outputs(1136));
    layer4_outputs(338) <= not(layer3_outputs(2210)) or (layer3_outputs(3919));
    layer4_outputs(339) <= not(layer3_outputs(2069)) or (layer3_outputs(2357));
    layer4_outputs(340) <= (layer3_outputs(1128)) and not (layer3_outputs(4074));
    layer4_outputs(341) <= layer3_outputs(1711);
    layer4_outputs(342) <= (layer3_outputs(4073)) and (layer3_outputs(1219));
    layer4_outputs(343) <= not(layer3_outputs(2375));
    layer4_outputs(344) <= not((layer3_outputs(1423)) and (layer3_outputs(4233)));
    layer4_outputs(345) <= not(layer3_outputs(4553));
    layer4_outputs(346) <= not(layer3_outputs(2544)) or (layer3_outputs(1548));
    layer4_outputs(347) <= layer3_outputs(529);
    layer4_outputs(348) <= not(layer3_outputs(3308));
    layer4_outputs(349) <= layer3_outputs(3793);
    layer4_outputs(350) <= (layer3_outputs(1181)) or (layer3_outputs(3697));
    layer4_outputs(351) <= not(layer3_outputs(1725));
    layer4_outputs(352) <= not((layer3_outputs(1739)) and (layer3_outputs(1916)));
    layer4_outputs(353) <= not(layer3_outputs(2707));
    layer4_outputs(354) <= not(layer3_outputs(766)) or (layer3_outputs(812));
    layer4_outputs(355) <= not(layer3_outputs(1074)) or (layer3_outputs(3243));
    layer4_outputs(356) <= (layer3_outputs(819)) and not (layer3_outputs(3557));
    layer4_outputs(357) <= not(layer3_outputs(1440));
    layer4_outputs(358) <= (layer3_outputs(1400)) and (layer3_outputs(4845));
    layer4_outputs(359) <= not(layer3_outputs(2726)) or (layer3_outputs(1890));
    layer4_outputs(360) <= (layer3_outputs(2323)) and not (layer3_outputs(2118));
    layer4_outputs(361) <= '0';
    layer4_outputs(362) <= (layer3_outputs(2857)) and not (layer3_outputs(4103));
    layer4_outputs(363) <= not((layer3_outputs(2623)) and (layer3_outputs(1383)));
    layer4_outputs(364) <= not(layer3_outputs(3929));
    layer4_outputs(365) <= (layer3_outputs(2408)) and (layer3_outputs(451));
    layer4_outputs(366) <= not(layer3_outputs(563));
    layer4_outputs(367) <= layer3_outputs(1089);
    layer4_outputs(368) <= not(layer3_outputs(18));
    layer4_outputs(369) <= not(layer3_outputs(153));
    layer4_outputs(370) <= layer3_outputs(4105);
    layer4_outputs(371) <= layer3_outputs(5019);
    layer4_outputs(372) <= layer3_outputs(2367);
    layer4_outputs(373) <= layer3_outputs(2063);
    layer4_outputs(374) <= (layer3_outputs(1997)) or (layer3_outputs(2094));
    layer4_outputs(375) <= layer3_outputs(2012);
    layer4_outputs(376) <= (layer3_outputs(1231)) or (layer3_outputs(3372));
    layer4_outputs(377) <= not(layer3_outputs(0));
    layer4_outputs(378) <= (layer3_outputs(3767)) and not (layer3_outputs(996));
    layer4_outputs(379) <= (layer3_outputs(910)) or (layer3_outputs(402));
    layer4_outputs(380) <= layer3_outputs(2970);
    layer4_outputs(381) <= (layer3_outputs(1582)) and not (layer3_outputs(23));
    layer4_outputs(382) <= not((layer3_outputs(3729)) and (layer3_outputs(3287)));
    layer4_outputs(383) <= layer3_outputs(2345);
    layer4_outputs(384) <= layer3_outputs(1648);
    layer4_outputs(385) <= (layer3_outputs(1471)) or (layer3_outputs(4626));
    layer4_outputs(386) <= not(layer3_outputs(3488));
    layer4_outputs(387) <= (layer3_outputs(3203)) or (layer3_outputs(2976));
    layer4_outputs(388) <= not((layer3_outputs(2723)) xor (layer3_outputs(4682)));
    layer4_outputs(389) <= layer3_outputs(346);
    layer4_outputs(390) <= not((layer3_outputs(2527)) or (layer3_outputs(3521)));
    layer4_outputs(391) <= layer3_outputs(4076);
    layer4_outputs(392) <= not(layer3_outputs(5078));
    layer4_outputs(393) <= layer3_outputs(1614);
    layer4_outputs(394) <= not(layer3_outputs(2816)) or (layer3_outputs(1194));
    layer4_outputs(395) <= layer3_outputs(4751);
    layer4_outputs(396) <= layer3_outputs(224);
    layer4_outputs(397) <= (layer3_outputs(2842)) and (layer3_outputs(1381));
    layer4_outputs(398) <= (layer3_outputs(172)) or (layer3_outputs(3021));
    layer4_outputs(399) <= not((layer3_outputs(2447)) or (layer3_outputs(4807)));
    layer4_outputs(400) <= not((layer3_outputs(891)) xor (layer3_outputs(611)));
    layer4_outputs(401) <= not((layer3_outputs(2702)) or (layer3_outputs(2556)));
    layer4_outputs(402) <= not(layer3_outputs(437));
    layer4_outputs(403) <= not((layer3_outputs(5069)) or (layer3_outputs(4864)));
    layer4_outputs(404) <= layer3_outputs(781);
    layer4_outputs(405) <= '0';
    layer4_outputs(406) <= (layer3_outputs(4685)) and (layer3_outputs(1392));
    layer4_outputs(407) <= not(layer3_outputs(1724));
    layer4_outputs(408) <= '0';
    layer4_outputs(409) <= '0';
    layer4_outputs(410) <= not(layer3_outputs(1531)) or (layer3_outputs(550));
    layer4_outputs(411) <= '1';
    layer4_outputs(412) <= not((layer3_outputs(17)) or (layer3_outputs(975)));
    layer4_outputs(413) <= not((layer3_outputs(102)) or (layer3_outputs(1608)));
    layer4_outputs(414) <= '0';
    layer4_outputs(415) <= layer3_outputs(1187);
    layer4_outputs(416) <= '1';
    layer4_outputs(417) <= layer3_outputs(596);
    layer4_outputs(418) <= not((layer3_outputs(175)) and (layer3_outputs(848)));
    layer4_outputs(419) <= layer3_outputs(1147);
    layer4_outputs(420) <= not(layer3_outputs(4148));
    layer4_outputs(421) <= not(layer3_outputs(2322));
    layer4_outputs(422) <= not(layer3_outputs(4080));
    layer4_outputs(423) <= not(layer3_outputs(2378));
    layer4_outputs(424) <= layer3_outputs(2156);
    layer4_outputs(425) <= (layer3_outputs(2480)) or (layer3_outputs(163));
    layer4_outputs(426) <= not(layer3_outputs(3657));
    layer4_outputs(427) <= layer3_outputs(1886);
    layer4_outputs(428) <= layer3_outputs(48);
    layer4_outputs(429) <= not(layer3_outputs(4701));
    layer4_outputs(430) <= not((layer3_outputs(2)) and (layer3_outputs(4110)));
    layer4_outputs(431) <= not((layer3_outputs(1052)) xor (layer3_outputs(2768)));
    layer4_outputs(432) <= (layer3_outputs(2829)) or (layer3_outputs(1803));
    layer4_outputs(433) <= not(layer3_outputs(484)) or (layer3_outputs(3757));
    layer4_outputs(434) <= (layer3_outputs(3001)) and not (layer3_outputs(4795));
    layer4_outputs(435) <= not((layer3_outputs(2617)) xor (layer3_outputs(2295)));
    layer4_outputs(436) <= not((layer3_outputs(578)) or (layer3_outputs(4591)));
    layer4_outputs(437) <= not(layer3_outputs(2851));
    layer4_outputs(438) <= not(layer3_outputs(2327));
    layer4_outputs(439) <= layer3_outputs(1123);
    layer4_outputs(440) <= layer3_outputs(3851);
    layer4_outputs(441) <= layer3_outputs(4497);
    layer4_outputs(442) <= (layer3_outputs(2273)) and (layer3_outputs(158));
    layer4_outputs(443) <= not(layer3_outputs(3505));
    layer4_outputs(444) <= layer3_outputs(1214);
    layer4_outputs(445) <= layer3_outputs(1111);
    layer4_outputs(446) <= not(layer3_outputs(3593)) or (layer3_outputs(568));
    layer4_outputs(447) <= layer3_outputs(4476);
    layer4_outputs(448) <= (layer3_outputs(3215)) and not (layer3_outputs(4086));
    layer4_outputs(449) <= (layer3_outputs(3528)) xor (layer3_outputs(2848));
    layer4_outputs(450) <= (layer3_outputs(5047)) and not (layer3_outputs(3111));
    layer4_outputs(451) <= not((layer3_outputs(2913)) and (layer3_outputs(4971)));
    layer4_outputs(452) <= not(layer3_outputs(3788));
    layer4_outputs(453) <= '1';
    layer4_outputs(454) <= (layer3_outputs(3469)) and not (layer3_outputs(352));
    layer4_outputs(455) <= layer3_outputs(2095);
    layer4_outputs(456) <= not(layer3_outputs(5082)) or (layer3_outputs(2274));
    layer4_outputs(457) <= not(layer3_outputs(2212));
    layer4_outputs(458) <= not(layer3_outputs(3359));
    layer4_outputs(459) <= '1';
    layer4_outputs(460) <= not(layer3_outputs(3906)) or (layer3_outputs(4447));
    layer4_outputs(461) <= not((layer3_outputs(1516)) or (layer3_outputs(2751)));
    layer4_outputs(462) <= not(layer3_outputs(2894));
    layer4_outputs(463) <= not(layer3_outputs(1755));
    layer4_outputs(464) <= not(layer3_outputs(4846));
    layer4_outputs(465) <= not(layer3_outputs(424));
    layer4_outputs(466) <= not(layer3_outputs(1867)) or (layer3_outputs(3538));
    layer4_outputs(467) <= (layer3_outputs(4679)) and (layer3_outputs(1700));
    layer4_outputs(468) <= (layer3_outputs(2404)) xor (layer3_outputs(1749));
    layer4_outputs(469) <= '0';
    layer4_outputs(470) <= not(layer3_outputs(3026));
    layer4_outputs(471) <= layer3_outputs(1638);
    layer4_outputs(472) <= not((layer3_outputs(167)) and (layer3_outputs(3274)));
    layer4_outputs(473) <= not(layer3_outputs(4577)) or (layer3_outputs(2127));
    layer4_outputs(474) <= not(layer3_outputs(728)) or (layer3_outputs(1962));
    layer4_outputs(475) <= '0';
    layer4_outputs(476) <= (layer3_outputs(2603)) or (layer3_outputs(4593));
    layer4_outputs(477) <= not((layer3_outputs(759)) and (layer3_outputs(299)));
    layer4_outputs(478) <= (layer3_outputs(1985)) and not (layer3_outputs(513));
    layer4_outputs(479) <= layer3_outputs(2545);
    layer4_outputs(480) <= not(layer3_outputs(3680));
    layer4_outputs(481) <= (layer3_outputs(3210)) and not (layer3_outputs(4068));
    layer4_outputs(482) <= not(layer3_outputs(3934)) or (layer3_outputs(540));
    layer4_outputs(483) <= (layer3_outputs(2874)) or (layer3_outputs(1744));
    layer4_outputs(484) <= not(layer3_outputs(3605)) or (layer3_outputs(3303));
    layer4_outputs(485) <= layer3_outputs(3761);
    layer4_outputs(486) <= (layer3_outputs(3072)) and not (layer3_outputs(1555));
    layer4_outputs(487) <= not((layer3_outputs(4125)) xor (layer3_outputs(2622)));
    layer4_outputs(488) <= not(layer3_outputs(241)) or (layer3_outputs(2622));
    layer4_outputs(489) <= not(layer3_outputs(2947));
    layer4_outputs(490) <= (layer3_outputs(3512)) and not (layer3_outputs(4490));
    layer4_outputs(491) <= not((layer3_outputs(3237)) and (layer3_outputs(5083)));
    layer4_outputs(492) <= layer3_outputs(4038);
    layer4_outputs(493) <= not((layer3_outputs(1232)) or (layer3_outputs(2232)));
    layer4_outputs(494) <= (layer3_outputs(1604)) and (layer3_outputs(4231));
    layer4_outputs(495) <= '1';
    layer4_outputs(496) <= layer3_outputs(1412);
    layer4_outputs(497) <= layer3_outputs(4468);
    layer4_outputs(498) <= (layer3_outputs(3409)) and not (layer3_outputs(4180));
    layer4_outputs(499) <= layer3_outputs(2298);
    layer4_outputs(500) <= '1';
    layer4_outputs(501) <= (layer3_outputs(2619)) or (layer3_outputs(3362));
    layer4_outputs(502) <= (layer3_outputs(261)) or (layer3_outputs(3003));
    layer4_outputs(503) <= (layer3_outputs(2638)) xor (layer3_outputs(4872));
    layer4_outputs(504) <= layer3_outputs(3891);
    layer4_outputs(505) <= not((layer3_outputs(3681)) xor (layer3_outputs(4191)));
    layer4_outputs(506) <= '0';
    layer4_outputs(507) <= not((layer3_outputs(39)) or (layer3_outputs(2869)));
    layer4_outputs(508) <= (layer3_outputs(1042)) and not (layer3_outputs(2838));
    layer4_outputs(509) <= '0';
    layer4_outputs(510) <= not(layer3_outputs(3983));
    layer4_outputs(511) <= layer3_outputs(3883);
    layer4_outputs(512) <= layer3_outputs(3821);
    layer4_outputs(513) <= not(layer3_outputs(453));
    layer4_outputs(514) <= not((layer3_outputs(3751)) or (layer3_outputs(3738)));
    layer4_outputs(515) <= not(layer3_outputs(1790)) or (layer3_outputs(3609));
    layer4_outputs(516) <= (layer3_outputs(2066)) or (layer3_outputs(1026));
    layer4_outputs(517) <= not(layer3_outputs(1578)) or (layer3_outputs(745));
    layer4_outputs(518) <= layer3_outputs(5107);
    layer4_outputs(519) <= (layer3_outputs(1003)) and not (layer3_outputs(3429));
    layer4_outputs(520) <= '1';
    layer4_outputs(521) <= layer3_outputs(3064);
    layer4_outputs(522) <= not(layer3_outputs(3602));
    layer4_outputs(523) <= layer3_outputs(121);
    layer4_outputs(524) <= layer3_outputs(4757);
    layer4_outputs(525) <= not(layer3_outputs(1641));
    layer4_outputs(526) <= not(layer3_outputs(2381));
    layer4_outputs(527) <= layer3_outputs(4698);
    layer4_outputs(528) <= (layer3_outputs(3080)) xor (layer3_outputs(632));
    layer4_outputs(529) <= (layer3_outputs(3967)) and not (layer3_outputs(4470));
    layer4_outputs(530) <= layer3_outputs(621);
    layer4_outputs(531) <= not(layer3_outputs(3291));
    layer4_outputs(532) <= not(layer3_outputs(4583));
    layer4_outputs(533) <= not(layer3_outputs(3253)) or (layer3_outputs(43));
    layer4_outputs(534) <= layer3_outputs(1882);
    layer4_outputs(535) <= not(layer3_outputs(2482)) or (layer3_outputs(3700));
    layer4_outputs(536) <= layer3_outputs(3664);
    layer4_outputs(537) <= not(layer3_outputs(1731)) or (layer3_outputs(2435));
    layer4_outputs(538) <= not(layer3_outputs(485));
    layer4_outputs(539) <= layer3_outputs(4357);
    layer4_outputs(540) <= not(layer3_outputs(619));
    layer4_outputs(541) <= not(layer3_outputs(1662));
    layer4_outputs(542) <= not((layer3_outputs(2218)) and (layer3_outputs(764)));
    layer4_outputs(543) <= layer3_outputs(3199);
    layer4_outputs(544) <= (layer3_outputs(4890)) and not (layer3_outputs(3800));
    layer4_outputs(545) <= layer3_outputs(1669);
    layer4_outputs(546) <= not(layer3_outputs(2975));
    layer4_outputs(547) <= not(layer3_outputs(949));
    layer4_outputs(548) <= (layer3_outputs(4075)) xor (layer3_outputs(738));
    layer4_outputs(549) <= layer3_outputs(2668);
    layer4_outputs(550) <= (layer3_outputs(4219)) and not (layer3_outputs(4037));
    layer4_outputs(551) <= layer3_outputs(2450);
    layer4_outputs(552) <= '1';
    layer4_outputs(553) <= (layer3_outputs(2626)) and not (layer3_outputs(5021));
    layer4_outputs(554) <= (layer3_outputs(2798)) and not (layer3_outputs(3808));
    layer4_outputs(555) <= layer3_outputs(2940);
    layer4_outputs(556) <= layer3_outputs(3932);
    layer4_outputs(557) <= not((layer3_outputs(1040)) or (layer3_outputs(2160)));
    layer4_outputs(558) <= not(layer3_outputs(29)) or (layer3_outputs(1874));
    layer4_outputs(559) <= '1';
    layer4_outputs(560) <= not(layer3_outputs(1414));
    layer4_outputs(561) <= not(layer3_outputs(3532));
    layer4_outputs(562) <= not(layer3_outputs(3810)) or (layer3_outputs(4930));
    layer4_outputs(563) <= (layer3_outputs(3635)) and not (layer3_outputs(806));
    layer4_outputs(564) <= not((layer3_outputs(4379)) or (layer3_outputs(3289)));
    layer4_outputs(565) <= layer3_outputs(4858);
    layer4_outputs(566) <= '0';
    layer4_outputs(567) <= not((layer3_outputs(668)) xor (layer3_outputs(3301)));
    layer4_outputs(568) <= layer3_outputs(4222);
    layer4_outputs(569) <= layer3_outputs(3011);
    layer4_outputs(570) <= layer3_outputs(941);
    layer4_outputs(571) <= layer3_outputs(5086);
    layer4_outputs(572) <= (layer3_outputs(4571)) and (layer3_outputs(1942));
    layer4_outputs(573) <= layer3_outputs(2062);
    layer4_outputs(574) <= not(layer3_outputs(901));
    layer4_outputs(575) <= layer3_outputs(2483);
    layer4_outputs(576) <= not(layer3_outputs(4482));
    layer4_outputs(577) <= not((layer3_outputs(4214)) or (layer3_outputs(2206)));
    layer4_outputs(578) <= not(layer3_outputs(1455)) or (layer3_outputs(2275));
    layer4_outputs(579) <= '1';
    layer4_outputs(580) <= layer3_outputs(211);
    layer4_outputs(581) <= not(layer3_outputs(3211));
    layer4_outputs(582) <= '1';
    layer4_outputs(583) <= (layer3_outputs(4628)) or (layer3_outputs(3826));
    layer4_outputs(584) <= not((layer3_outputs(2810)) xor (layer3_outputs(5097)));
    layer4_outputs(585) <= layer3_outputs(3583);
    layer4_outputs(586) <= layer3_outputs(4160);
    layer4_outputs(587) <= not(layer3_outputs(4367));
    layer4_outputs(588) <= (layer3_outputs(4660)) and not (layer3_outputs(4967));
    layer4_outputs(589) <= layer3_outputs(1905);
    layer4_outputs(590) <= not(layer3_outputs(3692)) or (layer3_outputs(3000));
    layer4_outputs(591) <= layer3_outputs(4913);
    layer4_outputs(592) <= '1';
    layer4_outputs(593) <= layer3_outputs(3358);
    layer4_outputs(594) <= '1';
    layer4_outputs(595) <= not(layer3_outputs(4648));
    layer4_outputs(596) <= '1';
    layer4_outputs(597) <= (layer3_outputs(1568)) and (layer3_outputs(767));
    layer4_outputs(598) <= not((layer3_outputs(281)) and (layer3_outputs(1433)));
    layer4_outputs(599) <= not(layer3_outputs(2894));
    layer4_outputs(600) <= not(layer3_outputs(2339)) or (layer3_outputs(2488));
    layer4_outputs(601) <= not(layer3_outputs(4378));
    layer4_outputs(602) <= not((layer3_outputs(3653)) or (layer3_outputs(2125)));
    layer4_outputs(603) <= '0';
    layer4_outputs(604) <= (layer3_outputs(4282)) or (layer3_outputs(4363));
    layer4_outputs(605) <= (layer3_outputs(4430)) and (layer3_outputs(804));
    layer4_outputs(606) <= not(layer3_outputs(554));
    layer4_outputs(607) <= layer3_outputs(4643);
    layer4_outputs(608) <= (layer3_outputs(3689)) and (layer3_outputs(3538));
    layer4_outputs(609) <= not(layer3_outputs(610));
    layer4_outputs(610) <= layer3_outputs(4607);
    layer4_outputs(611) <= layer3_outputs(2411);
    layer4_outputs(612) <= not(layer3_outputs(389)) or (layer3_outputs(1635));
    layer4_outputs(613) <= not(layer3_outputs(1272)) or (layer3_outputs(3899));
    layer4_outputs(614) <= not(layer3_outputs(3536));
    layer4_outputs(615) <= (layer3_outputs(3292)) and not (layer3_outputs(4551));
    layer4_outputs(616) <= not(layer3_outputs(3753)) or (layer3_outputs(3304));
    layer4_outputs(617) <= (layer3_outputs(519)) and (layer3_outputs(2731));
    layer4_outputs(618) <= layer3_outputs(751);
    layer4_outputs(619) <= not(layer3_outputs(702));
    layer4_outputs(620) <= not((layer3_outputs(4641)) or (layer3_outputs(663)));
    layer4_outputs(621) <= layer3_outputs(4026);
    layer4_outputs(622) <= not(layer3_outputs(3766));
    layer4_outputs(623) <= not(layer3_outputs(882));
    layer4_outputs(624) <= not(layer3_outputs(2466));
    layer4_outputs(625) <= (layer3_outputs(2497)) and not (layer3_outputs(861));
    layer4_outputs(626) <= not((layer3_outputs(3380)) or (layer3_outputs(4560)));
    layer4_outputs(627) <= layer3_outputs(376);
    layer4_outputs(628) <= not(layer3_outputs(5104)) or (layer3_outputs(4911));
    layer4_outputs(629) <= not((layer3_outputs(1837)) or (layer3_outputs(3888)));
    layer4_outputs(630) <= (layer3_outputs(1595)) and (layer3_outputs(1860));
    layer4_outputs(631) <= not(layer3_outputs(4778));
    layer4_outputs(632) <= layer3_outputs(1747);
    layer4_outputs(633) <= not((layer3_outputs(4823)) and (layer3_outputs(1294)));
    layer4_outputs(634) <= '0';
    layer4_outputs(635) <= layer3_outputs(3790);
    layer4_outputs(636) <= not((layer3_outputs(4785)) or (layer3_outputs(965)));
    layer4_outputs(637) <= (layer3_outputs(3979)) or (layer3_outputs(4765));
    layer4_outputs(638) <= not(layer3_outputs(1829));
    layer4_outputs(639) <= '1';
    layer4_outputs(640) <= not(layer3_outputs(1237));
    layer4_outputs(641) <= (layer3_outputs(1659)) or (layer3_outputs(4280));
    layer4_outputs(642) <= (layer3_outputs(2928)) and not (layer3_outputs(1069));
    layer4_outputs(643) <= not((layer3_outputs(3655)) or (layer3_outputs(2655)));
    layer4_outputs(644) <= layer3_outputs(2538);
    layer4_outputs(645) <= (layer3_outputs(2455)) xor (layer3_outputs(3005));
    layer4_outputs(646) <= not(layer3_outputs(2554));
    layer4_outputs(647) <= layer3_outputs(4437);
    layer4_outputs(648) <= not(layer3_outputs(3518));
    layer4_outputs(649) <= not(layer3_outputs(4919));
    layer4_outputs(650) <= layer3_outputs(2174);
    layer4_outputs(651) <= not((layer3_outputs(1651)) xor (layer3_outputs(3282)));
    layer4_outputs(652) <= layer3_outputs(947);
    layer4_outputs(653) <= not((layer3_outputs(1949)) or (layer3_outputs(1373)));
    layer4_outputs(654) <= '1';
    layer4_outputs(655) <= not(layer3_outputs(2641)) or (layer3_outputs(1598));
    layer4_outputs(656) <= not(layer3_outputs(4200)) or (layer3_outputs(3788));
    layer4_outputs(657) <= not(layer3_outputs(2459));
    layer4_outputs(658) <= not((layer3_outputs(1611)) or (layer3_outputs(4166)));
    layer4_outputs(659) <= (layer3_outputs(1108)) and (layer3_outputs(4939));
    layer4_outputs(660) <= layer3_outputs(778);
    layer4_outputs(661) <= (layer3_outputs(1824)) or (layer3_outputs(1908));
    layer4_outputs(662) <= not(layer3_outputs(474));
    layer4_outputs(663) <= not((layer3_outputs(3148)) xor (layer3_outputs(2470)));
    layer4_outputs(664) <= not(layer3_outputs(3327)) or (layer3_outputs(857));
    layer4_outputs(665) <= (layer3_outputs(194)) and (layer3_outputs(3107));
    layer4_outputs(666) <= layer3_outputs(2787);
    layer4_outputs(667) <= not(layer3_outputs(206)) or (layer3_outputs(1699));
    layer4_outputs(668) <= not((layer3_outputs(2280)) xor (layer3_outputs(1316)));
    layer4_outputs(669) <= not(layer3_outputs(2427));
    layer4_outputs(670) <= layer3_outputs(4505);
    layer4_outputs(671) <= '1';
    layer4_outputs(672) <= layer3_outputs(1892);
    layer4_outputs(673) <= '1';
    layer4_outputs(674) <= layer3_outputs(2147);
    layer4_outputs(675) <= '0';
    layer4_outputs(676) <= not(layer3_outputs(4506));
    layer4_outputs(677) <= not(layer3_outputs(817));
    layer4_outputs(678) <= (layer3_outputs(5073)) and (layer3_outputs(3325));
    layer4_outputs(679) <= (layer3_outputs(2559)) and not (layer3_outputs(3772));
    layer4_outputs(680) <= layer3_outputs(4901);
    layer4_outputs(681) <= layer3_outputs(3104);
    layer4_outputs(682) <= not(layer3_outputs(3915));
    layer4_outputs(683) <= not(layer3_outputs(177)) or (layer3_outputs(4200));
    layer4_outputs(684) <= not(layer3_outputs(3912)) or (layer3_outputs(2705));
    layer4_outputs(685) <= not(layer3_outputs(2839));
    layer4_outputs(686) <= not(layer3_outputs(4825));
    layer4_outputs(687) <= not(layer3_outputs(1371)) or (layer3_outputs(502));
    layer4_outputs(688) <= (layer3_outputs(4609)) and (layer3_outputs(355));
    layer4_outputs(689) <= layer3_outputs(1452);
    layer4_outputs(690) <= (layer3_outputs(3023)) and not (layer3_outputs(4449));
    layer4_outputs(691) <= '0';
    layer4_outputs(692) <= (layer3_outputs(1010)) and (layer3_outputs(892));
    layer4_outputs(693) <= not(layer3_outputs(4553));
    layer4_outputs(694) <= (layer3_outputs(3293)) xor (layer3_outputs(1930));
    layer4_outputs(695) <= (layer3_outputs(4677)) or (layer3_outputs(742));
    layer4_outputs(696) <= not((layer3_outputs(1335)) and (layer3_outputs(397)));
    layer4_outputs(697) <= not(layer3_outputs(3278)) or (layer3_outputs(4771));
    layer4_outputs(698) <= not(layer3_outputs(2360)) or (layer3_outputs(4081));
    layer4_outputs(699) <= not(layer3_outputs(3421)) or (layer3_outputs(2456));
    layer4_outputs(700) <= not(layer3_outputs(4667));
    layer4_outputs(701) <= layer3_outputs(2567);
    layer4_outputs(702) <= not((layer3_outputs(4058)) and (layer3_outputs(4755)));
    layer4_outputs(703) <= layer3_outputs(2358);
    layer4_outputs(704) <= '1';
    layer4_outputs(705) <= not(layer3_outputs(635));
    layer4_outputs(706) <= '1';
    layer4_outputs(707) <= layer3_outputs(795);
    layer4_outputs(708) <= not(layer3_outputs(1809));
    layer4_outputs(709) <= layer3_outputs(4749);
    layer4_outputs(710) <= not((layer3_outputs(3717)) xor (layer3_outputs(4595)));
    layer4_outputs(711) <= not((layer3_outputs(155)) xor (layer3_outputs(762)));
    layer4_outputs(712) <= not(layer3_outputs(189));
    layer4_outputs(713) <= layer3_outputs(4546);
    layer4_outputs(714) <= not(layer3_outputs(2811)) or (layer3_outputs(3230));
    layer4_outputs(715) <= not(layer3_outputs(642));
    layer4_outputs(716) <= (layer3_outputs(4727)) xor (layer3_outputs(4269));
    layer4_outputs(717) <= not((layer3_outputs(3515)) and (layer3_outputs(871)));
    layer4_outputs(718) <= not(layer3_outputs(663)) or (layer3_outputs(3467));
    layer4_outputs(719) <= not(layer3_outputs(2444)) or (layer3_outputs(5000));
    layer4_outputs(720) <= not((layer3_outputs(4382)) xor (layer3_outputs(2057)));
    layer4_outputs(721) <= layer3_outputs(205);
    layer4_outputs(722) <= layer3_outputs(1460);
    layer4_outputs(723) <= not(layer3_outputs(3997));
    layer4_outputs(724) <= '1';
    layer4_outputs(725) <= layer3_outputs(4419);
    layer4_outputs(726) <= layer3_outputs(4529);
    layer4_outputs(727) <= not(layer3_outputs(1437));
    layer4_outputs(728) <= not(layer3_outputs(3579));
    layer4_outputs(729) <= not(layer3_outputs(1637)) or (layer3_outputs(4981));
    layer4_outputs(730) <= layer3_outputs(1817);
    layer4_outputs(731) <= '0';
    layer4_outputs(732) <= not(layer3_outputs(685));
    layer4_outputs(733) <= layer3_outputs(504);
    layer4_outputs(734) <= not(layer3_outputs(510));
    layer4_outputs(735) <= layer3_outputs(758);
    layer4_outputs(736) <= not(layer3_outputs(171)) or (layer3_outputs(196));
    layer4_outputs(737) <= (layer3_outputs(2062)) and not (layer3_outputs(2318));
    layer4_outputs(738) <= '1';
    layer4_outputs(739) <= (layer3_outputs(2440)) and (layer3_outputs(2669));
    layer4_outputs(740) <= not(layer3_outputs(3777));
    layer4_outputs(741) <= layer3_outputs(4365);
    layer4_outputs(742) <= not(layer3_outputs(2867));
    layer4_outputs(743) <= not(layer3_outputs(5061));
    layer4_outputs(744) <= (layer3_outputs(2337)) and (layer3_outputs(269));
    layer4_outputs(745) <= layer3_outputs(1920);
    layer4_outputs(746) <= not(layer3_outputs(4284));
    layer4_outputs(747) <= not((layer3_outputs(1071)) xor (layer3_outputs(4384)));
    layer4_outputs(748) <= not((layer3_outputs(310)) xor (layer3_outputs(3654)));
    layer4_outputs(749) <= layer3_outputs(3573);
    layer4_outputs(750) <= not(layer3_outputs(318));
    layer4_outputs(751) <= (layer3_outputs(679)) or (layer3_outputs(2583));
    layer4_outputs(752) <= '0';
    layer4_outputs(753) <= not(layer3_outputs(794)) or (layer3_outputs(373));
    layer4_outputs(754) <= not((layer3_outputs(1408)) or (layer3_outputs(1862)));
    layer4_outputs(755) <= not(layer3_outputs(445)) or (layer3_outputs(2869));
    layer4_outputs(756) <= (layer3_outputs(4809)) and (layer3_outputs(3421));
    layer4_outputs(757) <= '0';
    layer4_outputs(758) <= layer3_outputs(3937);
    layer4_outputs(759) <= (layer3_outputs(5026)) and not (layer3_outputs(2519));
    layer4_outputs(760) <= not((layer3_outputs(1026)) and (layer3_outputs(327)));
    layer4_outputs(761) <= not((layer3_outputs(1880)) and (layer3_outputs(1065)));
    layer4_outputs(762) <= layer3_outputs(2946);
    layer4_outputs(763) <= layer3_outputs(3844);
    layer4_outputs(764) <= (layer3_outputs(4049)) and not (layer3_outputs(1674));
    layer4_outputs(765) <= (layer3_outputs(343)) or (layer3_outputs(1202));
    layer4_outputs(766) <= layer3_outputs(1746);
    layer4_outputs(767) <= (layer3_outputs(1801)) and (layer3_outputs(893));
    layer4_outputs(768) <= not(layer3_outputs(3352));
    layer4_outputs(769) <= (layer3_outputs(445)) and (layer3_outputs(3529));
    layer4_outputs(770) <= layer3_outputs(304);
    layer4_outputs(771) <= (layer3_outputs(2809)) and (layer3_outputs(4119));
    layer4_outputs(772) <= (layer3_outputs(903)) and (layer3_outputs(3958));
    layer4_outputs(773) <= (layer3_outputs(3839)) and not (layer3_outputs(809));
    layer4_outputs(774) <= (layer3_outputs(4304)) and not (layer3_outputs(1102));
    layer4_outputs(775) <= not(layer3_outputs(1728));
    layer4_outputs(776) <= (layer3_outputs(3405)) or (layer3_outputs(273));
    layer4_outputs(777) <= layer3_outputs(2666);
    layer4_outputs(778) <= layer3_outputs(1624);
    layer4_outputs(779) <= not(layer3_outputs(3694));
    layer4_outputs(780) <= (layer3_outputs(4955)) and (layer3_outputs(2916));
    layer4_outputs(781) <= not(layer3_outputs(64));
    layer4_outputs(782) <= not((layer3_outputs(2324)) and (layer3_outputs(3323)));
    layer4_outputs(783) <= layer3_outputs(849);
    layer4_outputs(784) <= (layer3_outputs(122)) and not (layer3_outputs(1278));
    layer4_outputs(785) <= (layer3_outputs(4892)) or (layer3_outputs(3804));
    layer4_outputs(786) <= not(layer3_outputs(4364));
    layer4_outputs(787) <= not(layer3_outputs(2833));
    layer4_outputs(788) <= not(layer3_outputs(4423));
    layer4_outputs(789) <= not((layer3_outputs(1759)) or (layer3_outputs(2615)));
    layer4_outputs(790) <= layer3_outputs(2695);
    layer4_outputs(791) <= not(layer3_outputs(2708)) or (layer3_outputs(351));
    layer4_outputs(792) <= not(layer3_outputs(1954));
    layer4_outputs(793) <= not((layer3_outputs(4454)) xor (layer3_outputs(4078)));
    layer4_outputs(794) <= not(layer3_outputs(1258));
    layer4_outputs(795) <= (layer3_outputs(1175)) and (layer3_outputs(1877));
    layer4_outputs(796) <= not(layer3_outputs(5101));
    layer4_outputs(797) <= not(layer3_outputs(4897)) or (layer3_outputs(2935));
    layer4_outputs(798) <= layer3_outputs(4692);
    layer4_outputs(799) <= not(layer3_outputs(4594));
    layer4_outputs(800) <= layer3_outputs(4218);
    layer4_outputs(801) <= not(layer3_outputs(1789));
    layer4_outputs(802) <= not((layer3_outputs(1173)) or (layer3_outputs(4320)));
    layer4_outputs(803) <= not(layer3_outputs(3032));
    layer4_outputs(804) <= (layer3_outputs(3413)) and not (layer3_outputs(2490));
    layer4_outputs(805) <= not(layer3_outputs(2523));
    layer4_outputs(806) <= '0';
    layer4_outputs(807) <= layer3_outputs(2824);
    layer4_outputs(808) <= not(layer3_outputs(4228));
    layer4_outputs(809) <= '1';
    layer4_outputs(810) <= not(layer3_outputs(686));
    layer4_outputs(811) <= layer3_outputs(3390);
    layer4_outputs(812) <= not(layer3_outputs(182));
    layer4_outputs(813) <= not(layer3_outputs(198));
    layer4_outputs(814) <= not(layer3_outputs(104)) or (layer3_outputs(3743));
    layer4_outputs(815) <= not(layer3_outputs(651));
    layer4_outputs(816) <= '0';
    layer4_outputs(817) <= not(layer3_outputs(3815));
    layer4_outputs(818) <= (layer3_outputs(3625)) and not (layer3_outputs(2540));
    layer4_outputs(819) <= not(layer3_outputs(220)) or (layer3_outputs(2235));
    layer4_outputs(820) <= not(layer3_outputs(3440));
    layer4_outputs(821) <= layer3_outputs(363);
    layer4_outputs(822) <= layer3_outputs(1932);
    layer4_outputs(823) <= not((layer3_outputs(311)) and (layer3_outputs(3109)));
    layer4_outputs(824) <= not(layer3_outputs(250));
    layer4_outputs(825) <= not(layer3_outputs(4801));
    layer4_outputs(826) <= not((layer3_outputs(3182)) xor (layer3_outputs(396)));
    layer4_outputs(827) <= (layer3_outputs(4487)) or (layer3_outputs(1170));
    layer4_outputs(828) <= not(layer3_outputs(3639)) or (layer3_outputs(17));
    layer4_outputs(829) <= not(layer3_outputs(2547));
    layer4_outputs(830) <= not((layer3_outputs(1643)) and (layer3_outputs(869)));
    layer4_outputs(831) <= not(layer3_outputs(3820)) or (layer3_outputs(4690));
    layer4_outputs(832) <= (layer3_outputs(2387)) or (layer3_outputs(744));
    layer4_outputs(833) <= not((layer3_outputs(5037)) or (layer3_outputs(2853)));
    layer4_outputs(834) <= (layer3_outputs(1476)) and not (layer3_outputs(626));
    layer4_outputs(835) <= not(layer3_outputs(4766));
    layer4_outputs(836) <= not((layer3_outputs(1622)) or (layer3_outputs(4579)));
    layer4_outputs(837) <= not((layer3_outputs(2020)) or (layer3_outputs(3286)));
    layer4_outputs(838) <= layer3_outputs(2213);
    layer4_outputs(839) <= '1';
    layer4_outputs(840) <= not(layer3_outputs(5112)) or (layer3_outputs(5078));
    layer4_outputs(841) <= not(layer3_outputs(2590));
    layer4_outputs(842) <= not(layer3_outputs(3137)) or (layer3_outputs(4728));
    layer4_outputs(843) <= not(layer3_outputs(1750));
    layer4_outputs(844) <= not(layer3_outputs(3424));
    layer4_outputs(845) <= (layer3_outputs(2842)) and not (layer3_outputs(552));
    layer4_outputs(846) <= not(layer3_outputs(1113));
    layer4_outputs(847) <= '1';
    layer4_outputs(848) <= (layer3_outputs(60)) and not (layer3_outputs(4411));
    layer4_outputs(849) <= (layer3_outputs(2220)) and (layer3_outputs(523));
    layer4_outputs(850) <= not(layer3_outputs(2828));
    layer4_outputs(851) <= (layer3_outputs(4190)) and (layer3_outputs(2158));
    layer4_outputs(852) <= (layer3_outputs(1192)) or (layer3_outputs(2472));
    layer4_outputs(853) <= (layer3_outputs(1206)) and not (layer3_outputs(2281));
    layer4_outputs(854) <= not((layer3_outputs(3093)) or (layer3_outputs(2038)));
    layer4_outputs(855) <= (layer3_outputs(2423)) and not (layer3_outputs(4460));
    layer4_outputs(856) <= layer3_outputs(3233);
    layer4_outputs(857) <= not(layer3_outputs(2602));
    layer4_outputs(858) <= not(layer3_outputs(4268));
    layer4_outputs(859) <= layer3_outputs(4634);
    layer4_outputs(860) <= layer3_outputs(4946);
    layer4_outputs(861) <= layer3_outputs(2043);
    layer4_outputs(862) <= (layer3_outputs(866)) or (layer3_outputs(1134));
    layer4_outputs(863) <= '1';
    layer4_outputs(864) <= (layer3_outputs(1720)) or (layer3_outputs(4834));
    layer4_outputs(865) <= not(layer3_outputs(779));
    layer4_outputs(866) <= not((layer3_outputs(4663)) or (layer3_outputs(4399)));
    layer4_outputs(867) <= '1';
    layer4_outputs(868) <= layer3_outputs(4715);
    layer4_outputs(869) <= not(layer3_outputs(1921));
    layer4_outputs(870) <= not(layer3_outputs(4306));
    layer4_outputs(871) <= not(layer3_outputs(4907));
    layer4_outputs(872) <= not((layer3_outputs(202)) and (layer3_outputs(2870)));
    layer4_outputs(873) <= (layer3_outputs(2545)) and not (layer3_outputs(4797));
    layer4_outputs(874) <= (layer3_outputs(1000)) and not (layer3_outputs(2286));
    layer4_outputs(875) <= layer3_outputs(2085);
    layer4_outputs(876) <= not(layer3_outputs(3970));
    layer4_outputs(877) <= (layer3_outputs(4805)) and not (layer3_outputs(998));
    layer4_outputs(878) <= not(layer3_outputs(3083)) or (layer3_outputs(1164));
    layer4_outputs(879) <= '0';
    layer4_outputs(880) <= not(layer3_outputs(367));
    layer4_outputs(881) <= not(layer3_outputs(2071));
    layer4_outputs(882) <= not(layer3_outputs(2966)) or (layer3_outputs(3343));
    layer4_outputs(883) <= '1';
    layer4_outputs(884) <= (layer3_outputs(3051)) and (layer3_outputs(3624));
    layer4_outputs(885) <= layer3_outputs(3228);
    layer4_outputs(886) <= '0';
    layer4_outputs(887) <= (layer3_outputs(3672)) and not (layer3_outputs(2825));
    layer4_outputs(888) <= not(layer3_outputs(1530));
    layer4_outputs(889) <= not((layer3_outputs(2167)) and (layer3_outputs(696)));
    layer4_outputs(890) <= not(layer3_outputs(3244));
    layer4_outputs(891) <= layer3_outputs(25);
    layer4_outputs(892) <= layer3_outputs(1969);
    layer4_outputs(893) <= not((layer3_outputs(4503)) and (layer3_outputs(692)));
    layer4_outputs(894) <= not((layer3_outputs(3411)) and (layer3_outputs(2154)));
    layer4_outputs(895) <= (layer3_outputs(69)) and (layer3_outputs(1101));
    layer4_outputs(896) <= (layer3_outputs(2860)) and not (layer3_outputs(584));
    layer4_outputs(897) <= layer3_outputs(4032);
    layer4_outputs(898) <= layer3_outputs(1927);
    layer4_outputs(899) <= (layer3_outputs(1629)) or (layer3_outputs(2660));
    layer4_outputs(900) <= layer3_outputs(2733);
    layer4_outputs(901) <= not((layer3_outputs(572)) and (layer3_outputs(3271)));
    layer4_outputs(902) <= (layer3_outputs(2503)) and (layer3_outputs(800));
    layer4_outputs(903) <= (layer3_outputs(4608)) xor (layer3_outputs(3800));
    layer4_outputs(904) <= '0';
    layer4_outputs(905) <= not(layer3_outputs(4515));
    layer4_outputs(906) <= layer3_outputs(2983);
    layer4_outputs(907) <= not((layer3_outputs(2786)) or (layer3_outputs(3143)));
    layer4_outputs(908) <= not(layer3_outputs(430));
    layer4_outputs(909) <= not(layer3_outputs(71));
    layer4_outputs(910) <= not(layer3_outputs(2251)) or (layer3_outputs(3409));
    layer4_outputs(911) <= not(layer3_outputs(3157));
    layer4_outputs(912) <= not(layer3_outputs(4464)) or (layer3_outputs(125));
    layer4_outputs(913) <= not(layer3_outputs(1467));
    layer4_outputs(914) <= not(layer3_outputs(235));
    layer4_outputs(915) <= layer3_outputs(2470);
    layer4_outputs(916) <= (layer3_outputs(1973)) and not (layer3_outputs(1417));
    layer4_outputs(917) <= not(layer3_outputs(2090));
    layer4_outputs(918) <= (layer3_outputs(1825)) and (layer3_outputs(3723));
    layer4_outputs(919) <= (layer3_outputs(3452)) and not (layer3_outputs(3633));
    layer4_outputs(920) <= not((layer3_outputs(2044)) and (layer3_outputs(4937)));
    layer4_outputs(921) <= not(layer3_outputs(2092));
    layer4_outputs(922) <= not(layer3_outputs(1499));
    layer4_outputs(923) <= layer3_outputs(31);
    layer4_outputs(924) <= layer3_outputs(2850);
    layer4_outputs(925) <= '0';
    layer4_outputs(926) <= layer3_outputs(1851);
    layer4_outputs(927) <= '1';
    layer4_outputs(928) <= not((layer3_outputs(3972)) or (layer3_outputs(2259)));
    layer4_outputs(929) <= (layer3_outputs(1553)) or (layer3_outputs(3331));
    layer4_outputs(930) <= '1';
    layer4_outputs(931) <= not(layer3_outputs(1740));
    layer4_outputs(932) <= not(layer3_outputs(1061));
    layer4_outputs(933) <= layer3_outputs(3492);
    layer4_outputs(934) <= not(layer3_outputs(4715));
    layer4_outputs(935) <= not((layer3_outputs(79)) and (layer3_outputs(646)));
    layer4_outputs(936) <= (layer3_outputs(1870)) and not (layer3_outputs(5028));
    layer4_outputs(937) <= '1';
    layer4_outputs(938) <= (layer3_outputs(2107)) and not (layer3_outputs(1240));
    layer4_outputs(939) <= '1';
    layer4_outputs(940) <= '0';
    layer4_outputs(941) <= (layer3_outputs(1409)) and not (layer3_outputs(1603));
    layer4_outputs(942) <= not(layer3_outputs(3823));
    layer4_outputs(943) <= layer3_outputs(1415);
    layer4_outputs(944) <= (layer3_outputs(4113)) and not (layer3_outputs(4745));
    layer4_outputs(945) <= layer3_outputs(2268);
    layer4_outputs(946) <= (layer3_outputs(2002)) xor (layer3_outputs(2433));
    layer4_outputs(947) <= not(layer3_outputs(2228));
    layer4_outputs(948) <= not(layer3_outputs(2030)) or (layer3_outputs(115));
    layer4_outputs(949) <= not((layer3_outputs(4000)) and (layer3_outputs(206)));
    layer4_outputs(950) <= not((layer3_outputs(2017)) xor (layer3_outputs(4222)));
    layer4_outputs(951) <= not((layer3_outputs(3196)) xor (layer3_outputs(419)));
    layer4_outputs(952) <= not(layer3_outputs(2658)) or (layer3_outputs(1686));
    layer4_outputs(953) <= (layer3_outputs(875)) and (layer3_outputs(414));
    layer4_outputs(954) <= layer3_outputs(2560);
    layer4_outputs(955) <= (layer3_outputs(2720)) or (layer3_outputs(1103));
    layer4_outputs(956) <= not(layer3_outputs(4973)) or (layer3_outputs(2543));
    layer4_outputs(957) <= not((layer3_outputs(2045)) or (layer3_outputs(4957)));
    layer4_outputs(958) <= layer3_outputs(4737);
    layer4_outputs(959) <= layer3_outputs(3065);
    layer4_outputs(960) <= (layer3_outputs(4011)) and (layer3_outputs(3175));
    layer4_outputs(961) <= not((layer3_outputs(244)) xor (layer3_outputs(1360)));
    layer4_outputs(962) <= layer3_outputs(1665);
    layer4_outputs(963) <= not((layer3_outputs(251)) xor (layer3_outputs(4316)));
    layer4_outputs(964) <= not((layer3_outputs(1813)) and (layer3_outputs(3723)));
    layer4_outputs(965) <= (layer3_outputs(1800)) and (layer3_outputs(4145));
    layer4_outputs(966) <= not(layer3_outputs(4478)) or (layer3_outputs(2700));
    layer4_outputs(967) <= '1';
    layer4_outputs(968) <= layer3_outputs(1566);
    layer4_outputs(969) <= not(layer3_outputs(2589));
    layer4_outputs(970) <= not((layer3_outputs(97)) and (layer3_outputs(1964)));
    layer4_outputs(971) <= (layer3_outputs(1189)) and not (layer3_outputs(2205));
    layer4_outputs(972) <= not(layer3_outputs(2448)) or (layer3_outputs(91));
    layer4_outputs(973) <= not(layer3_outputs(3704));
    layer4_outputs(974) <= layer3_outputs(3915);
    layer4_outputs(975) <= layer3_outputs(3733);
    layer4_outputs(976) <= '1';
    layer4_outputs(977) <= '0';
    layer4_outputs(978) <= '0';
    layer4_outputs(979) <= not(layer3_outputs(3583));
    layer4_outputs(980) <= not(layer3_outputs(212));
    layer4_outputs(981) <= not(layer3_outputs(1262)) or (layer3_outputs(3076));
    layer4_outputs(982) <= (layer3_outputs(4864)) or (layer3_outputs(2261));
    layer4_outputs(983) <= not((layer3_outputs(239)) and (layer3_outputs(471)));
    layer4_outputs(984) <= layer3_outputs(20);
    layer4_outputs(985) <= (layer3_outputs(1082)) or (layer3_outputs(1268));
    layer4_outputs(986) <= not(layer3_outputs(3686));
    layer4_outputs(987) <= (layer3_outputs(5108)) or (layer3_outputs(3701));
    layer4_outputs(988) <= (layer3_outputs(562)) and not (layer3_outputs(2130));
    layer4_outputs(989) <= (layer3_outputs(3560)) or (layer3_outputs(4520));
    layer4_outputs(990) <= '0';
    layer4_outputs(991) <= not(layer3_outputs(1264));
    layer4_outputs(992) <= not(layer3_outputs(4243));
    layer4_outputs(993) <= layer3_outputs(1881);
    layer4_outputs(994) <= layer3_outputs(2637);
    layer4_outputs(995) <= not(layer3_outputs(3944));
    layer4_outputs(996) <= layer3_outputs(4611);
    layer4_outputs(997) <= '0';
    layer4_outputs(998) <= (layer3_outputs(4919)) and not (layer3_outputs(442));
    layer4_outputs(999) <= not(layer3_outputs(4099));
    layer4_outputs(1000) <= not(layer3_outputs(277)) or (layer3_outputs(4706));
    layer4_outputs(1001) <= not(layer3_outputs(4866)) or (layer3_outputs(5051));
    layer4_outputs(1002) <= not(layer3_outputs(460));
    layer4_outputs(1003) <= not(layer3_outputs(4294));
    layer4_outputs(1004) <= not(layer3_outputs(2818));
    layer4_outputs(1005) <= '1';
    layer4_outputs(1006) <= not(layer3_outputs(1431));
    layer4_outputs(1007) <= not(layer3_outputs(4434));
    layer4_outputs(1008) <= not((layer3_outputs(5112)) xor (layer3_outputs(930)));
    layer4_outputs(1009) <= not(layer3_outputs(896));
    layer4_outputs(1010) <= layer3_outputs(3219);
    layer4_outputs(1011) <= '1';
    layer4_outputs(1012) <= not(layer3_outputs(394)) or (layer3_outputs(1891));
    layer4_outputs(1013) <= not(layer3_outputs(522));
    layer4_outputs(1014) <= not((layer3_outputs(2431)) or (layer3_outputs(636)));
    layer4_outputs(1015) <= (layer3_outputs(2616)) and (layer3_outputs(1841));
    layer4_outputs(1016) <= layer3_outputs(2575);
    layer4_outputs(1017) <= (layer3_outputs(1426)) and not (layer3_outputs(2770));
    layer4_outputs(1018) <= layer3_outputs(2790);
    layer4_outputs(1019) <= layer3_outputs(4746);
    layer4_outputs(1020) <= layer3_outputs(1514);
    layer4_outputs(1021) <= not(layer3_outputs(1940));
    layer4_outputs(1022) <= '1';
    layer4_outputs(1023) <= not(layer3_outputs(268)) or (layer3_outputs(3741));
    layer4_outputs(1024) <= not((layer3_outputs(2697)) or (layer3_outputs(1213)));
    layer4_outputs(1025) <= layer3_outputs(466);
    layer4_outputs(1026) <= layer3_outputs(4269);
    layer4_outputs(1027) <= layer3_outputs(3985);
    layer4_outputs(1028) <= '1';
    layer4_outputs(1029) <= layer3_outputs(3473);
    layer4_outputs(1030) <= not(layer3_outputs(4704));
    layer4_outputs(1031) <= not((layer3_outputs(2129)) xor (layer3_outputs(2673)));
    layer4_outputs(1032) <= not(layer3_outputs(4954)) or (layer3_outputs(4665));
    layer4_outputs(1033) <= (layer3_outputs(4215)) and not (layer3_outputs(935));
    layer4_outputs(1034) <= not(layer3_outputs(2184)) or (layer3_outputs(5065));
    layer4_outputs(1035) <= (layer3_outputs(2049)) and not (layer3_outputs(4009));
    layer4_outputs(1036) <= (layer3_outputs(4187)) and not (layer3_outputs(3748));
    layer4_outputs(1037) <= not(layer3_outputs(2937)) or (layer3_outputs(2905));
    layer4_outputs(1038) <= not((layer3_outputs(1330)) xor (layer3_outputs(1727)));
    layer4_outputs(1039) <= not(layer3_outputs(2415));
    layer4_outputs(1040) <= layer3_outputs(3407);
    layer4_outputs(1041) <= layer3_outputs(3509);
    layer4_outputs(1042) <= not((layer3_outputs(3382)) and (layer3_outputs(1088)));
    layer4_outputs(1043) <= not(layer3_outputs(4861));
    layer4_outputs(1044) <= (layer3_outputs(1141)) and not (layer3_outputs(3414));
    layer4_outputs(1045) <= (layer3_outputs(974)) and (layer3_outputs(4221));
    layer4_outputs(1046) <= (layer3_outputs(3801)) or (layer3_outputs(4617));
    layer4_outputs(1047) <= '1';
    layer4_outputs(1048) <= (layer3_outputs(68)) and (layer3_outputs(4768));
    layer4_outputs(1049) <= not(layer3_outputs(4518));
    layer4_outputs(1050) <= not(layer3_outputs(3217));
    layer4_outputs(1051) <= layer3_outputs(3526);
    layer4_outputs(1052) <= layer3_outputs(2441);
    layer4_outputs(1053) <= not(layer3_outputs(2866));
    layer4_outputs(1054) <= not(layer3_outputs(2745)) or (layer3_outputs(2614));
    layer4_outputs(1055) <= not(layer3_outputs(407));
    layer4_outputs(1056) <= not((layer3_outputs(3693)) or (layer3_outputs(2383)));
    layer4_outputs(1057) <= not(layer3_outputs(2389));
    layer4_outputs(1058) <= (layer3_outputs(1290)) and not (layer3_outputs(959));
    layer4_outputs(1059) <= not((layer3_outputs(1100)) and (layer3_outputs(2571)));
    layer4_outputs(1060) <= not((layer3_outputs(3136)) and (layer3_outputs(3824)));
    layer4_outputs(1061) <= '0';
    layer4_outputs(1062) <= (layer3_outputs(5074)) and (layer3_outputs(1444));
    layer4_outputs(1063) <= layer3_outputs(2761);
    layer4_outputs(1064) <= not(layer3_outputs(4367));
    layer4_outputs(1065) <= layer3_outputs(329);
    layer4_outputs(1066) <= '0';
    layer4_outputs(1067) <= (layer3_outputs(4492)) or (layer3_outputs(2711));
    layer4_outputs(1068) <= not(layer3_outputs(860));
    layer4_outputs(1069) <= (layer3_outputs(2121)) or (layer3_outputs(4489));
    layer4_outputs(1070) <= layer3_outputs(1281);
    layer4_outputs(1071) <= layer3_outputs(1000);
    layer4_outputs(1072) <= '1';
    layer4_outputs(1073) <= not(layer3_outputs(1773));
    layer4_outputs(1074) <= (layer3_outputs(740)) xor (layer3_outputs(4406));
    layer4_outputs(1075) <= layer3_outputs(2814);
    layer4_outputs(1076) <= not(layer3_outputs(2365));
    layer4_outputs(1077) <= not((layer3_outputs(4676)) and (layer3_outputs(2728)));
    layer4_outputs(1078) <= (layer3_outputs(2868)) or (layer3_outputs(867));
    layer4_outputs(1079) <= not(layer3_outputs(3989));
    layer4_outputs(1080) <= '1';
    layer4_outputs(1081) <= layer3_outputs(4232);
    layer4_outputs(1082) <= '1';
    layer4_outputs(1083) <= layer3_outputs(4534);
    layer4_outputs(1084) <= (layer3_outputs(4232)) and not (layer3_outputs(3736));
    layer4_outputs(1085) <= not(layer3_outputs(1868));
    layer4_outputs(1086) <= '0';
    layer4_outputs(1087) <= not((layer3_outputs(313)) and (layer3_outputs(2587)));
    layer4_outputs(1088) <= not(layer3_outputs(2455));
    layer4_outputs(1089) <= (layer3_outputs(408)) or (layer3_outputs(350));
    layer4_outputs(1090) <= (layer3_outputs(2051)) and not (layer3_outputs(3960));
    layer4_outputs(1091) <= '1';
    layer4_outputs(1092) <= layer3_outputs(3252);
    layer4_outputs(1093) <= not(layer3_outputs(2845));
    layer4_outputs(1094) <= not(layer3_outputs(4644));
    layer4_outputs(1095) <= layer3_outputs(4056);
    layer4_outputs(1096) <= not(layer3_outputs(427)) or (layer3_outputs(479));
    layer4_outputs(1097) <= layer3_outputs(3117);
    layer4_outputs(1098) <= (layer3_outputs(2239)) and not (layer3_outputs(3397));
    layer4_outputs(1099) <= (layer3_outputs(2676)) and (layer3_outputs(3751));
    layer4_outputs(1100) <= not(layer3_outputs(1223));
    layer4_outputs(1101) <= not(layer3_outputs(899)) or (layer3_outputs(3314));
    layer4_outputs(1102) <= not(layer3_outputs(4417));
    layer4_outputs(1103) <= layer3_outputs(2652);
    layer4_outputs(1104) <= not(layer3_outputs(2860)) or (layer3_outputs(1950));
    layer4_outputs(1105) <= layer3_outputs(2531);
    layer4_outputs(1106) <= not(layer3_outputs(832));
    layer4_outputs(1107) <= not(layer3_outputs(4332)) or (layer3_outputs(4658));
    layer4_outputs(1108) <= '0';
    layer4_outputs(1109) <= (layer3_outputs(2397)) and not (layer3_outputs(2813));
    layer4_outputs(1110) <= not((layer3_outputs(1807)) and (layer3_outputs(3599)));
    layer4_outputs(1111) <= '1';
    layer4_outputs(1112) <= (layer3_outputs(271)) or (layer3_outputs(1768));
    layer4_outputs(1113) <= not(layer3_outputs(2758));
    layer4_outputs(1114) <= not((layer3_outputs(3406)) or (layer3_outputs(5007)));
    layer4_outputs(1115) <= not(layer3_outputs(3426)) or (layer3_outputs(3675));
    layer4_outputs(1116) <= not((layer3_outputs(1999)) or (layer3_outputs(2690)));
    layer4_outputs(1117) <= not((layer3_outputs(2647)) or (layer3_outputs(3772)));
    layer4_outputs(1118) <= '1';
    layer4_outputs(1119) <= not(layer3_outputs(4853));
    layer4_outputs(1120) <= not(layer3_outputs(2066)) or (layer3_outputs(320));
    layer4_outputs(1121) <= not((layer3_outputs(1701)) xor (layer3_outputs(1235)));
    layer4_outputs(1122) <= (layer3_outputs(3310)) and not (layer3_outputs(4170));
    layer4_outputs(1123) <= '1';
    layer4_outputs(1124) <= '0';
    layer4_outputs(1125) <= layer3_outputs(2083);
    layer4_outputs(1126) <= (layer3_outputs(3430)) and not (layer3_outputs(268));
    layer4_outputs(1127) <= not(layer3_outputs(2376));
    layer4_outputs(1128) <= not(layer3_outputs(4437));
    layer4_outputs(1129) <= layer3_outputs(3149);
    layer4_outputs(1130) <= not(layer3_outputs(1609));
    layer4_outputs(1131) <= layer3_outputs(4557);
    layer4_outputs(1132) <= not(layer3_outputs(1444)) or (layer3_outputs(295));
    layer4_outputs(1133) <= not(layer3_outputs(80));
    layer4_outputs(1134) <= (layer3_outputs(2618)) or (layer3_outputs(88));
    layer4_outputs(1135) <= not((layer3_outputs(4335)) and (layer3_outputs(2353)));
    layer4_outputs(1136) <= layer3_outputs(2799);
    layer4_outputs(1137) <= (layer3_outputs(2929)) or (layer3_outputs(2209));
    layer4_outputs(1138) <= '1';
    layer4_outputs(1139) <= not(layer3_outputs(2111));
    layer4_outputs(1140) <= not((layer3_outputs(3067)) and (layer3_outputs(2254)));
    layer4_outputs(1141) <= not(layer3_outputs(1207));
    layer4_outputs(1142) <= not((layer3_outputs(4908)) or (layer3_outputs(1758)));
    layer4_outputs(1143) <= layer3_outputs(2658);
    layer4_outputs(1144) <= (layer3_outputs(652)) xor (layer3_outputs(1439));
    layer4_outputs(1145) <= '0';
    layer4_outputs(1146) <= (layer3_outputs(4954)) and (layer3_outputs(4198));
    layer4_outputs(1147) <= not(layer3_outputs(3506)) or (layer3_outputs(3394));
    layer4_outputs(1148) <= not(layer3_outputs(980));
    layer4_outputs(1149) <= layer3_outputs(4910);
    layer4_outputs(1150) <= not((layer3_outputs(2236)) or (layer3_outputs(928)));
    layer4_outputs(1151) <= (layer3_outputs(4951)) xor (layer3_outputs(2144));
    layer4_outputs(1152) <= not((layer3_outputs(3206)) xor (layer3_outputs(3101)));
    layer4_outputs(1153) <= layer3_outputs(2574);
    layer4_outputs(1154) <= layer3_outputs(1364);
    layer4_outputs(1155) <= not(layer3_outputs(3543));
    layer4_outputs(1156) <= not((layer3_outputs(1096)) or (layer3_outputs(1640)));
    layer4_outputs(1157) <= not(layer3_outputs(3943)) or (layer3_outputs(1723));
    layer4_outputs(1158) <= not(layer3_outputs(3243));
    layer4_outputs(1159) <= (layer3_outputs(2074)) and not (layer3_outputs(223));
    layer4_outputs(1160) <= (layer3_outputs(2994)) and (layer3_outputs(3992));
    layer4_outputs(1161) <= not(layer3_outputs(961));
    layer4_outputs(1162) <= not(layer3_outputs(4360));
    layer4_outputs(1163) <= not(layer3_outputs(2832)) or (layer3_outputs(4702));
    layer4_outputs(1164) <= (layer3_outputs(1322)) and (layer3_outputs(19));
    layer4_outputs(1165) <= layer3_outputs(2513);
    layer4_outputs(1166) <= not(layer3_outputs(4633));
    layer4_outputs(1167) <= (layer3_outputs(4791)) and not (layer3_outputs(623));
    layer4_outputs(1168) <= not(layer3_outputs(4618));
    layer4_outputs(1169) <= (layer3_outputs(3057)) and (layer3_outputs(4504));
    layer4_outputs(1170) <= (layer3_outputs(4828)) and (layer3_outputs(4714));
    layer4_outputs(1171) <= not(layer3_outputs(1769));
    layer4_outputs(1172) <= (layer3_outputs(153)) and (layer3_outputs(2113));
    layer4_outputs(1173) <= (layer3_outputs(4157)) xor (layer3_outputs(4568));
    layer4_outputs(1174) <= not(layer3_outputs(2592)) or (layer3_outputs(1182));
    layer4_outputs(1175) <= '0';
    layer4_outputs(1176) <= layer3_outputs(1125);
    layer4_outputs(1177) <= not((layer3_outputs(3795)) and (layer3_outputs(3168)));
    layer4_outputs(1178) <= not(layer3_outputs(4402));
    layer4_outputs(1179) <= layer3_outputs(634);
    layer4_outputs(1180) <= layer3_outputs(2464);
    layer4_outputs(1181) <= not(layer3_outputs(783));
    layer4_outputs(1182) <= not((layer3_outputs(4804)) or (layer3_outputs(3094)));
    layer4_outputs(1183) <= layer3_outputs(783);
    layer4_outputs(1184) <= (layer3_outputs(79)) and not (layer3_outputs(2308));
    layer4_outputs(1185) <= (layer3_outputs(4872)) and not (layer3_outputs(1490));
    layer4_outputs(1186) <= layer3_outputs(3877);
    layer4_outputs(1187) <= not(layer3_outputs(2584));
    layer4_outputs(1188) <= layer3_outputs(205);
    layer4_outputs(1189) <= not((layer3_outputs(2608)) and (layer3_outputs(1685)));
    layer4_outputs(1190) <= not(layer3_outputs(4739));
    layer4_outputs(1191) <= layer3_outputs(4902);
    layer4_outputs(1192) <= not(layer3_outputs(329));
    layer4_outputs(1193) <= layer3_outputs(1592);
    layer4_outputs(1194) <= not(layer3_outputs(3817));
    layer4_outputs(1195) <= layer3_outputs(3497);
    layer4_outputs(1196) <= layer3_outputs(3013);
    layer4_outputs(1197) <= not(layer3_outputs(634)) or (layer3_outputs(4653));
    layer4_outputs(1198) <= not((layer3_outputs(1679)) xor (layer3_outputs(4976)));
    layer4_outputs(1199) <= not(layer3_outputs(2939)) or (layer3_outputs(1885));
    layer4_outputs(1200) <= (layer3_outputs(2677)) and not (layer3_outputs(4896));
    layer4_outputs(1201) <= not(layer3_outputs(4788)) or (layer3_outputs(3893));
    layer4_outputs(1202) <= '0';
    layer4_outputs(1203) <= not(layer3_outputs(1550));
    layer4_outputs(1204) <= not((layer3_outputs(1276)) or (layer3_outputs(2014)));
    layer4_outputs(1205) <= (layer3_outputs(3829)) and (layer3_outputs(1521));
    layer4_outputs(1206) <= not(layer3_outputs(2659));
    layer4_outputs(1207) <= not(layer3_outputs(38));
    layer4_outputs(1208) <= not(layer3_outputs(2249)) or (layer3_outputs(1458));
    layer4_outputs(1209) <= not(layer3_outputs(515)) or (layer3_outputs(1807));
    layer4_outputs(1210) <= layer3_outputs(3719);
    layer4_outputs(1211) <= (layer3_outputs(4778)) or (layer3_outputs(3713));
    layer4_outputs(1212) <= (layer3_outputs(1917)) or (layer3_outputs(4095));
    layer4_outputs(1213) <= not(layer3_outputs(2586));
    layer4_outputs(1214) <= (layer3_outputs(799)) and not (layer3_outputs(1716));
    layer4_outputs(1215) <= (layer3_outputs(3841)) and not (layer3_outputs(2756));
    layer4_outputs(1216) <= layer3_outputs(1210);
    layer4_outputs(1217) <= not(layer3_outputs(3536));
    layer4_outputs(1218) <= not(layer3_outputs(1714));
    layer4_outputs(1219) <= not(layer3_outputs(1663));
    layer4_outputs(1220) <= layer3_outputs(2611);
    layer4_outputs(1221) <= not((layer3_outputs(2953)) and (layer3_outputs(4578)));
    layer4_outputs(1222) <= (layer3_outputs(1670)) and (layer3_outputs(3570));
    layer4_outputs(1223) <= layer3_outputs(4773);
    layer4_outputs(1224) <= layer3_outputs(3255);
    layer4_outputs(1225) <= layer3_outputs(1403);
    layer4_outputs(1226) <= not(layer3_outputs(1117)) or (layer3_outputs(2175));
    layer4_outputs(1227) <= layer3_outputs(2048);
    layer4_outputs(1228) <= not(layer3_outputs(1500));
    layer4_outputs(1229) <= (layer3_outputs(4965)) and (layer3_outputs(3581));
    layer4_outputs(1230) <= (layer3_outputs(4329)) xor (layer3_outputs(3643));
    layer4_outputs(1231) <= layer3_outputs(2796);
    layer4_outputs(1232) <= not(layer3_outputs(3046)) or (layer3_outputs(1325));
    layer4_outputs(1233) <= not(layer3_outputs(461));
    layer4_outputs(1234) <= not(layer3_outputs(2800));
    layer4_outputs(1235) <= (layer3_outputs(2413)) and (layer3_outputs(1722));
    layer4_outputs(1236) <= not((layer3_outputs(4097)) xor (layer3_outputs(4799)));
    layer4_outputs(1237) <= (layer3_outputs(1320)) and (layer3_outputs(4030));
    layer4_outputs(1238) <= '1';
    layer4_outputs(1239) <= not((layer3_outputs(1650)) and (layer3_outputs(3798)));
    layer4_outputs(1240) <= not(layer3_outputs(1709));
    layer4_outputs(1241) <= not(layer3_outputs(1230));
    layer4_outputs(1242) <= (layer3_outputs(922)) and not (layer3_outputs(2039));
    layer4_outputs(1243) <= '1';
    layer4_outputs(1244) <= layer3_outputs(1347);
    layer4_outputs(1245) <= not((layer3_outputs(1360)) xor (layer3_outputs(2834)));
    layer4_outputs(1246) <= not(layer3_outputs(3902));
    layer4_outputs(1247) <= '0';
    layer4_outputs(1248) <= '1';
    layer4_outputs(1249) <= layer3_outputs(1558);
    layer4_outputs(1250) <= not(layer3_outputs(618));
    layer4_outputs(1251) <= (layer3_outputs(4041)) and not (layer3_outputs(3945));
    layer4_outputs(1252) <= layer3_outputs(4216);
    layer4_outputs(1253) <= not(layer3_outputs(2344));
    layer4_outputs(1254) <= not((layer3_outputs(3192)) or (layer3_outputs(4328)));
    layer4_outputs(1255) <= not(layer3_outputs(2139)) or (layer3_outputs(1772));
    layer4_outputs(1256) <= '1';
    layer4_outputs(1257) <= (layer3_outputs(590)) and not (layer3_outputs(1176));
    layer4_outputs(1258) <= (layer3_outputs(4721)) or (layer3_outputs(3319));
    layer4_outputs(1259) <= not(layer3_outputs(2767));
    layer4_outputs(1260) <= '1';
    layer4_outputs(1261) <= (layer3_outputs(3885)) and (layer3_outputs(1831));
    layer4_outputs(1262) <= layer3_outputs(4681);
    layer4_outputs(1263) <= not(layer3_outputs(2921));
    layer4_outputs(1264) <= layer3_outputs(4688);
    layer4_outputs(1265) <= layer3_outputs(2019);
    layer4_outputs(1266) <= layer3_outputs(4432);
    layer4_outputs(1267) <= not(layer3_outputs(4537));
    layer4_outputs(1268) <= not(layer3_outputs(1781)) or (layer3_outputs(454));
    layer4_outputs(1269) <= not(layer3_outputs(756));
    layer4_outputs(1270) <= '0';
    layer4_outputs(1271) <= not(layer3_outputs(4040));
    layer4_outputs(1272) <= not((layer3_outputs(3365)) xor (layer3_outputs(4796)));
    layer4_outputs(1273) <= layer3_outputs(2180);
    layer4_outputs(1274) <= not(layer3_outputs(1374));
    layer4_outputs(1275) <= not(layer3_outputs(2865));
    layer4_outputs(1276) <= not(layer3_outputs(991));
    layer4_outputs(1277) <= not((layer3_outputs(625)) and (layer3_outputs(1507)));
    layer4_outputs(1278) <= not(layer3_outputs(1844));
    layer4_outputs(1279) <= (layer3_outputs(319)) and not (layer3_outputs(2680));
    layer4_outputs(1280) <= not((layer3_outputs(3832)) xor (layer3_outputs(4605)));
    layer4_outputs(1281) <= '0';
    layer4_outputs(1282) <= not(layer3_outputs(372));
    layer4_outputs(1283) <= not(layer3_outputs(468)) or (layer3_outputs(2299));
    layer4_outputs(1284) <= layer3_outputs(3116);
    layer4_outputs(1285) <= not((layer3_outputs(3649)) and (layer3_outputs(424)));
    layer4_outputs(1286) <= layer3_outputs(3719);
    layer4_outputs(1287) <= layer3_outputs(3158);
    layer4_outputs(1288) <= not((layer3_outputs(1952)) or (layer3_outputs(3731)));
    layer4_outputs(1289) <= not(layer3_outputs(4720));
    layer4_outputs(1290) <= not(layer3_outputs(2355));
    layer4_outputs(1291) <= not(layer3_outputs(5024));
    layer4_outputs(1292) <= layer3_outputs(968);
    layer4_outputs(1293) <= layer3_outputs(1334);
    layer4_outputs(1294) <= not((layer3_outputs(2168)) or (layer3_outputs(798)));
    layer4_outputs(1295) <= not(layer3_outputs(453));
    layer4_outputs(1296) <= not(layer3_outputs(1276));
    layer4_outputs(1297) <= not((layer3_outputs(3078)) or (layer3_outputs(809)));
    layer4_outputs(1298) <= not(layer3_outputs(1270));
    layer4_outputs(1299) <= (layer3_outputs(1118)) and (layer3_outputs(4060));
    layer4_outputs(1300) <= not((layer3_outputs(1646)) xor (layer3_outputs(2465)));
    layer4_outputs(1301) <= '1';
    layer4_outputs(1302) <= not((layer3_outputs(3886)) or (layer3_outputs(1975)));
    layer4_outputs(1303) <= layer3_outputs(222);
    layer4_outputs(1304) <= not((layer3_outputs(489)) xor (layer3_outputs(3152)));
    layer4_outputs(1305) <= not((layer3_outputs(3178)) xor (layer3_outputs(2380)));
    layer4_outputs(1306) <= (layer3_outputs(2578)) and (layer3_outputs(4921));
    layer4_outputs(1307) <= not((layer3_outputs(2727)) or (layer3_outputs(1171)));
    layer4_outputs(1308) <= '0';
    layer4_outputs(1309) <= not(layer3_outputs(1267));
    layer4_outputs(1310) <= not(layer3_outputs(1765)) or (layer3_outputs(960));
    layer4_outputs(1311) <= (layer3_outputs(70)) and (layer3_outputs(4033));
    layer4_outputs(1312) <= '1';
    layer4_outputs(1313) <= '0';
    layer4_outputs(1314) <= not(layer3_outputs(290));
    layer4_outputs(1315) <= not(layer3_outputs(1716)) or (layer3_outputs(2330));
    layer4_outputs(1316) <= not(layer3_outputs(1419));
    layer4_outputs(1317) <= '0';
    layer4_outputs(1318) <= not(layer3_outputs(2120));
    layer4_outputs(1319) <= layer3_outputs(2644);
    layer4_outputs(1320) <= (layer3_outputs(69)) and not (layer3_outputs(1802));
    layer4_outputs(1321) <= (layer3_outputs(733)) and not (layer3_outputs(839));
    layer4_outputs(1322) <= not(layer3_outputs(798)) or (layer3_outputs(782));
    layer4_outputs(1323) <= layer3_outputs(995);
    layer4_outputs(1324) <= not(layer3_outputs(4800));
    layer4_outputs(1325) <= '0';
    layer4_outputs(1326) <= not(layer3_outputs(1659)) or (layer3_outputs(4629));
    layer4_outputs(1327) <= not(layer3_outputs(4458));
    layer4_outputs(1328) <= not(layer3_outputs(1946));
    layer4_outputs(1329) <= not(layer3_outputs(4999)) or (layer3_outputs(4735));
    layer4_outputs(1330) <= layer3_outputs(4901);
    layer4_outputs(1331) <= (layer3_outputs(3122)) and (layer3_outputs(72));
    layer4_outputs(1332) <= (layer3_outputs(145)) and not (layer3_outputs(1821));
    layer4_outputs(1333) <= not((layer3_outputs(3089)) or (layer3_outputs(4878)));
    layer4_outputs(1334) <= layer3_outputs(1476);
    layer4_outputs(1335) <= (layer3_outputs(5081)) and not (layer3_outputs(815));
    layer4_outputs(1336) <= '1';
    layer4_outputs(1337) <= not((layer3_outputs(2403)) or (layer3_outputs(359)));
    layer4_outputs(1338) <= not(layer3_outputs(4959));
    layer4_outputs(1339) <= not((layer3_outputs(842)) and (layer3_outputs(175)));
    layer4_outputs(1340) <= not(layer3_outputs(1805));
    layer4_outputs(1341) <= not(layer3_outputs(1044));
    layer4_outputs(1342) <= layer3_outputs(4718);
    layer4_outputs(1343) <= (layer3_outputs(1956)) or (layer3_outputs(2262));
    layer4_outputs(1344) <= layer3_outputs(3929);
    layer4_outputs(1345) <= not(layer3_outputs(1140));
    layer4_outputs(1346) <= layer3_outputs(1800);
    layer4_outputs(1347) <= (layer3_outputs(1733)) or (layer3_outputs(1962));
    layer4_outputs(1348) <= '1';
    layer4_outputs(1349) <= layer3_outputs(97);
    layer4_outputs(1350) <= layer3_outputs(4118);
    layer4_outputs(1351) <= '1';
    layer4_outputs(1352) <= layer3_outputs(2911);
    layer4_outputs(1353) <= layer3_outputs(4313);
    layer4_outputs(1354) <= layer3_outputs(4444);
    layer4_outputs(1355) <= not(layer3_outputs(4668));
    layer4_outputs(1356) <= '0';
    layer4_outputs(1357) <= layer3_outputs(1610);
    layer4_outputs(1358) <= not(layer3_outputs(2315));
    layer4_outputs(1359) <= layer3_outputs(4960);
    layer4_outputs(1360) <= layer3_outputs(443);
    layer4_outputs(1361) <= not(layer3_outputs(4181)) or (layer3_outputs(1025));
    layer4_outputs(1362) <= not(layer3_outputs(907));
    layer4_outputs(1363) <= not(layer3_outputs(4877));
    layer4_outputs(1364) <= (layer3_outputs(771)) and not (layer3_outputs(1577));
    layer4_outputs(1365) <= '0';
    layer4_outputs(1366) <= not(layer3_outputs(1686));
    layer4_outputs(1367) <= layer3_outputs(4146);
    layer4_outputs(1368) <= not((layer3_outputs(1506)) and (layer3_outputs(3530)));
    layer4_outputs(1369) <= '1';
    layer4_outputs(1370) <= (layer3_outputs(586)) and not (layer3_outputs(1880));
    layer4_outputs(1371) <= not(layer3_outputs(3336)) or (layer3_outputs(227));
    layer4_outputs(1372) <= (layer3_outputs(1415)) and (layer3_outputs(2917));
    layer4_outputs(1373) <= (layer3_outputs(2314)) or (layer3_outputs(4852));
    layer4_outputs(1374) <= (layer3_outputs(1625)) xor (layer3_outputs(497));
    layer4_outputs(1375) <= (layer3_outputs(3079)) xor (layer3_outputs(4002));
    layer4_outputs(1376) <= (layer3_outputs(13)) and not (layer3_outputs(1160));
    layer4_outputs(1377) <= (layer3_outputs(3388)) and not (layer3_outputs(1450));
    layer4_outputs(1378) <= '1';
    layer4_outputs(1379) <= not(layer3_outputs(4136)) or (layer3_outputs(4753));
    layer4_outputs(1380) <= not((layer3_outputs(1884)) or (layer3_outputs(1774)));
    layer4_outputs(1381) <= not((layer3_outputs(4583)) xor (layer3_outputs(2836)));
    layer4_outputs(1382) <= (layer3_outputs(787)) or (layer3_outputs(4233));
    layer4_outputs(1383) <= not(layer3_outputs(357));
    layer4_outputs(1384) <= not(layer3_outputs(1234));
    layer4_outputs(1385) <= (layer3_outputs(4418)) or (layer3_outputs(1053));
    layer4_outputs(1386) <= (layer3_outputs(2766)) and not (layer3_outputs(2110));
    layer4_outputs(1387) <= not(layer3_outputs(3391));
    layer4_outputs(1388) <= not((layer3_outputs(1049)) and (layer3_outputs(3180)));
    layer4_outputs(1389) <= not(layer3_outputs(2617));
    layer4_outputs(1390) <= '1';
    layer4_outputs(1391) <= (layer3_outputs(1024)) and (layer3_outputs(3031));
    layer4_outputs(1392) <= (layer3_outputs(3000)) and not (layer3_outputs(582));
    layer4_outputs(1393) <= (layer3_outputs(2695)) or (layer3_outputs(4356));
    layer4_outputs(1394) <= layer3_outputs(93);
    layer4_outputs(1395) <= layer3_outputs(1499);
    layer4_outputs(1396) <= (layer3_outputs(554)) and not (layer3_outputs(2744));
    layer4_outputs(1397) <= (layer3_outputs(4929)) and (layer3_outputs(4585));
    layer4_outputs(1398) <= not((layer3_outputs(3910)) xor (layer3_outputs(3319)));
    layer4_outputs(1399) <= (layer3_outputs(3831)) and not (layer3_outputs(1234));
    layer4_outputs(1400) <= not(layer3_outputs(5058)) or (layer3_outputs(3739));
    layer4_outputs(1401) <= layer3_outputs(2046);
    layer4_outputs(1402) <= (layer3_outputs(3604)) and (layer3_outputs(3773));
    layer4_outputs(1403) <= not(layer3_outputs(3401));
    layer4_outputs(1404) <= not(layer3_outputs(4514));
    layer4_outputs(1405) <= not((layer3_outputs(1428)) and (layer3_outputs(99)));
    layer4_outputs(1406) <= (layer3_outputs(3753)) xor (layer3_outputs(3937));
    layer4_outputs(1407) <= not(layer3_outputs(1921));
    layer4_outputs(1408) <= not(layer3_outputs(5054));
    layer4_outputs(1409) <= not((layer3_outputs(65)) xor (layer3_outputs(890)));
    layer4_outputs(1410) <= layer3_outputs(56);
    layer4_outputs(1411) <= (layer3_outputs(313)) and not (layer3_outputs(500));
    layer4_outputs(1412) <= not(layer3_outputs(1928)) or (layer3_outputs(966));
    layer4_outputs(1413) <= '1';
    layer4_outputs(1414) <= (layer3_outputs(1938)) xor (layer3_outputs(1280));
    layer4_outputs(1415) <= (layer3_outputs(2671)) and not (layer3_outputs(3852));
    layer4_outputs(1416) <= layer3_outputs(4143);
    layer4_outputs(1417) <= (layer3_outputs(1438)) xor (layer3_outputs(2023));
    layer4_outputs(1418) <= layer3_outputs(3987);
    layer4_outputs(1419) <= (layer3_outputs(0)) and not (layer3_outputs(2805));
    layer4_outputs(1420) <= not((layer3_outputs(779)) or (layer3_outputs(1707)));
    layer4_outputs(1421) <= not(layer3_outputs(3185));
    layer4_outputs(1422) <= not(layer3_outputs(4956));
    layer4_outputs(1423) <= (layer3_outputs(2807)) and not (layer3_outputs(2164));
    layer4_outputs(1424) <= not(layer3_outputs(1283));
    layer4_outputs(1425) <= not((layer3_outputs(580)) or (layer3_outputs(386)));
    layer4_outputs(1426) <= layer3_outputs(5081);
    layer4_outputs(1427) <= layer3_outputs(900);
    layer4_outputs(1428) <= not((layer3_outputs(2129)) xor (layer3_outputs(600)));
    layer4_outputs(1429) <= layer3_outputs(1252);
    layer4_outputs(1430) <= layer3_outputs(5040);
    layer4_outputs(1431) <= layer3_outputs(3095);
    layer4_outputs(1432) <= (layer3_outputs(2597)) xor (layer3_outputs(2948));
    layer4_outputs(1433) <= not(layer3_outputs(2476)) or (layer3_outputs(1790));
    layer4_outputs(1434) <= not(layer3_outputs(4817));
    layer4_outputs(1435) <= not(layer3_outputs(2887));
    layer4_outputs(1436) <= not(layer3_outputs(3600));
    layer4_outputs(1437) <= not(layer3_outputs(4849));
    layer4_outputs(1438) <= not(layer3_outputs(1477));
    layer4_outputs(1439) <= not(layer3_outputs(4848)) or (layer3_outputs(3217));
    layer4_outputs(1440) <= not((layer3_outputs(5093)) or (layer3_outputs(3943)));
    layer4_outputs(1441) <= not(layer3_outputs(4542));
    layer4_outputs(1442) <= (layer3_outputs(4922)) and not (layer3_outputs(3342));
    layer4_outputs(1443) <= not(layer3_outputs(1656));
    layer4_outputs(1444) <= layer3_outputs(2321);
    layer4_outputs(1445) <= (layer3_outputs(4925)) and not (layer3_outputs(2370));
    layer4_outputs(1446) <= layer3_outputs(4042);
    layer4_outputs(1447) <= layer3_outputs(197);
    layer4_outputs(1448) <= layer3_outputs(1996);
    layer4_outputs(1449) <= (layer3_outputs(2236)) or (layer3_outputs(4775));
    layer4_outputs(1450) <= '0';
    layer4_outputs(1451) <= (layer3_outputs(4793)) and not (layer3_outputs(8));
    layer4_outputs(1452) <= (layer3_outputs(3397)) and not (layer3_outputs(4544));
    layer4_outputs(1453) <= not((layer3_outputs(1376)) and (layer3_outputs(3894)));
    layer4_outputs(1454) <= '0';
    layer4_outputs(1455) <= (layer3_outputs(5020)) or (layer3_outputs(4865));
    layer4_outputs(1456) <= layer3_outputs(4491);
    layer4_outputs(1457) <= not(layer3_outputs(3979));
    layer4_outputs(1458) <= not(layer3_outputs(4140));
    layer4_outputs(1459) <= not(layer3_outputs(4246));
    layer4_outputs(1460) <= not(layer3_outputs(1469));
    layer4_outputs(1461) <= not((layer3_outputs(3792)) or (layer3_outputs(4724)));
    layer4_outputs(1462) <= not(layer3_outputs(1201));
    layer4_outputs(1463) <= not(layer3_outputs(2227));
    layer4_outputs(1464) <= not(layer3_outputs(1883));
    layer4_outputs(1465) <= not((layer3_outputs(5023)) and (layer3_outputs(1203)));
    layer4_outputs(1466) <= (layer3_outputs(2338)) and not (layer3_outputs(1338));
    layer4_outputs(1467) <= layer3_outputs(4780);
    layer4_outputs(1468) <= (layer3_outputs(3225)) xor (layer3_outputs(3230));
    layer4_outputs(1469) <= layer3_outputs(243);
    layer4_outputs(1470) <= not(layer3_outputs(1226));
    layer4_outputs(1471) <= not((layer3_outputs(2494)) xor (layer3_outputs(2120)));
    layer4_outputs(1472) <= layer3_outputs(2857);
    layer4_outputs(1473) <= not(layer3_outputs(3769));
    layer4_outputs(1474) <= layer3_outputs(4287);
    layer4_outputs(1475) <= layer3_outputs(4088);
    layer4_outputs(1476) <= not((layer3_outputs(3334)) and (layer3_outputs(503)));
    layer4_outputs(1477) <= '1';
    layer4_outputs(1478) <= not(layer3_outputs(1112)) or (layer3_outputs(517));
    layer4_outputs(1479) <= not(layer3_outputs(688));
    layer4_outputs(1480) <= not(layer3_outputs(379));
    layer4_outputs(1481) <= layer3_outputs(4389);
    layer4_outputs(1482) <= layer3_outputs(1915);
    layer4_outputs(1483) <= layer3_outputs(2883);
    layer4_outputs(1484) <= not(layer3_outputs(4804));
    layer4_outputs(1485) <= not(layer3_outputs(4014));
    layer4_outputs(1486) <= (layer3_outputs(4816)) or (layer3_outputs(4144));
    layer4_outputs(1487) <= (layer3_outputs(3036)) or (layer3_outputs(3640));
    layer4_outputs(1488) <= not(layer3_outputs(2473));
    layer4_outputs(1489) <= not(layer3_outputs(2741)) or (layer3_outputs(3724));
    layer4_outputs(1490) <= layer3_outputs(2488);
    layer4_outputs(1491) <= not(layer3_outputs(293));
    layer4_outputs(1492) <= layer3_outputs(4508);
    layer4_outputs(1493) <= layer3_outputs(2284);
    layer4_outputs(1494) <= not(layer3_outputs(3419));
    layer4_outputs(1495) <= not(layer3_outputs(2533));
    layer4_outputs(1496) <= not(layer3_outputs(5115)) or (layer3_outputs(1020));
    layer4_outputs(1497) <= (layer3_outputs(291)) and (layer3_outputs(4164));
    layer4_outputs(1498) <= not(layer3_outputs(475));
    layer4_outputs(1499) <= layer3_outputs(2765);
    layer4_outputs(1500) <= not((layer3_outputs(3045)) or (layer3_outputs(4205)));
    layer4_outputs(1501) <= not((layer3_outputs(3404)) xor (layer3_outputs(666)));
    layer4_outputs(1502) <= not(layer3_outputs(2134)) or (layer3_outputs(718));
    layer4_outputs(1503) <= not(layer3_outputs(3459));
    layer4_outputs(1504) <= layer3_outputs(791);
    layer4_outputs(1505) <= not((layer3_outputs(2997)) and (layer3_outputs(1653)));
    layer4_outputs(1506) <= (layer3_outputs(4947)) and not (layer3_outputs(2532));
    layer4_outputs(1507) <= layer3_outputs(3883);
    layer4_outputs(1508) <= layer3_outputs(4165);
    layer4_outputs(1509) <= layer3_outputs(4388);
    layer4_outputs(1510) <= (layer3_outputs(1850)) and not (layer3_outputs(4427));
    layer4_outputs(1511) <= not(layer3_outputs(950)) or (layer3_outputs(3073));
    layer4_outputs(1512) <= not(layer3_outputs(2754));
    layer4_outputs(1513) <= not((layer3_outputs(2820)) and (layer3_outputs(1292)));
    layer4_outputs(1514) <= not(layer3_outputs(4749));
    layer4_outputs(1515) <= (layer3_outputs(1458)) xor (layer3_outputs(3262));
    layer4_outputs(1516) <= '0';
    layer4_outputs(1517) <= not((layer3_outputs(1058)) and (layer3_outputs(780)));
    layer4_outputs(1518) <= not(layer3_outputs(188));
    layer4_outputs(1519) <= layer3_outputs(1372);
    layer4_outputs(1520) <= '1';
    layer4_outputs(1521) <= layer3_outputs(2361);
    layer4_outputs(1522) <= (layer3_outputs(40)) and not (layer3_outputs(680));
    layer4_outputs(1523) <= not(layer3_outputs(3398)) or (layer3_outputs(3927));
    layer4_outputs(1524) <= (layer3_outputs(1064)) and not (layer3_outputs(4139));
    layer4_outputs(1525) <= not((layer3_outputs(1060)) or (layer3_outputs(168)));
    layer4_outputs(1526) <= not((layer3_outputs(3018)) or (layer3_outputs(819)));
    layer4_outputs(1527) <= '1';
    layer4_outputs(1528) <= not(layer3_outputs(821));
    layer4_outputs(1529) <= '1';
    layer4_outputs(1530) <= not(layer3_outputs(3004)) or (layer3_outputs(4137));
    layer4_outputs(1531) <= layer3_outputs(30);
    layer4_outputs(1532) <= '1';
    layer4_outputs(1533) <= layer3_outputs(3024);
    layer4_outputs(1534) <= not(layer3_outputs(1019));
    layer4_outputs(1535) <= layer3_outputs(1657);
    layer4_outputs(1536) <= layer3_outputs(3651);
    layer4_outputs(1537) <= layer3_outputs(2173);
    layer4_outputs(1538) <= not((layer3_outputs(3942)) or (layer3_outputs(3974)));
    layer4_outputs(1539) <= layer3_outputs(4105);
    layer4_outputs(1540) <= not((layer3_outputs(2798)) and (layer3_outputs(3)));
    layer4_outputs(1541) <= (layer3_outputs(3165)) or (layer3_outputs(211));
    layer4_outputs(1542) <= '0';
    layer4_outputs(1543) <= (layer3_outputs(984)) and not (layer3_outputs(4629));
    layer4_outputs(1544) <= not(layer3_outputs(283)) or (layer3_outputs(2361));
    layer4_outputs(1545) <= layer3_outputs(1978);
    layer4_outputs(1546) <= '1';
    layer4_outputs(1547) <= not(layer3_outputs(2128));
    layer4_outputs(1548) <= layer3_outputs(3782);
    layer4_outputs(1549) <= not(layer3_outputs(909));
    layer4_outputs(1550) <= not((layer3_outputs(1108)) or (layer3_outputs(2307)));
    layer4_outputs(1551) <= '1';
    layer4_outputs(1552) <= not(layer3_outputs(4880));
    layer4_outputs(1553) <= layer3_outputs(3298);
    layer4_outputs(1554) <= '0';
    layer4_outputs(1555) <= (layer3_outputs(2075)) or (layer3_outputs(3619));
    layer4_outputs(1556) <= not(layer3_outputs(3644));
    layer4_outputs(1557) <= '1';
    layer4_outputs(1558) <= not((layer3_outputs(801)) or (layer3_outputs(2501)));
    layer4_outputs(1559) <= (layer3_outputs(847)) and not (layer3_outputs(2709));
    layer4_outputs(1560) <= not(layer3_outputs(3241));
    layer4_outputs(1561) <= not(layer3_outputs(2723)) or (layer3_outputs(3688));
    layer4_outputs(1562) <= (layer3_outputs(3499)) or (layer3_outputs(2999));
    layer4_outputs(1563) <= '1';
    layer4_outputs(1564) <= (layer3_outputs(3975)) or (layer3_outputs(2625));
    layer4_outputs(1565) <= not(layer3_outputs(214));
    layer4_outputs(1566) <= not(layer3_outputs(653));
    layer4_outputs(1567) <= (layer3_outputs(3980)) and not (layer3_outputs(2243));
    layer4_outputs(1568) <= (layer3_outputs(2223)) and not (layer3_outputs(3950));
    layer4_outputs(1569) <= not(layer3_outputs(504)) or (layer3_outputs(2034));
    layer4_outputs(1570) <= layer3_outputs(699);
    layer4_outputs(1571) <= (layer3_outputs(2970)) or (layer3_outputs(1167));
    layer4_outputs(1572) <= layer3_outputs(2568);
    layer4_outputs(1573) <= '0';
    layer4_outputs(1574) <= '1';
    layer4_outputs(1575) <= not((layer3_outputs(3895)) and (layer3_outputs(784)));
    layer4_outputs(1576) <= (layer3_outputs(4146)) and not (layer3_outputs(4363));
    layer4_outputs(1577) <= not(layer3_outputs(723)) or (layer3_outputs(3187));
    layer4_outputs(1578) <= not(layer3_outputs(3322));
    layer4_outputs(1579) <= layer3_outputs(3655);
    layer4_outputs(1580) <= not(layer3_outputs(5029));
    layer4_outputs(1581) <= not(layer3_outputs(3516)) or (layer3_outputs(3214));
    layer4_outputs(1582) <= (layer3_outputs(3186)) and (layer3_outputs(1573));
    layer4_outputs(1583) <= '0';
    layer4_outputs(1584) <= not(layer3_outputs(3897)) or (layer3_outputs(1615));
    layer4_outputs(1585) <= layer3_outputs(3444);
    layer4_outputs(1586) <= not(layer3_outputs(5040)) or (layer3_outputs(3169));
    layer4_outputs(1587) <= not(layer3_outputs(2912)) or (layer3_outputs(423));
    layer4_outputs(1588) <= not(layer3_outputs(176)) or (layer3_outputs(4844));
    layer4_outputs(1589) <= not((layer3_outputs(588)) xor (layer3_outputs(3893)));
    layer4_outputs(1590) <= not(layer3_outputs(3588));
    layer4_outputs(1591) <= layer3_outputs(235);
    layer4_outputs(1592) <= layer3_outputs(4883);
    layer4_outputs(1593) <= layer3_outputs(4293);
    layer4_outputs(1594) <= not(layer3_outputs(1362)) or (layer3_outputs(4541));
    layer4_outputs(1595) <= not((layer3_outputs(3207)) or (layer3_outputs(3517)));
    layer4_outputs(1596) <= layer3_outputs(3726);
    layer4_outputs(1597) <= not(layer3_outputs(667)) or (layer3_outputs(3099));
    layer4_outputs(1598) <= layer3_outputs(36);
    layer4_outputs(1599) <= (layer3_outputs(2205)) or (layer3_outputs(228));
    layer4_outputs(1600) <= layer3_outputs(3510);
    layer4_outputs(1601) <= (layer3_outputs(2060)) xor (layer3_outputs(4092));
    layer4_outputs(1602) <= not((layer3_outputs(4870)) and (layer3_outputs(730)));
    layer4_outputs(1603) <= not(layer3_outputs(2844));
    layer4_outputs(1604) <= (layer3_outputs(4418)) and not (layer3_outputs(3068));
    layer4_outputs(1605) <= not(layer3_outputs(5039));
    layer4_outputs(1606) <= layer3_outputs(2410);
    layer4_outputs(1607) <= not((layer3_outputs(436)) xor (layer3_outputs(464)));
    layer4_outputs(1608) <= layer3_outputs(1768);
    layer4_outputs(1609) <= not(layer3_outputs(34)) or (layer3_outputs(4016));
    layer4_outputs(1610) <= not((layer3_outputs(3832)) xor (layer3_outputs(5068)));
    layer4_outputs(1611) <= (layer3_outputs(897)) and (layer3_outputs(1730));
    layer4_outputs(1612) <= '0';
    layer4_outputs(1613) <= (layer3_outputs(1337)) and (layer3_outputs(1405));
    layer4_outputs(1614) <= (layer3_outputs(3891)) or (layer3_outputs(651));
    layer4_outputs(1615) <= (layer3_outputs(1229)) and not (layer3_outputs(4968));
    layer4_outputs(1616) <= not((layer3_outputs(3463)) and (layer3_outputs(3450)));
    layer4_outputs(1617) <= (layer3_outputs(4895)) and not (layer3_outputs(1773));
    layer4_outputs(1618) <= '0';
    layer4_outputs(1619) <= not(layer3_outputs(4636));
    layer4_outputs(1620) <= (layer3_outputs(4915)) xor (layer3_outputs(856));
    layer4_outputs(1621) <= (layer3_outputs(4711)) and (layer3_outputs(1858));
    layer4_outputs(1622) <= not(layer3_outputs(5106));
    layer4_outputs(1623) <= not(layer3_outputs(1259));
    layer4_outputs(1624) <= not((layer3_outputs(4036)) and (layer3_outputs(12)));
    layer4_outputs(1625) <= layer3_outputs(5003);
    layer4_outputs(1626) <= not((layer3_outputs(84)) and (layer3_outputs(42)));
    layer4_outputs(1627) <= '1';
    layer4_outputs(1628) <= '1';
    layer4_outputs(1629) <= layer3_outputs(1767);
    layer4_outputs(1630) <= not(layer3_outputs(3168)) or (layer3_outputs(3863));
    layer4_outputs(1631) <= (layer3_outputs(3991)) and (layer3_outputs(3164));
    layer4_outputs(1632) <= not((layer3_outputs(3344)) and (layer3_outputs(26)));
    layer4_outputs(1633) <= (layer3_outputs(2972)) or (layer3_outputs(1593));
    layer4_outputs(1634) <= (layer3_outputs(2760)) and not (layer3_outputs(1192));
    layer4_outputs(1635) <= layer3_outputs(1059);
    layer4_outputs(1636) <= not((layer3_outputs(1105)) and (layer3_outputs(2945)));
    layer4_outputs(1637) <= not(layer3_outputs(2151));
    layer4_outputs(1638) <= not((layer3_outputs(4011)) and (layer3_outputs(2091)));
    layer4_outputs(1639) <= not((layer3_outputs(1795)) or (layer3_outputs(68)));
    layer4_outputs(1640) <= (layer3_outputs(2678)) or (layer3_outputs(2925));
    layer4_outputs(1641) <= not((layer3_outputs(4893)) and (layer3_outputs(1547)));
    layer4_outputs(1642) <= not(layer3_outputs(2033)) or (layer3_outputs(1839));
    layer4_outputs(1643) <= not(layer3_outputs(3910));
    layer4_outputs(1644) <= not(layer3_outputs(2145));
    layer4_outputs(1645) <= (layer3_outputs(4837)) or (layer3_outputs(4813));
    layer4_outputs(1646) <= not((layer3_outputs(4862)) xor (layer3_outputs(4293)));
    layer4_outputs(1647) <= not(layer3_outputs(2252));
    layer4_outputs(1648) <= (layer3_outputs(2497)) and not (layer3_outputs(2873));
    layer4_outputs(1649) <= not(layer3_outputs(2824)) or (layer3_outputs(2217));
    layer4_outputs(1650) <= not((layer3_outputs(976)) and (layer3_outputs(2267)));
    layer4_outputs(1651) <= layer3_outputs(1208);
    layer4_outputs(1652) <= not(layer3_outputs(835)) or (layer3_outputs(489));
    layer4_outputs(1653) <= (layer3_outputs(4289)) and not (layer3_outputs(4637));
    layer4_outputs(1654) <= (layer3_outputs(3523)) or (layer3_outputs(4381));
    layer4_outputs(1655) <= not((layer3_outputs(3914)) and (layer3_outputs(473)));
    layer4_outputs(1656) <= layer3_outputs(1056);
    layer4_outputs(1657) <= layer3_outputs(2632);
    layer4_outputs(1658) <= not((layer3_outputs(4803)) and (layer3_outputs(1971)));
    layer4_outputs(1659) <= not(layer3_outputs(3261)) or (layer3_outputs(4307));
    layer4_outputs(1660) <= (layer3_outputs(2402)) and not (layer3_outputs(2906));
    layer4_outputs(1661) <= (layer3_outputs(3109)) and not (layer3_outputs(412));
    layer4_outputs(1662) <= layer3_outputs(1584);
    layer4_outputs(1663) <= not(layer3_outputs(782));
    layer4_outputs(1664) <= (layer3_outputs(4920)) or (layer3_outputs(1083));
    layer4_outputs(1665) <= not((layer3_outputs(5043)) or (layer3_outputs(860)));
    layer4_outputs(1666) <= (layer3_outputs(883)) or (layer3_outputs(1297));
    layer4_outputs(1667) <= not(layer3_outputs(908)) or (layer3_outputs(3940));
    layer4_outputs(1668) <= '0';
    layer4_outputs(1669) <= (layer3_outputs(2899)) xor (layer3_outputs(3706));
    layer4_outputs(1670) <= (layer3_outputs(952)) and not (layer3_outputs(3898));
    layer4_outputs(1671) <= (layer3_outputs(2706)) and not (layer3_outputs(550));
    layer4_outputs(1672) <= layer3_outputs(3663);
    layer4_outputs(1673) <= not(layer3_outputs(4533));
    layer4_outputs(1674) <= not(layer3_outputs(4895)) or (layer3_outputs(185));
    layer4_outputs(1675) <= layer3_outputs(1753);
    layer4_outputs(1676) <= (layer3_outputs(265)) and not (layer3_outputs(4395));
    layer4_outputs(1677) <= layer3_outputs(314);
    layer4_outputs(1678) <= layer3_outputs(3811);
    layer4_outputs(1679) <= not(layer3_outputs(953));
    layer4_outputs(1680) <= layer3_outputs(1083);
    layer4_outputs(1681) <= (layer3_outputs(2256)) and (layer3_outputs(2738));
    layer4_outputs(1682) <= layer3_outputs(3678);
    layer4_outputs(1683) <= not(layer3_outputs(3219));
    layer4_outputs(1684) <= not(layer3_outputs(2394));
    layer4_outputs(1685) <= (layer3_outputs(2194)) and not (layer3_outputs(4085));
    layer4_outputs(1686) <= not(layer3_outputs(4168));
    layer4_outputs(1687) <= (layer3_outputs(74)) and not (layer3_outputs(5009));
    layer4_outputs(1688) <= (layer3_outputs(1708)) or (layer3_outputs(3227));
    layer4_outputs(1689) <= not(layer3_outputs(4210));
    layer4_outputs(1690) <= layer3_outputs(683);
    layer4_outputs(1691) <= not((layer3_outputs(741)) and (layer3_outputs(2390)));
    layer4_outputs(1692) <= '0';
    layer4_outputs(1693) <= (layer3_outputs(142)) and not (layer3_outputs(1601));
    layer4_outputs(1694) <= not(layer3_outputs(2634));
    layer4_outputs(1695) <= layer3_outputs(3090);
    layer4_outputs(1696) <= layer3_outputs(2142);
    layer4_outputs(1697) <= not((layer3_outputs(4860)) xor (layer3_outputs(1918)));
    layer4_outputs(1698) <= not(layer3_outputs(2612));
    layer4_outputs(1699) <= layer3_outputs(1140);
    layer4_outputs(1700) <= not(layer3_outputs(1731));
    layer4_outputs(1701) <= layer3_outputs(86);
    layer4_outputs(1702) <= not(layer3_outputs(3867));
    layer4_outputs(1703) <= not(layer3_outputs(1959));
    layer4_outputs(1704) <= not(layer3_outputs(4690));
    layer4_outputs(1705) <= not(layer3_outputs(2519)) or (layer3_outputs(1657));
    layer4_outputs(1706) <= not((layer3_outputs(221)) or (layer3_outputs(4149)));
    layer4_outputs(1707) <= not((layer3_outputs(1910)) and (layer3_outputs(406)));
    layer4_outputs(1708) <= not(layer3_outputs(685));
    layer4_outputs(1709) <= layer3_outputs(2940);
    layer4_outputs(1710) <= layer3_outputs(4858);
    layer4_outputs(1711) <= (layer3_outputs(2632)) and (layer3_outputs(1729));
    layer4_outputs(1712) <= '1';
    layer4_outputs(1713) <= layer3_outputs(4260);
    layer4_outputs(1714) <= not((layer3_outputs(534)) and (layer3_outputs(11)));
    layer4_outputs(1715) <= layer3_outputs(2549);
    layer4_outputs(1716) <= layer3_outputs(2108);
    layer4_outputs(1717) <= not((layer3_outputs(3576)) or (layer3_outputs(4085)));
    layer4_outputs(1718) <= not(layer3_outputs(51));
    layer4_outputs(1719) <= not(layer3_outputs(4452));
    layer4_outputs(1720) <= '1';
    layer4_outputs(1721) <= not((layer3_outputs(4481)) and (layer3_outputs(1607)));
    layer4_outputs(1722) <= not(layer3_outputs(4197));
    layer4_outputs(1723) <= '1';
    layer4_outputs(1724) <= not(layer3_outputs(676));
    layer4_outputs(1725) <= not((layer3_outputs(4576)) and (layer3_outputs(1127)));
    layer4_outputs(1726) <= (layer3_outputs(4091)) and not (layer3_outputs(1673));
    layer4_outputs(1727) <= not((layer3_outputs(2859)) and (layer3_outputs(3491)));
    layer4_outputs(1728) <= not((layer3_outputs(2507)) or (layer3_outputs(4563)));
    layer4_outputs(1729) <= '1';
    layer4_outputs(1730) <= not((layer3_outputs(1193)) and (layer3_outputs(4077)));
    layer4_outputs(1731) <= not(layer3_outputs(3861));
    layer4_outputs(1732) <= '0';
    layer4_outputs(1733) <= (layer3_outputs(62)) and not (layer3_outputs(1812));
    layer4_outputs(1734) <= not(layer3_outputs(4334)) or (layer3_outputs(4776));
    layer4_outputs(1735) <= (layer3_outputs(5049)) or (layer3_outputs(1445));
    layer4_outputs(1736) <= (layer3_outputs(3196)) and (layer3_outputs(631));
    layer4_outputs(1737) <= layer3_outputs(2772);
    layer4_outputs(1738) <= (layer3_outputs(4899)) or (layer3_outputs(1483));
    layer4_outputs(1739) <= not(layer3_outputs(1177)) or (layer3_outputs(4240));
    layer4_outputs(1740) <= not((layer3_outputs(2920)) or (layer3_outputs(4292)));
    layer4_outputs(1741) <= (layer3_outputs(2302)) and not (layer3_outputs(488));
    layer4_outputs(1742) <= layer3_outputs(4886);
    layer4_outputs(1743) <= not(layer3_outputs(3269));
    layer4_outputs(1744) <= '0';
    layer4_outputs(1745) <= (layer3_outputs(2338)) and (layer3_outputs(4589));
    layer4_outputs(1746) <= not(layer3_outputs(4934));
    layer4_outputs(1747) <= layer3_outputs(3823);
    layer4_outputs(1748) <= not(layer3_outputs(2616));
    layer4_outputs(1749) <= not(layer3_outputs(2766)) or (layer3_outputs(3849));
    layer4_outputs(1750) <= not((layer3_outputs(1689)) or (layer3_outputs(612)));
    layer4_outputs(1751) <= not(layer3_outputs(1618));
    layer4_outputs(1752) <= not(layer3_outputs(1311)) or (layer3_outputs(1368));
    layer4_outputs(1753) <= (layer3_outputs(4157)) and (layer3_outputs(2773));
    layer4_outputs(1754) <= layer3_outputs(772);
    layer4_outputs(1755) <= layer3_outputs(4750);
    layer4_outputs(1756) <= not(layer3_outputs(805));
    layer4_outputs(1757) <= (layer3_outputs(2636)) and (layer3_outputs(4857));
    layer4_outputs(1758) <= layer3_outputs(1688);
    layer4_outputs(1759) <= layer3_outputs(1924);
    layer4_outputs(1760) <= not(layer3_outputs(980)) or (layer3_outputs(3713));
    layer4_outputs(1761) <= layer3_outputs(4256);
    layer4_outputs(1762) <= not(layer3_outputs(2680));
    layer4_outputs(1763) <= not(layer3_outputs(4677));
    layer4_outputs(1764) <= '1';
    layer4_outputs(1765) <= (layer3_outputs(3495)) and (layer3_outputs(638));
    layer4_outputs(1766) <= not(layer3_outputs(5039)) or (layer3_outputs(1602));
    layer4_outputs(1767) <= not(layer3_outputs(4974));
    layer4_outputs(1768) <= '1';
    layer4_outputs(1769) <= layer3_outputs(4385);
    layer4_outputs(1770) <= layer3_outputs(4281);
    layer4_outputs(1771) <= not(layer3_outputs(138));
    layer4_outputs(1772) <= not((layer3_outputs(2863)) xor (layer3_outputs(1582)));
    layer4_outputs(1773) <= not((layer3_outputs(343)) and (layer3_outputs(4023)));
    layer4_outputs(1774) <= not(layer3_outputs(4632));
    layer4_outputs(1775) <= not((layer3_outputs(4718)) and (layer3_outputs(3084)));
    layer4_outputs(1776) <= not((layer3_outputs(1215)) and (layer3_outputs(1642)));
    layer4_outputs(1777) <= not(layer3_outputs(4484)) or (layer3_outputs(4888));
    layer4_outputs(1778) <= '0';
    layer4_outputs(1779) <= layer3_outputs(2681);
    layer4_outputs(1780) <= not((layer3_outputs(668)) and (layer3_outputs(2181)));
    layer4_outputs(1781) <= not(layer3_outputs(420));
    layer4_outputs(1782) <= (layer3_outputs(590)) and not (layer3_outputs(4661));
    layer4_outputs(1783) <= not(layer3_outputs(2550));
    layer4_outputs(1784) <= not(layer3_outputs(3385)) or (layer3_outputs(2603));
    layer4_outputs(1785) <= layer3_outputs(729);
    layer4_outputs(1786) <= layer3_outputs(1195);
    layer4_outputs(1787) <= not(layer3_outputs(1620)) or (layer3_outputs(5044));
    layer4_outputs(1788) <= '0';
    layer4_outputs(1789) <= (layer3_outputs(4714)) and not (layer3_outputs(2984));
    layer4_outputs(1790) <= layer3_outputs(3301);
    layer4_outputs(1791) <= not(layer3_outputs(4578)) or (layer3_outputs(496));
    layer4_outputs(1792) <= not(layer3_outputs(301));
    layer4_outputs(1793) <= layer3_outputs(3174);
    layer4_outputs(1794) <= (layer3_outputs(4421)) and not (layer3_outputs(2930));
    layer4_outputs(1795) <= layer3_outputs(4936);
    layer4_outputs(1796) <= not(layer3_outputs(1977));
    layer4_outputs(1797) <= layer3_outputs(1963);
    layer4_outputs(1798) <= (layer3_outputs(4342)) and not (layer3_outputs(4160));
    layer4_outputs(1799) <= (layer3_outputs(1522)) and (layer3_outputs(854));
    layer4_outputs(1800) <= '1';
    layer4_outputs(1801) <= layer3_outputs(1497);
    layer4_outputs(1802) <= '0';
    layer4_outputs(1803) <= layer3_outputs(1818);
    layer4_outputs(1804) <= not(layer3_outputs(2775));
    layer4_outputs(1805) <= not((layer3_outputs(1845)) and (layer3_outputs(2576)));
    layer4_outputs(1806) <= (layer3_outputs(3591)) or (layer3_outputs(4272));
    layer4_outputs(1807) <= not(layer3_outputs(4396));
    layer4_outputs(1808) <= layer3_outputs(4828);
    layer4_outputs(1809) <= layer3_outputs(393);
    layer4_outputs(1810) <= not((layer3_outputs(1359)) xor (layer3_outputs(738)));
    layer4_outputs(1811) <= not((layer3_outputs(4559)) and (layer3_outputs(3584)));
    layer4_outputs(1812) <= layer3_outputs(3630);
    layer4_outputs(1813) <= not(layer3_outputs(1782));
    layer4_outputs(1814) <= (layer3_outputs(81)) or (layer3_outputs(1983));
    layer4_outputs(1815) <= layer3_outputs(1911);
    layer4_outputs(1816) <= layer3_outputs(1449);
    layer4_outputs(1817) <= not((layer3_outputs(945)) and (layer3_outputs(2579)));
    layer4_outputs(1818) <= layer3_outputs(3560);
    layer4_outputs(1819) <= not(layer3_outputs(736)) or (layer3_outputs(2720));
    layer4_outputs(1820) <= layer3_outputs(1988);
    layer4_outputs(1821) <= '0';
    layer4_outputs(1822) <= not(layer3_outputs(157));
    layer4_outputs(1823) <= (layer3_outputs(1142)) and not (layer3_outputs(1139));
    layer4_outputs(1824) <= (layer3_outputs(4055)) and not (layer3_outputs(571));
    layer4_outputs(1825) <= (layer3_outputs(174)) xor (layer3_outputs(3126));
    layer4_outputs(1826) <= (layer3_outputs(315)) and (layer3_outputs(4738));
    layer4_outputs(1827) <= not((layer3_outputs(493)) or (layer3_outputs(3994)));
    layer4_outputs(1828) <= not(layer3_outputs(2396));
    layer4_outputs(1829) <= layer3_outputs(4674);
    layer4_outputs(1830) <= (layer3_outputs(2054)) and not (layer3_outputs(2253));
    layer4_outputs(1831) <= not((layer3_outputs(2537)) or (layer3_outputs(389)));
    layer4_outputs(1832) <= not(layer3_outputs(2202)) or (layer3_outputs(2424));
    layer4_outputs(1833) <= not(layer3_outputs(486));
    layer4_outputs(1834) <= not((layer3_outputs(2193)) xor (layer3_outputs(2165)));
    layer4_outputs(1835) <= not((layer3_outputs(1491)) and (layer3_outputs(3687)));
    layer4_outputs(1836) <= not((layer3_outputs(606)) or (layer3_outputs(1571)));
    layer4_outputs(1837) <= '1';
    layer4_outputs(1838) <= (layer3_outputs(537)) and (layer3_outputs(4428));
    layer4_outputs(1839) <= not(layer3_outputs(1612)) or (layer3_outputs(1802));
    layer4_outputs(1840) <= (layer3_outputs(753)) or (layer3_outputs(723));
    layer4_outputs(1841) <= '1';
    layer4_outputs(1842) <= layer3_outputs(521);
    layer4_outputs(1843) <= '0';
    layer4_outputs(1844) <= layer3_outputs(4185);
    layer4_outputs(1845) <= (layer3_outputs(2251)) or (layer3_outputs(2893));
    layer4_outputs(1846) <= not(layer3_outputs(92)) or (layer3_outputs(4038));
    layer4_outputs(1847) <= not((layer3_outputs(3446)) and (layer3_outputs(2540)));
    layer4_outputs(1848) <= '1';
    layer4_outputs(1849) <= not((layer3_outputs(2613)) and (layer3_outputs(3183)));
    layer4_outputs(1850) <= (layer3_outputs(3922)) and not (layer3_outputs(1404));
    layer4_outputs(1851) <= (layer3_outputs(3553)) and not (layer3_outputs(2140));
    layer4_outputs(1852) <= not(layer3_outputs(2264));
    layer4_outputs(1853) <= (layer3_outputs(2364)) and not (layer3_outputs(3785));
    layer4_outputs(1854) <= layer3_outputs(3139);
    layer4_outputs(1855) <= '0';
    layer4_outputs(1856) <= not(layer3_outputs(1631)) or (layer3_outputs(1720));
    layer4_outputs(1857) <= not(layer3_outputs(3178)) or (layer3_outputs(1534));
    layer4_outputs(1858) <= (layer3_outputs(304)) and not (layer3_outputs(5093));
    layer4_outputs(1859) <= (layer3_outputs(4506)) and (layer3_outputs(528));
    layer4_outputs(1860) <= '0';
    layer4_outputs(1861) <= (layer3_outputs(987)) and not (layer3_outputs(2303));
    layer4_outputs(1862) <= layer3_outputs(1457);
    layer4_outputs(1863) <= (layer3_outputs(259)) and (layer3_outputs(992));
    layer4_outputs(1864) <= '0';
    layer4_outputs(1865) <= not(layer3_outputs(885));
    layer4_outputs(1866) <= (layer3_outputs(2729)) and not (layer3_outputs(4473));
    layer4_outputs(1867) <= not((layer3_outputs(3635)) and (layer3_outputs(3320)));
    layer4_outputs(1868) <= (layer3_outputs(3310)) or (layer3_outputs(3638));
    layer4_outputs(1869) <= not(layer3_outputs(3078));
    layer4_outputs(1870) <= not(layer3_outputs(2152));
    layer4_outputs(1871) <= layer3_outputs(3703);
    layer4_outputs(1872) <= layer3_outputs(2343);
    layer4_outputs(1873) <= '1';
    layer4_outputs(1874) <= not((layer3_outputs(286)) and (layer3_outputs(3234)));
    layer4_outputs(1875) <= layer3_outputs(3626);
    layer4_outputs(1876) <= not(layer3_outputs(2931));
    layer4_outputs(1877) <= (layer3_outputs(358)) and (layer3_outputs(5044));
    layer4_outputs(1878) <= layer3_outputs(647);
    layer4_outputs(1879) <= (layer3_outputs(748)) or (layer3_outputs(1478));
    layer4_outputs(1880) <= not((layer3_outputs(2031)) and (layer3_outputs(4511)));
    layer4_outputs(1881) <= (layer3_outputs(151)) xor (layer3_outputs(4304));
    layer4_outputs(1882) <= layer3_outputs(3119);
    layer4_outputs(1883) <= not(layer3_outputs(838));
    layer4_outputs(1884) <= layer3_outputs(4388);
    layer4_outputs(1885) <= (layer3_outputs(1664)) and not (layer3_outputs(3793));
    layer4_outputs(1886) <= (layer3_outputs(2109)) and not (layer3_outputs(2539));
    layer4_outputs(1887) <= (layer3_outputs(2687)) and not (layer3_outputs(4210));
    layer4_outputs(1888) <= not((layer3_outputs(3131)) and (layer3_outputs(3967)));
    layer4_outputs(1889) <= not(layer3_outputs(3073));
    layer4_outputs(1890) <= not(layer3_outputs(2613));
    layer4_outputs(1891) <= (layer3_outputs(4091)) and not (layer3_outputs(103));
    layer4_outputs(1892) <= not(layer3_outputs(1607)) or (layer3_outputs(1109));
    layer4_outputs(1893) <= not(layer3_outputs(4185));
    layer4_outputs(1894) <= (layer3_outputs(3523)) and (layer3_outputs(1339));
    layer4_outputs(1895) <= not(layer3_outputs(262)) or (layer3_outputs(1302));
    layer4_outputs(1896) <= layer3_outputs(1698);
    layer4_outputs(1897) <= '0';
    layer4_outputs(1898) <= not(layer3_outputs(4741));
    layer4_outputs(1899) <= layer3_outputs(1501);
    layer4_outputs(1900) <= not(layer3_outputs(1384));
    layer4_outputs(1901) <= not((layer3_outputs(2234)) and (layer3_outputs(3783)));
    layer4_outputs(1902) <= not(layer3_outputs(604));
    layer4_outputs(1903) <= not((layer3_outputs(2324)) and (layer3_outputs(4321)));
    layer4_outputs(1904) <= '1';
    layer4_outputs(1905) <= layer3_outputs(3541);
    layer4_outputs(1906) <= not((layer3_outputs(4465)) or (layer3_outputs(3702)));
    layer4_outputs(1907) <= '1';
    layer4_outputs(1908) <= not((layer3_outputs(31)) and (layer3_outputs(2721)));
    layer4_outputs(1909) <= not(layer3_outputs(1304));
    layer4_outputs(1910) <= (layer3_outputs(1014)) xor (layer3_outputs(635));
    layer4_outputs(1911) <= '1';
    layer4_outputs(1912) <= layer3_outputs(5008);
    layer4_outputs(1913) <= not((layer3_outputs(4726)) or (layer3_outputs(2261)));
    layer4_outputs(1914) <= '0';
    layer4_outputs(1915) <= not(layer3_outputs(3997));
    layer4_outputs(1916) <= '0';
    layer4_outputs(1917) <= not(layer3_outputs(3952)) or (layer3_outputs(1784));
    layer4_outputs(1918) <= not(layer3_outputs(1922)) or (layer3_outputs(3086));
    layer4_outputs(1919) <= not(layer3_outputs(1166)) or (layer3_outputs(1263));
    layer4_outputs(1920) <= not((layer3_outputs(914)) or (layer3_outputs(748)));
    layer4_outputs(1921) <= not((layer3_outputs(4383)) xor (layer3_outputs(948)));
    layer4_outputs(1922) <= not((layer3_outputs(811)) and (layer3_outputs(21)));
    layer4_outputs(1923) <= not(layer3_outputs(3283)) or (layer3_outputs(4060));
    layer4_outputs(1924) <= '0';
    layer4_outputs(1925) <= (layer3_outputs(4539)) xor (layer3_outputs(4962));
    layer4_outputs(1926) <= layer3_outputs(1455);
    layer4_outputs(1927) <= (layer3_outputs(1435)) and not (layer3_outputs(1798));
    layer4_outputs(1928) <= not(layer3_outputs(383));
    layer4_outputs(1929) <= '1';
    layer4_outputs(1930) <= layer3_outputs(4314);
    layer4_outputs(1931) <= not(layer3_outputs(660));
    layer4_outputs(1932) <= '0';
    layer4_outputs(1933) <= (layer3_outputs(4079)) and not (layer3_outputs(2026));
    layer4_outputs(1934) <= '1';
    layer4_outputs(1935) <= (layer3_outputs(3312)) and (layer3_outputs(3221));
    layer4_outputs(1936) <= not(layer3_outputs(581));
    layer4_outputs(1937) <= (layer3_outputs(4247)) and not (layer3_outputs(3141));
    layer4_outputs(1938) <= not(layer3_outputs(2862));
    layer4_outputs(1939) <= layer3_outputs(2843);
    layer4_outputs(1940) <= (layer3_outputs(1442)) or (layer3_outputs(1583));
    layer4_outputs(1941) <= '1';
    layer4_outputs(1942) <= layer3_outputs(2438);
    layer4_outputs(1943) <= not(layer3_outputs(2643)) or (layer3_outputs(4540));
    layer4_outputs(1944) <= layer3_outputs(4806);
    layer4_outputs(1945) <= not(layer3_outputs(1523));
    layer4_outputs(1946) <= not((layer3_outputs(3279)) and (layer3_outputs(3857)));
    layer4_outputs(1947) <= not(layer3_outputs(2649));
    layer4_outputs(1948) <= (layer3_outputs(2428)) and (layer3_outputs(4786));
    layer4_outputs(1949) <= layer3_outputs(3099);
    layer4_outputs(1950) <= (layer3_outputs(3804)) and not (layer3_outputs(3959));
    layer4_outputs(1951) <= (layer3_outputs(4530)) or (layer3_outputs(1935));
    layer4_outputs(1952) <= layer3_outputs(4347);
    layer4_outputs(1953) <= (layer3_outputs(3866)) and not (layer3_outputs(2683));
    layer4_outputs(1954) <= layer3_outputs(3103);
    layer4_outputs(1955) <= (layer3_outputs(1890)) and not (layer3_outputs(4540));
    layer4_outputs(1956) <= not((layer3_outputs(3689)) and (layer3_outputs(385)));
    layer4_outputs(1957) <= '1';
    layer4_outputs(1958) <= not((layer3_outputs(971)) and (layer3_outputs(3294)));
    layer4_outputs(1959) <= (layer3_outputs(978)) xor (layer3_outputs(4800));
    layer4_outputs(1960) <= layer3_outputs(2105);
    layer4_outputs(1961) <= layer3_outputs(3864);
    layer4_outputs(1962) <= '0';
    layer4_outputs(1963) <= not(layer3_outputs(1633));
    layer4_outputs(1964) <= (layer3_outputs(490)) xor (layer3_outputs(3852));
    layer4_outputs(1965) <= layer3_outputs(3882);
    layer4_outputs(1966) <= not(layer3_outputs(366));
    layer4_outputs(1967) <= not((layer3_outputs(1365)) and (layer3_outputs(467)));
    layer4_outputs(1968) <= (layer3_outputs(566)) and (layer3_outputs(1426));
    layer4_outputs(1969) <= (layer3_outputs(3849)) and not (layer3_outputs(4196));
    layer4_outputs(1970) <= not(layer3_outputs(3588)) or (layer3_outputs(2601));
    layer4_outputs(1971) <= '0';
    layer4_outputs(1972) <= layer3_outputs(681);
    layer4_outputs(1973) <= layer3_outputs(3034);
    layer4_outputs(1974) <= (layer3_outputs(4818)) and not (layer3_outputs(1595));
    layer4_outputs(1975) <= layer3_outputs(5117);
    layer4_outputs(1976) <= not(layer3_outputs(4441));
    layer4_outputs(1977) <= '0';
    layer4_outputs(1978) <= '0';
    layer4_outputs(1979) <= (layer3_outputs(3690)) and not (layer3_outputs(3101));
    layer4_outputs(1980) <= not((layer3_outputs(4155)) or (layer3_outputs(5011)));
    layer4_outputs(1981) <= layer3_outputs(2675);
    layer4_outputs(1982) <= '1';
    layer4_outputs(1983) <= not(layer3_outputs(300)) or (layer3_outputs(4549));
    layer4_outputs(1984) <= not(layer3_outputs(4673));
    layer4_outputs(1985) <= (layer3_outputs(3996)) and not (layer3_outputs(2926));
    layer4_outputs(1986) <= not(layer3_outputs(2018));
    layer4_outputs(1987) <= '1';
    layer4_outputs(1988) <= (layer3_outputs(3974)) or (layer3_outputs(3035));
    layer4_outputs(1989) <= '0';
    layer4_outputs(1990) <= layer3_outputs(3173);
    layer4_outputs(1991) <= (layer3_outputs(4315)) and (layer3_outputs(3715));
    layer4_outputs(1992) <= layer3_outputs(756);
    layer4_outputs(1993) <= layer3_outputs(416);
    layer4_outputs(1994) <= (layer3_outputs(1667)) and (layer3_outputs(4529));
    layer4_outputs(1995) <= not((layer3_outputs(2177)) and (layer3_outputs(3767)));
    layer4_outputs(1996) <= not((layer3_outputs(4784)) xor (layer3_outputs(2793)));
    layer4_outputs(1997) <= (layer3_outputs(516)) and not (layer3_outputs(2191));
    layer4_outputs(1998) <= layer3_outputs(4792);
    layer4_outputs(1999) <= not((layer3_outputs(3754)) and (layer3_outputs(4165)));
    layer4_outputs(2000) <= (layer3_outputs(2199)) and (layer3_outputs(3525));
    layer4_outputs(2001) <= (layer3_outputs(800)) and not (layer3_outputs(2852));
    layer4_outputs(2002) <= (layer3_outputs(3085)) and not (layer3_outputs(419));
    layer4_outputs(2003) <= layer3_outputs(3647);
    layer4_outputs(2004) <= not(layer3_outputs(1352)) or (layer3_outputs(3288));
    layer4_outputs(2005) <= not((layer3_outputs(3033)) or (layer3_outputs(1920)));
    layer4_outputs(2006) <= layer3_outputs(3851);
    layer4_outputs(2007) <= (layer3_outputs(1619)) or (layer3_outputs(360));
    layer4_outputs(2008) <= layer3_outputs(3790);
    layer4_outputs(2009) <= not(layer3_outputs(5057));
    layer4_outputs(2010) <= not(layer3_outputs(4155));
    layer4_outputs(2011) <= '1';
    layer4_outputs(2012) <= not((layer3_outputs(4772)) and (layer3_outputs(991)));
    layer4_outputs(2013) <= not(layer3_outputs(3088));
    layer4_outputs(2014) <= layer3_outputs(3939);
    layer4_outputs(2015) <= not((layer3_outputs(67)) xor (layer3_outputs(541)));
    layer4_outputs(2016) <= (layer3_outputs(1509)) and (layer3_outputs(4218));
    layer4_outputs(2017) <= not(layer3_outputs(585)) or (layer3_outputs(4228));
    layer4_outputs(2018) <= not(layer3_outputs(1752)) or (layer3_outputs(450));
    layer4_outputs(2019) <= layer3_outputs(4202);
    layer4_outputs(2020) <= (layer3_outputs(151)) and not (layer3_outputs(4881));
    layer4_outputs(2021) <= (layer3_outputs(342)) and (layer3_outputs(4111));
    layer4_outputs(2022) <= layer3_outputs(2517);
    layer4_outputs(2023) <= (layer3_outputs(2358)) and not (layer3_outputs(4088));
    layer4_outputs(2024) <= not(layer3_outputs(4533));
    layer4_outputs(2025) <= layer3_outputs(3440);
    layer4_outputs(2026) <= not(layer3_outputs(3281));
    layer4_outputs(2027) <= (layer3_outputs(602)) and (layer3_outputs(3141));
    layer4_outputs(2028) <= not(layer3_outputs(1039));
    layer4_outputs(2029) <= not(layer3_outputs(3533));
    layer4_outputs(2030) <= layer3_outputs(4779);
    layer4_outputs(2031) <= layer3_outputs(4416);
    layer4_outputs(2032) <= layer3_outputs(1003);
    layer4_outputs(2033) <= layer3_outputs(393);
    layer4_outputs(2034) <= layer3_outputs(1154);
    layer4_outputs(2035) <= not(layer3_outputs(607)) or (layer3_outputs(2923));
    layer4_outputs(2036) <= not(layer3_outputs(1783));
    layer4_outputs(2037) <= layer3_outputs(1265);
    layer4_outputs(2038) <= not((layer3_outputs(4435)) xor (layer3_outputs(638)));
    layer4_outputs(2039) <= (layer3_outputs(1157)) and (layer3_outputs(2100));
    layer4_outputs(2040) <= (layer3_outputs(2042)) or (layer3_outputs(3549));
    layer4_outputs(2041) <= layer3_outputs(284);
    layer4_outputs(2042) <= layer3_outputs(1750);
    layer4_outputs(2043) <= not((layer3_outputs(201)) or (layer3_outputs(4862)));
    layer4_outputs(2044) <= not((layer3_outputs(4820)) and (layer3_outputs(1406)));
    layer4_outputs(2045) <= layer3_outputs(2967);
    layer4_outputs(2046) <= (layer3_outputs(8)) and not (layer3_outputs(2430));
    layer4_outputs(2047) <= (layer3_outputs(1251)) or (layer3_outputs(2346));
    layer4_outputs(2048) <= (layer3_outputs(1585)) and not (layer3_outputs(2541));
    layer4_outputs(2049) <= layer3_outputs(4099);
    layer4_outputs(2050) <= not(layer3_outputs(186)) or (layer3_outputs(4873));
    layer4_outputs(2051) <= layer3_outputs(5017);
    layer4_outputs(2052) <= not(layer3_outputs(4328));
    layer4_outputs(2053) <= (layer3_outputs(1255)) and not (layer3_outputs(4564));
    layer4_outputs(2054) <= layer3_outputs(1677);
    layer4_outputs(2055) <= not(layer3_outputs(2638)) or (layer3_outputs(2875));
    layer4_outputs(2056) <= layer3_outputs(2001);
    layer4_outputs(2057) <= not(layer3_outputs(1340));
    layer4_outputs(2058) <= (layer3_outputs(2974)) and (layer3_outputs(345));
    layer4_outputs(2059) <= not(layer3_outputs(3314)) or (layer3_outputs(2825));
    layer4_outputs(2060) <= not(layer3_outputs(2352));
    layer4_outputs(2061) <= layer3_outputs(958);
    layer4_outputs(2062) <= '1';
    layer4_outputs(2063) <= not(layer3_outputs(3576));
    layer4_outputs(2064) <= (layer3_outputs(4941)) and (layer3_outputs(3687));
    layer4_outputs(2065) <= (layer3_outputs(3474)) or (layer3_outputs(77));
    layer4_outputs(2066) <= layer3_outputs(2560);
    layer4_outputs(2067) <= layer3_outputs(1371);
    layer4_outputs(2068) <= not((layer3_outputs(539)) or (layer3_outputs(1819)));
    layer4_outputs(2069) <= (layer3_outputs(1846)) and not (layer3_outputs(1853));
    layer4_outputs(2070) <= (layer3_outputs(615)) and not (layer3_outputs(3700));
    layer4_outputs(2071) <= '1';
    layer4_outputs(2072) <= not(layer3_outputs(3328));
    layer4_outputs(2073) <= layer3_outputs(2354);
    layer4_outputs(2074) <= not(layer3_outputs(2301));
    layer4_outputs(2075) <= (layer3_outputs(3709)) xor (layer3_outputs(4375));
    layer4_outputs(2076) <= not(layer3_outputs(2276)) or (layer3_outputs(2348));
    layer4_outputs(2077) <= not((layer3_outputs(3820)) and (layer3_outputs(3282)));
    layer4_outputs(2078) <= layer3_outputs(1116);
    layer4_outputs(2079) <= not((layer3_outputs(1314)) and (layer3_outputs(2406)));
    layer4_outputs(2080) <= not(layer3_outputs(3580));
    layer4_outputs(2081) <= (layer3_outputs(1787)) or (layer3_outputs(532));
    layer4_outputs(2082) <= not(layer3_outputs(1001)) or (layer3_outputs(1295));
    layer4_outputs(2083) <= not(layer3_outputs(4636)) or (layer3_outputs(2744));
    layer4_outputs(2084) <= layer3_outputs(4392);
    layer4_outputs(2085) <= not(layer3_outputs(1321));
    layer4_outputs(2086) <= (layer3_outputs(4453)) xor (layer3_outputs(1621));
    layer4_outputs(2087) <= (layer3_outputs(1310)) and (layer3_outputs(625));
    layer4_outputs(2088) <= layer3_outputs(208);
    layer4_outputs(2089) <= not(layer3_outputs(833));
    layer4_outputs(2090) <= not(layer3_outputs(3202));
    layer4_outputs(2091) <= not(layer3_outputs(4291));
    layer4_outputs(2092) <= not((layer3_outputs(3071)) or (layer3_outputs(4634)));
    layer4_outputs(2093) <= not(layer3_outputs(1446)) or (layer3_outputs(1165));
    layer4_outputs(2094) <= not(layer3_outputs(2012));
    layer4_outputs(2095) <= layer3_outputs(1597);
    layer4_outputs(2096) <= layer3_outputs(2731);
    layer4_outputs(2097) <= not(layer3_outputs(3032));
    layer4_outputs(2098) <= not((layer3_outputs(4572)) and (layer3_outputs(2398)));
    layer4_outputs(2099) <= (layer3_outputs(4433)) or (layer3_outputs(3312));
    layer4_outputs(2100) <= not((layer3_outputs(470)) or (layer3_outputs(4808)));
    layer4_outputs(2101) <= layer3_outputs(2653);
    layer4_outputs(2102) <= layer3_outputs(2375);
    layer4_outputs(2103) <= (layer3_outputs(4821)) xor (layer3_outputs(655));
    layer4_outputs(2104) <= (layer3_outputs(2794)) and not (layer3_outputs(3338));
    layer4_outputs(2105) <= not(layer3_outputs(3673));
    layer4_outputs(2106) <= layer3_outputs(3248);
    layer4_outputs(2107) <= layer3_outputs(1759);
    layer4_outputs(2108) <= not(layer3_outputs(641));
    layer4_outputs(2109) <= layer3_outputs(4761);
    layer4_outputs(2110) <= (layer3_outputs(3914)) or (layer3_outputs(2064));
    layer4_outputs(2111) <= not(layer3_outputs(1047)) or (layer3_outputs(4355));
    layer4_outputs(2112) <= layer3_outputs(2770);
    layer4_outputs(2113) <= not(layer3_outputs(1967));
    layer4_outputs(2114) <= (layer3_outputs(3125)) and (layer3_outputs(2100));
    layer4_outputs(2115) <= not(layer3_outputs(2843));
    layer4_outputs(2116) <= not(layer3_outputs(1473)) or (layer3_outputs(3855));
    layer4_outputs(2117) <= '0';
    layer4_outputs(2118) <= layer3_outputs(195);
    layer4_outputs(2119) <= (layer3_outputs(4581)) and not (layer3_outputs(2148));
    layer4_outputs(2120) <= '0';
    layer4_outputs(2121) <= layer3_outputs(1061);
    layer4_outputs(2122) <= not(layer3_outputs(981)) or (layer3_outputs(4125));
    layer4_outputs(2123) <= not(layer3_outputs(2388)) or (layer3_outputs(516));
    layer4_outputs(2124) <= not((layer3_outputs(176)) and (layer3_outputs(3356)));
    layer4_outputs(2125) <= not((layer3_outputs(2585)) xor (layer3_outputs(3882)));
    layer4_outputs(2126) <= not(layer3_outputs(4720));
    layer4_outputs(2127) <= not(layer3_outputs(2932)) or (layer3_outputs(139));
    layer4_outputs(2128) <= not((layer3_outputs(59)) or (layer3_outputs(4457)));
    layer4_outputs(2129) <= not(layer3_outputs(1022));
    layer4_outputs(2130) <= layer3_outputs(4692);
    layer4_outputs(2131) <= not(layer3_outputs(701));
    layer4_outputs(2132) <= not(layer3_outputs(390));
    layer4_outputs(2133) <= '1';
    layer4_outputs(2134) <= not(layer3_outputs(4777)) or (layer3_outputs(5119));
    layer4_outputs(2135) <= (layer3_outputs(3691)) xor (layer3_outputs(3616));
    layer4_outputs(2136) <= not((layer3_outputs(2737)) or (layer3_outputs(305)));
    layer4_outputs(2137) <= not(layer3_outputs(2748));
    layer4_outputs(2138) <= not(layer3_outputs(1808));
    layer4_outputs(2139) <= not(layer3_outputs(4600));
    layer4_outputs(2140) <= (layer3_outputs(2605)) and not (layer3_outputs(4550));
    layer4_outputs(2141) <= not(layer3_outputs(1257));
    layer4_outputs(2142) <= not(layer3_outputs(1940));
    layer4_outputs(2143) <= (layer3_outputs(2390)) and (layer3_outputs(4932));
    layer4_outputs(2144) <= '1';
    layer4_outputs(2145) <= not(layer3_outputs(2461));
    layer4_outputs(2146) <= (layer3_outputs(2208)) and (layer3_outputs(2325));
    layer4_outputs(2147) <= layer3_outputs(173);
    layer4_outputs(2148) <= '0';
    layer4_outputs(2149) <= not((layer3_outputs(3189)) xor (layer3_outputs(3192)));
    layer4_outputs(2150) <= not(layer3_outputs(2599));
    layer4_outputs(2151) <= layer3_outputs(609);
    layer4_outputs(2152) <= (layer3_outputs(55)) and not (layer3_outputs(1483));
    layer4_outputs(2153) <= '1';
    layer4_outputs(2154) <= not(layer3_outputs(3796)) or (layer3_outputs(1216));
    layer4_outputs(2155) <= (layer3_outputs(4928)) or (layer3_outputs(4461));
    layer4_outputs(2156) <= (layer3_outputs(2511)) or (layer3_outputs(272));
    layer4_outputs(2157) <= not((layer3_outputs(2039)) or (layer3_outputs(3456)));
    layer4_outputs(2158) <= layer3_outputs(5066);
    layer4_outputs(2159) <= '0';
    layer4_outputs(2160) <= not(layer3_outputs(1314));
    layer4_outputs(2161) <= layer3_outputs(2933);
    layer4_outputs(2162) <= layer3_outputs(1285);
    layer4_outputs(2163) <= '1';
    layer4_outputs(2164) <= not((layer3_outputs(4130)) or (layer3_outputs(4178)));
    layer4_outputs(2165) <= (layer3_outputs(4442)) xor (layer3_outputs(1592));
    layer4_outputs(2166) <= not(layer3_outputs(728));
    layer4_outputs(2167) <= layer3_outputs(3679);
    layer4_outputs(2168) <= (layer3_outputs(210)) and (layer3_outputs(1905));
    layer4_outputs(2169) <= not((layer3_outputs(3240)) and (layer3_outputs(808)));
    layer4_outputs(2170) <= layer3_outputs(1518);
    layer4_outputs(2171) <= not(layer3_outputs(1875));
    layer4_outputs(2172) <= (layer3_outputs(1390)) and not (layer3_outputs(212));
    layer4_outputs(2173) <= '1';
    layer4_outputs(2174) <= (layer3_outputs(4717)) and not (layer3_outputs(1087));
    layer4_outputs(2175) <= (layer3_outputs(1182)) and (layer3_outputs(283));
    layer4_outputs(2176) <= not(layer3_outputs(4996));
    layer4_outputs(2177) <= not(layer3_outputs(4879));
    layer4_outputs(2178) <= not(layer3_outputs(972));
    layer4_outputs(2179) <= '1';
    layer4_outputs(2180) <= layer3_outputs(75);
    layer4_outputs(2181) <= not((layer3_outputs(4584)) or (layer3_outputs(2968)));
    layer4_outputs(2182) <= (layer3_outputs(4776)) and not (layer3_outputs(3957));
    layer4_outputs(2183) <= not(layer3_outputs(4624));
    layer4_outputs(2184) <= not(layer3_outputs(260)) or (layer3_outputs(353));
    layer4_outputs(2185) <= layer3_outputs(2493);
    layer4_outputs(2186) <= not((layer3_outputs(3145)) and (layer3_outputs(1130)));
    layer4_outputs(2187) <= not((layer3_outputs(759)) or (layer3_outputs(1412)));
    layer4_outputs(2188) <= not((layer3_outputs(4702)) or (layer3_outputs(2246)));
    layer4_outputs(2189) <= '0';
    layer4_outputs(2190) <= not(layer3_outputs(411)) or (layer3_outputs(1788));
    layer4_outputs(2191) <= (layer3_outputs(1898)) xor (layer3_outputs(2156));
    layer4_outputs(2192) <= not(layer3_outputs(1655)) or (layer3_outputs(352));
    layer4_outputs(2193) <= layer3_outputs(1524);
    layer4_outputs(2194) <= not((layer3_outputs(117)) xor (layer3_outputs(3708)));
    layer4_outputs(2195) <= (layer3_outputs(3075)) and (layer3_outputs(4047));
    layer4_outputs(2196) <= not(layer3_outputs(3734));
    layer4_outputs(2197) <= (layer3_outputs(4176)) or (layer3_outputs(521));
    layer4_outputs(2198) <= not(layer3_outputs(3220));
    layer4_outputs(2199) <= (layer3_outputs(3960)) and not (layer3_outputs(2729));
    layer4_outputs(2200) <= (layer3_outputs(4239)) and not (layer3_outputs(4873));
    layer4_outputs(2201) <= (layer3_outputs(2804)) and not (layer3_outputs(2193));
    layer4_outputs(2202) <= (layer3_outputs(144)) and (layer3_outputs(1965));
    layer4_outputs(2203) <= (layer3_outputs(2878)) or (layer3_outputs(1473));
    layer4_outputs(2204) <= not((layer3_outputs(4708)) or (layer3_outputs(101)));
    layer4_outputs(2205) <= not((layer3_outputs(2391)) and (layer3_outputs(1210)));
    layer4_outputs(2206) <= (layer3_outputs(238)) and (layer3_outputs(1576));
    layer4_outputs(2207) <= layer3_outputs(1852);
    layer4_outputs(2208) <= not(layer3_outputs(483));
    layer4_outputs(2209) <= layer3_outputs(1564);
    layer4_outputs(2210) <= not(layer3_outputs(55));
    layer4_outputs(2211) <= not(layer3_outputs(4148)) or (layer3_outputs(3503));
    layer4_outputs(2212) <= not((layer3_outputs(2181)) and (layer3_outputs(1617)));
    layer4_outputs(2213) <= (layer3_outputs(888)) or (layer3_outputs(240));
    layer4_outputs(2214) <= not(layer3_outputs(795)) or (layer3_outputs(4931));
    layer4_outputs(2215) <= not(layer3_outputs(2083));
    layer4_outputs(2216) <= (layer3_outputs(2783)) and not (layer3_outputs(316));
    layer4_outputs(2217) <= '1';
    layer4_outputs(2218) <= (layer3_outputs(3948)) and not (layer3_outputs(1593));
    layer4_outputs(2219) <= (layer3_outputs(1201)) or (layer3_outputs(1494));
    layer4_outputs(2220) <= '0';
    layer4_outputs(2221) <= layer3_outputs(359);
    layer4_outputs(2222) <= not((layer3_outputs(1876)) and (layer3_outputs(4102)));
    layer4_outputs(2223) <= not(layer3_outputs(1266)) or (layer3_outputs(731));
    layer4_outputs(2224) <= not(layer3_outputs(1047));
    layer4_outputs(2225) <= (layer3_outputs(1332)) xor (layer3_outputs(632));
    layer4_outputs(2226) <= layer3_outputs(3661);
    layer4_outputs(2227) <= not(layer3_outputs(3502));
    layer4_outputs(2228) <= not(layer3_outputs(2487)) or (layer3_outputs(3841));
    layer4_outputs(2229) <= layer3_outputs(1576);
    layer4_outputs(2230) <= not(layer3_outputs(56));
    layer4_outputs(2231) <= not(layer3_outputs(1470)) or (layer3_outputs(3273));
    layer4_outputs(2232) <= layer3_outputs(4490);
    layer4_outputs(2233) <= not(layer3_outputs(2149));
    layer4_outputs(2234) <= not(layer3_outputs(1380)) or (layer3_outputs(869));
    layer4_outputs(2235) <= not(layer3_outputs(4689)) or (layer3_outputs(1949));
    layer4_outputs(2236) <= not(layer3_outputs(5077)) or (layer3_outputs(1909));
    layer4_outputs(2237) <= not((layer3_outputs(4251)) and (layer3_outputs(2044)));
    layer4_outputs(2238) <= (layer3_outputs(4655)) or (layer3_outputs(1156));
    layer4_outputs(2239) <= not(layer3_outputs(1658)) or (layer3_outputs(5038));
    layer4_outputs(2240) <= (layer3_outputs(1387)) or (layer3_outputs(4850));
    layer4_outputs(2241) <= not(layer3_outputs(1849)) or (layer3_outputs(4050));
    layer4_outputs(2242) <= not(layer3_outputs(549));
    layer4_outputs(2243) <= '0';
    layer4_outputs(2244) <= layer3_outputs(2345);
    layer4_outputs(2245) <= not(layer3_outputs(2959)) or (layer3_outputs(4052));
    layer4_outputs(2246) <= (layer3_outputs(2914)) xor (layer3_outputs(2304));
    layer4_outputs(2247) <= (layer3_outputs(1079)) and not (layer3_outputs(954));
    layer4_outputs(2248) <= not((layer3_outputs(29)) or (layer3_outputs(1684)));
    layer4_outputs(2249) <= layer3_outputs(2085);
    layer4_outputs(2250) <= (layer3_outputs(2891)) xor (layer3_outputs(2594));
    layer4_outputs(2251) <= (layer3_outputs(702)) and not (layer3_outputs(1307));
    layer4_outputs(2252) <= not((layer3_outputs(3744)) and (layer3_outputs(3702)));
    layer4_outputs(2253) <= not(layer3_outputs(384));
    layer4_outputs(2254) <= not(layer3_outputs(4359)) or (layer3_outputs(3063));
    layer4_outputs(2255) <= not(layer3_outputs(587));
    layer4_outputs(2256) <= (layer3_outputs(52)) and not (layer3_outputs(4683));
    layer4_outputs(2257) <= not(layer3_outputs(1018));
    layer4_outputs(2258) <= (layer3_outputs(1546)) and not (layer3_outputs(2211));
    layer4_outputs(2259) <= not(layer3_outputs(4874)) or (layer3_outputs(4822));
    layer4_outputs(2260) <= not(layer3_outputs(2740));
    layer4_outputs(2261) <= not(layer3_outputs(3254)) or (layer3_outputs(5114));
    layer4_outputs(2262) <= '1';
    layer4_outputs(2263) <= layer3_outputs(5096);
    layer4_outputs(2264) <= (layer3_outputs(2058)) and (layer3_outputs(3442));
    layer4_outputs(2265) <= (layer3_outputs(2224)) or (layer3_outputs(1224));
    layer4_outputs(2266) <= layer3_outputs(2281);
    layer4_outputs(2267) <= layer3_outputs(2466);
    layer4_outputs(2268) <= not(layer3_outputs(4070));
    layer4_outputs(2269) <= (layer3_outputs(4689)) xor (layer3_outputs(2672));
    layer4_outputs(2270) <= layer3_outputs(1078);
    layer4_outputs(2271) <= (layer3_outputs(2499)) or (layer3_outputs(2016));
    layer4_outputs(2272) <= not(layer3_outputs(1932));
    layer4_outputs(2273) <= not((layer3_outputs(4508)) xor (layer3_outputs(3115)));
    layer4_outputs(2274) <= '1';
    layer4_outputs(2275) <= not((layer3_outputs(163)) and (layer3_outputs(1450)));
    layer4_outputs(2276) <= layer3_outputs(3272);
    layer4_outputs(2277) <= layer3_outputs(3455);
    layer4_outputs(2278) <= not(layer3_outputs(4923)) or (layer3_outputs(438));
    layer4_outputs(2279) <= not(layer3_outputs(619));
    layer4_outputs(2280) <= '1';
    layer4_outputs(2281) <= layer3_outputs(2000);
    layer4_outputs(2282) <= (layer3_outputs(3592)) xor (layer3_outputs(4664));
    layer4_outputs(2283) <= '1';
    layer4_outputs(2284) <= layer3_outputs(4881);
    layer4_outputs(2285) <= not(layer3_outputs(1482));
    layer4_outputs(2286) <= not(layer3_outputs(3340));
    layer4_outputs(2287) <= layer3_outputs(1687);
    layer4_outputs(2288) <= (layer3_outputs(1271)) xor (layer3_outputs(3313));
    layer4_outputs(2289) <= (layer3_outputs(1014)) and not (layer3_outputs(2172));
    layer4_outputs(2290) <= (layer3_outputs(2047)) and not (layer3_outputs(4466));
    layer4_outputs(2291) <= (layer3_outputs(2296)) or (layer3_outputs(3371));
    layer4_outputs(2292) <= not((layer3_outputs(1754)) xor (layer3_outputs(3737)));
    layer4_outputs(2293) <= not(layer3_outputs(3520)) or (layer3_outputs(4826));
    layer4_outputs(2294) <= (layer3_outputs(1313)) and (layer3_outputs(1296));
    layer4_outputs(2295) <= (layer3_outputs(3346)) or (layer3_outputs(1094));
    layer4_outputs(2296) <= (layer3_outputs(1793)) and (layer3_outputs(2049));
    layer4_outputs(2297) <= not(layer3_outputs(2966)) or (layer3_outputs(3682));
    layer4_outputs(2298) <= '1';
    layer4_outputs(2299) <= layer3_outputs(3410);
    layer4_outputs(2300) <= not((layer3_outputs(3995)) or (layer3_outputs(4654)));
    layer4_outputs(2301) <= (layer3_outputs(501)) and (layer3_outputs(2688));
    layer4_outputs(2302) <= (layer3_outputs(4241)) and not (layer3_outputs(2881));
    layer4_outputs(2303) <= not(layer3_outputs(4053)) or (layer3_outputs(4113));
    layer4_outputs(2304) <= not(layer3_outputs(2279));
    layer4_outputs(2305) <= (layer3_outputs(3568)) xor (layer3_outputs(3464));
    layer4_outputs(2306) <= layer3_outputs(1006);
    layer4_outputs(2307) <= layer3_outputs(3049);
    layer4_outputs(2308) <= layer3_outputs(3268);
    layer4_outputs(2309) <= not((layer3_outputs(2546)) and (layer3_outputs(905)));
    layer4_outputs(2310) <= not((layer3_outputs(2256)) or (layer3_outputs(3399)));
    layer4_outputs(2311) <= '0';
    layer4_outputs(2312) <= not(layer3_outputs(3364));
    layer4_outputs(2313) <= (layer3_outputs(1736)) xor (layer3_outputs(649));
    layer4_outputs(2314) <= not(layer3_outputs(518)) or (layer3_outputs(4434));
    layer4_outputs(2315) <= not((layer3_outputs(859)) and (layer3_outputs(4818)));
    layer4_outputs(2316) <= not(layer3_outputs(5115)) or (layer3_outputs(2665));
    layer4_outputs(2317) <= (layer3_outputs(2675)) and not (layer3_outputs(2569));
    layer4_outputs(2318) <= not((layer3_outputs(3496)) or (layer3_outputs(2831)));
    layer4_outputs(2319) <= (layer3_outputs(4659)) or (layer3_outputs(1533));
    layer4_outputs(2320) <= (layer3_outputs(2230)) or (layer3_outputs(2403));
    layer4_outputs(2321) <= not((layer3_outputs(4835)) and (layer3_outputs(1893)));
    layer4_outputs(2322) <= (layer3_outputs(3256)) and not (layer3_outputs(864));
    layer4_outputs(2323) <= layer3_outputs(2136);
    layer4_outputs(2324) <= not(layer3_outputs(1306));
    layer4_outputs(2325) <= not(layer3_outputs(3691));
    layer4_outputs(2326) <= not((layer3_outputs(80)) and (layer3_outputs(2948)));
    layer4_outputs(2327) <= not(layer3_outputs(1694));
    layer4_outputs(2328) <= not(layer3_outputs(713)) or (layer3_outputs(2588));
    layer4_outputs(2329) <= (layer3_outputs(492)) and not (layer3_outputs(3201));
    layer4_outputs(2330) <= not(layer3_outputs(3037)) or (layer3_outputs(473));
    layer4_outputs(2331) <= (layer3_outputs(3950)) or (layer3_outputs(2169));
    layer4_outputs(2332) <= layer3_outputs(2557);
    layer4_outputs(2333) <= (layer3_outputs(1960)) and (layer3_outputs(2331));
    layer4_outputs(2334) <= (layer3_outputs(879)) and not (layer3_outputs(2432));
    layer4_outputs(2335) <= not(layer3_outputs(964));
    layer4_outputs(2336) <= (layer3_outputs(78)) or (layer3_outputs(1832));
    layer4_outputs(2337) <= (layer3_outputs(4837)) or (layer3_outputs(2555));
    layer4_outputs(2338) <= layer3_outputs(2299);
    layer4_outputs(2339) <= not(layer3_outputs(4422)) or (layer3_outputs(152));
    layer4_outputs(2340) <= not((layer3_outputs(2630)) and (layer3_outputs(2221)));
    layer4_outputs(2341) <= layer3_outputs(4742);
    layer4_outputs(2342) <= not((layer3_outputs(2682)) xor (layer3_outputs(3420)));
    layer4_outputs(2343) <= (layer3_outputs(535)) xor (layer3_outputs(1573));
    layer4_outputs(2344) <= (layer3_outputs(1255)) and not (layer3_outputs(334));
    layer4_outputs(2345) <= layer3_outputs(4350);
    layer4_outputs(2346) <= layer3_outputs(2763);
    layer4_outputs(2347) <= '0';
    layer4_outputs(2348) <= (layer3_outputs(2080)) and (layer3_outputs(5100));
    layer4_outputs(2349) <= not(layer3_outputs(4074));
    layer4_outputs(2350) <= (layer3_outputs(1776)) and (layer3_outputs(1518));
    layer4_outputs(2351) <= not((layer3_outputs(3054)) and (layer3_outputs(2405)));
    layer4_outputs(2352) <= not(layer3_outputs(2503)) or (layer3_outputs(997));
    layer4_outputs(2353) <= not((layer3_outputs(137)) or (layer3_outputs(1896)));
    layer4_outputs(2354) <= '1';
    layer4_outputs(2355) <= (layer3_outputs(3123)) and not (layer3_outputs(1143));
    layer4_outputs(2356) <= (layer3_outputs(1191)) and not (layer3_outputs(2498));
    layer4_outputs(2357) <= not(layer3_outputs(2258)) or (layer3_outputs(1015));
    layer4_outputs(2358) <= '0';
    layer4_outputs(2359) <= layer3_outputs(575);
    layer4_outputs(2360) <= layer3_outputs(498);
    layer4_outputs(2361) <= not((layer3_outputs(627)) xor (layer3_outputs(5076)));
    layer4_outputs(2362) <= not((layer3_outputs(3165)) and (layer3_outputs(4570)));
    layer4_outputs(2363) <= (layer3_outputs(528)) and not (layer3_outputs(5041));
    layer4_outputs(2364) <= layer3_outputs(4391);
    layer4_outputs(2365) <= layer3_outputs(714);
    layer4_outputs(2366) <= layer3_outputs(1613);
    layer4_outputs(2367) <= not(layer3_outputs(3940));
    layer4_outputs(2368) <= not((layer3_outputs(1799)) xor (layer3_outputs(2023)));
    layer4_outputs(2369) <= not(layer3_outputs(2530));
    layer4_outputs(2370) <= not(layer3_outputs(4663));
    layer4_outputs(2371) <= layer3_outputs(1249);
    layer4_outputs(2372) <= not(layer3_outputs(3204)) or (layer3_outputs(1981));
    layer4_outputs(2373) <= layer3_outputs(4248);
    layer4_outputs(2374) <= (layer3_outputs(4725)) and (layer3_outputs(3182));
    layer4_outputs(2375) <= not(layer3_outputs(1847)) or (layer3_outputs(3285));
    layer4_outputs(2376) <= (layer3_outputs(3535)) or (layer3_outputs(4805));
    layer4_outputs(2377) <= '1';
    layer4_outputs(2378) <= not(layer3_outputs(1163));
    layer4_outputs(2379) <= (layer3_outputs(4601)) and not (layer3_outputs(392));
    layer4_outputs(2380) <= not(layer3_outputs(1504));
    layer4_outputs(2381) <= (layer3_outputs(1018)) and not (layer3_outputs(1113));
    layer4_outputs(2382) <= not(layer3_outputs(3377));
    layer4_outputs(2383) <= (layer3_outputs(4575)) and not (layer3_outputs(865));
    layer4_outputs(2384) <= not(layer3_outputs(979));
    layer4_outputs(2385) <= not((layer3_outputs(4907)) or (layer3_outputs(1420)));
    layer4_outputs(2386) <= not(layer3_outputs(4062));
    layer4_outputs(2387) <= not(layer3_outputs(2564)) or (layer3_outputs(1980));
    layer4_outputs(2388) <= (layer3_outputs(4558)) and (layer3_outputs(2551));
    layer4_outputs(2389) <= layer3_outputs(5118);
    layer4_outputs(2390) <= layer3_outputs(44);
    layer4_outputs(2391) <= not(layer3_outputs(3140)) or (layer3_outputs(3224));
    layer4_outputs(2392) <= (layer3_outputs(4874)) xor (layer3_outputs(1545));
    layer4_outputs(2393) <= '0';
    layer4_outputs(2394) <= layer3_outputs(4982);
    layer4_outputs(2395) <= not(layer3_outputs(1089));
    layer4_outputs(2396) <= not(layer3_outputs(747)) or (layer3_outputs(1480));
    layer4_outputs(2397) <= not(layer3_outputs(4346));
    layer4_outputs(2398) <= not(layer3_outputs(4738));
    layer4_outputs(2399) <= not(layer3_outputs(4405)) or (layer3_outputs(3425));
    layer4_outputs(2400) <= not(layer3_outputs(961));
    layer4_outputs(2401) <= layer3_outputs(3266);
    layer4_outputs(2402) <= not(layer3_outputs(898)) or (layer3_outputs(323));
    layer4_outputs(2403) <= not(layer3_outputs(1150));
    layer4_outputs(2404) <= not((layer3_outputs(3789)) or (layer3_outputs(717)));
    layer4_outputs(2405) <= layer3_outputs(4512);
    layer4_outputs(2406) <= not(layer3_outputs(1098)) or (layer3_outputs(4971));
    layer4_outputs(2407) <= '1';
    layer4_outputs(2408) <= '0';
    layer4_outputs(2409) <= (layer3_outputs(3004)) and not (layer3_outputs(1187));
    layer4_outputs(2410) <= not((layer3_outputs(1154)) xor (layer3_outputs(3118)));
    layer4_outputs(2411) <= (layer3_outputs(3981)) and not (layer3_outputs(292));
    layer4_outputs(2412) <= layer3_outputs(508);
    layer4_outputs(2413) <= (layer3_outputs(3066)) and (layer3_outputs(4031));
    layer4_outputs(2414) <= (layer3_outputs(4917)) and not (layer3_outputs(2310));
    layer4_outputs(2415) <= layer3_outputs(1874);
    layer4_outputs(2416) <= '1';
    layer4_outputs(2417) <= not(layer3_outputs(4071));
    layer4_outputs(2418) <= not(layer3_outputs(1815));
    layer4_outputs(2419) <= (layer3_outputs(578)) and not (layer3_outputs(1468));
    layer4_outputs(2420) <= layer3_outputs(3928);
    layer4_outputs(2421) <= not(layer3_outputs(2789));
    layer4_outputs(2422) <= layer3_outputs(4144);
    layer4_outputs(2423) <= not(layer3_outputs(4285)) or (layer3_outputs(3748));
    layer4_outputs(2424) <= layer3_outputs(1696);
    layer4_outputs(2425) <= layer3_outputs(2692);
    layer4_outputs(2426) <= not(layer3_outputs(517)) or (layer3_outputs(3771));
    layer4_outputs(2427) <= not(layer3_outputs(1939));
    layer4_outputs(2428) <= not(layer3_outputs(3364)) or (layer3_outputs(447));
    layer4_outputs(2429) <= not((layer3_outputs(337)) xor (layer3_outputs(2263)));
    layer4_outputs(2430) <= not(layer3_outputs(1136));
    layer4_outputs(2431) <= layer3_outputs(2419);
    layer4_outputs(2432) <= layer3_outputs(2137);
    layer4_outputs(2433) <= not(layer3_outputs(149)) or (layer3_outputs(1133));
    layer4_outputs(2434) <= not((layer3_outputs(4223)) or (layer3_outputs(4382)));
    layer4_outputs(2435) <= not(layer3_outputs(1365));
    layer4_outputs(2436) <= not(layer3_outputs(477)) or (layer3_outputs(1066));
    layer4_outputs(2437) <= layer3_outputs(766);
    layer4_outputs(2438) <= not(layer3_outputs(4412));
    layer4_outputs(2439) <= layer3_outputs(2027);
    layer4_outputs(2440) <= not(layer3_outputs(4684));
    layer4_outputs(2441) <= (layer3_outputs(4310)) and not (layer3_outputs(2755));
    layer4_outputs(2442) <= (layer3_outputs(3163)) and not (layer3_outputs(320));
    layer4_outputs(2443) <= not(layer3_outputs(986));
    layer4_outputs(2444) <= not(layer3_outputs(2908));
    layer4_outputs(2445) <= not(layer3_outputs(1671)) or (layer3_outputs(4327));
    layer4_outputs(2446) <= layer3_outputs(1652);
    layer4_outputs(2447) <= layer3_outputs(370);
    layer4_outputs(2448) <= layer3_outputs(3990);
    layer4_outputs(2449) <= layer3_outputs(1279);
    layer4_outputs(2450) <= not(layer3_outputs(904));
    layer4_outputs(2451) <= not(layer3_outputs(1517));
    layer4_outputs(2452) <= not((layer3_outputs(479)) and (layer3_outputs(1120)));
    layer4_outputs(2453) <= not((layer3_outputs(48)) or (layer3_outputs(696)));
    layer4_outputs(2454) <= (layer3_outputs(2237)) and (layer3_outputs(2010));
    layer4_outputs(2455) <= not(layer3_outputs(884)) or (layer3_outputs(4471));
    layer4_outputs(2456) <= not(layer3_outputs(4423));
    layer4_outputs(2457) <= layer3_outputs(192);
    layer4_outputs(2458) <= not(layer3_outputs(4267));
    layer4_outputs(2459) <= not(layer3_outputs(3352));
    layer4_outputs(2460) <= '1';
    layer4_outputs(2461) <= not(layer3_outputs(4531));
    layer4_outputs(2462) <= layer3_outputs(4809);
    layer4_outputs(2463) <= layer3_outputs(3903);
    layer4_outputs(2464) <= layer3_outputs(1627);
    layer4_outputs(2465) <= not(layer3_outputs(2829)) or (layer3_outputs(3781));
    layer4_outputs(2466) <= not(layer3_outputs(4743)) or (layer3_outputs(877));
    layer4_outputs(2467) <= not(layer3_outputs(4271)) or (layer3_outputs(3758));
    layer4_outputs(2468) <= (layer3_outputs(4562)) xor (layer3_outputs(1957));
    layer4_outputs(2469) <= layer3_outputs(1050);
    layer4_outputs(2470) <= not(layer3_outputs(378)) or (layer3_outputs(4194));
    layer4_outputs(2471) <= '1';
    layer4_outputs(2472) <= '1';
    layer4_outputs(2473) <= (layer3_outputs(643)) or (layer3_outputs(22));
    layer4_outputs(2474) <= '0';
    layer4_outputs(2475) <= (layer3_outputs(1578)) and (layer3_outputs(4080));
    layer4_outputs(2476) <= not((layer3_outputs(4168)) xor (layer3_outputs(2396)));
    layer4_outputs(2477) <= '0';
    layer4_outputs(2478) <= layer3_outputs(835);
    layer4_outputs(2479) <= not(layer3_outputs(4710));
    layer4_outputs(2480) <= (layer3_outputs(377)) or (layer3_outputs(3779));
    layer4_outputs(2481) <= '1';
    layer4_outputs(2482) <= not((layer3_outputs(2015)) xor (layer3_outputs(4027)));
    layer4_outputs(2483) <= not(layer3_outputs(1370));
    layer4_outputs(2484) <= (layer3_outputs(2749)) xor (layer3_outputs(5022));
    layer4_outputs(2485) <= layer3_outputs(361);
    layer4_outputs(2486) <= not(layer3_outputs(3449)) or (layer3_outputs(1106));
    layer4_outputs(2487) <= layer3_outputs(1164);
    layer4_outputs(2488) <= layer3_outputs(1375);
    layer4_outputs(2489) <= not(layer3_outputs(1076));
    layer4_outputs(2490) <= not((layer3_outputs(4237)) or (layer3_outputs(4404)));
    layer4_outputs(2491) <= '0';
    layer4_outputs(2492) <= layer3_outputs(2925);
    layer4_outputs(2493) <= not(layer3_outputs(2188)) or (layer3_outputs(4682));
    layer4_outputs(2494) <= (layer3_outputs(1318)) and (layer3_outputs(2173));
    layer4_outputs(2495) <= not(layer3_outputs(2415));
    layer4_outputs(2496) <= not(layer3_outputs(2722));
    layer4_outputs(2497) <= not(layer3_outputs(1126));
    layer4_outputs(2498) <= layer3_outputs(846);
    layer4_outputs(2499) <= not((layer3_outputs(2844)) and (layer3_outputs(3166)));
    layer4_outputs(2500) <= (layer3_outputs(2426)) xor (layer3_outputs(1480));
    layer4_outputs(2501) <= not((layer3_outputs(701)) or (layer3_outputs(4560)));
    layer4_outputs(2502) <= not(layer3_outputs(421));
    layer4_outputs(2503) <= (layer3_outputs(3022)) and not (layer3_outputs(1645));
    layer4_outputs(2504) <= not((layer3_outputs(5103)) and (layer3_outputs(2454)));
    layer4_outputs(2505) <= not(layer3_outputs(1270));
    layer4_outputs(2506) <= not(layer3_outputs(284));
    layer4_outputs(2507) <= (layer3_outputs(1721)) or (layer3_outputs(4924));
    layer4_outputs(2508) <= not((layer3_outputs(3404)) xor (layer3_outputs(2572)));
    layer4_outputs(2509) <= not((layer3_outputs(3290)) and (layer3_outputs(469)));
    layer4_outputs(2510) <= not((layer3_outputs(1965)) and (layer3_outputs(956)));
    layer4_outputs(2511) <= (layer3_outputs(4631)) and (layer3_outputs(4263));
    layer4_outputs(2512) <= not(layer3_outputs(1570));
    layer4_outputs(2513) <= layer3_outputs(4516);
    layer4_outputs(2514) <= (layer3_outputs(2437)) and (layer3_outputs(460));
    layer4_outputs(2515) <= not(layer3_outputs(950));
    layer4_outputs(2516) <= not(layer3_outputs(1438));
    layer4_outputs(2517) <= (layer3_outputs(858)) and not (layer3_outputs(3931));
    layer4_outputs(2518) <= not(layer3_outputs(1301));
    layer4_outputs(2519) <= layer3_outputs(4763);
    layer4_outputs(2520) <= layer3_outputs(1293);
    layer4_outputs(2521) <= layer3_outputs(3918);
    layer4_outputs(2522) <= (layer3_outputs(3382)) and not (layer3_outputs(1715));
    layer4_outputs(2523) <= not(layer3_outputs(2513)) or (layer3_outputs(1934));
    layer4_outputs(2524) <= not(layer3_outputs(3432)) or (layer3_outputs(5080));
    layer4_outputs(2525) <= not((layer3_outputs(1922)) xor (layer3_outputs(4348)));
    layer4_outputs(2526) <= layer3_outputs(114);
    layer4_outputs(2527) <= (layer3_outputs(1023)) and not (layer3_outputs(3188));
    layer4_outputs(2528) <= not(layer3_outputs(2270)) or (layer3_outputs(1054));
    layer4_outputs(2529) <= (layer3_outputs(4994)) and (layer3_outputs(487));
    layer4_outputs(2530) <= not((layer3_outputs(2567)) and (layer3_outputs(27)));
    layer4_outputs(2531) <= (layer3_outputs(2889)) xor (layer3_outputs(2830));
    layer4_outputs(2532) <= not((layer3_outputs(3144)) and (layer3_outputs(1253)));
    layer4_outputs(2533) <= not(layer3_outputs(1417));
    layer4_outputs(2534) <= not(layer3_outputs(1726));
    layer4_outputs(2535) <= not((layer3_outputs(1296)) and (layer3_outputs(1966)));
    layer4_outputs(2536) <= not(layer3_outputs(4499)) or (layer3_outputs(4614));
    layer4_outputs(2537) <= '1';
    layer4_outputs(2538) <= not(layer3_outputs(1891)) or (layer3_outputs(3868));
    layer4_outputs(2539) <= not(layer3_outputs(4056));
    layer4_outputs(2540) <= not((layer3_outputs(2098)) or (layer3_outputs(3195)));
    layer4_outputs(2541) <= not(layer3_outputs(4552));
    layer4_outputs(2542) <= (layer3_outputs(2189)) or (layer3_outputs(926));
    layer4_outputs(2543) <= (layer3_outputs(3725)) and not (layer3_outputs(123));
    layer4_outputs(2544) <= layer3_outputs(4128);
    layer4_outputs(2545) <= layer3_outputs(1033);
    layer4_outputs(2546) <= not((layer3_outputs(3590)) and (layer3_outputs(540)));
    layer4_outputs(2547) <= (layer3_outputs(3471)) and (layer3_outputs(2328));
    layer4_outputs(2548) <= not((layer3_outputs(2389)) or (layer3_outputs(1989)));
    layer4_outputs(2549) <= not((layer3_outputs(1861)) xor (layer3_outputs(2938)));
    layer4_outputs(2550) <= not(layer3_outputs(5));
    layer4_outputs(2551) <= not(layer3_outputs(1030));
    layer4_outputs(2552) <= layer3_outputs(4697);
    layer4_outputs(2553) <= not(layer3_outputs(3385));
    layer4_outputs(2554) <= not(layer3_outputs(3859)) or (layer3_outputs(2326));
    layer4_outputs(2555) <= not(layer3_outputs(905));
    layer4_outputs(2556) <= layer3_outputs(1830);
    layer4_outputs(2557) <= layer3_outputs(3638);
    layer4_outputs(2558) <= not(layer3_outputs(4697));
    layer4_outputs(2559) <= not(layer3_outputs(3354));
    layer4_outputs(2560) <= (layer3_outputs(3054)) and not (layer3_outputs(2393));
    layer4_outputs(2561) <= (layer3_outputs(514)) and (layer3_outputs(2649));
    layer4_outputs(2562) <= layer3_outputs(2747);
    layer4_outputs(2563) <= (layer3_outputs(3531)) and (layer3_outputs(116));
    layer4_outputs(2564) <= not(layer3_outputs(257));
    layer4_outputs(2565) <= not(layer3_outputs(655)) or (layer3_outputs(298));
    layer4_outputs(2566) <= (layer3_outputs(4987)) or (layer3_outputs(4930));
    layer4_outputs(2567) <= (layer3_outputs(108)) or (layer3_outputs(410));
    layer4_outputs(2568) <= '0';
    layer4_outputs(2569) <= not((layer3_outputs(2074)) and (layer3_outputs(4090)));
    layer4_outputs(2570) <= not(layer3_outputs(2849)) or (layer3_outputs(1027));
    layer4_outputs(2571) <= (layer3_outputs(2817)) and not (layer3_outputs(46));
    layer4_outputs(2572) <= layer3_outputs(1200);
    layer4_outputs(2573) <= not(layer3_outputs(4496));
    layer4_outputs(2574) <= '0';
    layer4_outputs(2575) <= not(layer3_outputs(3058));
    layer4_outputs(2576) <= not((layer3_outputs(3250)) xor (layer3_outputs(247)));
    layer4_outputs(2577) <= layer3_outputs(1555);
    layer4_outputs(2578) <= not(layer3_outputs(3173)) or (layer3_outputs(3));
    layer4_outputs(2579) <= not(layer3_outputs(3435));
    layer4_outputs(2580) <= (layer3_outputs(2819)) and not (layer3_outputs(1610));
    layer4_outputs(2581) <= not(layer3_outputs(4627));
    layer4_outputs(2582) <= not(layer3_outputs(2510));
    layer4_outputs(2583) <= not(layer3_outputs(1586));
    layer4_outputs(2584) <= not(layer3_outputs(4966));
    layer4_outputs(2585) <= not((layer3_outputs(2269)) or (layer3_outputs(3083)));
    layer4_outputs(2586) <= (layer3_outputs(2515)) and (layer3_outputs(2159));
    layer4_outputs(2587) <= (layer3_outputs(53)) and (layer3_outputs(4112));
    layer4_outputs(2588) <= '1';
    layer4_outputs(2589) <= layer3_outputs(3928);
    layer4_outputs(2590) <= not(layer3_outputs(341)) or (layer3_outputs(3544));
    layer4_outputs(2591) <= '1';
    layer4_outputs(2592) <= not((layer3_outputs(3658)) and (layer3_outputs(3064)));
    layer4_outputs(2593) <= not(layer3_outputs(4256));
    layer4_outputs(2594) <= not(layer3_outputs(1250));
    layer4_outputs(2595) <= not(layer3_outputs(4581)) or (layer3_outputs(2278));
    layer4_outputs(2596) <= (layer3_outputs(3286)) and not (layer3_outputs(1405));
    layer4_outputs(2597) <= not((layer3_outputs(3780)) or (layer3_outputs(5004)));
    layer4_outputs(2598) <= (layer3_outputs(1959)) and (layer3_outputs(2655));
    layer4_outputs(2599) <= '1';
    layer4_outputs(2600) <= layer3_outputs(1563);
    layer4_outputs(2601) <= (layer3_outputs(5020)) and (layer3_outputs(4236));
    layer4_outputs(2602) <= not((layer3_outputs(1321)) and (layer3_outputs(3353)));
    layer4_outputs(2603) <= (layer3_outputs(4309)) and not (layer3_outputs(2634));
    layer4_outputs(2604) <= '0';
    layer4_outputs(2605) <= not(layer3_outputs(2826));
    layer4_outputs(2606) <= not(layer3_outputs(4251));
    layer4_outputs(2607) <= not(layer3_outputs(3434)) or (layer3_outputs(2971));
    layer4_outputs(2608) <= (layer3_outputs(338)) and not (layer3_outputs(736));
    layer4_outputs(2609) <= (layer3_outputs(3846)) and not (layer3_outputs(665));
    layer4_outputs(2610) <= layer3_outputs(3545);
    layer4_outputs(2611) <= (layer3_outputs(1043)) and not (layer3_outputs(538));
    layer4_outputs(2612) <= layer3_outputs(2783);
    layer4_outputs(2613) <= layer3_outputs(1695);
    layer4_outputs(2614) <= not((layer3_outputs(1097)) or (layer3_outputs(2780)));
    layer4_outputs(2615) <= (layer3_outputs(2863)) and (layer3_outputs(1005));
    layer4_outputs(2616) <= not(layer3_outputs(1147)) or (layer3_outputs(4605));
    layer4_outputs(2617) <= not(layer3_outputs(3490));
    layer4_outputs(2618) <= not((layer3_outputs(2807)) and (layer3_outputs(4227)));
    layer4_outputs(2619) <= layer3_outputs(4174);
    layer4_outputs(2620) <= (layer3_outputs(3304)) and not (layer3_outputs(4141));
    layer4_outputs(2621) <= not(layer3_outputs(3673));
    layer4_outputs(2622) <= layer3_outputs(742);
    layer4_outputs(2623) <= layer3_outputs(327);
    layer4_outputs(2624) <= '1';
    layer4_outputs(2625) <= (layer3_outputs(4077)) and not (layer3_outputs(1964));
    layer4_outputs(2626) <= not((layer3_outputs(4124)) xor (layer3_outputs(4288)));
    layer4_outputs(2627) <= not(layer3_outputs(4678));
    layer4_outputs(2628) <= not(layer3_outputs(1760)) or (layer3_outputs(918));
    layer4_outputs(2629) <= not((layer3_outputs(3511)) or (layer3_outputs(1549)));
    layer4_outputs(2630) <= not((layer3_outputs(955)) or (layer3_outputs(2949)));
    layer4_outputs(2631) <= not(layer3_outputs(4297));
    layer4_outputs(2632) <= '0';
    layer4_outputs(2633) <= not(layer3_outputs(4129));
    layer4_outputs(2634) <= not(layer3_outputs(4640));
    layer4_outputs(2635) <= (layer3_outputs(1695)) xor (layer3_outputs(3902));
    layer4_outputs(2636) <= not((layer3_outputs(837)) or (layer3_outputs(159)));
    layer4_outputs(2637) <= not(layer3_outputs(317));
    layer4_outputs(2638) <= (layer3_outputs(2376)) and not (layer3_outputs(2341));
    layer4_outputs(2639) <= layer3_outputs(1447);
    layer4_outputs(2640) <= '0';
    layer4_outputs(2641) <= not((layer3_outputs(2641)) xor (layer3_outputs(3548)));
    layer4_outputs(2642) <= layer3_outputs(3968);
    layer4_outputs(2643) <= not(layer3_outputs(1732));
    layer4_outputs(2644) <= not(layer3_outputs(2446));
    layer4_outputs(2645) <= layer3_outputs(4393);
    layer4_outputs(2646) <= not(layer3_outputs(4599));
    layer4_outputs(2647) <= (layer3_outputs(4493)) xor (layer3_outputs(4268));
    layer4_outputs(2648) <= layer3_outputs(3632);
    layer4_outputs(2649) <= not(layer3_outputs(1626));
    layer4_outputs(2650) <= not(layer3_outputs(3718));
    layer4_outputs(2651) <= layer3_outputs(3557);
    layer4_outputs(2652) <= not(layer3_outputs(1801));
    layer4_outputs(2653) <= (layer3_outputs(3006)) and not (layer3_outputs(2596));
    layer4_outputs(2654) <= layer3_outputs(3760);
    layer4_outputs(2655) <= layer3_outputs(3739);
    layer4_outputs(2656) <= not(layer3_outputs(4403));
    layer4_outputs(2657) <= not(layer3_outputs(592));
    layer4_outputs(2658) <= not((layer3_outputs(1531)) xor (layer3_outputs(5087)));
    layer4_outputs(2659) <= not(layer3_outputs(1994));
    layer4_outputs(2660) <= not(layer3_outputs(3056));
    layer4_outputs(2661) <= (layer3_outputs(1901)) and not (layer3_outputs(5012));
    layer4_outputs(2662) <= not(layer3_outputs(274)) or (layer3_outputs(2386));
    layer4_outputs(2663) <= (layer3_outputs(2030)) and not (layer3_outputs(2138));
    layer4_outputs(2664) <= not(layer3_outputs(2620));
    layer4_outputs(2665) <= not(layer3_outputs(2892)) or (layer3_outputs(2876));
    layer4_outputs(2666) <= not((layer3_outputs(1343)) and (layer3_outputs(1551)));
    layer4_outputs(2667) <= not(layer3_outputs(3485));
    layer4_outputs(2668) <= not(layer3_outputs(4857));
    layer4_outputs(2669) <= not(layer3_outputs(502));
    layer4_outputs(2670) <= layer3_outputs(1881);
    layer4_outputs(2671) <= layer3_outputs(3869);
    layer4_outputs(2672) <= layer3_outputs(2772);
    layer4_outputs(2673) <= layer3_outputs(2786);
    layer4_outputs(2674) <= layer3_outputs(3082);
    layer4_outputs(2675) <= (layer3_outputs(3309)) and not (layer3_outputs(4098));
    layer4_outputs(2676) <= not(layer3_outputs(4345)) or (layer3_outputs(2386));
    layer4_outputs(2677) <= layer3_outputs(224);
    layer4_outputs(2678) <= not(layer3_outputs(1827));
    layer4_outputs(2679) <= not(layer3_outputs(3140)) or (layer3_outputs(4172));
    layer4_outputs(2680) <= layer3_outputs(324);
    layer4_outputs(2681) <= not(layer3_outputs(4703));
    layer4_outputs(2682) <= not(layer3_outputs(5013)) or (layer3_outputs(1674));
    layer4_outputs(2683) <= layer3_outputs(3014);
    layer4_outputs(2684) <= layer3_outputs(1974);
    layer4_outputs(2685) <= not(layer3_outputs(3802));
    layer4_outputs(2686) <= not((layer3_outputs(4517)) and (layer3_outputs(239)));
    layer4_outputs(2687) <= layer3_outputs(3952);
    layer4_outputs(2688) <= layer3_outputs(3477);
    layer4_outputs(2689) <= layer3_outputs(3116);
    layer4_outputs(2690) <= not(layer3_outputs(3103));
    layer4_outputs(2691) <= '1';
    layer4_outputs(2692) <= layer3_outputs(308);
    layer4_outputs(2693) <= not(layer3_outputs(1510)) or (layer3_outputs(2547));
    layer4_outputs(2694) <= not(layer3_outputs(4671));
    layer4_outputs(2695) <= (layer3_outputs(2818)) and not (layer3_outputs(841));
    layer4_outputs(2696) <= '0';
    layer4_outputs(2697) <= not(layer3_outputs(1158));
    layer4_outputs(2698) <= not(layer3_outputs(650)) or (layer3_outputs(1512));
    layer4_outputs(2699) <= layer3_outputs(2034);
    layer4_outputs(2700) <= (layer3_outputs(2420)) xor (layer3_outputs(4970));
    layer4_outputs(2701) <= (layer3_outputs(683)) and not (layer3_outputs(3837));
    layer4_outputs(2702) <= not(layer3_outputs(1220));
    layer4_outputs(2703) <= (layer3_outputs(3160)) and (layer3_outputs(512));
    layer4_outputs(2704) <= (layer3_outputs(2528)) and (layer3_outputs(1291));
    layer4_outputs(2705) <= (layer3_outputs(1811)) and not (layer3_outputs(1822));
    layer4_outputs(2706) <= (layer3_outputs(2401)) and not (layer3_outputs(3019));
    layer4_outputs(2707) <= (layer3_outputs(5009)) and (layer3_outputs(4754));
    layer4_outputs(2708) <= not(layer3_outputs(1846));
    layer4_outputs(2709) <= not((layer3_outputs(127)) or (layer3_outputs(3714)));
    layer4_outputs(2710) <= not(layer3_outputs(2942));
    layer4_outputs(2711) <= (layer3_outputs(3865)) and (layer3_outputs(3279));
    layer4_outputs(2712) <= '0';
    layer4_outputs(2713) <= '1';
    layer4_outputs(2714) <= layer3_outputs(1854);
    layer4_outputs(2715) <= (layer3_outputs(3992)) xor (layer3_outputs(3027));
    layer4_outputs(2716) <= not((layer3_outputs(1456)) or (layer3_outputs(3716)));
    layer4_outputs(2717) <= layer3_outputs(3395);
    layer4_outputs(2718) <= not(layer3_outputs(3229));
    layer4_outputs(2719) <= (layer3_outputs(4713)) and (layer3_outputs(1618));
    layer4_outputs(2720) <= (layer3_outputs(777)) xor (layer3_outputs(1568));
    layer4_outputs(2721) <= not(layer3_outputs(2769));
    layer4_outputs(2722) <= not(layer3_outputs(2022)) or (layer3_outputs(3953));
    layer4_outputs(2723) <= not(layer3_outputs(793));
    layer4_outputs(2724) <= layer3_outputs(303);
    layer4_outputs(2725) <= not((layer3_outputs(3985)) xor (layer3_outputs(2306)));
    layer4_outputs(2726) <= (layer3_outputs(3406)) or (layer3_outputs(565));
    layer4_outputs(2727) <= layer3_outputs(4642);
    layer4_outputs(2728) <= (layer3_outputs(4827)) or (layer3_outputs(5099));
    layer4_outputs(2729) <= layer3_outputs(1312);
    layer4_outputs(2730) <= '0';
    layer4_outputs(2731) <= (layer3_outputs(1903)) and (layer3_outputs(3613));
    layer4_outputs(2732) <= (layer3_outputs(3174)) xor (layer3_outputs(21));
    layer4_outputs(2733) <= not(layer3_outputs(3624)) or (layer3_outputs(4242));
    layer4_outputs(2734) <= layer3_outputs(4686);
    layer4_outputs(2735) <= not(layer3_outputs(1260));
    layer4_outputs(2736) <= not(layer3_outputs(2320));
    layer4_outputs(2737) <= not((layer3_outputs(4832)) or (layer3_outputs(1005)));
    layer4_outputs(2738) <= '1';
    layer4_outputs(2739) <= not(layer3_outputs(4811));
    layer4_outputs(2740) <= not(layer3_outputs(4192));
    layer4_outputs(2741) <= (layer3_outputs(3636)) and (layer3_outputs(147));
    layer4_outputs(2742) <= layer3_outputs(1553);
    layer4_outputs(2743) <= layer3_outputs(3579);
    layer4_outputs(2744) <= layer3_outputs(1099);
    layer4_outputs(2745) <= layer3_outputs(3735);
    layer4_outputs(2746) <= not(layer3_outputs(3053));
    layer4_outputs(2747) <= (layer3_outputs(602)) and not (layer3_outputs(4848));
    layer4_outputs(2748) <= not(layer3_outputs(4703));
    layer4_outputs(2749) <= not(layer3_outputs(1467)) or (layer3_outputs(2124));
    layer4_outputs(2750) <= '0';
    layer4_outputs(2751) <= (layer3_outputs(4890)) and not (layer3_outputs(2518));
    layer4_outputs(2752) <= layer3_outputs(2462);
    layer4_outputs(2753) <= (layer3_outputs(1091)) and (layer3_outputs(4163));
    layer4_outputs(2754) <= layer3_outputs(3276);
    layer4_outputs(2755) <= (layer3_outputs(3729)) and not (layer3_outputs(531));
    layer4_outputs(2756) <= not(layer3_outputs(371));
    layer4_outputs(2757) <= (layer3_outputs(2957)) and (layer3_outputs(4208));
    layer4_outputs(2758) <= not(layer3_outputs(2297)) or (layer3_outputs(375));
    layer4_outputs(2759) <= not((layer3_outputs(2359)) and (layer3_outputs(4494)));
    layer4_outputs(2760) <= (layer3_outputs(203)) and not (layer3_outputs(1866));
    layer4_outputs(2761) <= not(layer3_outputs(880));
    layer4_outputs(2762) <= (layer3_outputs(5089)) and (layer3_outputs(1676));
    layer4_outputs(2763) <= not(layer3_outputs(2816)) or (layer3_outputs(4912));
    layer4_outputs(2764) <= not((layer3_outputs(294)) and (layer3_outputs(2414)));
    layer4_outputs(2765) <= (layer3_outputs(4810)) and (layer3_outputs(3972));
    layer4_outputs(2766) <= layer3_outputs(4829);
    layer4_outputs(2767) <= (layer3_outputs(446)) xor (layer3_outputs(4640));
    layer4_outputs(2768) <= (layer3_outputs(2169)) or (layer3_outputs(2294));
    layer4_outputs(2769) <= (layer3_outputs(4993)) and (layer3_outputs(814));
    layer4_outputs(2770) <= layer3_outputs(4369);
    layer4_outputs(2771) <= (layer3_outputs(2840)) and not (layer3_outputs(3106));
    layer4_outputs(2772) <= not((layer3_outputs(4644)) and (layer3_outputs(236)));
    layer4_outputs(2773) <= not((layer3_outputs(589)) and (layer3_outputs(3872)));
    layer4_outputs(2774) <= not(layer3_outputs(336)) or (layer3_outputs(786));
    layer4_outputs(2775) <= (layer3_outputs(5006)) and not (layer3_outputs(3467));
    layer4_outputs(2776) <= '0';
    layer4_outputs(2777) <= not(layer3_outputs(2225)) or (layer3_outputs(3497));
    layer4_outputs(2778) <= layer3_outputs(761);
    layer4_outputs(2779) <= '1';
    layer4_outputs(2780) <= (layer3_outputs(3905)) or (layer3_outputs(3242));
    layer4_outputs(2781) <= '1';
    layer4_outputs(2782) <= (layer3_outputs(2691)) and (layer3_outputs(1930));
    layer4_outputs(2783) <= not(layer3_outputs(3085));
    layer4_outputs(2784) <= not(layer3_outputs(4510));
    layer4_outputs(2785) <= (layer3_outputs(4362)) and not (layer3_outputs(1902));
    layer4_outputs(2786) <= not(layer3_outputs(4936));
    layer4_outputs(2787) <= not((layer3_outputs(2689)) or (layer3_outputs(4707)));
    layer4_outputs(2788) <= layer3_outputs(2631);
    layer4_outputs(2789) <= '1';
    layer4_outputs(2790) <= not((layer3_outputs(2347)) and (layer3_outputs(4843)));
    layer4_outputs(2791) <= layer3_outputs(1907);
    layer4_outputs(2792) <= not((layer3_outputs(3899)) or (layer3_outputs(3448)));
    layer4_outputs(2793) <= layer3_outputs(3662);
    layer4_outputs(2794) <= '0';
    layer4_outputs(2795) <= not(layer3_outputs(4998));
    layer4_outputs(2796) <= (layer3_outputs(4049)) and not (layer3_outputs(2615));
    layer4_outputs(2797) <= not((layer3_outputs(2853)) xor (layer3_outputs(3420)));
    layer4_outputs(2798) <= not(layer3_outputs(4722)) or (layer3_outputs(3887));
    layer4_outputs(2799) <= layer3_outputs(545);
    layer4_outputs(2800) <= layer3_outputs(1529);
    layer4_outputs(2801) <= not((layer3_outputs(833)) xor (layer3_outputs(3461)));
    layer4_outputs(2802) <= (layer3_outputs(433)) and not (layer3_outputs(1356));
    layer4_outputs(2803) <= not(layer3_outputs(2989));
    layer4_outputs(2804) <= not((layer3_outputs(4635)) and (layer3_outputs(3592)));
    layer4_outputs(2805) <= (layer3_outputs(2029)) xor (layer3_outputs(4766));
    layer4_outputs(2806) <= layer3_outputs(2344);
    layer4_outputs(2807) <= not(layer3_outputs(3584));
    layer4_outputs(2808) <= not(layer3_outputs(4983));
    layer4_outputs(2809) <= (layer3_outputs(5111)) and not (layer3_outputs(3750));
    layer4_outputs(2810) <= not(layer3_outputs(4536)) or (layer3_outputs(3438));
    layer4_outputs(2811) <= (layer3_outputs(2153)) and (layer3_outputs(2253));
    layer4_outputs(2812) <= not(layer3_outputs(2788));
    layer4_outputs(2813) <= not((layer3_outputs(3738)) xor (layer3_outputs(839)));
    layer4_outputs(2814) <= not(layer3_outputs(4084)) or (layer3_outputs(3072));
    layer4_outputs(2815) <= not(layer3_outputs(469));
    layer4_outputs(2816) <= (layer3_outputs(3685)) xor (layer3_outputs(182));
    layer4_outputs(2817) <= not((layer3_outputs(1783)) and (layer3_outputs(3661)));
    layer4_outputs(2818) <= layer3_outputs(4094);
    layer4_outputs(2819) <= layer3_outputs(89);
    layer4_outputs(2820) <= layer3_outputs(1149);
    layer4_outputs(2821) <= (layer3_outputs(4669)) and (layer3_outputs(1173));
    layer4_outputs(2822) <= not(layer3_outputs(3437));
    layer4_outputs(2823) <= layer3_outputs(2635);
    layer4_outputs(2824) <= '0';
    layer4_outputs(2825) <= not((layer3_outputs(221)) or (layer3_outputs(2239)));
    layer4_outputs(2826) <= layer3_outputs(912);
    layer4_outputs(2827) <= '1';
    layer4_outputs(2828) <= not((layer3_outputs(998)) xor (layer3_outputs(1793)));
    layer4_outputs(2829) <= (layer3_outputs(4794)) and (layer3_outputs(219));
    layer4_outputs(2830) <= layer3_outputs(3532);
    layer4_outputs(2831) <= not((layer3_outputs(5021)) and (layer3_outputs(2536)));
    layer4_outputs(2832) <= (layer3_outputs(852)) and not (layer3_outputs(3251));
    layer4_outputs(2833) <= layer3_outputs(1519);
    layer4_outputs(2834) <= not((layer3_outputs(4095)) or (layer3_outputs(3850)));
    layer4_outputs(2835) <= layer3_outputs(4695);
    layer4_outputs(2836) <= (layer3_outputs(3982)) or (layer3_outputs(3746));
    layer4_outputs(2837) <= layer3_outputs(4883);
    layer4_outputs(2838) <= layer3_outputs(2879);
    layer4_outputs(2839) <= '0';
    layer4_outputs(2840) <= not((layer3_outputs(1712)) or (layer3_outputs(1914)));
    layer4_outputs(2841) <= '0';
    layer4_outputs(2842) <= not((layer3_outputs(824)) xor (layer3_outputs(1092)));
    layer4_outputs(2843) <= not(layer3_outputs(4229));
    layer4_outputs(2844) <= not(layer3_outputs(3904)) or (layer3_outputs(1590));
    layer4_outputs(2845) <= (layer3_outputs(832)) and (layer3_outputs(1630));
    layer4_outputs(2846) <= (layer3_outputs(1765)) or (layer3_outputs(2990));
    layer4_outputs(2847) <= '0';
    layer4_outputs(2848) <= layer3_outputs(1177);
    layer4_outputs(2849) <= (layer3_outputs(2791)) or (layer3_outputs(4566));
    layer4_outputs(2850) <= not(layer3_outputs(3251)) or (layer3_outputs(2628));
    layer4_outputs(2851) <= '0';
    layer4_outputs(2852) <= not((layer3_outputs(1401)) or (layer3_outputs(4313)));
    layer4_outputs(2853) <= '0';
    layer4_outputs(2854) <= layer3_outputs(4472);
    layer4_outputs(2855) <= not(layer3_outputs(3794)) or (layer3_outputs(3129));
    layer4_outputs(2856) <= not((layer3_outputs(1104)) and (layer3_outputs(1566)));
    layer4_outputs(2857) <= '0';
    layer4_outputs(2858) <= layer3_outputs(3566);
    layer4_outputs(2859) <= not(layer3_outputs(2700));
    layer4_outputs(2860) <= (layer3_outputs(2309)) or (layer3_outputs(2537));
    layer4_outputs(2861) <= layer3_outputs(812);
    layer4_outputs(2862) <= (layer3_outputs(2756)) and not (layer3_outputs(1822));
    layer4_outputs(2863) <= not(layer3_outputs(4528));
    layer4_outputs(2864) <= layer3_outputs(2237);
    layer4_outputs(2865) <= not(layer3_outputs(4324));
    layer4_outputs(2866) <= not((layer3_outputs(291)) and (layer3_outputs(2070)));
    layer4_outputs(2867) <= '0';
    layer4_outputs(2868) <= (layer3_outputs(3935)) and not (layer3_outputs(1389));
    layer4_outputs(2869) <= (layer3_outputs(4184)) and (layer3_outputs(2758));
    layer4_outputs(2870) <= (layer3_outputs(2608)) and not (layer3_outputs(4154));
    layer4_outputs(2871) <= not(layer3_outputs(1402));
    layer4_outputs(2872) <= not(layer3_outputs(807)) or (layer3_outputs(697));
    layer4_outputs(2873) <= not(layer3_outputs(1373)) or (layer3_outputs(240));
    layer4_outputs(2874) <= not((layer3_outputs(1335)) xor (layer3_outputs(1917)));
    layer4_outputs(2875) <= not((layer3_outputs(4292)) xor (layer3_outputs(852)));
    layer4_outputs(2876) <= not(layer3_outputs(2078));
    layer4_outputs(2877) <= not(layer3_outputs(2642));
    layer4_outputs(2878) <= '0';
    layer4_outputs(2879) <= not((layer3_outputs(1889)) xor (layer3_outputs(483)));
    layer4_outputs(2880) <= not(layer3_outputs(3890)) or (layer3_outputs(1809));
    layer4_outputs(2881) <= (layer3_outputs(767)) and not (layer3_outputs(2294));
    layer4_outputs(2882) <= not(layer3_outputs(4133));
    layer4_outputs(2883) <= (layer3_outputs(2117)) or (layer3_outputs(2469));
    layer4_outputs(2884) <= not(layer3_outputs(1973));
    layer4_outputs(2885) <= not((layer3_outputs(4666)) and (layer3_outputs(5053)));
    layer4_outputs(2886) <= (layer3_outputs(285)) xor (layer3_outputs(4832));
    layer4_outputs(2887) <= not(layer3_outputs(640));
    layer4_outputs(2888) <= (layer3_outputs(4042)) or (layer3_outputs(4345));
    layer4_outputs(2889) <= (layer3_outputs(1995)) and not (layer3_outputs(2439));
    layer4_outputs(2890) <= (layer3_outputs(1707)) and not (layer3_outputs(2426));
    layer4_outputs(2891) <= (layer3_outputs(3130)) and not (layer3_outputs(2243));
    layer4_outputs(2892) <= (layer3_outputs(3690)) and (layer3_outputs(3707));
    layer4_outputs(2893) <= not(layer3_outputs(2065));
    layer4_outputs(2894) <= not(layer3_outputs(3615));
    layer4_outputs(2895) <= not((layer3_outputs(4407)) or (layer3_outputs(1198)));
    layer4_outputs(2896) <= not(layer3_outputs(4926));
    layer4_outputs(2897) <= layer3_outputs(5091);
    layer4_outputs(2898) <= not(layer3_outputs(1325));
    layer4_outputs(2899) <= layer3_outputs(4024);
    layer4_outputs(2900) <= not(layer3_outputs(1952));
    layer4_outputs(2901) <= (layer3_outputs(3763)) and not (layer3_outputs(2852));
    layer4_outputs(2902) <= (layer3_outputs(3529)) or (layer3_outputs(1857));
    layer4_outputs(2903) <= (layer3_outputs(3473)) or (layer3_outputs(1138));
    layer4_outputs(2904) <= layer3_outputs(2507);
    layer4_outputs(2905) <= not(layer3_outputs(789));
    layer4_outputs(2906) <= not(layer3_outputs(1011));
    layer4_outputs(2907) <= not(layer3_outputs(477)) or (layer3_outputs(3198));
    layer4_outputs(2908) <= not(layer3_outputs(4400)) or (layer3_outputs(2916));
    layer4_outputs(2909) <= '0';
    layer4_outputs(2910) <= not(layer3_outputs(3023));
    layer4_outputs(2911) <= not((layer3_outputs(1214)) or (layer3_outputs(536)));
    layer4_outputs(2912) <= layer3_outputs(2353);
    layer4_outputs(2913) <= (layer3_outputs(1993)) xor (layer3_outputs(2516));
    layer4_outputs(2914) <= not(layer3_outputs(3003));
    layer4_outputs(2915) <= layer3_outputs(2297);
    layer4_outputs(2916) <= not((layer3_outputs(3818)) or (layer3_outputs(3674)));
    layer4_outputs(2917) <= not(layer3_outputs(4370)) or (layer3_outputs(3308));
    layer4_outputs(2918) <= layer3_outputs(3008);
    layer4_outputs(2919) <= '1';
    layer4_outputs(2920) <= '0';
    layer4_outputs(2921) <= layer3_outputs(3086);
    layer4_outputs(2922) <= '0';
    layer4_outputs(2923) <= (layer3_outputs(3316)) and (layer3_outputs(4941));
    layer4_outputs(2924) <= (layer3_outputs(4120)) and (layer3_outputs(2394));
    layer4_outputs(2925) <= (layer3_outputs(1722)) or (layer3_outputs(2053));
    layer4_outputs(2926) <= not((layer3_outputs(3052)) or (layer3_outputs(3266)));
    layer4_outputs(2927) <= not(layer3_outputs(2440)) or (layer3_outputs(4549));
    layer4_outputs(2928) <= layer3_outputs(4773);
    layer4_outputs(2929) <= '0';
    layer4_outputs(2930) <= (layer3_outputs(4948)) or (layer3_outputs(1640));
    layer4_outputs(2931) <= not(layer3_outputs(1711));
    layer4_outputs(2932) <= (layer3_outputs(3374)) and not (layer3_outputs(3969));
    layer4_outputs(2933) <= not((layer3_outputs(4979)) xor (layer3_outputs(4624)));
    layer4_outputs(2934) <= layer3_outputs(4463);
    layer4_outputs(2935) <= '1';
    layer4_outputs(2936) <= not((layer3_outputs(3708)) and (layer3_outputs(3993)));
    layer4_outputs(2937) <= not(layer3_outputs(3699));
    layer4_outputs(2938) <= '0';
    layer4_outputs(2939) <= not((layer3_outputs(2980)) or (layer3_outputs(2421)));
    layer4_outputs(2940) <= layer3_outputs(3451);
    layer4_outputs(2941) <= (layer3_outputs(3046)) and not (layer3_outputs(3627));
    layer4_outputs(2942) <= (layer3_outputs(1323)) and not (layer3_outputs(472));
    layer4_outputs(2943) <= not((layer3_outputs(4353)) and (layer3_outputs(1923)));
    layer4_outputs(2944) <= layer3_outputs(4620);
    layer4_outputs(2945) <= not(layer3_outputs(3924));
    layer4_outputs(2946) <= not(layer3_outputs(719));
    layer4_outputs(2947) <= not((layer3_outputs(677)) or (layer3_outputs(4989)));
    layer4_outputs(2948) <= layer3_outputs(1084);
    layer4_outputs(2949) <= not((layer3_outputs(846)) or (layer3_outputs(3916)));
    layer4_outputs(2950) <= (layer3_outputs(1633)) and not (layer3_outputs(2080));
    layer4_outputs(2951) <= not(layer3_outputs(4387));
    layer4_outputs(2952) <= '0';
    layer4_outputs(2953) <= layer3_outputs(3226);
    layer4_outputs(2954) <= (layer3_outputs(496)) and not (layer3_outputs(2877));
    layer4_outputs(2955) <= layer3_outputs(2444);
    layer4_outputs(2956) <= not(layer3_outputs(2177)) or (layer3_outputs(64));
    layer4_outputs(2957) <= layer3_outputs(3939);
    layer4_outputs(2958) <= not(layer3_outputs(4278));
    layer4_outputs(2959) <= layer3_outputs(3028);
    layer4_outputs(2960) <= '0';
    layer4_outputs(2961) <= not(layer3_outputs(5050));
    layer4_outputs(2962) <= (layer3_outputs(3329)) and not (layer3_outputs(170));
    layer4_outputs(2963) <= layer3_outputs(3388);
    layer4_outputs(2964) <= '0';
    layer4_outputs(2965) <= not(layer3_outputs(3459)) or (layer3_outputs(2332));
    layer4_outputs(2966) <= '1';
    layer4_outputs(2967) <= (layer3_outputs(3539)) and (layer3_outputs(1814));
    layer4_outputs(2968) <= '1';
    layer4_outputs(2969) <= layer3_outputs(1831);
    layer4_outputs(2970) <= not(layer3_outputs(2011));
    layer4_outputs(2971) <= layer3_outputs(1572);
    layer4_outputs(2972) <= (layer3_outputs(911)) and not (layer3_outputs(1481));
    layer4_outputs(2973) <= layer3_outputs(2026);
    layer4_outputs(2974) <= (layer3_outputs(1161)) and not (layer3_outputs(4706));
    layer4_outputs(2975) <= not(layer3_outputs(405)) or (layer3_outputs(3134));
    layer4_outputs(2976) <= not((layer3_outputs(4670)) and (layer3_outputs(4630)));
    layer4_outputs(2977) <= (layer3_outputs(2713)) xor (layer3_outputs(4997));
    layer4_outputs(2978) <= (layer3_outputs(4261)) and not (layer3_outputs(3582));
    layer4_outputs(2979) <= not((layer3_outputs(3363)) xor (layer3_outputs(3887)));
    layer4_outputs(2980) <= not((layer3_outputs(2897)) and (layer3_outputs(890)));
    layer4_outputs(2981) <= not(layer3_outputs(3688));
    layer4_outputs(2982) <= (layer3_outputs(4732)) and not (layer3_outputs(5104));
    layer4_outputs(2983) <= layer3_outputs(4192);
    layer4_outputs(2984) <= not(layer3_outputs(3222));
    layer4_outputs(2985) <= not(layer3_outputs(1247));
    layer4_outputs(2986) <= layer3_outputs(1378);
    layer4_outputs(2987) <= not(layer3_outputs(2048)) or (layer3_outputs(4318));
    layer4_outputs(2988) <= not((layer3_outputs(4352)) and (layer3_outputs(840)));
    layer4_outputs(2989) <= (layer3_outputs(1048)) and not (layer3_outputs(4485));
    layer4_outputs(2990) <= not(layer3_outputs(4220)) or (layer3_outputs(2956));
    layer4_outputs(2991) <= layer3_outputs(3903);
    layer4_outputs(2992) <= layer3_outputs(1418);
    layer4_outputs(2993) <= (layer3_outputs(2227)) xor (layer3_outputs(4752));
    layer4_outputs(2994) <= layer3_outputs(1746);
    layer4_outputs(2995) <= not(layer3_outputs(881));
    layer4_outputs(2996) <= layer3_outputs(693);
    layer4_outputs(2997) <= not(layer3_outputs(4410));
    layer4_outputs(2998) <= layer3_outputs(4783);
    layer4_outputs(2999) <= not((layer3_outputs(1838)) xor (layer3_outputs(2363)));
    layer4_outputs(3000) <= layer3_outputs(2964);
    layer4_outputs(3001) <= not(layer3_outputs(2724));
    layer4_outputs(3002) <= (layer3_outputs(4723)) or (layer3_outputs(2840));
    layer4_outputs(3003) <= not(layer3_outputs(4372));
    layer4_outputs(3004) <= layer3_outputs(4333);
    layer4_outputs(3005) <= (layer3_outputs(1144)) and not (layer3_outputs(1209));
    layer4_outputs(3006) <= layer3_outputs(3742);
    layer4_outputs(3007) <= layer3_outputs(1080);
    layer4_outputs(3008) <= not(layer3_outputs(3418));
    layer4_outputs(3009) <= (layer3_outputs(3803)) and (layer3_outputs(1009));
    layer4_outputs(3010) <= (layer3_outputs(1933)) and (layer3_outputs(2870));
    layer4_outputs(3011) <= not((layer3_outputs(5063)) or (layer3_outputs(5097)));
    layer4_outputs(3012) <= (layer3_outputs(2401)) xor (layer3_outputs(1413));
    layer4_outputs(3013) <= (layer3_outputs(1838)) and (layer3_outputs(2784));
    layer4_outputs(3014) <= '1';
    layer4_outputs(3015) <= (layer3_outputs(6)) and (layer3_outputs(1123));
    layer4_outputs(3016) <= (layer3_outputs(612)) xor (layer3_outputs(3458));
    layer4_outputs(3017) <= not(layer3_outputs(726));
    layer4_outputs(3018) <= not(layer3_outputs(41));
    layer4_outputs(3019) <= layer3_outputs(946);
    layer4_outputs(3020) <= '1';
    layer4_outputs(3021) <= '0';
    layer4_outputs(3022) <= (layer3_outputs(4975)) and not (layer3_outputs(4467));
    layer4_outputs(3023) <= layer3_outputs(3439);
    layer4_outputs(3024) <= not(layer3_outputs(1622)) or (layer3_outputs(2725));
    layer4_outputs(3025) <= layer3_outputs(4609);
    layer4_outputs(3026) <= layer3_outputs(1096);
    layer4_outputs(3027) <= not(layer3_outputs(2919));
    layer4_outputs(3028) <= not(layer3_outputs(3300));
    layer4_outputs(3029) <= '0';
    layer4_outputs(3030) <= not(layer3_outputs(4219));
    layer4_outputs(3031) <= not(layer3_outputs(1660));
    layer4_outputs(3032) <= (layer3_outputs(1230)) and (layer3_outputs(1072));
    layer4_outputs(3033) <= not(layer3_outputs(2244));
    layer4_outputs(3034) <= not((layer3_outputs(2341)) or (layer3_outputs(4349)));
    layer4_outputs(3035) <= layer3_outputs(3917);
    layer4_outputs(3036) <= not((layer3_outputs(2348)) and (layer3_outputs(1366)));
    layer4_outputs(3037) <= not((layer3_outputs(3285)) or (layer3_outputs(2696)));
    layer4_outputs(3038) <= not(layer3_outputs(3457)) or (layer3_outputs(3468));
    layer4_outputs(3039) <= layer3_outputs(555);
    layer4_outputs(3040) <= not(layer3_outputs(3925)) or (layer3_outputs(126));
    layer4_outputs(3041) <= not(layer3_outputs(1336)) or (layer3_outputs(243));
    layer4_outputs(3042) <= (layer3_outputs(2362)) and not (layer3_outputs(146));
    layer4_outputs(3043) <= layer3_outputs(4945);
    layer4_outputs(3044) <= '0';
    layer4_outputs(3045) <= not((layer3_outputs(3303)) and (layer3_outputs(207)));
    layer4_outputs(3046) <= '1';
    layer4_outputs(3047) <= (layer3_outputs(1041)) and not (layer3_outputs(3865));
    layer4_outputs(3048) <= not((layer3_outputs(4694)) and (layer3_outputs(3156)));
    layer4_outputs(3049) <= (layer3_outputs(2112)) and not (layer3_outputs(4409));
    layer4_outputs(3050) <= not(layer3_outputs(726));
    layer4_outputs(3051) <= not(layer3_outputs(2333)) or (layer3_outputs(5085));
    layer4_outputs(3052) <= not(layer3_outputs(2996));
    layer4_outputs(3053) <= (layer3_outputs(4413)) or (layer3_outputs(3627));
    layer4_outputs(3054) <= (layer3_outputs(1725)) xor (layer3_outputs(1400));
    layer4_outputs(3055) <= not(layer3_outputs(3545));
    layer4_outputs(3056) <= (layer3_outputs(4855)) and (layer3_outputs(4645));
    layer4_outputs(3057) <= (layer3_outputs(1931)) or (layer3_outputs(1379));
    layer4_outputs(3058) <= not(layer3_outputs(1085));
    layer4_outputs(3059) <= not(layer3_outputs(3416));
    layer4_outputs(3060) <= (layer3_outputs(418)) and (layer3_outputs(3670));
    layer4_outputs(3061) <= (layer3_outputs(2371)) and not (layer3_outputs(2934));
    layer4_outputs(3062) <= (layer3_outputs(2661)) and (layer3_outputs(2648));
    layer4_outputs(3063) <= (layer3_outputs(999)) and not (layer3_outputs(765));
    layer4_outputs(3064) <= layer3_outputs(3307);
    layer4_outputs(3065) <= not(layer3_outputs(1351));
    layer4_outputs(3066) <= not(layer3_outputs(739));
    layer4_outputs(3067) <= (layer3_outputs(4826)) and not (layer3_outputs(855));
    layer4_outputs(3068) <= '0';
    layer4_outputs(3069) <= (layer3_outputs(4729)) or (layer3_outputs(4072));
    layer4_outputs(3070) <= not(layer3_outputs(3402));
    layer4_outputs(3071) <= (layer3_outputs(4244)) or (layer3_outputs(601));
    layer4_outputs(3072) <= not(layer3_outputs(3077));
    layer4_outputs(3073) <= layer3_outputs(519);
    layer4_outputs(3074) <= layer3_outputs(1363);
    layer4_outputs(3075) <= not(layer3_outputs(1138));
    layer4_outputs(3076) <= (layer3_outputs(3096)) and not (layer3_outputs(962));
    layer4_outputs(3077) <= layer3_outputs(2139);
    layer4_outputs(3078) <= not(layer3_outputs(476)) or (layer3_outputs(3884));
    layer4_outputs(3079) <= (layer3_outputs(2019)) and not (layer3_outputs(2041));
    layer4_outputs(3080) <= not(layer3_outputs(3603));
    layer4_outputs(3081) <= layer3_outputs(1262);
    layer4_outputs(3082) <= (layer3_outputs(3838)) xor (layer3_outputs(2381));
    layer4_outputs(3083) <= '0';
    layer4_outputs(3084) <= not(layer3_outputs(1532)) or (layer3_outputs(2677));
    layer4_outputs(3085) <= not(layer3_outputs(1297)) or (layer3_outputs(3878));
    layer4_outputs(3086) <= not(layer3_outputs(4409));
    layer4_outputs(3087) <= '0';
    layer4_outputs(3088) <= not(layer3_outputs(3138));
    layer4_outputs(3089) <= (layer3_outputs(242)) or (layer3_outputs(3315));
    layer4_outputs(3090) <= not(layer3_outputs(4488));
    layer4_outputs(3091) <= not((layer3_outputs(2575)) or (layer3_outputs(4456)));
    layer4_outputs(3092) <= layer3_outputs(458);
    layer4_outputs(3093) <= not(layer3_outputs(4051));
    layer4_outputs(3094) <= not(layer3_outputs(178));
    layer4_outputs(3095) <= (layer3_outputs(1945)) and not (layer3_outputs(4330));
    layer4_outputs(3096) <= not(layer3_outputs(3941)) or (layer3_outputs(1226));
    layer4_outputs(3097) <= not(layer3_outputs(4579));
    layer4_outputs(3098) <= not(layer3_outputs(2819)) or (layer3_outputs(2171));
    layer4_outputs(3099) <= not(layer3_outputs(587)) or (layer3_outputs(4772));
    layer4_outputs(3100) <= layer3_outputs(5054);
    layer4_outputs(3101) <= not((layer3_outputs(4861)) and (layer3_outputs(2915)));
    layer4_outputs(3102) <= not((layer3_outputs(801)) and (layer3_outputs(932)));
    layer4_outputs(3103) <= not(layer3_outputs(3597));
    layer4_outputs(3104) <= not((layer3_outputs(2694)) or (layer3_outputs(4613)));
    layer4_outputs(3105) <= layer3_outputs(1539);
    layer4_outputs(3106) <= not(layer3_outputs(2774));
    layer4_outputs(3107) <= layer3_outputs(330);
    layer4_outputs(3108) <= '1';
    layer4_outputs(3109) <= (layer3_outputs(2710)) xor (layer3_outputs(993));
    layer4_outputs(3110) <= layer3_outputs(1878);
    layer4_outputs(3111) <= (layer3_outputs(4066)) or (layer3_outputs(328));
    layer4_outputs(3112) <= not(layer3_outputs(1195)) or (layer3_outputs(1305));
    layer4_outputs(3113) <= not(layer3_outputs(2099)) or (layer3_outputs(734));
    layer4_outputs(3114) <= not((layer3_outputs(1484)) or (layer3_outputs(3650)));
    layer4_outputs(3115) <= '0';
    layer4_outputs(3116) <= not((layer3_outputs(1428)) xor (layer3_outputs(3880)));
    layer4_outputs(3117) <= not(layer3_outputs(923));
    layer4_outputs(3118) <= (layer3_outputs(1093)) and not (layer3_outputs(321));
    layer4_outputs(3119) <= layer3_outputs(3715);
    layer4_outputs(3120) <= not(layer3_outputs(2362)) or (layer3_outputs(104));
    layer4_outputs(3121) <= (layer3_outputs(1786)) and (layer3_outputs(2962));
    layer4_outputs(3122) <= (layer3_outputs(132)) and (layer3_outputs(1572));
    layer4_outputs(3123) <= (layer3_outputs(241)) and not (layer3_outputs(2421));
    layer4_outputs(3124) <= not(layer3_outputs(1833));
    layer4_outputs(3125) <= not(layer3_outputs(2072));
    layer4_outputs(3126) <= not(layer3_outputs(3623));
    layer4_outputs(3127) <= layer3_outputs(1209);
    layer4_outputs(3128) <= not(layer3_outputs(894)) or (layer3_outputs(3798));
    layer4_outputs(3129) <= layer3_outputs(939);
    layer4_outputs(3130) <= not(layer3_outputs(4931)) or (layer3_outputs(5046));
    layer4_outputs(3131) <= (layer3_outputs(3976)) or (layer3_outputs(3980));
    layer4_outputs(3132) <= (layer3_outputs(822)) or (layer3_outputs(4462));
    layer4_outputs(3133) <= not(layer3_outputs(2377)) or (layer3_outputs(1654));
    layer4_outputs(3134) <= not(layer3_outputs(467));
    layer4_outputs(3135) <= not(layer3_outputs(2116));
    layer4_outputs(3136) <= (layer3_outputs(277)) and not (layer3_outputs(4769));
    layer4_outputs(3137) <= layer3_outputs(2611);
    layer4_outputs(3138) <= not(layer3_outputs(1056));
    layer4_outputs(3139) <= layer3_outputs(3094);
    layer4_outputs(3140) <= not((layer3_outputs(2170)) xor (layer3_outputs(1397)));
    layer4_outputs(3141) <= not((layer3_outputs(3296)) and (layer3_outputs(1289)));
    layer4_outputs(3142) <= not(layer3_outputs(431));
    layer4_outputs(3143) <= layer3_outputs(2625);
    layer4_outputs(3144) <= not(layer3_outputs(2032)) or (layer3_outputs(275));
    layer4_outputs(3145) <= not(layer3_outputs(1867));
    layer4_outputs(3146) <= not((layer3_outputs(1792)) or (layer3_outputs(840)));
    layer4_outputs(3147) <= not(layer3_outputs(810));
    layer4_outputs(3148) <= (layer3_outputs(3746)) xor (layer3_outputs(1107));
    layer4_outputs(3149) <= not(layer3_outputs(4741)) or (layer3_outputs(3144));
    layer4_outputs(3150) <= (layer3_outputs(2662)) or (layer3_outputs(2329));
    layer4_outputs(3151) <= not(layer3_outputs(218));
    layer4_outputs(3152) <= '1';
    layer4_outputs(3153) <= '1';
    layer4_outputs(3154) <= (layer3_outputs(1969)) and not (layer3_outputs(3599));
    layer4_outputs(3155) <= layer3_outputs(3620);
    layer4_outputs(3156) <= not((layer3_outputs(4564)) or (layer3_outputs(1287)));
    layer4_outputs(3157) <= layer3_outputs(4359);
    layer4_outputs(3158) <= not(layer3_outputs(2452)) or (layer3_outputs(599));
    layer4_outputs(3159) <= not(layer3_outputs(3908));
    layer4_outputs(3160) <= (layer3_outputs(2721)) or (layer3_outputs(2578));
    layer4_outputs(3161) <= not(layer3_outputs(4856));
    layer4_outputs(3162) <= (layer3_outputs(377)) and not (layer3_outputs(4453));
    layer4_outputs(3163) <= (layer3_outputs(3460)) or (layer3_outputs(4914));
    layer4_outputs(3164) <= not((layer3_outputs(988)) and (layer3_outputs(2572)));
    layer4_outputs(3165) <= layer3_outputs(629);
    layer4_outputs(3166) <= not(layer3_outputs(462)) or (layer3_outputs(2955));
    layer4_outputs(3167) <= not(layer3_outputs(3177));
    layer4_outputs(3168) <= layer3_outputs(2782);
    layer4_outputs(3169) <= (layer3_outputs(1820)) and not (layer3_outputs(3041));
    layer4_outputs(3170) <= not(layer3_outputs(123));
    layer4_outputs(3171) <= (layer3_outputs(1958)) and not (layer3_outputs(870));
    layer4_outputs(3172) <= not(layer3_outputs(1713));
    layer4_outputs(3173) <= not(layer3_outputs(4545));
    layer4_outputs(3174) <= not(layer3_outputs(1697));
    layer4_outputs(3175) <= not((layer3_outputs(1233)) or (layer3_outputs(2279)));
    layer4_outputs(3176) <= (layer3_outputs(3645)) and (layer3_outputs(2432));
    layer4_outputs(3177) <= not(layer3_outputs(2286));
    layer4_outputs(3178) <= not(layer3_outputs(1399)) or (layer3_outputs(5085));
    layer4_outputs(3179) <= layer3_outputs(1956);
    layer4_outputs(3180) <= not((layer3_outputs(2150)) or (layer3_outputs(1982)));
    layer4_outputs(3181) <= not(layer3_outputs(803));
    layer4_outputs(3182) <= layer3_outputs(5041);
    layer4_outputs(3183) <= (layer3_outputs(2456)) or (layer3_outputs(2183));
    layer4_outputs(3184) <= layer3_outputs(2462);
    layer4_outputs(3185) <= not(layer3_outputs(71));
    layer4_outputs(3186) <= layer3_outputs(3100);
    layer4_outputs(3187) <= not((layer3_outputs(2900)) or (layer3_outputs(4972)));
    layer4_outputs(3188) <= layer3_outputs(4744);
    layer4_outputs(3189) <= layer3_outputs(3328);
    layer4_outputs(3190) <= not(layer3_outputs(2514));
    layer4_outputs(3191) <= not((layer3_outputs(3273)) or (layer3_outputs(1413)));
    layer4_outputs(3192) <= not(layer3_outputs(4662)) or (layer3_outputs(2379));
    layer4_outputs(3193) <= not(layer3_outputs(285));
    layer4_outputs(3194) <= layer3_outputs(2885);
    layer4_outputs(3195) <= (layer3_outputs(2336)) and (layer3_outputs(276));
    layer4_outputs(3196) <= (layer3_outputs(3965)) and not (layer3_outputs(4880));
    layer4_outputs(3197) <= '1';
    layer4_outputs(3198) <= not(layer3_outputs(2167));
    layer4_outputs(3199) <= (layer3_outputs(4263)) and not (layer3_outputs(2670));
    layer4_outputs(3200) <= not((layer3_outputs(1485)) xor (layer3_outputs(1894)));
    layer4_outputs(3201) <= not(layer3_outputs(1035));
    layer4_outputs(3202) <= not(layer3_outputs(1169));
    layer4_outputs(3203) <= (layer3_outputs(1275)) xor (layer3_outputs(3791));
    layer4_outputs(3204) <= (layer3_outputs(4730)) and not (layer3_outputs(2947));
    layer4_outputs(3205) <= (layer3_outputs(1944)) and not (layer3_outputs(2089));
    layer4_outputs(3206) <= not(layer3_outputs(2963)) or (layer3_outputs(4403));
    layer4_outputs(3207) <= '0';
    layer4_outputs(3208) <= '0';
    layer4_outputs(3209) <= not(layer3_outputs(3115));
    layer4_outputs(3210) <= not(layer3_outputs(4458)) or (layer3_outputs(967));
    layer4_outputs(3211) <= (layer3_outputs(1525)) and (layer3_outputs(4661));
    layer4_outputs(3212) <= not(layer3_outputs(1076));
    layer4_outputs(3213) <= not(layer3_outputs(5048));
    layer4_outputs(3214) <= (layer3_outputs(1208)) and not (layer3_outputs(3254));
    layer4_outputs(3215) <= not(layer3_outputs(3926));
    layer4_outputs(3216) <= (layer3_outputs(4943)) and not (layer3_outputs(2366));
    layer4_outputs(3217) <= not(layer3_outputs(1656)) or (layer3_outputs(256));
    layer4_outputs(3218) <= (layer3_outputs(4005)) and (layer3_outputs(4756));
    layer4_outputs(3219) <= not((layer3_outputs(2202)) or (layer3_outputs(280)));
    layer4_outputs(3220) <= (layer3_outputs(2108)) and not (layer3_outputs(1277));
    layer4_outputs(3221) <= not(layer3_outputs(2040));
    layer4_outputs(3222) <= not((layer3_outputs(4570)) xor (layer3_outputs(3179)));
    layer4_outputs(3223) <= not(layer3_outputs(3789));
    layer4_outputs(3224) <= not((layer3_outputs(4436)) or (layer3_outputs(348)));
    layer4_outputs(3225) <= layer3_outputs(1684);
    layer4_outputs(3226) <= not((layer3_outputs(1552)) or (layer3_outputs(1816)));
    layer4_outputs(3227) <= (layer3_outputs(4332)) and not (layer3_outputs(2938));
    layer4_outputs(3228) <= not(layer3_outputs(4569));
    layer4_outputs(3229) <= not((layer3_outputs(2918)) or (layer3_outputs(3600)));
    layer4_outputs(3230) <= not(layer3_outputs(141));
    layer4_outputs(3231) <= not(layer3_outputs(633));
    layer4_outputs(3232) <= '0';
    layer4_outputs(3233) <= not((layer3_outputs(2423)) or (layer3_outputs(2184)));
    layer4_outputs(3234) <= (layer3_outputs(718)) or (layer3_outputs(4513));
    layer4_outputs(3235) <= not(layer3_outputs(919)) or (layer3_outputs(1239));
    layer4_outputs(3236) <= '0';
    layer4_outputs(3237) <= not(layer3_outputs(3833));
    layer4_outputs(3238) <= not(layer3_outputs(3333));
    layer4_outputs(3239) <= not(layer3_outputs(1168));
    layer4_outputs(3240) <= layer3_outputs(4646);
    layer4_outputs(3241) <= (layer3_outputs(3211)) and (layer3_outputs(2368));
    layer4_outputs(3242) <= layer3_outputs(2178);
    layer4_outputs(3243) <= '0';
    layer4_outputs(3244) <= not(layer3_outputs(1705));
    layer4_outputs(3245) <= (layer3_outputs(3069)) and not (layer3_outputs(4372));
    layer4_outputs(3246) <= layer3_outputs(3749);
    layer4_outputs(3247) <= layer3_outputs(3546);
    layer4_outputs(3248) <= (layer3_outputs(506)) or (layer3_outputs(1037));
    layer4_outputs(3249) <= (layer3_outputs(388)) and not (layer3_outputs(2318));
    layer4_outputs(3250) <= not(layer3_outputs(924));
    layer4_outputs(3251) <= (layer3_outputs(2410)) or (layer3_outputs(3885));
    layer4_outputs(3252) <= not(layer3_outputs(2903));
    layer4_outputs(3253) <= not(layer3_outputs(2506));
    layer4_outputs(3254) <= not(layer3_outputs(2548)) or (layer3_outputs(2384));
    layer4_outputs(3255) <= (layer3_outputs(4376)) or (layer3_outputs(4607));
    layer4_outputs(3256) <= layer3_outputs(2742);
    layer4_outputs(3257) <= not(layer3_outputs(2315)) or (layer3_outputs(725));
    layer4_outputs(3258) <= not(layer3_outputs(3996)) or (layer3_outputs(2510));
    layer4_outputs(3259) <= not((layer3_outputs(2204)) or (layer3_outputs(1547)));
    layer4_outputs(3260) <= not(layer3_outputs(2118)) or (layer3_outputs(546));
    layer4_outputs(3261) <= not(layer3_outputs(4863)) or (layer3_outputs(4716));
    layer4_outputs(3262) <= (layer3_outputs(87)) or (layer3_outputs(1242));
    layer4_outputs(3263) <= layer3_outputs(1343);
    layer4_outputs(3264) <= layer3_outputs(3068);
    layer4_outputs(3265) <= (layer3_outputs(4696)) or (layer3_outputs(215));
    layer4_outputs(3266) <= not(layer3_outputs(3034)) or (layer3_outputs(94));
    layer4_outputs(3267) <= (layer3_outputs(4286)) xor (layer3_outputs(3665));
    layer4_outputs(3268) <= layer3_outputs(3901);
    layer4_outputs(3269) <= (layer3_outputs(4212)) xor (layer3_outputs(2469));
    layer4_outputs(3270) <= not((layer3_outputs(3092)) and (layer3_outputs(4764)));
    layer4_outputs(3271) <= not((layer3_outputs(2827)) xor (layer3_outputs(3407)));
    layer4_outputs(3272) <= (layer3_outputs(3257)) or (layer3_outputs(3093));
    layer4_outputs(3273) <= (layer3_outputs(1655)) and not (layer3_outputs(4782));
    layer4_outputs(3274) <= not(layer3_outputs(593));
    layer4_outputs(3275) <= not(layer3_outputs(3225));
    layer4_outputs(3276) <= (layer3_outputs(2892)) xor (layer3_outputs(762));
    layer4_outputs(3277) <= (layer3_outputs(223)) and not (layer3_outputs(3324));
    layer4_outputs(3278) <= (layer3_outputs(4956)) xor (layer3_outputs(2191));
    layer4_outputs(3279) <= layer3_outputs(1162);
    layer4_outputs(3280) <= not(layer3_outputs(3339));
    layer4_outputs(3281) <= (layer3_outputs(2337)) xor (layer3_outputs(2704));
    layer4_outputs(3282) <= layer3_outputs(3235);
    layer4_outputs(3283) <= '1';
    layer4_outputs(3284) <= not((layer3_outputs(2994)) and (layer3_outputs(444)));
    layer4_outputs(3285) <= '0';
    layer4_outputs(3286) <= not((layer3_outputs(557)) or (layer3_outputs(2854)));
    layer4_outputs(3287) <= not(layer3_outputs(2978));
    layer4_outputs(3288) <= (layer3_outputs(1561)) or (layer3_outputs(3031));
    layer4_outputs(3289) <= layer3_outputs(2137);
    layer4_outputs(3290) <= not(layer3_outputs(84)) or (layer3_outputs(2265));
    layer4_outputs(3291) <= not(layer3_outputs(3552));
    layer4_outputs(3292) <= layer3_outputs(1528);
    layer4_outputs(3293) <= not((layer3_outputs(4054)) or (layer3_outputs(4658)));
    layer4_outputs(3294) <= not((layer3_outputs(3356)) or (layer3_outputs(1375)));
    layer4_outputs(3295) <= (layer3_outputs(2449)) and not (layer3_outputs(4128));
    layer4_outputs(3296) <= not(layer3_outputs(4315));
    layer4_outputs(3297) <= not(layer3_outputs(2499));
    layer4_outputs(3298) <= not(layer3_outputs(4010));
    layer4_outputs(3299) <= not(layer3_outputs(1202)) or (layer3_outputs(1155));
    layer4_outputs(3300) <= layer3_outputs(583);
    layer4_outputs(3301) <= not(layer3_outputs(4097));
    layer4_outputs(3302) <= (layer3_outputs(3508)) or (layer3_outputs(3373));
    layer4_outputs(3303) <= layer3_outputs(404);
    layer4_outputs(3304) <= not(layer3_outputs(4485));
    layer4_outputs(3305) <= (layer3_outputs(2493)) and not (layer3_outputs(4687));
    layer4_outputs(3306) <= '1';
    layer4_outputs(3307) <= (layer3_outputs(2133)) and not (layer3_outputs(1066));
    layer4_outputs(3308) <= not(layer3_outputs(667));
    layer4_outputs(3309) <= not(layer3_outputs(493));
    layer4_outputs(3310) <= not(layer3_outputs(3711));
    layer4_outputs(3311) <= not(layer3_outputs(3232)) or (layer3_outputs(4439));
    layer4_outputs(3312) <= not((layer3_outputs(2271)) or (layer3_outputs(4358)));
    layer4_outputs(3313) <= not(layer3_outputs(2326));
    layer4_outputs(3314) <= not(layer3_outputs(126));
    layer4_outputs(3315) <= not(layer3_outputs(1631)) or (layer3_outputs(3039));
    layer4_outputs(3316) <= layer3_outputs(4768);
    layer4_outputs(3317) <= not(layer3_outputs(3727));
    layer4_outputs(3318) <= not(layer3_outputs(2504));
    layer4_outputs(3319) <= not(layer3_outputs(593));
    layer4_outputs(3320) <= (layer3_outputs(474)) and not (layer3_outputs(1976));
    layer4_outputs(3321) <= (layer3_outputs(1251)) and (layer3_outputs(3581));
    layer4_outputs(3322) <= not((layer3_outputs(2607)) or (layer3_outputs(5034)));
    layer4_outputs(3323) <= not((layer3_outputs(1597)) xor (layer3_outputs(4344)));
    layer4_outputs(3324) <= not((layer3_outputs(618)) or (layer3_outputs(2935)));
    layer4_outputs(3325) <= layer3_outputs(3900);
    layer4_outputs(3326) <= not((layer3_outputs(689)) or (layer3_outputs(420)));
    layer4_outputs(3327) <= layer3_outputs(1355);
    layer4_outputs(3328) <= layer3_outputs(3774);
    layer4_outputs(3329) <= '1';
    layer4_outputs(3330) <= not((layer3_outputs(2802)) or (layer3_outputs(3797)));
    layer4_outputs(3331) <= '0';
    layer4_outputs(3332) <= layer3_outputs(1097);
    layer4_outputs(3333) <= not(layer3_outputs(1558));
    layer4_outputs(3334) <= (layer3_outputs(99)) or (layer3_outputs(164));
    layer4_outputs(3335) <= layer3_outputs(2054);
    layer4_outputs(3336) <= (layer3_outputs(605)) and not (layer3_outputs(3989));
    layer4_outputs(3337) <= layer3_outputs(1560);
    layer4_outputs(3338) <= (layer3_outputs(230)) and (layer3_outputs(1283));
    layer4_outputs(3339) <= (layer3_outputs(4572)) and not (layer3_outputs(391));
    layer4_outputs(3340) <= not(layer3_outputs(2187));
    layer4_outputs(3341) <= layer3_outputs(4264);
    layer4_outputs(3342) <= (layer3_outputs(1970)) or (layer3_outputs(4959));
    layer4_outputs(3343) <= not(layer3_outputs(1122)) or (layer3_outputs(1124));
    layer4_outputs(3344) <= not((layer3_outputs(2413)) and (layer3_outputs(3803)));
    layer4_outputs(3345) <= '0';
    layer4_outputs(3346) <= layer3_outputs(3493);
    layer4_outputs(3347) <= (layer3_outputs(4258)) xor (layer3_outputs(2864));
    layer4_outputs(3348) <= (layer3_outputs(4137)) or (layer3_outputs(3531));
    layer4_outputs(3349) <= not(layer3_outputs(4135)) or (layer3_outputs(1632));
    layer4_outputs(3350) <= not(layer3_outputs(233));
    layer4_outputs(3351) <= not((layer3_outputs(1167)) or (layer3_outputs(4206)));
    layer4_outputs(3352) <= not(layer3_outputs(4908));
    layer4_outputs(3353) <= not((layer3_outputs(579)) or (layer3_outputs(2628)));
    layer4_outputs(3354) <= not(layer3_outputs(4249));
    layer4_outputs(3355) <= layer3_outputs(2939);
    layer4_outputs(3356) <= not((layer3_outputs(2749)) and (layer3_outputs(2670)));
    layer4_outputs(3357) <= (layer3_outputs(1139)) or (layer3_outputs(3792));
    layer4_outputs(3358) <= layer3_outputs(4751);
    layer4_outputs(3359) <= layer3_outputs(1267);
    layer4_outputs(3360) <= not((layer3_outputs(3821)) and (layer3_outputs(4504)));
    layer4_outputs(3361) <= not((layer3_outputs(5030)) xor (layer3_outputs(3227)));
    layer4_outputs(3362) <= not(layer3_outputs(4336));
    layer4_outputs(3363) <= not(layer3_outputs(3834)) or (layer3_outputs(2200));
    layer4_outputs(3364) <= (layer3_outputs(82)) and not (layer3_outputs(1086));
    layer4_outputs(3365) <= not(layer3_outputs(370));
    layer4_outputs(3366) <= layer3_outputs(1359);
    layer4_outputs(3367) <= (layer3_outputs(407)) and not (layer3_outputs(308));
    layer4_outputs(3368) <= (layer3_outputs(1496)) or (layer3_outputs(3147));
    layer4_outputs(3369) <= layer3_outputs(1672);
    layer4_outputs(3370) <= '1';
    layer4_outputs(3371) <= not(layer3_outputs(1080)) or (layer3_outputs(676));
    layer4_outputs(3372) <= (layer3_outputs(4394)) and (layer3_outputs(2549));
    layer4_outputs(3373) <= not(layer3_outputs(3412));
    layer4_outputs(3374) <= '1';
    layer4_outputs(3375) <= not((layer3_outputs(3815)) xor (layer3_outputs(2121)));
    layer4_outputs(3376) <= '0';
    layer4_outputs(3377) <= (layer3_outputs(107)) or (layer3_outputs(3712));
    layer4_outputs(3378) <= (layer3_outputs(4503)) and not (layer3_outputs(4208));
    layer4_outputs(3379) <= layer3_outputs(921);
    layer4_outputs(3380) <= layer3_outputs(710);
    layer4_outputs(3381) <= not(layer3_outputs(278));
    layer4_outputs(3382) <= (layer3_outputs(2418)) and (layer3_outputs(4815));
    layer4_outputs(3383) <= (layer3_outputs(3454)) and not (layer3_outputs(4733));
    layer4_outputs(3384) <= not(layer3_outputs(385)) or (layer3_outputs(4350));
    layer4_outputs(3385) <= not((layer3_outputs(1782)) or (layer3_outputs(4381)));
    layer4_outputs(3386) <= not(layer3_outputs(3623));
    layer4_outputs(3387) <= not(layer3_outputs(1692));
    layer4_outputs(3388) <= (layer3_outputs(2743)) and (layer3_outputs(4156));
    layer4_outputs(3389) <= layer3_outputs(1409);
    layer4_outputs(3390) <= not(layer3_outputs(1168));
    layer4_outputs(3391) <= not(layer3_outputs(4408));
    layer4_outputs(3392) <= not(layer3_outputs(4008)) or (layer3_outputs(3558));
    layer4_outputs(3393) <= not((layer3_outputs(3055)) or (layer3_outputs(3633)));
    layer4_outputs(3394) <= not(layer3_outputs(4694)) or (layer3_outputs(2431));
    layer4_outputs(3395) <= not(layer3_outputs(4502));
    layer4_outputs(3396) <= not(layer3_outputs(269)) or (layer3_outputs(3271));
    layer4_outputs(3397) <= (layer3_outputs(5031)) and not (layer3_outputs(979));
    layer4_outputs(3398) <= (layer3_outputs(1924)) or (layer3_outputs(1653));
    layer4_outputs(3399) <= layer3_outputs(434);
    layer4_outputs(3400) <= not(layer3_outputs(1227));
    layer4_outputs(3401) <= not((layer3_outputs(4856)) and (layer3_outputs(5045)));
    layer4_outputs(3402) <= not(layer3_outputs(2067));
    layer4_outputs(3403) <= '0';
    layer4_outputs(3404) <= not((layer3_outputs(3740)) and (layer3_outputs(3170)));
    layer4_outputs(3405) <= layer3_outputs(4934);
    layer4_outputs(3406) <= not(layer3_outputs(774)) or (layer3_outputs(933));
    layer4_outputs(3407) <= not(layer3_outputs(3183)) or (layer3_outputs(4492));
    layer4_outputs(3408) <= (layer3_outputs(4019)) xor (layer3_outputs(4827));
    layer4_outputs(3409) <= not(layer3_outputs(322)) or (layer3_outputs(3848));
    layer4_outputs(3410) <= not((layer3_outputs(3782)) or (layer3_outputs(4179)));
    layer4_outputs(3411) <= not(layer3_outputs(3877));
    layer4_outputs(3412) <= (layer3_outputs(917)) and not (layer3_outputs(4651));
    layer4_outputs(3413) <= (layer3_outputs(480)) and (layer3_outputs(1007));
    layer4_outputs(3414) <= layer3_outputs(2794);
    layer4_outputs(3415) <= layer3_outputs(2188);
    layer4_outputs(3416) <= '1';
    layer4_outputs(3417) <= (layer3_outputs(1948)) and not (layer3_outputs(3842));
    layer4_outputs(3418) <= (layer3_outputs(3228)) and (layer3_outputs(2812));
    layer4_outputs(3419) <= not(layer3_outputs(2110));
    layer4_outputs(3420) <= (layer3_outputs(560)) and (layer3_outputs(3900));
    layer4_outputs(3421) <= layer3_outputs(2884);
    layer4_outputs(3422) <= (layer3_outputs(3730)) and not (layer3_outputs(1385));
    layer4_outputs(3423) <= (layer3_outputs(1128)) and (layer3_outputs(3446));
    layer4_outputs(3424) <= layer3_outputs(2119);
    layer4_outputs(3425) <= '0';
    layer4_outputs(3426) <= (layer3_outputs(2774)) or (layer3_outputs(4130));
    layer4_outputs(3427) <= not(layer3_outputs(1617));
    layer4_outputs(3428) <= not(layer3_outputs(3133));
    layer4_outputs(3429) <= not(layer3_outputs(90));
    layer4_outputs(3430) <= (layer3_outputs(4421)) and not (layer3_outputs(654));
    layer4_outputs(3431) <= layer3_outputs(3873);
    layer4_outputs(3432) <= (layer3_outputs(1238)) and not (layer3_outputs(2888));
    layer4_outputs(3433) <= (layer3_outputs(3088)) or (layer3_outputs(1623));
    layer4_outputs(3434) <= not(layer3_outputs(844));
    layer4_outputs(3435) <= not(layer3_outputs(3484));
    layer4_outputs(3436) <= (layer3_outputs(2123)) and not (layer3_outputs(3232));
    layer4_outputs(3437) <= (layer3_outputs(4152)) and not (layer3_outputs(3806));
    layer4_outputs(3438) <= (layer3_outputs(3834)) and not (layer3_outputs(1419));
    layer4_outputs(3439) <= (layer3_outputs(4648)) and not (layer3_outputs(1529));
    layer4_outputs(3440) <= layer3_outputs(3747);
    layer4_outputs(3441) <= '1';
    layer4_outputs(3442) <= (layer3_outputs(4048)) and not (layer3_outputs(4153));
    layer4_outputs(3443) <= not(layer3_outputs(5015));
    layer4_outputs(3444) <= not(layer3_outputs(4059));
    layer4_outputs(3445) <= (layer3_outputs(4984)) or (layer3_outputs(2882));
    layer4_outputs(3446) <= not((layer3_outputs(735)) or (layer3_outputs(2229)));
    layer4_outputs(3447) <= not((layer3_outputs(3563)) or (layer3_outputs(3620)));
    layer4_outputs(3448) <= '0';
    layer4_outputs(3449) <= layer3_outputs(3668);
    layer4_outputs(3450) <= not(layer3_outputs(3056));
    layer4_outputs(3451) <= not(layer3_outputs(5001));
    layer4_outputs(3452) <= (layer3_outputs(4783)) and (layer3_outputs(3629));
    layer4_outputs(3453) <= (layer3_outputs(1982)) or (layer3_outputs(2832));
    layer4_outputs(3454) <= not(layer3_outputs(2763));
    layer4_outputs(3455) <= not(layer3_outputs(4254)) or (layer3_outputs(2528));
    layer4_outputs(3456) <= not(layer3_outputs(3223));
    layer4_outputs(3457) <= not(layer3_outputs(199)) or (layer3_outputs(3696));
    layer4_outputs(3458) <= layer3_outputs(3238);
    layer4_outputs(3459) <= (layer3_outputs(1029)) or (layer3_outputs(2201));
    layer4_outputs(3460) <= layer3_outputs(4707);
    layer4_outputs(3461) <= '0';
    layer4_outputs(3462) <= not(layer3_outputs(1989));
    layer4_outputs(3463) <= not(layer3_outputs(1058));
    layer4_outputs(3464) <= layer3_outputs(3487);
    layer4_outputs(3465) <= not(layer3_outputs(2223));
    layer4_outputs(3466) <= layer3_outputs(4451);
    layer4_outputs(3467) <= not((layer3_outputs(3235)) xor (layer3_outputs(1197)));
    layer4_outputs(3468) <= layer3_outputs(1048);
    layer4_outputs(3469) <= layer3_outputs(4145);
    layer4_outputs(3470) <= not((layer3_outputs(1436)) or (layer3_outputs(1212)));
    layer4_outputs(3471) <= (layer3_outputs(1535)) and not (layer3_outputs(1821));
    layer4_outputs(3472) <= not((layer3_outputs(2471)) xor (layer3_outputs(2593)));
    layer4_outputs(3473) <= not(layer3_outputs(4619));
    layer4_outputs(3474) <= layer3_outputs(1148);
    layer4_outputs(3475) <= '0';
    layer4_outputs(3476) <= (layer3_outputs(4100)) or (layer3_outputs(1614));
    layer4_outputs(3477) <= layer3_outputs(2801);
    layer4_outputs(3478) <= not(layer3_outputs(450));
    layer4_outputs(3479) <= '1';
    layer4_outputs(3480) <= (layer3_outputs(2334)) and not (layer3_outputs(2577));
    layer4_outputs(3481) <= not(layer3_outputs(1346));
    layer4_outputs(3482) <= (layer3_outputs(3631)) or (layer3_outputs(2621));
    layer4_outputs(3483) <= (layer3_outputs(2149)) and not (layer3_outputs(628));
    layer4_outputs(3484) <= not(layer3_outputs(3448));
    layer4_outputs(3485) <= not(layer3_outputs(2453)) or (layer3_outputs(743));
    layer4_outputs(3486) <= layer3_outputs(1291);
    layer4_outputs(3487) <= layer3_outputs(3361);
    layer4_outputs(3488) <= '1';
    layer4_outputs(3489) <= not((layer3_outputs(4035)) and (layer3_outputs(2776)));
    layer4_outputs(3490) <= not(layer3_outputs(1931));
    layer4_outputs(3491) <= (layer3_outputs(670)) or (layer3_outputs(946));
    layer4_outputs(3492) <= not((layer3_outputs(3640)) and (layer3_outputs(4480)));
    layer4_outputs(3493) <= not(layer3_outputs(3424));
    layer4_outputs(3494) <= not(layer3_outputs(2694)) or (layer3_outputs(5035));
    layer4_outputs(3495) <= not(layer3_outputs(2446)) or (layer3_outputs(1498));
    layer4_outputs(3496) <= not(layer3_outputs(5053));
    layer4_outputs(3497) <= not(layer3_outputs(2364));
    layer4_outputs(3498) <= not(layer3_outputs(2646));
    layer4_outputs(3499) <= layer3_outputs(956);
    layer4_outputs(3500) <= not((layer3_outputs(165)) and (layer3_outputs(2487)));
    layer4_outputs(3501) <= (layer3_outputs(4780)) and not (layer3_outputs(2087));
    layer4_outputs(3502) <= not((layer3_outputs(485)) and (layer3_outputs(100)));
    layer4_outputs(3503) <= (layer3_outputs(1179)) and not (layer3_outputs(4957));
    layer4_outputs(3504) <= not(layer3_outputs(405));
    layer4_outputs(3505) <= (layer3_outputs(2964)) and (layer3_outputs(1737));
    layer4_outputs(3506) <= not(layer3_outputs(4067));
    layer4_outputs(3507) <= '1';
    layer4_outputs(3508) <= not(layer3_outputs(505));
    layer4_outputs(3509) <= layer3_outputs(1194);
    layer4_outputs(3510) <= not((layer3_outputs(3129)) or (layer3_outputs(3040)));
    layer4_outputs(3511) <= not(layer3_outputs(2673));
    layer4_outputs(3512) <= not(layer3_outputs(2201)) or (layer3_outputs(4234));
    layer4_outputs(3513) <= not(layer3_outputs(1560));
    layer4_outputs(3514) <= (layer3_outputs(4481)) and not (layer3_outputs(3197));
    layer4_outputs(3515) <= not(layer3_outputs(4402));
    layer4_outputs(3516) <= not((layer3_outputs(2759)) and (layer3_outputs(1327)));
    layer4_outputs(3517) <= '0';
    layer4_outputs(3518) <= not(layer3_outputs(3365)) or (layer3_outputs(216));
    layer4_outputs(3519) <= not(layer3_outputs(990));
    layer4_outputs(3520) <= layer3_outputs(1979);
    layer4_outputs(3521) <= not((layer3_outputs(9)) and (layer3_outputs(3615)));
    layer4_outputs(3522) <= '0';
    layer4_outputs(3523) <= not(layer3_outputs(3318));
    layer4_outputs(3524) <= layer3_outputs(1495);
    layer4_outputs(3525) <= (layer3_outputs(1654)) and not (layer3_outputs(530));
    layer4_outputs(3526) <= (layer3_outputs(2417)) or (layer3_outputs(2104));
    layer4_outputs(3527) <= not(layer3_outputs(1478)) or (layer3_outputs(4373));
    layer4_outputs(3528) <= (layer3_outputs(1330)) xor (layer3_outputs(4462));
    layer4_outputs(3529) <= not((layer3_outputs(3317)) or (layer3_outputs(761)));
    layer4_outputs(3530) <= not(layer3_outputs(4159));
    layer4_outputs(3531) <= (layer3_outputs(3341)) and (layer3_outputs(915));
    layer4_outputs(3532) <= not(layer3_outputs(1452));
    layer4_outputs(3533) <= (layer3_outputs(1704)) xor (layer3_outputs(3876));
    layer4_outputs(3534) <= not(layer3_outputs(4036));
    layer4_outputs(3535) <= not(layer3_outputs(4212)) or (layer3_outputs(604));
    layer4_outputs(3536) <= not(layer3_outputs(1878));
    layer4_outputs(3537) <= not((layer3_outputs(983)) or (layer3_outputs(4884)));
    layer4_outputs(3538) <= not(layer3_outputs(3061));
    layer4_outputs(3539) <= not(layer3_outputs(2623));
    layer4_outputs(3540) <= not(layer3_outputs(4513));
    layer4_outputs(3541) <= layer3_outputs(2942);
    layer4_outputs(3542) <= layer3_outputs(130);
    layer4_outputs(3543) <= layer3_outputs(5033);
    layer4_outputs(3544) <= layer3_outputs(4598);
    layer4_outputs(3545) <= (layer3_outputs(4331)) and (layer3_outputs(4538));
    layer4_outputs(3546) <= not(layer3_outputs(3566));
    layer4_outputs(3547) <= layer3_outputs(3191);
    layer4_outputs(3548) <= not(layer3_outputs(4329));
    layer4_outputs(3549) <= (layer3_outputs(2917)) and (layer3_outputs(845));
    layer4_outputs(3550) <= layer3_outputs(4810);
    layer4_outputs(3551) <= not(layer3_outputs(3445));
    layer4_outputs(3552) <= (layer3_outputs(2821)) and not (layer3_outputs(2999));
    layer4_outputs(3553) <= not(layer3_outputs(4438));
    layer4_outputs(3554) <= layer3_outputs(165);
    layer4_outputs(3555) <= layer3_outputs(442);
    layer4_outputs(3556) <= not(layer3_outputs(4448)) or (layer3_outputs(2321));
    layer4_outputs(3557) <= not(layer3_outputs(4446)) or (layer3_outputs(1356));
    layer4_outputs(3558) <= (layer3_outputs(2654)) and (layer3_outputs(3343));
    layer4_outputs(3559) <= layer3_outputs(4274);
    layer4_outputs(3560) <= '0';
    layer4_outputs(3561) <= layer3_outputs(1146);
    layer4_outputs(3562) <= not(layer3_outputs(2004));
    layer4_outputs(3563) <= not((layer3_outputs(288)) and (layer3_outputs(3606)));
    layer4_outputs(3564) <= not(layer3_outputs(2268));
    layer4_outputs(3565) <= layer3_outputs(4567);
    layer4_outputs(3566) <= '1';
    layer4_outputs(3567) <= layer3_outputs(3590);
    layer4_outputs(3568) <= '1';
    layer4_outputs(3569) <= layer3_outputs(4257);
    layer4_outputs(3570) <= (layer3_outputs(629)) and (layer3_outputs(5087));
    layer4_outputs(3571) <= layer3_outputs(4121);
    layer4_outputs(3572) <= not(layer3_outputs(7));
    layer4_outputs(3573) <= not(layer3_outputs(3119));
    layer4_outputs(3574) <= layer3_outputs(739);
    layer4_outputs(3575) <= (layer3_outputs(627)) or (layer3_outputs(197));
    layer4_outputs(3576) <= not(layer3_outputs(4044));
    layer4_outputs(3577) <= not((layer3_outputs(4575)) and (layer3_outputs(4393)));
    layer4_outputs(3578) <= not((layer3_outputs(4147)) or (layer3_outputs(3181)));
    layer4_outputs(3579) <= layer3_outputs(1451);
    layer4_outputs(3580) <= not(layer3_outputs(3013));
    layer4_outputs(3581) <= layer3_outputs(912);
    layer4_outputs(3582) <= '1';
    layer4_outputs(3583) <= layer3_outputs(2932);
    layer4_outputs(3584) <= not(layer3_outputs(3569)) or (layer3_outputs(4227));
    layer4_outputs(3585) <= (layer3_outputs(4294)) and not (layer3_outputs(3322));
    layer4_outputs(3586) <= '0';
    layer4_outputs(3587) <= not(layer3_outputs(2347)) or (layer3_outputs(360));
    layer4_outputs(3588) <= (layer3_outputs(3671)) and (layer3_outputs(3912));
    layer4_outputs(3589) <= (layer3_outputs(4482)) and (layer3_outputs(121));
    layer4_outputs(3590) <= not(layer3_outputs(1425));
    layer4_outputs(3591) <= not(layer3_outputs(3886));
    layer4_outputs(3592) <= not((layer3_outputs(429)) and (layer3_outputs(1913)));
    layer4_outputs(3593) <= layer3_outputs(4277);
    layer4_outputs(3594) <= not(layer3_outputs(2106));
    layer4_outputs(3595) <= layer3_outputs(3504);
    layer4_outputs(3596) <= layer3_outputs(1743);
    layer4_outputs(3597) <= '0';
    layer4_outputs(3598) <= layer3_outputs(4392);
    layer4_outputs(3599) <= not(layer3_outputs(2052));
    layer4_outputs(3600) <= (layer3_outputs(3932)) and not (layer3_outputs(4167));
    layer4_outputs(3601) <= not(layer3_outputs(2823));
    layer4_outputs(3602) <= not((layer3_outputs(3755)) xor (layer3_outputs(2923)));
    layer4_outputs(3603) <= '1';
    layer4_outputs(3604) <= not(layer3_outputs(2679));
    layer4_outputs(3605) <= not(layer3_outputs(1388)) or (layer3_outputs(2821));
    layer4_outputs(3606) <= (layer3_outputs(1979)) or (layer3_outputs(432));
    layer4_outputs(3607) <= layer3_outputs(4742);
    layer4_outputs(3608) <= layer3_outputs(2461);
    layer4_outputs(3609) <= not(layer3_outputs(4424));
    layer4_outputs(3610) <= layer3_outputs(2718);
    layer4_outputs(3611) <= not(layer3_outputs(4387)) or (layer3_outputs(232));
    layer4_outputs(3612) <= (layer3_outputs(2215)) xor (layer3_outputs(2238));
    layer4_outputs(3613) <= '0';
    layer4_outputs(3614) <= not(layer3_outputs(1081));
    layer4_outputs(3615) <= not((layer3_outputs(42)) or (layer3_outputs(4075)));
    layer4_outputs(3616) <= not(layer3_outputs(2313)) or (layer3_outputs(5070));
    layer4_outputs(3617) <= not(layer3_outputs(1290)) or (layer3_outputs(1211));
    layer4_outputs(3618) <= not(layer3_outputs(4151)) or (layer3_outputs(290));
    layer4_outputs(3619) <= not(layer3_outputs(4477));
    layer4_outputs(3620) <= layer3_outputs(931);
    layer4_outputs(3621) <= not(layer3_outputs(3284));
    layer4_outputs(3622) <= '1';
    layer4_outputs(3623) <= (layer3_outputs(4612)) and not (layer3_outputs(3441));
    layer4_outputs(3624) <= '0';
    layer4_outputs(3625) <= '0';
    layer4_outputs(3626) <= (layer3_outputs(1967)) and (layer3_outputs(652));
    layer4_outputs(3627) <= '0';
    layer4_outputs(3628) <= not(layer3_outputs(4334)) or (layer3_outputs(989));
    layer4_outputs(3629) <= (layer3_outputs(920)) and (layer3_outputs(3180));
    layer4_outputs(3630) <= (layer3_outputs(1258)) and (layer3_outputs(4995));
    layer4_outputs(3631) <= not(layer3_outputs(3157));
    layer4_outputs(3632) <= '0';
    layer4_outputs(3633) <= not(layer3_outputs(2003));
    layer4_outputs(3634) <= not(layer3_outputs(1843)) or (layer3_outputs(307));
    layer4_outputs(3635) <= (layer3_outputs(639)) or (layer3_outputs(386));
    layer4_outputs(3636) <= layer3_outputs(572);
    layer4_outputs(3637) <= (layer3_outputs(551)) and not (layer3_outputs(3456));
    layer4_outputs(3638) <= not(layer3_outputs(1261)) or (layer3_outputs(1130));
    layer4_outputs(3639) <= (layer3_outputs(2412)) and not (layer3_outputs(1222));
    layer4_outputs(3640) <= layer3_outputs(957);
    layer4_outputs(3641) <= not((layer3_outputs(4939)) or (layer3_outputs(286)));
    layer4_outputs(3642) <= not((layer3_outputs(1682)) or (layer3_outputs(4735)));
    layer4_outputs(3643) <= not(layer3_outputs(996));
    layer4_outputs(3644) <= layer3_outputs(4510);
    layer4_outputs(3645) <= not(layer3_outputs(4499));
    layer4_outputs(3646) <= not(layer3_outputs(2521));
    layer4_outputs(3647) <= not((layer3_outputs(1856)) and (layer3_outputs(1984)));
    layer4_outputs(3648) <= layer3_outputs(3212);
    layer4_outputs(3649) <= (layer3_outputs(4541)) and not (layer3_outputs(2179));
    layer4_outputs(3650) <= not(layer3_outputs(1823));
    layer4_outputs(3651) <= (layer3_outputs(4291)) and not (layer3_outputs(1955));
    layer4_outputs(3652) <= (layer3_outputs(4976)) xor (layer3_outputs(288));
    layer4_outputs(3653) <= not(layer3_outputs(949)) or (layer3_outputs(242));
    layer4_outputs(3654) <= (layer3_outputs(4561)) or (layer3_outputs(575));
    layer4_outputs(3655) <= layer3_outputs(948);
    layer4_outputs(3656) <= not(layer3_outputs(1344)) or (layer3_outputs(637));
    layer4_outputs(3657) <= (layer3_outputs(2726)) or (layer3_outputs(3481));
    layer4_outputs(3658) <= not((layer3_outputs(3200)) and (layer3_outputs(1971)));
    layer4_outputs(3659) <= not((layer3_outputs(1537)) and (layer3_outputs(1495)));
    layer4_outputs(3660) <= '0';
    layer4_outputs(3661) <= layer3_outputs(4836);
    layer4_outputs(3662) <= not(layer3_outputs(4326)) or (layer3_outputs(2166));
    layer4_outputs(3663) <= layer3_outputs(4764);
    layer4_outputs(3664) <= not(layer3_outputs(1309));
    layer4_outputs(3665) <= not(layer3_outputs(3816)) or (layer3_outputs(541));
    layer4_outputs(3666) <= not(layer3_outputs(3612));
    layer4_outputs(3667) <= (layer3_outputs(5107)) and not (layer3_outputs(2092));
    layer4_outputs(3668) <= layer3_outputs(1204);
    layer4_outputs(3669) <= (layer3_outputs(4265)) or (layer3_outputs(1694));
    layer4_outputs(3670) <= not((layer3_outputs(4613)) or (layer3_outputs(2922)));
    layer4_outputs(3671) <= not((layer3_outputs(721)) and (layer3_outputs(1820)));
    layer4_outputs(3672) <= '1';
    layer4_outputs(3673) <= (layer3_outputs(4598)) and not (layer3_outputs(98));
    layer4_outputs(3674) <= layer3_outputs(2778);
    layer4_outputs(3675) <= not((layer3_outputs(4534)) or (layer3_outputs(1863)));
    layer4_outputs(3676) <= '0';
    layer4_outputs(3677) <= layer3_outputs(1307);
    layer4_outputs(3678) <= (layer3_outputs(383)) and (layer3_outputs(2538));
    layer4_outputs(3679) <= (layer3_outputs(381)) and not (layer3_outputs(2007));
    layer4_outputs(3680) <= not(layer3_outputs(594));
    layer4_outputs(3681) <= not(layer3_outputs(4789)) or (layer3_outputs(3216));
    layer4_outputs(3682) <= not(layer3_outputs(2926));
    layer4_outputs(3683) <= layer3_outputs(236);
    layer4_outputs(3684) <= layer3_outputs(346);
    layer4_outputs(3685) <= not(layer3_outputs(4361)) or (layer3_outputs(1282));
    layer4_outputs(3686) <= (layer3_outputs(3856)) or (layer3_outputs(3315));
    layer4_outputs(3687) <= not(layer3_outputs(1033));
    layer4_outputs(3688) <= '0';
    layer4_outputs(3689) <= layer3_outputs(943);
    layer4_outputs(3690) <= (layer3_outputs(2320)) and (layer3_outputs(2303));
    layer4_outputs(3691) <= not(layer3_outputs(2089)) or (layer3_outputs(4301));
    layer4_outputs(3692) <= '0';
    layer4_outputs(3693) <= layer3_outputs(4207);
    layer4_outputs(3694) <= (layer3_outputs(98)) and not (layer3_outputs(769));
    layer4_outputs(3695) <= (layer3_outputs(1570)) and not (layer3_outputs(2427));
    layer4_outputs(3696) <= not(layer3_outputs(3516));
    layer4_outputs(3697) <= not((layer3_outputs(3561)) xor (layer3_outputs(2752)));
    layer4_outputs(3698) <= not(layer3_outputs(2157));
    layer4_outputs(3699) <= layer3_outputs(1311);
    layer4_outputs(3700) <= (layer3_outputs(4333)) and (layer3_outputs(4107));
    layer4_outputs(3701) <= not(layer3_outputs(3947));
    layer4_outputs(3702) <= (layer3_outputs(1166)) xor (layer3_outputs(2899));
    layer4_outputs(3703) <= (layer3_outputs(2220)) and (layer3_outputs(161));
    layer4_outputs(3704) <= layer3_outputs(712);
    layer4_outputs(3705) <= (layer3_outputs(864)) and not (layer3_outputs(4986));
    layer4_outputs(3706) <= layer3_outputs(2458);
    layer4_outputs(3707) <= not((layer3_outputs(4443)) or (layer3_outputs(229)));
    layer4_outputs(3708) <= not((layer3_outputs(3208)) or (layer3_outputs(881)));
    layer4_outputs(3709) <= not(layer3_outputs(4452));
    layer4_outputs(3710) <= not((layer3_outputs(4982)) or (layer3_outputs(2573)));
    layer4_outputs(3711) <= (layer3_outputs(1266)) and (layer3_outputs(2535));
    layer4_outputs(3712) <= (layer3_outputs(4622)) and not (layer3_outputs(2082));
    layer4_outputs(3713) <= (layer3_outputs(2065)) and not (layer3_outputs(2949));
    layer4_outputs(3714) <= not(layer3_outputs(2789));
    layer4_outputs(3715) <= not(layer3_outputs(2859));
    layer4_outputs(3716) <= layer3_outputs(1755);
    layer4_outputs(3717) <= not(layer3_outputs(4719));
    layer4_outputs(3718) <= (layer3_outputs(246)) and (layer3_outputs(2734));
    layer4_outputs(3719) <= layer3_outputs(3843);
    layer4_outputs(3720) <= '1';
    layer4_outputs(3721) <= not(layer3_outputs(2018)) or (layer3_outputs(4150));
    layer4_outputs(3722) <= not(layer3_outputs(1660)) or (layer3_outputs(1030));
    layer4_outputs(3723) <= not(layer3_outputs(581));
    layer4_outputs(3724) <= layer3_outputs(1744);
    layer4_outputs(3725) <= not(layer3_outputs(3574));
    layer4_outputs(3726) <= not(layer3_outputs(631));
    layer4_outputs(3727) <= '1';
    layer4_outputs(3728) <= layer3_outputs(936);
    layer4_outputs(3729) <= (layer3_outputs(2751)) and (layer3_outputs(4216));
    layer4_outputs(3730) <= layer3_outputs(4025);
    layer4_outputs(3731) <= '0';
    layer4_outputs(3732) <= (layer3_outputs(430)) and (layer3_outputs(4968));
    layer4_outputs(3733) <= not(layer3_outputs(4118));
    layer4_outputs(3734) <= '1';
    layer4_outputs(3735) <= '1';
    layer4_outputs(3736) <= '1';
    layer4_outputs(3737) <= (layer3_outputs(3205)) or (layer3_outputs(4302));
    layer4_outputs(3738) <= layer3_outputs(1430);
    layer4_outputs(3739) <= (layer3_outputs(4998)) or (layer3_outputs(561));
    layer4_outputs(3740) <= not(layer3_outputs(1544));
    layer4_outputs(3741) <= (layer3_outputs(836)) xor (layer3_outputs(1449));
    layer4_outputs(3742) <= (layer3_outputs(4942)) and (layer3_outputs(2739));
    layer4_outputs(3743) <= not((layer3_outputs(2621)) xor (layer3_outputs(4532)));
    layer4_outputs(3744) <= not((layer3_outputs(2589)) and (layer3_outputs(1856)));
    layer4_outputs(3745) <= (layer3_outputs(2276)) and (layer3_outputs(2011));
    layer4_outputs(3746) <= not(layer3_outputs(3784));
    layer4_outputs(3747) <= layer3_outputs(5056);
    layer4_outputs(3748) <= not(layer3_outputs(2090)) or (layer3_outputs(954));
    layer4_outputs(3749) <= layer3_outputs(3783);
    layer4_outputs(3750) <= layer3_outputs(4116);
    layer4_outputs(3751) <= not((layer3_outputs(2895)) or (layer3_outputs(2088)));
    layer4_outputs(3752) <= not(layer3_outputs(4349)) or (layer3_outputs(1590));
    layer4_outputs(3753) <= not((layer3_outputs(349)) or (layer3_outputs(2270)));
    layer4_outputs(3754) <= not(layer3_outputs(4404));
    layer4_outputs(3755) <= layer3_outputs(2482);
    layer4_outputs(3756) <= not(layer3_outputs(2468)) or (layer3_outputs(4652));
    layer4_outputs(3757) <= (layer3_outputs(4847)) xor (layer3_outputs(1828));
    layer4_outputs(3758) <= layer3_outputs(1501);
    layer4_outputs(3759) <= layer3_outputs(4618);
    layer4_outputs(3760) <= (layer3_outputs(828)) xor (layer3_outputs(47));
    layer4_outputs(3761) <= (layer3_outputs(2480)) and not (layer3_outputs(1358));
    layer4_outputs(3762) <= (layer3_outputs(3207)) xor (layer3_outputs(4196));
    layer4_outputs(3763) <= layer3_outputs(563);
    layer4_outputs(3764) <= (layer3_outputs(1830)) and not (layer3_outputs(3311));
    layer4_outputs(3765) <= (layer3_outputs(1544)) and (layer3_outputs(2897));
    layer4_outputs(3766) <= not((layer3_outputs(1634)) or (layer3_outputs(2312)));
    layer4_outputs(3767) <= not((layer3_outputs(1569)) and (layer3_outputs(400)));
    layer4_outputs(3768) <= not(layer3_outputs(4280)) or (layer3_outputs(4717));
    layer4_outputs(3769) <= layer3_outputs(5);
    layer4_outputs(3770) <= layer3_outputs(3043);
    layer4_outputs(3771) <= layer3_outputs(5055);
    layer4_outputs(3772) <= not(layer3_outputs(1812));
    layer4_outputs(3773) <= not(layer3_outputs(1284));
    layer4_outputs(3774) <= layer3_outputs(4336);
    layer4_outputs(3775) <= (layer3_outputs(2247)) and (layer3_outputs(1588));
    layer4_outputs(3776) <= (layer3_outputs(1037)) and not (layer3_outputs(495));
    layer4_outputs(3777) <= (layer3_outputs(2553)) or (layer3_outputs(3964));
    layer4_outputs(3778) <= not((layer3_outputs(439)) xor (layer3_outputs(3074)));
    layer4_outputs(3779) <= not((layer3_outputs(2888)) and (layer3_outputs(4590)));
    layer4_outputs(3780) <= layer3_outputs(657);
    layer4_outputs(3781) <= not(layer3_outputs(1306));
    layer4_outputs(3782) <= not(layer3_outputs(4763));
    layer4_outputs(3783) <= layer3_outputs(4906);
    layer4_outputs(3784) <= layer3_outputs(2668);
    layer4_outputs(3785) <= layer3_outputs(4391);
    layer4_outputs(3786) <= '0';
    layer4_outputs(3787) <= layer3_outputs(3618);
    layer4_outputs(3788) <= layer3_outputs(3962);
    layer4_outputs(3789) <= '1';
    layer4_outputs(3790) <= '0';
    layer4_outputs(3791) <= (layer3_outputs(1652)) and not (layer3_outputs(1491));
    layer4_outputs(3792) <= (layer3_outputs(4468)) and not (layer3_outputs(3554));
    layer4_outputs(3793) <= layer3_outputs(38);
    layer4_outputs(3794) <= (layer3_outputs(225)) and not (layer3_outputs(3069));
    layer4_outputs(3795) <= not((layer3_outputs(3059)) xor (layer3_outputs(1315)));
    layer4_outputs(3796) <= layer3_outputs(3375);
    layer4_outputs(3797) <= not(layer3_outputs(1869));
    layer4_outputs(3798) <= not(layer3_outputs(3586));
    layer4_outputs(3799) <= not((layer3_outputs(3945)) and (layer3_outputs(2053)));
    layer4_outputs(3800) <= not((layer3_outputs(1274)) and (layer3_outputs(1580)));
    layer4_outputs(3801) <= not(layer3_outputs(2262)) or (layer3_outputs(3097));
    layer4_outputs(3802) <= (layer3_outputs(4018)) and (layer3_outputs(325));
    layer4_outputs(3803) <= layer3_outputs(3895);
    layer4_outputs(3804) <= not((layer3_outputs(1151)) xor (layer3_outputs(2024)));
    layer4_outputs(3805) <= not((layer3_outputs(3242)) or (layer3_outputs(2533)));
    layer4_outputs(3806) <= layer3_outputs(4202);
    layer4_outputs(3807) <= layer3_outputs(3208);
    layer4_outputs(3808) <= (layer3_outputs(3295)) and not (layer3_outputs(1761));
    layer4_outputs(3809) <= not(layer3_outputs(5077));
    layer4_outputs(3810) <= not((layer3_outputs(658)) xor (layer3_outputs(3010)));
    layer4_outputs(3811) <= '1';
    layer4_outputs(3812) <= (layer3_outputs(2159)) and not (layer3_outputs(2392));
    layer4_outputs(3813) <= not(layer3_outputs(1575)) or (layer3_outputs(1086));
    layer4_outputs(3814) <= (layer3_outputs(4014)) xor (layer3_outputs(4407));
    layer4_outputs(3815) <= (layer3_outputs(3028)) and not (layer3_outputs(4779));
    layer4_outputs(3816) <= (layer3_outputs(3329)) and not (layer3_outputs(2781));
    layer4_outputs(3817) <= not(layer3_outputs(435));
    layer4_outputs(3818) <= (layer3_outputs(1868)) and (layer3_outputs(964));
    layer4_outputs(3819) <= layer3_outputs(4254);
    layer4_outputs(3820) <= layer3_outputs(162);
    layer4_outputs(3821) <= not((layer3_outputs(4562)) or (layer3_outputs(3892)));
    layer4_outputs(3822) <= layer3_outputs(2313);
    layer4_outputs(3823) <= not((layer3_outputs(1349)) or (layer3_outputs(443)));
    layer4_outputs(3824) <= layer3_outputs(751);
    layer4_outputs(3825) <= not((layer3_outputs(4638)) or (layer3_outputs(2319)));
    layer4_outputs(3826) <= (layer3_outputs(1346)) and not (layer3_outputs(4684));
    layer4_outputs(3827) <= not((layer3_outputs(1477)) xor (layer3_outputs(2902)));
    layer4_outputs(3828) <= layer3_outputs(3367);
    layer4_outputs(3829) <= '0';
    layer4_outputs(3830) <= layer3_outputs(1241);
    layer4_outputs(3831) <= layer3_outputs(57);
    layer4_outputs(3832) <= not((layer3_outputs(1791)) and (layer3_outputs(2109)));
    layer4_outputs(3833) <= layer3_outputs(1709);
    layer4_outputs(3834) <= (layer3_outputs(4576)) and not (layer3_outputs(2495));
    layer4_outputs(3835) <= (layer3_outputs(2350)) and (layer3_outputs(2451));
    layer4_outputs(3836) <= not(layer3_outputs(4927)) or (layer3_outputs(1527));
    layer4_outputs(3837) <= (layer3_outputs(524)) and (layer3_outputs(1004));
    layer4_outputs(3838) <= not(layer3_outputs(1599));
    layer4_outputs(3839) <= not(layer3_outputs(3844));
    layer4_outputs(3840) <= layer3_outputs(4224);
    layer4_outputs(3841) <= (layer3_outputs(1947)) and not (layer3_outputs(1342));
    layer4_outputs(3842) <= '0';
    layer4_outputs(3843) <= (layer3_outputs(1186)) and not (layer3_outputs(2663));
    layer4_outputs(3844) <= '0';
    layer4_outputs(3845) <= (layer3_outputs(2746)) and (layer3_outputs(3096));
    layer4_outputs(3846) <= layer3_outputs(2453);
    layer4_outputs(3847) <= not(layer3_outputs(3892));
    layer4_outputs(3848) <= layer3_outputs(441);
    layer4_outputs(3849) <= not((layer3_outputs(771)) and (layer3_outputs(4295)));
    layer4_outputs(3850) <= not(layer3_outputs(2593));
    layer4_outputs(3851) <= (layer3_outputs(4615)) and not (layer3_outputs(325));
    layer4_outputs(3852) <= not(layer3_outputs(1109));
    layer4_outputs(3853) <= layer3_outputs(128);
    layer4_outputs(3854) <= not(layer3_outputs(936)) or (layer3_outputs(1241));
    layer4_outputs(3855) <= (layer3_outputs(132)) and not (layer3_outputs(1023));
    layer4_outputs(3856) <= not((layer3_outputs(3961)) xor (layer3_outputs(836)));
    layer4_outputs(3857) <= not(layer3_outputs(4849));
    layer4_outputs(3858) <= layer3_outputs(892);
    layer4_outputs(3859) <= layer3_outputs(2750);
    layer4_outputs(3860) <= '1';
    layer4_outputs(3861) <= (layer3_outputs(4604)) and not (layer3_outputs(1669));
    layer4_outputs(3862) <= layer3_outputs(155);
    layer4_outputs(3863) <= not(layer3_outputs(1398)) or (layer3_outputs(4573));
    layer4_outputs(3864) <= not(layer3_outputs(1345)) or (layer3_outputs(2858));
    layer4_outputs(3865) <= '1';
    layer4_outputs(3866) <= (layer3_outputs(3400)) and (layer3_outputs(83));
    layer4_outputs(3867) <= layer3_outputs(1795);
    layer4_outputs(3868) <= '1';
    layer4_outputs(3869) <= not(layer3_outputs(1046));
    layer4_outputs(3870) <= not(layer3_outputs(2598)) or (layer3_outputs(3744));
    layer4_outputs(3871) <= layer3_outputs(399);
    layer4_outputs(3872) <= not((layer3_outputs(4610)) and (layer3_outputs(4910)));
    layer4_outputs(3873) <= not((layer3_outputs(1205)) xor (layer3_outputs(2960)));
    layer4_outputs(3874) <= not(layer3_outputs(498));
    layer4_outputs(3875) <= (layer3_outputs(2833)) or (layer3_outputs(4383));
    layer4_outputs(3876) <= (layer3_outputs(3861)) and not (layer3_outputs(1986));
    layer4_outputs(3877) <= (layer3_outputs(3780)) and not (layer3_outputs(2692));
    layer4_outputs(3878) <= not((layer3_outputs(853)) xor (layer3_outputs(2738)));
    layer4_outputs(3879) <= not(layer3_outputs(28));
    layer4_outputs(3880) <= not(layer3_outputs(4823));
    layer4_outputs(3881) <= not(layer3_outputs(1548));
    layer4_outputs(3882) <= not(layer3_outputs(2242));
    layer4_outputs(3883) <= not(layer3_outputs(3461));
    layer4_outputs(3884) <= not(layer3_outputs(258));
    layer4_outputs(3885) <= not((layer3_outputs(1803)) or (layer3_outputs(3164)));
    layer4_outputs(3886) <= '0';
    layer4_outputs(3887) <= not(layer3_outputs(292)) or (layer3_outputs(4991));
    layer4_outputs(3888) <= layer3_outputs(560);
    layer4_outputs(3889) <= (layer3_outputs(3814)) and (layer3_outputs(2492));
    layer4_outputs(3890) <= not((layer3_outputs(1552)) or (layer3_outputs(2659)));
    layer4_outputs(3891) <= not(layer3_outputs(2645));
    layer4_outputs(3892) <= '0';
    layer4_outputs(3893) <= layer3_outputs(395);
    layer4_outputs(3894) <= not(layer3_outputs(2742));
    layer4_outputs(3895) <= not(layer3_outputs(3381)) or (layer3_outputs(5004));
    layer4_outputs(3896) <= not((layer3_outputs(4840)) or (layer3_outputs(2791)));
    layer4_outputs(3897) <= not(layer3_outputs(4281));
    layer4_outputs(3898) <= (layer3_outputs(1035)) and (layer3_outputs(780));
    layer4_outputs(3899) <= not(layer3_outputs(2479)) or (layer3_outputs(5025));
    layer4_outputs(3900) <= not((layer3_outputs(3710)) and (layer3_outputs(645)));
    layer4_outputs(3901) <= not((layer3_outputs(4111)) and (layer3_outputs(374)));
    layer4_outputs(3902) <= '1';
    layer4_outputs(3903) <= (layer3_outputs(4193)) or (layer3_outputs(219));
    layer4_outputs(3904) <= not(layer3_outputs(2234));
    layer4_outputs(3905) <= not((layer3_outputs(4863)) xor (layer3_outputs(4360)));
    layer4_outputs(3906) <= layer3_outputs(1919);
    layer4_outputs(3907) <= (layer3_outputs(1265)) and not (layer3_outputs(4015));
    layer4_outputs(3908) <= layer3_outputs(3001);
    layer4_outputs(3909) <= layer3_outputs(4020);
    layer4_outputs(3910) <= layer3_outputs(2998);
    layer4_outputs(3911) <= '0';
    layer4_outputs(3912) <= layer3_outputs(3791);
    layer4_outputs(3913) <= layer3_outputs(1185);
    layer4_outputs(3914) <= not(layer3_outputs(138));
    layer4_outputs(3915) <= (layer3_outputs(4712)) xor (layer3_outputs(2982));
    layer4_outputs(3916) <= not((layer3_outputs(3722)) and (layer3_outputs(3070)));
    layer4_outputs(3917) <= layer3_outputs(3551);
    layer4_outputs(3918) <= (layer3_outputs(526)) xor (layer3_outputs(820));
    layer4_outputs(3919) <= (layer3_outputs(2284)) and not (layer3_outputs(4436));
    layer4_outputs(3920) <= not(layer3_outputs(1792));
    layer4_outputs(3921) <= not(layer3_outputs(2882)) or (layer3_outputs(3264));
    layer4_outputs(3922) <= (layer3_outputs(2103)) and (layer3_outputs(2087));
    layer4_outputs(3923) <= not((layer3_outputs(882)) xor (layer3_outputs(3629)));
    layer4_outputs(3924) <= '0';
    layer4_outputs(3925) <= (layer3_outputs(4996)) and not (layer3_outputs(1152));
    layer4_outputs(3926) <= (layer3_outputs(2282)) xor (layer3_outputs(4180));
    layer4_outputs(3927) <= layer3_outputs(4398);
    layer4_outputs(3928) <= (layer3_outputs(5058)) or (layer3_outputs(1968));
    layer4_outputs(3929) <= layer3_outputs(1395);
    layer4_outputs(3930) <= not((layer3_outputs(3855)) and (layer3_outputs(3383)));
    layer4_outputs(3931) <= layer3_outputs(1132);
    layer4_outputs(3932) <= not(layer3_outputs(187));
    layer4_outputs(3933) <= not(layer3_outputs(3856)) or (layer3_outputs(433));
    layer4_outputs(3934) <= not(layer3_outputs(3283));
    layer4_outputs(3935) <= not((layer3_outputs(4477)) and (layer3_outputs(972)));
    layer4_outputs(3936) <= not(layer3_outputs(3881)) or (layer3_outputs(623));
    layer4_outputs(3937) <= layer3_outputs(3837);
    layer4_outputs(3938) <= '1';
    layer4_outputs(3939) <= layer3_outputs(293);
    layer4_outputs(3940) <= (layer3_outputs(3826)) or (layer3_outputs(1540));
    layer4_outputs(3941) <= not(layer3_outputs(1280));
    layer4_outputs(3942) <= (layer3_outputs(1012)) xor (layer3_outputs(345));
    layer4_outputs(3943) <= '0';
    layer4_outputs(3944) <= (layer3_outputs(5048)) and not (layer3_outputs(4275));
    layer4_outputs(3945) <= layer3_outputs(1092);
    layer4_outputs(3946) <= (layer3_outputs(1172)) and not (layer3_outputs(4868));
    layer4_outputs(3947) <= not(layer3_outputs(3321));
    layer4_outputs(3948) <= (layer3_outputs(968)) and (layer3_outputs(2898));
    layer4_outputs(3949) <= '0';
    layer4_outputs(3950) <= (layer3_outputs(1205)) or (layer3_outputs(1954));
    layer4_outputs(3951) <= (layer3_outputs(1508)) or (layer3_outputs(2806));
    layer4_outputs(3952) <= not((layer3_outputs(4724)) xor (layer3_outputs(3249)));
    layer4_outputs(3953) <= (layer3_outputs(1240)) and (layer3_outputs(1748));
    layer4_outputs(3954) <= not(layer3_outputs(1849));
    layer4_outputs(3955) <= not((layer3_outputs(494)) or (layer3_outputs(746)));
    layer4_outputs(3956) <= '1';
    layer4_outputs(3957) <= '1';
    layer4_outputs(3958) <= (layer3_outputs(2835)) and not (layer3_outputs(4623));
    layer4_outputs(3959) <= layer3_outputs(3586);
    layer4_outputs(3960) <= not((layer3_outputs(4410)) or (layer3_outputs(3530)));
    layer4_outputs(3961) <= (layer3_outputs(3112)) and not (layer3_outputs(3907));
    layer4_outputs(3962) <= not(layer3_outputs(788)) or (layer3_outputs(2508));
    layer4_outputs(3963) <= '0';
    layer4_outputs(3964) <= (layer3_outputs(2735)) and (layer3_outputs(3128));
    layer4_outputs(3965) <= not(layer3_outputs(3201));
    layer4_outputs(3966) <= (layer3_outputs(1309)) and not (layer3_outputs(4622));
    layer4_outputs(3967) <= (layer3_outputs(4830)) and (layer3_outputs(1887));
    layer4_outputs(3968) <= not((layer3_outputs(2536)) and (layer3_outputs(5092)));
    layer4_outputs(3969) <= (layer3_outputs(3504)) and (layer3_outputs(709));
    layer4_outputs(3970) <= '0';
    layer4_outputs(3971) <= (layer3_outputs(3431)) and (layer3_outputs(1007));
    layer4_outputs(3972) <= (layer3_outputs(3295)) and not (layer3_outputs(1876));
    layer4_outputs(3973) <= not(layer3_outputs(1512));
    layer4_outputs(3974) <= layer3_outputs(5028);
    layer4_outputs(3975) <= not(layer3_outputs(1994));
    layer4_outputs(3976) <= not(layer3_outputs(1341));
    layer4_outputs(3977) <= not(layer3_outputs(4435));
    layer4_outputs(3978) <= (layer3_outputs(2710)) and not (layer3_outputs(3773));
    layer4_outputs(3979) <= not(layer3_outputs(3377)) or (layer3_outputs(4933));
    layer4_outputs(3980) <= '1';
    layer4_outputs(3981) <= (layer3_outputs(3667)) and (layer3_outputs(2476));
    layer4_outputs(3982) <= not((layer3_outputs(1006)) and (layer3_outputs(54)));
    layer4_outputs(3983) <= (layer3_outputs(4311)) and (layer3_outputs(448));
    layer4_outputs(3984) <= layer3_outputs(4933);
    layer4_outputs(3985) <= not(layer3_outputs(2644)) or (layer3_outputs(3431));
    layer4_outputs(3986) <= not(layer3_outputs(3016));
    layer4_outputs(3987) <= '0';
    layer4_outputs(3988) <= not(layer3_outputs(2831)) or (layer3_outputs(2696));
    layer4_outputs(3989) <= layer3_outputs(543);
    layer4_outputs(3990) <= layer3_outputs(1988);
    layer4_outputs(3991) <= (layer3_outputs(1115)) and not (layer3_outputs(3976));
    layer4_outputs(3992) <= (layer3_outputs(3682)) and not (layer3_outputs(1676));
    layer4_outputs(3993) <= not((layer3_outputs(4377)) and (layer3_outputs(3190)));
    layer4_outputs(3994) <= not((layer3_outputs(1723)) and (layer3_outputs(895)));
    layer4_outputs(3995) <= layer3_outputs(4182);
    layer4_outputs(3996) <= (layer3_outputs(1888)) and not (layer3_outputs(4852));
    layer4_outputs(3997) <= (layer3_outputs(4296)) and not (layer3_outputs(2383));
    layer4_outputs(3998) <= not(layer3_outputs(1985));
    layer4_outputs(3999) <= '0';
    layer4_outputs(4000) <= not(layer3_outputs(475));
    layer4_outputs(4001) <= not(layer3_outputs(2133));
    layer4_outputs(4002) <= not(layer3_outputs(624));
    layer4_outputs(4003) <= (layer3_outputs(3535)) and not (layer3_outputs(3261));
    layer4_outputs(4004) <= not(layer3_outputs(4705));
    layer4_outputs(4005) <= not(layer3_outputs(2909));
    layer4_outputs(4006) <= not(layer3_outputs(617));
    layer4_outputs(4007) <= '0';
    layer4_outputs(4008) <= (layer3_outputs(1556)) and not (layer3_outputs(1826));
    layer4_outputs(4009) <= layer3_outputs(1992);
    layer4_outputs(4010) <= not(layer3_outputs(818));
    layer4_outputs(4011) <= not((layer3_outputs(1443)) xor (layer3_outputs(3889)));
    layer4_outputs(4012) <= (layer3_outputs(4217)) and not (layer3_outputs(815));
    layer4_outputs(4013) <= not((layer3_outputs(1925)) xor (layer3_outputs(3936)));
    layer4_outputs(4014) <= '0';
    layer4_outputs(4015) <= (layer3_outputs(2702)) and (layer3_outputs(3657));
    layer4_outputs(4016) <= not(layer3_outputs(3553));
    layer4_outputs(4017) <= not(layer3_outputs(2035)) or (layer3_outputs(874));
    layer4_outputs(4018) <= layer3_outputs(316);
    layer4_outputs(4019) <= '1';
    layer4_outputs(4020) <= not(layer3_outputs(2585)) or (layer3_outputs(4426));
    layer4_outputs(4021) <= layer3_outputs(4204);
    layer4_outputs(4022) <= '1';
    layer4_outputs(4023) <= (layer3_outputs(4348)) and not (layer3_outputs(957));
    layer4_outputs(4024) <= not(layer3_outputs(1456));
    layer4_outputs(4025) <= not(layer3_outputs(4224)) or (layer3_outputs(2293));
    layer4_outputs(4026) <= layer3_outputs(1680);
    layer4_outputs(4027) <= not(layer3_outputs(3954)) or (layer3_outputs(1530));
    layer4_outputs(4028) <= layer3_outputs(1424);
    layer4_outputs(4029) <= not(layer3_outputs(3025)) or (layer3_outputs(125));
    layer4_outputs(4030) <= (layer3_outputs(4057)) and not (layer3_outputs(166));
    layer4_outputs(4031) <= not((layer3_outputs(244)) or (layer3_outputs(2157)));
    layer4_outputs(4032) <= not(layer3_outputs(506));
    layer4_outputs(4033) <= not((layer3_outputs(1300)) and (layer3_outputs(4043)));
    layer4_outputs(4034) <= (layer3_outputs(4986)) and (layer3_outputs(1050));
    layer4_outputs(4035) <= not(layer3_outputs(27)) or (layer3_outputs(1898));
    layer4_outputs(4036) <= layer3_outputs(1383);
    layer4_outputs(4037) <= (layer3_outputs(3370)) or (layer3_outputs(85));
    layer4_outputs(4038) <= layer3_outputs(806);
    layer4_outputs(4039) <= layer3_outputs(559);
    layer4_outputs(4040) <= (layer3_outputs(987)) or (layer3_outputs(3127));
    layer4_outputs(4041) <= layer3_outputs(2316);
    layer4_outputs(4042) <= layer3_outputs(3686);
    layer4_outputs(4043) <= layer3_outputs(3656);
    layer4_outputs(4044) <= (layer3_outputs(3475)) or (layer3_outputs(698));
    layer4_outputs(4045) <= not((layer3_outputs(5023)) xor (layer3_outputs(3323)));
    layer4_outputs(4046) <= layer3_outputs(3346);
    layer4_outputs(4047) <= (layer3_outputs(3593)) and (layer3_outputs(3549));
    layer4_outputs(4048) <= (layer3_outputs(3002)) and not (layer3_outputs(2551));
    layer4_outputs(4049) <= not(layer3_outputs(1416));
    layer4_outputs(4050) <= layer3_outputs(3488);
    layer4_outputs(4051) <= not(layer3_outputs(4914));
    layer4_outputs(4052) <= (layer3_outputs(580)) and not (layer3_outputs(1503));
    layer4_outputs(4053) <= not(layer3_outputs(878)) or (layer3_outputs(682));
    layer4_outputs(4054) <= not(layer3_outputs(872)) or (layer3_outputs(2657));
    layer4_outputs(4055) <= layer3_outputs(4323);
    layer4_outputs(4056) <= not(layer3_outputs(2522));
    layer4_outputs(4057) <= (layer3_outputs(792)) and (layer3_outputs(1900));
    layer4_outputs(4058) <= layer3_outputs(3616);
    layer4_outputs(4059) <= not(layer3_outputs(4732));
    layer4_outputs(4060) <= not(layer3_outputs(366)) or (layer3_outputs(1561));
    layer4_outputs(4061) <= layer3_outputs(1769);
    layer4_outputs(4062) <= not(layer3_outputs(3843));
    layer4_outputs(4063) <= not(layer3_outputs(2800)) or (layer3_outputs(2594));
    layer4_outputs(4064) <= layer3_outputs(74);
    layer4_outputs(4065) <= layer3_outputs(4865);
    layer4_outputs(4066) <= not(layer3_outputs(237)) or (layer3_outputs(4486));
    layer4_outputs(4067) <= (layer3_outputs(1706)) or (layer3_outputs(4992));
    layer4_outputs(4068) <= not((layer3_outputs(5094)) and (layer3_outputs(3894)));
    layer4_outputs(4069) <= '0';
    layer4_outputs(4070) <= (layer3_outputs(2730)) or (layer3_outputs(70));
    layer4_outputs(4071) <= (layer3_outputs(3489)) and not (layer3_outputs(4946));
    layer4_outputs(4072) <= (layer3_outputs(25)) and not (layer3_outputs(2815));
    layer4_outputs(4073) <= (layer3_outputs(3305)) and (layer3_outputs(3752));
    layer4_outputs(4074) <= (layer3_outputs(3651)) or (layer3_outputs(4061));
    layer4_outputs(4075) <= '1';
    layer4_outputs(4076) <= layer3_outputs(1042);
    layer4_outputs(4077) <= (layer3_outputs(2566)) xor (layer3_outputs(183));
    layer4_outputs(4078) <= not((layer3_outputs(1017)) xor (layer3_outputs(1757)));
    layer4_outputs(4079) <= not((layer3_outputs(553)) and (layer3_outputs(1535)));
    layer4_outputs(4080) <= not(layer3_outputs(2458));
    layer4_outputs(4081) <= (layer3_outputs(3246)) and (layer3_outputs(2041));
    layer4_outputs(4082) <= layer3_outputs(4885);
    layer4_outputs(4083) <= layer3_outputs(1332);
    layer4_outputs(4084) <= layer3_outputs(3847);
    layer4_outputs(4085) <= layer3_outputs(3327);
    layer4_outputs(4086) <= (layer3_outputs(4325)) and (layer3_outputs(3190));
    layer4_outputs(4087) <= layer3_outputs(1119);
    layer4_outputs(4088) <= (layer3_outputs(4514)) xor (layer3_outputs(113));
    layer4_outputs(4089) <= layer3_outputs(1475);
    layer4_outputs(4090) <= layer3_outputs(4561);
    layer4_outputs(4091) <= not((layer3_outputs(2924)) and (layer3_outputs(660)));
    layer4_outputs(4092) <= not((layer3_outputs(396)) or (layer3_outputs(2911)));
    layer4_outputs(4093) <= not((layer3_outputs(2086)) and (layer3_outputs(1604)));
    layer4_outputs(4094) <= not((layer3_outputs(4961)) xor (layer3_outputs(4127)));
    layer4_outputs(4095) <= layer3_outputs(4686);
    layer4_outputs(4096) <= (layer3_outputs(5042)) and not (layer3_outputs(4338));
    layer4_outputs(4097) <= layer3_outputs(2998);
    layer4_outputs(4098) <= (layer3_outputs(3231)) and not (layer3_outputs(3896));
    layer4_outputs(4099) <= layer3_outputs(5110);
    layer4_outputs(4100) <= not(layer3_outputs(522));
    layer4_outputs(4101) <= (layer3_outputs(3762)) and not (layer3_outputs(4156));
    layer4_outputs(4102) <= (layer3_outputs(101)) and (layer3_outputs(20));
    layer4_outputs(4103) <= not((layer3_outputs(4623)) and (layer3_outputs(4695)));
    layer4_outputs(4104) <= layer3_outputs(4611);
    layer4_outputs(4105) <= layer3_outputs(1840);
    layer4_outputs(4106) <= not(layer3_outputs(4374));
    layer4_outputs(4107) <= (layer3_outputs(598)) and not (layer3_outputs(2185));
    layer4_outputs(4108) <= layer3_outputs(4963);
    layer4_outputs(4109) <= not(layer3_outputs(3172));
    layer4_outputs(4110) <= layer3_outputs(814);
    layer4_outputs(4111) <= layer3_outputs(640);
    layer4_outputs(4112) <= '1';
    layer4_outputs(4113) <= not((layer3_outputs(3666)) and (layer3_outputs(3608)));
    layer4_outputs(4114) <= (layer3_outputs(2588)) and not (layer3_outputs(4131));
    layer4_outputs(4115) <= (layer3_outputs(2084)) and (layer3_outputs(3736));
    layer4_outputs(4116) <= not(layer3_outputs(4535)) or (layer3_outputs(3375));
    layer4_outputs(4117) <= not((layer3_outputs(2225)) and (layer3_outputs(4469)));
    layer4_outputs(4118) <= not((layer3_outputs(4230)) xor (layer3_outputs(1098)));
    layer4_outputs(4119) <= (layer3_outputs(3035)) and not (layer3_outputs(5117));
    layer4_outputs(4120) <= layer3_outputs(2599);
    layer4_outputs(4121) <= (layer3_outputs(4150)) and not (layer3_outputs(255));
    layer4_outputs(4122) <= (layer3_outputs(2730)) and not (layer3_outputs(542));
    layer4_outputs(4123) <= layer3_outputs(3683);
    layer4_outputs(4124) <= (layer3_outputs(457)) or (layer3_outputs(3858));
    layer4_outputs(4125) <= '0';
    layer4_outputs(4126) <= not(layer3_outputs(1032));
    layer4_outputs(4127) <= not(layer3_outputs(1366)) or (layer3_outputs(5079));
    layer4_outputs(4128) <= layer3_outputs(3193);
    layer4_outputs(4129) <= layer3_outputs(2823);
    layer4_outputs(4130) <= layer3_outputs(2035);
    layer4_outputs(4131) <= not(layer3_outputs(3487));
    layer4_outputs(4132) <= layer3_outputs(2336);
    layer4_outputs(4133) <= '0';
    layer4_outputs(4134) <= not(layer3_outputs(4487));
    layer4_outputs(4135) <= not((layer3_outputs(3679)) or (layer3_outputs(3345)));
    layer4_outputs(4136) <= layer3_outputs(4290);
    layer4_outputs(4137) <= (layer3_outputs(1472)) and (layer3_outputs(2322));
    layer4_outputs(4138) <= not((layer3_outputs(3801)) or (layer3_outputs(3447)));
    layer4_outputs(4139) <= not(layer3_outputs(4918));
    layer4_outputs(4140) <= (layer3_outputs(1675)) and (layer3_outputs(1357));
    layer4_outputs(4141) <= layer3_outputs(3663);
    layer4_outputs(4142) <= not((layer3_outputs(2185)) and (layer3_outputs(4374)));
    layer4_outputs(4143) <= not(layer3_outputs(2827));
    layer4_outputs(4144) <= not(layer3_outputs(4034));
    layer4_outputs(4145) <= not((layer3_outputs(2991)) and (layer3_outputs(3806)));
    layer4_outputs(4146) <= '1';
    layer4_outputs(4147) <= not(layer3_outputs(1507)) or (layer3_outputs(1567));
    layer4_outputs(4148) <= '1';
    layer4_outputs(4149) <= (layer3_outputs(3811)) and (layer3_outputs(4948));
    layer4_outputs(4150) <= '1';
    layer4_outputs(4151) <= (layer3_outputs(2189)) xor (layer3_outputs(2555));
    layer4_outputs(4152) <= '0';
    layer4_outputs(4153) <= layer3_outputs(1340);
    layer4_outputs(4154) <= (layer3_outputs(2272)) or (layer3_outputs(282));
    layer4_outputs(4155) <= not((layer3_outputs(2171)) and (layer3_outputs(1199)));
    layer4_outputs(4156) <= layer3_outputs(3733);
    layer4_outputs(4157) <= not(layer3_outputs(4337));
    layer4_outputs(4158) <= (layer3_outputs(2612)) xor (layer3_outputs(2298));
    layer4_outputs(4159) <= not(layer3_outputs(350));
    layer4_outputs(4160) <= not(layer3_outputs(3654));
    layer4_outputs(4161) <= layer3_outputs(799);
    layer4_outputs(4162) <= not(layer3_outputs(135));
    layer4_outputs(4163) <= not(layer3_outputs(5108));
    layer4_outputs(4164) <= '0';
    layer4_outputs(4165) <= (layer3_outputs(4924)) and (layer3_outputs(4474));
    layer4_outputs(4166) <= '0';
    layer4_outputs(4167) <= not(layer3_outputs(940));
    layer4_outputs(4168) <= not((layer3_outputs(2988)) or (layer3_outputs(2841)));
    layer4_outputs(4169) <= not(layer3_outputs(368));
    layer4_outputs(4170) <= (layer3_outputs(838)) and not (layer3_outputs(2245));
    layer4_outputs(4171) <= not((layer3_outputs(4509)) xor (layer3_outputs(3758)));
    layer4_outputs(4172) <= '0';
    layer4_outputs(4173) <= not(layer3_outputs(544)) or (layer3_outputs(2365));
    layer4_outputs(4174) <= layer3_outputs(4117);
    layer4_outputs(4175) <= '1';
    layer4_outputs(4176) <= not(layer3_outputs(2485));
    layer4_outputs(4177) <= (layer3_outputs(2024)) and (layer3_outputs(1537));
    layer4_outputs(4178) <= not(layer3_outputs(2408));
    layer4_outputs(4179) <= layer3_outputs(2357);
    layer4_outputs(4180) <= (layer3_outputs(4296)) and not (layer3_outputs(1286));
    layer4_outputs(4181) <= (layer3_outputs(1347)) and (layer3_outputs(4040));
    layer4_outputs(4182) <= (layer3_outputs(1246)) or (layer3_outputs(169));
    layer4_outputs(4183) <= '1';
    layer4_outputs(4184) <= not(layer3_outputs(2531));
    layer4_outputs(4185) <= (layer3_outputs(1469)) and (layer3_outputs(4425));
    layer4_outputs(4186) <= '1';
    layer4_outputs(4187) <= (layer3_outputs(4126)) and not (layer3_outputs(3712));
    layer4_outputs(4188) <= not(layer3_outputs(1639)) or (layer3_outputs(1200));
    layer4_outputs(4189) <= (layer3_outputs(1539)) and not (layer3_outputs(3796));
    layer4_outputs(4190) <= (layer3_outputs(417)) and (layer3_outputs(3018));
    layer4_outputs(4191) <= (layer3_outputs(5030)) and not (layer3_outputs(1649));
    layer4_outputs(4192) <= layer3_outputs(4502);
    layer4_outputs(4193) <= (layer3_outputs(3951)) and (layer3_outputs(19));
    layer4_outputs(4194) <= layer3_outputs(1775);
    layer4_outputs(4195) <= not(layer3_outputs(1484));
    layer4_outputs(4196) <= (layer3_outputs(354)) and not (layer3_outputs(3155));
    layer4_outputs(4197) <= (layer3_outputs(2327)) or (layer3_outputs(57));
    layer4_outputs(4198) <= layer3_outputs(3858);
    layer4_outputs(4199) <= layer3_outputs(4719);
    layer4_outputs(4200) <= not((layer3_outputs(3577)) xor (layer3_outputs(4793)));
    layer4_outputs(4201) <= not(layer3_outputs(700));
    layer4_outputs(4202) <= not(layer3_outputs(2775));
    layer4_outputs(4203) <= layer3_outputs(4226);
    layer4_outputs(4204) <= layer3_outputs(229);
    layer4_outputs(4205) <= not((layer3_outputs(3024)) or (layer3_outputs(2140)));
    layer4_outputs(4206) <= not(layer3_outputs(4963));
    layer4_outputs(4207) <= not(layer3_outputs(1063));
    layer4_outputs(4208) <= not(layer3_outputs(4603));
    layer4_outputs(4209) <= (layer3_outputs(3302)) and not (layer3_outputs(1432));
    layer4_outputs(4210) <= not(layer3_outputs(310));
    layer4_outputs(4211) <= not(layer3_outputs(4470));
    layer4_outputs(4212) <= (layer3_outputs(1505)) and (layer3_outputs(5109));
    layer4_outputs(4213) <= (layer3_outputs(4693)) xor (layer3_outputs(2374));
    layer4_outputs(4214) <= '1';
    layer4_outputs(4215) <= not(layer3_outputs(4569));
    layer4_outputs(4216) <= (layer3_outputs(4664)) and not (layer3_outputs(3218));
    layer4_outputs(4217) <= layer3_outputs(2855);
    layer4_outputs(4218) <= not(layer3_outputs(177));
    layer4_outputs(4219) <= not((layer3_outputs(4419)) and (layer3_outputs(447)));
    layer4_outputs(4220) <= not((layer3_outputs(2372)) xor (layer3_outputs(4712)));
    layer4_outputs(4221) <= layer3_outputs(3896);
    layer4_outputs(4222) <= not((layer3_outputs(897)) and (layer3_outputs(1520)));
    layer4_outputs(4223) <= not((layer3_outputs(830)) and (layer3_outputs(413)));
    layer4_outputs(4224) <= not(layer3_outputs(1250)) or (layer3_outputs(4496));
    layer4_outputs(4225) <= not(layer3_outputs(2246));
    layer4_outputs(4226) <= '0';
    layer4_outputs(4227) <= '1';
    layer4_outputs(4228) <= not((layer3_outputs(1174)) and (layer3_outputs(2745)));
    layer4_outputs(4229) <= '0';
    layer4_outputs(4230) <= '1';
    layer4_outputs(4231) <= '0';
    layer4_outputs(4232) <= not((layer3_outputs(1522)) xor (layer3_outputs(3632)));
    layer4_outputs(4233) <= '0';
    layer4_outputs(4234) <= not(layer3_outputs(4159));
    layer4_outputs(4235) <= not((layer3_outputs(1364)) and (layer3_outputs(3272)));
    layer4_outputs(4236) <= not(layer3_outputs(1051));
    layer4_outputs(4237) <= (layer3_outputs(2352)) and not (layer3_outputs(1411));
    layer4_outputs(4238) <= (layer3_outputs(2155)) or (layer3_outputs(4277));
    layer4_outputs(4239) <= layer3_outputs(2180);
    layer4_outputs(4240) <= not(layer3_outputs(4841));
    layer4_outputs(4241) <= (layer3_outputs(5069)) xor (layer3_outputs(2905));
    layer4_outputs(4242) <= not(layer3_outputs(1703));
    layer4_outputs(4243) <= layer3_outputs(2094);
    layer4_outputs(4244) <= (layer3_outputs(611)) and (layer3_outputs(4851));
    layer4_outputs(4245) <= layer3_outputs(2475);
    layer4_outputs(4246) <= not(layer3_outputs(1742));
    layer4_outputs(4247) <= not(layer3_outputs(3604));
    layer4_outputs(4248) <= '1';
    layer4_outputs(4249) <= layer3_outputs(468);
    layer4_outputs(4250) <= layer3_outputs(4351);
    layer4_outputs(4251) <= (layer3_outputs(2304)) and (layer3_outputs(3188));
    layer4_outputs(4252) <= layer3_outputs(3878);
    layer4_outputs(4253) <= (layer3_outputs(4792)) or (layer3_outputs(1031));
    layer4_outputs(4254) <= not(layer3_outputs(3097));
    layer4_outputs(4255) <= not(layer3_outputs(134));
    layer4_outputs(4256) <= not(layer3_outputs(3332));
    layer4_outputs(4257) <= (layer3_outputs(2931)) and not (layer3_outputs(2277));
    layer4_outputs(4258) <= layer3_outputs(117);
    layer4_outputs(4259) <= layer3_outputs(1049);
    layer4_outputs(4260) <= not(layer3_outputs(2082));
    layer4_outputs(4261) <= layer3_outputs(3202);
    layer4_outputs(4262) <= (layer3_outputs(4966)) and (layer3_outputs(1482));
    layer4_outputs(4263) <= (layer3_outputs(1427)) and not (layer3_outputs(3155));
    layer4_outputs(4264) <= (layer3_outputs(295)) and not (layer3_outputs(3664));
    layer4_outputs(4265) <= not(layer3_outputs(4601));
    layer4_outputs(4266) <= not((layer3_outputs(190)) and (layer3_outputs(4051)));
    layer4_outputs(4267) <= not((layer3_outputs(3041)) xor (layer3_outputs(2099)));
    layer4_outputs(4268) <= '0';
    layer4_outputs(4269) <= layer3_outputs(364);
    layer4_outputs(4270) <= not((layer3_outputs(4854)) and (layer3_outputs(1505)));
    layer4_outputs(4271) <= not(layer3_outputs(5018)) or (layer3_outputs(1510));
    layer4_outputs(4272) <= layer3_outputs(425);
    layer4_outputs(4273) <= not(layer3_outputs(821));
    layer4_outputs(4274) <= (layer3_outputs(4020)) xor (layer3_outputs(3114));
    layer4_outputs(4275) <= not((layer3_outputs(567)) xor (layer3_outputs(2957)));
    layer4_outputs(4276) <= not((layer3_outputs(4081)) or (layer3_outputs(653)));
    layer4_outputs(4277) <= layer3_outputs(1993);
    layer4_outputs(4278) <= not(layer3_outputs(1747));
    layer4_outputs(4279) <= not(layer3_outputs(775));
    layer4_outputs(4280) <= not((layer3_outputs(3360)) and (layer3_outputs(1024)));
    layer4_outputs(4281) <= not((layer3_outputs(3813)) and (layer3_outputs(601)));
    layer4_outputs(4282) <= not(layer3_outputs(2669));
    layer4_outputs(4283) <= layer3_outputs(2289);
    layer4_outputs(4284) <= not(layer3_outputs(2914)) or (layer3_outputs(2068));
    layer4_outputs(4285) <= (layer3_outputs(1834)) xor (layer3_outputs(164));
    layer4_outputs(4286) <= '0';
    layer4_outputs(4287) <= layer3_outputs(552);
    layer4_outputs(4288) <= not(layer3_outputs(3920));
    layer4_outputs(4289) <= layer3_outputs(1986);
    layer4_outputs(4290) <= not(layer3_outputs(3435));
    layer4_outputs(4291) <= not(layer3_outputs(760));
    layer4_outputs(4292) <= layer3_outputs(2565);
    layer4_outputs(4293) <= (layer3_outputs(1163)) and not (layer3_outputs(3355));
    layer4_outputs(4294) <= layer3_outputs(3626);
    layer4_outputs(4295) <= layer3_outputs(5027);
    layer4_outputs(4296) <= layer3_outputs(3277);
    layer4_outputs(4297) <= '1';
    layer4_outputs(4298) <= (layer3_outputs(1)) and (layer3_outputs(549));
    layer4_outputs(4299) <= (layer3_outputs(775)) and (layer3_outputs(4316));
    layer4_outputs(4300) <= not((layer3_outputs(788)) xor (layer3_outputs(4456)));
    layer4_outputs(4301) <= layer3_outputs(2477);
    layer4_outputs(4302) <= (layer3_outputs(3160)) and not (layer3_outputs(1611));
    layer4_outputs(4303) <= layer3_outputs(3819);
    layer4_outputs(4304) <= '1';
    layer4_outputs(4305) <= layer3_outputs(2416);
    layer4_outputs(4306) <= layer3_outputs(89);
    layer4_outputs(4307) <= not(layer3_outputs(2586));
    layer4_outputs(4308) <= layer3_outputs(2778);
    layer4_outputs(4309) <= (layer3_outputs(716)) and (layer3_outputs(4139));
    layer4_outputs(4310) <= not(layer3_outputs(1298));
    layer4_outputs(4311) <= not((layer3_outputs(4266)) or (layer3_outputs(4497)));
    layer4_outputs(4312) <= not(layer3_outputs(4275));
    layer4_outputs(4313) <= '0';
    layer4_outputs(4314) <= not(layer3_outputs(4798)) or (layer3_outputs(2554));
    layer4_outputs(4315) <= '0';
    layer4_outputs(4316) <= not(layer3_outputs(4868));
    layer4_outputs(4317) <= not(layer3_outputs(2192));
    layer4_outputs(4318) <= not(layer3_outputs(2837));
    layer4_outputs(4319) <= not(layer3_outputs(435));
    layer4_outputs(4320) <= not(layer3_outputs(1855));
    layer4_outputs(4321) <= not(layer3_outputs(976));
    layer4_outputs(4322) <= (layer3_outputs(4962)) and (layer3_outputs(1126));
    layer4_outputs(4323) <= (layer3_outputs(544)) and not (layer3_outputs(1114));
    layer4_outputs(4324) <= layer3_outputs(909);
    layer4_outputs(4325) <= (layer3_outputs(2224)) or (layer3_outputs(1847));
    layer4_outputs(4326) <= layer3_outputs(3927);
    layer4_outputs(4327) <= '0';
    layer4_outputs(4328) <= layer3_outputs(1780);
    layer4_outputs(4329) <= not(layer3_outputs(54));
    layer4_outputs(4330) <= (layer3_outputs(1075)) and not (layer3_outputs(423));
    layer4_outputs(4331) <= not(layer3_outputs(228));
    layer4_outputs(4332) <= not(layer3_outputs(451));
    layer4_outputs(4333) <= (layer3_outputs(4807)) and not (layer3_outputs(2342));
    layer4_outputs(4334) <= '0';
    layer4_outputs(4335) <= not((layer3_outputs(3850)) and (layer3_outputs(4021)));
    layer4_outputs(4336) <= '0';
    layer4_outputs(4337) <= (layer3_outputs(4597)) or (layer3_outputs(3621));
    layer4_outputs(4338) <= layer3_outputs(2955);
    layer4_outputs(4339) <= not((layer3_outputs(963)) xor (layer3_outputs(1798)));
    layer4_outputs(4340) <= layer3_outputs(1046);
    layer4_outputs(4341) <= not(layer3_outputs(895)) or (layer3_outputs(4444));
    layer4_outputs(4342) <= not((layer3_outputs(1923)) or (layer3_outputs(1698)));
    layer4_outputs(4343) <= (layer3_outputs(3476)) or (layer3_outputs(672));
    layer4_outputs(4344) <= not(layer3_outputs(547));
    layer4_outputs(4345) <= layer3_outputs(3062);
    layer4_outputs(4346) <= '0';
    layer4_outputs(4347) <= not(layer3_outputs(4262));
    layer4_outputs(4348) <= not(layer3_outputs(3381));
    layer4_outputs(4349) <= not((layer3_outputs(3993)) or (layer3_outputs(873)));
    layer4_outputs(4350) <= not(layer3_outputs(2830));
    layer4_outputs(4351) <= layer3_outputs(1580);
    layer4_outputs(4352) <= layer3_outputs(2534);
    layer4_outputs(4353) <= (layer3_outputs(4079)) and (layer3_outputs(1936));
    layer4_outputs(4354) <= not(layer3_outputs(883));
    layer4_outputs(4355) <= not(layer3_outputs(3016));
    layer4_outputs(4356) <= (layer3_outputs(3874)) and (layer3_outputs(231));
    layer4_outputs(4357) <= (layer3_outputs(1377)) and not (layer3_outputs(3797));
    layer4_outputs(4358) <= (layer3_outputs(4174)) or (layer3_outputs(75));
    layer4_outputs(4359) <= not((layer3_outputs(4319)) or (layer3_outputs(4944)));
    layer4_outputs(4360) <= layer3_outputs(4822);
    layer4_outputs(4361) <= (layer3_outputs(2114)) or (layer3_outputs(354));
    layer4_outputs(4362) <= not(layer3_outputs(3732));
    layer4_outputs(4363) <= not(layer3_outputs(2406));
    layer4_outputs(4364) <= not(layer3_outputs(1916));
    layer4_outputs(4365) <= not((layer3_outputs(3863)) or (layer3_outputs(1571)));
    layer4_outputs(4366) <= (layer3_outputs(374)) or (layer3_outputs(871));
    layer4_outputs(4367) <= not(layer3_outputs(4186));
    layer4_outputs(4368) <= (layer3_outputs(4473)) or (layer3_outputs(1433));
    layer4_outputs(4369) <= not(layer3_outputs(4891));
    layer4_outputs(4370) <= not((layer3_outputs(3703)) or (layer3_outputs(1756)));
    layer4_outputs(4371) <= not(layer3_outputs(1317)) or (layer3_outputs(2287));
    layer4_outputs(4372) <= layer3_outputs(3477);
    layer4_outputs(4373) <= layer3_outputs(680);
    layer4_outputs(4374) <= (layer3_outputs(569)) and (layer3_outputs(4781));
    layer4_outputs(4375) <= (layer3_outputs(3263)) and not (layer3_outputs(4302));
    layer4_outputs(4376) <= not((layer3_outputs(724)) or (layer3_outputs(2587)));
    layer4_outputs(4377) <= (layer3_outputs(2448)) and not (layer3_outputs(66));
    layer4_outputs(4378) <= not((layer3_outputs(3483)) and (layer3_outputs(2936)));
    layer4_outputs(4379) <= not(layer3_outputs(1845));
    layer4_outputs(4380) <= layer3_outputs(4653);
    layer4_outputs(4381) <= (layer3_outputs(2081)) xor (layer3_outputs(4639));
    layer4_outputs(4382) <= layer3_outputs(2043);
    layer4_outputs(4383) <= not(layer3_outputs(1556));
    layer4_outputs(4384) <= not(layer3_outputs(2779));
    layer4_outputs(4385) <= layer3_outputs(906);
    layer4_outputs(4386) <= layer3_outputs(267);
    layer4_outputs(4387) <= not(layer3_outputs(3869));
    layer4_outputs(4388) <= (layer3_outputs(1344)) and not (layer3_outputs(3422));
    layer4_outputs(4389) <= not(layer3_outputs(1399));
    layer4_outputs(4390) <= (layer3_outputs(1479)) and (layer3_outputs(1367));
    layer4_outputs(4391) <= not((layer3_outputs(204)) and (layer3_outputs(1227)));
    layer4_outputs(4392) <= (layer3_outputs(4584)) or (layer3_outputs(204));
    layer4_outputs(4393) <= layer3_outputs(4853);
    layer4_outputs(4394) <= (layer3_outputs(4265)) xor (layer3_outputs(3118));
    layer4_outputs(4395) <= not((layer3_outputs(3475)) or (layer3_outputs(2069)));
    layer4_outputs(4396) <= layer3_outputs(1462);
    layer4_outputs(4397) <= not(layer3_outputs(2921));
    layer4_outputs(4398) <= not((layer3_outputs(716)) and (layer3_outputs(2527)));
    layer4_outputs(4399) <= layer3_outputs(309);
    layer4_outputs(4400) <= layer3_outputs(2985);
    layer4_outputs(4401) <= not(layer3_outputs(398));
    layer4_outputs(4402) <= layer3_outputs(2502);
    layer4_outputs(4403) <= layer3_outputs(1328);
    layer4_outputs(4404) <= not(layer3_outputs(503)) or (layer3_outputs(1885));
    layer4_outputs(4405) <= not(layer3_outputs(3670)) or (layer3_outputs(5099));
    layer4_outputs(4406) <= not(layer3_outputs(3925));
    layer4_outputs(4407) <= not(layer3_outputs(4894));
    layer4_outputs(4408) <= layer3_outputs(3631);
    layer4_outputs(4409) <= (layer3_outputs(4003)) or (layer3_outputs(2477));
    layer4_outputs(4410) <= (layer3_outputs(1333)) and (layer3_outputs(1337));
    layer4_outputs(4411) <= '1';
    layer4_outputs(4412) <= (layer3_outputs(1463)) and not (layer3_outputs(4812));
    layer4_outputs(4413) <= not(layer3_outputs(3934));
    layer4_outputs(4414) <= (layer3_outputs(4013)) or (layer3_outputs(4922));
    layer4_outputs(4415) <= layer3_outputs(1286);
    layer4_outputs(4416) <= not((layer3_outputs(4339)) and (layer3_outputs(2595)));
    layer4_outputs(4417) <= not(layer3_outputs(3809));
    layer4_outputs(4418) <= not(layer3_outputs(1116));
    layer4_outputs(4419) <= not(layer3_outputs(4142)) or (layer3_outputs(1511));
    layer4_outputs(4420) <= '0';
    layer4_outputs(4421) <= not((layer3_outputs(1668)) and (layer3_outputs(482)));
    layer4_outputs(4422) <= '0';
    layer4_outputs(4423) <= not((layer3_outputs(4903)) xor (layer3_outputs(1094)));
    layer4_outputs(4424) <= not((layer3_outputs(1186)) xor (layer3_outputs(2484)));
    layer4_outputs(4425) <= not(layer3_outputs(1341));
    layer4_outputs(4426) <= not(layer3_outputs(2409));
    layer4_outputs(4427) <= (layer3_outputs(4489)) and (layer3_outputs(4501));
    layer4_outputs(4428) <= not(layer3_outputs(2754));
    layer4_outputs(4429) <= layer3_outputs(2285);
    layer4_outputs(4430) <= (layer3_outputs(3659)) and not (layer3_outputs(4108));
    layer4_outputs(4431) <= not((layer3_outputs(2579)) or (layer3_outputs(3162)));
    layer4_outputs(4432) <= not((layer3_outputs(2454)) or (layer3_outputs(3888)));
    layer4_outputs(4433) <= layer3_outputs(4543);
    layer4_outputs(4434) <= not((layer3_outputs(1536)) xor (layer3_outputs(1423)));
    layer4_outputs(4435) <= (layer3_outputs(324)) and (layer3_outputs(3193));
    layer4_outputs(4436) <= layer3_outputs(5074);
    layer4_outputs(4437) <= (layer3_outputs(1815)) or (layer3_outputs(1013));
    layer4_outputs(4438) <= layer3_outputs(3938);
    layer4_outputs(4439) <= layer3_outputs(1410);
    layer4_outputs(4440) <= '1';
    layer4_outputs(4441) <= layer3_outputs(2761);
    layer4_outputs(4442) <= not((layer3_outputs(1085)) and (layer3_outputs(3466)));
    layer4_outputs(4443) <= not(layer3_outputs(2871));
    layer4_outputs(4444) <= not(layer3_outputs(4953));
    layer4_outputs(4445) <= not(layer3_outputs(2712)) or (layer3_outputs(1879));
    layer4_outputs(4446) <= not(layer3_outputs(4916));
    layer4_outputs(4447) <= not((layer3_outputs(870)) and (layer3_outputs(2773)));
    layer4_outputs(4448) <= (layer3_outputs(1422)) and (layer3_outputs(4344));
    layer4_outputs(4449) <= layer3_outputs(1754);
    layer4_outputs(4450) <= layer3_outputs(4667);
    layer4_outputs(4451) <= layer3_outputs(2046);
    layer4_outputs(4452) <= not((layer3_outputs(4760)) or (layer3_outputs(3383)));
    layer4_outputs(4453) <= not(layer3_outputs(4464));
    layer4_outputs(4454) <= layer3_outputs(392);
    layer4_outputs(4455) <= not(layer3_outputs(1600));
    layer4_outputs(4456) <= layer3_outputs(4126);
    layer4_outputs(4457) <= (layer3_outputs(5026)) xor (layer3_outputs(3296));
    layer4_outputs(4458) <= not((layer3_outputs(4745)) and (layer3_outputs(3037)));
    layer4_outputs(4459) <= (layer3_outputs(3400)) and not (layer3_outputs(4132));
    layer4_outputs(4460) <= not((layer3_outputs(109)) or (layer3_outputs(3012)));
    layer4_outputs(4461) <= layer3_outputs(2561);
    layer4_outputs(4462) <= not(layer3_outputs(3675));
    layer4_outputs(4463) <= '1';
    layer4_outputs(4464) <= not(layer3_outputs(3121));
    layer4_outputs(4465) <= (layer3_outputs(3662)) and (layer3_outputs(4290));
    layer4_outputs(4466) <= layer3_outputs(700);
    layer4_outputs(4467) <= '0';
    layer4_outputs(4468) <= not(layer3_outputs(113));
    layer4_outputs(4469) <= not((layer3_outputs(974)) or (layer3_outputs(891)));
    layer4_outputs(4470) <= layer3_outputs(1393);
    layer4_outputs(4471) <= not(layer3_outputs(1472));
    layer4_outputs(4472) <= layer3_outputs(3901);
    layer4_outputs(4473) <= not(layer3_outputs(823)) or (layer3_outputs(3777));
    layer4_outputs(4474) <= (layer3_outputs(226)) and not (layer3_outputs(261));
    layer4_outputs(4475) <= not((layer3_outputs(3537)) or (layer3_outputs(2307)));
    layer4_outputs(4476) <= not((layer3_outputs(2233)) and (layer3_outputs(669)));
    layer4_outputs(4477) <= not(layer3_outputs(2164));
    layer4_outputs(4478) <= '0';
    layer4_outputs(4479) <= not(layer3_outputs(382));
    layer4_outputs(4480) <= not(layer3_outputs(862));
    layer4_outputs(4481) <= layer3_outputs(3668);
    layer4_outputs(4482) <= (layer3_outputs(1714)) and not (layer3_outputs(2280));
    layer4_outputs(4483) <= not(layer3_outputs(1389));
    layer4_outputs(4484) <= not(layer3_outputs(3126));
    layer4_outputs(4485) <= not(layer3_outputs(2195));
    layer4_outputs(4486) <= not(layer3_outputs(2732));
    layer4_outputs(4487) <= (layer3_outputs(568)) or (layer3_outputs(1591));
    layer4_outputs(4488) <= not((layer3_outputs(4347)) or (layer3_outputs(148)));
    layer4_outputs(4489) <= (layer3_outputs(2875)) and (layer3_outputs(1155));
    layer4_outputs(4490) <= not(layer3_outputs(711));
    layer4_outputs(4491) <= (layer3_outputs(914)) or (layer3_outputs(361));
    layer4_outputs(4492) <= not((layer3_outputs(3040)) or (layer3_outputs(3288)));
    layer4_outputs(4493) <= layer3_outputs(4211);
    layer4_outputs(4494) <= not(layer3_outputs(1779));
    layer4_outputs(4495) <= not(layer3_outputs(3854));
    layer4_outputs(4496) <= (layer3_outputs(2663)) and not (layer3_outputs(994));
    layer4_outputs(4497) <= (layer3_outputs(3681)) and not (layer3_outputs(1301));
    layer4_outputs(4498) <= '1';
    layer4_outputs(4499) <= '0';
    layer4_outputs(4500) <= not(layer3_outputs(1391));
    layer4_outputs(4501) <= not(layer3_outputs(2806)) or (layer3_outputs(3513));
    layer4_outputs(4502) <= not(layer3_outputs(768));
    layer4_outputs(4503) <= '1';
    layer4_outputs(4504) <= '0';
    layer4_outputs(4505) <= not(layer3_outputs(4147)) or (layer3_outputs(4985));
    layer4_outputs(4506) <= '1';
    layer4_outputs(4507) <= not(layer3_outputs(1465)) or (layer3_outputs(1515));
    layer4_outputs(4508) <= not(layer3_outputs(1036)) or (layer3_outputs(4248));
    layer4_outputs(4509) <= not((layer3_outputs(3280)) xor (layer3_outputs(3150)));
    layer4_outputs(4510) <= layer3_outputs(3936);
    layer4_outputs(4511) <= (layer3_outputs(3982)) or (layer3_outputs(1717));
    layer4_outputs(4512) <= layer3_outputs(1581);
    layer4_outputs(4513) <= not(layer3_outputs(3731));
    layer4_outputs(4514) <= layer3_outputs(1019);
    layer4_outputs(4515) <= (layer3_outputs(2707)) and not (layer3_outputs(4022));
    layer4_outputs(4516) <= (layer3_outputs(230)) and (layer3_outputs(3389));
    layer4_outputs(4517) <= (layer3_outputs(4536)) and not (layer3_outputs(3184));
    layer4_outputs(4518) <= not(layer3_outputs(1853)) or (layer3_outputs(4008));
    layer4_outputs(4519) <= '1';
    layer4_outputs(4520) <= (layer3_outputs(3618)) and (layer3_outputs(1425));
    layer4_outputs(4521) <= (layer3_outputs(2283)) and (layer3_outputs(1841));
    layer4_outputs(4522) <= layer3_outputs(796);
    layer4_outputs(4523) <= (layer3_outputs(2713)) and (layer3_outputs(3384));
    layer4_outputs(4524) <= not(layer3_outputs(5091));
    layer4_outputs(4525) <= layer3_outputs(1700);
    layer4_outputs(4526) <= layer3_outputs(4034);
    layer4_outputs(4527) <= not(layer3_outputs(4368));
    layer4_outputs(4528) <= '1';
    layer4_outputs(4529) <= layer3_outputs(2903);
    layer4_outputs(4530) <= (layer3_outputs(3011)) and not (layer3_outputs(1760));
    layer4_outputs(4531) <= not(layer3_outputs(610));
    layer4_outputs(4532) <= not(layer3_outputs(624));
    layer4_outputs(4533) <= not(layer3_outputs(2422)) or (layer3_outputs(2687));
    layer4_outputs(4534) <= not(layer3_outputs(942));
    layer4_outputs(4535) <= not(layer3_outputs(2762)) or (layer3_outputs(2652));
    layer4_outputs(4536) <= not(layer3_outputs(1673));
    layer4_outputs(4537) <= (layer3_outputs(3372)) or (layer3_outputs(2850));
    layer4_outputs(4538) <= not((layer3_outputs(4362)) and (layer3_outputs(2479)));
    layer4_outputs(4539) <= layer3_outputs(2112);
    layer4_outputs(4540) <= (layer3_outputs(5010)) or (layer3_outputs(5092));
    layer4_outputs(4541) <= '0';
    layer4_outputs(4542) <= not(layer3_outputs(2033)) or (layer3_outputs(3539));
    layer4_outputs(4543) <= not(layer3_outputs(2500));
    layer4_outputs(4544) <= layer3_outputs(4842);
    layer4_outputs(4545) <= layer3_outputs(5089);
    layer4_outputs(4546) <= not((layer3_outputs(2267)) xor (layer3_outputs(353)));
    layer4_outputs(4547) <= (layer3_outputs(1448)) and not (layer3_outputs(664));
    layer4_outputs(4548) <= '0';
    layer4_outputs(4549) <= layer3_outputs(3081);
    layer4_outputs(4550) <= not(layer3_outputs(2952)) or (layer3_outputs(76));
    layer4_outputs(4551) <= not(layer3_outputs(2795));
    layer4_outputs(4552) <= '1';
    layer4_outputs(4553) <= not(layer3_outputs(3334)) or (layer3_outputs(3415));
    layer4_outputs(4554) <= not((layer3_outputs(4092)) or (layer3_outputs(2287)));
    layer4_outputs(4555) <= not(layer3_outputs(2828)) or (layer3_outputs(536));
    layer4_outputs(4556) <= layer3_outputs(4454);
    layer4_outputs(4557) <= layer3_outputs(1430);
    layer4_outputs(4558) <= (layer3_outputs(2407)) or (layer3_outputs(2719));
    layer4_outputs(4559) <= (layer3_outputs(2542)) and (layer3_outputs(3039));
    layer4_outputs(4560) <= layer3_outputs(1112);
    layer4_outputs(4561) <= not(layer3_outputs(3326));
    layer4_outputs(4562) <= '0';
    layer4_outputs(4563) <= not((layer3_outputs(4288)) xor (layer3_outputs(2198)));
    layer4_outputs(4564) <= '1';
    layer4_outputs(4565) <= not(layer3_outputs(2060));
    layer4_outputs(4566) <= '0';
    layer4_outputs(4567) <= (layer3_outputs(818)) xor (layer3_outputs(4450));
    layer4_outputs(4568) <= (layer3_outputs(4725)) and not (layer3_outputs(1031));
    layer4_outputs(4569) <= not(layer3_outputs(3125)) or (layer3_outputs(911));
    layer4_outputs(4570) <= not(layer3_outputs(3698)) or (layer3_outputs(3907));
    layer4_outputs(4571) <= '1';
    layer4_outputs(4572) <= not(layer3_outputs(1950));
    layer4_outputs(4573) <= not((layer3_outputs(2081)) or (layer3_outputs(5011)));
    layer4_outputs(4574) <= '0';
    layer4_outputs(4575) <= not((layer3_outputs(4029)) or (layer3_outputs(1948)));
    layer4_outputs(4576) <= '1';
    layer4_outputs(4577) <= layer3_outputs(3215);
    layer4_outputs(4578) <= layer3_outputs(4657);
    layer4_outputs(4579) <= layer3_outputs(866);
    layer4_outputs(4580) <= layer3_outputs(1176);
    layer4_outputs(4581) <= (layer3_outputs(661)) and not (layer3_outputs(328));
    layer4_outputs(4582) <= not((layer3_outputs(754)) and (layer3_outputs(3809)));
    layer4_outputs(4583) <= not(layer3_outputs(3479)) or (layer3_outputs(4245));
    layer4_outputs(4584) <= not(layer3_outputs(2231));
    layer4_outputs(4585) <= '1';
    layer4_outputs(4586) <= layer3_outputs(1293);
    layer4_outputs(4587) <= (layer3_outputs(2093)) and not (layer3_outputs(1160));
    layer4_outputs(4588) <= '0';
    layer4_outputs(4589) <= (layer3_outputs(1888)) or (layer3_outputs(720));
    layer4_outputs(4590) <= not(layer3_outputs(1705));
    layer4_outputs(4591) <= not(layer3_outputs(2055));
    layer4_outputs(4592) <= not(layer3_outputs(24));
    layer4_outputs(4593) <= not((layer3_outputs(1059)) xor (layer3_outputs(2977)));
    layer4_outputs(4594) <= not(layer3_outputs(3873)) or (layer3_outputs(2061));
    layer4_outputs(4595) <= layer3_outputs(105);
    layer4_outputs(4596) <= not((layer3_outputs(5027)) and (layer3_outputs(3458)));
    layer4_outputs(4597) <= (layer3_outputs(1579)) and not (layer3_outputs(837));
    layer4_outputs(4598) <= not((layer3_outputs(2971)) or (layer3_outputs(4241)));
    layer4_outputs(4599) <= not((layer3_outputs(152)) and (layer3_outputs(2951)));
    layer4_outputs(4600) <= not((layer3_outputs(3176)) or (layer3_outputs(5014)));
    layer4_outputs(4601) <= (layer3_outputs(4153)) and (layer3_outputs(4721));
    layer4_outputs(4602) <= not(layer3_outputs(4547));
    layer4_outputs(4603) <= layer3_outputs(3522);
    layer4_outputs(4604) <= not(layer3_outputs(3491));
    layer4_outputs(4605) <= not(layer3_outputs(3642)) or (layer3_outputs(4380));
    layer4_outputs(4606) <= (layer3_outputs(2582)) or (layer3_outputs(5095));
    layer4_outputs(4607) <= (layer3_outputs(2445)) and not (layer3_outputs(3198));
    layer4_outputs(4608) <= not((layer3_outputs(1152)) and (layer3_outputs(4357)));
    layer4_outputs(4609) <= not(layer3_outputs(495));
    layer4_outputs(4610) <= (layer3_outputs(1777)) and not (layer3_outputs(4958));
    layer4_outputs(4611) <= not((layer3_outputs(884)) and (layer3_outputs(2648)));
    layer4_outputs(4612) <= (layer3_outputs(986)) and not (layer3_outputs(7));
    layer4_outputs(4613) <= (layer3_outputs(4187)) and not (layer3_outputs(2618));
    layer4_outputs(4614) <= '1';
    layer4_outputs(4615) <= layer3_outputs(1110);
    layer4_outputs(4616) <= '1';
    layer4_outputs(4617) <= not(layer3_outputs(4066)) or (layer3_outputs(2788));
    layer4_outputs(4618) <= (layer3_outputs(843)) and not (layer3_outputs(1627));
    layer4_outputs(4619) <= '0';
    layer4_outputs(4620) <= layer3_outputs(1324);
    layer4_outputs(4621) <= not((layer3_outputs(3154)) and (layer3_outputs(4743)));
    layer4_outputs(4622) <= not(layer3_outputs(3570)) or (layer3_outputs(3824));
    layer4_outputs(4623) <= not(layer3_outputs(4500));
    layer4_outputs(4624) <= (layer3_outputs(3595)) and (layer3_outputs(3817));
    layer4_outputs(4625) <= not(layer3_outputs(2693));
    layer4_outputs(4626) <= layer3_outputs(2556);
    layer4_outputs(4627) <= not(layer3_outputs(4902));
    layer4_outputs(4628) <= not(layer3_outputs(4834));
    layer4_outputs(4629) <= (layer3_outputs(4417)) and (layer3_outputs(907));
    layer4_outputs(4630) <= not((layer3_outputs(673)) xor (layer3_outputs(4824)));
    layer4_outputs(4631) <= '0';
    layer4_outputs(4632) <= layer3_outputs(2342);
    layer4_outputs(4633) <= (layer3_outputs(2813)) and (layer3_outputs(3968));
    layer4_outputs(4634) <= not(layer3_outputs(2521)) or (layer3_outputs(1016));
    layer4_outputs(4635) <= layer3_outputs(4100);
    layer4_outputs(4636) <= layer3_outputs(1145);
    layer4_outputs(4637) <= not((layer3_outputs(4234)) and (layer3_outputs(4469)));
    layer4_outputs(4638) <= layer3_outputs(598);
    layer4_outputs(4639) <= (layer3_outputs(40)) and not (layer3_outputs(2563));
    layer4_outputs(4640) <= layer3_outputs(3645);
    layer4_outputs(4641) <= not((layer3_outputs(1369)) or (layer3_outputs(4632)));
    layer4_outputs(4642) <= not(layer3_outputs(1302));
    layer4_outputs(4643) <= (layer3_outputs(2978)) and not (layer3_outputs(3540));
    layer4_outputs(4644) <= (layer3_outputs(349)) and not (layer3_outputs(1791));
    layer4_outputs(4645) <= (layer3_outputs(4691)) or (layer3_outputs(3956));
    layer4_outputs(4646) <= not(layer3_outputs(3577));
    layer4_outputs(4647) <= not(layer3_outputs(1825)) or (layer3_outputs(2051));
    layer4_outputs(4648) <= layer3_outputs(1796);
    layer4_outputs(4649) <= not(layer3_outputs(703));
    layer4_outputs(4650) <= '0';
    layer4_outputs(4651) <= layer3_outputs(4246);
    layer4_outputs(4652) <= not((layer3_outputs(3029)) and (layer3_outputs(4057)));
    layer4_outputs(4653) <= layer3_outputs(3275);
    layer4_outputs(4654) <= not(layer3_outputs(1207));
    layer4_outputs(4655) <= not(layer3_outputs(32));
    layer4_outputs(4656) <= layer3_outputs(906);
    layer4_outputs(4657) <= layer3_outputs(2143);
    layer4_outputs(4658) <= (layer3_outputs(2207)) and not (layer3_outputs(1411));
    layer4_outputs(4659) <= layer3_outputs(1095);
    layer4_outputs(4660) <= layer3_outputs(1719);
    layer4_outputs(4661) <= not(layer3_outputs(3828));
    layer4_outputs(4662) <= layer3_outputs(5006);
    layer4_outputs(4663) <= not(layer3_outputs(713)) or (layer3_outputs(3742));
    layer4_outputs(4664) <= not((layer3_outputs(2757)) and (layer3_outputs(3816)));
    layer4_outputs(4665) <= not(layer3_outputs(4757)) or (layer3_outputs(3392));
    layer4_outputs(4666) <= layer3_outputs(3971);
    layer4_outputs(4667) <= not((layer3_outputs(2835)) and (layer3_outputs(3871)));
    layer4_outputs(4668) <= (layer3_outputs(3825)) or (layer3_outputs(3917));
    layer4_outputs(4669) <= not(layer3_outputs(2411));
    layer4_outputs(4670) <= (layer3_outputs(4912)) and not (layer3_outputs(4386));
    layer4_outputs(4671) <= not(layer3_outputs(2650)) or (layer3_outputs(1436));
    layer4_outputs(4672) <= not((layer3_outputs(3836)) xor (layer3_outputs(4449)));
    layer4_outputs(4673) <= not(layer3_outputs(4831));
    layer4_outputs(4674) <= not((layer3_outputs(691)) and (layer3_outputs(1331)));
    layer4_outputs(4675) <= (layer3_outputs(3357)) and not (layer3_outputs(4253));
    layer4_outputs(4676) <= layer3_outputs(5014);
    layer4_outputs(4677) <= (layer3_outputs(2877)) and not (layer3_outputs(3571));
    layer4_outputs(4678) <= not(layer3_outputs(3755)) or (layer3_outputs(2414));
    layer4_outputs(4679) <= layer3_outputs(3676);
    layer4_outputs(4680) <= not(layer3_outputs(2214));
    layer4_outputs(4681) <= (layer3_outputs(3973)) and (layer3_outputs(4261));
    layer4_outputs(4682) <= not(layer3_outputs(2145));
    layer4_outputs(4683) <= layer3_outputs(1632);
    layer4_outputs(4684) <= layer3_outputs(1269);
    layer4_outputs(4685) <= (layer3_outputs(2796)) and not (layer3_outputs(2958));
    layer4_outputs(4686) <= (layer3_outputs(4635)) and (layer3_outputs(4176));
    layer4_outputs(4687) <= '1';
    layer4_outputs(4688) <= layer3_outputs(3015);
    layer4_outputs(4689) <= (layer3_outputs(362)) and not (layer3_outputs(399));
    layer4_outputs(4690) <= layer3_outputs(3276);
    layer4_outputs(4691) <= (layer3_outputs(4041)) or (layer3_outputs(2273));
    layer4_outputs(4692) <= not(layer3_outputs(886));
    layer4_outputs(4693) <= not((layer3_outputs(4339)) xor (layer3_outputs(2514)));
    layer4_outputs(4694) <= not((layer3_outputs(3156)) and (layer3_outputs(4273)));
    layer4_outputs(4695) <= not(layer3_outputs(3949));
    layer4_outputs(4696) <= (layer3_outputs(3695)) and (layer3_outputs(535));
    layer4_outputs(4697) <= (layer3_outputs(41)) or (layer3_outputs(2395));
    layer4_outputs(4698) <= (layer3_outputs(1724)) or (layer3_outputs(2529));
    layer4_outputs(4699) <= layer3_outputs(1162);
    layer4_outputs(4700) <= '0';
    layer4_outputs(4701) <= layer3_outputs(196);
    layer4_outputs(4702) <= not(layer3_outputs(4990));
    layer4_outputs(4703) <= (layer3_outputs(1441)) or (layer3_outputs(3933));
    layer4_outputs(4704) <= (layer3_outputs(3291)) and not (layer3_outputs(1647));
    layer4_outputs(4705) <= not(layer3_outputs(2475));
    layer4_outputs(4706) <= not(layer3_outputs(251));
    layer4_outputs(4707) <= layer3_outputs(2192);
    layer4_outputs(4708) <= not(layer3_outputs(3135));
    layer4_outputs(4709) <= (layer3_outputs(3745)) and not (layer3_outputs(2485));
    layer4_outputs(4710) <= (layer3_outputs(4340)) and not (layer3_outputs(3637));
    layer4_outputs(4711) <= not(layer3_outputs(1398));
    layer4_outputs(4712) <= not((layer3_outputs(1873)) or (layer3_outputs(1355)));
    layer4_outputs(4713) <= not(layer3_outputs(2561));
    layer4_outputs(4714) <= layer3_outputs(4186);
    layer4_outputs(4715) <= not(layer3_outputs(1928));
    layer4_outputs(4716) <= not(layer3_outputs(4258)) or (layer3_outputs(464));
    layer4_outputs(4717) <= not(layer3_outputs(289));
    layer4_outputs(4718) <= not(layer3_outputs(3762));
    layer4_outputs(4719) <= not(layer3_outputs(4547)) or (layer3_outputs(335));
    layer4_outputs(4720) <= (layer3_outputs(2004)) or (layer3_outputs(3890));
    layer4_outputs(4721) <= not(layer3_outputs(3961));
    layer4_outputs(4722) <= '1';
    layer4_outputs(4723) <= (layer3_outputs(2377)) or (layer3_outputs(2096));
    layer4_outputs(4724) <= not(layer3_outputs(298));
    layer4_outputs(4725) <= not(layer3_outputs(3948));
    layer4_outputs(4726) <= (layer3_outputs(4298)) and not (layer3_outputs(3778));
    layer4_outputs(4727) <= (layer3_outputs(4838)) and not (layer3_outputs(746));
    layer4_outputs(4728) <= (layer3_outputs(3768)) and not (layer3_outputs(4839));
    layer4_outputs(4729) <= (layer3_outputs(3084)) xor (layer3_outputs(2679));
    layer4_outputs(4730) <= (layer3_outputs(3294)) and (layer3_outputs(4769));
    layer4_outputs(4731) <= not((layer3_outputs(4197)) and (layer3_outputs(3608)));
    layer4_outputs(4732) <= layer3_outputs(3457);
    layer4_outputs(4733) <= not((layer3_outputs(3768)) or (layer3_outputs(4103)));
    layer4_outputs(4734) <= not((layer3_outputs(3387)) and (layer3_outputs(1766)));
    layer4_outputs(4735) <= not(layer3_outputs(193)) or (layer3_outputs(2509));
    layer4_outputs(4736) <= not((layer3_outputs(2885)) xor (layer3_outputs(951)));
    layer4_outputs(4737) <= (layer3_outputs(3181)) xor (layer3_outputs(1021));
    layer4_outputs(4738) <= layer3_outputs(36);
    layer4_outputs(4739) <= (layer3_outputs(4460)) and not (layer3_outputs(1264));
    layer4_outputs(4740) <= (layer3_outputs(4969)) xor (layer3_outputs(2214));
    layer4_outputs(4741) <= not(layer3_outputs(3297));
    layer4_outputs(4742) <= not((layer3_outputs(4521)) or (layer3_outputs(4699)));
    layer4_outputs(4743) <= not(layer3_outputs(662));
    layer4_outputs(4744) <= layer3_outputs(303);
    layer4_outputs(4745) <= layer3_outputs(263);
    layer4_outputs(4746) <= not((layer3_outputs(863)) or (layer3_outputs(1859)));
    layer4_outputs(4747) <= not(layer3_outputs(3353));
    layer4_outputs(4748) <= (layer3_outputs(805)) and not (layer3_outputs(144));
    layer4_outputs(4749) <= layer3_outputs(3669);
    layer4_outputs(4750) <= not((layer3_outputs(1318)) and (layer3_outputs(1095)));
    layer4_outputs(4751) <= (layer3_outputs(641)) and not (layer3_outputs(1016));
    layer4_outputs(4752) <= (layer3_outputs(2010)) and (layer3_outputs(916));
    layer4_outputs(4753) <= (layer3_outputs(4445)) or (layer3_outputs(4425));
    layer4_outputs(4754) <= '0';
    layer4_outputs(4755) <= (layer3_outputs(326)) xor (layer3_outputs(140));
    layer4_outputs(4756) <= (layer3_outputs(5062)) and not (layer3_outputs(4921));
    layer4_outputs(4757) <= (layer3_outputs(3408)) and not (layer3_outputs(3047));
    layer4_outputs(4758) <= (layer3_outputs(1396)) and not (layer3_outputs(4279));
    layer4_outputs(4759) <= (layer3_outputs(1734)) and not (layer3_outputs(3909));
    layer4_outputs(4760) <= (layer3_outputs(1738)) and not (layer3_outputs(356));
    layer4_outputs(4761) <= layer3_outputs(1864);
    layer4_outputs(4762) <= not(layer3_outputs(4750));
    layer4_outputs(4763) <= not((layer3_outputs(2428)) or (layer3_outputs(2867)));
    layer4_outputs(4764) <= not((layer3_outputs(2443)) or (layer3_outputs(1299)));
    layer4_outputs(4765) <= not((layer3_outputs(5000)) and (layer3_outputs(4459)));
    layer4_outputs(4766) <= layer3_outputs(2481);
    layer4_outputs(4767) <= layer3_outputs(784);
    layer4_outputs(4768) <= not((layer3_outputs(4507)) xor (layer3_outputs(4158)));
    layer4_outputs(4769) <= (layer3_outputs(2544)) and not (layer3_outputs(35));
    layer4_outputs(4770) <= not(layer3_outputs(3589));
    layer4_outputs(4771) <= not(layer3_outputs(3799)) or (layer3_outputs(3921));
    layer4_outputs(4772) <= not(layer3_outputs(3220));
    layer4_outputs(4773) <= not(layer3_outputs(4585));
    layer4_outputs(4774) <= '0';
    layer4_outputs(4775) <= layer3_outputs(1911);
    layer4_outputs(4776) <= layer3_outputs(1273);
    layer4_outputs(4777) <= not(layer3_outputs(2552));
    layer4_outputs(4778) <= layer3_outputs(3909);
    layer4_outputs(4779) <= (layer3_outputs(2206)) and (layer3_outputs(994));
    layer4_outputs(4780) <= layer3_outputs(3578);
    layer4_outputs(4781) <= not(layer3_outputs(741));
    layer4_outputs(4782) <= not(layer3_outputs(1463)) or (layer3_outputs(694));
    layer4_outputs(4783) <= not((layer3_outputs(478)) or (layer3_outputs(456)));
    layer4_outputs(4784) <= layer3_outputs(4824);
    layer4_outputs(4785) <= not(layer3_outputs(3509));
    layer4_outputs(4786) <= layer3_outputs(848);
    layer4_outputs(4787) <= not(layer3_outputs(2762));
    layer4_outputs(4788) <= (layer3_outputs(4925)) and not (layer3_outputs(1392));
    layer4_outputs(4789) <= not(layer3_outputs(2927));
    layer4_outputs(4790) <= (layer3_outputs(289)) and (layer3_outputs(719));
    layer4_outputs(4791) <= not(layer3_outputs(3595));
    layer4_outputs(4792) <= layer3_outputs(2302);
    layer4_outputs(4793) <= not(layer3_outputs(1322));
    layer4_outputs(4794) <= not((layer3_outputs(4044)) xor (layer3_outputs(3831)));
    layer4_outputs(4795) <= '1';
    layer4_outputs(4796) <= (layer3_outputs(129)) and not (layer3_outputs(3120));
    layer4_outputs(4797) <= not((layer3_outputs(88)) and (layer3_outputs(4672)));
    layer4_outputs(4798) <= (layer3_outputs(1779)) or (layer3_outputs(4244));
    layer4_outputs(4799) <= not(layer3_outputs(4978)) or (layer3_outputs(3373));
    layer4_outputs(4800) <= '0';
    layer4_outputs(4801) <= (layer3_outputs(1608)) and not (layer3_outputs(4882));
    layer4_outputs(4802) <= layer3_outputs(4566);
    layer4_outputs(4803) <= not((layer3_outputs(2429)) and (layer3_outputs(49)));
    layer4_outputs(4804) <= not(layer3_outputs(4678)) or (layer3_outputs(4207));
    layer4_outputs(4805) <= layer3_outputs(2933);
    layer4_outputs(4806) <= '0';
    layer4_outputs(4807) <= '0';
    layer4_outputs(4808) <= (layer3_outputs(202)) and not (layer3_outputs(3522));
    layer4_outputs(4809) <= not(layer3_outputs(1615)) or (layer3_outputs(5025));
    layer4_outputs(4810) <= '0';
    layer4_outputs(4811) <= layer3_outputs(1361);
    layer4_outputs(4812) <= layer3_outputs(2737);
    layer4_outputs(4813) <= not(layer3_outputs(225)) or (layer3_outputs(213));
    layer4_outputs(4814) <= '1';
    layer4_outputs(4815) <= layer3_outputs(645);
    layer4_outputs(4816) <= (layer3_outputs(4740)) and (layer3_outputs(365));
    layer4_outputs(4817) <= (layer3_outputs(3179)) and not (layer3_outputs(3274));
    layer4_outputs(4818) <= not(layer3_outputs(1134)) or (layer3_outputs(245));
    layer4_outputs(4819) <= (layer3_outputs(2714)) and not (layer3_outputs(1015));
    layer4_outputs(4820) <= not((layer3_outputs(4083)) and (layer3_outputs(4762)));
    layer4_outputs(4821) <= layer3_outputs(4544);
    layer4_outputs(4822) <= (layer3_outputs(1361)) and not (layer3_outputs(3540));
    layer4_outputs(4823) <= not(layer3_outputs(3656)) or (layer3_outputs(3022));
    layer4_outputs(4824) <= not(layer3_outputs(1408));
    layer4_outputs(4825) <= not((layer3_outputs(1852)) and (layer3_outputs(2712)));
    layer4_outputs(4826) <= not(layer3_outputs(542));
    layer4_outputs(4827) <= layer3_outputs(3630);
    layer4_outputs(4828) <= '0';
    layer4_outputs(4829) <= (layer3_outputs(4680)) and (layer3_outputs(2600));
    layer4_outputs(4830) <= (layer3_outputs(3081)) xor (layer3_outputs(3840));
    layer4_outputs(4831) <= not((layer3_outputs(2464)) and (layer3_outputs(647)));
    layer4_outputs(4832) <= (layer3_outputs(52)) and (layer3_outputs(3697));
    layer4_outputs(4833) <= layer3_outputs(3430);
    layer4_outputs(4834) <= layer3_outputs(5062);
    layer4_outputs(4835) <= not(layer3_outputs(1679)) or (layer3_outputs(3184));
    layer4_outputs(4836) <= (layer3_outputs(525)) and not (layer3_outputs(1287));
    layer4_outputs(4837) <= not(layer3_outputs(856));
    layer4_outputs(4838) <= not((layer3_outputs(1118)) or (layer3_outputs(3110)));
    layer4_outputs(4839) <= not(layer3_outputs(797));
    layer4_outputs(4840) <= '0';
    layer4_outputs(4841) <= not(layer3_outputs(3544)) or (layer3_outputs(2566));
    layer4_outputs(4842) <= not((layer3_outputs(3741)) xor (layer3_outputs(1519)));
    layer4_outputs(4843) <= not((layer3_outputs(4681)) and (layer3_outputs(1933)));
    layer4_outputs(4844) <= layer3_outputs(1675);
    layer4_outputs(4845) <= '0';
    layer4_outputs(4846) <= not(layer3_outputs(459));
    layer4_outputs(4847) <= '0';
    layer4_outputs(4848) <= not(layer3_outputs(4543));
    layer4_outputs(4849) <= not(layer3_outputs(1300)) or (layer3_outputs(3062));
    layer4_outputs(4850) <= layer3_outputs(2230);
    layer4_outputs(4851) <= not(layer3_outputs(131));
    layer4_outputs(4852) <= not(layer3_outputs(2354)) or (layer3_outputs(3774));
    layer4_outputs(4853) <= '1';
    layer4_outputs(4854) <= not(layer3_outputs(3239));
    layer4_outputs(4855) <= (layer3_outputs(2419)) xor (layer3_outputs(4413));
    layer4_outputs(4856) <= not((layer3_outputs(4592)) and (layer3_outputs(2463)));
    layer4_outputs(4857) <= not(layer3_outputs(2355));
    layer4_outputs(4858) <= (layer3_outputs(4479)) and not (layer3_outputs(4354));
    layer4_outputs(4859) <= (layer3_outputs(2187)) and not (layer3_outputs(4162));
    layer4_outputs(4860) <= layer3_outputs(2530);
    layer4_outputs(4861) <= layer3_outputs(1374);
    layer4_outputs(4862) <= not((layer3_outputs(614)) xor (layer3_outputs(5109)));
    layer4_outputs(4863) <= not(layer3_outputs(4704));
    layer4_outputs(4864) <= (layer3_outputs(61)) xor (layer3_outputs(1189));
    layer4_outputs(4865) <= (layer3_outputs(5046)) and not (layer3_outputs(4842));
    layer4_outputs(4866) <= layer3_outputs(1013);
    layer4_outputs(4867) <= not(layer3_outputs(1045));
    layer4_outputs(4868) <= layer3_outputs(1504);
    layer4_outputs(4869) <= layer3_outputs(4625);
    layer4_outputs(4870) <= not((layer3_outputs(3872)) or (layer3_outputs(2459)));
    layer4_outputs(4871) <= not(layer3_outputs(1354));
    layer4_outputs(4872) <= (layer3_outputs(3537)) and not (layer3_outputs(1879));
    layer4_outputs(4873) <= not((layer3_outputs(4838)) and (layer3_outputs(191)));
    layer4_outputs(4874) <= layer3_outputs(1110);
    layer4_outputs(4875) <= layer3_outputs(3926);
    layer4_outputs(4876) <= not((layer3_outputs(3245)) or (layer3_outputs(3453)));
    layer4_outputs(4877) <= (layer3_outputs(2165)) xor (layer3_outputs(1333));
    layer4_outputs(4878) <= not(layer3_outputs(973));
    layer4_outputs(4879) <= not((layer3_outputs(2866)) xor (layer3_outputs(1613)));
    layer4_outputs(4880) <= layer3_outputs(1777);
    layer4_outputs(4881) <= not(layer3_outputs(482));
    layer4_outputs(4882) <= layer3_outputs(4052);
    layer4_outputs(4883) <= not(layer3_outputs(2115));
    layer4_outputs(4884) <= not(layer3_outputs(1161)) or (layer3_outputs(1601));
    layer4_outputs(4885) <= not((layer3_outputs(1228)) xor (layer3_outputs(5016)));
    layer4_outputs(4886) <= layer3_outputs(2095);
    layer4_outputs(4887) <= not((layer3_outputs(1072)) or (layer3_outputs(4107)));
    layer4_outputs(4888) <= '1';
    layer4_outputs(4889) <= layer3_outputs(2715);
    layer4_outputs(4890) <= not(layer3_outputs(2055));
    layer4_outputs(4891) <= (layer3_outputs(899)) and (layer3_outputs(3460));
    layer4_outputs(4892) <= not((layer3_outputs(134)) and (layer3_outputs(4573)));
    layer4_outputs(4893) <= not((layer3_outputs(422)) and (layer3_outputs(1151)));
    layer4_outputs(4894) <= '1';
    layer4_outputs(4895) <= layer3_outputs(943);
    layer4_outputs(4896) <= layer3_outputs(858);
    layer4_outputs(4897) <= layer3_outputs(1470);
    layer4_outputs(4898) <= layer3_outputs(299);
    layer4_outputs(4899) <= not((layer3_outputs(4010)) or (layer3_outputs(2134)));
    layer4_outputs(4900) <= layer3_outputs(5016);
    layer4_outputs(4901) <= (layer3_outputs(1859)) xor (layer3_outputs(3596));
    layer4_outputs(4902) <= not(layer3_outputs(1677));
    layer4_outputs(4903) <= layer3_outputs(1557);
    layer4_outputs(4904) <= (layer3_outputs(4400)) xor (layer3_outputs(4790));
    layer4_outputs(4905) <= layer3_outputs(23);
    layer4_outputs(4906) <= not(layer3_outputs(4759));
    layer4_outputs(4907) <= not(layer3_outputs(3622));
    layer4_outputs(4908) <= (layer3_outputs(3745)) or (layer3_outputs(1172));
    layer4_outputs(4909) <= not(layer3_outputs(3194));
    layer4_outputs(4910) <= (layer3_outputs(3998)) and not (layer3_outputs(1237));
    layer4_outputs(4911) <= not(layer3_outputs(1638));
    layer4_outputs(4912) <= layer3_outputs(3087);
    layer4_outputs(4913) <= not((layer3_outputs(3848)) and (layer3_outputs(1457)));
    layer4_outputs(4914) <= not(layer3_outputs(3562)) or (layer3_outputs(708));
    layer4_outputs(4915) <= '1';
    layer4_outputs(4916) <= layer3_outputs(1474);
    layer4_outputs(4917) <= '1';
    layer4_outputs(4918) <= not(layer3_outputs(4493));
    layer4_outputs(4919) <= (layer3_outputs(2563)) or (layer3_outputs(4151));
    layer4_outputs(4920) <= (layer3_outputs(4026)) or (layer3_outputs(1188));
    layer4_outputs(4921) <= not(layer3_outputs(3802)) or (layer3_outputs(2203));
    layer4_outputs(4922) <= not(layer3_outputs(3221));
    layer4_outputs(4923) <= layer3_outputs(112);
    layer4_outputs(4924) <= not(layer3_outputs(1927));
    layer4_outputs(4925) <= not(layer3_outputs(4215)) or (layer3_outputs(1263));
    layer4_outputs(4926) <= layer3_outputs(514);
    layer4_outputs(4927) <= not(layer3_outputs(989));
    layer4_outputs(4928) <= not(layer3_outputs(1972)) or (layer3_outputs(1835));
    layer4_outputs(4929) <= not(layer3_outputs(3336));
    layer4_outputs(4930) <= not(layer3_outputs(380));
    layer4_outputs(4931) <= layer3_outputs(3527);
    layer4_outputs(4932) <= '1';
    layer4_outputs(4933) <= (layer3_outputs(977)) or (layer3_outputs(4201));
    layer4_outputs(4934) <= not(layer3_outputs(4432)) or (layer3_outputs(1432));
    layer4_outputs(4935) <= not((layer3_outputs(2148)) and (layer3_outputs(571)));
    layer4_outputs(4936) <= layer3_outputs(1481);
    layer4_outputs(4937) <= not(layer3_outputs(1002));
    layer4_outputs(4938) <= layer3_outputs(4321);
    layer4_outputs(4939) <= not(layer3_outputs(2969)) or (layer3_outputs(3565));
    layer4_outputs(4940) <= (layer3_outputs(3986)) xor (layer3_outputs(4030));
    layer4_outputs(4941) <= not(layer3_outputs(4512));
    layer4_outputs(4942) <= (layer3_outputs(3368)) xor (layer3_outputs(3524));
    layer4_outputs(4943) <= (layer3_outputs(3470)) and not (layer3_outputs(16));
    layer4_outputs(4944) <= not(layer3_outputs(2370)) or (layer3_outputs(675));
    layer4_outputs(4945) <= not(layer3_outputs(1998)) or (layer3_outputs(4935));
    layer4_outputs(4946) <= not(layer3_outputs(4465)) or (layer3_outputs(3267));
    layer4_outputs(4947) <= layer3_outputs(2478);
    layer4_outputs(4948) <= not(layer3_outputs(3414));
    layer4_outputs(4949) <= '0';
    layer4_outputs(4950) <= not(layer3_outputs(4608));
    layer4_outputs(4951) <= (layer3_outputs(4466)) and (layer3_outputs(1939));
    layer4_outputs(4952) <= (layer3_outputs(1065)) and (layer3_outputs(4846));
    layer4_outputs(4953) <= not(layer3_outputs(2128));
    layer4_outputs(4954) <= (layer3_outputs(1159)) and not (layer3_outputs(3875));
    layer4_outputs(4955) <= (layer3_outputs(938)) xor (layer3_outputs(4866));
    layer4_outputs(4956) <= '0';
    layer4_outputs(4957) <= layer3_outputs(5031);
    layer4_outputs(4958) <= not(layer3_outputs(2826));
    layer4_outputs(4959) <= (layer3_outputs(1511)) or (layer3_outputs(2684));
    layer4_outputs(4960) <= not((layer3_outputs(3405)) and (layer3_outputs(170)));
    layer4_outputs(4961) <= not(layer3_outputs(3970));
    layer4_outputs(4962) <= layer3_outputs(3959);
    layer4_outputs(4963) <= '1';
    layer4_outputs(4964) <= not(layer3_outputs(4716));
    layer4_outputs(4965) <= not(layer3_outputs(3648)) or (layer3_outputs(259));
    layer4_outputs(4966) <= layer3_outputs(100);
    layer4_outputs(4967) <= (layer3_outputs(1288)) or (layer3_outputs(83));
    layer4_outputs(4968) <= layer3_outputs(3969);
    layer4_outputs(4969) <= (layer3_outputs(4211)) and not (layer3_outputs(3110));
    layer4_outputs(4970) <= layer3_outputs(4938);
    layer4_outputs(4971) <= (layer3_outputs(670)) or (layer3_outputs(3725));
    layer4_outputs(4972) <= not(layer3_outputs(3290));
    layer4_outputs(4973) <= (layer3_outputs(1687)) xor (layer3_outputs(1308));
    layer4_outputs(4974) <= not(layer3_outputs(1493));
    layer4_outputs(4975) <= not(layer3_outputs(1261));
    layer4_outputs(4976) <= not(layer3_outputs(646));
    layer4_outputs(4977) <= layer3_outputs(1836);
    layer4_outputs(4978) <= not(layer3_outputs(2368));
    layer4_outputs(4979) <= layer3_outputs(4520);
    layer4_outputs(4980) <= (layer3_outputs(402)) and not (layer3_outputs(171));
    layer4_outputs(4981) <= layer3_outputs(1937);
    layer4_outputs(4982) <= layer3_outputs(4001);
    layer4_outputs(4983) <= not((layer3_outputs(2029)) or (layer3_outputs(3259)));
    layer4_outputs(4984) <= not((layer3_outputs(2250)) and (layer3_outputs(2260)));
    layer4_outputs(4985) <= layer3_outputs(86);
    layer4_outputs(4986) <= layer3_outputs(4498);
    layer4_outputs(4987) <= (layer3_outputs(3052)) and not (layer3_outputs(1143));
    layer4_outputs(4988) <= (layer3_outputs(1620)) xor (layer3_outputs(4871));
    layer4_outputs(4989) <= not((layer3_outputs(209)) and (layer3_outputs(440)));
    layer4_outputs(4990) <= not((layer3_outputs(4991)) xor (layer3_outputs(4774)));
    layer4_outputs(4991) <= layer3_outputs(1745);
    layer4_outputs(4992) <= not((layer3_outputs(4524)) xor (layer3_outputs(4491)));
    layer4_outputs(4993) <= layer3_outputs(2221);
    layer4_outputs(4994) <= (layer3_outputs(3042)) and (layer3_outputs(1785));
    layer4_outputs(4995) <= not((layer3_outputs(3510)) xor (layer3_outputs(2022)));
    layer4_outputs(4996) <= layer3_outputs(2768);
    layer4_outputs(4997) <= layer3_outputs(4660);
    layer4_outputs(4998) <= layer3_outputs(1991);
    layer4_outputs(4999) <= not((layer3_outputs(143)) xor (layer3_outputs(4646)));
    layer4_outputs(5000) <= (layer3_outputs(3135)) xor (layer3_outputs(173));
    layer4_outputs(5001) <= layer3_outputs(335);
    layer4_outputs(5002) <= '1';
    layer4_outputs(5003) <= (layer3_outputs(480)) xor (layer3_outputs(4972));
    layer4_outputs(5004) <= layer3_outputs(2409);
    layer4_outputs(5005) <= layer3_outputs(740);
    layer4_outputs(5006) <= not((layer3_outputs(3154)) and (layer3_outputs(3728)));
    layer4_outputs(5007) <= layer3_outputs(5111);
    layer4_outputs(5008) <= layer3_outputs(1594);
    layer4_outputs(5009) <= (layer3_outputs(2404)) and (layer3_outputs(2822));
    layer4_outputs(5010) <= (layer3_outputs(1129)) or (layer3_outputs(681));
    layer4_outputs(5011) <= layer3_outputs(3498);
    layer4_outputs(5012) <= layer3_outputs(564);
    layer4_outputs(5013) <= (layer3_outputs(3597)) and not (layer3_outputs(234));
    layer4_outputs(5014) <= not(layer3_outputs(637));
    layer4_outputs(5015) <= not((layer3_outputs(2295)) and (layer3_outputs(4337)));
    layer4_outputs(5016) <= (layer3_outputs(1527)) and not (layer3_outputs(472));
    layer4_outputs(5017) <= not((layer3_outputs(384)) and (layer3_outputs(2927)));
    layer4_outputs(5018) <= layer3_outputs(1106);
    layer4_outputs(5019) <= '0';
    layer4_outputs(5020) <= layer3_outputs(2245);
    layer4_outputs(5021) <= (layer3_outputs(1259)) or (layer3_outputs(4696));
    layer4_outputs(5022) <= not(layer3_outputs(3362));
    layer4_outputs(5023) <= not((layer3_outputs(874)) and (layer3_outputs(412)));
    layer4_outputs(5024) <= (layer3_outputs(2624)) and not (layer3_outputs(490));
    layer4_outputs(5025) <= not(layer3_outputs(4588));
    layer4_outputs(5026) <= layer3_outputs(2494);
    layer4_outputs(5027) <= (layer3_outputs(227)) xor (layer3_outputs(1708));
    layer4_outputs(5028) <= not(layer3_outputs(2356));
    layer4_outputs(5029) <= (layer3_outputs(4043)) and (layer3_outputs(3574));
    layer4_outputs(5030) <= not((layer3_outputs(934)) or (layer3_outputs(1918)));
    layer4_outputs(5031) <= not((layer3_outputs(3957)) or (layer3_outputs(1348)));
    layer4_outputs(5032) <= (layer3_outputs(2633)) xor (layer3_outputs(880));
    layer4_outputs(5033) <= not((layer3_outputs(3641)) and (layer3_outputs(1668)));
    layer4_outputs(5034) <= (layer3_outputs(2122)) and (layer3_outputs(2001));
    layer4_outputs(5035) <= not(layer3_outputs(520));
    layer4_outputs(5036) <= not(layer3_outputs(4602));
    layer4_outputs(5037) <= not(layer3_outputs(558));
    layer4_outputs(5038) <= not(layer3_outputs(4300));
    layer4_outputs(5039) <= (layer3_outputs(4242)) or (layer3_outputs(3378));
    layer4_outputs(5040) <= not(layer3_outputs(4366)) or (layer3_outputs(620));
    layer4_outputs(5041) <= not(layer3_outputs(209));
    layer4_outputs(5042) <= (layer3_outputs(3822)) and (layer3_outputs(4016));
    layer4_outputs(5043) <= not(layer3_outputs(1737));
    layer4_outputs(5044) <= '1';
    layer4_outputs(5045) <= not(layer3_outputs(3177)) or (layer3_outputs(4867));
    layer4_outputs(5046) <= (layer3_outputs(512)) and not (layer3_outputs(2591));
    layer4_outputs(5047) <= not(layer3_outputs(2086));
    layer4_outputs(5048) <= layer3_outputs(5114);
    layer4_outputs(5049) <= '1';
    layer4_outputs(5050) <= (layer3_outputs(378)) and not (layer3_outputs(2965));
    layer4_outputs(5051) <= layer3_outputs(1680);
    layer4_outputs(5052) <= '0';
    layer4_outputs(5053) <= layer3_outputs(2037);
    layer4_outputs(5054) <= not(layer3_outputs(984)) or (layer3_outputs(1886));
    layer4_outputs(5055) <= not(layer3_outputs(5118));
    layer4_outputs(5056) <= not((layer3_outputs(4046)) or (layer3_outputs(2580)));
    layer4_outputs(5057) <= '1';
    layer4_outputs(5058) <= (layer3_outputs(3680)) and (layer3_outputs(1978));
    layer4_outputs(5059) <= '0';
    layer4_outputs(5060) <= not(layer3_outputs(1054));
    layer4_outputs(5061) <= not(layer3_outputs(1771));
    layer4_outputs(5062) <= (layer3_outputs(3309)) and not (layer3_outputs(5101));
    layer4_outputs(5063) <= not((layer3_outputs(3047)) xor (layer3_outputs(4089)));
    layer4_outputs(5064) <= not(layer3_outputs(263));
    layer4_outputs(5065) <= not(layer3_outputs(2520));
    layer4_outputs(5066) <= not(layer3_outputs(3050));
    layer4_outputs(5067) <= layer3_outputs(518);
    layer4_outputs(5068) <= (layer3_outputs(2834)) xor (layer3_outputs(1379));
    layer4_outputs(5069) <= (layer3_outputs(1770)) and not (layer3_outputs(930));
    layer4_outputs(5070) <= not(layer3_outputs(1236)) or (layer3_outputs(2750));
    layer4_outputs(5071) <= '1';
    layer4_outputs(5072) <= not((layer3_outputs(5098)) and (layer3_outputs(904)));
    layer4_outputs(5073) <= layer3_outputs(3756);
    layer4_outputs(5074) <= not((layer3_outputs(3994)) or (layer3_outputs(180)));
    layer4_outputs(5075) <= not(layer3_outputs(4478));
    layer4_outputs(5076) <= layer3_outputs(3962);
    layer4_outputs(5077) <= layer3_outputs(931);
    layer4_outputs(5078) <= not(layer3_outputs(426)) or (layer3_outputs(793));
    layer4_outputs(5079) <= layer3_outputs(421);
    layer4_outputs(5080) <= not(layer3_outputs(3061));
    layer4_outputs(5081) <= not(layer3_outputs(1348));
    layer4_outputs(5082) <= (layer3_outputs(776)) and not (layer3_outputs(3252));
    layer4_outputs(5083) <= layer3_outputs(2146);
    layer4_outputs(5084) <= '1';
    layer4_outputs(5085) <= (layer3_outputs(797)) and (layer3_outputs(2058));
    layer4_outputs(5086) <= not(layer3_outputs(3378)) or (layer3_outputs(315));
    layer4_outputs(5087) <= not(layer3_outputs(1915)) or (layer3_outputs(3145));
    layer4_outputs(5088) <= (layer3_outputs(5005)) and (layer3_outputs(3150));
    layer4_outputs(5089) <= not((layer3_outputs(1447)) xor (layer3_outputs(4229)));
    layer4_outputs(5090) <= not(layer3_outputs(3386)) or (layer3_outputs(452));
    layer4_outputs(5091) <= layer3_outputs(231);
    layer4_outputs(5092) <= '1';
    layer4_outputs(5093) <= layer3_outputs(4515);
    layer4_outputs(5094) <= '1';
    layer4_outputs(5095) <= not(layer3_outputs(4816)) or (layer3_outputs(5096));
    layer4_outputs(5096) <= not(layer3_outputs(5103));
    layer4_outputs(5097) <= (layer3_outputs(4977)) and not (layer3_outputs(4330));
    layer4_outputs(5098) <= (layer3_outputs(1238)) and (layer3_outputs(172));
    layer4_outputs(5099) <= not((layer3_outputs(3260)) and (layer3_outputs(2976)));
    layer4_outputs(5100) <= '1';
    layer4_outputs(5101) <= (layer3_outputs(1218)) and not (layer3_outputs(1691));
    layer4_outputs(5102) <= (layer3_outputs(1327)) and (layer3_outputs(2667));
    layer4_outputs(5103) <= layer3_outputs(1839);
    layer4_outputs(5104) <= layer3_outputs(3147);
    layer4_outputs(5105) <= (layer3_outputs(3908)) and not (layer3_outputs(2972));
    layer4_outputs(5106) <= '0';
    layer4_outputs(5107) <= layer3_outputs(4173);
    layer4_outputs(5108) <= '1';
    layer4_outputs(5109) <= not(layer3_outputs(686)) or (layer3_outputs(413));
    layer4_outputs(5110) <= layer3_outputs(3534);
    layer4_outputs(5111) <= (layer3_outputs(4135)) xor (layer3_outputs(1893));
    layer4_outputs(5112) <= not(layer3_outputs(4440));
    layer4_outputs(5113) <= layer3_outputs(4203);
    layer4_outputs(5114) <= layer3_outputs(4973);
    layer4_outputs(5115) <= not((layer3_outputs(4308)) or (layer3_outputs(3827)));
    layer4_outputs(5116) <= (layer3_outputs(1970)) and not (layer3_outputs(4898));
    layer4_outputs(5117) <= layer3_outputs(247);
    layer4_outputs(5118) <= (layer3_outputs(2429)) and (layer3_outputs(1813));
    layer4_outputs(5119) <= not(layer3_outputs(4546)) or (layer3_outputs(2050));
    layer5_outputs(0) <= layer4_outputs(936);
    layer5_outputs(1) <= (layer4_outputs(515)) and not (layer4_outputs(2675));
    layer5_outputs(2) <= layer4_outputs(3808);
    layer5_outputs(3) <= not(layer4_outputs(4210)) or (layer4_outputs(3570));
    layer5_outputs(4) <= (layer4_outputs(892)) and (layer4_outputs(2766));
    layer5_outputs(5) <= not(layer4_outputs(475));
    layer5_outputs(6) <= (layer4_outputs(1625)) and (layer4_outputs(4758));
    layer5_outputs(7) <= not((layer4_outputs(2465)) and (layer4_outputs(2548)));
    layer5_outputs(8) <= layer4_outputs(702);
    layer5_outputs(9) <= (layer4_outputs(2482)) or (layer4_outputs(726));
    layer5_outputs(10) <= layer4_outputs(1341);
    layer5_outputs(11) <= not(layer4_outputs(2678)) or (layer4_outputs(3066));
    layer5_outputs(12) <= layer4_outputs(2281);
    layer5_outputs(13) <= not(layer4_outputs(1129));
    layer5_outputs(14) <= not(layer4_outputs(2483));
    layer5_outputs(15) <= (layer4_outputs(904)) and not (layer4_outputs(3260));
    layer5_outputs(16) <= not(layer4_outputs(1581));
    layer5_outputs(17) <= not((layer4_outputs(4051)) or (layer4_outputs(3726)));
    layer5_outputs(18) <= not((layer4_outputs(2044)) and (layer4_outputs(2600)));
    layer5_outputs(19) <= '1';
    layer5_outputs(20) <= not(layer4_outputs(2266)) or (layer4_outputs(3382));
    layer5_outputs(21) <= not((layer4_outputs(67)) xor (layer4_outputs(3385)));
    layer5_outputs(22) <= not(layer4_outputs(3587));
    layer5_outputs(23) <= '0';
    layer5_outputs(24) <= (layer4_outputs(4332)) and not (layer4_outputs(1660));
    layer5_outputs(25) <= layer4_outputs(3730);
    layer5_outputs(26) <= not(layer4_outputs(1399));
    layer5_outputs(27) <= layer4_outputs(2648);
    layer5_outputs(28) <= '1';
    layer5_outputs(29) <= layer4_outputs(3581);
    layer5_outputs(30) <= not((layer4_outputs(725)) or (layer4_outputs(3472)));
    layer5_outputs(31) <= (layer4_outputs(2225)) and (layer4_outputs(3950));
    layer5_outputs(32) <= layer4_outputs(4193);
    layer5_outputs(33) <= layer4_outputs(440);
    layer5_outputs(34) <= not(layer4_outputs(3716));
    layer5_outputs(35) <= (layer4_outputs(1924)) and (layer4_outputs(875));
    layer5_outputs(36) <= (layer4_outputs(2954)) and (layer4_outputs(4828));
    layer5_outputs(37) <= not(layer4_outputs(1688));
    layer5_outputs(38) <= not(layer4_outputs(1855));
    layer5_outputs(39) <= (layer4_outputs(466)) xor (layer4_outputs(1787));
    layer5_outputs(40) <= not((layer4_outputs(894)) xor (layer4_outputs(4760)));
    layer5_outputs(41) <= not(layer4_outputs(4156)) or (layer4_outputs(2723));
    layer5_outputs(42) <= (layer4_outputs(535)) or (layer4_outputs(2538));
    layer5_outputs(43) <= (layer4_outputs(1527)) and not (layer4_outputs(4709));
    layer5_outputs(44) <= layer4_outputs(4061);
    layer5_outputs(45) <= not(layer4_outputs(634)) or (layer4_outputs(2478));
    layer5_outputs(46) <= (layer4_outputs(701)) and not (layer4_outputs(1283));
    layer5_outputs(47) <= not(layer4_outputs(4021));
    layer5_outputs(48) <= not(layer4_outputs(3026)) or (layer4_outputs(3992));
    layer5_outputs(49) <= (layer4_outputs(3666)) or (layer4_outputs(4085));
    layer5_outputs(50) <= not(layer4_outputs(1915));
    layer5_outputs(51) <= (layer4_outputs(1613)) and not (layer4_outputs(4869));
    layer5_outputs(52) <= '1';
    layer5_outputs(53) <= (layer4_outputs(64)) and not (layer4_outputs(4263));
    layer5_outputs(54) <= layer4_outputs(898);
    layer5_outputs(55) <= (layer4_outputs(1343)) and not (layer4_outputs(914));
    layer5_outputs(56) <= layer4_outputs(2051);
    layer5_outputs(57) <= not(layer4_outputs(4250));
    layer5_outputs(58) <= layer4_outputs(1417);
    layer5_outputs(59) <= not(layer4_outputs(2708));
    layer5_outputs(60) <= (layer4_outputs(1664)) and (layer4_outputs(1905));
    layer5_outputs(61) <= layer4_outputs(4538);
    layer5_outputs(62) <= (layer4_outputs(1546)) or (layer4_outputs(4087));
    layer5_outputs(63) <= '0';
    layer5_outputs(64) <= not(layer4_outputs(841));
    layer5_outputs(65) <= layer4_outputs(3813);
    layer5_outputs(66) <= layer4_outputs(1805);
    layer5_outputs(67) <= not(layer4_outputs(2356)) or (layer4_outputs(4517));
    layer5_outputs(68) <= layer4_outputs(2590);
    layer5_outputs(69) <= layer4_outputs(4786);
    layer5_outputs(70) <= not((layer4_outputs(1505)) xor (layer4_outputs(1608)));
    layer5_outputs(71) <= not(layer4_outputs(3363)) or (layer4_outputs(4677));
    layer5_outputs(72) <= layer4_outputs(3913);
    layer5_outputs(73) <= '0';
    layer5_outputs(74) <= not(layer4_outputs(1031));
    layer5_outputs(75) <= not((layer4_outputs(2584)) and (layer4_outputs(4511)));
    layer5_outputs(76) <= layer4_outputs(460);
    layer5_outputs(77) <= layer4_outputs(2590);
    layer5_outputs(78) <= layer4_outputs(601);
    layer5_outputs(79) <= layer4_outputs(3609);
    layer5_outputs(80) <= layer4_outputs(3097);
    layer5_outputs(81) <= not((layer4_outputs(1679)) xor (layer4_outputs(1703)));
    layer5_outputs(82) <= not(layer4_outputs(3433)) or (layer4_outputs(305));
    layer5_outputs(83) <= layer4_outputs(1323);
    layer5_outputs(84) <= (layer4_outputs(2502)) and not (layer4_outputs(82));
    layer5_outputs(85) <= not(layer4_outputs(4733)) or (layer4_outputs(4925));
    layer5_outputs(86) <= not(layer4_outputs(2955));
    layer5_outputs(87) <= not((layer4_outputs(230)) xor (layer4_outputs(3086)));
    layer5_outputs(88) <= layer4_outputs(1334);
    layer5_outputs(89) <= not(layer4_outputs(2736));
    layer5_outputs(90) <= layer4_outputs(4511);
    layer5_outputs(91) <= '1';
    layer5_outputs(92) <= not((layer4_outputs(2373)) and (layer4_outputs(4016)));
    layer5_outputs(93) <= layer4_outputs(4680);
    layer5_outputs(94) <= layer4_outputs(268);
    layer5_outputs(95) <= not(layer4_outputs(3848)) or (layer4_outputs(4751));
    layer5_outputs(96) <= not(layer4_outputs(4182));
    layer5_outputs(97) <= (layer4_outputs(2608)) and not (layer4_outputs(3478));
    layer5_outputs(98) <= (layer4_outputs(3394)) xor (layer4_outputs(1438));
    layer5_outputs(99) <= '1';
    layer5_outputs(100) <= not(layer4_outputs(4931));
    layer5_outputs(101) <= not(layer4_outputs(2292));
    layer5_outputs(102) <= (layer4_outputs(3910)) and not (layer4_outputs(497));
    layer5_outputs(103) <= not(layer4_outputs(1960));
    layer5_outputs(104) <= '1';
    layer5_outputs(105) <= not(layer4_outputs(1912));
    layer5_outputs(106) <= layer4_outputs(3621);
    layer5_outputs(107) <= (layer4_outputs(5018)) and not (layer4_outputs(2637));
    layer5_outputs(108) <= (layer4_outputs(1124)) and not (layer4_outputs(2900));
    layer5_outputs(109) <= '0';
    layer5_outputs(110) <= not(layer4_outputs(4744));
    layer5_outputs(111) <= not(layer4_outputs(2761));
    layer5_outputs(112) <= (layer4_outputs(3255)) and not (layer4_outputs(4827));
    layer5_outputs(113) <= layer4_outputs(1906);
    layer5_outputs(114) <= not((layer4_outputs(26)) or (layer4_outputs(2109)));
    layer5_outputs(115) <= not((layer4_outputs(2814)) xor (layer4_outputs(917)));
    layer5_outputs(116) <= not(layer4_outputs(2664)) or (layer4_outputs(4142));
    layer5_outputs(117) <= '1';
    layer5_outputs(118) <= not(layer4_outputs(3638)) or (layer4_outputs(5079));
    layer5_outputs(119) <= (layer4_outputs(4798)) and (layer4_outputs(4953));
    layer5_outputs(120) <= '1';
    layer5_outputs(121) <= not(layer4_outputs(1660)) or (layer4_outputs(651));
    layer5_outputs(122) <= layer4_outputs(3805);
    layer5_outputs(123) <= layer4_outputs(4189);
    layer5_outputs(124) <= not(layer4_outputs(1348));
    layer5_outputs(125) <= layer4_outputs(1330);
    layer5_outputs(126) <= layer4_outputs(497);
    layer5_outputs(127) <= layer4_outputs(3601);
    layer5_outputs(128) <= layer4_outputs(2421);
    layer5_outputs(129) <= '1';
    layer5_outputs(130) <= layer4_outputs(2634);
    layer5_outputs(131) <= layer4_outputs(5092);
    layer5_outputs(132) <= layer4_outputs(406);
    layer5_outputs(133) <= not(layer4_outputs(2521));
    layer5_outputs(134) <= (layer4_outputs(4105)) xor (layer4_outputs(4915));
    layer5_outputs(135) <= not((layer4_outputs(1270)) and (layer4_outputs(2930)));
    layer5_outputs(136) <= not((layer4_outputs(3539)) or (layer4_outputs(2547)));
    layer5_outputs(137) <= layer4_outputs(2130);
    layer5_outputs(138) <= not(layer4_outputs(2696)) or (layer4_outputs(111));
    layer5_outputs(139) <= not(layer4_outputs(4993));
    layer5_outputs(140) <= layer4_outputs(4442);
    layer5_outputs(141) <= '0';
    layer5_outputs(142) <= not(layer4_outputs(3275));
    layer5_outputs(143) <= layer4_outputs(5101);
    layer5_outputs(144) <= layer4_outputs(3765);
    layer5_outputs(145) <= (layer4_outputs(180)) and not (layer4_outputs(1508));
    layer5_outputs(146) <= layer4_outputs(1040);
    layer5_outputs(147) <= layer4_outputs(4559);
    layer5_outputs(148) <= (layer4_outputs(3806)) and not (layer4_outputs(4912));
    layer5_outputs(149) <= layer4_outputs(4472);
    layer5_outputs(150) <= (layer4_outputs(860)) and not (layer4_outputs(674));
    layer5_outputs(151) <= layer4_outputs(206);
    layer5_outputs(152) <= (layer4_outputs(1201)) and not (layer4_outputs(1684));
    layer5_outputs(153) <= not((layer4_outputs(1928)) and (layer4_outputs(3122)));
    layer5_outputs(154) <= not(layer4_outputs(4389)) or (layer4_outputs(2802));
    layer5_outputs(155) <= not(layer4_outputs(4709));
    layer5_outputs(156) <= not(layer4_outputs(299));
    layer5_outputs(157) <= not(layer4_outputs(3951));
    layer5_outputs(158) <= not((layer4_outputs(3057)) or (layer4_outputs(146)));
    layer5_outputs(159) <= (layer4_outputs(1043)) xor (layer4_outputs(5005));
    layer5_outputs(160) <= layer4_outputs(1759);
    layer5_outputs(161) <= not((layer4_outputs(3417)) and (layer4_outputs(1883)));
    layer5_outputs(162) <= not((layer4_outputs(299)) or (layer4_outputs(2731)));
    layer5_outputs(163) <= not(layer4_outputs(3172));
    layer5_outputs(164) <= not((layer4_outputs(1372)) xor (layer4_outputs(4636)));
    layer5_outputs(165) <= not((layer4_outputs(3631)) or (layer4_outputs(3756)));
    layer5_outputs(166) <= '0';
    layer5_outputs(167) <= not(layer4_outputs(4179));
    layer5_outputs(168) <= not(layer4_outputs(2519));
    layer5_outputs(169) <= (layer4_outputs(665)) and not (layer4_outputs(1333));
    layer5_outputs(170) <= '1';
    layer5_outputs(171) <= (layer4_outputs(1178)) and not (layer4_outputs(3045));
    layer5_outputs(172) <= layer4_outputs(4330);
    layer5_outputs(173) <= layer4_outputs(119);
    layer5_outputs(174) <= '0';
    layer5_outputs(175) <= layer4_outputs(4417);
    layer5_outputs(176) <= not(layer4_outputs(1036)) or (layer4_outputs(1750));
    layer5_outputs(177) <= (layer4_outputs(1516)) xor (layer4_outputs(2007));
    layer5_outputs(178) <= not((layer4_outputs(1319)) xor (layer4_outputs(3452)));
    layer5_outputs(179) <= not(layer4_outputs(777));
    layer5_outputs(180) <= not(layer4_outputs(1433)) or (layer4_outputs(4069));
    layer5_outputs(181) <= layer4_outputs(809);
    layer5_outputs(182) <= not(layer4_outputs(5035));
    layer5_outputs(183) <= layer4_outputs(3653);
    layer5_outputs(184) <= not(layer4_outputs(3554)) or (layer4_outputs(4186));
    layer5_outputs(185) <= layer4_outputs(2013);
    layer5_outputs(186) <= not(layer4_outputs(1696)) or (layer4_outputs(2964));
    layer5_outputs(187) <= not(layer4_outputs(3102)) or (layer4_outputs(3049));
    layer5_outputs(188) <= '1';
    layer5_outputs(189) <= not(layer4_outputs(909));
    layer5_outputs(190) <= layer4_outputs(4784);
    layer5_outputs(191) <= not(layer4_outputs(181));
    layer5_outputs(192) <= not(layer4_outputs(1102));
    layer5_outputs(193) <= '1';
    layer5_outputs(194) <= layer4_outputs(2125);
    layer5_outputs(195) <= not((layer4_outputs(4544)) xor (layer4_outputs(1111)));
    layer5_outputs(196) <= (layer4_outputs(4452)) xor (layer4_outputs(2238));
    layer5_outputs(197) <= not(layer4_outputs(3823)) or (layer4_outputs(4886));
    layer5_outputs(198) <= not((layer4_outputs(4265)) xor (layer4_outputs(189)));
    layer5_outputs(199) <= layer4_outputs(2755);
    layer5_outputs(200) <= layer4_outputs(387);
    layer5_outputs(201) <= layer4_outputs(28);
    layer5_outputs(202) <= not((layer4_outputs(3032)) xor (layer4_outputs(3778)));
    layer5_outputs(203) <= not(layer4_outputs(1314));
    layer5_outputs(204) <= not((layer4_outputs(1354)) xor (layer4_outputs(3127)));
    layer5_outputs(205) <= layer4_outputs(2090);
    layer5_outputs(206) <= not(layer4_outputs(366));
    layer5_outputs(207) <= not(layer4_outputs(4382));
    layer5_outputs(208) <= (layer4_outputs(626)) xor (layer4_outputs(4693));
    layer5_outputs(209) <= (layer4_outputs(4577)) and not (layer4_outputs(3317));
    layer5_outputs(210) <= not(layer4_outputs(2710));
    layer5_outputs(211) <= not(layer4_outputs(2512));
    layer5_outputs(212) <= (layer4_outputs(4262)) or (layer4_outputs(2778));
    layer5_outputs(213) <= layer4_outputs(1030);
    layer5_outputs(214) <= not((layer4_outputs(322)) or (layer4_outputs(3924)));
    layer5_outputs(215) <= layer4_outputs(2576);
    layer5_outputs(216) <= not(layer4_outputs(1783)) or (layer4_outputs(4445));
    layer5_outputs(217) <= not(layer4_outputs(4152)) or (layer4_outputs(1072));
    layer5_outputs(218) <= (layer4_outputs(776)) or (layer4_outputs(1901));
    layer5_outputs(219) <= not(layer4_outputs(2397));
    layer5_outputs(220) <= not(layer4_outputs(5081));
    layer5_outputs(221) <= '1';
    layer5_outputs(222) <= not(layer4_outputs(3179));
    layer5_outputs(223) <= not((layer4_outputs(4554)) or (layer4_outputs(3379)));
    layer5_outputs(224) <= layer4_outputs(463);
    layer5_outputs(225) <= not(layer4_outputs(3412)) or (layer4_outputs(30));
    layer5_outputs(226) <= (layer4_outputs(5086)) and not (layer4_outputs(4856));
    layer5_outputs(227) <= layer4_outputs(7);
    layer5_outputs(228) <= not(layer4_outputs(2970));
    layer5_outputs(229) <= not(layer4_outputs(2755));
    layer5_outputs(230) <= (layer4_outputs(2411)) xor (layer4_outputs(5082));
    layer5_outputs(231) <= not(layer4_outputs(2038));
    layer5_outputs(232) <= '0';
    layer5_outputs(233) <= (layer4_outputs(5015)) or (layer4_outputs(5034));
    layer5_outputs(234) <= layer4_outputs(1690);
    layer5_outputs(235) <= not((layer4_outputs(4407)) or (layer4_outputs(4154)));
    layer5_outputs(236) <= layer4_outputs(3935);
    layer5_outputs(237) <= not(layer4_outputs(3658));
    layer5_outputs(238) <= not((layer4_outputs(2303)) or (layer4_outputs(2856)));
    layer5_outputs(239) <= not(layer4_outputs(2151));
    layer5_outputs(240) <= (layer4_outputs(632)) and not (layer4_outputs(3540));
    layer5_outputs(241) <= not(layer4_outputs(694));
    layer5_outputs(242) <= (layer4_outputs(3066)) and not (layer4_outputs(2460));
    layer5_outputs(243) <= layer4_outputs(5036);
    layer5_outputs(244) <= (layer4_outputs(4405)) and (layer4_outputs(203));
    layer5_outputs(245) <= not(layer4_outputs(3503));
    layer5_outputs(246) <= layer4_outputs(2772);
    layer5_outputs(247) <= (layer4_outputs(2180)) xor (layer4_outputs(3635));
    layer5_outputs(248) <= layer4_outputs(2818);
    layer5_outputs(249) <= layer4_outputs(2519);
    layer5_outputs(250) <= not(layer4_outputs(3850));
    layer5_outputs(251) <= (layer4_outputs(254)) and not (layer4_outputs(4801));
    layer5_outputs(252) <= '0';
    layer5_outputs(253) <= layer4_outputs(2922);
    layer5_outputs(254) <= '0';
    layer5_outputs(255) <= not((layer4_outputs(2442)) xor (layer4_outputs(3210)));
    layer5_outputs(256) <= not(layer4_outputs(212));
    layer5_outputs(257) <= not(layer4_outputs(2696));
    layer5_outputs(258) <= not((layer4_outputs(1852)) or (layer4_outputs(329)));
    layer5_outputs(259) <= (layer4_outputs(3604)) xor (layer4_outputs(164));
    layer5_outputs(260) <= (layer4_outputs(4656)) and not (layer4_outputs(4018));
    layer5_outputs(261) <= not((layer4_outputs(1060)) or (layer4_outputs(4467)));
    layer5_outputs(262) <= layer4_outputs(4602);
    layer5_outputs(263) <= not(layer4_outputs(3541));
    layer5_outputs(264) <= layer4_outputs(1864);
    layer5_outputs(265) <= not(layer4_outputs(1275));
    layer5_outputs(266) <= layer4_outputs(1057);
    layer5_outputs(267) <= not((layer4_outputs(3900)) xor (layer4_outputs(3413)));
    layer5_outputs(268) <= not((layer4_outputs(757)) and (layer4_outputs(944)));
    layer5_outputs(269) <= not((layer4_outputs(5041)) and (layer4_outputs(2641)));
    layer5_outputs(270) <= not((layer4_outputs(756)) xor (layer4_outputs(4804)));
    layer5_outputs(271) <= '1';
    layer5_outputs(272) <= layer4_outputs(2314);
    layer5_outputs(273) <= layer4_outputs(3386);
    layer5_outputs(274) <= not(layer4_outputs(2882));
    layer5_outputs(275) <= (layer4_outputs(3111)) or (layer4_outputs(1995));
    layer5_outputs(276) <= layer4_outputs(3869);
    layer5_outputs(277) <= '1';
    layer5_outputs(278) <= not((layer4_outputs(628)) or (layer4_outputs(4582)));
    layer5_outputs(279) <= not(layer4_outputs(3335)) or (layer4_outputs(97));
    layer5_outputs(280) <= (layer4_outputs(529)) and not (layer4_outputs(3218));
    layer5_outputs(281) <= not(layer4_outputs(2852));
    layer5_outputs(282) <= (layer4_outputs(2125)) and (layer4_outputs(59));
    layer5_outputs(283) <= not(layer4_outputs(1168));
    layer5_outputs(284) <= (layer4_outputs(3600)) xor (layer4_outputs(87));
    layer5_outputs(285) <= layer4_outputs(1171);
    layer5_outputs(286) <= not(layer4_outputs(2355));
    layer5_outputs(287) <= not(layer4_outputs(2263));
    layer5_outputs(288) <= not(layer4_outputs(2643));
    layer5_outputs(289) <= not(layer4_outputs(3355)) or (layer4_outputs(4892));
    layer5_outputs(290) <= (layer4_outputs(4779)) and (layer4_outputs(3036));
    layer5_outputs(291) <= not(layer4_outputs(3483)) or (layer4_outputs(479));
    layer5_outputs(292) <= not((layer4_outputs(1422)) xor (layer4_outputs(4845)));
    layer5_outputs(293) <= not(layer4_outputs(783));
    layer5_outputs(294) <= not((layer4_outputs(4508)) and (layer4_outputs(3454)));
    layer5_outputs(295) <= (layer4_outputs(87)) and (layer4_outputs(3243));
    layer5_outputs(296) <= not(layer4_outputs(2625));
    layer5_outputs(297) <= layer4_outputs(2235);
    layer5_outputs(298) <= not(layer4_outputs(3022)) or (layer4_outputs(1823));
    layer5_outputs(299) <= layer4_outputs(2172);
    layer5_outputs(300) <= not(layer4_outputs(2397));
    layer5_outputs(301) <= not(layer4_outputs(1035));
    layer5_outputs(302) <= (layer4_outputs(904)) or (layer4_outputs(2249));
    layer5_outputs(303) <= (layer4_outputs(2295)) or (layer4_outputs(2634));
    layer5_outputs(304) <= not(layer4_outputs(3050));
    layer5_outputs(305) <= not(layer4_outputs(1521));
    layer5_outputs(306) <= layer4_outputs(81);
    layer5_outputs(307) <= not((layer4_outputs(3834)) and (layer4_outputs(469)));
    layer5_outputs(308) <= (layer4_outputs(2200)) and (layer4_outputs(3740));
    layer5_outputs(309) <= layer4_outputs(2112);
    layer5_outputs(310) <= not(layer4_outputs(2351));
    layer5_outputs(311) <= (layer4_outputs(2429)) or (layer4_outputs(1864));
    layer5_outputs(312) <= layer4_outputs(580);
    layer5_outputs(313) <= (layer4_outputs(2722)) and not (layer4_outputs(3221));
    layer5_outputs(314) <= (layer4_outputs(1409)) xor (layer4_outputs(2121));
    layer5_outputs(315) <= not((layer4_outputs(3269)) xor (layer4_outputs(2047)));
    layer5_outputs(316) <= not(layer4_outputs(4104));
    layer5_outputs(317) <= not((layer4_outputs(505)) xor (layer4_outputs(1618)));
    layer5_outputs(318) <= not(layer4_outputs(1205));
    layer5_outputs(319) <= (layer4_outputs(444)) and not (layer4_outputs(4147));
    layer5_outputs(320) <= not(layer4_outputs(2223)) or (layer4_outputs(2775));
    layer5_outputs(321) <= not(layer4_outputs(4881));
    layer5_outputs(322) <= layer4_outputs(5069);
    layer5_outputs(323) <= (layer4_outputs(5059)) and not (layer4_outputs(1385));
    layer5_outputs(324) <= not(layer4_outputs(3733));
    layer5_outputs(325) <= layer4_outputs(1553);
    layer5_outputs(326) <= not(layer4_outputs(2106)) or (layer4_outputs(1134));
    layer5_outputs(327) <= (layer4_outputs(4586)) or (layer4_outputs(4838));
    layer5_outputs(328) <= not(layer4_outputs(1315)) or (layer4_outputs(1609));
    layer5_outputs(329) <= (layer4_outputs(3392)) or (layer4_outputs(2180));
    layer5_outputs(330) <= layer4_outputs(4878);
    layer5_outputs(331) <= not(layer4_outputs(4572));
    layer5_outputs(332) <= layer4_outputs(4894);
    layer5_outputs(333) <= not(layer4_outputs(3095));
    layer5_outputs(334) <= layer4_outputs(4403);
    layer5_outputs(335) <= layer4_outputs(4321);
    layer5_outputs(336) <= not((layer4_outputs(480)) or (layer4_outputs(3103)));
    layer5_outputs(337) <= layer4_outputs(396);
    layer5_outputs(338) <= layer4_outputs(2481);
    layer5_outputs(339) <= layer4_outputs(4991);
    layer5_outputs(340) <= not(layer4_outputs(2942));
    layer5_outputs(341) <= layer4_outputs(3093);
    layer5_outputs(342) <= not(layer4_outputs(4413));
    layer5_outputs(343) <= not((layer4_outputs(3632)) xor (layer4_outputs(4805)));
    layer5_outputs(344) <= not(layer4_outputs(1440));
    layer5_outputs(345) <= not(layer4_outputs(4366));
    layer5_outputs(346) <= not(layer4_outputs(3707)) or (layer4_outputs(4776));
    layer5_outputs(347) <= layer4_outputs(2596);
    layer5_outputs(348) <= layer4_outputs(3595);
    layer5_outputs(349) <= not((layer4_outputs(4350)) or (layer4_outputs(2633)));
    layer5_outputs(350) <= layer4_outputs(1456);
    layer5_outputs(351) <= not((layer4_outputs(2692)) and (layer4_outputs(3762)));
    layer5_outputs(352) <= (layer4_outputs(525)) and (layer4_outputs(2728));
    layer5_outputs(353) <= layer4_outputs(1562);
    layer5_outputs(354) <= layer4_outputs(1440);
    layer5_outputs(355) <= layer4_outputs(5080);
    layer5_outputs(356) <= layer4_outputs(1261);
    layer5_outputs(357) <= not(layer4_outputs(2201));
    layer5_outputs(358) <= (layer4_outputs(2484)) and not (layer4_outputs(185));
    layer5_outputs(359) <= '1';
    layer5_outputs(360) <= layer4_outputs(400);
    layer5_outputs(361) <= '1';
    layer5_outputs(362) <= (layer4_outputs(1750)) and not (layer4_outputs(515));
    layer5_outputs(363) <= not(layer4_outputs(1434));
    layer5_outputs(364) <= layer4_outputs(2688);
    layer5_outputs(365) <= not(layer4_outputs(3915));
    layer5_outputs(366) <= not(layer4_outputs(4059)) or (layer4_outputs(4980));
    layer5_outputs(367) <= (layer4_outputs(2178)) and (layer4_outputs(1418));
    layer5_outputs(368) <= layer4_outputs(1872);
    layer5_outputs(369) <= not(layer4_outputs(2056));
    layer5_outputs(370) <= not(layer4_outputs(4090));
    layer5_outputs(371) <= layer4_outputs(1797);
    layer5_outputs(372) <= layer4_outputs(2510);
    layer5_outputs(373) <= (layer4_outputs(2298)) or (layer4_outputs(1322));
    layer5_outputs(374) <= (layer4_outputs(3772)) or (layer4_outputs(4242));
    layer5_outputs(375) <= not(layer4_outputs(2443));
    layer5_outputs(376) <= '0';
    layer5_outputs(377) <= layer4_outputs(2800);
    layer5_outputs(378) <= layer4_outputs(527);
    layer5_outputs(379) <= (layer4_outputs(3129)) and (layer4_outputs(844));
    layer5_outputs(380) <= not((layer4_outputs(3547)) xor (layer4_outputs(390)));
    layer5_outputs(381) <= layer4_outputs(2707);
    layer5_outputs(382) <= layer4_outputs(3097);
    layer5_outputs(383) <= not(layer4_outputs(3493));
    layer5_outputs(384) <= layer4_outputs(1251);
    layer5_outputs(385) <= not(layer4_outputs(2387));
    layer5_outputs(386) <= not(layer4_outputs(1028));
    layer5_outputs(387) <= layer4_outputs(180);
    layer5_outputs(388) <= layer4_outputs(292);
    layer5_outputs(389) <= (layer4_outputs(1365)) xor (layer4_outputs(3185));
    layer5_outputs(390) <= not(layer4_outputs(89));
    layer5_outputs(391) <= (layer4_outputs(4958)) and (layer4_outputs(6));
    layer5_outputs(392) <= not(layer4_outputs(3474));
    layer5_outputs(393) <= not(layer4_outputs(4473));
    layer5_outputs(394) <= (layer4_outputs(2372)) and (layer4_outputs(2360));
    layer5_outputs(395) <= not(layer4_outputs(1970));
    layer5_outputs(396) <= not(layer4_outputs(2267));
    layer5_outputs(397) <= layer4_outputs(5115);
    layer5_outputs(398) <= layer4_outputs(3464);
    layer5_outputs(399) <= not(layer4_outputs(773));
    layer5_outputs(400) <= not((layer4_outputs(3656)) or (layer4_outputs(2413)));
    layer5_outputs(401) <= not(layer4_outputs(2718));
    layer5_outputs(402) <= layer4_outputs(2291);
    layer5_outputs(403) <= layer4_outputs(3415);
    layer5_outputs(404) <= not((layer4_outputs(1889)) and (layer4_outputs(3256)));
    layer5_outputs(405) <= not(layer4_outputs(116));
    layer5_outputs(406) <= not((layer4_outputs(1143)) xor (layer4_outputs(2838)));
    layer5_outputs(407) <= not((layer4_outputs(4795)) and (layer4_outputs(4318)));
    layer5_outputs(408) <= not((layer4_outputs(3239)) xor (layer4_outputs(4479)));
    layer5_outputs(409) <= not(layer4_outputs(218));
    layer5_outputs(410) <= layer4_outputs(1467);
    layer5_outputs(411) <= not(layer4_outputs(3580)) or (layer4_outputs(886));
    layer5_outputs(412) <= layer4_outputs(5099);
    layer5_outputs(413) <= not(layer4_outputs(871));
    layer5_outputs(414) <= not(layer4_outputs(3072));
    layer5_outputs(415) <= not(layer4_outputs(1977));
    layer5_outputs(416) <= not((layer4_outputs(842)) xor (layer4_outputs(2323)));
    layer5_outputs(417) <= layer4_outputs(260);
    layer5_outputs(418) <= layer4_outputs(2795);
    layer5_outputs(419) <= (layer4_outputs(2095)) or (layer4_outputs(1555));
    layer5_outputs(420) <= (layer4_outputs(1979)) or (layer4_outputs(3661));
    layer5_outputs(421) <= not(layer4_outputs(4352));
    layer5_outputs(422) <= (layer4_outputs(2671)) and not (layer4_outputs(1581));
    layer5_outputs(423) <= layer4_outputs(204);
    layer5_outputs(424) <= not(layer4_outputs(2019));
    layer5_outputs(425) <= (layer4_outputs(4038)) or (layer4_outputs(5011));
    layer5_outputs(426) <= layer4_outputs(1435);
    layer5_outputs(427) <= (layer4_outputs(1136)) and not (layer4_outputs(4917));
    layer5_outputs(428) <= layer4_outputs(1808);
    layer5_outputs(429) <= layer4_outputs(3863);
    layer5_outputs(430) <= not(layer4_outputs(509));
    layer5_outputs(431) <= not((layer4_outputs(2393)) or (layer4_outputs(986)));
    layer5_outputs(432) <= layer4_outputs(460);
    layer5_outputs(433) <= not((layer4_outputs(3714)) or (layer4_outputs(1772)));
    layer5_outputs(434) <= not((layer4_outputs(905)) xor (layer4_outputs(626)));
    layer5_outputs(435) <= layer4_outputs(3429);
    layer5_outputs(436) <= not((layer4_outputs(2455)) xor (layer4_outputs(751)));
    layer5_outputs(437) <= not(layer4_outputs(198));
    layer5_outputs(438) <= (layer4_outputs(1888)) xor (layer4_outputs(2456));
    layer5_outputs(439) <= not(layer4_outputs(1478));
    layer5_outputs(440) <= layer4_outputs(816);
    layer5_outputs(441) <= (layer4_outputs(4686)) or (layer4_outputs(2033));
    layer5_outputs(442) <= not(layer4_outputs(3857));
    layer5_outputs(443) <= (layer4_outputs(1879)) and not (layer4_outputs(1611));
    layer5_outputs(444) <= layer4_outputs(2503);
    layer5_outputs(445) <= layer4_outputs(1526);
    layer5_outputs(446) <= not(layer4_outputs(4580));
    layer5_outputs(447) <= not(layer4_outputs(1044));
    layer5_outputs(448) <= (layer4_outputs(994)) and not (layer4_outputs(788));
    layer5_outputs(449) <= layer4_outputs(2577);
    layer5_outputs(450) <= (layer4_outputs(84)) and (layer4_outputs(2946));
    layer5_outputs(451) <= layer4_outputs(4055);
    layer5_outputs(452) <= (layer4_outputs(3526)) and not (layer4_outputs(3553));
    layer5_outputs(453) <= layer4_outputs(5067);
    layer5_outputs(454) <= (layer4_outputs(1640)) or (layer4_outputs(1949));
    layer5_outputs(455) <= not(layer4_outputs(4506));
    layer5_outputs(456) <= not(layer4_outputs(3216));
    layer5_outputs(457) <= not((layer4_outputs(2404)) xor (layer4_outputs(4578)));
    layer5_outputs(458) <= layer4_outputs(4477);
    layer5_outputs(459) <= not(layer4_outputs(4592));
    layer5_outputs(460) <= layer4_outputs(4278);
    layer5_outputs(461) <= not(layer4_outputs(76)) or (layer4_outputs(239));
    layer5_outputs(462) <= not(layer4_outputs(91));
    layer5_outputs(463) <= layer4_outputs(4155);
    layer5_outputs(464) <= (layer4_outputs(2983)) and not (layer4_outputs(1430));
    layer5_outputs(465) <= not(layer4_outputs(3242));
    layer5_outputs(466) <= (layer4_outputs(4401)) and (layer4_outputs(2367));
    layer5_outputs(467) <= (layer4_outputs(3411)) and not (layer4_outputs(1739));
    layer5_outputs(468) <= not(layer4_outputs(2588));
    layer5_outputs(469) <= not((layer4_outputs(2376)) and (layer4_outputs(4539)));
    layer5_outputs(470) <= layer4_outputs(1076);
    layer5_outputs(471) <= layer4_outputs(143);
    layer5_outputs(472) <= (layer4_outputs(3512)) and (layer4_outputs(2318));
    layer5_outputs(473) <= not(layer4_outputs(4194));
    layer5_outputs(474) <= not((layer4_outputs(1010)) xor (layer4_outputs(2235)));
    layer5_outputs(475) <= '1';
    layer5_outputs(476) <= not((layer4_outputs(1804)) or (layer4_outputs(434)));
    layer5_outputs(477) <= '0';
    layer5_outputs(478) <= (layer4_outputs(188)) or (layer4_outputs(324));
    layer5_outputs(479) <= (layer4_outputs(1850)) xor (layer4_outputs(5050));
    layer5_outputs(480) <= (layer4_outputs(3259)) and not (layer4_outputs(752));
    layer5_outputs(481) <= (layer4_outputs(2217)) xor (layer4_outputs(640));
    layer5_outputs(482) <= '0';
    layer5_outputs(483) <= not(layer4_outputs(3657));
    layer5_outputs(484) <= not(layer4_outputs(45));
    layer5_outputs(485) <= layer4_outputs(2194);
    layer5_outputs(486) <= (layer4_outputs(710)) and not (layer4_outputs(5068));
    layer5_outputs(487) <= not(layer4_outputs(5024));
    layer5_outputs(488) <= not(layer4_outputs(511));
    layer5_outputs(489) <= layer4_outputs(3989);
    layer5_outputs(490) <= '0';
    layer5_outputs(491) <= (layer4_outputs(3947)) or (layer4_outputs(727));
    layer5_outputs(492) <= not(layer4_outputs(1041));
    layer5_outputs(493) <= not((layer4_outputs(758)) or (layer4_outputs(2240)));
    layer5_outputs(494) <= layer4_outputs(2761);
    layer5_outputs(495) <= not(layer4_outputs(300));
    layer5_outputs(496) <= not((layer4_outputs(2256)) xor (layer4_outputs(3212)));
    layer5_outputs(497) <= not(layer4_outputs(1722));
    layer5_outputs(498) <= not((layer4_outputs(3422)) and (layer4_outputs(4814)));
    layer5_outputs(499) <= not(layer4_outputs(3157));
    layer5_outputs(500) <= not(layer4_outputs(2415));
    layer5_outputs(501) <= layer4_outputs(1453);
    layer5_outputs(502) <= not(layer4_outputs(2937)) or (layer4_outputs(984));
    layer5_outputs(503) <= (layer4_outputs(499)) and (layer4_outputs(1072));
    layer5_outputs(504) <= layer4_outputs(2912);
    layer5_outputs(505) <= not(layer4_outputs(390));
    layer5_outputs(506) <= layer4_outputs(2024);
    layer5_outputs(507) <= layer4_outputs(3831);
    layer5_outputs(508) <= not((layer4_outputs(320)) xor (layer4_outputs(5064)));
    layer5_outputs(509) <= layer4_outputs(1954);
    layer5_outputs(510) <= not(layer4_outputs(1042));
    layer5_outputs(511) <= (layer4_outputs(1401)) and (layer4_outputs(1667));
    layer5_outputs(512) <= not((layer4_outputs(3494)) and (layer4_outputs(866)));
    layer5_outputs(513) <= (layer4_outputs(2442)) and not (layer4_outputs(2328));
    layer5_outputs(514) <= (layer4_outputs(225)) and (layer4_outputs(1222));
    layer5_outputs(515) <= not(layer4_outputs(1519));
    layer5_outputs(516) <= layer4_outputs(1710);
    layer5_outputs(517) <= not(layer4_outputs(4732));
    layer5_outputs(518) <= not(layer4_outputs(2728));
    layer5_outputs(519) <= not(layer4_outputs(3575));
    layer5_outputs(520) <= '0';
    layer5_outputs(521) <= not((layer4_outputs(159)) xor (layer4_outputs(4112)));
    layer5_outputs(522) <= layer4_outputs(2756);
    layer5_outputs(523) <= not((layer4_outputs(834)) xor (layer4_outputs(1921)));
    layer5_outputs(524) <= not(layer4_outputs(3081));
    layer5_outputs(525) <= (layer4_outputs(840)) xor (layer4_outputs(4243));
    layer5_outputs(526) <= '0';
    layer5_outputs(527) <= not(layer4_outputs(2841)) or (layer4_outputs(2386));
    layer5_outputs(528) <= not(layer4_outputs(1947));
    layer5_outputs(529) <= (layer4_outputs(1510)) or (layer4_outputs(2350));
    layer5_outputs(530) <= not((layer4_outputs(5076)) xor (layer4_outputs(4747)));
    layer5_outputs(531) <= not((layer4_outputs(1520)) and (layer4_outputs(3467)));
    layer5_outputs(532) <= (layer4_outputs(4876)) xor (layer4_outputs(680));
    layer5_outputs(533) <= (layer4_outputs(426)) and (layer4_outputs(5039));
    layer5_outputs(534) <= (layer4_outputs(868)) and not (layer4_outputs(862));
    layer5_outputs(535) <= layer4_outputs(3268);
    layer5_outputs(536) <= layer4_outputs(617);
    layer5_outputs(537) <= not((layer4_outputs(1659)) xor (layer4_outputs(3229)));
    layer5_outputs(538) <= (layer4_outputs(4455)) and not (layer4_outputs(1776));
    layer5_outputs(539) <= layer4_outputs(239);
    layer5_outputs(540) <= (layer4_outputs(3409)) xor (layer4_outputs(3899));
    layer5_outputs(541) <= not(layer4_outputs(4824)) or (layer4_outputs(1083));
    layer5_outputs(542) <= '0';
    layer5_outputs(543) <= not(layer4_outputs(789));
    layer5_outputs(544) <= (layer4_outputs(137)) and not (layer4_outputs(4674));
    layer5_outputs(545) <= (layer4_outputs(486)) and not (layer4_outputs(34));
    layer5_outputs(546) <= layer4_outputs(253);
    layer5_outputs(547) <= layer4_outputs(1683);
    layer5_outputs(548) <= (layer4_outputs(2349)) and not (layer4_outputs(1836));
    layer5_outputs(549) <= not(layer4_outputs(4940));
    layer5_outputs(550) <= layer4_outputs(4705);
    layer5_outputs(551) <= not(layer4_outputs(4602)) or (layer4_outputs(1650));
    layer5_outputs(552) <= layer4_outputs(4521);
    layer5_outputs(553) <= not(layer4_outputs(378)) or (layer4_outputs(3020));
    layer5_outputs(554) <= layer4_outputs(2956);
    layer5_outputs(555) <= layer4_outputs(3959);
    layer5_outputs(556) <= (layer4_outputs(4354)) and not (layer4_outputs(3354));
    layer5_outputs(557) <= layer4_outputs(4065);
    layer5_outputs(558) <= not(layer4_outputs(3389));
    layer5_outputs(559) <= not(layer4_outputs(1040));
    layer5_outputs(560) <= not(layer4_outputs(1549));
    layer5_outputs(561) <= layer4_outputs(50);
    layer5_outputs(562) <= layer4_outputs(3532);
    layer5_outputs(563) <= (layer4_outputs(2115)) xor (layer4_outputs(105));
    layer5_outputs(564) <= layer4_outputs(1179);
    layer5_outputs(565) <= layer4_outputs(4282);
    layer5_outputs(566) <= (layer4_outputs(3094)) and not (layer4_outputs(700));
    layer5_outputs(567) <= (layer4_outputs(1373)) xor (layer4_outputs(2848));
    layer5_outputs(568) <= '1';
    layer5_outputs(569) <= layer4_outputs(4624);
    layer5_outputs(570) <= (layer4_outputs(2088)) or (layer4_outputs(2747));
    layer5_outputs(571) <= not(layer4_outputs(730));
    layer5_outputs(572) <= not((layer4_outputs(4162)) and (layer4_outputs(467)));
    layer5_outputs(573) <= not(layer4_outputs(4329));
    layer5_outputs(574) <= layer4_outputs(1088);
    layer5_outputs(575) <= not(layer4_outputs(3561));
    layer5_outputs(576) <= (layer4_outputs(2967)) xor (layer4_outputs(394));
    layer5_outputs(577) <= layer4_outputs(503);
    layer5_outputs(578) <= not(layer4_outputs(3264));
    layer5_outputs(579) <= layer4_outputs(3085);
    layer5_outputs(580) <= (layer4_outputs(3793)) and not (layer4_outputs(1600));
    layer5_outputs(581) <= (layer4_outputs(4936)) xor (layer4_outputs(3316));
    layer5_outputs(582) <= not(layer4_outputs(3155));
    layer5_outputs(583) <= not((layer4_outputs(354)) or (layer4_outputs(4911)));
    layer5_outputs(584) <= layer4_outputs(570);
    layer5_outputs(585) <= not(layer4_outputs(350));
    layer5_outputs(586) <= not((layer4_outputs(4317)) and (layer4_outputs(1364)));
    layer5_outputs(587) <= (layer4_outputs(2599)) or (layer4_outputs(3043));
    layer5_outputs(588) <= not(layer4_outputs(1189));
    layer5_outputs(589) <= (layer4_outputs(4519)) and not (layer4_outputs(166));
    layer5_outputs(590) <= (layer4_outputs(245)) xor (layer4_outputs(2415));
    layer5_outputs(591) <= not(layer4_outputs(216));
    layer5_outputs(592) <= (layer4_outputs(596)) xor (layer4_outputs(1119));
    layer5_outputs(593) <= not(layer4_outputs(2232));
    layer5_outputs(594) <= not(layer4_outputs(3331));
    layer5_outputs(595) <= not(layer4_outputs(610));
    layer5_outputs(596) <= layer4_outputs(3118);
    layer5_outputs(597) <= not(layer4_outputs(131));
    layer5_outputs(598) <= not(layer4_outputs(32));
    layer5_outputs(599) <= layer4_outputs(59);
    layer5_outputs(600) <= layer4_outputs(3484);
    layer5_outputs(601) <= (layer4_outputs(3933)) and (layer4_outputs(2275));
    layer5_outputs(602) <= layer4_outputs(2256);
    layer5_outputs(603) <= (layer4_outputs(3359)) and not (layer4_outputs(2172));
    layer5_outputs(604) <= not((layer4_outputs(4028)) or (layer4_outputs(551)));
    layer5_outputs(605) <= layer4_outputs(4321);
    layer5_outputs(606) <= '1';
    layer5_outputs(607) <= '0';
    layer5_outputs(608) <= layer4_outputs(1265);
    layer5_outputs(609) <= (layer4_outputs(4247)) and not (layer4_outputs(304));
    layer5_outputs(610) <= not((layer4_outputs(3041)) xor (layer4_outputs(1450)));
    layer5_outputs(611) <= (layer4_outputs(4451)) and not (layer4_outputs(4211));
    layer5_outputs(612) <= not((layer4_outputs(4162)) xor (layer4_outputs(3714)));
    layer5_outputs(613) <= not((layer4_outputs(2012)) and (layer4_outputs(2315)));
    layer5_outputs(614) <= (layer4_outputs(3099)) or (layer4_outputs(4726));
    layer5_outputs(615) <= not(layer4_outputs(3940));
    layer5_outputs(616) <= not(layer4_outputs(1936));
    layer5_outputs(617) <= not(layer4_outputs(4116));
    layer5_outputs(618) <= not(layer4_outputs(4694));
    layer5_outputs(619) <= not(layer4_outputs(2605));
    layer5_outputs(620) <= not(layer4_outputs(2034));
    layer5_outputs(621) <= not(layer4_outputs(1204));
    layer5_outputs(622) <= (layer4_outputs(1482)) and not (layer4_outputs(4064));
    layer5_outputs(623) <= layer4_outputs(3030);
    layer5_outputs(624) <= (layer4_outputs(1472)) xor (layer4_outputs(1692));
    layer5_outputs(625) <= layer4_outputs(4340);
    layer5_outputs(626) <= layer4_outputs(4485);
    layer5_outputs(627) <= '1';
    layer5_outputs(628) <= not(layer4_outputs(920));
    layer5_outputs(629) <= layer4_outputs(4220);
    layer5_outputs(630) <= not(layer4_outputs(2869));
    layer5_outputs(631) <= layer4_outputs(2433);
    layer5_outputs(632) <= not(layer4_outputs(1952)) or (layer4_outputs(2241));
    layer5_outputs(633) <= not(layer4_outputs(1910));
    layer5_outputs(634) <= layer4_outputs(1416);
    layer5_outputs(635) <= (layer4_outputs(1966)) and (layer4_outputs(3583));
    layer5_outputs(636) <= layer4_outputs(3874);
    layer5_outputs(637) <= not(layer4_outputs(100)) or (layer4_outputs(5106));
    layer5_outputs(638) <= not((layer4_outputs(2237)) xor (layer4_outputs(1413)));
    layer5_outputs(639) <= (layer4_outputs(3836)) or (layer4_outputs(3507));
    layer5_outputs(640) <= not((layer4_outputs(4309)) xor (layer4_outputs(3524)));
    layer5_outputs(641) <= not((layer4_outputs(657)) and (layer4_outputs(2039)));
    layer5_outputs(642) <= not(layer4_outputs(4096));
    layer5_outputs(643) <= (layer4_outputs(3630)) and not (layer4_outputs(151));
    layer5_outputs(644) <= not(layer4_outputs(3858)) or (layer4_outputs(2402));
    layer5_outputs(645) <= (layer4_outputs(1064)) and not (layer4_outputs(4524));
    layer5_outputs(646) <= layer4_outputs(1531);
    layer5_outputs(647) <= (layer4_outputs(3250)) and not (layer4_outputs(3843));
    layer5_outputs(648) <= (layer4_outputs(1888)) and not (layer4_outputs(4785));
    layer5_outputs(649) <= layer4_outputs(3501);
    layer5_outputs(650) <= not(layer4_outputs(4268));
    layer5_outputs(651) <= (layer4_outputs(4492)) and not (layer4_outputs(2486));
    layer5_outputs(652) <= layer4_outputs(1469);
    layer5_outputs(653) <= not(layer4_outputs(4727));
    layer5_outputs(654) <= layer4_outputs(874);
    layer5_outputs(655) <= (layer4_outputs(4551)) or (layer4_outputs(377));
    layer5_outputs(656) <= (layer4_outputs(2444)) and not (layer4_outputs(4327));
    layer5_outputs(657) <= layer4_outputs(3083);
    layer5_outputs(658) <= not((layer4_outputs(3818)) or (layer4_outputs(3123)));
    layer5_outputs(659) <= layer4_outputs(717);
    layer5_outputs(660) <= (layer4_outputs(3548)) or (layer4_outputs(888));
    layer5_outputs(661) <= not((layer4_outputs(4809)) and (layer4_outputs(5056)));
    layer5_outputs(662) <= (layer4_outputs(3442)) and not (layer4_outputs(3048));
    layer5_outputs(663) <= (layer4_outputs(114)) and not (layer4_outputs(4255));
    layer5_outputs(664) <= not((layer4_outputs(1396)) and (layer4_outputs(5)));
    layer5_outputs(665) <= layer4_outputs(1448);
    layer5_outputs(666) <= not((layer4_outputs(343)) and (layer4_outputs(3497)));
    layer5_outputs(667) <= not((layer4_outputs(4117)) xor (layer4_outputs(579)));
    layer5_outputs(668) <= layer4_outputs(3769);
    layer5_outputs(669) <= not(layer4_outputs(3652));
    layer5_outputs(670) <= '1';
    layer5_outputs(671) <= not(layer4_outputs(4293));
    layer5_outputs(672) <= layer4_outputs(1455);
    layer5_outputs(673) <= not(layer4_outputs(2906));
    layer5_outputs(674) <= not((layer4_outputs(1399)) or (layer4_outputs(4864)));
    layer5_outputs(675) <= layer4_outputs(1392);
    layer5_outputs(676) <= (layer4_outputs(4199)) or (layer4_outputs(4423));
    layer5_outputs(677) <= not(layer4_outputs(2921));
    layer5_outputs(678) <= layer4_outputs(1572);
    layer5_outputs(679) <= layer4_outputs(3041);
    layer5_outputs(680) <= not(layer4_outputs(971));
    layer5_outputs(681) <= (layer4_outputs(4312)) or (layer4_outputs(2029));
    layer5_outputs(682) <= layer4_outputs(155);
    layer5_outputs(683) <= not(layer4_outputs(2016));
    layer5_outputs(684) <= (layer4_outputs(2994)) and not (layer4_outputs(236));
    layer5_outputs(685) <= layer4_outputs(3046);
    layer5_outputs(686) <= layer4_outputs(3827);
    layer5_outputs(687) <= layer4_outputs(3507);
    layer5_outputs(688) <= not(layer4_outputs(3912));
    layer5_outputs(689) <= not((layer4_outputs(4625)) xor (layer4_outputs(3141)));
    layer5_outputs(690) <= (layer4_outputs(4061)) and not (layer4_outputs(2425));
    layer5_outputs(691) <= not((layer4_outputs(1108)) and (layer4_outputs(4474)));
    layer5_outputs(692) <= (layer4_outputs(4792)) and not (layer4_outputs(3125));
    layer5_outputs(693) <= not(layer4_outputs(659));
    layer5_outputs(694) <= (layer4_outputs(1829)) or (layer4_outputs(1524));
    layer5_outputs(695) <= layer4_outputs(3648);
    layer5_outputs(696) <= layer4_outputs(4384);
    layer5_outputs(697) <= layer4_outputs(1882);
    layer5_outputs(698) <= (layer4_outputs(1883)) and not (layer4_outputs(1308));
    layer5_outputs(699) <= (layer4_outputs(2865)) and (layer4_outputs(3253));
    layer5_outputs(700) <= not(layer4_outputs(1327)) or (layer4_outputs(2203));
    layer5_outputs(701) <= layer4_outputs(2135);
    layer5_outputs(702) <= layer4_outputs(1905);
    layer5_outputs(703) <= (layer4_outputs(4948)) and not (layer4_outputs(4450));
    layer5_outputs(704) <= not(layer4_outputs(3800));
    layer5_outputs(705) <= layer4_outputs(2358);
    layer5_outputs(706) <= '1';
    layer5_outputs(707) <= not(layer4_outputs(1293)) or (layer4_outputs(522));
    layer5_outputs(708) <= (layer4_outputs(2435)) and not (layer4_outputs(4249));
    layer5_outputs(709) <= not(layer4_outputs(2468));
    layer5_outputs(710) <= layer4_outputs(3699);
    layer5_outputs(711) <= layer4_outputs(672);
    layer5_outputs(712) <= (layer4_outputs(757)) and not (layer4_outputs(906));
    layer5_outputs(713) <= not(layer4_outputs(2033));
    layer5_outputs(714) <= not(layer4_outputs(3337)) or (layer4_outputs(4925));
    layer5_outputs(715) <= layer4_outputs(4553);
    layer5_outputs(716) <= layer4_outputs(4659);
    layer5_outputs(717) <= (layer4_outputs(2862)) xor (layer4_outputs(2688));
    layer5_outputs(718) <= not((layer4_outputs(3753)) xor (layer4_outputs(1560)));
    layer5_outputs(719) <= not(layer4_outputs(1136));
    layer5_outputs(720) <= layer4_outputs(4909);
    layer5_outputs(721) <= not(layer4_outputs(1561)) or (layer4_outputs(4649));
    layer5_outputs(722) <= not(layer4_outputs(429)) or (layer4_outputs(1213));
    layer5_outputs(723) <= not((layer4_outputs(3)) xor (layer4_outputs(3662)));
    layer5_outputs(724) <= (layer4_outputs(5034)) xor (layer4_outputs(1664));
    layer5_outputs(725) <= not(layer4_outputs(1836));
    layer5_outputs(726) <= layer4_outputs(4668);
    layer5_outputs(727) <= not((layer4_outputs(1013)) or (layer4_outputs(1385)));
    layer5_outputs(728) <= layer4_outputs(3172);
    layer5_outputs(729) <= not(layer4_outputs(518));
    layer5_outputs(730) <= not(layer4_outputs(4026));
    layer5_outputs(731) <= not(layer4_outputs(1654)) or (layer4_outputs(3304));
    layer5_outputs(732) <= (layer4_outputs(1081)) and not (layer4_outputs(814));
    layer5_outputs(733) <= (layer4_outputs(4322)) and not (layer4_outputs(2903));
    layer5_outputs(734) <= '0';
    layer5_outputs(735) <= not(layer4_outputs(335)) or (layer4_outputs(946));
    layer5_outputs(736) <= (layer4_outputs(262)) and not (layer4_outputs(502));
    layer5_outputs(737) <= not(layer4_outputs(4399));
    layer5_outputs(738) <= (layer4_outputs(2700)) and not (layer4_outputs(3881));
    layer5_outputs(739) <= layer4_outputs(4534);
    layer5_outputs(740) <= not((layer4_outputs(3477)) xor (layer4_outputs(4879)));
    layer5_outputs(741) <= not(layer4_outputs(5056)) or (layer4_outputs(3788));
    layer5_outputs(742) <= (layer4_outputs(1747)) or (layer4_outputs(4633));
    layer5_outputs(743) <= '0';
    layer5_outputs(744) <= layer4_outputs(4108);
    layer5_outputs(745) <= layer4_outputs(3262);
    layer5_outputs(746) <= not(layer4_outputs(106));
    layer5_outputs(747) <= not(layer4_outputs(2076)) or (layer4_outputs(2401));
    layer5_outputs(748) <= layer4_outputs(1383);
    layer5_outputs(749) <= layer4_outputs(1762);
    layer5_outputs(750) <= '1';
    layer5_outputs(751) <= (layer4_outputs(1027)) and (layer4_outputs(4417));
    layer5_outputs(752) <= not((layer4_outputs(2492)) or (layer4_outputs(271)));
    layer5_outputs(753) <= not(layer4_outputs(2915));
    layer5_outputs(754) <= not(layer4_outputs(2581));
    layer5_outputs(755) <= not(layer4_outputs(4076));
    layer5_outputs(756) <= layer4_outputs(2837);
    layer5_outputs(757) <= not(layer4_outputs(2850));
    layer5_outputs(758) <= not(layer4_outputs(487));
    layer5_outputs(759) <= layer4_outputs(4120);
    layer5_outputs(760) <= not((layer4_outputs(4123)) xor (layer4_outputs(533)));
    layer5_outputs(761) <= not(layer4_outputs(4101));
    layer5_outputs(762) <= layer4_outputs(1756);
    layer5_outputs(763) <= not(layer4_outputs(2087));
    layer5_outputs(764) <= not(layer4_outputs(265));
    layer5_outputs(765) <= layer4_outputs(231);
    layer5_outputs(766) <= not((layer4_outputs(1089)) or (layer4_outputs(3656)));
    layer5_outputs(767) <= (layer4_outputs(2359)) xor (layer4_outputs(386));
    layer5_outputs(768) <= not(layer4_outputs(2074));
    layer5_outputs(769) <= not(layer4_outputs(2212));
    layer5_outputs(770) <= (layer4_outputs(1841)) and not (layer4_outputs(4983));
    layer5_outputs(771) <= layer4_outputs(1687);
    layer5_outputs(772) <= layer4_outputs(3613);
    layer5_outputs(773) <= (layer4_outputs(746)) and not (layer4_outputs(1342));
    layer5_outputs(774) <= not(layer4_outputs(4159));
    layer5_outputs(775) <= not(layer4_outputs(48));
    layer5_outputs(776) <= layer4_outputs(3521);
    layer5_outputs(777) <= layer4_outputs(4225);
    layer5_outputs(778) <= not(layer4_outputs(4694));
    layer5_outputs(779) <= (layer4_outputs(2542)) or (layer4_outputs(80));
    layer5_outputs(780) <= (layer4_outputs(652)) and not (layer4_outputs(4375));
    layer5_outputs(781) <= not(layer4_outputs(2646));
    layer5_outputs(782) <= (layer4_outputs(3605)) or (layer4_outputs(1055));
    layer5_outputs(783) <= not(layer4_outputs(2461)) or (layer4_outputs(2233));
    layer5_outputs(784) <= (layer4_outputs(2757)) and not (layer4_outputs(1631));
    layer5_outputs(785) <= (layer4_outputs(542)) or (layer4_outputs(2320));
    layer5_outputs(786) <= layer4_outputs(2677);
    layer5_outputs(787) <= (layer4_outputs(417)) xor (layer4_outputs(1867));
    layer5_outputs(788) <= layer4_outputs(4778);
    layer5_outputs(789) <= not((layer4_outputs(531)) xor (layer4_outputs(3285)));
    layer5_outputs(790) <= layer4_outputs(5018);
    layer5_outputs(791) <= layer4_outputs(4009);
    layer5_outputs(792) <= layer4_outputs(2749);
    layer5_outputs(793) <= not(layer4_outputs(1228));
    layer5_outputs(794) <= not(layer4_outputs(274));
    layer5_outputs(795) <= not((layer4_outputs(3329)) and (layer4_outputs(374)));
    layer5_outputs(796) <= (layer4_outputs(1459)) xor (layer4_outputs(5040));
    layer5_outputs(797) <= not(layer4_outputs(1241));
    layer5_outputs(798) <= not((layer4_outputs(3554)) and (layer4_outputs(2544)));
    layer5_outputs(799) <= not(layer4_outputs(957));
    layer5_outputs(800) <= layer4_outputs(2558);
    layer5_outputs(801) <= (layer4_outputs(2900)) and not (layer4_outputs(97));
    layer5_outputs(802) <= layer4_outputs(1125);
    layer5_outputs(803) <= layer4_outputs(1218);
    layer5_outputs(804) <= (layer4_outputs(2143)) and (layer4_outputs(2488));
    layer5_outputs(805) <= (layer4_outputs(3525)) and (layer4_outputs(1411));
    layer5_outputs(806) <= layer4_outputs(4192);
    layer5_outputs(807) <= not(layer4_outputs(2661));
    layer5_outputs(808) <= layer4_outputs(1245);
    layer5_outputs(809) <= layer4_outputs(3314);
    layer5_outputs(810) <= layer4_outputs(1937);
    layer5_outputs(811) <= (layer4_outputs(2312)) and (layer4_outputs(4494));
    layer5_outputs(812) <= layer4_outputs(52);
    layer5_outputs(813) <= not(layer4_outputs(2065)) or (layer4_outputs(1993));
    layer5_outputs(814) <= layer4_outputs(1513);
    layer5_outputs(815) <= layer4_outputs(2621);
    layer5_outputs(816) <= not((layer4_outputs(3436)) xor (layer4_outputs(1344)));
    layer5_outputs(817) <= not(layer4_outputs(2792));
    layer5_outputs(818) <= not(layer4_outputs(4347));
    layer5_outputs(819) <= layer4_outputs(1461);
    layer5_outputs(820) <= not(layer4_outputs(3427));
    layer5_outputs(821) <= (layer4_outputs(3743)) and not (layer4_outputs(4405));
    layer5_outputs(822) <= layer4_outputs(4646);
    layer5_outputs(823) <= layer4_outputs(4083);
    layer5_outputs(824) <= layer4_outputs(1564);
    layer5_outputs(825) <= layer4_outputs(2010);
    layer5_outputs(826) <= not(layer4_outputs(303));
    layer5_outputs(827) <= not(layer4_outputs(4370));
    layer5_outputs(828) <= not(layer4_outputs(3981));
    layer5_outputs(829) <= (layer4_outputs(2305)) and not (layer4_outputs(1563));
    layer5_outputs(830) <= not(layer4_outputs(2684));
    layer5_outputs(831) <= layer4_outputs(2188);
    layer5_outputs(832) <= not(layer4_outputs(1436));
    layer5_outputs(833) <= layer4_outputs(2);
    layer5_outputs(834) <= layer4_outputs(1833);
    layer5_outputs(835) <= (layer4_outputs(1550)) or (layer4_outputs(3500));
    layer5_outputs(836) <= not(layer4_outputs(824));
    layer5_outputs(837) <= layer4_outputs(252);
    layer5_outputs(838) <= not(layer4_outputs(268));
    layer5_outputs(839) <= not(layer4_outputs(4676));
    layer5_outputs(840) <= not((layer4_outputs(4093)) or (layer4_outputs(3401)));
    layer5_outputs(841) <= layer4_outputs(3273);
    layer5_outputs(842) <= layer4_outputs(1525);
    layer5_outputs(843) <= not(layer4_outputs(2041)) or (layer4_outputs(1781));
    layer5_outputs(844) <= not((layer4_outputs(1983)) and (layer4_outputs(2272)));
    layer5_outputs(845) <= not(layer4_outputs(3952)) or (layer4_outputs(4830));
    layer5_outputs(846) <= not(layer4_outputs(1316));
    layer5_outputs(847) <= not((layer4_outputs(2573)) or (layer4_outputs(2098)));
    layer5_outputs(848) <= not(layer4_outputs(4791));
    layer5_outputs(849) <= not(layer4_outputs(4827));
    layer5_outputs(850) <= not(layer4_outputs(2153));
    layer5_outputs(851) <= not((layer4_outputs(4537)) and (layer4_outputs(2964)));
    layer5_outputs(852) <= not(layer4_outputs(4587));
    layer5_outputs(853) <= (layer4_outputs(101)) and not (layer4_outputs(654));
    layer5_outputs(854) <= (layer4_outputs(1284)) and not (layer4_outputs(4979));
    layer5_outputs(855) <= layer4_outputs(509);
    layer5_outputs(856) <= layer4_outputs(983);
    layer5_outputs(857) <= not(layer4_outputs(668));
    layer5_outputs(858) <= layer4_outputs(799);
    layer5_outputs(859) <= layer4_outputs(2102);
    layer5_outputs(860) <= layer4_outputs(1709);
    layer5_outputs(861) <= layer4_outputs(3289);
    layer5_outputs(862) <= not(layer4_outputs(4090));
    layer5_outputs(863) <= not((layer4_outputs(3225)) and (layer4_outputs(641)));
    layer5_outputs(864) <= not(layer4_outputs(2419)) or (layer4_outputs(124));
    layer5_outputs(865) <= layer4_outputs(3082);
    layer5_outputs(866) <= (layer4_outputs(1138)) and not (layer4_outputs(1908));
    layer5_outputs(867) <= layer4_outputs(1673);
    layer5_outputs(868) <= not((layer4_outputs(11)) xor (layer4_outputs(1056)));
    layer5_outputs(869) <= (layer4_outputs(2712)) xor (layer4_outputs(196));
    layer5_outputs(870) <= layer4_outputs(2382);
    layer5_outputs(871) <= not(layer4_outputs(3152)) or (layer4_outputs(1584));
    layer5_outputs(872) <= layer4_outputs(1381);
    layer5_outputs(873) <= not(layer4_outputs(3018)) or (layer4_outputs(3818));
    layer5_outputs(874) <= not((layer4_outputs(462)) and (layer4_outputs(283)));
    layer5_outputs(875) <= not((layer4_outputs(1267)) and (layer4_outputs(4651)));
    layer5_outputs(876) <= layer4_outputs(3723);
    layer5_outputs(877) <= layer4_outputs(2636);
    layer5_outputs(878) <= not((layer4_outputs(2001)) or (layer4_outputs(4035)));
    layer5_outputs(879) <= not(layer4_outputs(603));
    layer5_outputs(880) <= not((layer4_outputs(2633)) xor (layer4_outputs(769)));
    layer5_outputs(881) <= layer4_outputs(1429);
    layer5_outputs(882) <= layer4_outputs(2979);
    layer5_outputs(883) <= layer4_outputs(2476);
    layer5_outputs(884) <= not(layer4_outputs(1700));
    layer5_outputs(885) <= not(layer4_outputs(3349));
    layer5_outputs(886) <= layer4_outputs(685);
    layer5_outputs(887) <= '1';
    layer5_outputs(888) <= layer4_outputs(415);
    layer5_outputs(889) <= not(layer4_outputs(4730)) or (layer4_outputs(4779));
    layer5_outputs(890) <= not(layer4_outputs(287));
    layer5_outputs(891) <= (layer4_outputs(947)) or (layer4_outputs(4091));
    layer5_outputs(892) <= not(layer4_outputs(1500));
    layer5_outputs(893) <= not(layer4_outputs(4119));
    layer5_outputs(894) <= not(layer4_outputs(576));
    layer5_outputs(895) <= not(layer4_outputs(581));
    layer5_outputs(896) <= not(layer4_outputs(470)) or (layer4_outputs(3196));
    layer5_outputs(897) <= not((layer4_outputs(1126)) xor (layer4_outputs(749)));
    layer5_outputs(898) <= '1';
    layer5_outputs(899) <= (layer4_outputs(1286)) and not (layer4_outputs(1261));
    layer5_outputs(900) <= (layer4_outputs(2337)) and not (layer4_outputs(294));
    layer5_outputs(901) <= not(layer4_outputs(4770));
    layer5_outputs(902) <= not(layer4_outputs(2072)) or (layer4_outputs(4607));
    layer5_outputs(903) <= layer4_outputs(4861);
    layer5_outputs(904) <= not(layer4_outputs(4625)) or (layer4_outputs(1001));
    layer5_outputs(905) <= not(layer4_outputs(2897));
    layer5_outputs(906) <= layer4_outputs(504);
    layer5_outputs(907) <= not(layer4_outputs(3824));
    layer5_outputs(908) <= layer4_outputs(1159);
    layer5_outputs(909) <= not(layer4_outputs(675));
    layer5_outputs(910) <= (layer4_outputs(3008)) and not (layer4_outputs(4007));
    layer5_outputs(911) <= not(layer4_outputs(2428));
    layer5_outputs(912) <= layer4_outputs(166);
    layer5_outputs(913) <= not(layer4_outputs(3722));
    layer5_outputs(914) <= not(layer4_outputs(4251));
    layer5_outputs(915) <= layer4_outputs(700);
    layer5_outputs(916) <= not(layer4_outputs(1320));
    layer5_outputs(917) <= not(layer4_outputs(3774)) or (layer4_outputs(2302));
    layer5_outputs(918) <= not(layer4_outputs(4626));
    layer5_outputs(919) <= layer4_outputs(487);
    layer5_outputs(920) <= (layer4_outputs(159)) xor (layer4_outputs(4433));
    layer5_outputs(921) <= not(layer4_outputs(4466));
    layer5_outputs(922) <= not(layer4_outputs(1041));
    layer5_outputs(923) <= not(layer4_outputs(1617));
    layer5_outputs(924) <= not(layer4_outputs(8));
    layer5_outputs(925) <= (layer4_outputs(1295)) xor (layer4_outputs(117));
    layer5_outputs(926) <= layer4_outputs(2715);
    layer5_outputs(927) <= layer4_outputs(2705);
    layer5_outputs(928) <= (layer4_outputs(1514)) or (layer4_outputs(413));
    layer5_outputs(929) <= not(layer4_outputs(1018));
    layer5_outputs(930) <= (layer4_outputs(1727)) and not (layer4_outputs(4439));
    layer5_outputs(931) <= layer4_outputs(541);
    layer5_outputs(932) <= not((layer4_outputs(652)) and (layer4_outputs(4218)));
    layer5_outputs(933) <= layer4_outputs(4471);
    layer5_outputs(934) <= not(layer4_outputs(4691));
    layer5_outputs(935) <= not(layer4_outputs(4938));
    layer5_outputs(936) <= layer4_outputs(2135);
    layer5_outputs(937) <= not(layer4_outputs(3090));
    layer5_outputs(938) <= (layer4_outputs(4941)) xor (layer4_outputs(3723));
    layer5_outputs(939) <= (layer4_outputs(1079)) xor (layer4_outputs(2363));
    layer5_outputs(940) <= not(layer4_outputs(1149));
    layer5_outputs(941) <= not(layer4_outputs(1120));
    layer5_outputs(942) <= (layer4_outputs(2803)) xor (layer4_outputs(1602));
    layer5_outputs(943) <= (layer4_outputs(4685)) and (layer4_outputs(3926));
    layer5_outputs(944) <= not((layer4_outputs(178)) xor (layer4_outputs(1318)));
    layer5_outputs(945) <= layer4_outputs(3598);
    layer5_outputs(946) <= not((layer4_outputs(1368)) xor (layer4_outputs(1409)));
    layer5_outputs(947) <= (layer4_outputs(4822)) xor (layer4_outputs(980));
    layer5_outputs(948) <= (layer4_outputs(118)) and not (layer4_outputs(1034));
    layer5_outputs(949) <= not(layer4_outputs(767));
    layer5_outputs(950) <= not(layer4_outputs(227));
    layer5_outputs(951) <= (layer4_outputs(567)) xor (layer4_outputs(1911));
    layer5_outputs(952) <= (layer4_outputs(760)) and (layer4_outputs(1729));
    layer5_outputs(953) <= '1';
    layer5_outputs(954) <= not(layer4_outputs(228));
    layer5_outputs(955) <= not((layer4_outputs(4706)) and (layer4_outputs(909)));
    layer5_outputs(956) <= layer4_outputs(2445);
    layer5_outputs(957) <= not((layer4_outputs(2965)) and (layer4_outputs(4273)));
    layer5_outputs(958) <= not(layer4_outputs(3508)) or (layer4_outputs(1655));
    layer5_outputs(959) <= not(layer4_outputs(64));
    layer5_outputs(960) <= layer4_outputs(4316);
    layer5_outputs(961) <= layer4_outputs(3305);
    layer5_outputs(962) <= (layer4_outputs(2604)) and not (layer4_outputs(1766));
    layer5_outputs(963) <= (layer4_outputs(2224)) or (layer4_outputs(257));
    layer5_outputs(964) <= not(layer4_outputs(4968));
    layer5_outputs(965) <= not((layer4_outputs(3299)) xor (layer4_outputs(2368)));
    layer5_outputs(966) <= not(layer4_outputs(4702));
    layer5_outputs(967) <= '1';
    layer5_outputs(968) <= not(layer4_outputs(1283));
    layer5_outputs(969) <= layer4_outputs(3759);
    layer5_outputs(970) <= layer4_outputs(4086);
    layer5_outputs(971) <= (layer4_outputs(2157)) and not (layer4_outputs(2857));
    layer5_outputs(972) <= (layer4_outputs(2455)) and (layer4_outputs(3274));
    layer5_outputs(973) <= not(layer4_outputs(782)) or (layer4_outputs(2710));
    layer5_outputs(974) <= not(layer4_outputs(3871));
    layer5_outputs(975) <= '1';
    layer5_outputs(976) <= layer4_outputs(1264);
    layer5_outputs(977) <= '1';
    layer5_outputs(978) <= layer4_outputs(46);
    layer5_outputs(979) <= not(layer4_outputs(4832));
    layer5_outputs(980) <= not((layer4_outputs(1195)) or (layer4_outputs(3976)));
    layer5_outputs(981) <= not(layer4_outputs(3280));
    layer5_outputs(982) <= not(layer4_outputs(4617));
    layer5_outputs(983) <= not((layer4_outputs(855)) or (layer4_outputs(4458)));
    layer5_outputs(984) <= layer4_outputs(427);
    layer5_outputs(985) <= layer4_outputs(4852);
    layer5_outputs(986) <= not(layer4_outputs(3640));
    layer5_outputs(987) <= layer4_outputs(3565);
    layer5_outputs(988) <= layer4_outputs(3005);
    layer5_outputs(989) <= not(layer4_outputs(4951)) or (layer4_outputs(2659));
    layer5_outputs(990) <= not(layer4_outputs(2734));
    layer5_outputs(991) <= '1';
    layer5_outputs(992) <= (layer4_outputs(2717)) xor (layer4_outputs(2950));
    layer5_outputs(993) <= layer4_outputs(2032);
    layer5_outputs(994) <= not(layer4_outputs(4868)) or (layer4_outputs(4336));
    layer5_outputs(995) <= (layer4_outputs(3717)) or (layer4_outputs(3075));
    layer5_outputs(996) <= not(layer4_outputs(2382));
    layer5_outputs(997) <= not(layer4_outputs(3201)) or (layer4_outputs(126));
    layer5_outputs(998) <= layer4_outputs(1578);
    layer5_outputs(999) <= '0';
    layer5_outputs(1000) <= not((layer4_outputs(712)) or (layer4_outputs(3257)));
    layer5_outputs(1001) <= not(layer4_outputs(2078));
    layer5_outputs(1002) <= (layer4_outputs(4214)) or (layer4_outputs(2343));
    layer5_outputs(1003) <= not((layer4_outputs(2525)) or (layer4_outputs(1423)));
    layer5_outputs(1004) <= '0';
    layer5_outputs(1005) <= not(layer4_outputs(3362)) or (layer4_outputs(911));
    layer5_outputs(1006) <= (layer4_outputs(4423)) and (layer4_outputs(1940));
    layer5_outputs(1007) <= not((layer4_outputs(4927)) xor (layer4_outputs(532)));
    layer5_outputs(1008) <= (layer4_outputs(2357)) and not (layer4_outputs(4234));
    layer5_outputs(1009) <= '1';
    layer5_outputs(1010) <= (layer4_outputs(553)) or (layer4_outputs(1949));
    layer5_outputs(1011) <= layer4_outputs(860);
    layer5_outputs(1012) <= '1';
    layer5_outputs(1013) <= not(layer4_outputs(1090));
    layer5_outputs(1014) <= not(layer4_outputs(4973)) or (layer4_outputs(4871));
    layer5_outputs(1015) <= not((layer4_outputs(4008)) and (layer4_outputs(4031)));
    layer5_outputs(1016) <= not(layer4_outputs(3230));
    layer5_outputs(1017) <= layer4_outputs(4436);
    layer5_outputs(1018) <= '1';
    layer5_outputs(1019) <= not((layer4_outputs(562)) and (layer4_outputs(4108)));
    layer5_outputs(1020) <= (layer4_outputs(2289)) and not (layer4_outputs(2814));
    layer5_outputs(1021) <= '0';
    layer5_outputs(1022) <= layer4_outputs(2516);
    layer5_outputs(1023) <= not(layer4_outputs(3504));
    layer5_outputs(1024) <= layer4_outputs(951);
    layer5_outputs(1025) <= (layer4_outputs(4681)) and not (layer4_outputs(3261));
    layer5_outputs(1026) <= (layer4_outputs(2933)) or (layer4_outputs(1926));
    layer5_outputs(1027) <= (layer4_outputs(1666)) and not (layer4_outputs(2207));
    layer5_outputs(1028) <= not(layer4_outputs(1824));
    layer5_outputs(1029) <= not(layer4_outputs(3291)) or (layer4_outputs(2669));
    layer5_outputs(1030) <= not(layer4_outputs(4692));
    layer5_outputs(1031) <= not(layer4_outputs(3059)) or (layer4_outputs(589));
    layer5_outputs(1032) <= (layer4_outputs(3302)) xor (layer4_outputs(2216));
    layer5_outputs(1033) <= not((layer4_outputs(5102)) xor (layer4_outputs(1279)));
    layer5_outputs(1034) <= not(layer4_outputs(1395));
    layer5_outputs(1035) <= '0';
    layer5_outputs(1036) <= layer4_outputs(3559);
    layer5_outputs(1037) <= layer4_outputs(1926);
    layer5_outputs(1038) <= layer4_outputs(1447);
    layer5_outputs(1039) <= not((layer4_outputs(1371)) xor (layer4_outputs(3333)));
    layer5_outputs(1040) <= not(layer4_outputs(4996)) or (layer4_outputs(1085));
    layer5_outputs(1041) <= not((layer4_outputs(560)) and (layer4_outputs(2830)));
    layer5_outputs(1042) <= not((layer4_outputs(3291)) and (layer4_outputs(3039)));
    layer5_outputs(1043) <= not(layer4_outputs(1644));
    layer5_outputs(1044) <= (layer4_outputs(2407)) xor (layer4_outputs(3425));
    layer5_outputs(1045) <= layer4_outputs(3808);
    layer5_outputs(1046) <= not((layer4_outputs(815)) xor (layer4_outputs(1853)));
    layer5_outputs(1047) <= layer4_outputs(561);
    layer5_outputs(1048) <= layer4_outputs(1916);
    layer5_outputs(1049) <= not(layer4_outputs(270));
    layer5_outputs(1050) <= layer4_outputs(1158);
    layer5_outputs(1051) <= not(layer4_outputs(3255));
    layer5_outputs(1052) <= not(layer4_outputs(210)) or (layer4_outputs(1197));
    layer5_outputs(1053) <= (layer4_outputs(4666)) and not (layer4_outputs(4296));
    layer5_outputs(1054) <= not((layer4_outputs(1742)) xor (layer4_outputs(95)));
    layer5_outputs(1055) <= layer4_outputs(4560);
    layer5_outputs(1056) <= not((layer4_outputs(385)) or (layer4_outputs(4446)));
    layer5_outputs(1057) <= (layer4_outputs(803)) and not (layer4_outputs(3036));
    layer5_outputs(1058) <= (layer4_outputs(4065)) and not (layer4_outputs(598));
    layer5_outputs(1059) <= '1';
    layer5_outputs(1060) <= not(layer4_outputs(2476));
    layer5_outputs(1061) <= not((layer4_outputs(3795)) and (layer4_outputs(3996)));
    layer5_outputs(1062) <= not(layer4_outputs(4968)) or (layer4_outputs(3947));
    layer5_outputs(1063) <= not(layer4_outputs(1738));
    layer5_outputs(1064) <= layer4_outputs(3807);
    layer5_outputs(1065) <= not(layer4_outputs(2820));
    layer5_outputs(1066) <= not(layer4_outputs(1849));
    layer5_outputs(1067) <= not((layer4_outputs(4992)) or (layer4_outputs(3993)));
    layer5_outputs(1068) <= layer4_outputs(3339);
    layer5_outputs(1069) <= not(layer4_outputs(2055)) or (layer4_outputs(4662));
    layer5_outputs(1070) <= not(layer4_outputs(4758)) or (layer4_outputs(5109));
    layer5_outputs(1071) <= layer4_outputs(4462);
    layer5_outputs(1072) <= layer4_outputs(4832);
    layer5_outputs(1073) <= (layer4_outputs(1270)) xor (layer4_outputs(1721));
    layer5_outputs(1074) <= layer4_outputs(4778);
    layer5_outputs(1075) <= not(layer4_outputs(788));
    layer5_outputs(1076) <= not(layer4_outputs(2527));
    layer5_outputs(1077) <= not(layer4_outputs(835));
    layer5_outputs(1078) <= (layer4_outputs(2438)) xor (layer4_outputs(4306));
    layer5_outputs(1079) <= layer4_outputs(3642);
    layer5_outputs(1080) <= not((layer4_outputs(3296)) and (layer4_outputs(4541)));
    layer5_outputs(1081) <= not(layer4_outputs(3871));
    layer5_outputs(1082) <= not(layer4_outputs(1828));
    layer5_outputs(1083) <= not((layer4_outputs(3724)) xor (layer4_outputs(938)));
    layer5_outputs(1084) <= not(layer4_outputs(2096));
    layer5_outputs(1085) <= layer4_outputs(2261);
    layer5_outputs(1086) <= not(layer4_outputs(4257));
    layer5_outputs(1087) <= not((layer4_outputs(3402)) and (layer4_outputs(2106)));
    layer5_outputs(1088) <= not(layer4_outputs(1100));
    layer5_outputs(1089) <= not(layer4_outputs(2503));
    layer5_outputs(1090) <= not(layer4_outputs(2544)) or (layer4_outputs(2745));
    layer5_outputs(1091) <= not(layer4_outputs(1991)) or (layer4_outputs(3547));
    layer5_outputs(1092) <= layer4_outputs(4770);
    layer5_outputs(1093) <= layer4_outputs(2208);
    layer5_outputs(1094) <= not(layer4_outputs(4970));
    layer5_outputs(1095) <= not((layer4_outputs(3228)) or (layer4_outputs(4670)));
    layer5_outputs(1096) <= layer4_outputs(3804);
    layer5_outputs(1097) <= layer4_outputs(2400);
    layer5_outputs(1098) <= not(layer4_outputs(4917)) or (layer4_outputs(4198));
    layer5_outputs(1099) <= layer4_outputs(3630);
    layer5_outputs(1100) <= not((layer4_outputs(2729)) or (layer4_outputs(3979)));
    layer5_outputs(1101) <= not(layer4_outputs(2800)) or (layer4_outputs(2790));
    layer5_outputs(1102) <= layer4_outputs(2157);
    layer5_outputs(1103) <= (layer4_outputs(2335)) or (layer4_outputs(222));
    layer5_outputs(1104) <= not(layer4_outputs(52));
    layer5_outputs(1105) <= (layer4_outputs(172)) and (layer4_outputs(3835));
    layer5_outputs(1106) <= layer4_outputs(1189);
    layer5_outputs(1107) <= not(layer4_outputs(2114)) or (layer4_outputs(310));
    layer5_outputs(1108) <= (layer4_outputs(2703)) xor (layer4_outputs(832));
    layer5_outputs(1109) <= (layer4_outputs(3110)) or (layer4_outputs(4160));
    layer5_outputs(1110) <= (layer4_outputs(638)) xor (layer4_outputs(3221));
    layer5_outputs(1111) <= not(layer4_outputs(2375)) or (layer4_outputs(3336));
    layer5_outputs(1112) <= not(layer4_outputs(2364));
    layer5_outputs(1113) <= (layer4_outputs(1689)) and not (layer4_outputs(4097));
    layer5_outputs(1114) <= (layer4_outputs(2065)) or (layer4_outputs(2143));
    layer5_outputs(1115) <= (layer4_outputs(2374)) or (layer4_outputs(833));
    layer5_outputs(1116) <= not((layer4_outputs(3100)) or (layer4_outputs(4939)));
    layer5_outputs(1117) <= not(layer4_outputs(1012)) or (layer4_outputs(3870));
    layer5_outputs(1118) <= (layer4_outputs(2960)) and not (layer4_outputs(3265));
    layer5_outputs(1119) <= '0';
    layer5_outputs(1120) <= not(layer4_outputs(1166)) or (layer4_outputs(4721));
    layer5_outputs(1121) <= not((layer4_outputs(3845)) or (layer4_outputs(4101)));
    layer5_outputs(1122) <= layer4_outputs(3516);
    layer5_outputs(1123) <= not(layer4_outputs(1767));
    layer5_outputs(1124) <= not(layer4_outputs(439)) or (layer4_outputs(1460));
    layer5_outputs(1125) <= layer4_outputs(4317);
    layer5_outputs(1126) <= not(layer4_outputs(139)) or (layer4_outputs(406));
    layer5_outputs(1127) <= '1';
    layer5_outputs(1128) <= not(layer4_outputs(241)) or (layer4_outputs(2115));
    layer5_outputs(1129) <= layer4_outputs(4712);
    layer5_outputs(1130) <= (layer4_outputs(3825)) and not (layer4_outputs(1163));
    layer5_outputs(1131) <= not(layer4_outputs(4033));
    layer5_outputs(1132) <= not(layer4_outputs(399));
    layer5_outputs(1133) <= (layer4_outputs(4728)) and (layer4_outputs(5097));
    layer5_outputs(1134) <= (layer4_outputs(696)) and (layer4_outputs(1691));
    layer5_outputs(1135) <= layer4_outputs(2474);
    layer5_outputs(1136) <= (layer4_outputs(3115)) and (layer4_outputs(1376));
    layer5_outputs(1137) <= (layer4_outputs(1885)) and (layer4_outputs(5116));
    layer5_outputs(1138) <= (layer4_outputs(3312)) xor (layer4_outputs(2479));
    layer5_outputs(1139) <= not(layer4_outputs(3274));
    layer5_outputs(1140) <= not(layer4_outputs(1445));
    layer5_outputs(1141) <= (layer4_outputs(2892)) and not (layer4_outputs(761));
    layer5_outputs(1142) <= layer4_outputs(849);
    layer5_outputs(1143) <= not(layer4_outputs(4568));
    layer5_outputs(1144) <= not(layer4_outputs(3578));
    layer5_outputs(1145) <= (layer4_outputs(3617)) xor (layer4_outputs(4257));
    layer5_outputs(1146) <= not(layer4_outputs(353));
    layer5_outputs(1147) <= not(layer4_outputs(958)) or (layer4_outputs(2226));
    layer5_outputs(1148) <= (layer4_outputs(1979)) and not (layer4_outputs(330));
    layer5_outputs(1149) <= not((layer4_outputs(4545)) or (layer4_outputs(1657)));
    layer5_outputs(1150) <= not(layer4_outputs(592));
    layer5_outputs(1151) <= '0';
    layer5_outputs(1152) <= '1';
    layer5_outputs(1153) <= (layer4_outputs(3319)) and not (layer4_outputs(2561));
    layer5_outputs(1154) <= not(layer4_outputs(4534));
    layer5_outputs(1155) <= layer4_outputs(2910);
    layer5_outputs(1156) <= not((layer4_outputs(4538)) and (layer4_outputs(2419)));
    layer5_outputs(1157) <= (layer4_outputs(2556)) and (layer4_outputs(2491));
    layer5_outputs(1158) <= (layer4_outputs(2467)) and not (layer4_outputs(4324));
    layer5_outputs(1159) <= not((layer4_outputs(423)) xor (layer4_outputs(3213)));
    layer5_outputs(1160) <= not(layer4_outputs(4271));
    layer5_outputs(1161) <= not((layer4_outputs(4918)) and (layer4_outputs(137)));
    layer5_outputs(1162) <= not(layer4_outputs(2514)) or (layer4_outputs(577));
    layer5_outputs(1163) <= (layer4_outputs(3930)) or (layer4_outputs(3875));
    layer5_outputs(1164) <= (layer4_outputs(4228)) or (layer4_outputs(2946));
    layer5_outputs(1165) <= layer4_outputs(3040);
    layer5_outputs(1166) <= not(layer4_outputs(1086));
    layer5_outputs(1167) <= layer4_outputs(4881);
    layer5_outputs(1168) <= not(layer4_outputs(4999));
    layer5_outputs(1169) <= (layer4_outputs(2809)) and (layer4_outputs(3978));
    layer5_outputs(1170) <= (layer4_outputs(2548)) or (layer4_outputs(3925));
    layer5_outputs(1171) <= not(layer4_outputs(4367));
    layer5_outputs(1172) <= '1';
    layer5_outputs(1173) <= not(layer4_outputs(4757));
    layer5_outputs(1174) <= not((layer4_outputs(3088)) xor (layer4_outputs(2343)));
    layer5_outputs(1175) <= (layer4_outputs(3649)) and (layer4_outputs(1156));
    layer5_outputs(1176) <= layer4_outputs(4149);
    layer5_outputs(1177) <= (layer4_outputs(2700)) and (layer4_outputs(4514));
    layer5_outputs(1178) <= layer4_outputs(3475);
    layer5_outputs(1179) <= not(layer4_outputs(1629));
    layer5_outputs(1180) <= not(layer4_outputs(3769));
    layer5_outputs(1181) <= layer4_outputs(2015);
    layer5_outputs(1182) <= layer4_outputs(2534);
    layer5_outputs(1183) <= layer4_outputs(1999);
    layer5_outputs(1184) <= layer4_outputs(5070);
    layer5_outputs(1185) <= not(layer4_outputs(4020)) or (layer4_outputs(2944));
    layer5_outputs(1186) <= (layer4_outputs(298)) or (layer4_outputs(1108));
    layer5_outputs(1187) <= not((layer4_outputs(1343)) xor (layer4_outputs(1535)));
    layer5_outputs(1188) <= not(layer4_outputs(2925));
    layer5_outputs(1189) <= not((layer4_outputs(353)) xor (layer4_outputs(960)));
    layer5_outputs(1190) <= not((layer4_outputs(3042)) xor (layer4_outputs(2100)));
    layer5_outputs(1191) <= not(layer4_outputs(1311));
    layer5_outputs(1192) <= not(layer4_outputs(3556));
    layer5_outputs(1193) <= '1';
    layer5_outputs(1194) <= layer4_outputs(1181);
    layer5_outputs(1195) <= not((layer4_outputs(1838)) or (layer4_outputs(455)));
    layer5_outputs(1196) <= not((layer4_outputs(555)) and (layer4_outputs(1643)));
    layer5_outputs(1197) <= not(layer4_outputs(3954));
    layer5_outputs(1198) <= not(layer4_outputs(4016));
    layer5_outputs(1199) <= layer4_outputs(276);
    layer5_outputs(1200) <= not((layer4_outputs(3150)) and (layer4_outputs(4114)));
    layer5_outputs(1201) <= (layer4_outputs(4572)) and not (layer4_outputs(3544));
    layer5_outputs(1202) <= not(layer4_outputs(3564)) or (layer4_outputs(3896));
    layer5_outputs(1203) <= (layer4_outputs(2389)) xor (layer4_outputs(2179));
    layer5_outputs(1204) <= not((layer4_outputs(4272)) and (layer4_outputs(2915)));
    layer5_outputs(1205) <= not(layer4_outputs(1381));
    layer5_outputs(1206) <= not((layer4_outputs(4571)) xor (layer4_outputs(1822)));
    layer5_outputs(1207) <= not((layer4_outputs(2603)) xor (layer4_outputs(4772)));
    layer5_outputs(1208) <= layer4_outputs(4821);
    layer5_outputs(1209) <= not(layer4_outputs(391));
    layer5_outputs(1210) <= not((layer4_outputs(3693)) or (layer4_outputs(3279)));
    layer5_outputs(1211) <= layer4_outputs(4961);
    layer5_outputs(1212) <= (layer4_outputs(4416)) or (layer4_outputs(1323));
    layer5_outputs(1213) <= not(layer4_outputs(4234));
    layer5_outputs(1214) <= not(layer4_outputs(426));
    layer5_outputs(1215) <= layer4_outputs(4110);
    layer5_outputs(1216) <= not(layer4_outputs(3999)) or (layer4_outputs(3290));
    layer5_outputs(1217) <= layer4_outputs(4044);
    layer5_outputs(1218) <= not(layer4_outputs(3204));
    layer5_outputs(1219) <= not((layer4_outputs(3576)) xor (layer4_outputs(1577)));
    layer5_outputs(1220) <= not(layer4_outputs(386));
    layer5_outputs(1221) <= (layer4_outputs(1325)) and (layer4_outputs(4325));
    layer5_outputs(1222) <= layer4_outputs(1670);
    layer5_outputs(1223) <= (layer4_outputs(3838)) xor (layer4_outputs(214));
    layer5_outputs(1224) <= layer4_outputs(1174);
    layer5_outputs(1225) <= layer4_outputs(4280);
    layer5_outputs(1226) <= (layer4_outputs(2630)) and not (layer4_outputs(3204));
    layer5_outputs(1227) <= layer4_outputs(3346);
    layer5_outputs(1228) <= layer4_outputs(1874);
    layer5_outputs(1229) <= layer4_outputs(221);
    layer5_outputs(1230) <= (layer4_outputs(4566)) or (layer4_outputs(347));
    layer5_outputs(1231) <= layer4_outputs(1547);
    layer5_outputs(1232) <= (layer4_outputs(2083)) and not (layer4_outputs(3853));
    layer5_outputs(1233) <= layer4_outputs(718);
    layer5_outputs(1234) <= not(layer4_outputs(996));
    layer5_outputs(1235) <= not(layer4_outputs(32));
    layer5_outputs(1236) <= (layer4_outputs(54)) and not (layer4_outputs(1718));
    layer5_outputs(1237) <= not(layer4_outputs(4095));
    layer5_outputs(1238) <= not(layer4_outputs(3174));
    layer5_outputs(1239) <= layer4_outputs(4740);
    layer5_outputs(1240) <= layer4_outputs(800);
    layer5_outputs(1241) <= not(layer4_outputs(624));
    layer5_outputs(1242) <= (layer4_outputs(2403)) and (layer4_outputs(476));
    layer5_outputs(1243) <= (layer4_outputs(4576)) and (layer4_outputs(643));
    layer5_outputs(1244) <= not(layer4_outputs(410));
    layer5_outputs(1245) <= layer4_outputs(179);
    layer5_outputs(1246) <= (layer4_outputs(3307)) or (layer4_outputs(3017));
    layer5_outputs(1247) <= not((layer4_outputs(4739)) xor (layer4_outputs(4696)));
    layer5_outputs(1248) <= (layer4_outputs(2159)) xor (layer4_outputs(550));
    layer5_outputs(1249) <= layer4_outputs(2448);
    layer5_outputs(1250) <= layer4_outputs(39);
    layer5_outputs(1251) <= layer4_outputs(2907);
    layer5_outputs(1252) <= (layer4_outputs(2786)) and (layer4_outputs(2632));
    layer5_outputs(1253) <= not(layer4_outputs(73));
    layer5_outputs(1254) <= not((layer4_outputs(4279)) or (layer4_outputs(232)));
    layer5_outputs(1255) <= not((layer4_outputs(2779)) or (layer4_outputs(764)));
    layer5_outputs(1256) <= layer4_outputs(1917);
    layer5_outputs(1257) <= not(layer4_outputs(619));
    layer5_outputs(1258) <= not((layer4_outputs(4305)) xor (layer4_outputs(4166)));
    layer5_outputs(1259) <= not(layer4_outputs(4759));
    layer5_outputs(1260) <= layer4_outputs(3278);
    layer5_outputs(1261) <= not(layer4_outputs(2432));
    layer5_outputs(1262) <= not(layer4_outputs(498)) or (layer4_outputs(3847));
    layer5_outputs(1263) <= '1';
    layer5_outputs(1264) <= '1';
    layer5_outputs(1265) <= '0';
    layer5_outputs(1266) <= '1';
    layer5_outputs(1267) <= not(layer4_outputs(1119));
    layer5_outputs(1268) <= not(layer4_outputs(3054));
    layer5_outputs(1269) <= layer4_outputs(2473);
    layer5_outputs(1270) <= not((layer4_outputs(4052)) or (layer4_outputs(4028)));
    layer5_outputs(1271) <= not(layer4_outputs(4444));
    layer5_outputs(1272) <= not(layer4_outputs(3137));
    layer5_outputs(1273) <= not(layer4_outputs(2187));
    layer5_outputs(1274) <= layer4_outputs(748);
    layer5_outputs(1275) <= (layer4_outputs(4181)) xor (layer4_outputs(4223));
    layer5_outputs(1276) <= not((layer4_outputs(3645)) or (layer4_outputs(4490)));
    layer5_outputs(1277) <= not((layer4_outputs(2586)) xor (layer4_outputs(2797)));
    layer5_outputs(1278) <= not((layer4_outputs(522)) xor (layer4_outputs(4518)));
    layer5_outputs(1279) <= (layer4_outputs(741)) and not (layer4_outputs(4703));
    layer5_outputs(1280) <= layer4_outputs(2175);
    layer5_outputs(1281) <= layer4_outputs(2720);
    layer5_outputs(1282) <= layer4_outputs(3348);
    layer5_outputs(1283) <= layer4_outputs(4250);
    layer5_outputs(1284) <= not(layer4_outputs(3007));
    layer5_outputs(1285) <= '0';
    layer5_outputs(1286) <= not(layer4_outputs(2999));
    layer5_outputs(1287) <= not(layer4_outputs(2893));
    layer5_outputs(1288) <= not(layer4_outputs(4747)) or (layer4_outputs(1391));
    layer5_outputs(1289) <= not((layer4_outputs(148)) and (layer4_outputs(4323)));
    layer5_outputs(1290) <= not((layer4_outputs(3052)) and (layer4_outputs(3909)));
    layer5_outputs(1291) <= '0';
    layer5_outputs(1292) <= layer4_outputs(3286);
    layer5_outputs(1293) <= not(layer4_outputs(1633));
    layer5_outputs(1294) <= (layer4_outputs(1221)) and not (layer4_outputs(4157));
    layer5_outputs(1295) <= layer4_outputs(1870);
    layer5_outputs(1296) <= not(layer4_outputs(710)) or (layer4_outputs(1442));
    layer5_outputs(1297) <= not(layer4_outputs(2559)) or (layer4_outputs(35));
    layer5_outputs(1298) <= (layer4_outputs(3390)) and not (layer4_outputs(978));
    layer5_outputs(1299) <= (layer4_outputs(2856)) and not (layer4_outputs(1930));
    layer5_outputs(1300) <= not(layer4_outputs(4100));
    layer5_outputs(1301) <= (layer4_outputs(4147)) or (layer4_outputs(4256));
    layer5_outputs(1302) <= (layer4_outputs(943)) xor (layer4_outputs(3929));
    layer5_outputs(1303) <= not((layer4_outputs(3144)) or (layer4_outputs(2331)));
    layer5_outputs(1304) <= layer4_outputs(2694);
    layer5_outputs(1305) <= (layer4_outputs(3182)) or (layer4_outputs(1540));
    layer5_outputs(1306) <= not(layer4_outputs(2827));
    layer5_outputs(1307) <= not(layer4_outputs(391));
    layer5_outputs(1308) <= layer4_outputs(4952);
    layer5_outputs(1309) <= (layer4_outputs(1925)) and not (layer4_outputs(3629));
    layer5_outputs(1310) <= not(layer4_outputs(4638));
    layer5_outputs(1311) <= (layer4_outputs(3225)) and not (layer4_outputs(203));
    layer5_outputs(1312) <= layer4_outputs(3329);
    layer5_outputs(1313) <= not((layer4_outputs(477)) xor (layer4_outputs(2052)));
    layer5_outputs(1314) <= not(layer4_outputs(1593));
    layer5_outputs(1315) <= layer4_outputs(2367);
    layer5_outputs(1316) <= not(layer4_outputs(3369));
    layer5_outputs(1317) <= not(layer4_outputs(761));
    layer5_outputs(1318) <= not(layer4_outputs(2898));
    layer5_outputs(1319) <= not(layer4_outputs(4289));
    layer5_outputs(1320) <= not(layer4_outputs(2405));
    layer5_outputs(1321) <= (layer4_outputs(1420)) or (layer4_outputs(1107));
    layer5_outputs(1322) <= layer4_outputs(1199);
    layer5_outputs(1323) <= not(layer4_outputs(3584));
    layer5_outputs(1324) <= layer4_outputs(131);
    layer5_outputs(1325) <= (layer4_outputs(3571)) and not (layer4_outputs(4092));
    layer5_outputs(1326) <= not(layer4_outputs(1193));
    layer5_outputs(1327) <= not((layer4_outputs(1430)) or (layer4_outputs(3362)));
    layer5_outputs(1328) <= layer4_outputs(4946);
    layer5_outputs(1329) <= layer4_outputs(2212);
    layer5_outputs(1330) <= not((layer4_outputs(2711)) or (layer4_outputs(3524)));
    layer5_outputs(1331) <= layer4_outputs(1329);
    layer5_outputs(1332) <= not(layer4_outputs(4821));
    layer5_outputs(1333) <= (layer4_outputs(2410)) and not (layer4_outputs(4487));
    layer5_outputs(1334) <= not(layer4_outputs(24));
    layer5_outputs(1335) <= not(layer4_outputs(2973));
    layer5_outputs(1336) <= (layer4_outputs(265)) and not (layer4_outputs(2880));
    layer5_outputs(1337) <= '1';
    layer5_outputs(1338) <= not(layer4_outputs(575)) or (layer4_outputs(5111));
    layer5_outputs(1339) <= not(layer4_outputs(207));
    layer5_outputs(1340) <= (layer4_outputs(332)) and not (layer4_outputs(96));
    layer5_outputs(1341) <= (layer4_outputs(1451)) xor (layer4_outputs(2843));
    layer5_outputs(1342) <= '0';
    layer5_outputs(1343) <= not(layer4_outputs(3688)) or (layer4_outputs(3462));
    layer5_outputs(1344) <= layer4_outputs(1492);
    layer5_outputs(1345) <= layer4_outputs(640);
    layer5_outputs(1346) <= layer4_outputs(871);
    layer5_outputs(1347) <= layer4_outputs(1084);
    layer5_outputs(1348) <= not((layer4_outputs(656)) or (layer4_outputs(1771)));
    layer5_outputs(1349) <= not(layer4_outputs(72));
    layer5_outputs(1350) <= not(layer4_outputs(1537));
    layer5_outputs(1351) <= not((layer4_outputs(4115)) xor (layer4_outputs(1208)));
    layer5_outputs(1352) <= not((layer4_outputs(2136)) and (layer4_outputs(1706)));
    layer5_outputs(1353) <= not(layer4_outputs(4892)) or (layer4_outputs(2282));
    layer5_outputs(1354) <= layer4_outputs(4504);
    layer5_outputs(1355) <= (layer4_outputs(3360)) and (layer4_outputs(4307));
    layer5_outputs(1356) <= layer4_outputs(1472);
    layer5_outputs(1357) <= layer4_outputs(3135);
    layer5_outputs(1358) <= not(layer4_outputs(3883)) or (layer4_outputs(577));
    layer5_outputs(1359) <= not((layer4_outputs(4496)) xor (layer4_outputs(2558)));
    layer5_outputs(1360) <= (layer4_outputs(3578)) and not (layer4_outputs(3937));
    layer5_outputs(1361) <= (layer4_outputs(3514)) and (layer4_outputs(1391));
    layer5_outputs(1362) <= not(layer4_outputs(118)) or (layer4_outputs(3681));
    layer5_outputs(1363) <= (layer4_outputs(2945)) and not (layer4_outputs(1150));
    layer5_outputs(1364) <= not((layer4_outputs(3754)) xor (layer4_outputs(2357)));
    layer5_outputs(1365) <= layer4_outputs(2754);
    layer5_outputs(1366) <= not((layer4_outputs(2932)) xor (layer4_outputs(1191)));
    layer5_outputs(1367) <= not((layer4_outputs(3531)) and (layer4_outputs(1567)));
    layer5_outputs(1368) <= layer4_outputs(4382);
    layer5_outputs(1369) <= layer4_outputs(2058);
    layer5_outputs(1370) <= layer4_outputs(2565);
    layer5_outputs(1371) <= layer4_outputs(839);
    layer5_outputs(1372) <= layer4_outputs(2787);
    layer5_outputs(1373) <= layer4_outputs(3974);
    layer5_outputs(1374) <= not(layer4_outputs(4126));
    layer5_outputs(1375) <= (layer4_outputs(4161)) and not (layer4_outputs(3077));
    layer5_outputs(1376) <= not(layer4_outputs(50));
    layer5_outputs(1377) <= not((layer4_outputs(5094)) and (layer4_outputs(1909)));
    layer5_outputs(1378) <= layer4_outputs(1357);
    layer5_outputs(1379) <= not(layer4_outputs(3651));
    layer5_outputs(1380) <= layer4_outputs(4973);
    layer5_outputs(1381) <= (layer4_outputs(3923)) and (layer4_outputs(2478));
    layer5_outputs(1382) <= not(layer4_outputs(4420));
    layer5_outputs(1383) <= (layer4_outputs(489)) and not (layer4_outputs(2839));
    layer5_outputs(1384) <= not((layer4_outputs(3673)) xor (layer4_outputs(4888)));
    layer5_outputs(1385) <= (layer4_outputs(5009)) or (layer4_outputs(4242));
    layer5_outputs(1386) <= (layer4_outputs(2549)) and not (layer4_outputs(3583));
    layer5_outputs(1387) <= not((layer4_outputs(2288)) and (layer4_outputs(4802)));
    layer5_outputs(1388) <= layer4_outputs(775);
    layer5_outputs(1389) <= not(layer4_outputs(956));
    layer5_outputs(1390) <= not(layer4_outputs(1405));
    layer5_outputs(1391) <= not(layer4_outputs(2122));
    layer5_outputs(1392) <= layer4_outputs(3016);
    layer5_outputs(1393) <= not(layer4_outputs(4062));
    layer5_outputs(1394) <= layer4_outputs(4299);
    layer5_outputs(1395) <= not((layer4_outputs(3396)) and (layer4_outputs(3687)));
    layer5_outputs(1396) <= layer4_outputs(2627);
    layer5_outputs(1397) <= not(layer4_outputs(188)) or (layer4_outputs(3860));
    layer5_outputs(1398) <= not(layer4_outputs(3011));
    layer5_outputs(1399) <= (layer4_outputs(4635)) xor (layer4_outputs(1967));
    layer5_outputs(1400) <= (layer4_outputs(1642)) xor (layer4_outputs(581));
    layer5_outputs(1401) <= layer4_outputs(3819);
    layer5_outputs(1402) <= layer4_outputs(1884);
    layer5_outputs(1403) <= not(layer4_outputs(4269)) or (layer4_outputs(3315));
    layer5_outputs(1404) <= not(layer4_outputs(3761)) or (layer4_outputs(1483));
    layer5_outputs(1405) <= not(layer4_outputs(323));
    layer5_outputs(1406) <= layer4_outputs(748);
    layer5_outputs(1407) <= not(layer4_outputs(1662));
    layer5_outputs(1408) <= not(layer4_outputs(2613));
    layer5_outputs(1409) <= (layer4_outputs(4006)) xor (layer4_outputs(4959));
    layer5_outputs(1410) <= layer4_outputs(678);
    layer5_outputs(1411) <= not(layer4_outputs(4576));
    layer5_outputs(1412) <= not((layer4_outputs(1126)) and (layer4_outputs(4259)));
    layer5_outputs(1413) <= (layer4_outputs(3134)) or (layer4_outputs(3646));
    layer5_outputs(1414) <= (layer4_outputs(2734)) and (layer4_outputs(2470));
    layer5_outputs(1415) <= (layer4_outputs(2585)) or (layer4_outputs(1787));
    layer5_outputs(1416) <= (layer4_outputs(4193)) or (layer4_outputs(2622));
    layer5_outputs(1417) <= not(layer4_outputs(4927)) or (layer4_outputs(67));
    layer5_outputs(1418) <= not((layer4_outputs(3736)) xor (layer4_outputs(1092)));
    layer5_outputs(1419) <= not(layer4_outputs(1025));
    layer5_outputs(1420) <= not(layer4_outputs(1844));
    layer5_outputs(1421) <= not(layer4_outputs(3309));
    layer5_outputs(1422) <= not(layer4_outputs(4252)) or (layer4_outputs(609));
    layer5_outputs(1423) <= layer4_outputs(3756);
    layer5_outputs(1424) <= layer4_outputs(4225);
    layer5_outputs(1425) <= (layer4_outputs(2469)) and not (layer4_outputs(3880));
    layer5_outputs(1426) <= '1';
    layer5_outputs(1427) <= not(layer4_outputs(3282));
    layer5_outputs(1428) <= not(layer4_outputs(3428));
    layer5_outputs(1429) <= (layer4_outputs(3571)) and (layer4_outputs(3245));
    layer5_outputs(1430) <= layer4_outputs(4283);
    layer5_outputs(1431) <= layer4_outputs(4596);
    layer5_outputs(1432) <= not(layer4_outputs(4239));
    layer5_outputs(1433) <= not(layer4_outputs(336));
    layer5_outputs(1434) <= layer4_outputs(636);
    layer5_outputs(1435) <= not(layer4_outputs(4615));
    layer5_outputs(1436) <= not(layer4_outputs(1731)) or (layer4_outputs(2663));
    layer5_outputs(1437) <= not(layer4_outputs(3002));
    layer5_outputs(1438) <= layer4_outputs(1886);
    layer5_outputs(1439) <= (layer4_outputs(202)) or (layer4_outputs(1209));
    layer5_outputs(1440) <= not(layer4_outputs(850));
    layer5_outputs(1441) <= not((layer4_outputs(1023)) xor (layer4_outputs(3846)));
    layer5_outputs(1442) <= not(layer4_outputs(2502));
    layer5_outputs(1443) <= (layer4_outputs(4553)) and not (layer4_outputs(1515));
    layer5_outputs(1444) <= not((layer4_outputs(1801)) and (layer4_outputs(2793)));
    layer5_outputs(1445) <= (layer4_outputs(2852)) or (layer4_outputs(258));
    layer5_outputs(1446) <= not((layer4_outputs(3369)) xor (layer4_outputs(1913)));
    layer5_outputs(1447) <= (layer4_outputs(1928)) and (layer4_outputs(20));
    layer5_outputs(1448) <= not(layer4_outputs(2942));
    layer5_outputs(1449) <= layer4_outputs(878);
    layer5_outputs(1450) <= not((layer4_outputs(3261)) or (layer4_outputs(2552)));
    layer5_outputs(1451) <= not((layer4_outputs(2373)) and (layer4_outputs(2016)));
    layer5_outputs(1452) <= not((layer4_outputs(500)) and (layer4_outputs(4246)));
    layer5_outputs(1453) <= not(layer4_outputs(362));
    layer5_outputs(1454) <= not(layer4_outputs(4486)) or (layer4_outputs(421));
    layer5_outputs(1455) <= not((layer4_outputs(1077)) or (layer4_outputs(2538)));
    layer5_outputs(1456) <= layer4_outputs(2255);
    layer5_outputs(1457) <= layer4_outputs(1831);
    layer5_outputs(1458) <= not(layer4_outputs(1880));
    layer5_outputs(1459) <= layer4_outputs(3765);
    layer5_outputs(1460) <= not((layer4_outputs(2930)) or (layer4_outputs(4436)));
    layer5_outputs(1461) <= not(layer4_outputs(2342)) or (layer4_outputs(2169));
    layer5_outputs(1462) <= not(layer4_outputs(2572));
    layer5_outputs(1463) <= (layer4_outputs(1856)) and (layer4_outputs(3188));
    layer5_outputs(1464) <= (layer4_outputs(2252)) xor (layer4_outputs(4386));
    layer5_outputs(1465) <= layer4_outputs(4788);
    layer5_outputs(1466) <= not(layer4_outputs(1705));
    layer5_outputs(1467) <= (layer4_outputs(1246)) or (layer4_outputs(3917));
    layer5_outputs(1468) <= (layer4_outputs(2028)) and (layer4_outputs(3872));
    layer5_outputs(1469) <= (layer4_outputs(2528)) and not (layer4_outputs(3981));
    layer5_outputs(1470) <= (layer4_outputs(3395)) and (layer4_outputs(1770));
    layer5_outputs(1471) <= layer4_outputs(540);
    layer5_outputs(1472) <= not(layer4_outputs(1839));
    layer5_outputs(1473) <= '1';
    layer5_outputs(1474) <= '1';
    layer5_outputs(1475) <= not((layer4_outputs(4977)) and (layer4_outputs(53)));
    layer5_outputs(1476) <= not((layer4_outputs(2845)) xor (layer4_outputs(1015)));
    layer5_outputs(1477) <= not(layer4_outputs(2552)) or (layer4_outputs(644));
    layer5_outputs(1478) <= layer4_outputs(3324);
    layer5_outputs(1479) <= layer4_outputs(456);
    layer5_outputs(1480) <= not(layer4_outputs(4689));
    layer5_outputs(1481) <= (layer4_outputs(3324)) or (layer4_outputs(2432));
    layer5_outputs(1482) <= not(layer4_outputs(1833));
    layer5_outputs(1483) <= not((layer4_outputs(1397)) and (layer4_outputs(982)));
    layer5_outputs(1484) <= layer4_outputs(2174);
    layer5_outputs(1485) <= (layer4_outputs(3973)) xor (layer4_outputs(1694));
    layer5_outputs(1486) <= layer4_outputs(1712);
    layer5_outputs(1487) <= not(layer4_outputs(1477));
    layer5_outputs(1488) <= layer4_outputs(3119);
    layer5_outputs(1489) <= not(layer4_outputs(3130)) or (layer4_outputs(1093));
    layer5_outputs(1490) <= (layer4_outputs(2921)) and not (layer4_outputs(1169));
    layer5_outputs(1491) <= (layer4_outputs(5021)) and not (layer4_outputs(4277));
    layer5_outputs(1492) <= not(layer4_outputs(585));
    layer5_outputs(1493) <= not(layer4_outputs(1992));
    layer5_outputs(1494) <= (layer4_outputs(3072)) xor (layer4_outputs(3739));
    layer5_outputs(1495) <= (layer4_outputs(895)) or (layer4_outputs(437));
    layer5_outputs(1496) <= not((layer4_outputs(974)) or (layer4_outputs(2067)));
    layer5_outputs(1497) <= not((layer4_outputs(2997)) or (layer4_outputs(1439)));
    layer5_outputs(1498) <= not(layer4_outputs(4360));
    layer5_outputs(1499) <= not(layer4_outputs(3793)) or (layer4_outputs(4299));
    layer5_outputs(1500) <= (layer4_outputs(1858)) or (layer4_outputs(3500));
    layer5_outputs(1501) <= (layer4_outputs(1426)) and not (layer4_outputs(4050));
    layer5_outputs(1502) <= (layer4_outputs(2748)) and not (layer4_outputs(4854));
    layer5_outputs(1503) <= not(layer4_outputs(1230));
    layer5_outputs(1504) <= '1';
    layer5_outputs(1505) <= layer4_outputs(2812);
    layer5_outputs(1506) <= (layer4_outputs(3095)) xor (layer4_outputs(2414));
    layer5_outputs(1507) <= not(layer4_outputs(5037));
    layer5_outputs(1508) <= not(layer4_outputs(276));
    layer5_outputs(1509) <= not((layer4_outputs(1336)) or (layer4_outputs(3151)));
    layer5_outputs(1510) <= layer4_outputs(2928);
    layer5_outputs(1511) <= not(layer4_outputs(1708));
    layer5_outputs(1512) <= not(layer4_outputs(481)) or (layer4_outputs(588));
    layer5_outputs(1513) <= layer4_outputs(885);
    layer5_outputs(1514) <= not(layer4_outputs(2412));
    layer5_outputs(1515) <= (layer4_outputs(841)) or (layer4_outputs(2179));
    layer5_outputs(1516) <= not((layer4_outputs(2355)) and (layer4_outputs(738)));
    layer5_outputs(1517) <= not((layer4_outputs(3516)) and (layer4_outputs(2594)));
    layer5_outputs(1518) <= layer4_outputs(584);
    layer5_outputs(1519) <= not(layer4_outputs(5065));
    layer5_outputs(1520) <= not((layer4_outputs(328)) xor (layer4_outputs(4717)));
    layer5_outputs(1521) <= layer4_outputs(4811);
    layer5_outputs(1522) <= not(layer4_outputs(1818));
    layer5_outputs(1523) <= (layer4_outputs(167)) xor (layer4_outputs(3910));
    layer5_outputs(1524) <= layer4_outputs(17);
    layer5_outputs(1525) <= layer4_outputs(2174);
    layer5_outputs(1526) <= not(layer4_outputs(3104));
    layer5_outputs(1527) <= layer4_outputs(1419);
    layer5_outputs(1528) <= (layer4_outputs(3752)) or (layer4_outputs(2499));
    layer5_outputs(1529) <= not((layer4_outputs(2981)) or (layer4_outputs(3195)));
    layer5_outputs(1530) <= layer4_outputs(1613);
    layer5_outputs(1531) <= not((layer4_outputs(2581)) or (layer4_outputs(3643)));
    layer5_outputs(1532) <= not(layer4_outputs(978));
    layer5_outputs(1533) <= (layer4_outputs(2675)) or (layer4_outputs(1762));
    layer5_outputs(1534) <= layer4_outputs(5103);
    layer5_outputs(1535) <= not(layer4_outputs(2783));
    layer5_outputs(1536) <= (layer4_outputs(2437)) xor (layer4_outputs(3625));
    layer5_outputs(1537) <= (layer4_outputs(2058)) xor (layer4_outputs(2464));
    layer5_outputs(1538) <= not((layer4_outputs(4797)) xor (layer4_outputs(398)));
    layer5_outputs(1539) <= not((layer4_outputs(4792)) xor (layer4_outputs(3942)));
    layer5_outputs(1540) <= not(layer4_outputs(861));
    layer5_outputs(1541) <= not((layer4_outputs(3266)) and (layer4_outputs(1424)));
    layer5_outputs(1542) <= (layer4_outputs(327)) and (layer4_outputs(1616));
    layer5_outputs(1543) <= not((layer4_outputs(3211)) xor (layer4_outputs(4253)));
    layer5_outputs(1544) <= (layer4_outputs(2484)) and (layer4_outputs(836));
    layer5_outputs(1545) <= layer4_outputs(3165);
    layer5_outputs(1546) <= (layer4_outputs(3193)) and not (layer4_outputs(3260));
    layer5_outputs(1547) <= (layer4_outputs(4738)) or (layer4_outputs(2023));
    layer5_outputs(1548) <= not(layer4_outputs(3914));
    layer5_outputs(1549) <= not((layer4_outputs(4904)) and (layer4_outputs(3147)));
    layer5_outputs(1550) <= not((layer4_outputs(2893)) xor (layer4_outputs(3359)));
    layer5_outputs(1551) <= '1';
    layer5_outputs(1552) <= not(layer4_outputs(2341));
    layer5_outputs(1553) <= (layer4_outputs(4484)) and not (layer4_outputs(1345));
    layer5_outputs(1554) <= '0';
    layer5_outputs(1555) <= not(layer4_outputs(3478));
    layer5_outputs(1556) <= '1';
    layer5_outputs(1557) <= not(layer4_outputs(4626));
    layer5_outputs(1558) <= layer4_outputs(4682);
    layer5_outputs(1559) <= not(layer4_outputs(5112));
    layer5_outputs(1560) <= not(layer4_outputs(805));
    layer5_outputs(1561) <= not(layer4_outputs(1460));
    layer5_outputs(1562) <= not(layer4_outputs(702));
    layer5_outputs(1563) <= (layer4_outputs(2028)) xor (layer4_outputs(4157));
    layer5_outputs(1564) <= not((layer4_outputs(499)) and (layer4_outputs(2337)));
    layer5_outputs(1565) <= '0';
    layer5_outputs(1566) <= layer4_outputs(4982);
    layer5_outputs(1567) <= not((layer4_outputs(1768)) xor (layer4_outputs(1313)));
    layer5_outputs(1568) <= not(layer4_outputs(3597)) or (layer4_outputs(2124));
    layer5_outputs(1569) <= layer4_outputs(2807);
    layer5_outputs(1570) <= not(layer4_outputs(735));
    layer5_outputs(1571) <= layer4_outputs(1287);
    layer5_outputs(1572) <= not((layer4_outputs(3876)) or (layer4_outputs(1955)));
    layer5_outputs(1573) <= (layer4_outputs(5050)) or (layer4_outputs(2279));
    layer5_outputs(1574) <= not(layer4_outputs(1363)) or (layer4_outputs(2936));
    layer5_outputs(1575) <= not((layer4_outputs(1171)) or (layer4_outputs(4350)));
    layer5_outputs(1576) <= '1';
    layer5_outputs(1577) <= '0';
    layer5_outputs(1578) <= not(layer4_outputs(3596));
    layer5_outputs(1579) <= not(layer4_outputs(931));
    layer5_outputs(1580) <= layer4_outputs(4088);
    layer5_outputs(1581) <= not(layer4_outputs(988)) or (layer4_outputs(1749));
    layer5_outputs(1582) <= layer4_outputs(1945);
    layer5_outputs(1583) <= layer4_outputs(3005);
    layer5_outputs(1584) <= layer4_outputs(1115);
    layer5_outputs(1585) <= (layer4_outputs(370)) and not (layer4_outputs(3796));
    layer5_outputs(1586) <= layer4_outputs(3814);
    layer5_outputs(1587) <= layer4_outputs(4326);
    layer5_outputs(1588) <= (layer4_outputs(1615)) or (layer4_outputs(388));
    layer5_outputs(1589) <= not(layer4_outputs(4343));
    layer5_outputs(1590) <= not(layer4_outputs(4345));
    layer5_outputs(1591) <= '0';
    layer5_outputs(1592) <= (layer4_outputs(264)) and (layer4_outputs(2059));
    layer5_outputs(1593) <= (layer4_outputs(1421)) or (layer4_outputs(530));
    layer5_outputs(1594) <= '0';
    layer5_outputs(1595) <= (layer4_outputs(1768)) and not (layer4_outputs(1352));
    layer5_outputs(1596) <= layer4_outputs(3648);
    layer5_outputs(1597) <= layer4_outputs(1095);
    layer5_outputs(1598) <= not((layer4_outputs(195)) or (layer4_outputs(4849)));
    layer5_outputs(1599) <= '1';
    layer5_outputs(1600) <= not(layer4_outputs(3288));
    layer5_outputs(1601) <= not(layer4_outputs(441));
    layer5_outputs(1602) <= layer4_outputs(4724);
    layer5_outputs(1603) <= (layer4_outputs(1969)) xor (layer4_outputs(3451));
    layer5_outputs(1604) <= not((layer4_outputs(1967)) or (layer4_outputs(3737)));
    layer5_outputs(1605) <= not(layer4_outputs(1181)) or (layer4_outputs(1820));
    layer5_outputs(1606) <= not(layer4_outputs(3750));
    layer5_outputs(1607) <= layer4_outputs(3889);
    layer5_outputs(1608) <= layer4_outputs(1976);
    layer5_outputs(1609) <= not(layer4_outputs(4283));
    layer5_outputs(1610) <= layer4_outputs(2785);
    layer5_outputs(1611) <= not((layer4_outputs(797)) xor (layer4_outputs(3819)));
    layer5_outputs(1612) <= not(layer4_outputs(2991));
    layer5_outputs(1613) <= (layer4_outputs(3177)) and not (layer4_outputs(2592));
    layer5_outputs(1614) <= (layer4_outputs(1714)) and (layer4_outputs(5014));
    layer5_outputs(1615) <= not((layer4_outputs(1366)) or (layer4_outputs(3696)));
    layer5_outputs(1616) <= layer4_outputs(1528);
    layer5_outputs(1617) <= layer4_outputs(2147);
    layer5_outputs(1618) <= (layer4_outputs(1262)) and (layer4_outputs(1666));
    layer5_outputs(1619) <= layer4_outputs(3100);
    layer5_outputs(1620) <= layer4_outputs(2970);
    layer5_outputs(1621) <= (layer4_outputs(3059)) xor (layer4_outputs(721));
    layer5_outputs(1622) <= layer4_outputs(4385);
    layer5_outputs(1623) <= '0';
    layer5_outputs(1624) <= not(layer4_outputs(5080));
    layer5_outputs(1625) <= not(layer4_outputs(2656)) or (layer4_outputs(2940));
    layer5_outputs(1626) <= not((layer4_outputs(4378)) or (layer4_outputs(5042)));
    layer5_outputs(1627) <= not(layer4_outputs(633));
    layer5_outputs(1628) <= (layer4_outputs(674)) and (layer4_outputs(4866));
    layer5_outputs(1629) <= (layer4_outputs(1130)) and not (layer4_outputs(291));
    layer5_outputs(1630) <= not((layer4_outputs(3698)) or (layer4_outputs(286)));
    layer5_outputs(1631) <= (layer4_outputs(3822)) and (layer4_outputs(4279));
    layer5_outputs(1632) <= (layer4_outputs(1862)) and not (layer4_outputs(4188));
    layer5_outputs(1633) <= not(layer4_outputs(1871));
    layer5_outputs(1634) <= not(layer4_outputs(4749));
    layer5_outputs(1635) <= not(layer4_outputs(5012));
    layer5_outputs(1636) <= not(layer4_outputs(3785));
    layer5_outputs(1637) <= layer4_outputs(3021);
    layer5_outputs(1638) <= not((layer4_outputs(2812)) xor (layer4_outputs(2929)));
    layer5_outputs(1639) <= not(layer4_outputs(1507)) or (layer4_outputs(4231));
    layer5_outputs(1640) <= not(layer4_outputs(1247)) or (layer4_outputs(43));
    layer5_outputs(1641) <= not((layer4_outputs(4326)) xor (layer4_outputs(316)));
    layer5_outputs(1642) <= not(layer4_outputs(4776)) or (layer4_outputs(1024));
    layer5_outputs(1643) <= not(layer4_outputs(597));
    layer5_outputs(1644) <= (layer4_outputs(40)) xor (layer4_outputs(961));
    layer5_outputs(1645) <= (layer4_outputs(1263)) and not (layer4_outputs(2090));
    layer5_outputs(1646) <= not(layer4_outputs(19));
    layer5_outputs(1647) <= not(layer4_outputs(2843));
    layer5_outputs(1648) <= (layer4_outputs(517)) or (layer4_outputs(3799));
    layer5_outputs(1649) <= (layer4_outputs(3751)) and not (layer4_outputs(4073));
    layer5_outputs(1650) <= not(layer4_outputs(1599)) or (layer4_outputs(4756));
    layer5_outputs(1651) <= not(layer4_outputs(4510));
    layer5_outputs(1652) <= layer4_outputs(1387);
    layer5_outputs(1653) <= (layer4_outputs(1398)) xor (layer4_outputs(3076));
    layer5_outputs(1654) <= not(layer4_outputs(2676));
    layer5_outputs(1655) <= not((layer4_outputs(4185)) and (layer4_outputs(2345)));
    layer5_outputs(1656) <= '1';
    layer5_outputs(1657) <= layer4_outputs(4002);
    layer5_outputs(1658) <= not(layer4_outputs(1150));
    layer5_outputs(1659) <= '1';
    layer5_outputs(1660) <= '0';
    layer5_outputs(1661) <= not(layer4_outputs(3567)) or (layer4_outputs(2279));
    layer5_outputs(1662) <= not(layer4_outputs(4438));
    layer5_outputs(1663) <= layer4_outputs(1922);
    layer5_outputs(1664) <= not(layer4_outputs(2488)) or (layer4_outputs(1509));
    layer5_outputs(1665) <= layer4_outputs(1164);
    layer5_outputs(1666) <= not(layer4_outputs(591));
    layer5_outputs(1667) <= (layer4_outputs(3491)) and not (layer4_outputs(4835));
    layer5_outputs(1668) <= not(layer4_outputs(3781));
    layer5_outputs(1669) <= layer4_outputs(4129);
    layer5_outputs(1670) <= not(layer4_outputs(765)) or (layer4_outputs(1622));
    layer5_outputs(1671) <= layer4_outputs(5032);
    layer5_outputs(1672) <= layer4_outputs(1632);
    layer5_outputs(1673) <= (layer4_outputs(4027)) and (layer4_outputs(271));
    layer5_outputs(1674) <= layer4_outputs(471);
    layer5_outputs(1675) <= layer4_outputs(2346);
    layer5_outputs(1676) <= (layer4_outputs(3948)) and (layer4_outputs(1789));
    layer5_outputs(1677) <= (layer4_outputs(257)) or (layer4_outputs(3443));
    layer5_outputs(1678) <= layer4_outputs(1099);
    layer5_outputs(1679) <= layer4_outputs(3923);
    layer5_outputs(1680) <= (layer4_outputs(820)) xor (layer4_outputs(2412));
    layer5_outputs(1681) <= not(layer4_outputs(4201)) or (layer4_outputs(1931));
    layer5_outputs(1682) <= layer4_outputs(2724);
    layer5_outputs(1683) <= not(layer4_outputs(2071)) or (layer4_outputs(993));
    layer5_outputs(1684) <= not(layer4_outputs(3271));
    layer5_outputs(1685) <= layer4_outputs(1745);
    layer5_outputs(1686) <= not(layer4_outputs(3955));
    layer5_outputs(1687) <= not((layer4_outputs(2322)) or (layer4_outputs(4373)));
    layer5_outputs(1688) <= not(layer4_outputs(3252)) or (layer4_outputs(2828));
    layer5_outputs(1689) <= not((layer4_outputs(1527)) xor (layer4_outputs(2255)));
    layer5_outputs(1690) <= not((layer4_outputs(2384)) or (layer4_outputs(1216)));
    layer5_outputs(1691) <= not(layer4_outputs(3638));
    layer5_outputs(1692) <= not((layer4_outputs(501)) or (layer4_outputs(4363)));
    layer5_outputs(1693) <= (layer4_outputs(3550)) and (layer4_outputs(3959));
    layer5_outputs(1694) <= (layer4_outputs(419)) and (layer4_outputs(3028));
    layer5_outputs(1695) <= not(layer4_outputs(3247)) or (layer4_outputs(108));
    layer5_outputs(1696) <= not(layer4_outputs(1149)) or (layer4_outputs(506));
    layer5_outputs(1697) <= (layer4_outputs(4499)) and not (layer4_outputs(4478));
    layer5_outputs(1698) <= not(layer4_outputs(617));
    layer5_outputs(1699) <= not(layer4_outputs(1158));
    layer5_outputs(1700) <= not((layer4_outputs(4337)) or (layer4_outputs(3049)));
    layer5_outputs(1701) <= layer4_outputs(2845);
    layer5_outputs(1702) <= not(layer4_outputs(4898));
    layer5_outputs(1703) <= layer4_outputs(1132);
    layer5_outputs(1704) <= not(layer4_outputs(2150));
    layer5_outputs(1705) <= (layer4_outputs(2299)) xor (layer4_outputs(1844));
    layer5_outputs(1706) <= not(layer4_outputs(3440)) or (layer4_outputs(2390));
    layer5_outputs(1707) <= not((layer4_outputs(4850)) and (layer4_outputs(2365)));
    layer5_outputs(1708) <= not(layer4_outputs(4362)) or (layer4_outputs(2004));
    layer5_outputs(1709) <= '1';
    layer5_outputs(1710) <= layer4_outputs(1663);
    layer5_outputs(1711) <= (layer4_outputs(2980)) xor (layer4_outputs(1964));
    layer5_outputs(1712) <= not(layer4_outputs(1314));
    layer5_outputs(1713) <= layer4_outputs(2268);
    layer5_outputs(1714) <= layer4_outputs(4745);
    layer5_outputs(1715) <= (layer4_outputs(319)) and (layer4_outputs(2289));
    layer5_outputs(1716) <= '1';
    layer5_outputs(1717) <= '0';
    layer5_outputs(1718) <= layer4_outputs(1887);
    layer5_outputs(1719) <= '0';
    layer5_outputs(1720) <= not((layer4_outputs(31)) xor (layer4_outputs(3302)));
    layer5_outputs(1721) <= '0';
    layer5_outputs(1722) <= layer4_outputs(637);
    layer5_outputs(1723) <= not(layer4_outputs(1930));
    layer5_outputs(1724) <= not((layer4_outputs(1064)) and (layer4_outputs(3146)));
    layer5_outputs(1725) <= layer4_outputs(4462);
    layer5_outputs(1726) <= not((layer4_outputs(4116)) or (layer4_outputs(3659)));
    layer5_outputs(1727) <= not(layer4_outputs(368));
    layer5_outputs(1728) <= not(layer4_outputs(1441));
    layer5_outputs(1729) <= not(layer4_outputs(2579));
    layer5_outputs(1730) <= '0';
    layer5_outputs(1731) <= layer4_outputs(459);
    layer5_outputs(1732) <= not((layer4_outputs(4228)) and (layer4_outputs(3222)));
    layer5_outputs(1733) <= layer4_outputs(1220);
    layer5_outputs(1734) <= (layer4_outputs(2509)) and not (layer4_outputs(625));
    layer5_outputs(1735) <= not((layer4_outputs(2447)) xor (layer4_outputs(1567)));
    layer5_outputs(1736) <= layer4_outputs(1908);
    layer5_outputs(1737) <= not(layer4_outputs(4170));
    layer5_outputs(1738) <= not(layer4_outputs(2210));
    layer5_outputs(1739) <= (layer4_outputs(141)) and not (layer4_outputs(2520));
    layer5_outputs(1740) <= (layer4_outputs(2137)) and not (layer4_outputs(1622));
    layer5_outputs(1741) <= layer4_outputs(4630);
    layer5_outputs(1742) <= (layer4_outputs(1733)) and not (layer4_outputs(4422));
    layer5_outputs(1743) <= layer4_outputs(3459);
    layer5_outputs(1744) <= not(layer4_outputs(4199));
    layer5_outputs(1745) <= layer4_outputs(1439);
    layer5_outputs(1746) <= layer4_outputs(1459);
    layer5_outputs(1747) <= layer4_outputs(4361);
    layer5_outputs(1748) <= (layer4_outputs(2140)) and not (layer4_outputs(4253));
    layer5_outputs(1749) <= (layer4_outputs(1977)) or (layer4_outputs(1846));
    layer5_outputs(1750) <= layer4_outputs(1659);
    layer5_outputs(1751) <= not(layer4_outputs(1379)) or (layer4_outputs(2002));
    layer5_outputs(1752) <= (layer4_outputs(1284)) and not (layer4_outputs(2990));
    layer5_outputs(1753) <= not(layer4_outputs(1803));
    layer5_outputs(1754) <= (layer4_outputs(2665)) or (layer4_outputs(801));
    layer5_outputs(1755) <= layer4_outputs(709);
    layer5_outputs(1756) <= (layer4_outputs(4258)) xor (layer4_outputs(4330));
    layer5_outputs(1757) <= layer4_outputs(418);
    layer5_outputs(1758) <= layer4_outputs(3003);
    layer5_outputs(1759) <= not(layer4_outputs(4176));
    layer5_outputs(1760) <= layer4_outputs(1752);
    layer5_outputs(1761) <= not(layer4_outputs(986));
    layer5_outputs(1762) <= (layer4_outputs(2711)) or (layer4_outputs(1678));
    layer5_outputs(1763) <= (layer4_outputs(1128)) and not (layer4_outputs(1486));
    layer5_outputs(1764) <= '0';
    layer5_outputs(1765) <= not(layer4_outputs(4132));
    layer5_outputs(1766) <= (layer4_outputs(905)) and (layer4_outputs(1948));
    layer5_outputs(1767) <= not(layer4_outputs(1612)) or (layer4_outputs(1031));
    layer5_outputs(1768) <= (layer4_outputs(4942)) xor (layer4_outputs(2586));
    layer5_outputs(1769) <= (layer4_outputs(481)) and not (layer4_outputs(3207));
    layer5_outputs(1770) <= not(layer4_outputs(4197));
    layer5_outputs(1771) <= not(layer4_outputs(2249)) or (layer4_outputs(5002));
    layer5_outputs(1772) <= (layer4_outputs(2299)) and not (layer4_outputs(1074));
    layer5_outputs(1773) <= not(layer4_outputs(169));
    layer5_outputs(1774) <= not(layer4_outputs(3975));
    layer5_outputs(1775) <= layer4_outputs(4559);
    layer5_outputs(1776) <= not(layer4_outputs(3469));
    layer5_outputs(1777) <= (layer4_outputs(2145)) xor (layer4_outputs(3542));
    layer5_outputs(1778) <= layer4_outputs(396);
    layer5_outputs(1779) <= layer4_outputs(910);
    layer5_outputs(1780) <= (layer4_outputs(490)) or (layer4_outputs(3620));
    layer5_outputs(1781) <= layer4_outputs(1159);
    layer5_outputs(1782) <= not((layer4_outputs(785)) or (layer4_outputs(3717)));
    layer5_outputs(1783) <= layer4_outputs(4742);
    layer5_outputs(1784) <= not(layer4_outputs(1917)) or (layer4_outputs(4245));
    layer5_outputs(1785) <= layer4_outputs(5003);
    layer5_outputs(1786) <= not((layer4_outputs(3286)) xor (layer4_outputs(2540)));
    layer5_outputs(1787) <= (layer4_outputs(3613)) xor (layer4_outputs(4924));
    layer5_outputs(1788) <= not((layer4_outputs(4708)) and (layer4_outputs(4860)));
    layer5_outputs(1789) <= layer4_outputs(2495);
    layer5_outputs(1790) <= '1';
    layer5_outputs(1791) <= layer4_outputs(2631);
    layer5_outputs(1792) <= not(layer4_outputs(2431));
    layer5_outputs(1793) <= layer4_outputs(3988);
    layer5_outputs(1794) <= not((layer4_outputs(135)) xor (layer4_outputs(275)));
    layer5_outputs(1795) <= '1';
    layer5_outputs(1796) <= (layer4_outputs(1595)) or (layer4_outputs(240));
    layer5_outputs(1797) <= not(layer4_outputs(482)) or (layer4_outputs(1895));
    layer5_outputs(1798) <= '0';
    layer5_outputs(1799) <= (layer4_outputs(1840)) or (layer4_outputs(1253));
    layer5_outputs(1800) <= not(layer4_outputs(2922)) or (layer4_outputs(1411));
    layer5_outputs(1801) <= not(layer4_outputs(4632));
    layer5_outputs(1802) <= not(layer4_outputs(622));
    layer5_outputs(1803) <= layer4_outputs(1921);
    layer5_outputs(1804) <= not(layer4_outputs(2161)) or (layer4_outputs(4936));
    layer5_outputs(1805) <= (layer4_outputs(2234)) and not (layer4_outputs(3214));
    layer5_outputs(1806) <= layer4_outputs(3850);
    layer5_outputs(1807) <= not(layer4_outputs(3846)) or (layer4_outputs(2395));
    layer5_outputs(1808) <= (layer4_outputs(3076)) and not (layer4_outputs(1704));
    layer5_outputs(1809) <= (layer4_outputs(3806)) and (layer4_outputs(3253));
    layer5_outputs(1810) <= not((layer4_outputs(770)) and (layer4_outputs(2918)));
    layer5_outputs(1811) <= layer4_outputs(1751);
    layer5_outputs(1812) <= not(layer4_outputs(3843));
    layer5_outputs(1813) <= not(layer4_outputs(3366)) or (layer4_outputs(4641));
    layer5_outputs(1814) <= not(layer4_outputs(4212));
    layer5_outputs(1815) <= not(layer4_outputs(1332));
    layer5_outputs(1816) <= not(layer4_outputs(3572));
    layer5_outputs(1817) <= (layer4_outputs(1743)) or (layer4_outputs(784));
    layer5_outputs(1818) <= not(layer4_outputs(3663));
    layer5_outputs(1819) <= not(layer4_outputs(3179));
    layer5_outputs(1820) <= not((layer4_outputs(692)) and (layer4_outputs(1554)));
    layer5_outputs(1821) <= layer4_outputs(4629);
    layer5_outputs(1822) <= not(layer4_outputs(4637)) or (layer4_outputs(1289));
    layer5_outputs(1823) <= (layer4_outputs(661)) and not (layer4_outputs(2614));
    layer5_outputs(1824) <= (layer4_outputs(3042)) xor (layer4_outputs(4957));
    layer5_outputs(1825) <= not(layer4_outputs(3378)) or (layer4_outputs(1997));
    layer5_outputs(1826) <= layer4_outputs(3619);
    layer5_outputs(1827) <= not(layer4_outputs(1729));
    layer5_outputs(1828) <= layer4_outputs(2010);
    layer5_outputs(1829) <= not((layer4_outputs(1310)) or (layer4_outputs(1528)));
    layer5_outputs(1830) <= layer4_outputs(2805);
    layer5_outputs(1831) <= not(layer4_outputs(3528));
    layer5_outputs(1832) <= (layer4_outputs(2926)) and not (layer4_outputs(2008));
    layer5_outputs(1833) <= layer4_outputs(2513);
    layer5_outputs(1834) <= (layer4_outputs(3672)) or (layer4_outputs(4809));
    layer5_outputs(1835) <= not((layer4_outputs(2768)) or (layer4_outputs(4388)));
    layer5_outputs(1836) <= '0';
    layer5_outputs(1837) <= (layer4_outputs(3982)) and not (layer4_outputs(2426));
    layer5_outputs(1838) <= (layer4_outputs(1019)) xor (layer4_outputs(3941));
    layer5_outputs(1839) <= layer4_outputs(3190);
    layer5_outputs(1840) <= '0';
    layer5_outputs(1841) <= (layer4_outputs(3526)) xor (layer4_outputs(3527));
    layer5_outputs(1842) <= layer4_outputs(3454);
    layer5_outputs(1843) <= not(layer4_outputs(1382));
    layer5_outputs(1844) <= (layer4_outputs(2882)) and not (layer4_outputs(2758));
    layer5_outputs(1845) <= (layer4_outputs(4991)) and not (layer4_outputs(1868));
    layer5_outputs(1846) <= layer4_outputs(4316);
    layer5_outputs(1847) <= layer4_outputs(4788);
    layer5_outputs(1848) <= layer4_outputs(2825);
    layer5_outputs(1849) <= not((layer4_outputs(2857)) and (layer4_outputs(1702)));
    layer5_outputs(1850) <= '0';
    layer5_outputs(1851) <= (layer4_outputs(3787)) and not (layer4_outputs(4482));
    layer5_outputs(1852) <= not(layer4_outputs(2846));
    layer5_outputs(1853) <= not((layer4_outputs(3448)) or (layer4_outputs(4177)));
    layer5_outputs(1854) <= layer4_outputs(2587);
    layer5_outputs(1855) <= not(layer4_outputs(2818));
    layer5_outputs(1856) <= not(layer4_outputs(2036));
    layer5_outputs(1857) <= (layer4_outputs(514)) and (layer4_outputs(2636));
    layer5_outputs(1858) <= '0';
    layer5_outputs(1859) <= '1';
    layer5_outputs(1860) <= layer4_outputs(5091);
    layer5_outputs(1861) <= not(layer4_outputs(1096));
    layer5_outputs(1862) <= not(layer4_outputs(4885));
    layer5_outputs(1863) <= not(layer4_outputs(3810));
    layer5_outputs(1864) <= (layer4_outputs(4394)) or (layer4_outputs(5068));
    layer5_outputs(1865) <= (layer4_outputs(2523)) or (layer4_outputs(4271));
    layer5_outputs(1866) <= layer4_outputs(4437);
    layer5_outputs(1867) <= not((layer4_outputs(1096)) xor (layer4_outputs(862)));
    layer5_outputs(1868) <= not((layer4_outputs(3390)) or (layer4_outputs(3967)));
    layer5_outputs(1869) <= not(layer4_outputs(1972));
    layer5_outputs(1870) <= not(layer4_outputs(2485));
    layer5_outputs(1871) <= not(layer4_outputs(1299));
    layer5_outputs(1872) <= layer4_outputs(2833);
    layer5_outputs(1873) <= not(layer4_outputs(1548));
    layer5_outputs(1874) <= not(layer4_outputs(4363));
    layer5_outputs(1875) <= (layer4_outputs(2444)) and (layer4_outputs(2844));
    layer5_outputs(1876) <= not(layer4_outputs(3591));
    layer5_outputs(1877) <= not(layer4_outputs(121)) or (layer4_outputs(3219));
    layer5_outputs(1878) <= layer4_outputs(2069);
    layer5_outputs(1879) <= layer4_outputs(2741);
    layer5_outputs(1880) <= not(layer4_outputs(2105));
    layer5_outputs(1881) <= (layer4_outputs(1253)) and not (layer4_outputs(3297));
    layer5_outputs(1882) <= not(layer4_outputs(836));
    layer5_outputs(1883) <= not(layer4_outputs(4919)) or (layer4_outputs(3798));
    layer5_outputs(1884) <= layer4_outputs(1564);
    layer5_outputs(1885) <= layer4_outputs(1359);
    layer5_outputs(1886) <= layer4_outputs(4862);
    layer5_outputs(1887) <= layer4_outputs(2422);
    layer5_outputs(1888) <= (layer4_outputs(278)) and (layer4_outputs(115));
    layer5_outputs(1889) <= not((layer4_outputs(200)) xor (layer4_outputs(2359)));
    layer5_outputs(1890) <= (layer4_outputs(3446)) or (layer4_outputs(2533));
    layer5_outputs(1891) <= not(layer4_outputs(3650));
    layer5_outputs(1892) <= not((layer4_outputs(3433)) xor (layer4_outputs(3445)));
    layer5_outputs(1893) <= (layer4_outputs(4909)) and not (layer4_outputs(393));
    layer5_outputs(1894) <= layer4_outputs(4570);
    layer5_outputs(1895) <= not(layer4_outputs(1213));
    layer5_outputs(1896) <= not(layer4_outputs(891));
    layer5_outputs(1897) <= not(layer4_outputs(1322));
    layer5_outputs(1898) <= not(layer4_outputs(4360)) or (layer4_outputs(4992));
    layer5_outputs(1899) <= (layer4_outputs(1658)) xor (layer4_outputs(12));
    layer5_outputs(1900) <= (layer4_outputs(4041)) xor (layer4_outputs(2948));
    layer5_outputs(1901) <= layer4_outputs(1849);
    layer5_outputs(1902) <= not(layer4_outputs(2141));
    layer5_outputs(1903) <= not(layer4_outputs(3687));
    layer5_outputs(1904) <= not((layer4_outputs(2855)) or (layer4_outputs(4585)));
    layer5_outputs(1905) <= not(layer4_outputs(1765));
    layer5_outputs(1906) <= layer4_outputs(728);
    layer5_outputs(1907) <= (layer4_outputs(2883)) or (layer4_outputs(513));
    layer5_outputs(1908) <= not((layer4_outputs(3685)) or (layer4_outputs(648)));
    layer5_outputs(1909) <= (layer4_outputs(2425)) and (layer4_outputs(2959));
    layer5_outputs(1910) <= layer4_outputs(4328);
    layer5_outputs(1911) <= layer4_outputs(4934);
    layer5_outputs(1912) <= layer4_outputs(5019);
    layer5_outputs(1913) <= (layer4_outputs(4062)) and not (layer4_outputs(4650));
    layer5_outputs(1914) <= not(layer4_outputs(523)) or (layer4_outputs(1339));
    layer5_outputs(1915) <= (layer4_outputs(401)) xor (layer4_outputs(5054));
    layer5_outputs(1916) <= not(layer4_outputs(1571)) or (layer4_outputs(4840));
    layer5_outputs(1917) <= layer4_outputs(1761);
    layer5_outputs(1918) <= layer4_outputs(3934);
    layer5_outputs(1919) <= not(layer4_outputs(4390));
    layer5_outputs(1920) <= '1';
    layer5_outputs(1921) <= not((layer4_outputs(2424)) or (layer4_outputs(3865)));
    layer5_outputs(1922) <= not(layer4_outputs(3798));
    layer5_outputs(1923) <= not(layer4_outputs(3962));
    layer5_outputs(1924) <= not(layer4_outputs(1531)) or (layer4_outputs(4567));
    layer5_outputs(1925) <= layer4_outputs(1957);
    layer5_outputs(1926) <= not(layer4_outputs(3333));
    layer5_outputs(1927) <= (layer4_outputs(2929)) or (layer4_outputs(34));
    layer5_outputs(1928) <= not(layer4_outputs(1354));
    layer5_outputs(1929) <= layer4_outputs(2089);
    layer5_outputs(1930) <= not(layer4_outputs(4217));
    layer5_outputs(1931) <= (layer4_outputs(1299)) and (layer4_outputs(4365));
    layer5_outputs(1932) <= not(layer4_outputs(4029)) or (layer4_outputs(1859));
    layer5_outputs(1933) <= '1';
    layer5_outputs(1934) <= layer4_outputs(1188);
    layer5_outputs(1935) <= layer4_outputs(4719);
    layer5_outputs(1936) <= not((layer4_outputs(2607)) xor (layer4_outputs(1866)));
    layer5_outputs(1937) <= not((layer4_outputs(3268)) and (layer4_outputs(1572)));
    layer5_outputs(1938) <= (layer4_outputs(1936)) or (layer4_outputs(2422));
    layer5_outputs(1939) <= not(layer4_outputs(3037));
    layer5_outputs(1940) <= not(layer4_outputs(3744));
    layer5_outputs(1941) <= (layer4_outputs(1641)) and not (layer4_outputs(2914));
    layer5_outputs(1942) <= (layer4_outputs(312)) xor (layer4_outputs(4354));
    layer5_outputs(1943) <= not(layer4_outputs(1676));
    layer5_outputs(1944) <= (layer4_outputs(5070)) xor (layer4_outputs(3489));
    layer5_outputs(1945) <= not((layer4_outputs(3314)) or (layer4_outputs(366)));
    layer5_outputs(1946) <= layer4_outputs(1973);
    layer5_outputs(1947) <= (layer4_outputs(100)) and (layer4_outputs(1146));
    layer5_outputs(1948) <= (layer4_outputs(4810)) and not (layer4_outputs(3616));
    layer5_outputs(1949) <= layer4_outputs(1998);
    layer5_outputs(1950) <= not(layer4_outputs(4531));
    layer5_outputs(1951) <= not((layer4_outputs(3432)) and (layer4_outputs(302)));
    layer5_outputs(1952) <= layer4_outputs(1523);
    layer5_outputs(1953) <= (layer4_outputs(1815)) or (layer4_outputs(4204));
    layer5_outputs(1954) <= layer4_outputs(4641);
    layer5_outputs(1955) <= layer4_outputs(3397);
    layer5_outputs(1956) <= (layer4_outputs(3031)) xor (layer4_outputs(1226));
    layer5_outputs(1957) <= not(layer4_outputs(308)) or (layer4_outputs(1037));
    layer5_outputs(1958) <= not(layer4_outputs(3304));
    layer5_outputs(1959) <= not((layer4_outputs(183)) or (layer4_outputs(3136)));
    layer5_outputs(1960) <= (layer4_outputs(1959)) and not (layer4_outputs(1207));
    layer5_outputs(1961) <= not((layer4_outputs(2286)) and (layer4_outputs(3888)));
    layer5_outputs(1962) <= not((layer4_outputs(2326)) xor (layer4_outputs(847)));
    layer5_outputs(1963) <= not(layer4_outputs(2370));
    layer5_outputs(1964) <= '0';
    layer5_outputs(1965) <= '0';
    layer5_outputs(1966) <= '0';
    layer5_outputs(1967) <= '1';
    layer5_outputs(1968) <= not(layer4_outputs(3760));
    layer5_outputs(1969) <= layer4_outputs(607);
    layer5_outputs(1970) <= not(layer4_outputs(2834));
    layer5_outputs(1971) <= not(layer4_outputs(1500)) or (layer4_outputs(797));
    layer5_outputs(1972) <= not((layer4_outputs(3455)) or (layer4_outputs(3201)));
    layer5_outputs(1973) <= not(layer4_outputs(4767));
    layer5_outputs(1974) <= (layer4_outputs(3768)) and not (layer4_outputs(3944));
    layer5_outputs(1975) <= not(layer4_outputs(1356)) or (layer4_outputs(2109));
    layer5_outputs(1976) <= not(layer4_outputs(1612));
    layer5_outputs(1977) <= '0';
    layer5_outputs(1978) <= not((layer4_outputs(182)) xor (layer4_outputs(1974)));
    layer5_outputs(1979) <= (layer4_outputs(4480)) and not (layer4_outputs(2515));
    layer5_outputs(1980) <= '0';
    layer5_outputs(1981) <= not(layer4_outputs(804));
    layer5_outputs(1982) <= not(layer4_outputs(1174)) or (layer4_outputs(4057));
    layer5_outputs(1983) <= not(layer4_outputs(1512));
    layer5_outputs(1984) <= not(layer4_outputs(5114));
    layer5_outputs(1985) <= not(layer4_outputs(4351));
    layer5_outputs(1986) <= layer4_outputs(1552);
    layer5_outputs(1987) <= not(layer4_outputs(259));
    layer5_outputs(1988) <= '0';
    layer5_outputs(1989) <= not(layer4_outputs(3654));
    layer5_outputs(1990) <= layer4_outputs(3668);
    layer5_outputs(1991) <= not((layer4_outputs(4248)) xor (layer4_outputs(1212)));
    layer5_outputs(1992) <= (layer4_outputs(4846)) and not (layer4_outputs(195));
    layer5_outputs(1993) <= not(layer4_outputs(2078));
    layer5_outputs(1994) <= layer4_outputs(5038);
    layer5_outputs(1995) <= not(layer4_outputs(4613));
    layer5_outputs(1996) <= not(layer4_outputs(3677));
    layer5_outputs(1997) <= not(layer4_outputs(1110)) or (layer4_outputs(1294));
    layer5_outputs(1998) <= not(layer4_outputs(461));
    layer5_outputs(1999) <= not(layer4_outputs(874));
    layer5_outputs(2000) <= not(layer4_outputs(3721)) or (layer4_outputs(318));
    layer5_outputs(2001) <= layer4_outputs(2955);
    layer5_outputs(2002) <= (layer4_outputs(1335)) and (layer4_outputs(527));
    layer5_outputs(2003) <= layer4_outputs(485);
    layer5_outputs(2004) <= not(layer4_outputs(3060));
    layer5_outputs(2005) <= not(layer4_outputs(175));
    layer5_outputs(2006) <= (layer4_outputs(1360)) and not (layer4_outputs(2095));
    layer5_outputs(2007) <= layer4_outputs(2687);
    layer5_outputs(2008) <= (layer4_outputs(1429)) or (layer4_outputs(5001));
    layer5_outputs(2009) <= layer4_outputs(382);
    layer5_outputs(2010) <= not(layer4_outputs(1769));
    layer5_outputs(2011) <= layer4_outputs(1133);
    layer5_outputs(2012) <= not(layer4_outputs(4699));
    layer5_outputs(2013) <= not(layer4_outputs(845)) or (layer4_outputs(3357));
    layer5_outputs(2014) <= not(layer4_outputs(2281));
    layer5_outputs(2015) <= (layer4_outputs(4327)) and not (layer4_outputs(4048));
    layer5_outputs(2016) <= not(layer4_outputs(4042)) or (layer4_outputs(2107));
    layer5_outputs(2017) <= '1';
    layer5_outputs(2018) <= not(layer4_outputs(2073));
    layer5_outputs(2019) <= layer4_outputs(4913);
    layer5_outputs(2020) <= not(layer4_outputs(3764));
    layer5_outputs(2021) <= layer4_outputs(4009);
    layer5_outputs(2022) <= not(layer4_outputs(4158));
    layer5_outputs(2023) <= (layer4_outputs(973)) and (layer4_outputs(3193));
    layer5_outputs(2024) <= not(layer4_outputs(2239));
    layer5_outputs(2025) <= not((layer4_outputs(1971)) and (layer4_outputs(1744)));
    layer5_outputs(2026) <= (layer4_outputs(2576)) and not (layer4_outputs(4203));
    layer5_outputs(2027) <= not((layer4_outputs(3198)) or (layer4_outputs(300)));
    layer5_outputs(2028) <= (layer4_outputs(3562)) and (layer4_outputs(1520));
    layer5_outputs(2029) <= layer4_outputs(4184);
    layer5_outputs(2030) <= not(layer4_outputs(1637));
    layer5_outputs(2031) <= '0';
    layer5_outputs(2032) <= layer4_outputs(4232);
    layer5_outputs(2033) <= layer4_outputs(5114);
    layer5_outputs(2034) <= layer4_outputs(2489);
    layer5_outputs(2035) <= (layer4_outputs(1952)) and not (layer4_outputs(2215));
    layer5_outputs(2036) <= not(layer4_outputs(5048));
    layer5_outputs(2037) <= (layer4_outputs(3306)) or (layer4_outputs(208));
    layer5_outputs(2038) <= not(layer4_outputs(4124));
    layer5_outputs(2039) <= layer4_outputs(3301);
    layer5_outputs(2040) <= layer4_outputs(2487);
    layer5_outputs(2041) <= not(layer4_outputs(1871)) or (layer4_outputs(2957));
    layer5_outputs(2042) <= not(layer4_outputs(1297));
    layer5_outputs(2043) <= layer4_outputs(4049);
    layer5_outputs(2044) <= not(layer4_outputs(787)) or (layer4_outputs(1812));
    layer5_outputs(2045) <= not(layer4_outputs(848)) or (layer4_outputs(5119));
    layer5_outputs(2046) <= not((layer4_outputs(142)) and (layer4_outputs(1737)));
    layer5_outputs(2047) <= not(layer4_outputs(3497));
    layer5_outputs(2048) <= (layer4_outputs(3148)) and not (layer4_outputs(4237));
    layer5_outputs(2049) <= not(layer4_outputs(1273));
    layer5_outputs(2050) <= not(layer4_outputs(2313));
    layer5_outputs(2051) <= not(layer4_outputs(5095));
    layer5_outputs(2052) <= layer4_outputs(1488);
    layer5_outputs(2053) <= not(layer4_outputs(3241));
    layer5_outputs(2054) <= not(layer4_outputs(2656));
    layer5_outputs(2055) <= not(layer4_outputs(4529));
    layer5_outputs(2056) <= '0';
    layer5_outputs(2057) <= not(layer4_outputs(1015));
    layer5_outputs(2058) <= (layer4_outputs(938)) xor (layer4_outputs(3929));
    layer5_outputs(2059) <= not(layer4_outputs(596));
    layer5_outputs(2060) <= layer4_outputs(3181);
    layer5_outputs(2061) <= layer4_outputs(4873);
    layer5_outputs(2062) <= '0';
    layer5_outputs(2063) <= not(layer4_outputs(403)) or (layer4_outputs(2595));
    layer5_outputs(2064) <= not(layer4_outputs(384));
    layer5_outputs(2065) <= not(layer4_outputs(635));
    layer5_outputs(2066) <= not(layer4_outputs(2545));
    layer5_outputs(2067) <= layer4_outputs(4802);
    layer5_outputs(2068) <= layer4_outputs(5055);
    layer5_outputs(2069) <= not((layer4_outputs(1125)) xor (layer4_outputs(3599)));
    layer5_outputs(2070) <= layer4_outputs(4017);
    layer5_outputs(2071) <= not(layer4_outputs(2606)) or (layer4_outputs(5058));
    layer5_outputs(2072) <= not(layer4_outputs(3385));
    layer5_outputs(2073) <= not(layer4_outputs(129));
    layer5_outputs(2074) <= (layer4_outputs(2234)) and not (layer4_outputs(4036));
    layer5_outputs(2075) <= (layer4_outputs(2226)) and not (layer4_outputs(1693));
    layer5_outputs(2076) <= '1';
    layer5_outputs(2077) <= not(layer4_outputs(4963));
    layer5_outputs(2078) <= (layer4_outputs(3803)) and not (layer4_outputs(2064));
    layer5_outputs(2079) <= not((layer4_outputs(1114)) and (layer4_outputs(4465)));
    layer5_outputs(2080) <= (layer4_outputs(3683)) or (layer4_outputs(1852));
    layer5_outputs(2081) <= not(layer4_outputs(805));
    layer5_outputs(2082) <= not(layer4_outputs(36)) or (layer4_outputs(1201));
    layer5_outputs(2083) <= (layer4_outputs(2534)) and not (layer4_outputs(673));
    layer5_outputs(2084) <= (layer4_outputs(1569)) and not (layer4_outputs(318));
    layer5_outputs(2085) <= (layer4_outputs(3181)) and (layer4_outputs(2457));
    layer5_outputs(2086) <= (layer4_outputs(3254)) xor (layer4_outputs(999));
    layer5_outputs(2087) <= not(layer4_outputs(1052));
    layer5_outputs(2088) <= '1';
    layer5_outputs(2089) <= (layer4_outputs(528)) or (layer4_outputs(3655));
    layer5_outputs(2090) <= layer4_outputs(2418);
    layer5_outputs(2091) <= not(layer4_outputs(4484));
    layer5_outputs(2092) <= (layer4_outputs(4320)) or (layer4_outputs(3384));
    layer5_outputs(2093) <= not(layer4_outputs(4441));
    layer5_outputs(2094) <= not(layer4_outputs(4409));
    layer5_outputs(2095) <= not(layer4_outputs(3445));
    layer5_outputs(2096) <= (layer4_outputs(3739)) or (layer4_outputs(1890));
    layer5_outputs(2097) <= not(layer4_outputs(4256)) or (layer4_outputs(2709));
    layer5_outputs(2098) <= not(layer4_outputs(3936));
    layer5_outputs(2099) <= not(layer4_outputs(759));
    layer5_outputs(2100) <= layer4_outputs(4207);
    layer5_outputs(2101) <= not(layer4_outputs(2396));
    layer5_outputs(2102) <= not(layer4_outputs(3603));
    layer5_outputs(2103) <= not((layer4_outputs(3969)) xor (layer4_outputs(3715)));
    layer5_outputs(2104) <= (layer4_outputs(3466)) and not (layer4_outputs(1094));
    layer5_outputs(2105) <= not((layer4_outputs(2313)) and (layer4_outputs(3977)));
    layer5_outputs(2106) <= layer4_outputs(1614);
    layer5_outputs(2107) <= not(layer4_outputs(3975));
    layer5_outputs(2108) <= not(layer4_outputs(711));
    layer5_outputs(2109) <= layer4_outputs(3313);
    layer5_outputs(2110) <= not(layer4_outputs(452)) or (layer4_outputs(2611));
    layer5_outputs(2111) <= '1';
    layer5_outputs(2112) <= not(layer4_outputs(3418));
    layer5_outputs(2113) <= layer4_outputs(5030);
    layer5_outputs(2114) <= (layer4_outputs(4267)) and not (layer4_outputs(4134));
    layer5_outputs(2115) <= layer4_outputs(1504);
    layer5_outputs(2116) <= (layer4_outputs(4099)) and not (layer4_outputs(1665));
    layer5_outputs(2117) <= (layer4_outputs(2259)) and not (layer4_outputs(2981));
    layer5_outputs(2118) <= not((layer4_outputs(725)) or (layer4_outputs(1913)));
    layer5_outputs(2119) <= layer4_outputs(4260);
    layer5_outputs(2120) <= not(layer4_outputs(3420));
    layer5_outputs(2121) <= not(layer4_outputs(2202)) or (layer4_outputs(1987));
    layer5_outputs(2122) <= not(layer4_outputs(1176));
    layer5_outputs(2123) <= not(layer4_outputs(3821));
    layer5_outputs(2124) <= not((layer4_outputs(3700)) and (layer4_outputs(2559)));
    layer5_outputs(2125) <= not((layer4_outputs(342)) or (layer4_outputs(576)));
    layer5_outputs(2126) <= (layer4_outputs(3234)) and (layer4_outputs(1680));
    layer5_outputs(2127) <= '1';
    layer5_outputs(2128) <= not(layer4_outputs(5006)) or (layer4_outputs(3832));
    layer5_outputs(2129) <= layer4_outputs(3157);
    layer5_outputs(2130) <= (layer4_outputs(5061)) and not (layer4_outputs(1111));
    layer5_outputs(2131) <= layer4_outputs(2607);
    layer5_outputs(2132) <= layer4_outputs(2380);
    layer5_outputs(2133) <= not(layer4_outputs(3991));
    layer5_outputs(2134) <= not(layer4_outputs(4918));
    layer5_outputs(2135) <= not(layer4_outputs(683)) or (layer4_outputs(1200));
    layer5_outputs(2136) <= not(layer4_outputs(591));
    layer5_outputs(2137) <= not((layer4_outputs(4224)) xor (layer4_outputs(1700)));
    layer5_outputs(2138) <= not(layer4_outputs(1095));
    layer5_outputs(2139) <= not((layer4_outputs(699)) xor (layer4_outputs(432)));
    layer5_outputs(2140) <= (layer4_outputs(686)) and not (layer4_outputs(5041));
    layer5_outputs(2141) <= not(layer4_outputs(912));
    layer5_outputs(2142) <= layer4_outputs(3079);
    layer5_outputs(2143) <= (layer4_outputs(4183)) and (layer4_outputs(1854));
    layer5_outputs(2144) <= not(layer4_outputs(2637));
    layer5_outputs(2145) <= layer4_outputs(2489);
    layer5_outputs(2146) <= (layer4_outputs(371)) and not (layer4_outputs(2690));
    layer5_outputs(2147) <= not((layer4_outputs(3957)) and (layer4_outputs(4977)));
    layer5_outputs(2148) <= layer4_outputs(2287);
    layer5_outputs(2149) <= layer4_outputs(385);
    layer5_outputs(2150) <= (layer4_outputs(389)) and (layer4_outputs(2902));
    layer5_outputs(2151) <= (layer4_outputs(2103)) and (layer4_outputs(3791));
    layer5_outputs(2152) <= not((layer4_outputs(2163)) xor (layer4_outputs(4488)));
    layer5_outputs(2153) <= not(layer4_outputs(48));
    layer5_outputs(2154) <= (layer4_outputs(897)) xor (layer4_outputs(3149));
    layer5_outputs(2155) <= (layer4_outputs(2594)) xor (layer4_outputs(2199));
    layer5_outputs(2156) <= '1';
    layer5_outputs(2157) <= (layer4_outputs(4922)) xor (layer4_outputs(3748));
    layer5_outputs(2158) <= not((layer4_outputs(4843)) xor (layer4_outputs(462)));
    layer5_outputs(2159) <= (layer4_outputs(1702)) and not (layer4_outputs(85));
    layer5_outputs(2160) <= not(layer4_outputs(3485));
    layer5_outputs(2161) <= not((layer4_outputs(2459)) or (layer4_outputs(1349)));
    layer5_outputs(2162) <= (layer4_outputs(2625)) xor (layer4_outputs(2719));
    layer5_outputs(2163) <= layer4_outputs(2802);
    layer5_outputs(2164) <= layer4_outputs(121);
    layer5_outputs(2165) <= not(layer4_outputs(4785));
    layer5_outputs(2166) <= layer4_outputs(2583);
    layer5_outputs(2167) <= layer4_outputs(3768);
    layer5_outputs(2168) <= (layer4_outputs(5088)) or (layer4_outputs(43));
    layer5_outputs(2169) <= (layer4_outputs(4774)) and not (layer4_outputs(823));
    layer5_outputs(2170) <= '0';
    layer5_outputs(2171) <= not(layer4_outputs(4595));
    layer5_outputs(2172) <= not(layer4_outputs(3010));
    layer5_outputs(2173) <= not(layer4_outputs(780)) or (layer4_outputs(4801));
    layer5_outputs(2174) <= not(layer4_outputs(4843));
    layer5_outputs(2175) <= not(layer4_outputs(2803));
    layer5_outputs(2176) <= not(layer4_outputs(3742));
    layer5_outputs(2177) <= layer4_outputs(3419);
    layer5_outputs(2178) <= not((layer4_outputs(927)) or (layer4_outputs(1914)));
    layer5_outputs(2179) <= (layer4_outputs(3633)) or (layer4_outputs(4882));
    layer5_outputs(2180) <= layer4_outputs(2630);
    layer5_outputs(2181) <= not((layer4_outputs(2816)) and (layer4_outputs(2477)));
    layer5_outputs(2182) <= not(layer4_outputs(4351));
    layer5_outputs(2183) <= (layer4_outputs(1631)) xor (layer4_outputs(3145));
    layer5_outputs(2184) <= not(layer4_outputs(3033)) or (layer4_outputs(2948));
    layer5_outputs(2185) <= layer4_outputs(4704);
    layer5_outputs(2186) <= not(layer4_outputs(609));
    layer5_outputs(2187) <= layer4_outputs(4408);
    layer5_outputs(2188) <= (layer4_outputs(1677)) and (layer4_outputs(2632));
    layer5_outputs(2189) <= not(layer4_outputs(4359));
    layer5_outputs(2190) <= (layer4_outputs(3883)) xor (layer4_outputs(1753));
    layer5_outputs(2191) <= not((layer4_outputs(2966)) or (layer4_outputs(3601)));
    layer5_outputs(2192) <= not((layer4_outputs(4089)) and (layer4_outputs(2165)));
    layer5_outputs(2193) <= not(layer4_outputs(2251)) or (layer4_outputs(1818));
    layer5_outputs(2194) <= (layer4_outputs(3025)) and (layer4_outputs(3407));
    layer5_outputs(2195) <= layer4_outputs(4481);
    layer5_outputs(2196) <= '0';
    layer5_outputs(2197) <= not(layer4_outputs(1022));
    layer5_outputs(2198) <= not(layer4_outputs(86));
    layer5_outputs(2199) <= layer4_outputs(194);
    layer5_outputs(2200) <= (layer4_outputs(140)) and (layer4_outputs(961));
    layer5_outputs(2201) <= (layer4_outputs(1152)) or (layer4_outputs(2578));
    layer5_outputs(2202) <= (layer4_outputs(2127)) and not (layer4_outputs(90));
    layer5_outputs(2203) <= (layer4_outputs(5025)) or (layer4_outputs(2470));
    layer5_outputs(2204) <= (layer4_outputs(2244)) and not (layer4_outputs(2370));
    layer5_outputs(2205) <= not(layer4_outputs(4573));
    layer5_outputs(2206) <= layer4_outputs(3405);
    layer5_outputs(2207) <= (layer4_outputs(2464)) and not (layer4_outputs(4600));
    layer5_outputs(2208) <= not((layer4_outputs(3212)) or (layer4_outputs(1898)));
    layer5_outputs(2209) <= layer4_outputs(2456);
    layer5_outputs(2210) <= layer4_outputs(1475);
    layer5_outputs(2211) <= not(layer4_outputs(1055));
    layer5_outputs(2212) <= '0';
    layer5_outputs(2213) <= not(layer4_outputs(2169)) or (layer4_outputs(1851));
    layer5_outputs(2214) <= layer4_outputs(3126);
    layer5_outputs(2215) <= layer4_outputs(1165);
    layer5_outputs(2216) <= (layer4_outputs(1610)) and not (layer4_outputs(2152));
    layer5_outputs(2217) <= layer4_outputs(3796);
    layer5_outputs(2218) <= (layer4_outputs(4588)) and not (layer4_outputs(3961));
    layer5_outputs(2219) <= not(layer4_outputs(2623));
    layer5_outputs(2220) <= not(layer4_outputs(2894));
    layer5_outputs(2221) <= '1';
    layer5_outputs(2222) <= layer4_outputs(1382);
    layer5_outputs(2223) <= (layer4_outputs(2987)) or (layer4_outputs(2547));
    layer5_outputs(2224) <= (layer4_outputs(1499)) xor (layer4_outputs(2156));
    layer5_outputs(2225) <= not(layer4_outputs(2651));
    layer5_outputs(2226) <= (layer4_outputs(2)) or (layer4_outputs(4689));
    layer5_outputs(2227) <= layer4_outputs(3297);
    layer5_outputs(2228) <= (layer4_outputs(3350)) and not (layer4_outputs(3292));
    layer5_outputs(2229) <= '0';
    layer5_outputs(2230) <= not((layer4_outputs(5016)) or (layer4_outputs(4873)));
    layer5_outputs(2231) <= not(layer4_outputs(2079));
    layer5_outputs(2232) <= not((layer4_outputs(362)) or (layer4_outputs(4051)));
    layer5_outputs(2233) <= '0';
    layer5_outputs(2234) <= '0';
    layer5_outputs(2235) <= not(layer4_outputs(1529)) or (layer4_outputs(3223));
    layer5_outputs(2236) <= not(layer4_outputs(5033));
    layer5_outputs(2237) <= not(layer4_outputs(4396));
    layer5_outputs(2238) <= (layer4_outputs(3731)) and not (layer4_outputs(317));
    layer5_outputs(2239) <= not(layer4_outputs(2532));
    layer5_outputs(2240) <= (layer4_outputs(4106)) and not (layer4_outputs(3978));
    layer5_outputs(2241) <= (layer4_outputs(538)) xor (layer4_outputs(4725));
    layer5_outputs(2242) <= layer4_outputs(4882);
    layer5_outputs(2243) <= (layer4_outputs(3367)) and not (layer4_outputs(55));
    layer5_outputs(2244) <= not(layer4_outputs(699));
    layer5_outputs(2245) <= layer4_outputs(3927);
    layer5_outputs(2246) <= (layer4_outputs(3081)) and not (layer4_outputs(4994));
    layer5_outputs(2247) <= layer4_outputs(4391);
    layer5_outputs(2248) <= not(layer4_outputs(1098)) or (layer4_outputs(4503));
    layer5_outputs(2249) <= layer4_outputs(536);
    layer5_outputs(2250) <= not((layer4_outputs(1157)) or (layer4_outputs(1336)));
    layer5_outputs(2251) <= layer4_outputs(3615);
    layer5_outputs(2252) <= (layer4_outputs(992)) and not (layer4_outputs(3139));
    layer5_outputs(2253) <= layer4_outputs(3592);
    layer5_outputs(2254) <= layer4_outputs(3786);
    layer5_outputs(2255) <= not(layer4_outputs(5033)) or (layer4_outputs(670));
    layer5_outputs(2256) <= not(layer4_outputs(4440)) or (layer4_outputs(3857));
    layer5_outputs(2257) <= layer4_outputs(2390);
    layer5_outputs(2258) <= (layer4_outputs(1875)) or (layer4_outputs(864));
    layer5_outputs(2259) <= (layer4_outputs(4438)) and not (layer4_outputs(2327));
    layer5_outputs(2260) <= not(layer4_outputs(764));
    layer5_outputs(2261) <= not(layer4_outputs(1819)) or (layer4_outputs(739));
    layer5_outputs(2262) <= not(layer4_outputs(163));
    layer5_outputs(2263) <= (layer4_outputs(3826)) xor (layer4_outputs(263));
    layer5_outputs(2264) <= layer4_outputs(4278);
    layer5_outputs(2265) <= not(layer4_outputs(1065));
    layer5_outputs(2266) <= not(layer4_outputs(4399)) or (layer4_outputs(1764));
    layer5_outputs(2267) <= not(layer4_outputs(2822));
    layer5_outputs(2268) <= (layer4_outputs(1734)) and (layer4_outputs(1433));
    layer5_outputs(2269) <= layer4_outputs(3858);
    layer5_outputs(2270) <= not(layer4_outputs(4163));
    layer5_outputs(2271) <= not((layer4_outputs(4543)) xor (layer4_outputs(2560)));
    layer5_outputs(2272) <= (layer4_outputs(1551)) and not (layer4_outputs(2360));
    layer5_outputs(2273) <= (layer4_outputs(2008)) or (layer4_outputs(3203));
    layer5_outputs(2274) <= (layer4_outputs(1312)) and (layer4_outputs(2925));
    layer5_outputs(2275) <= layer4_outputs(4207);
    layer5_outputs(2276) <= not(layer4_outputs(4473));
    layer5_outputs(2277) <= not(layer4_outputs(4656));
    layer5_outputs(2278) <= layer4_outputs(3411);
    layer5_outputs(2279) <= layer4_outputs(2545);
    layer5_outputs(2280) <= '0';
    layer5_outputs(2281) <= not((layer4_outputs(65)) or (layer4_outputs(2860)));
    layer5_outputs(2282) <= (layer4_outputs(4171)) and not (layer4_outputs(1681));
    layer5_outputs(2283) <= '0';
    layer5_outputs(2284) <= (layer4_outputs(3388)) and not (layer4_outputs(4146));
    layer5_outputs(2285) <= not(layer4_outputs(2521));
    layer5_outputs(2286) <= (layer4_outputs(2334)) xor (layer4_outputs(3339));
    layer5_outputs(2287) <= (layer4_outputs(2897)) or (layer4_outputs(2496));
    layer5_outputs(2288) <= layer4_outputs(4007);
    layer5_outputs(2289) <= layer4_outputs(2767);
    layer5_outputs(2290) <= (layer4_outputs(2277)) and not (layer4_outputs(1432));
    layer5_outputs(2291) <= layer4_outputs(2704);
    layer5_outputs(2292) <= layer4_outputs(1749);
    layer5_outputs(2293) <= (layer4_outputs(14)) or (layer4_outputs(4094));
    layer5_outputs(2294) <= layer4_outputs(4429);
    layer5_outputs(2295) <= (layer4_outputs(2325)) or (layer4_outputs(572));
    layer5_outputs(2296) <= (layer4_outputs(2798)) and (layer4_outputs(4371));
    layer5_outputs(2297) <= not((layer4_outputs(900)) and (layer4_outputs(1422)));
    layer5_outputs(2298) <= (layer4_outputs(1272)) and not (layer4_outputs(127));
    layer5_outputs(2299) <= (layer4_outputs(3624)) xor (layer4_outputs(4180));
    layer5_outputs(2300) <= '1';
    layer5_outputs(2301) <= (layer4_outputs(4971)) and not (layer4_outputs(369));
    layer5_outputs(2302) <= not((layer4_outputs(3903)) and (layer4_outputs(4464)));
    layer5_outputs(2303) <= not(layer4_outputs(3725)) or (layer4_outputs(889));
    layer5_outputs(2304) <= not(layer4_outputs(1848)) or (layer4_outputs(4510));
    layer5_outputs(2305) <= layer4_outputs(471);
    layer5_outputs(2306) <= not((layer4_outputs(873)) or (layer4_outputs(284)));
    layer5_outputs(2307) <= (layer4_outputs(3087)) and not (layer4_outputs(2112));
    layer5_outputs(2308) <= (layer4_outputs(3812)) and not (layer4_outputs(4237));
    layer5_outputs(2309) <= not(layer4_outputs(1060)) or (layer4_outputs(4597));
    layer5_outputs(2310) <= not(layer4_outputs(1709)) or (layer4_outputs(2739));
    layer5_outputs(2311) <= (layer4_outputs(2009)) xor (layer4_outputs(4227));
    layer5_outputs(2312) <= not(layer4_outputs(843));
    layer5_outputs(2313) <= (layer4_outputs(630)) and (layer4_outputs(4246));
    layer5_outputs(2314) <= (layer4_outputs(1328)) and (layer4_outputs(4289));
    layer5_outputs(2315) <= (layer4_outputs(2628)) xor (layer4_outputs(3453));
    layer5_outputs(2316) <= (layer4_outputs(1154)) and (layer4_outputs(1393));
    layer5_outputs(2317) <= '0';
    layer5_outputs(2318) <= not(layer4_outputs(502));
    layer5_outputs(2319) <= (layer4_outputs(1379)) and (layer4_outputs(3430));
    layer5_outputs(2320) <= (layer4_outputs(3938)) and not (layer4_outputs(2873));
    layer5_outputs(2321) <= layer4_outputs(2941);
    layer5_outputs(2322) <= '0';
    layer5_outputs(2323) <= not(layer4_outputs(854));
    layer5_outputs(2324) <= layer4_outputs(1289);
    layer5_outputs(2325) <= not(layer4_outputs(145));
    layer5_outputs(2326) <= (layer4_outputs(2246)) or (layer4_outputs(1682));
    layer5_outputs(2327) <= (layer4_outputs(1160)) and not (layer4_outputs(2273));
    layer5_outputs(2328) <= not(layer4_outputs(916));
    layer5_outputs(2329) <= not(layer4_outputs(4249));
    layer5_outputs(2330) <= layer4_outputs(102);
    layer5_outputs(2331) <= layer4_outputs(569);
    layer5_outputs(2332) <= not(layer4_outputs(1601));
    layer5_outputs(2333) <= not(layer4_outputs(249));
    layer5_outputs(2334) <= (layer4_outputs(438)) xor (layer4_outputs(5040));
    layer5_outputs(2335) <= (layer4_outputs(3689)) and not (layer4_outputs(2824));
    layer5_outputs(2336) <= layer4_outputs(964);
    layer5_outputs(2337) <= not(layer4_outputs(2646)) or (layer4_outputs(4355));
    layer5_outputs(2338) <= '1';
    layer5_outputs(2339) <= not(layer4_outputs(1645)) or (layer4_outputs(4210));
    layer5_outputs(2340) <= layer4_outputs(3321);
    layer5_outputs(2341) <= layer4_outputs(2131);
    layer5_outputs(2342) <= not((layer4_outputs(4353)) or (layer4_outputs(1065)));
    layer5_outputs(2343) <= (layer4_outputs(2727)) or (layer4_outputs(4797));
    layer5_outputs(2344) <= layer4_outputs(744);
    layer5_outputs(2345) <= not(layer4_outputs(2450));
    layer5_outputs(2346) <= not(layer4_outputs(1404));
    layer5_outputs(2347) <= not(layer4_outputs(3543));
    layer5_outputs(2348) <= not(layer4_outputs(510)) or (layer4_outputs(4502));
    layer5_outputs(2349) <= layer4_outputs(3186);
    layer5_outputs(2350) <= not(layer4_outputs(4217));
    layer5_outputs(2351) <= (layer4_outputs(1465)) and not (layer4_outputs(2366));
    layer5_outputs(2352) <= (layer4_outputs(3347)) or (layer4_outputs(651));
    layer5_outputs(2353) <= not(layer4_outputs(9));
    layer5_outputs(2354) <= not(layer4_outputs(1317));
    layer5_outputs(2355) <= not(layer4_outputs(370));
    layer5_outputs(2356) <= '1';
    layer5_outputs(2357) <= layer4_outputs(2458);
    layer5_outputs(2358) <= not(layer4_outputs(4767));
    layer5_outputs(2359) <= not(layer4_outputs(1272));
    layer5_outputs(2360) <= not(layer4_outputs(4871));
    layer5_outputs(2361) <= layer4_outputs(3867);
    layer5_outputs(2362) <= not(layer4_outputs(2228));
    layer5_outputs(2363) <= not(layer4_outputs(2697));
    layer5_outputs(2364) <= (layer4_outputs(3096)) and not (layer4_outputs(3134));
    layer5_outputs(2365) <= (layer4_outputs(724)) and (layer4_outputs(3315));
    layer5_outputs(2366) <= layer4_outputs(3282);
    layer5_outputs(2367) <= (layer4_outputs(3062)) and (layer4_outputs(1757));
    layer5_outputs(2368) <= layer4_outputs(1231);
    layer5_outputs(2369) <= not(layer4_outputs(942));
    layer5_outputs(2370) <= not(layer4_outputs(4034)) or (layer4_outputs(4336));
    layer5_outputs(2371) <= not(layer4_outputs(1960));
    layer5_outputs(2372) <= not(layer4_outputs(1252));
    layer5_outputs(2373) <= not(layer4_outputs(792));
    layer5_outputs(2374) <= not((layer4_outputs(2601)) xor (layer4_outputs(5105)));
    layer5_outputs(2375) <= not((layer4_outputs(4367)) and (layer4_outputs(3927)));
    layer5_outputs(2376) <= (layer4_outputs(2081)) xor (layer4_outputs(201));
    layer5_outputs(2377) <= layer4_outputs(1326);
    layer5_outputs(2378) <= not(layer4_outputs(3199));
    layer5_outputs(2379) <= '0';
    layer5_outputs(2380) <= layer4_outputs(1811);
    layer5_outputs(2381) <= (layer4_outputs(484)) or (layer4_outputs(4019));
    layer5_outputs(2382) <= not(layer4_outputs(1933)) or (layer4_outputs(910));
    layer5_outputs(2383) <= (layer4_outputs(2537)) and (layer4_outputs(4598));
    layer5_outputs(2384) <= not(layer4_outputs(4737));
    layer5_outputs(2385) <= (layer4_outputs(1958)) and (layer4_outputs(1585));
    layer5_outputs(2386) <= not(layer4_outputs(1545)) or (layer4_outputs(2146));
    layer5_outputs(2387) <= not(layer4_outputs(2678));
    layer5_outputs(2388) <= layer4_outputs(3906);
    layer5_outputs(2389) <= '1';
    layer5_outputs(2390) <= not(layer4_outputs(1350));
    layer5_outputs(2391) <= not((layer4_outputs(4195)) and (layer4_outputs(4798)));
    layer5_outputs(2392) <= layer4_outputs(1898);
    layer5_outputs(2393) <= layer4_outputs(5013);
    layer5_outputs(2394) <= not((layer4_outputs(1042)) xor (layer4_outputs(4863)));
    layer5_outputs(2395) <= not(layer4_outputs(1708));
    layer5_outputs(2396) <= not(layer4_outputs(2829)) or (layer4_outputs(3169));
    layer5_outputs(2397) <= not(layer4_outputs(1475));
    layer5_outputs(2398) <= (layer4_outputs(1662)) and not (layer4_outputs(51));
    layer5_outputs(2399) <= not(layer4_outputs(2712)) or (layer4_outputs(322));
    layer5_outputs(2400) <= (layer4_outputs(3116)) and (layer4_outputs(4428));
    layer5_outputs(2401) <= not(layer4_outputs(4211));
    layer5_outputs(2402) <= not(layer4_outputs(3472));
    layer5_outputs(2403) <= not(layer4_outputs(4748));
    layer5_outputs(2404) <= not(layer4_outputs(1981));
    layer5_outputs(2405) <= not(layer4_outputs(326));
    layer5_outputs(2406) <= (layer4_outputs(2194)) and (layer4_outputs(3241));
    layer5_outputs(2407) <= (layer4_outputs(2681)) xor (layer4_outputs(1554));
    layer5_outputs(2408) <= (layer4_outputs(4566)) xor (layer4_outputs(606));
    layer5_outputs(2409) <= layer4_outputs(2196);
    layer5_outputs(2410) <= (layer4_outputs(2566)) xor (layer4_outputs(2085));
    layer5_outputs(2411) <= not(layer4_outputs(4010));
    layer5_outputs(2412) <= (layer4_outputs(4695)) and (layer4_outputs(2480));
    layer5_outputs(2413) <= not(layer4_outputs(235));
    layer5_outputs(2414) <= (layer4_outputs(1959)) xor (layer4_outputs(1925));
    layer5_outputs(2415) <= not(layer4_outputs(2936));
    layer5_outputs(2416) <= not(layer4_outputs(2296)) or (layer4_outputs(3364));
    layer5_outputs(2417) <= (layer4_outputs(1765)) and not (layer4_outputs(1224));
    layer5_outputs(2418) <= not(layer4_outputs(3486));
    layer5_outputs(2419) <= layer4_outputs(977);
    layer5_outputs(2420) <= (layer4_outputs(94)) xor (layer4_outputs(1206));
    layer5_outputs(2421) <= (layer4_outputs(4831)) and not (layer4_outputs(4750));
    layer5_outputs(2422) <= '1';
    layer5_outputs(2423) <= '0';
    layer5_outputs(2424) <= not(layer4_outputs(915));
    layer5_outputs(2425) <= (layer4_outputs(3295)) or (layer4_outputs(3567));
    layer5_outputs(2426) <= not(layer4_outputs(4050)) or (layer4_outputs(1012));
    layer5_outputs(2427) <= not(layer4_outputs(3189));
    layer5_outputs(2428) <= not(layer4_outputs(4869));
    layer5_outputs(2429) <= not(layer4_outputs(885));
    layer5_outputs(2430) <= (layer4_outputs(1292)) and not (layer4_outputs(4516));
    layer5_outputs(2431) <= not(layer4_outputs(1842));
    layer5_outputs(2432) <= layer4_outputs(669);
    layer5_outputs(2433) <= not((layer4_outputs(2477)) or (layer4_outputs(4308)));
    layer5_outputs(2434) <= layer4_outputs(3874);
    layer5_outputs(2435) <= not(layer4_outputs(2562)) or (layer4_outputs(923));
    layer5_outputs(2436) <= layer4_outputs(3674);
    layer5_outputs(2437) <= layer4_outputs(1791);
    layer5_outputs(2438) <= not(layer4_outputs(3566));
    layer5_outputs(2439) <= not((layer4_outputs(4126)) and (layer4_outputs(2406)));
    layer5_outputs(2440) <= not(layer4_outputs(2617)) or (layer4_outputs(395));
    layer5_outputs(2441) <= not(layer4_outputs(4834));
    layer5_outputs(2442) <= (layer4_outputs(2138)) or (layer4_outputs(4400));
    layer5_outputs(2443) <= not((layer4_outputs(1533)) and (layer4_outputs(456)));
    layer5_outputs(2444) <= not(layer4_outputs(383));
    layer5_outputs(2445) <= (layer4_outputs(4490)) xor (layer4_outputs(1736));
    layer5_outputs(2446) <= (layer4_outputs(976)) and not (layer4_outputs(5113));
    layer5_outputs(2447) <= layer4_outputs(3949);
    layer5_outputs(2448) <= (layer4_outputs(1557)) and not (layer4_outputs(2626));
    layer5_outputs(2449) <= not(layer4_outputs(3381));
    layer5_outputs(2450) <= (layer4_outputs(3758)) and not (layer4_outputs(181));
    layer5_outputs(2451) <= layer4_outputs(3435);
    layer5_outputs(2452) <= (layer4_outputs(3480)) and (layer4_outputs(4115));
    layer5_outputs(2453) <= layer4_outputs(3558);
    layer5_outputs(2454) <= (layer4_outputs(4344)) or (layer4_outputs(2308));
    layer5_outputs(2455) <= layer4_outputs(4282);
    layer5_outputs(2456) <= layer4_outputs(81);
    layer5_outputs(2457) <= layer4_outputs(2214);
    layer5_outputs(2458) <= not(layer4_outputs(4308));
    layer5_outputs(2459) <= layer4_outputs(3098);
    layer5_outputs(2460) <= (layer4_outputs(2517)) or (layer4_outputs(3965));
    layer5_outputs(2461) <= layer4_outputs(4111);
    layer5_outputs(2462) <= (layer4_outputs(2953)) and not (layer4_outputs(291));
    layer5_outputs(2463) <= layer4_outputs(2822);
    layer5_outputs(2464) <= not(layer4_outputs(2032)) or (layer4_outputs(4307));
    layer5_outputs(2465) <= not((layer4_outputs(5083)) xor (layer4_outputs(4826)));
    layer5_outputs(2466) <= (layer4_outputs(109)) and (layer4_outputs(1337));
    layer5_outputs(2467) <= not((layer4_outputs(1246)) xor (layer4_outputs(2645)));
    layer5_outputs(2468) <= not(layer4_outputs(715)) or (layer4_outputs(4755));
    layer5_outputs(2469) <= not(layer4_outputs(3465));
    layer5_outputs(2470) <= layer4_outputs(2574);
    layer5_outputs(2471) <= not(layer4_outputs(566));
    layer5_outputs(2472) <= layer4_outputs(1812);
    layer5_outputs(2473) <= (layer4_outputs(2697)) or (layer4_outputs(1760));
    layer5_outputs(2474) <= not(layer4_outputs(1128));
    layer5_outputs(2475) <= layer4_outputs(2026);
    layer5_outputs(2476) <= not(layer4_outputs(2555));
    layer5_outputs(2477) <= not(layer4_outputs(3901));
    layer5_outputs(2478) <= not((layer4_outputs(763)) or (layer4_outputs(1817)));
    layer5_outputs(2479) <= not((layer4_outputs(3958)) xor (layer4_outputs(4220)));
    layer5_outputs(2480) <= not((layer4_outputs(4431)) xor (layer4_outputs(3171)));
    layer5_outputs(2481) <= (layer4_outputs(1153)) xor (layer4_outputs(3830));
    layer5_outputs(2482) <= layer4_outputs(2780);
    layer5_outputs(2483) <= layer4_outputs(297);
    layer5_outputs(2484) <= layer4_outputs(4143);
    layer5_outputs(2485) <= (layer4_outputs(4615)) and not (layer4_outputs(1758));
    layer5_outputs(2486) <= (layer4_outputs(605)) and not (layer4_outputs(2075));
    layer5_outputs(2487) <= (layer4_outputs(811)) and not (layer4_outputs(1746));
    layer5_outputs(2488) <= not(layer4_outputs(4335));
    layer5_outputs(2489) <= layer4_outputs(5110);
    layer5_outputs(2490) <= not(layer4_outputs(969));
    layer5_outputs(2491) <= (layer4_outputs(1566)) and not (layer4_outputs(3615));
    layer5_outputs(2492) <= not(layer4_outputs(3525));
    layer5_outputs(2493) <= (layer4_outputs(1053)) and not (layer4_outputs(4969));
    layer5_outputs(2494) <= not(layer4_outputs(371));
    layer5_outputs(2495) <= not(layer4_outputs(4358));
    layer5_outputs(2496) <= not((layer4_outputs(3579)) xor (layer4_outputs(3660)));
    layer5_outputs(2497) <= (layer4_outputs(1130)) and not (layer4_outputs(1107));
    layer5_outputs(2498) <= (layer4_outputs(2318)) and not (layer4_outputs(1434));
    layer5_outputs(2499) <= not(layer4_outputs(2771));
    layer5_outputs(2500) <= not((layer4_outputs(1617)) and (layer4_outputs(4046)));
    layer5_outputs(2501) <= not((layer4_outputs(3574)) or (layer4_outputs(2643)));
    layer5_outputs(2502) <= (layer4_outputs(755)) xor (layer4_outputs(2629));
    layer5_outputs(2503) <= not(layer4_outputs(2048)) or (layer4_outputs(4205));
    layer5_outputs(2504) <= layer4_outputs(3657);
    layer5_outputs(2505) <= (layer4_outputs(1522)) or (layer4_outputs(1779));
    layer5_outputs(2506) <= not((layer4_outputs(3622)) xor (layer4_outputs(4075)));
    layer5_outputs(2507) <= '0';
    layer5_outputs(2508) <= (layer4_outputs(2294)) and (layer4_outputs(2420));
    layer5_outputs(2509) <= not(layer4_outputs(3703));
    layer5_outputs(2510) <= (layer4_outputs(2329)) and (layer4_outputs(800));
    layer5_outputs(2511) <= (layer4_outputs(4889)) xor (layer4_outputs(4964));
    layer5_outputs(2512) <= (layer4_outputs(2549)) and (layer4_outputs(459));
    layer5_outputs(2513) <= (layer4_outputs(447)) and (layer4_outputs(813));
    layer5_outputs(2514) <= (layer4_outputs(2282)) xor (layer4_outputs(607));
    layer5_outputs(2515) <= not(layer4_outputs(2798)) or (layer4_outputs(1845));
    layer5_outputs(2516) <= not(layer4_outputs(3551));
    layer5_outputs(2517) <= not(layer4_outputs(3544)) or (layer4_outputs(3380));
    layer5_outputs(2518) <= not(layer4_outputs(4167));
    layer5_outputs(2519) <= layer4_outputs(569);
    layer5_outputs(2520) <= not(layer4_outputs(1723)) or (layer4_outputs(5087));
    layer5_outputs(2521) <= layer4_outputs(4886);
    layer5_outputs(2522) <= layer4_outputs(4529);
    layer5_outputs(2523) <= (layer4_outputs(4948)) or (layer4_outputs(1755));
    layer5_outputs(2524) <= layer4_outputs(465);
    layer5_outputs(2525) <= not(layer4_outputs(346));
    layer5_outputs(2526) <= layer4_outputs(4086);
    layer5_outputs(2527) <= '1';
    layer5_outputs(2528) <= layer4_outputs(4276);
    layer5_outputs(2529) <= layer4_outputs(1367);
    layer5_outputs(2530) <= layer4_outputs(3706);
    layer5_outputs(2531) <= not(layer4_outputs(601)) or (layer4_outputs(2790));
    layer5_outputs(2532) <= not((layer4_outputs(3162)) or (layer4_outputs(317)));
    layer5_outputs(2533) <= not((layer4_outputs(3893)) xor (layer4_outputs(4376)));
    layer5_outputs(2534) <= layer4_outputs(2097);
    layer5_outputs(2535) <= layer4_outputs(3664);
    layer5_outputs(2536) <= layer4_outputs(1257);
    layer5_outputs(2537) <= not(layer4_outputs(2473)) or (layer4_outputs(1779));
    layer5_outputs(2538) <= not((layer4_outputs(3270)) and (layer4_outputs(966)));
    layer5_outputs(2539) <= not(layer4_outputs(2718));
    layer5_outputs(2540) <= (layer4_outputs(1978)) or (layer4_outputs(2835));
    layer5_outputs(2541) <= (layer4_outputs(2268)) or (layer4_outputs(2427));
    layer5_outputs(2542) <= layer4_outputs(2736);
    layer5_outputs(2543) <= not((layer4_outputs(2170)) or (layer4_outputs(4731)));
    layer5_outputs(2544) <= (layer4_outputs(854)) and not (layer4_outputs(3737));
    layer5_outputs(2545) <= (layer4_outputs(683)) xor (layer4_outputs(1062));
    layer5_outputs(2546) <= layer4_outputs(2050);
    layer5_outputs(2547) <= not(layer4_outputs(4192));
    layer5_outputs(2548) <= not(layer4_outputs(3142));
    layer5_outputs(2549) <= layer4_outputs(3135);
    layer5_outputs(2550) <= layer4_outputs(4328);
    layer5_outputs(2551) <= not((layer4_outputs(3392)) xor (layer4_outputs(3303)));
    layer5_outputs(2552) <= not(layer4_outputs(4614));
    layer5_outputs(2553) <= not(layer4_outputs(3939));
    layer5_outputs(2554) <= (layer4_outputs(4755)) and not (layer4_outputs(3414));
    layer5_outputs(2555) <= not(layer4_outputs(1819));
    layer5_outputs(2556) <= layer4_outputs(984);
    layer5_outputs(2557) <= layer4_outputs(1842);
    layer5_outputs(2558) <= (layer4_outputs(2430)) xor (layer4_outputs(2719));
    layer5_outputs(2559) <= not(layer4_outputs(821));
    layer5_outputs(2560) <= not((layer4_outputs(2907)) or (layer4_outputs(772)));
    layer5_outputs(2561) <= not(layer4_outputs(4390));
    layer5_outputs(2562) <= (layer4_outputs(4204)) and not (layer4_outputs(1603));
    layer5_outputs(2563) <= (layer4_outputs(2909)) and (layer4_outputs(3586));
    layer5_outputs(2564) <= layer4_outputs(2132);
    layer5_outputs(2565) <= layer4_outputs(754);
    layer5_outputs(2566) <= layer4_outputs(2205);
    layer5_outputs(2567) <= (layer4_outputs(314)) and (layer4_outputs(2616));
    layer5_outputs(2568) <= (layer4_outputs(760)) or (layer4_outputs(4812));
    layer5_outputs(2569) <= not((layer4_outputs(3476)) xor (layer4_outputs(2290)));
    layer5_outputs(2570) <= layer4_outputs(3941);
    layer5_outputs(2571) <= not(layer4_outputs(4787));
    layer5_outputs(2572) <= not((layer4_outputs(3372)) xor (layer4_outputs(3176)));
    layer5_outputs(2573) <= not((layer4_outputs(2244)) or (layer4_outputs(2551)));
    layer5_outputs(2574) <= not((layer4_outputs(3523)) or (layer4_outputs(1499)));
    layer5_outputs(2575) <= (layer4_outputs(3107)) or (layer4_outputs(2616));
    layer5_outputs(2576) <= '0';
    layer5_outputs(2577) <= not(layer4_outputs(2457)) or (layer4_outputs(4729));
    layer5_outputs(2578) <= not((layer4_outputs(4863)) and (layer4_outputs(1503)));
    layer5_outputs(2579) <= not(layer4_outputs(3082));
    layer5_outputs(2580) <= not(layer4_outputs(796)) or (layer4_outputs(165));
    layer5_outputs(2581) <= layer4_outputs(129);
    layer5_outputs(2582) <= not(layer4_outputs(2076)) or (layer4_outputs(2740));
    layer5_outputs(2583) <= layer4_outputs(4794);
    layer5_outputs(2584) <= not(layer4_outputs(3728));
    layer5_outputs(2585) <= layer4_outputs(3257);
    layer5_outputs(2586) <= (layer4_outputs(3823)) and not (layer4_outputs(430));
    layer5_outputs(2587) <= layer4_outputs(898);
    layer5_outputs(2588) <= layer4_outputs(1647);
    layer5_outputs(2589) <= (layer4_outputs(3138)) and not (layer4_outputs(4830));
    layer5_outputs(2590) <= (layer4_outputs(4903)) and (layer4_outputs(3009));
    layer5_outputs(2591) <= not(layer4_outputs(3639));
    layer5_outputs(2592) <= (layer4_outputs(1578)) and not (layer4_outputs(1));
    layer5_outputs(2593) <= not(layer4_outputs(3307));
    layer5_outputs(2594) <= layer4_outputs(4777);
    layer5_outputs(2595) <= not((layer4_outputs(1402)) xor (layer4_outputs(495)));
    layer5_outputs(2596) <= not(layer4_outputs(218));
    layer5_outputs(2597) <= not(layer4_outputs(4697));
    layer5_outputs(2598) <= not((layer4_outputs(4002)) xor (layer4_outputs(1454)));
    layer5_outputs(2599) <= layer4_outputs(2068);
    layer5_outputs(2600) <= not(layer4_outputs(2165)) or (layer4_outputs(2819));
    layer5_outputs(2601) <= layer4_outputs(4109);
    layer5_outputs(2602) <= not(layer4_outputs(4739));
    layer5_outputs(2603) <= not(layer4_outputs(1980)) or (layer4_outputs(3851));
    layer5_outputs(2604) <= (layer4_outputs(796)) xor (layer4_outputs(2420));
    layer5_outputs(2605) <= (layer4_outputs(4562)) and not (layer4_outputs(2739));
    layer5_outputs(2606) <= layer4_outputs(779);
    layer5_outputs(2607) <= not(layer4_outputs(1748));
    layer5_outputs(2608) <= '1';
    layer5_outputs(2609) <= not(layer4_outputs(3428));
    layer5_outputs(2610) <= (layer4_outputs(241)) and (layer4_outputs(4837));
    layer5_outputs(2611) <= layer4_outputs(1736);
    layer5_outputs(2612) <= not(layer4_outputs(4690));
    layer5_outputs(2613) <= (layer4_outputs(5005)) and not (layer4_outputs(2986));
    layer5_outputs(2614) <= layer4_outputs(4565);
    layer5_outputs(2615) <= (layer4_outputs(3967)) and not (layer4_outputs(5084));
    layer5_outputs(2616) <= (layer4_outputs(4890)) and (layer4_outputs(856));
    layer5_outputs(2617) <= layer4_outputs(4074);
    layer5_outputs(2618) <= not((layer4_outputs(4183)) xor (layer4_outputs(4612)));
    layer5_outputs(2619) <= (layer4_outputs(1435)) and not (layer4_outputs(2750));
    layer5_outputs(2620) <= layer4_outputs(2353);
    layer5_outputs(2621) <= not(layer4_outputs(3409));
    layer5_outputs(2622) <= (layer4_outputs(3323)) and (layer4_outputs(216));
    layer5_outputs(2623) <= '1';
    layer5_outputs(2624) <= not((layer4_outputs(1285)) and (layer4_outputs(798)));
    layer5_outputs(2625) <= not(layer4_outputs(3586)) or (layer4_outputs(4479));
    layer5_outputs(2626) <= not(layer4_outputs(705));
    layer5_outputs(2627) <= not(layer4_outputs(2724));
    layer5_outputs(2628) <= layer4_outputs(4272);
    layer5_outputs(2629) <= not(layer4_outputs(36)) or (layer4_outputs(2770));
    layer5_outputs(2630) <= layer4_outputs(4201);
    layer5_outputs(2631) <= (layer4_outputs(2674)) xor (layer4_outputs(2218));
    layer5_outputs(2632) <= (layer4_outputs(2197)) or (layer4_outputs(3322));
    layer5_outputs(2633) <= not(layer4_outputs(3063)) or (layer4_outputs(2978));
    layer5_outputs(2634) <= (layer4_outputs(1135)) and not (layer4_outputs(3695));
    layer5_outputs(2635) <= (layer4_outputs(2943)) and not (layer4_outputs(1790));
    layer5_outputs(2636) <= layer4_outputs(3198);
    layer5_outputs(2637) <= layer4_outputs(4682);
    layer5_outputs(2638) <= (layer4_outputs(3124)) and (layer4_outputs(1438));
    layer5_outputs(2639) <= (layer4_outputs(730)) and not (layer4_outputs(1142));
    layer5_outputs(2640) <= not((layer4_outputs(2133)) xor (layer4_outputs(1182)));
    layer5_outputs(2641) <= layer4_outputs(1203);
    layer5_outputs(2642) <= layer4_outputs(2391);
    layer5_outputs(2643) <= (layer4_outputs(272)) xor (layer4_outputs(693));
    layer5_outputs(2644) <= layer4_outputs(552);
    layer5_outputs(2645) <= (layer4_outputs(3781)) and (layer4_outputs(677));
    layer5_outputs(2646) <= not(layer4_outputs(4107));
    layer5_outputs(2647) <= (layer4_outputs(1371)) or (layer4_outputs(1530));
    layer5_outputs(2648) <= '1';
    layer5_outputs(2649) <= layer4_outputs(1324);
    layer5_outputs(2650) <= (layer4_outputs(1605)) xor (layer4_outputs(2211));
    layer5_outputs(2651) <= (layer4_outputs(2953)) and not (layer4_outputs(582));
    layer5_outputs(2652) <= layer4_outputs(1716);
    layer5_outputs(2653) <= not(layer4_outputs(4141));
    layer5_outputs(2654) <= layer4_outputs(1058);
    layer5_outputs(2655) <= layer4_outputs(158);
    layer5_outputs(2656) <= not((layer4_outputs(1876)) xor (layer4_outputs(3933)));
    layer5_outputs(2657) <= not(layer4_outputs(647));
    layer5_outputs(2658) <= (layer4_outputs(2070)) or (layer4_outputs(35));
    layer5_outputs(2659) <= not(layer4_outputs(2195));
    layer5_outputs(2660) <= not(layer4_outputs(1362)) or (layer4_outputs(4414));
    layer5_outputs(2661) <= layer4_outputs(3863);
    layer5_outputs(2662) <= (layer4_outputs(171)) and (layer4_outputs(1753));
    layer5_outputs(2663) <= layer4_outputs(1558);
    layer5_outputs(2664) <= not(layer4_outputs(1607));
    layer5_outputs(2665) <= layer4_outputs(2087);
    layer5_outputs(2666) <= layer4_outputs(284);
    layer5_outputs(2667) <= not((layer4_outputs(1310)) and (layer4_outputs(4645)));
    layer5_outputs(2668) <= not((layer4_outputs(1032)) or (layer4_outputs(2619)));
    layer5_outputs(2669) <= (layer4_outputs(1648)) or (layer4_outputs(4613));
    layer5_outputs(2670) <= '1';
    layer5_outputs(2671) <= not(layer4_outputs(3750)) or (layer4_outputs(1017));
    layer5_outputs(2672) <= not(layer4_outputs(2271)) or (layer4_outputs(4701));
    layer5_outputs(2673) <= not(layer4_outputs(3957));
    layer5_outputs(2674) <= '0';
    layer5_outputs(2675) <= not((layer4_outputs(3092)) or (layer4_outputs(3088)));
    layer5_outputs(2676) <= not(layer4_outputs(2437));
    layer5_outputs(2677) <= not(layer4_outputs(5055));
    layer5_outputs(2678) <= (layer4_outputs(246)) xor (layer4_outputs(3206));
    layer5_outputs(2679) <= not((layer4_outputs(3573)) or (layer4_outputs(4893)));
    layer5_outputs(2680) <= (layer4_outputs(4671)) or (layer4_outputs(3262));
    layer5_outputs(2681) <= not((layer4_outputs(4981)) and (layer4_outputs(1683)));
    layer5_outputs(2682) <= not(layer4_outputs(1338)) or (layer4_outputs(941));
    layer5_outputs(2683) <= not(layer4_outputs(5027)) or (layer4_outputs(559));
    layer5_outputs(2684) <= not(layer4_outputs(3809));
    layer5_outputs(2685) <= not(layer4_outputs(3439));
    layer5_outputs(2686) <= layer4_outputs(1521);
    layer5_outputs(2687) <= not(layer4_outputs(3890)) or (layer4_outputs(847));
    layer5_outputs(2688) <= not(layer4_outputs(1807));
    layer5_outputs(2689) <= layer4_outputs(3313);
    layer5_outputs(2690) <= '0';
    layer5_outputs(2691) <= (layer4_outputs(1938)) or (layer4_outputs(3375));
    layer5_outputs(2692) <= layer4_outputs(192);
    layer5_outputs(2693) <= not((layer4_outputs(681)) xor (layer4_outputs(2413)));
    layer5_outputs(2694) <= not((layer4_outputs(3797)) and (layer4_outputs(4923)));
    layer5_outputs(2695) <= not((layer4_outputs(536)) or (layer4_outputs(4824)));
    layer5_outputs(2696) <= not(layer4_outputs(357));
    layer5_outputs(2697) <= (layer4_outputs(1142)) xor (layer4_outputs(3374));
    layer5_outputs(2698) <= not(layer4_outputs(1802)) or (layer4_outputs(1633));
    layer5_outputs(2699) <= (layer4_outputs(2500)) or (layer4_outputs(2054));
    layer5_outputs(2700) <= not(layer4_outputs(4787));
    layer5_outputs(2701) <= layer4_outputs(1389);
    layer5_outputs(2702) <= not(layer4_outputs(3156)) or (layer4_outputs(2057));
    layer5_outputs(2703) <= layer4_outputs(4468);
    layer5_outputs(2704) <= layer4_outputs(539);
    layer5_outputs(2705) <= layer4_outputs(2126);
    layer5_outputs(2706) <= not(layer4_outputs(1568)) or (layer4_outputs(2972));
    layer5_outputs(2707) <= '0';
    layer5_outputs(2708) <= '0';
    layer5_outputs(2709) <= not(layer4_outputs(269)) or (layer4_outputs(105));
    layer5_outputs(2710) <= (layer4_outputs(3112)) and not (layer4_outputs(1919));
    layer5_outputs(2711) <= not(layer4_outputs(1458));
    layer5_outputs(2712) <= not(layer4_outputs(2006));
    layer5_outputs(2713) <= not((layer4_outputs(3521)) and (layer4_outputs(3284)));
    layer5_outputs(2714) <= not((layer4_outputs(38)) or (layer4_outputs(4139)));
    layer5_outputs(2715) <= layer4_outputs(3364);
    layer5_outputs(2716) <= layer4_outputs(2271);
    layer5_outputs(2717) <= (layer4_outputs(3150)) and not (layer4_outputs(2849));
    layer5_outputs(2718) <= (layer4_outputs(2354)) and not (layer4_outputs(4789));
    layer5_outputs(2719) <= layer4_outputs(3774);
    layer5_outputs(2720) <= not((layer4_outputs(706)) xor (layer4_outputs(3766)));
    layer5_outputs(2721) <= not(layer4_outputs(3459)) or (layer4_outputs(1295));
    layer5_outputs(2722) <= layer4_outputs(4762);
    layer5_outputs(2723) <= not((layer4_outputs(2924)) and (layer4_outputs(2807)));
    layer5_outputs(2724) <= layer4_outputs(3387);
    layer5_outputs(2725) <= not(layer4_outputs(4861));
    layer5_outputs(2726) <= (layer4_outputs(3233)) or (layer4_outputs(54));
    layer5_outputs(2727) <= (layer4_outputs(2974)) and not (layer4_outputs(3608));
    layer5_outputs(2728) <= layer4_outputs(3803);
    layer5_outputs(2729) <= layer4_outputs(1339);
    layer5_outputs(2730) <= layer4_outputs(4461);
    layer5_outputs(2731) <= (layer4_outputs(533)) and not (layer4_outputs(3000));
    layer5_outputs(2732) <= (layer4_outputs(5046)) and (layer4_outputs(3123));
    layer5_outputs(2733) <= not(layer4_outputs(4780));
    layer5_outputs(2734) <= not((layer4_outputs(756)) or (layer4_outputs(4990)));
    layer5_outputs(2735) <= not(layer4_outputs(3440));
    layer5_outputs(2736) <= layer4_outputs(2689);
    layer5_outputs(2737) <= not(layer4_outputs(2050));
    layer5_outputs(2738) <= (layer4_outputs(4153)) and not (layer4_outputs(4530));
    layer5_outputs(2739) <= not(layer4_outputs(2821));
    layer5_outputs(2740) <= layer4_outputs(3216);
    layer5_outputs(2741) <= not(layer4_outputs(2292)) or (layer4_outputs(1740));
    layer5_outputs(2742) <= not(layer4_outputs(575));
    layer5_outputs(2743) <= not(layer4_outputs(827)) or (layer4_outputs(3146));
    layer5_outputs(2744) <= not((layer4_outputs(1758)) xor (layer4_outputs(1194)));
    layer5_outputs(2745) <= (layer4_outputs(15)) or (layer4_outputs(2603));
    layer5_outputs(2746) <= layer4_outputs(3237);
    layer5_outputs(2747) <= not(layer4_outputs(1845));
    layer5_outputs(2748) <= not(layer4_outputs(1222));
    layer5_outputs(2749) <= (layer4_outputs(1671)) and not (layer4_outputs(2884));
    layer5_outputs(2750) <= (layer4_outputs(381)) and not (layer4_outputs(2847));
    layer5_outputs(2751) <= (layer4_outputs(4620)) and not (layer4_outputs(1419));
    layer5_outputs(2752) <= (layer4_outputs(4915)) or (layer4_outputs(3610));
    layer5_outputs(2753) <= not((layer4_outputs(2725)) and (layer4_outputs(463)));
    layer5_outputs(2754) <= layer4_outputs(4113);
    layer5_outputs(2755) <= not(layer4_outputs(2041));
    layer5_outputs(2756) <= layer4_outputs(4169);
    layer5_outputs(2757) <= not(layer4_outputs(2205));
    layer5_outputs(2758) <= layer4_outputs(2107);
    layer5_outputs(2759) <= not((layer4_outputs(1121)) xor (layer4_outputs(2651)));
    layer5_outputs(2760) <= not(layer4_outputs(2879));
    layer5_outputs(2761) <= not(layer4_outputs(301)) or (layer4_outputs(3568));
    layer5_outputs(2762) <= (layer4_outputs(3045)) xor (layer4_outputs(1540));
    layer5_outputs(2763) <= not(layer4_outputs(4732));
    layer5_outputs(2764) <= (layer4_outputs(1733)) xor (layer4_outputs(4713));
    layer5_outputs(2765) <= not(layer4_outputs(2666)) or (layer4_outputs(3418));
    layer5_outputs(2766) <= layer4_outputs(1817);
    layer5_outputs(2767) <= (layer4_outputs(1103)) and not (layer4_outputs(2320));
    layer5_outputs(2768) <= (layer4_outputs(4455)) or (layer4_outputs(383));
    layer5_outputs(2769) <= not((layer4_outputs(4396)) xor (layer4_outputs(4807)));
    layer5_outputs(2770) <= layer4_outputs(2097);
    layer5_outputs(2771) <= not((layer4_outputs(1774)) or (layer4_outputs(2049)));
    layer5_outputs(2772) <= not(layer4_outputs(3725)) or (layer4_outputs(2402));
    layer5_outputs(2773) <= (layer4_outputs(4434)) and not (layer4_outputs(1704));
    layer5_outputs(2774) <= not(layer4_outputs(633));
    layer5_outputs(2775) <= not(layer4_outputs(3389)) or (layer4_outputs(1992));
    layer5_outputs(2776) <= (layer4_outputs(806)) and (layer4_outputs(1748));
    layer5_outputs(2777) <= not(layer4_outputs(3044)) or (layer4_outputs(681));
    layer5_outputs(2778) <= layer4_outputs(5073);
    layer5_outputs(2779) <= (layer4_outputs(3593)) xor (layer4_outputs(3748));
    layer5_outputs(2780) <= (layer4_outputs(1745)) and not (layer4_outputs(3920));
    layer5_outputs(2781) <= layer4_outputs(2237);
    layer5_outputs(2782) <= layer4_outputs(4240);
    layer5_outputs(2783) <= (layer4_outputs(1009)) xor (layer4_outputs(646));
    layer5_outputs(2784) <= layer4_outputs(2080);
    layer5_outputs(2785) <= not((layer4_outputs(4255)) xor (layer4_outputs(3785)));
    layer5_outputs(2786) <= (layer4_outputs(63)) and not (layer4_outputs(3602));
    layer5_outputs(2787) <= not((layer4_outputs(877)) or (layer4_outputs(1961)));
    layer5_outputs(2788) <= not(layer4_outputs(3782)) or (layer4_outputs(1957));
    layer5_outputs(2789) <= (layer4_outputs(1994)) xor (layer4_outputs(4013));
    layer5_outputs(2790) <= not(layer4_outputs(3741));
    layer5_outputs(2791) <= layer4_outputs(3878);
    layer5_outputs(2792) <= layer4_outputs(3686);
    layer5_outputs(2793) <= (layer4_outputs(3690)) xor (layer4_outputs(3058));
    layer5_outputs(2794) <= layer4_outputs(448);
    layer5_outputs(2795) <= layer4_outputs(3155);
    layer5_outputs(2796) <= not((layer4_outputs(4520)) and (layer4_outputs(2164)));
    layer5_outputs(2797) <= not((layer4_outputs(2863)) and (layer4_outputs(114)));
    layer5_outputs(2798) <= (layer4_outputs(18)) and not (layer4_outputs(2781));
    layer5_outputs(2799) <= not((layer4_outputs(237)) or (layer4_outputs(701)));
    layer5_outputs(2800) <= '1';
    layer5_outputs(2801) <= not(layer4_outputs(1293));
    layer5_outputs(2802) <= layer4_outputs(2324);
    layer5_outputs(2803) <= not(layer4_outputs(3912));
    layer5_outputs(2804) <= not((layer4_outputs(4464)) xor (layer4_outputs(3816)));
    layer5_outputs(2805) <= not((layer4_outputs(5029)) and (layer4_outputs(3488)));
    layer5_outputs(2806) <= not(layer4_outputs(4557));
    layer5_outputs(2807) <= layer4_outputs(2699);
    layer5_outputs(2808) <= not(layer4_outputs(4905));
    layer5_outputs(2809) <= (layer4_outputs(4080)) xor (layer4_outputs(1139));
    layer5_outputs(2810) <= layer4_outputs(1140);
    layer5_outputs(2811) <= not(layer4_outputs(76));
    layer5_outputs(2812) <= not(layer4_outputs(4793));
    layer5_outputs(2813) <= not((layer4_outputs(718)) or (layer4_outputs(4413)));
    layer5_outputs(2814) <= not((layer4_outputs(4874)) xor (layer4_outputs(457)));
    layer5_outputs(2815) <= (layer4_outputs(1351)) or (layer4_outputs(4072));
    layer5_outputs(2816) <= not(layer4_outputs(2797));
    layer5_outputs(2817) <= not((layer4_outputs(1202)) xor (layer4_outputs(219)));
    layer5_outputs(2818) <= (layer4_outputs(1669)) and not (layer4_outputs(1582));
    layer5_outputs(2819) <= not(layer4_outputs(4188));
    layer5_outputs(2820) <= layer4_outputs(3589);
    layer5_outputs(2821) <= (layer4_outputs(2920)) or (layer4_outputs(3183));
    layer5_outputs(2822) <= layer4_outputs(1598);
    layer5_outputs(2823) <= not(layer4_outputs(2164));
    layer5_outputs(2824) <= not(layer4_outputs(2914)) or (layer4_outputs(3435));
    layer5_outputs(2825) <= not(layer4_outputs(1264));
    layer5_outputs(2826) <= not(layer4_outputs(4238)) or (layer4_outputs(3870));
    layer5_outputs(2827) <= layer4_outputs(2262);
    layer5_outputs(2828) <= not(layer4_outputs(3594)) or (layer4_outputs(3237));
    layer5_outputs(2829) <= not(layer4_outputs(144));
    layer5_outputs(2830) <= not((layer4_outputs(4542)) xor (layer4_outputs(2347)));
    layer5_outputs(2831) <= layer4_outputs(3719);
    layer5_outputs(2832) <= layer4_outputs(99);
    layer5_outputs(2833) <= not(layer4_outputs(2740));
    layer5_outputs(2834) <= not((layer4_outputs(3351)) xor (layer4_outputs(4665)));
    layer5_outputs(2835) <= (layer4_outputs(5062)) and (layer4_outputs(4608));
    layer5_outputs(2836) <= layer4_outputs(2206);
    layer5_outputs(2837) <= not(layer4_outputs(2053));
    layer5_outputs(2838) <= not(layer4_outputs(96));
    layer5_outputs(2839) <= '0';
    layer5_outputs(2840) <= not(layer4_outputs(4920)) or (layer4_outputs(57));
    layer5_outputs(2841) <= not(layer4_outputs(2702));
    layer5_outputs(2842) <= layer4_outputs(2250);
    layer5_outputs(2843) <= '0';
    layer5_outputs(2844) <= layer4_outputs(2661);
    layer5_outputs(2845) <= not(layer4_outputs(4247));
    layer5_outputs(2846) <= layer4_outputs(631);
    layer5_outputs(2847) <= layer4_outputs(4672);
    layer5_outputs(2848) <= not(layer4_outputs(1792));
    layer5_outputs(2849) <= not((layer4_outputs(3775)) xor (layer4_outputs(500)));
    layer5_outputs(2850) <= not(layer4_outputs(4924));
    layer5_outputs(2851) <= layer4_outputs(2795);
    layer5_outputs(2852) <= layer4_outputs(295);
    layer5_outputs(2853) <= '0';
    layer5_outputs(2854) <= not(layer4_outputs(1240));
    layer5_outputs(2855) <= layer4_outputs(1680);
    layer5_outputs(2856) <= (layer4_outputs(1942)) xor (layer4_outputs(101));
    layer5_outputs(2857) <= layer4_outputs(3575);
    layer5_outputs(2858) <= not((layer4_outputs(2339)) and (layer4_outputs(1101)));
    layer5_outputs(2859) <= not((layer4_outputs(359)) or (layer4_outputs(1874)));
    layer5_outputs(2860) <= '1';
    layer5_outputs(2861) <= not(layer4_outputs(4485));
    layer5_outputs(2862) <= not(layer4_outputs(822));
    layer5_outputs(2863) <= not(layer4_outputs(2365));
    layer5_outputs(2864) <= not((layer4_outputs(398)) or (layer4_outputs(2592)));
    layer5_outputs(2865) <= layer4_outputs(2873);
    layer5_outputs(2866) <= layer4_outputs(573);
    layer5_outputs(2867) <= (layer4_outputs(1066)) and (layer4_outputs(3200));
    layer5_outputs(2868) <= not(layer4_outputs(2091));
    layer5_outputs(2869) <= not((layer4_outputs(266)) or (layer4_outputs(1810)));
    layer5_outputs(2870) <= not((layer4_outputs(3826)) xor (layer4_outputs(650)));
    layer5_outputs(2871) <= (layer4_outputs(2388)) and (layer4_outputs(4093));
    layer5_outputs(2872) <= layer4_outputs(4890);
    layer5_outputs(2873) <= not(layer4_outputs(3738));
    layer5_outputs(2874) <= not(layer4_outputs(769));
    layer5_outputs(2875) <= '0';
    layer5_outputs(2876) <= not((layer4_outputs(4569)) xor (layer4_outputs(3990)));
    layer5_outputs(2877) <= layer4_outputs(382);
    layer5_outputs(2878) <= not(layer4_outputs(4826));
    layer5_outputs(2879) <= layer4_outputs(1697);
    layer5_outputs(2880) <= not(layer4_outputs(809));
    layer5_outputs(2881) <= not((layer4_outputs(5030)) and (layer4_outputs(443)));
    layer5_outputs(2882) <= (layer4_outputs(3757)) or (layer4_outputs(3906));
    layer5_outputs(2883) <= layer4_outputs(3027);
    layer5_outputs(2884) <= (layer4_outputs(3563)) and (layer4_outputs(2185));
    layer5_outputs(2885) <= not(layer4_outputs(2901));
    layer5_outputs(2886) <= not((layer4_outputs(1954)) and (layer4_outputs(3482)));
    layer5_outputs(2887) <= (layer4_outputs(2723)) and (layer4_outputs(4064));
    layer5_outputs(2888) <= not(layer4_outputs(4922));
    layer5_outputs(2889) <= layer4_outputs(611);
    layer5_outputs(2890) <= not(layer4_outputs(3294));
    layer5_outputs(2891) <= not(layer4_outputs(1568)) or (layer4_outputs(750));
    layer5_outputs(2892) <= not(layer4_outputs(336)) or (layer4_outputs(168));
    layer5_outputs(2893) <= layer4_outputs(1524);
    layer5_outputs(2894) <= layer4_outputs(379);
    layer5_outputs(2895) <= layer4_outputs(1461);
    layer5_outputs(2896) <= not(layer4_outputs(4480));
    layer5_outputs(2897) <= not(layer4_outputs(4309));
    layer5_outputs(2898) <= (layer4_outputs(3626)) and not (layer4_outputs(1278));
    layer5_outputs(2899) <= (layer4_outputs(4419)) and (layer4_outputs(3070));
    layer5_outputs(2900) <= not(layer4_outputs(807));
    layer5_outputs(2901) <= layer4_outputs(2261);
    layer5_outputs(2902) <= not(layer4_outputs(408)) or (layer4_outputs(1006));
    layer5_outputs(2903) <= not((layer4_outputs(5011)) or (layer4_outputs(2297)));
    layer5_outputs(2904) <= not(layer4_outputs(351)) or (layer4_outputs(3436));
    layer5_outputs(2905) <= not((layer4_outputs(1410)) xor (layer4_outputs(1007)));
    layer5_outputs(2906) <= '1';
    layer5_outputs(2907) <= (layer4_outputs(3486)) and not (layer4_outputs(4489));
    layer5_outputs(2908) <= (layer4_outputs(1271)) and (layer4_outputs(1415));
    layer5_outputs(2909) <= not(layer4_outputs(1712)) or (layer4_outputs(3214));
    layer5_outputs(2910) <= not(layer4_outputs(1501));
    layer5_outputs(2911) <= (layer4_outputs(2847)) and (layer4_outputs(4975));
    layer5_outputs(2912) <= not(layer4_outputs(3968));
    layer5_outputs(2913) <= not(layer4_outputs(1498));
    layer5_outputs(2914) <= (layer4_outputs(660)) or (layer4_outputs(364));
    layer5_outputs(2915) <= layer4_outputs(537);
    layer5_outputs(2916) <= layer4_outputs(901);
    layer5_outputs(2917) <= (layer4_outputs(3109)) or (layer4_outputs(2971));
    layer5_outputs(2918) <= layer4_outputs(3112);
    layer5_outputs(2919) <= not(layer4_outputs(3976));
    layer5_outputs(2920) <= not(layer4_outputs(3332)) or (layer4_outputs(1194));
    layer5_outputs(2921) <= (layer4_outputs(256)) and not (layer4_outputs(1557));
    layer5_outputs(2922) <= not(layer4_outputs(2411));
    layer5_outputs(2923) <= not(layer4_outputs(3272));
    layer5_outputs(2924) <= layer4_outputs(206);
    layer5_outputs(2925) <= not(layer4_outputs(4292));
    layer5_outputs(2926) <= (layer4_outputs(4084)) xor (layer4_outputs(365));
    layer5_outputs(2927) <= (layer4_outputs(4825)) and not (layer4_outputs(1832));
    layer5_outputs(2928) <= '1';
    layer5_outputs(2929) <= '1';
    layer5_outputs(2930) <= not(layer4_outputs(1815));
    layer5_outputs(2931) <= not(layer4_outputs(1996));
    layer5_outputs(2932) <= not((layer4_outputs(5061)) xor (layer4_outputs(2848)));
    layer5_outputs(2933) <= not(layer4_outputs(2650));
    layer5_outputs(2934) <= not(layer4_outputs(4887));
    layer5_outputs(2935) <= layer4_outputs(3907);
    layer5_outputs(2936) <= layer4_outputs(341);
    layer5_outputs(2937) <= (layer4_outputs(777)) xor (layer4_outputs(2889));
    layer5_outputs(2938) <= layer4_outputs(3308);
    layer5_outputs(2939) <= (layer4_outputs(2923)) xor (layer4_outputs(4098));
    layer5_outputs(2940) <= not((layer4_outputs(1813)) or (layer4_outputs(4574)));
    layer5_outputs(2941) <= not(layer4_outputs(4548));
    layer5_outputs(2942) <= not((layer4_outputs(1616)) or (layer4_outputs(664)));
    layer5_outputs(2943) <= layer4_outputs(4135);
    layer5_outputs(2944) <= (layer4_outputs(3311)) or (layer4_outputs(1129));
    layer5_outputs(2945) <= not(layer4_outputs(1809)) or (layer4_outputs(3231));
    layer5_outputs(2946) <= not(layer4_outputs(3400));
    layer5_outputs(2947) <= not((layer4_outputs(877)) xor (layer4_outputs(1583)));
    layer5_outputs(2948) <= not((layer4_outputs(3375)) or (layer4_outputs(3278)));
    layer5_outputs(2949) <= not(layer4_outputs(513)) or (layer4_outputs(1813));
    layer5_outputs(2950) <= (layer4_outputs(546)) and not (layer4_outputs(3674));
    layer5_outputs(2951) <= '1';
    layer5_outputs(2952) <= (layer4_outputs(1780)) and (layer4_outputs(4932));
    layer5_outputs(2953) <= layer4_outputs(2052);
    layer5_outputs(2954) <= layer4_outputs(1511);
    layer5_outputs(2955) <= not(layer4_outputs(1900));
    layer5_outputs(2956) <= layer4_outputs(2515);
    layer5_outputs(2957) <= not(layer4_outputs(357));
    layer5_outputs(2958) <= (layer4_outputs(3394)) and not (layer4_outputs(1043));
    layer5_outputs(2959) <= not(layer4_outputs(1340));
    layer5_outputs(2960) <= not(layer4_outputs(3541));
    layer5_outputs(2961) <= not(layer4_outputs(4627));
    layer5_outputs(2962) <= layer4_outputs(2644);
    layer5_outputs(2963) <= (layer4_outputs(4447)) and (layer4_outputs(1899));
    layer5_outputs(2964) <= layer4_outputs(2898);
    layer5_outputs(2965) <= layer4_outputs(2556);
    layer5_outputs(2966) <= not((layer4_outputs(4938)) and (layer4_outputs(4078)));
    layer5_outputs(2967) <= '1';
    layer5_outputs(2968) <= not((layer4_outputs(4588)) and (layer4_outputs(3911)));
    layer5_outputs(2969) <= '1';
    layer5_outputs(2970) <= layer4_outputs(3105);
    layer5_outputs(2971) <= not((layer4_outputs(3477)) xor (layer4_outputs(3358)));
    layer5_outputs(2972) <= layer4_outputs(5051);
    layer5_outputs(2973) <= not(layer4_outputs(2606));
    layer5_outputs(2974) <= layer4_outputs(3318);
    layer5_outputs(2975) <= layer4_outputs(138);
    layer5_outputs(2976) <= not(layer4_outputs(4373));
    layer5_outputs(2977) <= not(layer4_outputs(1032));
    layer5_outputs(2978) <= (layer4_outputs(4667)) and not (layer4_outputs(3371));
    layer5_outputs(2979) <= not(layer4_outputs(3520)) or (layer4_outputs(2417));
    layer5_outputs(2980) <= (layer4_outputs(4476)) and not (layer4_outputs(324));
    layer5_outputs(2981) <= not(layer4_outputs(4445));
    layer5_outputs(2982) <= layer4_outputs(3170);
    layer5_outputs(2983) <= '0';
    layer5_outputs(2984) <= not(layer4_outputs(921));
    layer5_outputs(2985) <= not(layer4_outputs(698));
    layer5_outputs(2986) <= not(layer4_outputs(4466));
    layer5_outputs(2987) <= layer4_outputs(1514);
    layer5_outputs(2988) <= (layer4_outputs(4226)) and (layer4_outputs(3429));
    layer5_outputs(2989) <= not(layer4_outputs(1816));
    layer5_outputs(2990) <= layer4_outputs(1675);
    layer5_outputs(2991) <= (layer4_outputs(558)) and not (layer4_outputs(3474));
    layer5_outputs(2992) <= layer4_outputs(1236);
    layer5_outputs(2993) <= not((layer4_outputs(1167)) and (layer4_outputs(4712)));
    layer5_outputs(2994) <= layer4_outputs(2605);
    layer5_outputs(2995) <= layer4_outputs(3904);
    layer5_outputs(2996) <= layer4_outputs(5028);
    layer5_outputs(2997) <= not(layer4_outputs(152)) or (layer4_outputs(237));
    layer5_outputs(2998) <= not((layer4_outputs(2221)) or (layer4_outputs(1038)));
    layer5_outputs(2999) <= not((layer4_outputs(548)) or (layer4_outputs(3065)));
    layer5_outputs(3000) <= not(layer4_outputs(3170));
    layer5_outputs(3001) <= not((layer4_outputs(2793)) and (layer4_outputs(3538)));
    layer5_outputs(3002) <= layer4_outputs(345);
    layer5_outputs(3003) <= not(layer4_outputs(496));
    layer5_outputs(3004) <= (layer4_outputs(1141)) and not (layer4_outputs(1620));
    layer5_outputs(3005) <= not((layer4_outputs(1995)) xor (layer4_outputs(4796)));
    layer5_outputs(3006) <= not(layer4_outputs(3821));
    layer5_outputs(3007) <= layer4_outputs(4919);
    layer5_outputs(3008) <= not((layer4_outputs(1238)) xor (layer4_outputs(1626)));
    layer5_outputs(3009) <= (layer4_outputs(3655)) or (layer4_outputs(2264));
    layer5_outputs(3010) <= not(layer4_outputs(2683));
    layer5_outputs(3011) <= not((layer4_outputs(1940)) or (layer4_outputs(821)));
    layer5_outputs(3012) <= (layer4_outputs(819)) and (layer4_outputs(1854));
    layer5_outputs(3013) <= (layer4_outputs(4610)) and (layer4_outputs(4430));
    layer5_outputs(3014) <= not(layer4_outputs(4895));
    layer5_outputs(3015) <= not(layer4_outputs(1140)) or (layer4_outputs(2466));
    layer5_outputs(3016) <= not((layer4_outputs(4947)) and (layer4_outputs(3205)));
    layer5_outputs(3017) <= not((layer4_outputs(1147)) xor (layer4_outputs(3952)));
    layer5_outputs(3018) <= layer4_outputs(2371);
    layer5_outputs(3019) <= not(layer4_outputs(134));
    layer5_outputs(3020) <= not(layer4_outputs(2988)) or (layer4_outputs(2743));
    layer5_outputs(3021) <= (layer4_outputs(3832)) or (layer4_outputs(1795));
    layer5_outputs(3022) <= (layer4_outputs(2447)) and (layer4_outputs(2655));
    layer5_outputs(3023) <= not(layer4_outputs(2611)) or (layer4_outputs(3988));
    layer5_outputs(3024) <= not(layer4_outputs(1805));
    layer5_outputs(3025) <= layer4_outputs(1576);
    layer5_outputs(3026) <= layer4_outputs(3557);
    layer5_outputs(3027) <= (layer4_outputs(182)) and not (layer4_outputs(3336));
    layer5_outputs(3028) <= (layer4_outputs(4443)) and not (layer4_outputs(3715));
    layer5_outputs(3029) <= not(layer4_outputs(1233));
    layer5_outputs(3030) <= (layer4_outputs(4403)) xor (layer4_outputs(4671));
    layer5_outputs(3031) <= not(layer4_outputs(5110));
    layer5_outputs(3032) <= (layer4_outputs(2872)) and not (layer4_outputs(2912));
    layer5_outputs(3033) <= not((layer4_outputs(2363)) or (layer4_outputs(887)));
    layer5_outputs(3034) <= (layer4_outputs(1255)) and (layer4_outputs(4526));
    layer5_outputs(3035) <= not(layer4_outputs(1420));
    layer5_outputs(3036) <= not(layer4_outputs(3506));
    layer5_outputs(3037) <= (layer4_outputs(4180)) and not (layer4_outputs(4381));
    layer5_outputs(3038) <= (layer4_outputs(3570)) and not (layer4_outputs(1048));
    layer5_outputs(3039) <= layer4_outputs(4087);
    layer5_outputs(3040) <= not(layer4_outputs(2445));
    layer5_outputs(3041) <= not(layer4_outputs(2495));
    layer5_outputs(3042) <= not(layer4_outputs(4471));
    layer5_outputs(3043) <= not(layer4_outputs(4205));
    layer5_outputs(3044) <= (layer4_outputs(4063)) and (layer4_outputs(2520));
    layer5_outputs(3045) <= not(layer4_outputs(3166));
    layer5_outputs(3046) <= layer4_outputs(3419);
    layer5_outputs(3047) <= not(layer4_outputs(521));
    layer5_outputs(3048) <= layer4_outputs(4377);
    layer5_outputs(3049) <= not(layer4_outputs(4119));
    layer5_outputs(3050) <= '1';
    layer5_outputs(3051) <= not((layer4_outputs(852)) or (layer4_outputs(599)));
    layer5_outputs(3052) <= layer4_outputs(4737);
    layer5_outputs(3053) <= not((layer4_outputs(655)) xor (layer4_outputs(2383)));
    layer5_outputs(3054) <= not((layer4_outputs(1116)) or (layer4_outputs(4074)));
    layer5_outputs(3055) <= not(layer4_outputs(918)) or (layer4_outputs(2969));
    layer5_outputs(3056) <= '0';
    layer5_outputs(3057) <= not(layer4_outputs(1221)) or (layer4_outputs(3206));
    layer5_outputs(3058) <= (layer4_outputs(4034)) and not (layer4_outputs(4604));
    layer5_outputs(3059) <= layer4_outputs(4645);
    layer5_outputs(3060) <= not((layer4_outputs(4483)) and (layer4_outputs(1481)));
    layer5_outputs(3061) <= (layer4_outputs(1652)) and not (layer4_outputs(325));
    layer5_outputs(3062) <= not(layer4_outputs(4208));
    layer5_outputs(3063) <= not(layer4_outputs(1014));
    layer5_outputs(3064) <= not((layer4_outputs(4688)) or (layer4_outputs(2747)));
    layer5_outputs(3065) <= layer4_outputs(5051);
    layer5_outputs(3066) <= not(layer4_outputs(1530)) or (layer4_outputs(33));
    layer5_outputs(3067) <= (layer4_outputs(988)) and not (layer4_outputs(4430));
    layer5_outputs(3068) <= not(layer4_outputs(407)) or (layer4_outputs(953));
    layer5_outputs(3069) <= not(layer4_outputs(1121));
    layer5_outputs(3070) <= layer4_outputs(264);
    layer5_outputs(3071) <= not((layer4_outputs(5066)) and (layer4_outputs(2626)));
    layer5_outputs(3072) <= not(layer4_outputs(2601));
    layer5_outputs(3073) <= layer4_outputs(2504);
    layer5_outputs(3074) <= not(layer4_outputs(4215));
    layer5_outputs(3075) <= layer4_outputs(380);
    layer5_outputs(3076) <= layer4_outputs(4036);
    layer5_outputs(3077) <= not(layer4_outputs(392)) or (layer4_outputs(2154));
    layer5_outputs(3078) <= layer4_outputs(1197);
    layer5_outputs(3079) <= layer4_outputs(1694);
    layer5_outputs(3080) <= not((layer4_outputs(4835)) or (layer4_outputs(4018)));
    layer5_outputs(3081) <= layer4_outputs(3090);
    layer5_outputs(3082) <= not(layer4_outputs(1570)) or (layer4_outputs(4999));
    layer5_outputs(3083) <= not(layer4_outputs(1595));
    layer5_outputs(3084) <= not((layer4_outputs(2434)) or (layer4_outputs(277)));
    layer5_outputs(3085) <= not((layer4_outputs(4111)) xor (layer4_outputs(3732)));
    layer5_outputs(3086) <= (layer4_outputs(2494)) or (layer4_outputs(247));
    layer5_outputs(3087) <= layer4_outputs(3148);
    layer5_outputs(3088) <= not(layer4_outputs(3421));
    layer5_outputs(3089) <= layer4_outputs(1968);
    layer5_outputs(3090) <= layer4_outputs(680);
    layer5_outputs(3091) <= not(layer4_outputs(4418));
    layer5_outputs(3092) <= layer4_outputs(3797);
    layer5_outputs(3093) <= layer4_outputs(3232);
    layer5_outputs(3094) <= '1';
    layer5_outputs(3095) <= (layer4_outputs(666)) or (layer4_outputs(3277));
    layer5_outputs(3096) <= not(layer4_outputs(4603));
    layer5_outputs(3097) <= not(layer4_outputs(2057));
    layer5_outputs(3098) <= not(layer4_outputs(27));
    layer5_outputs(3099) <= not(layer4_outputs(2383));
    layer5_outputs(3100) <= layer4_outputs(4203);
    layer5_outputs(3101) <= not(layer4_outputs(4648));
    layer5_outputs(3102) <= layer4_outputs(224);
    layer5_outputs(3103) <= not(layer4_outputs(2658));
    layer5_outputs(3104) <= not(layer4_outputs(4391)) or (layer4_outputs(2463));
    layer5_outputs(3105) <= not(layer4_outputs(3187));
    layer5_outputs(3106) <= (layer4_outputs(3349)) or (layer4_outputs(1403));
    layer5_outputs(3107) <= not(layer4_outputs(1639)) or (layer4_outputs(4023));
    layer5_outputs(3108) <= (layer4_outputs(735)) and not (layer4_outputs(1317));
    layer5_outputs(3109) <= layer4_outputs(4672);
    layer5_outputs(3110) <= not(layer4_outputs(3023));
    layer5_outputs(3111) <= layer4_outputs(21);
    layer5_outputs(3112) <= '0';
    layer5_outputs(3113) <= layer4_outputs(1192);
    layer5_outputs(3114) <= not(layer4_outputs(3875)) or (layer4_outputs(3449));
    layer5_outputs(3115) <= layer4_outputs(4528);
    layer5_outputs(3116) <= (layer4_outputs(3470)) xor (layer4_outputs(384));
    layer5_outputs(3117) <= (layer4_outputs(5091)) and (layer4_outputs(2344));
    layer5_outputs(3118) <= not(layer4_outputs(1280));
    layer5_outputs(3119) <= layer4_outputs(3345);
    layer5_outputs(3120) <= '1';
    layer5_outputs(3121) <= layer4_outputs(3288);
    layer5_outputs(3122) <= '1';
    layer5_outputs(3123) <= not((layer4_outputs(704)) xor (layer4_outputs(510)));
    layer5_outputs(3124) <= not(layer4_outputs(4899));
    layer5_outputs(3125) <= layer4_outputs(4846);
    layer5_outputs(3126) <= not((layer4_outputs(3911)) and (layer4_outputs(1356)));
    layer5_outputs(3127) <= (layer4_outputs(2689)) and not (layer4_outputs(886));
    layer5_outputs(3128) <= not(layer4_outputs(2763)) or (layer4_outputs(3098));
    layer5_outputs(3129) <= not(layer4_outputs(1594));
    layer5_outputs(3130) <= layer4_outputs(2506);
    layer5_outputs(3131) <= not((layer4_outputs(251)) xor (layer4_outputs(3577)));
    layer5_outputs(3132) <= not(layer4_outputs(2375));
    layer5_outputs(3133) <= (layer4_outputs(1164)) or (layer4_outputs(2077));
    layer5_outputs(3134) <= (layer4_outputs(4408)) and not (layer4_outputs(879));
    layer5_outputs(3135) <= not(layer4_outputs(2039)) or (layer4_outputs(4975));
    layer5_outputs(3136) <= not(layer4_outputs(799));
    layer5_outputs(3137) <= not((layer4_outputs(4071)) or (layer4_outputs(3483)));
    layer5_outputs(3138) <= not(layer4_outputs(2374));
    layer5_outputs(3139) <= layer4_outputs(2834);
    layer5_outputs(3140) <= not((layer4_outputs(4761)) and (layer4_outputs(4144)));
    layer5_outputs(3141) <= (layer4_outputs(4491)) and (layer4_outputs(2815));
    layer5_outputs(3142) <= (layer4_outputs(4893)) or (layer4_outputs(1431));
    layer5_outputs(3143) <= (layer4_outputs(3303)) and not (layer4_outputs(567));
    layer5_outputs(3144) <= not(layer4_outputs(2704));
    layer5_outputs(3145) <= not((layer4_outputs(3632)) xor (layer4_outputs(4301)));
    layer5_outputs(3146) <= layer4_outputs(1428);
    layer5_outputs(3147) <= (layer4_outputs(858)) and (layer4_outputs(2440));
    layer5_outputs(3148) <= layer4_outputs(223);
    layer5_outputs(3149) <= not((layer4_outputs(2672)) and (layer4_outputs(2229)));
    layer5_outputs(3150) <= not((layer4_outputs(230)) xor (layer4_outputs(2919)));
    layer5_outputs(3151) <= not((layer4_outputs(1826)) and (layer4_outputs(3446)));
    layer5_outputs(3152) <= (layer4_outputs(2806)) xor (layer4_outputs(4164));
    layer5_outputs(3153) <= not(layer4_outputs(758));
    layer5_outputs(3154) <= '1';
    layer5_outputs(3155) <= layer4_outputs(3089);
    layer5_outputs(3156) <= not((layer4_outputs(3133)) and (layer4_outputs(3684)));
    layer5_outputs(3157) <= layer4_outputs(2905);
    layer5_outputs(3158) <= not(layer4_outputs(3250)) or (layer4_outputs(4891));
    layer5_outputs(3159) <= not(layer4_outputs(2823));
    layer5_outputs(3160) <= '0';
    layer5_outputs(3161) <= not(layer4_outputs(3828));
    layer5_outputs(3162) <= layer4_outputs(676);
    layer5_outputs(3163) <= '1';
    layer5_outputs(3164) <= layer4_outputs(1896);
    layer5_outputs(3165) <= layer4_outputs(3239);
    layer5_outputs(3166) <= not((layer4_outputs(4599)) xor (layer4_outputs(2077)));
    layer5_outputs(3167) <= layer4_outputs(4654);
    layer5_outputs(3168) <= layer4_outputs(4285);
    layer5_outputs(3169) <= not(layer4_outputs(2084));
    layer5_outputs(3170) <= not(layer4_outputs(3628)) or (layer4_outputs(2832));
    layer5_outputs(3171) <= not((layer4_outputs(88)) and (layer4_outputs(2504)));
    layer5_outputs(3172) <= not(layer4_outputs(3777));
    layer5_outputs(3173) <= not(layer4_outputs(4401));
    layer5_outputs(3174) <= not((layer4_outputs(2031)) or (layer4_outputs(2214)));
    layer5_outputs(3175) <= not(layer4_outputs(2137)) or (layer4_outputs(3400));
    layer5_outputs(3176) <= not(layer4_outputs(4395)) or (layer4_outputs(1624));
    layer5_outputs(3177) <= '1';
    layer5_outputs(3178) <= not((layer4_outputs(1309)) and (layer4_outputs(2595)));
    layer5_outputs(3179) <= (layer4_outputs(3325)) and not (layer4_outputs(3791));
    layer5_outputs(3180) <= layer4_outputs(4933);
    layer5_outputs(3181) <= not((layer4_outputs(826)) or (layer4_outputs(452)));
    layer5_outputs(3182) <= not(layer4_outputs(3444)) or (layer4_outputs(2858));
    layer5_outputs(3183) <= not(layer4_outputs(554));
    layer5_outputs(3184) <= not((layer4_outputs(4094)) or (layer4_outputs(122)));
    layer5_outputs(3185) <= not((layer4_outputs(2314)) xor (layer4_outputs(3631)));
    layer5_outputs(3186) <= not((layer4_outputs(3691)) xor (layer4_outputs(58)));
    layer5_outputs(3187) <= (layer4_outputs(4434)) or (layer4_outputs(3784));
    layer5_outputs(3188) <= (layer4_outputs(2949)) xor (layer4_outputs(4516));
    layer5_outputs(3189) <= not(layer4_outputs(1013));
    layer5_outputs(3190) <= (layer4_outputs(3496)) xor (layer4_outputs(304));
    layer5_outputs(3191) <= not(layer4_outputs(4097));
    layer5_outputs(3192) <= not((layer4_outputs(2750)) and (layer4_outputs(2434)));
    layer5_outputs(3193) <= not((layer4_outputs(4895)) or (layer4_outputs(3706)));
    layer5_outputs(3194) <= not(layer4_outputs(4855)) or (layer4_outputs(4005));
    layer5_outputs(3195) <= '0';
    layer5_outputs(3196) <= not(layer4_outputs(4063));
    layer5_outputs(3197) <= not(layer4_outputs(4885));
    layer5_outputs(3198) <= not((layer4_outputs(2303)) and (layer4_outputs(3982)));
    layer5_outputs(3199) <= layer4_outputs(1063);
    layer5_outputs(3200) <= not(layer4_outputs(4914)) or (layer4_outputs(117));
    layer5_outputs(3201) <= not(layer4_outputs(4046)) or (layer4_outputs(3833));
    layer5_outputs(3202) <= '0';
    layer5_outputs(3203) <= (layer4_outputs(2869)) and not (layer4_outputs(3782));
    layer5_outputs(3204) <= '0';
    layer5_outputs(3205) <= not(layer4_outputs(4935)) or (layer4_outputs(4022));
    layer5_outputs(3206) <= layer4_outputs(866);
    layer5_outputs(3207) <= not((layer4_outputs(1502)) and (layer4_outputs(1342)));
    layer5_outputs(3208) <= not(layer4_outputs(355));
    layer5_outputs(3209) <= layer4_outputs(4664);
    layer5_outputs(3210) <= (layer4_outputs(2842)) xor (layer4_outputs(891));
    layer5_outputs(3211) <= not(layer4_outputs(3960));
    layer5_outputs(3212) <= not((layer4_outputs(512)) and (layer4_outputs(2621)));
    layer5_outputs(3213) <= not(layer4_outputs(3919));
    layer5_outputs(3214) <= not(layer4_outputs(475)) or (layer4_outputs(3248));
    layer5_outputs(3215) <= (layer4_outputs(1453)) and not (layer4_outputs(80));
    layer5_outputs(3216) <= layer4_outputs(732);
    layer5_outputs(3217) <= not((layer4_outputs(2732)) or (layer4_outputs(3404)));
    layer5_outputs(3218) <= layer4_outputs(4319);
    layer5_outputs(3219) <= not(layer4_outputs(288)) or (layer4_outputs(454));
    layer5_outputs(3220) <= not((layer4_outputs(813)) and (layer4_outputs(991)));
    layer5_outputs(3221) <= '0';
    layer5_outputs(3222) <= layer4_outputs(1792);
    layer5_outputs(3223) <= (layer4_outputs(4675)) or (layer4_outputs(1891));
    layer5_outputs(3224) <= '0';
    layer5_outputs(3225) <= layer4_outputs(793);
    layer5_outputs(3226) <= layer4_outputs(2161);
    layer5_outputs(3227) <= layer4_outputs(1333);
    layer5_outputs(3228) <= not((layer4_outputs(2003)) xor (layer4_outputs(600)));
    layer5_outputs(3229) <= layer4_outputs(1449);
    layer5_outputs(3230) <= (layer4_outputs(2306)) or (layer4_outputs(1963));
    layer5_outputs(3231) <= not(layer4_outputs(1672));
    layer5_outputs(3232) <= not(layer4_outputs(321)) or (layer4_outputs(5072));
    layer5_outputs(3233) <= not(layer4_outputs(834)) or (layer4_outputs(1714));
    layer5_outputs(3234) <= not(layer4_outputs(439)) or (layer4_outputs(1254));
    layer5_outputs(3235) <= not(layer4_outputs(1727));
    layer5_outputs(3236) <= layer4_outputs(2248);
    layer5_outputs(3237) <= (layer4_outputs(4741)) or (layer4_outputs(2147));
    layer5_outputs(3238) <= not((layer4_outputs(4780)) or (layer4_outputs(1495)));
    layer5_outputs(3239) <= not(layer4_outputs(2452)) or (layer4_outputs(2829));
    layer5_outputs(3240) <= layer4_outputs(3322);
    layer5_outputs(3241) <= (layer4_outputs(340)) and (layer4_outputs(1950));
    layer5_outputs(3242) <= not(layer4_outputs(1539));
    layer5_outputs(3243) <= not((layer4_outputs(4812)) and (layer4_outputs(2701)));
    layer5_outputs(3244) <= (layer4_outputs(3117)) and not (layer4_outputs(903));
    layer5_outputs(3245) <= (layer4_outputs(1271)) and not (layer4_outputs(143));
    layer5_outputs(3246) <= not(layer4_outputs(472));
    layer5_outputs(3247) <= not(layer4_outputs(1008));
    layer5_outputs(3248) <= (layer4_outputs(853)) and not (layer4_outputs(1846));
    layer5_outputs(3249) <= not(layer4_outputs(4950)) or (layer4_outputs(14));
    layer5_outputs(3250) <= not(layer4_outputs(4290)) or (layer4_outputs(153));
    layer5_outputs(3251) <= (layer4_outputs(759)) xor (layer4_outputs(4906));
    layer5_outputs(3252) <= not(layer4_outputs(3102));
    layer5_outputs(3253) <= not(layer4_outputs(4319));
    layer5_outputs(3254) <= '0';
    layer5_outputs(3255) <= (layer4_outputs(1258)) xor (layer4_outputs(5060));
    layer5_outputs(3256) <= not(layer4_outputs(306));
    layer5_outputs(3257) <= not(layer4_outputs(198));
    layer5_outputs(3258) <= layer4_outputs(2508);
    layer5_outputs(3259) <= not(layer4_outputs(305));
    layer5_outputs(3260) <= layer4_outputs(3986);
    layer5_outputs(3261) <= not(layer4_outputs(4038));
    layer5_outputs(3262) <= '0';
    layer5_outputs(3263) <= '0';
    layer5_outputs(3264) <= not((layer4_outputs(911)) or (layer4_outputs(133)));
    layer5_outputs(3265) <= not(layer4_outputs(2532));
    layer5_outputs(3266) <= not(layer4_outputs(687));
    layer5_outputs(3267) <= (layer4_outputs(150)) and (layer4_outputs(3718));
    layer5_outputs(3268) <= (layer4_outputs(3007)) and not (layer4_outputs(2403));
    layer5_outputs(3269) <= (layer4_outputs(2691)) or (layer4_outputs(1671));
    layer5_outputs(3270) <= not(layer4_outputs(3464));
    layer5_outputs(3271) <= layer4_outputs(3716);
    layer5_outputs(3272) <= (layer4_outputs(2123)) xor (layer4_outputs(2254));
    layer5_outputs(3273) <= not(layer4_outputs(4987)) or (layer4_outputs(219));
    layer5_outputs(3274) <= not((layer4_outputs(1276)) xor (layer4_outputs(4440)));
    layer5_outputs(3275) <= layer4_outputs(2330);
    layer5_outputs(3276) <= not(layer4_outputs(1835)) or (layer4_outputs(3158));
    layer5_outputs(3277) <= layer4_outputs(445);
    layer5_outputs(3278) <= not(layer4_outputs(1619));
    layer5_outputs(3279) <= not((layer4_outputs(1640)) and (layer4_outputs(2025)));
    layer5_outputs(3280) <= not(layer4_outputs(5045)) or (layer4_outputs(2531));
    layer5_outputs(3281) <= (layer4_outputs(2836)) xor (layer4_outputs(914));
    layer5_outputs(3282) <= not(layer4_outputs(890)) or (layer4_outputs(3689));
    layer5_outputs(3283) <= layer4_outputs(2705);
    layer5_outputs(3284) <= layer4_outputs(3953);
    layer5_outputs(3285) <= not(layer4_outputs(1552));
    layer5_outputs(3286) <= layer4_outputs(4653);
    layer5_outputs(3287) <= layer4_outputs(908);
    layer5_outputs(3288) <= layer4_outputs(2871);
    layer5_outputs(3289) <= (layer4_outputs(1742)) xor (layer4_outputs(1243));
    layer5_outputs(3290) <= '1';
    layer5_outputs(3291) <= layer4_outputs(3393);
    layer5_outputs(3292) <= layer4_outputs(418);
    layer5_outputs(3293) <= not(layer4_outputs(173)) or (layer4_outputs(199));
    layer5_outputs(3294) <= not(layer4_outputs(3530));
    layer5_outputs(3295) <= not(layer4_outputs(3699));
    layer5_outputs(3296) <= layer4_outputs(2227);
    layer5_outputs(3297) <= not(layer4_outputs(2984));
    layer5_outputs(3298) <= not(layer4_outputs(1298));
    layer5_outputs(3299) <= layer4_outputs(1223);
    layer5_outputs(3300) <= layer4_outputs(4144);
    layer5_outputs(3301) <= layer4_outputs(1719);
    layer5_outputs(3302) <= '0';
    layer5_outputs(3303) <= (layer4_outputs(2259)) and not (layer4_outputs(2756));
    layer5_outputs(3304) <= (layer4_outputs(367)) and not (layer4_outputs(1240));
    layer5_outputs(3305) <= not(layer4_outputs(1644));
    layer5_outputs(3306) <= not((layer4_outputs(3555)) xor (layer4_outputs(173)));
    layer5_outputs(3307) <= (layer4_outputs(1918)) and not (layer4_outputs(2053));
    layer5_outputs(3308) <= not(layer4_outputs(3438));
    layer5_outputs(3309) <= not(layer4_outputs(3593));
    layer5_outputs(3310) <= layer4_outputs(3636);
    layer5_outputs(3311) <= '0';
    layer5_outputs(3312) <= (layer4_outputs(4003)) xor (layer4_outputs(260));
    layer5_outputs(3313) <= not(layer4_outputs(3730));
    layer5_outputs(3314) <= layer4_outputs(792);
    layer5_outputs(3315) <= '1';
    layer5_outputs(3316) <= layer4_outputs(1663);
    layer5_outputs(3317) <= not(layer4_outputs(750)) or (layer4_outputs(5107));
    layer5_outputs(3318) <= not(layer4_outputs(1506));
    layer5_outputs(3319) <= layer4_outputs(4765);
    layer5_outputs(3320) <= layer4_outputs(3560);
    layer5_outputs(3321) <= (layer4_outputs(3242)) and not (layer4_outputs(3103));
    layer5_outputs(3322) <= (layer4_outputs(1445)) or (layer4_outputs(1348));
    layer5_outputs(3323) <= layer4_outputs(4385);
    layer5_outputs(3324) <= not(layer4_outputs(987));
    layer5_outputs(3325) <= not(layer4_outputs(1668));
    layer5_outputs(3326) <= (layer4_outputs(3377)) xor (layer4_outputs(0));
    layer5_outputs(3327) <= layer4_outputs(3335);
    layer5_outputs(3328) <= not(layer4_outputs(1186));
    layer5_outputs(3329) <= (layer4_outputs(829)) and not (layer4_outputs(2257));
    layer5_outputs(3330) <= '1';
    layer5_outputs(3331) <= layer4_outputs(3222);
    layer5_outputs(3332) <= layer4_outputs(3729);
    layer5_outputs(3333) <= '0';
    layer5_outputs(3334) <= not(layer4_outputs(2140));
    layer5_outputs(3335) <= layer4_outputs(4577);
    layer5_outputs(3336) <= not((layer4_outputs(2602)) xor (layer4_outputs(2101)));
    layer5_outputs(3337) <= layer4_outputs(4777);
    layer5_outputs(3338) <= not(layer4_outputs(2854)) or (layer4_outputs(2472));
    layer5_outputs(3339) <= layer4_outputs(3856);
    layer5_outputs(3340) <= (layer4_outputs(189)) and (layer4_outputs(846));
    layer5_outputs(3341) <= not(layer4_outputs(3745)) or (layer4_outputs(1772));
    layer5_outputs(3342) <= (layer4_outputs(974)) and not (layer4_outputs(2777));
    layer5_outputs(3343) <= not(layer4_outputs(4369));
    layer5_outputs(3344) <= not(layer4_outputs(4930));
    layer5_outputs(3345) <= '0';
    layer5_outputs(3346) <= layer4_outputs(4197);
    layer5_outputs(3347) <= layer4_outputs(274);
    layer5_outputs(3348) <= (layer4_outputs(253)) or (layer4_outputs(1998));
    layer5_outputs(3349) <= (layer4_outputs(3218)) and (layer4_outputs(2589));
    layer5_outputs(3350) <= not(layer4_outputs(5023));
    layer5_outputs(3351) <= not(layer4_outputs(4610));
    layer5_outputs(3352) <= (layer4_outputs(3659)) and not (layer4_outputs(1569));
    layer5_outputs(3353) <= not(layer4_outputs(1021));
    layer5_outputs(3354) <= layer4_outputs(2944);
    layer5_outputs(3355) <= '1';
    layer5_outputs(3356) <= not(layer4_outputs(2267));
    layer5_outputs(3357) <= layer4_outputs(2208);
    layer5_outputs(3358) <= not(layer4_outputs(2985));
    layer5_outputs(3359) <= (layer4_outputs(3518)) or (layer4_outputs(4489));
    layer5_outputs(3360) <= (layer4_outputs(4453)) and not (layer4_outputs(2221));
    layer5_outputs(3361) <= not(layer4_outputs(3228));
    layer5_outputs(3362) <= not(layer4_outputs(4746)) or (layer4_outputs(3639));
    layer5_outputs(3363) <= not(layer4_outputs(639)) or (layer4_outputs(2966));
    layer5_outputs(3364) <= (layer4_outputs(1807)) xor (layer4_outputs(4008));
    layer5_outputs(3365) <= not((layer4_outputs(3626)) or (layer4_outputs(2699)));
    layer5_outputs(3366) <= layer4_outputs(2110);
    layer5_outputs(3367) <= not(layer4_outputs(4535));
    layer5_outputs(3368) <= not(layer4_outputs(3733));
    layer5_outputs(3369) <= layer4_outputs(1777);
    layer5_outputs(3370) <= not(layer4_outputs(4174)) or (layer4_outputs(837));
    layer5_outputs(3371) <= (layer4_outputs(4179)) and not (layer4_outputs(4556));
    layer5_outputs(3372) <= not((layer4_outputs(3720)) or (layer4_outputs(1878)));
    layer5_outputs(3373) <= not(layer4_outputs(3772)) or (layer4_outputs(4590));
    layer5_outputs(3374) <= layer4_outputs(3034);
    layer5_outputs(3375) <= (layer4_outputs(77)) xor (layer4_outputs(3969));
    layer5_outputs(3376) <= (layer4_outputs(4716)) and (layer4_outputs(1506));
    layer5_outputs(3377) <= layer4_outputs(1057);
    layer5_outputs(3378) <= not(layer4_outputs(535));
    layer5_outputs(3379) <= (layer4_outputs(1649)) and not (layer4_outputs(1579));
    layer5_outputs(3380) <= (layer4_outputs(2024)) and not (layer4_outputs(169));
    layer5_outputs(3381) <= layer4_outputs(1254);
    layer5_outputs(3382) <= not(layer4_outputs(3498));
    layer5_outputs(3383) <= not(layer4_outputs(3759));
    layer5_outputs(3384) <= (layer4_outputs(339)) and not (layer4_outputs(4121));
    layer5_outputs(3385) <= not((layer4_outputs(5099)) or (layer4_outputs(1046)));
    layer5_outputs(3386) <= not(layer4_outputs(3427));
    layer5_outputs(3387) <= not((layer4_outputs(464)) xor (layer4_outputs(1001)));
    layer5_outputs(3388) <= layer4_outputs(1008);
    layer5_outputs(3389) <= not((layer4_outputs(638)) or (layer4_outputs(3757)));
    layer5_outputs(3390) <= (layer4_outputs(3623)) and (layer4_outputs(2339));
    layer5_outputs(3391) <= not(layer4_outputs(4397)) or (layer4_outputs(4691));
    layer5_outputs(3392) <= layer4_outputs(1923);
    layer5_outputs(3393) <= layer4_outputs(2815);
    layer5_outputs(3394) <= layer4_outputs(3719);
    layer5_outputs(3395) <= not(layer4_outputs(44));
    layer5_outputs(3396) <= layer4_outputs(4642);
    layer5_outputs(3397) <= not(layer4_outputs(2758));
    layer5_outputs(3398) <= '1';
    layer5_outputs(3399) <= not(layer4_outputs(4393));
    layer5_outputs(3400) <= layer4_outputs(5119);
    layer5_outputs(3401) <= not((layer4_outputs(2436)) xor (layer4_outputs(4634)));
    layer5_outputs(3402) <= (layer4_outputs(4853)) and not (layer4_outputs(4270));
    layer5_outputs(3403) <= not(layer4_outputs(4667));
    layer5_outputs(3404) <= layer4_outputs(4258);
    layer5_outputs(3405) <= (layer4_outputs(3154)) and (layer4_outputs(3320));
    layer5_outputs(3406) <= not(layer4_outputs(947));
    layer5_outputs(3407) <= layer4_outputs(966);
    layer5_outputs(3408) <= layer4_outputs(2879);
    layer5_outputs(3409) <= layer4_outputs(2185);
    layer5_outputs(3410) <= not(layer4_outputs(1939));
    layer5_outputs(3411) <= (layer4_outputs(3343)) or (layer4_outputs(2040));
    layer5_outputs(3412) <= not(layer4_outputs(3499)) or (layer4_outputs(1075));
    layer5_outputs(3413) <= (layer4_outputs(3006)) and (layer4_outputs(3207));
    layer5_outputs(3414) <= layer4_outputs(1903);
    layer5_outputs(3415) <= layer4_outputs(2579);
    layer5_outputs(3416) <= (layer4_outputs(2142)) or (layer4_outputs(4532));
    layer5_outputs(3417) <= (layer4_outputs(4700)) xor (layer4_outputs(753));
    layer5_outputs(3418) <= (layer4_outputs(4731)) and not (layer4_outputs(2223));
    layer5_outputs(3419) <= layer4_outputs(1593);
    layer5_outputs(3420) <= layer4_outputs(2506);
    layer5_outputs(3421) <= (layer4_outputs(4219)) and not (layer4_outputs(714));
    layer5_outputs(3422) <= not((layer4_outputs(4392)) and (layer4_outputs(2546)));
    layer5_outputs(3423) <= layer4_outputs(3383);
    layer5_outputs(3424) <= layer4_outputs(3501);
    layer5_outputs(3425) <= (layer4_outputs(4679)) and (layer4_outputs(2386));
    layer5_outputs(3426) <= layer4_outputs(1443);
    layer5_outputs(3427) <= (layer4_outputs(4721)) or (layer4_outputs(3449));
    layer5_outputs(3428) <= not(layer4_outputs(2067)) or (layer4_outputs(5087));
    layer5_outputs(3429) <= layer4_outputs(2753);
    layer5_outputs(3430) <= (layer4_outputs(3111)) or (layer4_outputs(3311));
    layer5_outputs(3431) <= (layer4_outputs(2399)) xor (layer4_outputs(4596));
    layer5_outputs(3432) <= layer4_outputs(4735);
    layer5_outputs(3433) <= '0';
    layer5_outputs(3434) <= not(layer4_outputs(4636));
    layer5_outputs(3435) <= not(layer4_outputs(4647));
    layer5_outputs(3436) <= (layer4_outputs(296)) and not (layer4_outputs(4286));
    layer5_outputs(3437) <= layer4_outputs(21);
    layer5_outputs(3438) <= layer4_outputs(377);
    layer5_outputs(3439) <= layer4_outputs(3610);
    layer5_outputs(3440) <= not((layer4_outputs(3951)) and (layer4_outputs(1258)));
    layer5_outputs(3441) <= not((layer4_outputs(1225)) and (layer4_outputs(4414)));
    layer5_outputs(3442) <= not(layer4_outputs(3960));
    layer5_outputs(3443) <= (layer4_outputs(882)) and not (layer4_outputs(3962));
    layer5_outputs(3444) <= layer4_outputs(1384);
    layer5_outputs(3445) <= not(layer4_outputs(4190));
    layer5_outputs(3446) <= '0';
    layer5_outputs(3447) <= (layer4_outputs(2012)) and not (layer4_outputs(4598));
    layer5_outputs(3448) <= layer4_outputs(3052);
    layer5_outputs(3449) <= layer4_outputs(4773);
    layer5_outputs(3450) <= layer4_outputs(1436);
    layer5_outputs(3451) <= not((layer4_outputs(1326)) and (layer4_outputs(3556)));
    layer5_outputs(3452) <= layer4_outputs(2714);
    layer5_outputs(3453) <= not(layer4_outputs(4870));
    layer5_outputs(3454) <= not(layer4_outputs(1113));
    layer5_outputs(3455) <= (layer4_outputs(4943)) and (layer4_outputs(4800));
    layer5_outputs(3456) <= (layer4_outputs(3015)) and not (layer4_outputs(1715));
    layer5_outputs(3457) <= (layer4_outputs(3143)) and (layer4_outputs(1405));
    layer5_outputs(3458) <= (layer4_outputs(1162)) and not (layer4_outputs(194));
    layer5_outputs(3459) <= layer4_outputs(2896);
    layer5_outputs(3460) <= not((layer4_outputs(4564)) or (layer4_outputs(3669)));
    layer5_outputs(3461) <= not(layer4_outputs(1623));
    layer5_outputs(3462) <= '0';
    layer5_outputs(3463) <= layer4_outputs(1561);
    layer5_outputs(3464) <= not((layer4_outputs(3697)) and (layer4_outputs(2647)));
    layer5_outputs(3465) <= layer4_outputs(4837);
    layer5_outputs(3466) <= not(layer4_outputs(4730));
    layer5_outputs(3467) <= (layer4_outputs(4859)) xor (layer4_outputs(1172));
    layer5_outputs(3468) <= not(layer4_outputs(1296));
    layer5_outputs(3469) <= not(layer4_outputs(1713));
    layer5_outputs(3470) <= not(layer4_outputs(3650));
    layer5_outputs(3471) <= layer4_outputs(2265);
    layer5_outputs(3472) <= '0';
    layer5_outputs(3473) <= not((layer4_outputs(806)) and (layer4_outputs(1280)));
    layer5_outputs(3474) <= layer4_outputs(676);
    layer5_outputs(3475) <= layer4_outputs(3353);
    layer5_outputs(3476) <= not(layer4_outputs(663));
    layer5_outputs(3477) <= not((layer4_outputs(1007)) xor (layer4_outputs(147)));
    layer5_outputs(3478) <= not(layer4_outputs(1544)) or (layer4_outputs(3680));
    layer5_outputs(3479) <= not(layer4_outputs(3363));
    layer5_outputs(3480) <= layer4_outputs(1518);
    layer5_outputs(3481) <= (layer4_outputs(4296)) and (layer4_outputs(1747));
    layer5_outputs(3482) <= not((layer4_outputs(2539)) or (layer4_outputs(1509)));
    layer5_outputs(3483) <= layer4_outputs(1059);
    layer5_outputs(3484) <= (layer4_outputs(4073)) and (layer4_outputs(2409));
    layer5_outputs(3485) <= not(layer4_outputs(56));
    layer5_outputs(3486) <= layer4_outputs(4081);
    layer5_outputs(3487) <= not(layer4_outputs(850));
    layer5_outputs(3488) <= '1';
    layer5_outputs(3489) <= not(layer4_outputs(4383));
    layer5_outputs(3490) <= (layer4_outputs(3468)) xor (layer4_outputs(73));
    layer5_outputs(3491) <= (layer4_outputs(765)) and not (layer4_outputs(1803));
    layer5_outputs(3492) <= not(layer4_outputs(3511));
    layer5_outputs(3493) <= layer4_outputs(307);
    layer5_outputs(3494) <= layer4_outputs(4103);
    layer5_outputs(3495) <= not(layer4_outputs(292));
    layer5_outputs(3496) <= layer4_outputs(2971);
    layer5_outputs(3497) <= (layer4_outputs(433)) xor (layer4_outputs(1061));
    layer5_outputs(3498) <= not(layer4_outputs(3564));
    layer5_outputs(3499) <= layer4_outputs(931);
    layer5_outputs(3500) <= (layer4_outputs(771)) and (layer4_outputs(2505));
    layer5_outputs(3501) <= layer4_outputs(716);
    layer5_outputs(3502) <= not(layer4_outputs(2105));
    layer5_outputs(3503) <= (layer4_outputs(4984)) or (layer4_outputs(2241));
    layer5_outputs(3504) <= not(layer4_outputs(1051));
    layer5_outputs(3505) <= not(layer4_outputs(344));
    layer5_outputs(3506) <= not((layer4_outputs(4023)) or (layer4_outputs(1970)));
    layer5_outputs(3507) <= not(layer4_outputs(4424)) or (layer4_outputs(4344));
    layer5_outputs(3508) <= (layer4_outputs(3217)) and not (layer4_outputs(3753));
    layer5_outputs(3509) <= layer4_outputs(3946);
    layer5_outputs(3510) <= not(layer4_outputs(4964));
    layer5_outputs(3511) <= (layer4_outputs(4359)) or (layer4_outputs(2014));
    layer5_outputs(3512) <= not((layer4_outputs(3672)) or (layer4_outputs(1087)));
    layer5_outputs(3513) <= not(layer4_outputs(1230));
    layer5_outputs(3514) <= (layer4_outputs(2213)) and not (layer4_outputs(1703));
    layer5_outputs(3515) <= layer4_outputs(351);
    layer5_outputs(3516) <= layer4_outputs(1347);
    layer5_outputs(3517) <= layer4_outputs(4593);
    layer5_outputs(3518) <= (layer4_outputs(932)) and not (layer4_outputs(4705));
    layer5_outputs(3519) <= not(layer4_outputs(4371));
    layer5_outputs(3520) <= layer4_outputs(4342);
    layer5_outputs(3521) <= layer4_outputs(869);
    layer5_outputs(3522) <= not(layer4_outputs(2551));
    layer5_outputs(3523) <= '1';
    layer5_outputs(3524) <= not((layer4_outputs(2242)) and (layer4_outputs(1490)));
    layer5_outputs(3525) <= layer4_outputs(1701);
    layer5_outputs(3526) <= layer4_outputs(3822);
    layer5_outputs(3527) <= (layer4_outputs(2629)) xor (layer4_outputs(4486));
    layer5_outputs(3528) <= not(layer4_outputs(583));
    layer5_outputs(3529) <= not(layer4_outputs(2733));
    layer5_outputs(3530) <= not(layer4_outputs(5109));
    layer5_outputs(3531) <= not(layer4_outputs(2439)) or (layer4_outputs(4274));
    layer5_outputs(3532) <= (layer4_outputs(2269)) and not (layer4_outputs(4836));
    layer5_outputs(3533) <= layer4_outputs(4719);
    layer5_outputs(3534) <= not(layer4_outputs(2322)) or (layer4_outputs(3864));
    layer5_outputs(3535) <= layer4_outputs(3618);
    layer5_outputs(3536) <= not(layer4_outputs(1879)) or (layer4_outputs(363));
    layer5_outputs(3537) <= (layer4_outputs(3489)) or (layer4_outputs(614));
    layer5_outputs(3538) <= not(layer4_outputs(2198));
    layer5_outputs(3539) <= not((layer4_outputs(894)) and (layer4_outputs(1641)));
    layer5_outputs(3540) <= (layer4_outputs(1793)) and not (layer4_outputs(1674));
    layer5_outputs(3541) <= not(layer4_outputs(2962));
    layer5_outputs(3542) <= layer4_outputs(1468);
    layer5_outputs(3543) <= layer4_outputs(4215);
    layer5_outputs(3544) <= not(layer4_outputs(158));
    layer5_outputs(3545) <= not(layer4_outputs(3611));
    layer5_outputs(3546) <= not(layer4_outputs(4714));
    layer5_outputs(3547) <= not(layer4_outputs(4790)) or (layer4_outputs(233));
    layer5_outputs(3548) <= not(layer4_outputs(93));
    layer5_outputs(3549) <= not(layer4_outputs(4930)) or (layer4_outputs(1378));
    layer5_outputs(3550) <= not(layer4_outputs(3990)) or (layer4_outputs(1118));
    layer5_outputs(3551) <= layer4_outputs(2831);
    layer5_outputs(3552) <= (layer4_outputs(1177)) and (layer4_outputs(2597));
    layer5_outputs(3553) <= (layer4_outputs(4655)) and (layer4_outputs(1860));
    layer5_outputs(3554) <= layer4_outputs(2177);
    layer5_outputs(3555) <= (layer4_outputs(3115)) and not (layer4_outputs(3493));
    layer5_outputs(3556) <= layer4_outputs(3740);
    layer5_outputs(3557) <= layer4_outputs(635);
    layer5_outputs(3558) <= not((layer4_outputs(3064)) or (layer4_outputs(3416)));
    layer5_outputs(3559) <= not(layer4_outputs(1830));
    layer5_outputs(3560) <= (layer4_outputs(1606)) or (layer4_outputs(4127));
    layer5_outputs(3561) <= layer4_outputs(3309);
    layer5_outputs(3562) <= not(layer4_outputs(156));
    layer5_outputs(3563) <= not((layer4_outputs(703)) xor (layer4_outputs(3083)));
    layer5_outputs(3564) <= not((layer4_outputs(4551)) xor (layer4_outputs(1649)));
    layer5_outputs(3565) <= not((layer4_outputs(314)) and (layer4_outputs(817)));
    layer5_outputs(3566) <= not(layer4_outputs(3752));
    layer5_outputs(3567) <= not(layer4_outputs(2116)) or (layer4_outputs(2996));
    layer5_outputs(3568) <= not(layer4_outputs(642));
    layer5_outputs(3569) <= layer4_outputs(1654);
    layer5_outputs(3570) <= '1';
    layer5_outputs(3571) <= not((layer4_outputs(1184)) and (layer4_outputs(3106)));
    layer5_outputs(3572) <= not(layer4_outputs(3540));
    layer5_outputs(3573) <= (layer4_outputs(4707)) and (layer4_outputs(1156));
    layer5_outputs(3574) <= layer4_outputs(2352);
    layer5_outputs(3575) <= layer4_outputs(4103);
    layer5_outputs(3576) <= (layer4_outputs(2662)) or (layer4_outputs(2738));
    layer5_outputs(3577) <= (layer4_outputs(4760)) xor (layer4_outputs(4001));
    layer5_outputs(3578) <= (layer4_outputs(3794)) and not (layer4_outputs(1865));
    layer5_outputs(3579) <= not(layer4_outputs(923));
    layer5_outputs(3580) <= not(layer4_outputs(3515)) or (layer4_outputs(5043));
    layer5_outputs(3581) <= not(layer4_outputs(3368));
    layer5_outputs(3582) <= not(layer4_outputs(4298)) or (layer4_outputs(3056));
    layer5_outputs(3583) <= '1';
    layer5_outputs(3584) <= layer4_outputs(1927);
    layer5_outputs(3585) <= not(layer4_outputs(1457)) or (layer4_outputs(3046));
    layer5_outputs(3586) <= (layer4_outputs(4160)) and (layer4_outputs(975));
    layer5_outputs(3587) <= layer4_outputs(3909);
    layer5_outputs(3588) <= layer4_outputs(4902);
    layer5_outputs(3589) <= (layer4_outputs(3579)) xor (layer4_outputs(2035));
    layer5_outputs(3590) <= layer4_outputs(3878);
    layer5_outputs(3591) <= not(layer4_outputs(837)) or (layer4_outputs(3197));
    layer5_outputs(3592) <= (layer4_outputs(1809)) and not (layer4_outputs(2972));
    layer5_outputs(3593) <= not(layer4_outputs(4669));
    layer5_outputs(3594) <= layer4_outputs(2596);
    layer5_outputs(3595) <= layer4_outputs(2744);
    layer5_outputs(3596) <= not(layer4_outputs(2126)) or (layer4_outputs(3078));
    layer5_outputs(3597) <= not(layer4_outputs(3160));
    layer5_outputs(3598) <= layer4_outputs(404);
    layer5_outputs(3599) <= layer4_outputs(3035);
    layer5_outputs(3600) <= not(layer4_outputs(2998));
    layer5_outputs(3601) <= layer4_outputs(4782);
    layer5_outputs(3602) <= (layer4_outputs(541)) and (layer4_outputs(4513));
    layer5_outputs(3603) <= not(layer4_outputs(3817));
    layer5_outputs(3604) <= not((layer4_outputs(3903)) and (layer4_outputs(942)));
    layer5_outputs(3605) <= layer4_outputs(2060);
    layer5_outputs(3606) <= not(layer4_outputs(5026));
    layer5_outputs(3607) <= (layer4_outputs(4627)) xor (layer4_outputs(293));
    layer5_outputs(3608) <= not(layer4_outputs(3530));
    layer5_outputs(3609) <= not((layer4_outputs(770)) xor (layer4_outputs(4851)));
    layer5_outputs(3610) <= (layer4_outputs(2035)) xor (layer4_outputs(1798));
    layer5_outputs(3611) <= '1';
    layer5_outputs(3612) <= (layer4_outputs(1877)) and not (layer4_outputs(4605));
    layer5_outputs(3613) <= (layer4_outputs(2404)) and not (layer4_outputs(4456));
    layer5_outputs(3614) <= not(layer4_outputs(1483));
    layer5_outputs(3615) <= not(layer4_outputs(2394));
    layer5_outputs(3616) <= (layer4_outputs(4481)) and not (layer4_outputs(2615));
    layer5_outputs(3617) <= (layer4_outputs(2913)) and not (layer4_outputs(675));
    layer5_outputs(3618) <= not((layer4_outputs(3048)) xor (layer4_outputs(2833)));
    layer5_outputs(3619) <= not((layer4_outputs(3872)) or (layer4_outputs(713)));
    layer5_outputs(3620) <= not(layer4_outputs(4648));
    layer5_outputs(3621) <= not((layer4_outputs(493)) and (layer4_outputs(4346)));
    layer5_outputs(3622) <= not(layer4_outputs(5));
    layer5_outputs(3623) <= layer4_outputs(2679);
    layer5_outputs(3624) <= not((layer4_outputs(3279)) and (layer4_outputs(857)));
    layer5_outputs(3625) <= layer4_outputs(511);
    layer5_outputs(3626) <= not(layer4_outputs(2155));
    layer5_outputs(3627) <= layer4_outputs(3145);
    layer5_outputs(3628) <= (layer4_outputs(2530)) and not (layer4_outputs(2746));
    layer5_outputs(3629) <= layer4_outputs(5077);
    layer5_outputs(3630) <= not(layer4_outputs(334));
    layer5_outputs(3631) <= (layer4_outputs(1244)) and not (layer4_outputs(529));
    layer5_outputs(3632) <= not(layer4_outputs(3185));
    layer5_outputs(3633) <= not(layer4_outputs(3743));
    layer5_outputs(3634) <= (layer4_outputs(356)) and not (layer4_outputs(3810));
    layer5_outputs(3635) <= layer4_outputs(3859);
    layer5_outputs(3636) <= layer4_outputs(682);
    layer5_outputs(3637) <= '0';
    layer5_outputs(3638) <= not((layer4_outputs(2451)) or (layer4_outputs(4523)));
    layer5_outputs(3639) <= layer4_outputs(1178);
    layer5_outputs(3640) <= layer4_outputs(287);
    layer5_outputs(3641) <= not(layer4_outputs(3820)) or (layer4_outputs(5083));
    layer5_outputs(3642) <= not((layer4_outputs(1471)) xor (layer4_outputs(2440)));
    layer5_outputs(3643) <= not(layer4_outputs(1575));
    layer5_outputs(3644) <= not(layer4_outputs(4980)) or (layer4_outputs(1268));
    layer5_outputs(3645) <= (layer4_outputs(1380)) xor (layer4_outputs(2269));
    layer5_outputs(3646) <= layer4_outputs(830);
    layer5_outputs(3647) <= layer4_outputs(2182);
    layer5_outputs(3648) <= not(layer4_outputs(1063));
    layer5_outputs(3649) <= not(layer4_outputs(1507));
    layer5_outputs(3650) <= not(layer4_outputs(368));
    layer5_outputs(3651) <= not((layer4_outputs(4095)) or (layer4_outputs(724)));
    layer5_outputs(3652) <= layer4_outputs(2638);
    layer5_outputs(3653) <= layer4_outputs(1639);
    layer5_outputs(3654) <= layer4_outputs(2876);
    layer5_outputs(3655) <= '0';
    layer5_outputs(3656) <= not(layer4_outputs(4749));
    layer5_outputs(3657) <= not(layer4_outputs(4011)) or (layer4_outputs(2667));
    layer5_outputs(3658) <= (layer4_outputs(4457)) and not (layer4_outputs(2767));
    layer5_outputs(3659) <= (layer4_outputs(2564)) and not (layer4_outputs(3678));
    layer5_outputs(3660) <= layer4_outputs(2753);
    layer5_outputs(3661) <= not(layer4_outputs(2714));
    layer5_outputs(3662) <= not((layer4_outputs(2518)) and (layer4_outputs(4238)));
    layer5_outputs(3663) <= not(layer4_outputs(4302)) or (layer4_outputs(4633));
    layer5_outputs(3664) <= (layer4_outputs(3029)) xor (layer4_outputs(432));
    layer5_outputs(3665) <= not(layer4_outputs(3341));
    layer5_outputs(3666) <= not(layer4_outputs(1834));
    layer5_outputs(3667) <= not((layer4_outputs(3640)) and (layer4_outputs(4498)));
    layer5_outputs(3668) <= not(layer4_outputs(127));
    layer5_outputs(3669) <= layer4_outputs(4236);
    layer5_outputs(3670) <= not((layer4_outputs(217)) or (layer4_outputs(1046)));
    layer5_outputs(3671) <= (layer4_outputs(1510)) xor (layer4_outputs(2048));
    layer5_outputs(3672) <= not((layer4_outputs(1421)) and (layer4_outputs(4137)));
    layer5_outputs(3673) <= not(layer4_outputs(4590));
    layer5_outputs(3674) <= not(layer4_outputs(4547));
    layer5_outputs(3675) <= not(layer4_outputs(2398)) or (layer4_outputs(4974));
    layer5_outputs(3676) <= layer4_outputs(5029);
    layer5_outputs(3677) <= (layer4_outputs(23)) and not (layer4_outputs(3230));
    layer5_outputs(3678) <= (layer4_outputs(1781)) or (layer4_outputs(2859));
    layer5_outputs(3679) <= not(layer4_outputs(2831));
    layer5_outputs(3680) <= not(layer4_outputs(2102));
    layer5_outputs(3681) <= '0';
    layer5_outputs(3682) <= not((layer4_outputs(3)) xor (layer4_outputs(1364)));
    layer5_outputs(3683) <= layer4_outputs(3520);
    layer5_outputs(3684) <= not(layer4_outputs(3807));
    layer5_outputs(3685) <= not((layer4_outputs(1361)) or (layer4_outputs(3908)));
    layer5_outputs(3686) <= not(layer4_outputs(3573));
    layer5_outputs(3687) <= not(layer4_outputs(1274));
    layer5_outputs(3688) <= not(layer4_outputs(270));
    layer5_outputs(3689) <= layer4_outputs(5012);
    layer5_outputs(3690) <= (layer4_outputs(4418)) and not (layer4_outputs(4168));
    layer5_outputs(3691) <= not(layer4_outputs(259));
    layer5_outputs(3692) <= not(layer4_outputs(4815));
    layer5_outputs(3693) <= not(layer4_outputs(1482));
    layer5_outputs(3694) <= layer4_outputs(4693);
    layer5_outputs(3695) <= '1';
    layer5_outputs(3696) <= not(layer4_outputs(3175));
    layer5_outputs(3697) <= (layer4_outputs(3342)) and (layer4_outputs(1123));
    layer5_outputs(3698) <= '0';
    layer5_outputs(3699) <= not(layer4_outputs(1093));
    layer5_outputs(3700) <= not(layer4_outputs(4854));
    layer5_outputs(3701) <= layer4_outputs(1365);
    layer5_outputs(3702) <= (layer4_outputs(624)) and (layer4_outputs(1211));
    layer5_outputs(3703) <= not(layer4_outputs(4384)) or (layer4_outputs(4129));
    layer5_outputs(3704) <= not(layer4_outputs(820));
    layer5_outputs(3705) <= (layer4_outputs(723)) and not (layer4_outputs(2379));
    layer5_outputs(3706) <= (layer4_outputs(4958)) and not (layer4_outputs(2332));
    layer5_outputs(3707) <= not(layer4_outputs(112));
    layer5_outputs(3708) <= not(layer4_outputs(1791)) or (layer4_outputs(3705));
    layer5_outputs(3709) <= layer4_outputs(128);
    layer5_outputs(3710) <= not(layer4_outputs(1485));
    layer5_outputs(3711) <= not(layer4_outputs(1795));
    layer5_outputs(3712) <= (layer4_outputs(544)) or (layer4_outputs(4130));
    layer5_outputs(3713) <= not(layer4_outputs(1183)) or (layer4_outputs(3937));
    layer5_outputs(3714) <= (layer4_outputs(768)) and not (layer4_outputs(2554));
    layer5_outputs(3715) <= '1';
    layer5_outputs(3716) <= (layer4_outputs(3682)) and not (layer4_outputs(1875));
    layer5_outputs(3717) <= (layer4_outputs(2781)) and not (layer4_outputs(2524));
    layer5_outputs(3718) <= not((layer4_outputs(454)) xor (layer4_outputs(2866)));
    layer5_outputs(3719) <= layer4_outputs(4573);
    layer5_outputs(3720) <= not(layer4_outputs(4976)) or (layer4_outputs(1355));
    layer5_outputs(3721) <= '1';
    layer5_outputs(3722) <= not((layer4_outputs(1934)) and (layer4_outputs(4380)));
    layer5_outputs(3723) <= layer4_outputs(1370);
    layer5_outputs(3724) <= layer4_outputs(3852);
    layer5_outputs(3725) <= (layer4_outputs(420)) and not (layer4_outputs(4676));
    layer5_outputs(3726) <= (layer4_outputs(5008)) xor (layer4_outputs(3258));
    layer5_outputs(3727) <= '0';
    layer5_outputs(3728) <= not(layer4_outputs(3249)) or (layer4_outputs(5104));
    layer5_outputs(3729) <= layer4_outputs(4236);
    layer5_outputs(3730) <= not(layer4_outputs(2142));
    layer5_outputs(3731) <= layer4_outputs(461);
    layer5_outputs(3732) <= not(layer4_outputs(1586));
    layer5_outputs(3733) <= not(layer4_outputs(1713));
    layer5_outputs(3734) <= not(layer4_outputs(286)) or (layer4_outputs(3966));
    layer5_outputs(3735) <= not(layer4_outputs(4212));
    layer5_outputs(3736) <= layer4_outputs(4035);
    layer5_outputs(3737) <= layer4_outputs(1743);
    layer5_outputs(3738) <= not(layer4_outputs(187));
    layer5_outputs(3739) <= layer4_outputs(107);
    layer5_outputs(3740) <= not((layer4_outputs(559)) and (layer4_outputs(2240)));
    layer5_outputs(3741) <= layer4_outputs(4781);
    layer5_outputs(3742) <= '1';
    layer5_outputs(3743) <= not(layer4_outputs(808));
    layer5_outputs(3744) <= not(layer4_outputs(2501));
    layer5_outputs(3745) <= not(layer4_outputs(1245));
    layer5_outputs(3746) <= (layer4_outputs(5023)) and not (layer4_outputs(952));
    layer5_outputs(3747) <= not(layer4_outputs(1882)) or (layer4_outputs(4816));
    layer5_outputs(3748) <= not(layer4_outputs(4495));
    layer5_outputs(3749) <= not(layer4_outputs(4383));
    layer5_outputs(3750) <= (layer4_outputs(1167)) and not (layer4_outputs(2917));
    layer5_outputs(3751) <= '1';
    layer5_outputs(3752) <= (layer4_outputs(4934)) or (layer4_outputs(1003));
    layer5_outputs(3753) <= layer4_outputs(4216);
    layer5_outputs(3754) <= layer4_outputs(3684);
    layer5_outputs(3755) <= (layer4_outputs(465)) and not (layer4_outputs(4743));
    layer5_outputs(3756) <= not(layer4_outputs(2609));
    layer5_outputs(3757) <= not(layer4_outputs(1866)) or (layer4_outputs(4040));
    layer5_outputs(3758) <= (layer4_outputs(4136)) xor (layer4_outputs(326));
    layer5_outputs(3759) <= (layer4_outputs(3557)) and not (layer4_outputs(4159));
    layer5_outputs(3760) <= layer4_outputs(4469);
    layer5_outputs(3761) <= not((layer4_outputs(2649)) or (layer4_outputs(2886)));
    layer5_outputs(3762) <= (layer4_outputs(4536)) or (layer4_outputs(4711));
    layer5_outputs(3763) <= not(layer4_outputs(3711));
    layer5_outputs(3764) <= (layer4_outputs(2380)) or (layer4_outputs(1661));
    layer5_outputs(3765) <= '1';
    layer5_outputs(3766) <= (layer4_outputs(1863)) or (layer4_outputs(2539));
    layer5_outputs(3767) <= (layer4_outputs(3898)) xor (layer4_outputs(1170));
    layer5_outputs(3768) <= layer4_outputs(4720);
    layer5_outputs(3769) <= not(layer4_outputs(708)) or (layer4_outputs(4736));
    layer5_outputs(3770) <= not((layer4_outputs(3387)) and (layer4_outputs(794)));
    layer5_outputs(3771) <= not(layer4_outputs(442)) or (layer4_outputs(3918));
    layer5_outputs(3772) <= not(layer4_outputs(177));
    layer5_outputs(3773) <= layer4_outputs(643);
    layer5_outputs(3774) <= layer4_outputs(1869);
    layer5_outputs(3775) <= (layer4_outputs(4368)) and not (layer4_outputs(1315));
    layer5_outputs(3776) <= not((layer4_outputs(929)) or (layer4_outputs(244)));
    layer5_outputs(3777) <= (layer4_outputs(2428)) xor (layer4_outputs(4561));
    layer5_outputs(3778) <= not(layer4_outputs(4584));
    layer5_outputs(3779) <= not(layer4_outputs(1838)) or (layer4_outputs(791));
    layer5_outputs(3780) <= not(layer4_outputs(919)) or (layer4_outputs(1081));
    layer5_outputs(3781) <= (layer4_outputs(817)) and not (layer4_outputs(5077));
    layer5_outputs(3782) <= not(layer4_outputs(3587));
    layer5_outputs(3783) <= (layer4_outputs(3877)) and not (layer4_outputs(507));
    layer5_outputs(3784) <= layer4_outputs(4080);
    layer5_outputs(3785) <= not((layer4_outputs(4742)) or (layer4_outputs(2250)));
    layer5_outputs(3786) <= not(layer4_outputs(3970));
    layer5_outputs(3787) <= layer4_outputs(4524);
    layer5_outputs(3788) <= layer4_outputs(369);
    layer5_outputs(3789) <= not((layer4_outputs(3345)) and (layer4_outputs(4058)));
    layer5_outputs(3790) <= layer4_outputs(807);
    layer5_outputs(3791) <= (layer4_outputs(4605)) and not (layer4_outputs(696));
    layer5_outputs(3792) <= (layer4_outputs(4449)) or (layer4_outputs(1206));
    layer5_outputs(3793) <= (layer4_outputs(1670)) and not (layer4_outputs(2889));
    layer5_outputs(3794) <= not((layer4_outputs(4903)) or (layer4_outputs(641)));
    layer5_outputs(3795) <= not((layer4_outputs(970)) and (layer4_outputs(1728)));
    layer5_outputs(3796) <= layer4_outputs(1050);
    layer5_outputs(3797) <= (layer4_outputs(1387)) and not (layer4_outputs(1827));
    layer5_outputs(3798) <= not(layer4_outputs(41));
    layer5_outputs(3799) <= layer4_outputs(147);
    layer5_outputs(3800) <= not(layer4_outputs(1481));
    layer5_outputs(3801) <= not(layer4_outputs(77)) or (layer4_outputs(4200));
    layer5_outputs(3802) <= not(layer4_outputs(2170));
    layer5_outputs(3803) <= not(layer4_outputs(4849));
    layer5_outputs(3804) <= (layer4_outputs(4024)) and not (layer4_outputs(2867));
    layer5_outputs(3805) <= layer4_outputs(627);
    layer5_outputs(3806) <= layer4_outputs(1980);
    layer5_outputs(3807) <= '0';
    layer5_outputs(3808) <= layer4_outputs(3669);
    layer5_outputs(3809) <= not(layer4_outputs(611)) or (layer4_outputs(1250));
    layer5_outputs(3810) <= (layer4_outputs(4432)) or (layer4_outputs(2191));
    layer5_outputs(3811) <= (layer4_outputs(4554)) and not (layer4_outputs(2396));
    layer5_outputs(3812) <= layer4_outputs(240);
    layer5_outputs(3813) <= not(layer4_outputs(1097));
    layer5_outputs(3814) <= '0';
    layer5_outputs(3815) <= layer4_outputs(4591);
    layer5_outputs(3816) <= not((layer4_outputs(4338)) and (layer4_outputs(3196)));
    layer5_outputs(3817) <= not(layer4_outputs(2132)) or (layer4_outputs(3562));
    layer5_outputs(3818) <= not(layer4_outputs(716));
    layer5_outputs(3819) <= '1';
    layer5_outputs(3820) <= not(layer4_outputs(1739));
    layer5_outputs(3821) <= (layer4_outputs(1357)) and not (layer4_outputs(258));
    layer5_outputs(3822) <= (layer4_outputs(3166)) and not (layer4_outputs(2369));
    layer5_outputs(3823) <= layer4_outputs(1058);
    layer5_outputs(3824) <= not(layer4_outputs(3114));
    layer5_outputs(3825) <= layer4_outputs(183);
    layer5_outputs(3826) <= not(layer4_outputs(2883));
    layer5_outputs(3827) <= not(layer4_outputs(1955)) or (layer4_outputs(1518));
    layer5_outputs(3828) <= not((layer4_outputs(4746)) and (layer4_outputs(4085)));
    layer5_outputs(3829) <= '0';
    layer5_outputs(3830) <= not(layer4_outputs(65)) or (layer4_outputs(4042));
    layer5_outputs(3831) <= not(layer4_outputs(4209));
    layer5_outputs(3832) <= layer4_outputs(2949);
    layer5_outputs(3833) <= not(layer4_outputs(5118)) or (layer4_outputs(2307));
    layer5_outputs(3834) <= layer4_outputs(1731);
    layer5_outputs(3835) <= not(layer4_outputs(1892));
    layer5_outputs(3836) <= layer4_outputs(2007);
    layer5_outputs(3837) <= not((layer4_outputs(1470)) and (layer4_outputs(1686)));
    layer5_outputs(3838) <= layer4_outputs(2037);
    layer5_outputs(3839) <= not((layer4_outputs(1716)) xor (layer4_outputs(1242)));
    layer5_outputs(3840) <= layer4_outputs(3087);
    layer5_outputs(3841) <= '1';
    layer5_outputs(3842) <= not(layer4_outputs(4412));
    layer5_outputs(3843) <= not(layer4_outputs(134));
    layer5_outputs(3844) <= not(layer4_outputs(4587));
    layer5_outputs(3845) <= not(layer4_outputs(1114));
    layer5_outputs(3846) <= '1';
    layer5_outputs(3847) <= not(layer4_outputs(1049)) or (layer4_outputs(2361));
    layer5_outputs(3848) <= not(layer4_outputs(4966));
    layer5_outputs(3849) <= (layer4_outputs(4643)) xor (layer4_outputs(2243));
    layer5_outputs(3850) <= (layer4_outputs(1580)) or (layer4_outputs(3886));
    layer5_outputs(3851) <= layer4_outputs(3741);
    layer5_outputs(3852) <= (layer4_outputs(3327)) xor (layer4_outputs(2804));
    layer5_outputs(3853) <= layer4_outputs(4261);
    layer5_outputs(3854) <= not(layer4_outputs(4677));
    layer5_outputs(3855) <= (layer4_outputs(1214)) xor (layer4_outputs(2686));
    layer5_outputs(3856) <= '0';
    layer5_outputs(3857) <= not(layer4_outputs(3747));
    layer5_outputs(3858) <= (layer4_outputs(1324)) and not (layer4_outputs(3779));
    layer5_outputs(3859) <= not((layer4_outputs(233)) and (layer4_outputs(3200)));
    layer5_outputs(3860) <= layer4_outputs(4263);
    layer5_outputs(3861) <= (layer4_outputs(1790)) and not (layer4_outputs(4398));
    layer5_outputs(3862) <= (layer4_outputs(3287)) or (layer4_outputs(4474));
    layer5_outputs(3863) <= layer4_outputs(4060);
    layer5_outputs(3864) <= not(layer4_outputs(5021));
    layer5_outputs(3865) <= (layer4_outputs(2715)) and (layer4_outputs(221));
    layer5_outputs(3866) <= (layer4_outputs(2247)) and (layer4_outputs(4978));
    layer5_outputs(3867) <= not(layer4_outputs(1769));
    layer5_outputs(3868) <= not((layer4_outputs(4743)) xor (layer4_outputs(1157)));
    layer5_outputs(3869) <= '0';
    layer5_outputs(3870) <= not(layer4_outputs(4387));
    layer5_outputs(3871) <= not(layer4_outputs(3580));
    layer5_outputs(3872) <= '1';
    layer5_outputs(3873) <= layer4_outputs(4163);
    layer5_outputs(3874) <= not(layer4_outputs(859));
    layer5_outputs(3875) <= not(layer4_outputs(199)) or (layer4_outputs(1090));
    layer5_outputs(3876) <= not(layer4_outputs(3964));
    layer5_outputs(3877) <= not(layer4_outputs(1204)) or (layer4_outputs(3192));
    layer5_outputs(3878) <= (layer4_outputs(1796)) and (layer4_outputs(1243));
    layer5_outputs(3879) <= layer4_outputs(2089);
    layer5_outputs(3880) <= not(layer4_outputs(2570)) or (layer4_outputs(4173));
    layer5_outputs(3881) <= not(layer4_outputs(3484));
    layer5_outputs(3882) <= not((layer4_outputs(2034)) and (layer4_outputs(1110)));
    layer5_outputs(3883) <= not(layer4_outputs(618));
    layer5_outputs(3884) <= not(layer4_outputs(2458));
    layer5_outputs(3885) <= (layer4_outputs(1187)) and not (layer4_outputs(1881));
    layer5_outputs(3886) <= not(layer4_outputs(3897));
    layer5_outputs(3887) <= layer4_outputs(3365);
    layer5_outputs(3888) <= (layer4_outputs(1397)) and not (layer4_outputs(3379));
    layer5_outputs(3889) <= (layer4_outputs(4102)) or (layer4_outputs(508));
    layer5_outputs(3890) <= (layer4_outputs(4628)) and not (layer4_outputs(4284));
    layer5_outputs(3891) <= not(layer4_outputs(3492)) or (layer4_outputs(3447));
    layer5_outputs(3892) <= not((layer4_outputs(4888)) xor (layer4_outputs(585)));
    layer5_outputs(3893) <= not(layer4_outputs(1388));
    layer5_outputs(3894) <= not(layer4_outputs(3763));
    layer5_outputs(3895) <= not(layer4_outputs(4291)) or (layer4_outputs(3698));
    layer5_outputs(3896) <= not((layer4_outputs(3067)) and (layer4_outputs(4273)));
    layer5_outputs(3897) <= not((layer4_outputs(1759)) or (layer4_outputs(3318)));
    layer5_outputs(3898) <= (layer4_outputs(2838)) and (layer4_outputs(3044));
    layer5_outputs(3899) <= not(layer4_outputs(3995));
    layer5_outputs(3900) <= not((layer4_outputs(411)) or (layer4_outputs(1091)));
    layer5_outputs(3901) <= not(layer4_outputs(4318));
    layer5_outputs(3902) <= not((layer4_outputs(3661)) or (layer4_outputs(3079)));
    layer5_outputs(3903) <= not(layer4_outputs(1497));
    layer5_outputs(3904) <= not((layer4_outputs(3766)) or (layer4_outputs(155)));
    layer5_outputs(3905) <= layer4_outputs(5090);
    layer5_outputs(3906) <= layer4_outputs(979);
    layer5_outputs(3907) <= not(layer4_outputs(3197)) or (layer4_outputs(44));
    layer5_outputs(3908) <= not((layer4_outputs(2298)) or (layer4_outputs(534)));
    layer5_outputs(3909) <= (layer4_outputs(2694)) or (layer4_outputs(5006));
    layer5_outputs(3910) <= layer4_outputs(2273);
    layer5_outputs(3911) <= not(layer4_outputs(2451));
    layer5_outputs(3912) <= layer4_outputs(4131);
    layer5_outputs(3913) <= not(layer4_outputs(3328)) or (layer4_outputs(4276));
    layer5_outputs(3914) <= not(layer4_outputs(3159));
    layer5_outputs(3915) <= layer4_outputs(2911);
    layer5_outputs(3916) <= not((layer4_outputs(3539)) and (layer4_outputs(2497)));
    layer5_outputs(3917) <= not(layer4_outputs(4649)) or (layer4_outputs(2842));
    layer5_outputs(3918) <= not(layer4_outputs(2405));
    layer5_outputs(3919) <= not(layer4_outputs(2796));
    layer5_outputs(3920) <= not(layer4_outputs(4678)) or (layer4_outputs(2219));
    layer5_outputs(3921) <= (layer4_outputs(2985)) and not (layer4_outputs(1963));
    layer5_outputs(3922) <= not(layer4_outputs(4066));
    layer5_outputs(3923) <= layer4_outputs(2644);
    layer5_outputs(3924) <= layer4_outputs(3132);
    layer5_outputs(3925) <= (layer4_outputs(4544)) xor (layer4_outputs(3180));
    layer5_outputs(3926) <= (layer4_outputs(1691)) and not (layer4_outputs(3401));
    layer5_outputs(3927) <= layer4_outputs(3175);
    layer5_outputs(3928) <= not(layer4_outputs(3612));
    layer5_outputs(3929) <= not((layer4_outputs(1534)) xor (layer4_outputs(5045)));
    layer5_outputs(3930) <= (layer4_outputs(3346)) and not (layer4_outputs(2783));
    layer5_outputs(3931) <= not(layer4_outputs(4202));
    layer5_outputs(3932) <= layer4_outputs(4287);
    layer5_outputs(3933) <= not(layer4_outputs(2183)) or (layer4_outputs(2353));
    layer5_outputs(3934) <= not((layer4_outputs(960)) xor (layer4_outputs(2297)));
    layer5_outputs(3935) <= not(layer4_outputs(2789));
    layer5_outputs(3936) <= not((layer4_outputs(4027)) and (layer4_outputs(2253)));
    layer5_outputs(3937) <= not(layer4_outputs(1191)) or (layer4_outputs(4475));
    layer5_outputs(3938) <= (layer4_outputs(484)) and not (layer4_outputs(4629));
    layer5_outputs(3939) <= (layer4_outputs(3071)) and not (layer4_outputs(2670));
    layer5_outputs(3940) <= layer4_outputs(4240);
    layer5_outputs(3941) <= not((layer4_outputs(1297)) or (layer4_outputs(3922)));
    layer5_outputs(3942) <= not(layer4_outputs(4341));
    layer5_outputs(3943) <= (layer4_outputs(1978)) or (layer4_outputs(1711));
    layer5_outputs(3944) <= not((layer4_outputs(4851)) xor (layer4_outputs(2284)));
    layer5_outputs(3945) <= layer4_outputs(662);
    layer5_outputs(3946) <= (layer4_outputs(2091)) or (layer4_outputs(659));
    layer5_outputs(3947) <= (layer4_outputs(3767)) xor (layer4_outputs(1358));
    layer5_outputs(3948) <= layer4_outputs(1861);
    layer5_outputs(3949) <= not(layer4_outputs(1447)) or (layer4_outputs(1210));
    layer5_outputs(3950) <= (layer4_outputs(1707)) and not (layer4_outputs(1721));
    layer5_outputs(3951) <= '1';
    layer5_outputs(3952) <= layer4_outputs(1556);
    layer5_outputs(3953) <= not(layer4_outputs(4206));
    layer5_outputs(3954) <= layer4_outputs(224);
    layer5_outputs(3955) <= (layer4_outputs(3817)) xor (layer4_outputs(964));
    layer5_outputs(3956) <= not(layer4_outputs(2754));
    layer5_outputs(3957) <= not(layer4_outputs(247));
    layer5_outputs(3958) <= not(layer4_outputs(2553));
    layer5_outputs(3959) <= not(layer4_outputs(1858));
    layer5_outputs(3960) <= (layer4_outputs(2868)) or (layer4_outputs(2300));
    layer5_outputs(3961) <= layer4_outputs(3973);
    layer5_outputs(3962) <= not((layer4_outputs(1198)) or (layer4_outputs(1016)));
    layer5_outputs(3963) <= layer4_outputs(1501);
    layer5_outputs(3964) <= (layer4_outputs(2891)) and (layer4_outputs(4134));
    layer5_outputs(3965) <= (layer4_outputs(2963)) and not (layer4_outputs(2044));
    layer5_outputs(3966) <= not(layer4_outputs(3641)) or (layer4_outputs(706));
    layer5_outputs(3967) <= not((layer4_outputs(1269)) xor (layer4_outputs(4908)));
    layer5_outputs(3968) <= (layer4_outputs(3078)) or (layer4_outputs(2885));
    layer5_outputs(3969) <= not(layer4_outputs(4465));
    layer5_outputs(3970) <= layer4_outputs(4658);
    layer5_outputs(3971) <= not(layer4_outputs(3876)) or (layer4_outputs(4683));
    layer5_outputs(3972) <= (layer4_outputs(69)) or (layer4_outputs(5047));
    layer5_outputs(3973) <= layer4_outputs(4320);
    layer5_outputs(3974) <= layer4_outputs(4206);
    layer5_outputs(3975) <= not(layer4_outputs(4264));
    layer5_outputs(3976) <= (layer4_outputs(859)) or (layer4_outputs(4435));
    layer5_outputs(3977) <= '1';
    layer5_outputs(3978) <= not((layer4_outputs(1182)) or (layer4_outputs(3882)));
    layer5_outputs(3979) <= (layer4_outputs(3773)) and (layer4_outputs(110));
    layer5_outputs(3980) <= not(layer4_outputs(985));
    layer5_outputs(3981) <= not((layer4_outputs(2884)) or (layer4_outputs(2701)));
    layer5_outputs(3982) <= not(layer4_outputs(1458));
    layer5_outputs(3983) <= not(layer4_outputs(136)) or (layer4_outputs(1328));
    layer5_outputs(3984) <= layer4_outputs(2345);
    layer5_outputs(3985) <= (layer4_outputs(1504)) and not (layer4_outputs(3108));
    layer5_outputs(3986) <= not((layer4_outputs(1918)) and (layer4_outputs(1517)));
    layer5_outputs(3987) <= not(layer4_outputs(4379));
    layer5_outputs(3988) <= (layer4_outputs(3403)) or (layer4_outputs(1358));
    layer5_outputs(3989) <= (layer4_outputs(922)) and (layer4_outputs(1735));
    layer5_outputs(3990) <= (layer4_outputs(4433)) or (layer4_outputs(2655));
    layer5_outputs(3991) <= not(layer4_outputs(649));
    layer5_outputs(3992) <= not(layer4_outputs(4823)) or (layer4_outputs(789));
    layer5_outputs(3993) <= layer4_outputs(4165);
    layer5_outputs(3994) <= layer4_outputs(1770);
    layer5_outputs(3995) <= '1';
    layer5_outputs(3996) <= not(layer4_outputs(82));
    layer5_outputs(3997) <= layer4_outputs(3862);
    layer5_outputs(3998) <= layer4_outputs(4791);
    layer5_outputs(3999) <= not(layer4_outputs(1588));
    layer5_outputs(4000) <= not(layer4_outputs(1151));
    layer5_outputs(4001) <= layer4_outputs(5079);
    layer5_outputs(4002) <= (layer4_outputs(3545)) xor (layer4_outputs(1715));
    layer5_outputs(4003) <= not((layer4_outputs(4421)) xor (layer4_outputs(2614)));
    layer5_outputs(4004) <= layer4_outputs(2450);
    layer5_outputs(4005) <= '1';
    layer5_outputs(4006) <= not(layer4_outputs(740));
    layer5_outputs(4007) <= not((layer4_outputs(1951)) and (layer4_outputs(4620)));
    layer5_outputs(4008) <= layer4_outputs(1367);
    layer5_outputs(4009) <= not(layer4_outputs(116));
    layer5_outputs(4010) <= layer4_outputs(3704);
    layer5_outputs(4011) <= layer4_outputs(1215);
    layer5_outputs(4012) <= not(layer4_outputs(4783));
    layer5_outputs(4013) <= (layer4_outputs(3946)) or (layer4_outputs(1857));
    layer5_outputs(4014) <= not(layer4_outputs(5113));
    layer5_outputs(4015) <= layer4_outputs(3510);
    layer5_outputs(4016) <= (layer4_outputs(3070)) and not (layer4_outputs(2193));
    layer5_outputs(4017) <= layer4_outputs(4751);
    layer5_outputs(4018) <= (layer4_outputs(2285)) and not (layer4_outputs(4512));
    layer5_outputs(4019) <= layer4_outputs(2513);
    layer5_outputs(4020) <= layer4_outputs(4450);
    layer5_outputs(4021) <= not((layer4_outputs(1344)) and (layer4_outputs(2449)));
    layer5_outputs(4022) <= not(layer4_outputs(4132));
    layer5_outputs(4023) <= (layer4_outputs(466)) and not (layer4_outputs(3563));
    layer5_outputs(4024) <= layer4_outputs(1943);
    layer5_outputs(4025) <= not(layer4_outputs(4098));
    layer5_outputs(4026) <= (layer4_outputs(438)) and (layer4_outputs(2156));
    layer5_outputs(4027) <= not(layer4_outputs(831));
    layer5_outputs(4028) <= (layer4_outputs(1441)) or (layer4_outputs(3273));
    layer5_outputs(4029) <= not(layer4_outputs(4910)) or (layer4_outputs(4550));
    layer5_outputs(4030) <= not(layer4_outputs(4214)) or (layer4_outputs(338));
    layer5_outputs(4031) <= layer4_outputs(22);
    layer5_outputs(4032) <= not(layer4_outputs(4500));
    layer5_outputs(4033) <= not(layer4_outputs(636)) or (layer4_outputs(1084));
    layer5_outputs(4034) <= '1';
    layer5_outputs(4035) <= '1';
    layer5_outputs(4036) <= layer4_outputs(1127);
    layer5_outputs(4037) <= not(layer4_outputs(2317)) or (layer4_outputs(4555));
    layer5_outputs(4038) <= not(layer4_outputs(279));
    layer5_outputs(4039) <= not(layer4_outputs(3437));
    layer5_outputs(4040) <= layer4_outputs(4622);
    layer5_outputs(4041) <= not((layer4_outputs(3376)) and (layer4_outputs(4764)));
    layer5_outputs(4042) <= layer4_outputs(1687);
    layer5_outputs(4043) <= (layer4_outputs(4783)) and not (layer4_outputs(1117));
    layer5_outputs(4044) <= layer4_outputs(1834);
    layer5_outputs(4045) <= layer4_outputs(3220);
    layer5_outputs(4046) <= (layer4_outputs(1894)) and not (layer4_outputs(2997));
    layer5_outputs(4047) <= (layer4_outputs(4619)) or (layer4_outputs(4190));
    layer5_outputs(4048) <= not(layer4_outputs(884)) or (layer4_outputs(4877));
    layer5_outputs(4049) <= not(layer4_outputs(2876));
    layer5_outputs(4050) <= (layer4_outputs(3537)) xor (layer4_outputs(4266));
    layer5_outputs(4051) <= (layer4_outputs(1437)) or (layer4_outputs(2553));
    layer5_outputs(4052) <= layer4_outputs(953);
    layer5_outputs(4053) <= not(layer4_outputs(4612)) or (layer4_outputs(3879));
    layer5_outputs(4054) <= not(layer4_outputs(4532));
    layer5_outputs(4055) <= (layer4_outputs(3523)) and not (layer4_outputs(2703));
    layer5_outputs(4056) <= layer4_outputs(2654);
    layer5_outputs(4057) <= (layer4_outputs(2992)) and (layer4_outputs(2134));
    layer5_outputs(4058) <= layer4_outputs(2940);
    layer5_outputs(4059) <= not(layer4_outputs(679));
    layer5_outputs(4060) <= (layer4_outputs(602)) and (layer4_outputs(4030));
    layer5_outputs(4061) <= layer4_outputs(4542);
    layer5_outputs(4062) <= layer4_outputs(2500);
    layer5_outputs(4063) <= (layer4_outputs(663)) and not (layer4_outputs(4422));
    layer5_outputs(4064) <= not(layer4_outputs(2215));
    layer5_outputs(4065) <= not(layer4_outputs(2499));
    layer5_outputs(4066) <= not(layer4_outputs(2659)) or (layer4_outputs(1646));
    layer5_outputs(4067) <= not((layer4_outputs(705)) and (layer4_outputs(3374)));
    layer5_outputs(4068) <= not(layer4_outputs(5108));
    layer5_outputs(4069) <= (layer4_outputs(3011)) or (layer4_outputs(2469));
    layer5_outputs(4070) <= not(layer4_outputs(948));
    layer5_outputs(4071) <= (layer4_outputs(4170)) and (layer4_outputs(2366));
    layer5_outputs(4072) <= layer4_outputs(2258);
    layer5_outputs(4073) <= (layer4_outputs(1105)) xor (layer4_outputs(453));
    layer5_outputs(4074) <= (layer4_outputs(2899)) and (layer4_outputs(3299));
    layer5_outputs(4075) <= (layer4_outputs(927)) and (layer4_outputs(2958));
    layer5_outputs(4076) <= not((layer4_outputs(642)) and (layer4_outputs(4231)));
    layer5_outputs(4077) <= not(layer4_outputs(4557));
    layer5_outputs(4078) <= layer4_outputs(2668);
    layer5_outputs(4079) <= not(layer4_outputs(3619));
    layer5_outputs(4080) <= layer4_outputs(496);
    layer5_outputs(4081) <= layer4_outputs(3050);
    layer5_outputs(4082) <= not(layer4_outputs(2236));
    layer5_outputs(4083) <= layer4_outputs(4856);
    layer5_outputs(4084) <= layer4_outputs(4508);
    layer5_outputs(4085) <= not(layer4_outputs(1018));
    layer5_outputs(4086) <= (layer4_outputs(4055)) and (layer4_outputs(3950));
    layer5_outputs(4087) <= not((layer4_outputs(1863)) or (layer4_outputs(4907)));
    layer5_outputs(4088) <= (layer4_outputs(1685)) and not (layer4_outputs(745));
    layer5_outputs(4089) <= layer4_outputs(2888);
    layer5_outputs(4090) <= '1';
    layer5_outputs(4091) <= not(layer4_outputs(107));
    layer5_outputs(4092) <= not(layer4_outputs(2427));
    layer5_outputs(4093) <= layer4_outputs(3069);
    layer5_outputs(4094) <= layer4_outputs(2340);
    layer5_outputs(4095) <= not(layer4_outputs(411));
    layer5_outputs(4096) <= not(layer4_outputs(896)) or (layer4_outputs(5062));
    layer5_outputs(4097) <= (layer4_outputs(1218)) and not (layer4_outputs(3683));
    layer5_outputs(4098) <= (layer4_outputs(1287)) or (layer4_outputs(2263));
    layer5_outputs(4099) <= not(layer4_outputs(186)) or (layer4_outputs(4592));
    layer5_outputs(4100) <= not(layer4_outputs(2536));
    layer5_outputs(4101) <= (layer4_outputs(2040)) and not (layer4_outputs(1073));
    layer5_outputs(4102) <= (layer4_outputs(3713)) and (layer4_outputs(338));
    layer5_outputs(4103) <= not(layer4_outputs(4458));
    layer5_outputs(4104) <= not((layer4_outputs(3868)) xor (layer4_outputs(3238)));
    layer5_outputs(4105) <= not(layer4_outputs(1452));
    layer5_outputs(4106) <= layer4_outputs(2880);
    layer5_outputs(4107) <= layer4_outputs(3353);
    layer5_outputs(4108) <= layer4_outputs(926);
    layer5_outputs(4109) <= not(layer4_outputs(311)) or (layer4_outputs(4463));
    layer5_outputs(4110) <= not(layer4_outputs(1755));
    layer5_outputs(4111) <= layer4_outputs(1763);
    layer5_outputs(4112) <= layer4_outputs(2572);
    layer5_outputs(4113) <= not(layer4_outputs(4734));
    layer5_outputs(4114) <= layer4_outputs(2986);
    layer5_outputs(4115) <= not(layer4_outputs(2379)) or (layer4_outputs(4664));
    layer5_outputs(4116) <= layer4_outputs(1395);
    layer5_outputs(4117) <= not((layer4_outputs(1741)) xor (layer4_outputs(3853)));
    layer5_outputs(4118) <= layer4_outputs(3577);
    layer5_outputs(4119) <= not(layer4_outputs(3143));
    layer5_outputs(4120) <= not((layer4_outputs(140)) xor (layer4_outputs(2580)));
    layer5_outputs(4121) <= not((layer4_outputs(3552)) or (layer4_outputs(3948)));
    layer5_outputs(4122) <= not((layer4_outputs(1646)) and (layer4_outputs(3696)));
    layer5_outputs(4123) <= (layer4_outputs(1449)) and not (layer4_outputs(3002));
    layer5_outputs(4124) <= layer4_outputs(3915);
    layer5_outputs(4125) <= not((layer4_outputs(49)) xor (layer4_outputs(825)));
    layer5_outputs(4126) <= not(layer4_outputs(985)) or (layer4_outputs(3763));
    layer5_outputs(4127) <= not((layer4_outputs(1051)) xor (layer4_outputs(3568)));
    layer5_outputs(4128) <= (layer4_outputs(2799)) or (layer4_outputs(1195));
    layer5_outputs(4129) <= layer4_outputs(2684);
    layer5_outputs(4130) <= (layer4_outputs(2639)) and not (layer4_outputs(2192));
    layer5_outputs(4131) <= layer4_outputs(3758);
    layer5_outputs(4132) <= (layer4_outputs(436)) and not (layer4_outputs(1396));
    layer5_outputs(4133) <= not((layer4_outputs(4945)) and (layer4_outputs(2301)));
    layer5_outputs(4134) <= layer4_outputs(3064);
    layer5_outputs(4135) <= layer4_outputs(132);
    layer5_outputs(4136) <= (layer4_outputs(2002)) xor (layer4_outputs(277));
    layer5_outputs(4137) <= not((layer4_outputs(145)) xor (layer4_outputs(622)));
    layer5_outputs(4138) <= not((layer4_outputs(4506)) or (layer4_outputs(378)));
    layer5_outputs(4139) <= not((layer4_outputs(1774)) or (layer4_outputs(2950)));
    layer5_outputs(4140) <= not((layer4_outputs(1277)) or (layer4_outputs(3492)));
    layer5_outputs(4141) <= not(layer4_outputs(2429)) or (layer4_outputs(1417));
    layer5_outputs(4142) <= not(layer4_outputs(4708));
    layer5_outputs(4143) <= layer4_outputs(5038);
    layer5_outputs(4144) <= layer4_outputs(1599);
    layer5_outputs(4145) <= not(layer4_outputs(1893));
    layer5_outputs(4146) <= (layer4_outputs(2448)) and (layer4_outputs(857));
    layer5_outputs(4147) <= not(layer4_outputs(5076));
    layer5_outputs(4148) <= (layer4_outputs(4808)) and not (layer4_outputs(1837));
    layer5_outputs(4149) <= (layer4_outputs(4447)) and not (layer4_outputs(3004));
    layer5_outputs(4150) <= not(layer4_outputs(5089));
    layer5_outputs(4151) <= layer4_outputs(779);
    layer5_outputs(4152) <= layer4_outputs(2735);
    layer5_outputs(4153) <= not(layer4_outputs(4025));
    layer5_outputs(4154) <= (layer4_outputs(3815)) and (layer4_outputs(473));
    layer5_outputs(4155) <= not(layer4_outputs(3517));
    layer5_outputs(4156) <= not(layer4_outputs(4443));
    layer5_outputs(4157) <= (layer4_outputs(2017)) xor (layer4_outputs(751));
    layer5_outputs(4158) <= not(layer4_outputs(1650)) or (layer4_outputs(1026));
    layer5_outputs(4159) <= layer4_outputs(1134);
    layer5_outputs(4160) <= (layer4_outputs(1584)) or (layer4_outputs(1252));
    layer5_outputs(4161) <= (layer4_outputs(4651)) and not (layer4_outputs(5074));
    layer5_outputs(4162) <= (layer4_outputs(1220)) and not (layer4_outputs(2716));
    layer5_outputs(4163) <= (layer4_outputs(200)) and not (layer4_outputs(2501));
    layer5_outputs(4164) <= layer4_outputs(594);
    layer5_outputs(4165) <= not(layer4_outputs(2304)) or (layer4_outputs(3895));
    layer5_outputs(4166) <= '1';
    layer5_outputs(4167) <= not((layer4_outputs(2319)) or (layer4_outputs(1724)));
    layer5_outputs(4168) <= layer4_outputs(1428);
    layer5_outputs(4169) <= layer4_outputs(865);
    layer5_outputs(4170) <= layer4_outputs(3932);
    layer5_outputs(4171) <= '0';
    layer5_outputs(4172) <= layer4_outputs(1728);
    layer5_outputs(4173) <= not(layer4_outputs(4429));
    layer5_outputs(4174) <= not(layer4_outputs(2707));
    layer5_outputs(4175) <= '0';
    layer5_outputs(4176) <= layer4_outputs(1699);
    layer5_outputs(4177) <= not(layer4_outputs(4838));
    layer5_outputs(4178) <= (layer4_outputs(2564)) and (layer4_outputs(3248));
    layer5_outputs(4179) <= not((layer4_outputs(1256)) xor (layer4_outputs(2305)));
    layer5_outputs(4180) <= not(layer4_outputs(3305)) or (layer4_outputs(4109));
    layer5_outputs(4181) <= not(layer4_outputs(940));
    layer5_outputs(4182) <= (layer4_outputs(2580)) and (layer4_outputs(954));
    layer5_outputs(4183) <= not(layer4_outputs(720));
    layer5_outputs(4184) <= not(layer4_outputs(2073));
    layer5_outputs(4185) <= layer4_outputs(2850);
    layer5_outputs(4186) <= '1';
    layer5_outputs(4187) <= not((layer4_outputs(68)) and (layer4_outputs(4500)));
    layer5_outputs(4188) <= (layer4_outputs(517)) or (layer4_outputs(4047));
    layer5_outputs(4189) <= layer4_outputs(3897);
    layer5_outputs(4190) <= (layer4_outputs(3776)) xor (layer4_outputs(1229));
    layer5_outputs(4191) <= not(layer4_outputs(1139)) or (layer4_outputs(1138));
    layer5_outputs(4192) <= (layer4_outputs(3529)) and not (layer4_outputs(557));
    layer5_outputs(4193) <= (layer4_outputs(2479)) xor (layer4_outputs(2296));
    layer5_outputs(4194) <= not((layer4_outputs(482)) xor (layer4_outputs(2300)));
    layer5_outputs(4195) <= '0';
    layer5_outputs(4196) <= not(layer4_outputs(2652));
    layer5_outputs(4197) <= (layer4_outputs(2183)) and not (layer4_outputs(3481));
    layer5_outputs(4198) <= not((layer4_outputs(3734)) xor (layer4_outputs(4264)));
    layer5_outputs(4199) <= (layer4_outputs(4570)) and not (layer4_outputs(833));
    layer5_outputs(4200) <= not(layer4_outputs(593));
    layer5_outputs(4201) <= layer4_outputs(3055);
    layer5_outputs(4202) <= layer4_outputs(1907);
    layer5_outputs(4203) <= (layer4_outputs(213)) xor (layer4_outputs(2274));
    layer5_outputs(4204) <= (layer4_outputs(356)) and not (layer4_outputs(1109));
    layer5_outputs(4205) <= layer4_outputs(4015);
    layer5_outputs(4206) <= '1';
    layer5_outputs(4207) <= not((layer4_outputs(5013)) xor (layer4_outputs(493)));
    layer5_outputs(4208) <= not(layer4_outputs(2813));
    layer5_outputs(4209) <= not(layer4_outputs(2610));
    layer5_outputs(4210) <= not((layer4_outputs(2369)) and (layer4_outputs(4222)));
    layer5_outputs(4211) <= layer4_outputs(1021);
    layer5_outputs(4212) <= not(layer4_outputs(825));
    layer5_outputs(4213) <= layer4_outputs(1495);
    layer5_outputs(4214) <= not(layer4_outputs(3139));
    layer5_outputs(4215) <= not(layer4_outputs(485));
    layer5_outputs(4216) <= not(layer4_outputs(4972));
    layer5_outputs(4217) <= layer4_outputs(3356);
    layer5_outputs(4218) <= layer4_outputs(1227);
    layer5_outputs(4219) <= not(layer4_outputs(3287));
    layer5_outputs(4220) <= not((layer4_outputs(3168)) or (layer4_outputs(4032)));
    layer5_outputs(4221) <= not((layer4_outputs(3913)) or (layer4_outputs(376)));
    layer5_outputs(4222) <= not(layer4_outputs(3209));
    layer5_outputs(4223) <= (layer4_outputs(937)) and (layer4_outputs(2943));
    layer5_outputs(4224) <= not(layer4_outputs(3572));
    layer5_outputs(4225) <= (layer4_outputs(2151)) and (layer4_outputs(3828));
    layer5_outputs(4226) <= not((layer4_outputs(4353)) and (layer4_outputs(3118)));
    layer5_outputs(4227) <= layer4_outputs(981);
    layer5_outputs(4228) <= not(layer4_outputs(3925));
    layer5_outputs(4229) <= layer4_outputs(2958);
    layer5_outputs(4230) <= layer4_outputs(715);
    layer5_outputs(4231) <= not(layer4_outputs(3373));
    layer5_outputs(4232) <= (layer4_outputs(2535)) and not (layer4_outputs(3354));
    layer5_outputs(4233) <= not(layer4_outputs(2025));
    layer5_outputs(4234) <= (layer4_outputs(4507)) and not (layer4_outputs(2888));
    layer5_outputs(4235) <= layer4_outputs(1446);
    layer5_outputs(4236) <= layer4_outputs(968);
    layer5_outputs(4237) <= layer4_outputs(1109);
    layer5_outputs(4238) <= not(layer4_outputs(3596));
    layer5_outputs(4239) <= layer4_outputs(2741);
    layer5_outputs(4240) <= not((layer4_outputs(693)) and (layer4_outputs(4926)));
    layer5_outputs(4241) <= not(layer4_outputs(3366));
    layer5_outputs(4242) <= not(layer4_outputs(4870));
    layer5_outputs(4243) <= not(layer4_outputs(1685));
    layer5_outputs(4244) <= layer4_outputs(4368);
    layer5_outputs(4245) <= (layer4_outputs(2020)) or (layer4_outputs(4014));
    layer5_outputs(4246) <= not(layer4_outputs(1629));
    layer5_outputs(4247) <= not((layer4_outputs(3080)) or (layer4_outputs(3735)));
    layer5_outputs(4248) <= not(layer4_outputs(4807)) or (layer4_outputs(4146));
    layer5_outputs(4249) <= (layer4_outputs(3246)) and not (layer4_outputs(4297));
    layer5_outputs(4250) <= not(layer4_outputs(3161));
    layer5_outputs(4251) <= layer4_outputs(4569);
    layer5_outputs(4252) <= not(layer4_outputs(3010)) or (layer4_outputs(995));
    layer5_outputs(4253) <= layer4_outputs(597);
    layer5_outputs(4254) <= not((layer4_outputs(3238)) and (layer4_outputs(352)));
    layer5_outputs(4255) <= (layer4_outputs(4929)) and (layer4_outputs(1073));
    layer5_outputs(4256) <= not(layer4_outputs(526));
    layer5_outputs(4257) <= (layer4_outputs(3024)) and (layer4_outputs(3662));
    layer5_outputs(4258) <= not((layer4_outputs(1920)) and (layer4_outputs(571)));
    layer5_outputs(4259) <= (layer4_outputs(2113)) and not (layer4_outputs(3665));
    layer5_outputs(4260) <= layer4_outputs(2670);
    layer5_outputs(4261) <= not((layer4_outputs(2533)) xor (layer4_outputs(3954)));
    layer5_outputs(4262) <= not(layer4_outputs(4793)) or (layer4_outputs(33));
    layer5_outputs(4263) <= not(layer4_outputs(1485)) or (layer4_outputs(2189));
    layer5_outputs(4264) <= (layer4_outputs(3829)) and not (layer4_outputs(540));
    layer5_outputs(4265) <= not(layer4_outputs(3713));
    layer5_outputs(4266) <= layer4_outputs(2227);
    layer5_outputs(4267) <= (layer4_outputs(4388)) xor (layer4_outputs(2550));
    layer5_outputs(4268) <= (layer4_outputs(3001)) and (layer4_outputs(4498));
    layer5_outputs(4269) <= not(layer4_outputs(1340));
    layer5_outputs(4270) <= not(layer4_outputs(4880));
    layer5_outputs(4271) <= layer4_outputs(467);
    layer5_outputs(4272) <= layer4_outputs(94);
    layer5_outputs(4273) <= layer4_outputs(3901);
    layer5_outputs(4274) <= not((layer4_outputs(3019)) or (layer4_outputs(941)));
    layer5_outputs(4275) <= not(layer4_outputs(1981));
    layer5_outputs(4276) <= (layer4_outputs(358)) and not (layer4_outputs(1835));
    layer5_outputs(4277) <= (layer4_outputs(296)) or (layer4_outputs(4574));
    layer5_outputs(4278) <= (layer4_outputs(19)) xor (layer4_outputs(2498));
    layer5_outputs(4279) <= not(layer4_outputs(729));
    layer5_outputs(4280) <= not(layer4_outputs(815));
    layer5_outputs(4281) <= (layer4_outputs(2841)) or (layer4_outputs(811));
    layer5_outputs(4282) <= layer4_outputs(1537);
    layer5_outputs(4283) <= not(layer4_outputs(2026));
    layer5_outputs(4284) <= (layer4_outputs(3749)) and not (layer4_outputs(102));
    layer5_outputs(4285) <= not(layer4_outputs(2905)) or (layer4_outputs(4361));
    layer5_outputs(4286) <= not(layer4_outputs(969));
    layer5_outputs(4287) <= not(layer4_outputs(3804));
    layer5_outputs(4288) <= not((layer4_outputs(3382)) xor (layer4_outputs(4077)));
    layer5_outputs(4289) <= (layer4_outputs(4143)) xor (layer4_outputs(2118));
    layer5_outputs(4290) <= not((layer4_outputs(538)) xor (layer4_outputs(3012)));
    layer5_outputs(4291) <= '1';
    layer5_outputs(4292) <= not(layer4_outputs(2687));
    layer5_outputs(4293) <= layer4_outputs(1771);
    layer5_outputs(4294) <= (layer4_outputs(4558)) and (layer4_outputs(1414));
    layer5_outputs(4295) <= not(layer4_outputs(955)) or (layer4_outputs(1544));
    layer5_outputs(4296) <= layer4_outputs(1964);
    layer5_outputs(4297) <= not((layer4_outputs(1647)) and (layer4_outputs(3644)));
    layer5_outputs(4298) <= not(layer4_outputs(1525));
    layer5_outputs(4299) <= (layer4_outputs(1154)) and not (layer4_outputs(4518));
    layer5_outputs(4300) <= layer4_outputs(429);
    layer5_outputs(4301) <= not(layer4_outputs(830));
    layer5_outputs(4302) <= (layer4_outputs(319)) and (layer4_outputs(1288));
    layer5_outputs(4303) <= not((layer4_outputs(251)) or (layer4_outputs(10)));
    layer5_outputs(4304) <= layer4_outputs(590);
    layer5_outputs(4305) <= (layer4_outputs(4789)) and (layer4_outputs(1005));
    layer5_outputs(4306) <= not((layer4_outputs(3588)) and (layer4_outputs(323)));
    layer5_outputs(4307) <= (layer4_outputs(3215)) and (layer4_outputs(2526));
    layer5_outputs(4308) <= (layer4_outputs(2759)) and not (layer4_outputs(776));
    layer5_outputs(4309) <= (layer4_outputs(2583)) xor (layer4_outputs(3634));
    layer5_outputs(4310) <= not((layer4_outputs(2418)) or (layer4_outputs(344)));
    layer5_outputs(4311) <= not(layer4_outputs(2725)) or (layer4_outputs(881));
    layer5_outputs(4312) <= not(layer4_outputs(719)) or (layer4_outputs(3325));
    layer5_outputs(4313) <= not(layer4_outputs(3644));
    layer5_outputs(4314) <= layer4_outputs(2965);
    layer5_outputs(4315) <= not((layer4_outputs(3294)) xor (layer4_outputs(4614)));
    layer5_outputs(4316) <= layer4_outputs(1965);
    layer5_outputs(4317) <= not(layer4_outputs(1386)) or (layer4_outputs(2789));
    layer5_outputs(4318) <= layer4_outputs(3704);
    layer5_outputs(4319) <= not((layer4_outputs(2785)) or (layer4_outputs(3513)));
    layer5_outputs(4320) <= layer4_outputs(70);
    layer5_outputs(4321) <= (layer4_outputs(4847)) and not (layer4_outputs(888));
    layer5_outputs(4322) <= layer4_outputs(879);
    layer5_outputs(4323) <= '0';
    layer5_outputs(4324) <= layer4_outputs(2219);
    layer5_outputs(4325) <= layer4_outputs(3884);
    layer5_outputs(4326) <= layer4_outputs(47);
    layer5_outputs(4327) <= not(layer4_outputs(3174));
    layer5_outputs(4328) <= not(layer4_outputs(3167));
    layer5_outputs(4329) <= not((layer4_outputs(649)) xor (layer4_outputs(4005)));
    layer5_outputs(4330) <= layer4_outputs(4868);
    layer5_outputs(4331) <= not((layer4_outputs(602)) and (layer4_outputs(1648)));
    layer5_outputs(4332) <= layer4_outputs(3356);
    layer5_outputs(4333) <= not((layer4_outputs(3508)) xor (layer4_outputs(3035)));
    layer5_outputs(4334) <= not(layer4_outputs(4400));
    layer5_outputs(4335) <= (layer4_outputs(3506)) or (layer4_outputs(205));
    layer5_outputs(4336) <= not((layer4_outputs(4646)) or (layer4_outputs(2868)));
    layer5_outputs(4337) <= layer4_outputs(444);
    layer5_outputs(4338) <= '1';
    layer5_outputs(4339) <= not((layer4_outputs(4078)) or (layer4_outputs(3918)));
    layer5_outputs(4340) <= not(layer4_outputs(842));
    layer5_outputs(4341) <= not(layer4_outputs(2462)) or (layer4_outputs(3316));
    layer5_outputs(4342) <= '1';
    layer5_outputs(4343) <= (layer4_outputs(2080)) and not (layer4_outputs(4454));
    layer5_outputs(4344) <= (layer4_outputs(687)) and not (layer4_outputs(928));
    layer5_outputs(4345) <= (layer4_outputs(530)) xor (layer4_outputs(261));
    layer5_outputs(4346) <= layer4_outputs(4571);
    layer5_outputs(4347) <= (layer4_outputs(3319)) xor (layer4_outputs(3745));
    layer5_outputs(4348) <= (layer4_outputs(2939)) and not (layer4_outputs(494));
    layer5_outputs(4349) <= layer4_outputs(4173);
    layer5_outputs(4350) <= not(layer4_outputs(2743));
    layer5_outputs(4351) <= layer4_outputs(1207);
    layer5_outputs(4352) <= not(layer4_outputs(3099)) or (layer4_outputs(3543));
    layer5_outputs(4353) <= (layer4_outputs(3971)) and not (layer4_outputs(1151));
    layer5_outputs(4354) <= (layer4_outputs(1257)) and not (layer4_outputs(1086));
    layer5_outputs(4355) <= not(layer4_outputs(774)) or (layer4_outputs(2003));
    layer5_outputs(4356) <= not(layer4_outputs(3272)) or (layer4_outputs(355));
    layer5_outputs(4357) <= not(layer4_outputs(5004)) or (layer4_outputs(1053));
    layer5_outputs(4358) <= layer4_outputs(873);
    layer5_outputs(4359) <= layer4_outputs(690);
    layer5_outputs(4360) <= not((layer4_outputs(104)) xor (layer4_outputs(4254)));
    layer5_outputs(4361) <= not((layer4_outputs(3834)) and (layer4_outputs(1248)));
    layer5_outputs(4362) <= not((layer4_outputs(4521)) or (layer4_outputs(4459)));
    layer5_outputs(4363) <= layer4_outputs(491);
    layer5_outputs(4364) <= '1';
    layer5_outputs(4365) <= not((layer4_outputs(2676)) xor (layer4_outputs(422)));
    layer5_outputs(4366) <= not(layer4_outputs(2328)) or (layer4_outputs(192));
    layer5_outputs(4367) <= (layer4_outputs(2528)) and not (layer4_outputs(2996));
    layer5_outputs(4368) <= (layer4_outputs(215)) and not (layer4_outputs(1309));
    layer5_outputs(4369) <= not((layer4_outputs(4897)) and (layer4_outputs(4640)));
    layer5_outputs(4370) <= not(layer4_outputs(5032));
    layer5_outputs(4371) <= not(layer4_outputs(589)) or (layer4_outputs(4171));
    layer5_outputs(4372) <= not((layer4_outputs(3209)) and (layer4_outputs(2983)));
    layer5_outputs(4373) <= (layer4_outputs(645)) xor (layer4_outputs(1570));
    layer5_outputs(4374) <= (layer4_outputs(204)) and not (layer4_outputs(2186));
    layer5_outputs(4375) <= not(layer4_outputs(435));
    layer5_outputs(4376) <= (layer4_outputs(2023)) and (layer4_outputs(1895));
    layer5_outputs(4377) <= layer4_outputs(447);
    layer5_outputs(4378) <= not(layer4_outputs(3922));
    layer5_outputs(4379) <= layer4_outputs(2589);
    layer5_outputs(4380) <= (layer4_outputs(4658)) and not (layer4_outputs(298));
    layer5_outputs(4381) <= (layer4_outputs(3598)) and (layer4_outputs(4784));
    layer5_outputs(4382) <= layer4_outputs(1948);
    layer5_outputs(4383) <= not(layer4_outputs(3744));
    layer5_outputs(4384) <= not(layer4_outputs(849)) or (layer4_outputs(3854));
    layer5_outputs(4385) <= layer4_outputs(1767);
    layer5_outputs(4386) <= layer4_outputs(435);
    layer5_outputs(4387) <= not((layer4_outputs(4187)) and (layer4_outputs(1547)));
    layer5_outputs(4388) <= not(layer4_outputs(4380));
    layer5_outputs(4389) <= not(layer4_outputs(908));
    layer5_outputs(4390) <= layer4_outputs(2232);
    layer5_outputs(4391) <= not(layer4_outputs(2485));
    layer5_outputs(4392) <= not(layer4_outputs(1437));
    layer5_outputs(4393) <= layer4_outputs(321);
    layer5_outputs(4394) <= layer4_outputs(570);
    layer5_outputs(4395) <= layer4_outputs(1503);
    layer5_outputs(4396) <= (layer4_outputs(380)) xor (layer4_outputs(1473));
    layer5_outputs(4397) <= not((layer4_outputs(558)) or (layer4_outputs(657)));
    layer5_outputs(4398) <= (layer4_outputs(3153)) xor (layer4_outputs(3067));
    layer5_outputs(4399) <= layer4_outputs(2775);
    layer5_outputs(4400) <= layer4_outputs(2894);
    layer5_outputs(4401) <= not((layer4_outputs(1953)) and (layer4_outputs(3383)));
    layer5_outputs(4402) <= not(layer4_outputs(4702)) or (layer4_outputs(1946));
    layer5_outputs(4403) <= not(layer4_outputs(5112));
    layer5_outputs(4404) <= not((layer4_outputs(4512)) and (layer4_outputs(1605)));
    layer5_outputs(4405) <= not((layer4_outputs(2782)) xor (layer4_outputs(1487)));
    layer5_outputs(4406) <= layer4_outputs(4836);
    layer5_outputs(4407) <= '0';
    layer5_outputs(4408) <= not(layer4_outputs(428));
    layer5_outputs(4409) <= not(layer4_outputs(2066)) or (layer4_outputs(1186));
    layer5_outputs(4410) <= layer4_outputs(573);
    layer5_outputs(4411) <= not((layer4_outputs(1508)) or (layer4_outputs(1235)));
    layer5_outputs(4412) <= not(layer4_outputs(3104));
    layer5_outputs(4413) <= not(layer4_outputs(3340));
    layer5_outputs(4414) <= not(layer4_outputs(1549)) or (layer4_outputs(2213));
    layer5_outputs(4415) <= (layer4_outputs(1775)) and not (layer4_outputs(2522));
    layer5_outputs(4416) <= (layer4_outputs(4637)) and not (layer4_outputs(4251));
    layer5_outputs(4417) <= not(layer4_outputs(1020));
    layer5_outputs(4418) <= (layer4_outputs(22)) and not (layer4_outputs(176));
    layer5_outputs(4419) <= not(layer4_outputs(267));
    layer5_outputs(4420) <= not(layer4_outputs(2945));
    layer5_outputs(4421) <= layer4_outputs(2461);
    layer5_outputs(4422) <= not(layer4_outputs(1237));
    layer5_outputs(4423) <= layer4_outputs(4260);
    layer5_outputs(4424) <= '1';
    layer5_outputs(4425) <= (layer4_outputs(2913)) xor (layer4_outputs(248));
    layer5_outputs(4426) <= '1';
    layer5_outputs(4427) <= layer4_outputs(5100);
    layer5_outputs(4428) <= (layer4_outputs(1577)) and (layer4_outputs(4366));
    layer5_outputs(4429) <= not(layer4_outputs(1922));
    layer5_outputs(4430) <= not((layer4_outputs(2808)) and (layer4_outputs(1223)));
    layer5_outputs(4431) <= layer4_outputs(1575);
    layer5_outputs(4432) <= '0';
    layer5_outputs(4433) <= (layer4_outputs(1582)) xor (layer4_outputs(4966));
    layer5_outputs(4434) <= not(layer4_outputs(3670));
    layer5_outputs(4435) <= not((layer4_outputs(3879)) and (layer4_outputs(4454)));
    layer5_outputs(4436) <= not((layer4_outputs(4295)) and (layer4_outputs(2160)));
    layer5_outputs(4437) <= layer4_outputs(3271);
    layer5_outputs(4438) <= layer4_outputs(1037);
    layer5_outputs(4439) <= not((layer4_outputs(1643)) and (layer4_outputs(1590)));
    layer5_outputs(4440) <= not(layer4_outputs(1797)) or (layer4_outputs(3292));
    layer5_outputs(4441) <= layer4_outputs(4406);
    layer5_outputs(4442) <= not(layer4_outputs(3518));
    layer5_outputs(4443) <= not(layer4_outputs(3270));
    layer5_outputs(4444) <= not(layer4_outputs(4638));
    layer5_outputs(4445) <= layer4_outputs(4267);
    layer5_outputs(4446) <= layer4_outputs(1296);
    layer5_outputs(4447) <= not(layer4_outputs(917)) or (layer4_outputs(1278));
    layer5_outputs(4448) <= not(layer4_outputs(1466));
    layer5_outputs(4449) <= not((layer4_outputs(4692)) or (layer4_outputs(4623)));
    layer5_outputs(4450) <= (layer4_outputs(193)) and (layer4_outputs(2166));
    layer5_outputs(4451) <= layer4_outputs(4535);
    layer5_outputs(4452) <= not((layer4_outputs(1956)) and (layer4_outputs(3219)));
    layer5_outputs(4453) <= layer4_outputs(4946);
    layer5_outputs(4454) <= layer4_outputs(2195);
    layer5_outputs(4455) <= (layer4_outputs(4145)) and (layer4_outputs(2673));
    layer5_outputs(4456) <= (layer4_outputs(2096)) xor (layer4_outputs(308));
    layer5_outputs(4457) <= not(layer4_outputs(3983));
    layer5_outputs(4458) <= not(layer4_outputs(2575));
    layer5_outputs(4459) <= not(layer4_outputs(4459)) or (layer4_outputs(3536));
    layer5_outputs(4460) <= not(layer4_outputs(1236));
    layer5_outputs(4461) <= not(layer4_outputs(2677)) or (layer4_outputs(870));
    layer5_outputs(4462) <= (layer4_outputs(4897)) and (layer4_outputs(1077));
    layer5_outputs(4463) <= (layer4_outputs(2225)) and not (layer4_outputs(1511));
    layer5_outputs(4464) <= not((layer4_outputs(4750)) or (layer4_outputs(1122)));
    layer5_outputs(4465) <= not(layer4_outputs(4456));
    layer5_outputs(4466) <= not((layer4_outputs(343)) or (layer4_outputs(1229)));
    layer5_outputs(4467) <= not(layer4_outputs(623));
    layer5_outputs(4468) <= (layer4_outputs(3251)) or (layer4_outputs(1851));
    layer5_outputs(4469) <= not(layer4_outputs(1403));
    layer5_outputs(4470) <= (layer4_outputs(4575)) xor (layer4_outputs(3370));
    layer5_outputs(4471) <= layer4_outputs(1180);
    layer5_outputs(4472) <= not(layer4_outputs(1316)) or (layer4_outputs(1571));
    layer5_outputs(4473) <= layer4_outputs(4901);
    layer5_outputs(4474) <= layer4_outputs(685);
    layer5_outputs(4475) <= layer4_outputs(1910);
    layer5_outputs(4476) <= not(layer4_outputs(936));
    layer5_outputs(4477) <= layer4_outputs(566);
    layer5_outputs(4478) <= (layer4_outputs(945)) xor (layer4_outputs(98));
    layer5_outputs(4479) <= (layer4_outputs(736)) xor (layer4_outputs(2038));
    layer5_outputs(4480) <= not(layer4_outputs(2414));
    layer5_outputs(4481) <= not((layer4_outputs(2805)) and (layer4_outputs(2657)));
    layer5_outputs(4482) <= not((layer4_outputs(1307)) or (layer4_outputs(3637)));
    layer5_outputs(4483) <= layer4_outputs(458);
    layer5_outputs(4484) <= not((layer4_outputs(1464)) and (layer4_outputs(4053)));
    layer5_outputs(4485) <= (layer4_outputs(4342)) or (layer4_outputs(3955));
    layer5_outputs(4486) <= not((layer4_outputs(4650)) xor (layer4_outputs(4107)));
    layer5_outputs(4487) <= not((layer4_outputs(1000)) and (layer4_outputs(3254)));
    layer5_outputs(4488) <= not(layer4_outputs(739)) or (layer4_outputs(1423));
    layer5_outputs(4489) <= not(layer4_outputs(3344)) or (layer4_outputs(3861));
    layer5_outputs(4490) <= (layer4_outputs(2593)) and not (layer4_outputs(1543));
    layer5_outputs(4491) <= layer4_outputs(4745);
    layer5_outputs(4492) <= not(layer4_outputs(4945));
    layer5_outputs(4493) <= not(layer4_outputs(4663));
    layer5_outputs(4494) <= not(layer4_outputs(4041)) or (layer4_outputs(2505));
    layer5_outputs(4495) <= not(layer4_outputs(2682));
    layer5_outputs(4496) <= (layer4_outputs(1541)) and (layer4_outputs(2017));
    layer5_outputs(4497) <= (layer4_outputs(178)) xor (layer4_outputs(1627));
    layer5_outputs(4498) <= (layer4_outputs(5097)) or (layer4_outputs(2110));
    layer5_outputs(4499) <= '0';
    layer5_outputs(4500) <= layer4_outputs(2511);
    layer5_outputs(4501) <= layer4_outputs(4713);
    layer5_outputs(4502) <= not(layer4_outputs(4335));
    layer5_outputs(4503) <= '1';
    layer5_outputs(4504) <= not((layer4_outputs(1990)) and (layer4_outputs(4004)));
    layer5_outputs(4505) <= not(layer4_outputs(1545));
    layer5_outputs(4506) <= not(layer4_outputs(1592));
    layer5_outputs(4507) <= layer4_outputs(3164);
    layer5_outputs(4508) <= layer4_outputs(712);
    layer5_outputs(4509) <= layer4_outputs(3994);
    layer5_outputs(4510) <= not(layer4_outputs(4998)) or (layer4_outputs(1091));
    layer5_outputs(4511) <= (layer4_outputs(177)) and not (layer4_outputs(1474));
    layer5_outputs(4512) <= not((layer4_outputs(415)) or (layer4_outputs(733)));
    layer5_outputs(4513) <= not(layer4_outputs(1163)) or (layer4_outputs(667));
    layer5_outputs(4514) <= not((layer4_outputs(1345)) and (layer4_outputs(2864)));
    layer5_outputs(4515) <= '0';
    layer5_outputs(4516) <= not(layer4_outputs(3393));
    layer5_outputs(4517) <= not((layer4_outputs(1082)) or (layer4_outputs(4723)));
    layer5_outputs(4518) <= layer4_outputs(2517);
    layer5_outputs(4519) <= not((layer4_outputs(4616)) xor (layer4_outputs(2490)));
    layer5_outputs(4520) <= (layer4_outputs(4013)) and not (layer4_outputs(1376));
    layer5_outputs(4521) <= not(layer4_outputs(1859));
    layer5_outputs(4522) <= layer4_outputs(1000);
    layer5_outputs(4523) <= (layer4_outputs(1675)) and not (layer4_outputs(2181));
    layer5_outputs(4524) <= (layer4_outputs(4012)) and not (layer4_outputs(1604));
    layer5_outputs(4525) <= not(layer4_outputs(795));
    layer5_outputs(4526) <= not(layer4_outputs(4657)) or (layer4_outputs(793));
    layer5_outputs(4527) <= not(layer4_outputs(1816));
    layer5_outputs(4528) <= not(layer4_outputs(1711));
    layer5_outputs(4529) <= '0';
    layer5_outputs(4530) <= layer4_outputs(281);
    layer5_outputs(4531) <= (layer4_outputs(4470)) and (layer4_outputs(3000));
    layer5_outputs(4532) <= layer4_outputs(2665);
    layer5_outputs(4533) <= not(layer4_outputs(416)) or (layer4_outputs(3131));
    layer5_outputs(4534) <= (layer4_outputs(3487)) xor (layer4_outputs(1966));
    layer5_outputs(4535) <= layer4_outputs(1301);
    layer5_outputs(4536) <= not(layer4_outputs(1892));
    layer5_outputs(4537) <= not(layer4_outputs(4865)) or (layer4_outputs(844));
    layer5_outputs(4538) <= (layer4_outputs(4531)) or (layer4_outputs(232));
    layer5_outputs(4539) <= not(layer4_outputs(5096));
    layer5_outputs(4540) <= not(layer4_outputs(4075)) or (layer4_outputs(4402));
    layer5_outputs(4541) <= layer4_outputs(3485);
    layer5_outputs(4542) <= not((layer4_outputs(1827)) xor (layer4_outputs(4334)));
    layer5_outputs(4543) <= (layer4_outputs(503)) and not (layer4_outputs(2018));
    layer5_outputs(4544) <= layer4_outputs(2098);
    layer5_outputs(4545) <= (layer4_outputs(4916)) and (layer4_outputs(476));
    layer5_outputs(4546) <= not(layer4_outputs(600));
    layer5_outputs(4547) <= layer4_outputs(4533);
    layer5_outputs(4548) <= '0';
    layer5_outputs(4549) <= not(layer4_outputs(458));
    layer5_outputs(4550) <= layer4_outputs(4428);
    layer5_outputs(4551) <= not(layer4_outputs(932));
    layer5_outputs(4552) <= (layer4_outputs(1984)) and not (layer4_outputs(545));
    layer5_outputs(4553) <= layer4_outputs(1141);
    layer5_outputs(4554) <= (layer4_outputs(723)) and not (layer4_outputs(2720));
    layer5_outputs(4555) <= (layer4_outputs(341)) and (layer4_outputs(4599));
    layer5_outputs(4556) <= not(layer4_outputs(161)) or (layer4_outputs(3480));
    layer5_outputs(4557) <= not(layer4_outputs(2381));
    layer5_outputs(4558) <= (layer4_outputs(3226)) and not (layer4_outputs(4178));
    layer5_outputs(4559) <= not(layer4_outputs(1678));
    layer5_outputs(4560) <= (layer4_outputs(2398)) and not (layer4_outputs(3495));
    layer5_outputs(4561) <= not(layer4_outputs(2870));
    layer5_outputs(4562) <= (layer4_outputs(2660)) and not (layer4_outputs(1241));
    layer5_outputs(4563) <= not(layer4_outputs(5004));
    layer5_outputs(4564) <= not(layer4_outputs(1548));
    layer5_outputs(4565) <= (layer4_outputs(505)) xor (layer4_outputs(3233));
    layer5_outputs(4566) <= layer4_outputs(5015);
    layer5_outputs(4567) <= layer4_outputs(5067);
    layer5_outputs(4568) <= not(layer4_outputs(2561)) or (layer4_outputs(1543));
    layer5_outputs(4569) <= not(layer4_outputs(416));
    layer5_outputs(4570) <= layer4_outputs(881);
    layer5_outputs(4571) <= not(layer4_outputs(1398));
    layer5_outputs(4572) <= not(layer4_outputs(4762));
    layer5_outputs(4573) <= not((layer4_outputs(912)) and (layer4_outputs(3055)));
    layer5_outputs(4574) <= not(layer4_outputs(2692));
    layer5_outputs(4575) <= (layer4_outputs(3030)) or (layer4_outputs(3033));
    layer5_outputs(4576) <= not(layer4_outputs(3023));
    layer5_outputs(4577) <= not(layer4_outputs(4754)) or (layer4_outputs(981));
    layer5_outputs(4578) <= (layer4_outputs(266)) and not (layer4_outputs(2059));
    layer5_outputs(4579) <= layer4_outputs(3431);
    layer5_outputs(4580) <= not((layer4_outputs(1665)) xor (layer4_outputs(1005)));
    layer5_outputs(4581) <= not((layer4_outputs(1693)) and (layer4_outputs(1830)));
    layer5_outputs(4582) <= (layer4_outputs(1512)) or (layer4_outputs(4642));
    layer5_outputs(4583) <= layer4_outputs(29);
    layer5_outputs(4584) <= (layer4_outputs(337)) and (layer4_outputs(3122));
    layer5_outputs(4585) <= not(layer4_outputs(315));
    layer5_outputs(4586) <= not(layer4_outputs(2963));
    layer5_outputs(4587) <= '0';
    layer5_outputs(4588) <= (layer4_outputs(3054)) and not (layer4_outputs(4810));
    layer5_outputs(4589) <= not(layer4_outputs(3778)) or (layer4_outputs(1710));
    layer5_outputs(4590) <= not((layer4_outputs(3113)) or (layer4_outputs(954)));
    layer5_outputs(4591) <= (layer4_outputs(3882)) or (layer4_outputs(1304));
    layer5_outputs(4592) <= not(layer4_outputs(3495)) or (layer4_outputs(512));
    layer5_outputs(4593) <= not((layer4_outputs(2162)) or (layer4_outputs(883)));
    layer5_outputs(4594) <= (layer4_outputs(1562)) and not (layer4_outputs(252));
    layer5_outputs(4595) <= not(layer4_outputs(490)) or (layer4_outputs(2377));
    layer5_outputs(4596) <= (layer4_outputs(60)) and (layer4_outputs(4663));
    layer5_outputs(4597) <= not(layer4_outputs(4643)) or (layer4_outputs(3177));
    layer5_outputs(4598) <= (layer4_outputs(3460)) and not (layer4_outputs(486));
    layer5_outputs(4599) <= not(layer4_outputs(2079));
    layer5_outputs(4600) <= not(layer4_outputs(4104));
    layer5_outputs(4601) <= (layer4_outputs(2228)) or (layer4_outputs(1597));
    layer5_outputs(4602) <= not(layer4_outputs(1462));
    layer5_outputs(4603) <= layer4_outputs(2657);
    layer5_outputs(4604) <= (layer4_outputs(3029)) and (layer4_outputs(3519));
    layer5_outputs(4605) <= not((layer4_outputs(2022)) and (layer4_outputs(3995)));
    layer5_outputs(4606) <= not(layer4_outputs(2349));
    layer5_outputs(4607) <= layer4_outputs(5078);
    layer5_outputs(4608) <= (layer4_outputs(1587)) and not (layer4_outputs(1989));
    layer5_outputs(4609) <= not(layer4_outputs(4039));
    layer5_outputs(4610) <= not(layer4_outputs(3450));
    layer5_outputs(4611) <= (layer4_outputs(2563)) and not (layer4_outputs(1773));
    layer5_outputs(4612) <= layer4_outputs(4981);
    layer5_outputs(4613) <= layer4_outputs(2410);
    layer5_outputs(4614) <= layer4_outputs(3202);
    layer5_outputs(4615) <= not(layer4_outputs(1938)) or (layer4_outputs(4149));
    layer5_outputs(4616) <= (layer4_outputs(2574)) and not (layer4_outputs(2127));
    layer5_outputs(4617) <= not(layer4_outputs(3735)) or (layer4_outputs(1068));
    layer5_outputs(4618) <= (layer4_outputs(2887)) xor (layer4_outputs(5081));
    layer5_outputs(4619) <= not(layer4_outputs(4221)) or (layer4_outputs(1804));
    layer5_outputs(4620) <= (layer4_outputs(2939)) and not (layer4_outputs(4155));
    layer5_outputs(4621) <= layer4_outputs(3494);
    layer5_outputs(4622) <= (layer4_outputs(661)) xor (layer4_outputs(3191));
    layer5_outputs(4623) <= not(layer4_outputs(656));
    layer5_outputs(4624) <= not(layer4_outputs(4425));
    layer5_outputs(4625) <= (layer4_outputs(5020)) xor (layer4_outputs(3227));
    layer5_outputs(4626) <= not(layer4_outputs(3498));
    layer5_outputs(4627) <= not(layer4_outputs(3833));
    layer5_outputs(4628) <= not((layer4_outputs(5085)) or (layer4_outputs(959)));
    layer5_outputs(4629) <= (layer4_outputs(3217)) and (layer4_outputs(4421));
    layer5_outputs(4630) <= layer4_outputs(4829);
    layer5_outputs(4631) <= (layer4_outputs(4230)) xor (layer4_outputs(1362));
    layer5_outputs(4632) <= (layer4_outputs(2270)) and not (layer4_outputs(4842));
    layer5_outputs(4633) <= layer4_outputs(4331);
    layer5_outputs(4634) <= not(layer4_outputs(4200));
    layer5_outputs(4635) <= not((layer4_outputs(4678)) or (layer4_outputs(473)));
    layer5_outputs(4636) <= (layer4_outputs(1010)) xor (layer4_outputs(2617));
    layer5_outputs(4637) <= not(layer4_outputs(2049));
    layer5_outputs(4638) <= not((layer4_outputs(2124)) and (layer4_outputs(972)));
    layer5_outputs(4639) <= layer4_outputs(3301);
    layer5_outputs(4640) <= not((layer4_outputs(3788)) or (layer4_outputs(2346)));
    layer5_outputs(4641) <= not(layer4_outputs(1594));
    layer5_outputs(4642) <= not(layer4_outputs(1889)) or (layer4_outputs(1070));
    layer5_outputs(4643) <= not(layer4_outputs(1148));
    layer5_outputs(4644) <= not(layer4_outputs(4000));
    layer5_outputs(4645) <= (layer4_outputs(1238)) and not (layer4_outputs(4530));
    layer5_outputs(4646) <= not((layer4_outputs(3786)) xor (layer4_outputs(1829)));
    layer5_outputs(4647) <= not(layer4_outputs(4640));
    layer5_outputs(4648) <= (layer4_outputs(4536)) and not (layer4_outputs(4033));
    layer5_outputs(4649) <= not(layer4_outputs(4970)) or (layer4_outputs(3475));
    layer5_outputs(4650) <= (layer4_outputs(1591)) and not (layer4_outputs(2760));
    layer5_outputs(4651) <= layer4_outputs(2887);
    layer5_outputs(4652) <= not((layer4_outputs(3259)) xor (layer4_outputs(209)));
    layer5_outputs(4653) <= layer4_outputs(753);
    layer5_outputs(4654) <= not(layer4_outputs(1962));
    layer5_outputs(4655) <= (layer4_outputs(3119)) xor (layer4_outputs(2938));
    layer5_outputs(4656) <= not(layer4_outputs(572)) or (layer4_outputs(4003));
    layer5_outputs(4657) <= not(layer4_outputs(5118)) or (layer4_outputs(2120));
    layer5_outputs(4658) <= layer4_outputs(1635);
    layer5_outputs(4659) <= (layer4_outputs(4983)) or (layer4_outputs(3060));
    layer5_outputs(4660) <= not((layer4_outputs(747)) and (layer4_outputs(3008)));
    layer5_outputs(4661) <= not(layer4_outputs(4887)) or (layer4_outputs(688));
    layer5_outputs(4662) <= (layer4_outputs(3361)) and not (layer4_outputs(691));
    layer5_outputs(4663) <= not(layer4_outputs(136));
    layer5_outputs(4664) <= layer4_outputs(1899);
    layer5_outputs(4665) <= '1';
    layer5_outputs(4666) <= layer4_outputs(1179);
    layer5_outputs(4667) <= not(layer4_outputs(306));
    layer5_outputs(4668) <= not((layer4_outputs(2401)) or (layer4_outputs(2158)));
    layer5_outputs(4669) <= layer4_outputs(174);
    layer5_outputs(4670) <= layer4_outputs(2685);
    layer5_outputs(4671) <= not(layer4_outputs(2575));
    layer5_outputs(4672) <= (layer4_outputs(2791)) and not (layer4_outputs(480));
    layer5_outputs(4673) <= layer4_outputs(1811);
    layer5_outputs(4674) <= layer4_outputs(900);
    layer5_outputs(4675) <= not(layer4_outputs(2622));
    layer5_outputs(4676) <= (layer4_outputs(4123)) xor (layer4_outputs(2129));
    layer5_outputs(4677) <= (layer4_outputs(1400)) and not (layer4_outputs(1991));
    layer5_outputs(4678) <= not((layer4_outputs(4365)) or (layer4_outputs(479)));
    layer5_outputs(4679) <= layer4_outputs(1210);
    layer5_outputs(4680) <= layer4_outputs(1162);
    layer5_outputs(4681) <= layer4_outputs(971);
    layer5_outputs(4682) <= layer4_outputs(2364);
    layer5_outputs(4683) <= not(layer4_outputs(1188));
    layer5_outputs(4684) <= not(layer4_outputs(1841));
    layer5_outputs(4685) <= (layer4_outputs(4900)) and not (layer4_outputs(2597));
    layer5_outputs(4686) <= not(layer4_outputs(27));
    layer5_outputs(4687) <= not(layer4_outputs(5111));
    layer5_outputs(4688) <= not(layer4_outputs(2881));
    layer5_outputs(4689) <= not((layer4_outputs(3062)) or (layer4_outputs(1861)));
    layer5_outputs(4690) <= layer4_outputs(431);
    layer5_outputs(4691) <= not(layer4_outputs(1796)) or (layer4_outputs(3784));
    layer5_outputs(4692) <= (layer4_outputs(2810)) and not (layer4_outputs(528));
    layer5_outputs(4693) <= not(layer4_outputs(4118));
    layer5_outputs(4694) <= (layer4_outputs(238)) xor (layer4_outputs(495));
    layer5_outputs(4695) <= not(layer4_outputs(39)) or (layer4_outputs(172));
    layer5_outputs(4696) <= not(layer4_outputs(2066)) or (layer4_outputs(3552));
    layer5_outputs(4697) <= layer4_outputs(1400);
    layer5_outputs(4698) <= not(layer4_outputs(5036)) or (layer4_outputs(2859));
    layer5_outputs(4699) <= not(layer4_outputs(1427));
    layer5_outputs(4700) <= not(layer4_outputs(548));
    layer5_outputs(4701) <= (layer4_outputs(45)) and (layer4_outputs(2764));
    layer5_outputs(4702) <= layer4_outputs(4744);
    layer5_outputs(4703) <= not(layer4_outputs(119)) or (layer4_outputs(1997));
    layer5_outputs(4704) <= '0';
    layer5_outputs(4705) <= not((layer4_outputs(3017)) xor (layer4_outputs(1907)));
    layer5_outputs(4706) <= '0';
    layer5_outputs(4707) <= '1';
    layer5_outputs(4708) <= (layer4_outputs(4010)) and not (layer4_outputs(3837));
    layer5_outputs(4709) <= (layer4_outputs(4304)) and not (layer4_outputs(0));
    layer5_outputs(4710) <= '0';
    layer5_outputs(4711) <= not(layer4_outputs(1193));
    layer5_outputs(4712) <= not(layer4_outputs(446)) or (layer4_outputs(1112));
    layer5_outputs(4713) <= layer4_outputs(2358);
    layer5_outputs(4714) <= not(layer4_outputs(3590));
    layer5_outputs(4715) <= layer4_outputs(4591);
    layer5_outputs(4716) <= (layer4_outputs(399)) and not (layer4_outputs(1444));
    layer5_outputs(4717) <= (layer4_outputs(4266)) and not (layer4_outputs(3265));
    layer5_outputs(4718) <= not((layer4_outputs(2708)) and (layer4_outputs(2270)));
    layer5_outputs(4719) <= not(layer4_outputs(4451));
    layer5_outputs(4720) <= not(layer4_outputs(3856)) or (layer4_outputs(1304));
    layer5_outputs(4721) <= (layer4_outputs(2631)) or (layer4_outputs(3001));
    layer5_outputs(4722) <= not(layer4_outputs(3958)) or (layer4_outputs(4960));
    layer5_outputs(4723) <= not(layer4_outputs(2784));
    layer5_outputs(4724) <= layer4_outputs(4720);
    layer5_outputs(4725) <= not(layer4_outputs(3972));
    layer5_outputs(4726) <= not(layer4_outputs(4017));
    layer5_outputs(4727) <= layer4_outputs(2669);
    layer5_outputs(4728) <= (layer4_outputs(470)) and (layer4_outputs(1265));
    layer5_outputs(4729) <= not(layer4_outputs(4284)) or (layer4_outputs(957));
    layer5_outputs(4730) <= not(layer4_outputs(3247));
    layer5_outputs(4731) <= not(layer4_outputs(3447));
    layer5_outputs(4732) <= layer4_outputs(1112);
    layer5_outputs(4733) <= layer4_outputs(2209);
    layer5_outputs(4734) <= (layer4_outputs(972)) or (layer4_outputs(4277));
    layer5_outputs(4735) <= (layer4_outputs(3671)) and not (layer4_outputs(4540));
    layer5_outputs(4736) <= (layer4_outputs(4632)) or (layer4_outputs(3012));
    layer5_outputs(4737) <= not(layer4_outputs(647));
    layer5_outputs(4738) <= '1';
    layer5_outputs(4739) <= not(layer4_outputs(4347));
    layer5_outputs(4740) <= not(layer4_outputs(15));
    layer5_outputs(4741) <= (layer4_outputs(2709)) and (layer4_outputs(1778));
    layer5_outputs(4742) <= (layer4_outputs(2351)) and not (layer4_outputs(3550));
    layer5_outputs(4743) <= layer4_outputs(1448);
    layer5_outputs(4744) <= layer4_outputs(587);
    layer5_outputs(4745) <= (layer4_outputs(3358)) and not (layer4_outputs(3862));
    layer5_outputs(4746) <= not((layer4_outputs(3542)) xor (layer4_outputs(3916)));
    layer5_outputs(4747) <= layer4_outputs(3513);
    layer5_outputs(4748) <= not(layer4_outputs(3240));
    layer5_outputs(4749) <= layer4_outputs(349);
    layer5_outputs(4750) <= layer4_outputs(1589);
    layer5_outputs(4751) <= layer4_outputs(309);
    layer5_outputs(4752) <= not((layer4_outputs(4245)) or (layer4_outputs(2706)));
    layer5_outputs(4753) <= layer4_outputs(1026);
    layer5_outputs(4754) <= not(layer4_outputs(4803));
    layer5_outputs(4755) <= '1';
    layer5_outputs(4756) <= layer4_outputs(170);
    layer5_outputs(4757) <= (layer4_outputs(3156)) xor (layer4_outputs(2117));
    layer5_outputs(4758) <= layer4_outputs(1105);
    layer5_outputs(4759) <= layer4_outputs(4567);
    layer5_outputs(4760) <= (layer4_outputs(1637)) and (layer4_outputs(3068));
    layer5_outputs(4761) <= not(layer4_outputs(1560)) or (layer4_outputs(3460));
    layer5_outputs(4762) <= not(layer4_outputs(1517));
    layer5_outputs(4763) <= not(layer4_outputs(1260));
    layer5_outputs(4764) <= layer4_outputs(2131);
    layer5_outputs(4765) <= '0';
    layer5_outputs(4766) <= (layer4_outputs(3607)) and not (layer4_outputs(3837));
    layer5_outputs(4767) <= layer4_outputs(3645);
    layer5_outputs(4768) <= not(layer4_outputs(1320)) or (layer4_outputs(2204));
    layer5_outputs(4769) <= (layer4_outputs(5014)) and not (layer4_outputs(2011));
    layer5_outputs(4770) <= not(layer4_outputs(2980)) or (layer4_outputs(3825));
    layer5_outputs(4771) <= not((layer4_outputs(2216)) and (layer4_outputs(1565)));
    layer5_outputs(4772) <= '0';
    layer5_outputs(4773) <= not((layer4_outputs(3019)) xor (layer4_outputs(4896)));
    layer5_outputs(4774) <= not((layer4_outputs(2100)) or (layer4_outputs(3298)));
    layer5_outputs(4775) <= (layer4_outputs(2388)) and (layer4_outputs(2019));
    layer5_outputs(4776) <= not((layer4_outputs(2827)) or (layer4_outputs(1078)));
    layer5_outputs(4777) <= not(layer4_outputs(1935));
    layer5_outputs(4778) <= not(layer4_outputs(3675)) or (layer4_outputs(4985));
    layer5_outputs(4779) <= layer4_outputs(3365);
    layer5_outputs(4780) <= not(layer4_outputs(2327));
    layer5_outputs(4781) <= (layer4_outputs(2875)) and not (layer4_outputs(4089));
    layer5_outputs(4782) <= not(layer4_outputs(1113)) or (layer4_outputs(1476));
    layer5_outputs(4783) <= '1';
    layer5_outputs(4784) <= layer4_outputs(2426);
    layer5_outputs(4785) <= (layer4_outputs(1740)) and not (layer4_outputs(4303));
    layer5_outputs(4786) <= '0';
    layer5_outputs(4787) <= not(layer4_outputs(3546));
    layer5_outputs(4788) <= (layer4_outputs(3953)) xor (layer4_outputs(4842));
    layer5_outputs(4789) <= layer4_outputs(1137);
    layer5_outputs(4790) <= not(layer4_outputs(3885));
    layer5_outputs(4791) <= layer4_outputs(2468);
    layer5_outputs(4792) <= not(layer4_outputs(775)) or (layer4_outputs(4718));
    layer5_outputs(4793) <= (layer4_outputs(1353)) and not (layer4_outputs(491));
    layer5_outputs(4794) <= layer4_outputs(1302);
    layer5_outputs(4795) <= not((layer4_outputs(2810)) xor (layer4_outputs(4711)));
    layer5_outputs(4796) <= layer4_outputs(3232);
    layer5_outputs(4797) <= not((layer4_outputs(965)) or (layer4_outputs(190)));
    layer5_outputs(4798) <= not(layer4_outputs(130));
    layer5_outputs(4799) <= not(layer4_outputs(682));
    layer5_outputs(4800) <= layer4_outputs(3173);
    layer5_outputs(4801) <= not((layer4_outputs(1263)) and (layer4_outputs(4699)));
    layer5_outputs(4802) <= (layer4_outputs(2995)) and not (layer4_outputs(2542));
    layer5_outputs(4803) <= not(layer4_outputs(3116));
    layer5_outputs(4804) <= (layer4_outputs(4628)) and not (layer4_outputs(4769));
    layer5_outputs(4805) <= '0';
    layer5_outputs(4806) <= not((layer4_outputs(2557)) xor (layer4_outputs(4141)));
    layer5_outputs(4807) <= layer4_outputs(851);
    layer5_outputs(4808) <= layer4_outputs(3780);
    layer5_outputs(4809) <= not(layer4_outputs(3537)) or (layer4_outputs(3151));
    layer5_outputs(4810) <= (layer4_outputs(3246)) xor (layer4_outputs(1944));
    layer5_outputs(4811) <= not(layer4_outputs(4019));
    layer5_outputs(4812) <= not(layer4_outputs(4161));
    layer5_outputs(4813) <= not(layer4_outputs(3609)) or (layer4_outputs(1375));
    layer5_outputs(4814) <= (layer4_outputs(3457)) xor (layer4_outputs(3943));
    layer5_outputs(4815) <= not(layer4_outputs(5052));
    layer5_outputs(4816) <= not(layer4_outputs(1915));
    layer5_outputs(4817) <= (layer4_outputs(434)) xor (layer4_outputs(2877));
    layer5_outputs(4818) <= '0';
    layer5_outputs(4819) <= (layer4_outputs(4202)) xor (layer4_outputs(5096));
    layer5_outputs(4820) <= '1';
    layer5_outputs(4821) <= layer4_outputs(1148);
    layer5_outputs(4822) <= not(layer4_outputs(331));
    layer5_outputs(4823) <= not(layer4_outputs(4916));
    layer5_outputs(4824) <= not(layer4_outputs(2530));
    layer5_outputs(4825) <= layer4_outputs(2531);
    layer5_outputs(4826) <= layer4_outputs(3405);
    layer5_outputs(4827) <= (layer4_outputs(610)) and (layer4_outputs(1375));
    layer5_outputs(4828) <= not(layer4_outputs(1719));
    layer5_outputs(4829) <= not(layer4_outputs(773));
    layer5_outputs(4830) <= not(layer4_outputs(2027));
    layer5_outputs(4831) <= layer4_outputs(861);
    layer5_outputs(4832) <= (layer4_outputs(4972)) and not (layer4_outputs(3991));
    layer5_outputs(4833) <= (layer4_outputs(1847)) or (layer4_outputs(4967));
    layer5_outputs(4834) <= not(layer4_outputs(549));
    layer5_outputs(4835) <= not(layer4_outputs(3077));
    layer5_outputs(4836) <= (layer4_outputs(732)) and not (layer4_outputs(737));
    layer5_outputs(4837) <= '1';
    layer5_outputs(4838) <= layer4_outputs(707);
    layer5_outputs(4839) <= not((layer4_outputs(2094)) xor (layer4_outputs(2308)));
    layer5_outputs(4840) <= '1';
    layer5_outputs(4841) <= layer4_outputs(3267);
    layer5_outputs(4842) <= not((layer4_outputs(2168)) and (layer4_outputs(992)));
    layer5_outputs(4843) <= not(layer4_outputs(4704)) or (layer4_outputs(2525));
    layer5_outputs(4844) <= (layer4_outputs(402)) xor (layer4_outputs(2177));
    layer5_outputs(4845) <= (layer4_outputs(1359)) and not (layer4_outputs(1082));
    layer5_outputs(4846) <= not(layer4_outputs(4340)) or (layer4_outputs(1288));
    layer5_outputs(4847) <= layer4_outputs(1290);
    layer5_outputs(4848) <= not(layer4_outputs(780));
    layer5_outputs(4849) <= not(layer4_outputs(3801));
    layer5_outputs(4850) <= (layer4_outputs(483)) xor (layer4_outputs(3126));
    layer5_outputs(4851) <= layer4_outputs(4652);
    layer5_outputs(4852) <= not(layer4_outputs(551));
    layer5_outputs(4853) <= not(layer4_outputs(1273)) or (layer4_outputs(5105));
    layer5_outputs(4854) <= not(layer4_outputs(4020));
    layer5_outputs(4855) <= not((layer4_outputs(1579)) and (layer4_outputs(1777)));
    layer5_outputs(4856) <= not(layer4_outputs(4660));
    layer5_outputs(4857) <= (layer4_outputs(4989)) and (layer4_outputs(4314));
    layer5_outputs(4858) <= (layer4_outputs(4244)) or (layer4_outputs(3306));
    layer5_outputs(4859) <= not(layer4_outputs(3811)) or (layer4_outputs(2608));
    layer5_outputs(4860) <= layer4_outputs(1635);
    layer5_outputs(4861) <= not(layer4_outputs(790));
    layer5_outputs(4862) <= not(layer4_outputs(4669));
    layer5_outputs(4863) <= (layer4_outputs(4071)) and not (layer4_outputs(4775));
    layer5_outputs(4864) <= not((layer4_outputs(2804)) xor (layer4_outputs(2452)));
    layer5_outputs(4865) <= (layer4_outputs(4153)) or (layer4_outputs(3223));
    layer5_outputs(4866) <= not(layer4_outputs(2653)) or (layer4_outputs(3013));
    layer5_outputs(4867) <= (layer4_outputs(2784)) or (layer4_outputs(4182));
    layer5_outputs(4868) <= not((layer4_outputs(2043)) xor (layer4_outputs(3549)));
    layer5_outputs(4869) <= not((layer4_outputs(1219)) and (layer4_outputs(2310)));
    layer5_outputs(4870) <= not((layer4_outputs(3670)) xor (layer4_outputs(13)));
    layer5_outputs(4871) <= not(layer4_outputs(4357));
    layer5_outputs(4872) <= layer4_outputs(2006);
    layer5_outputs(4873) <= (layer4_outputs(1267)) and not (layer4_outputs(376));
    layer5_outputs(4874) <= (layer4_outputs(4044)) or (layer4_outputs(4914));
    layer5_outputs(4875) <= not(layer4_outputs(2813));
    layer5_outputs(4876) <= '1';
    layer5_outputs(4877) <= (layer4_outputs(562)) xor (layer4_outputs(810));
    layer5_outputs(4878) <= not((layer4_outputs(367)) and (layer4_outputs(4329)));
    layer5_outputs(4879) <= layer4_outputs(3621);
    layer5_outputs(4880) <= layer4_outputs(1920);
    layer5_outputs(4881) <= not(layer4_outputs(3809));
    layer5_outputs(4882) <= layer4_outputs(4606);
    layer5_outputs(4883) <= (layer4_outputs(568)) and not (layer4_outputs(4698));
    layer5_outputs(4884) <= layer4_outputs(2896);
    layer5_outputs(4885) <= not((layer4_outputs(2569)) xor (layer4_outputs(3732)));
    layer5_outputs(4886) <= not(layer4_outputs(4208));
    layer5_outputs(4887) <= layer4_outputs(26);
    layer5_outputs(4888) <= not(layer4_outputs(4154));
    layer5_outputs(4889) <= (layer4_outputs(2891)) and not (layer4_outputs(2721));
    layer5_outputs(4890) <= not(layer4_outputs(1350));
    layer5_outputs(4891) <= (layer4_outputs(4564)) and (layer4_outputs(4312));
    layer5_outputs(4892) <= not((layer4_outputs(3859)) or (layer4_outputs(3080)));
    layer5_outputs(4893) <= (layer4_outputs(2092)) and (layer4_outputs(3904));
    layer5_outputs(4894) <= not(layer4_outputs(994));
    layer5_outputs(4895) <= '1';
    layer5_outputs(4896) <= not(layer4_outputs(4710));
    layer5_outputs(4897) <= (layer4_outputs(3210)) and not (layer4_outputs(2555));
    layer5_outputs(4898) <= '0';
    layer5_outputs(4899) <= layer4_outputs(754);
    layer5_outputs(4900) <= not(layer4_outputs(4857)) or (layer4_outputs(1788));
    layer5_outputs(4901) <= (layer4_outputs(2742)) and (layer4_outputs(1806));
    layer5_outputs(4902) <= not(layer4_outputs(4172));
    layer5_outputs(4903) <= not(layer4_outputs(3972));
    layer5_outputs(4904) <= not(layer4_outputs(1855));
    layer5_outputs(4905) <= layer4_outputs(4410);
    layer5_outputs(4906) <= layer4_outputs(828);
    layer5_outputs(4907) <= not(layer4_outputs(2976));
    layer5_outputs(4908) <= layer4_outputs(2395);
    layer5_outputs(4909) <= layer4_outputs(526);
    layer5_outputs(4910) <= not(layer4_outputs(120));
    layer5_outputs(4911) <= not(layer4_outputs(2114)) or (layer4_outputs(604));
    layer5_outputs(4912) <= layer4_outputs(3018);
    layer5_outputs(4913) <= not((layer4_outputs(3986)) xor (layer4_outputs(25)));
    layer5_outputs(4914) <= not((layer4_outputs(2001)) or (layer4_outputs(125)));
    layer5_outputs(4915) <= layer4_outputs(3503);
    layer5_outputs(4916) <= not(layer4_outputs(3998));
    layer5_outputs(4917) <= (layer4_outputs(2072)) and (layer4_outputs(5086));
    layer5_outputs(4918) <= layer4_outputs(580);
    layer5_outputs(4919) <= not(layer4_outputs(3153));
    layer5_outputs(4920) <= not((layer4_outputs(3771)) and (layer4_outputs(4156)));
    layer5_outputs(4921) <= layer4_outputs(4772);
    layer5_outputs(4922) <= not(layer4_outputs(3636));
    layer5_outputs(4923) <= (layer4_outputs(477)) and (layer4_outputs(4604));
    layer5_outputs(4924) <= not(layer4_outputs(1249)) or (layer4_outputs(3195));
    layer5_outputs(4925) <= layer4_outputs(3519);
    layer5_outputs(4926) <= (layer4_outputs(468)) and (layer4_outputs(2086));
    layer5_outputs(4927) <= layer4_outputs(154);
    layer5_outputs(4928) <= not(layer4_outputs(2854));
    layer5_outputs(4929) <= not(layer4_outputs(4668));
    layer5_outputs(4930) <= not(layer4_outputs(4191));
    layer5_outputs(4931) <= layer4_outputs(3654);
    layer5_outputs(4932) <= layer4_outputs(4879);
    layer5_outputs(4933) <= not(layer4_outputs(2385));
    layer5_outputs(4934) <= layer4_outputs(1699);
    layer5_outputs(4935) <= not((layer4_outputs(3679)) or (layer4_outputs(627)));
    layer5_outputs(4936) <= not(layer4_outputs(5024));
    layer5_outputs(4937) <= not(layer4_outputs(2329)) or (layer4_outputs(4364));
    layer5_outputs(4938) <= not(layer4_outputs(5047)) or (layer4_outputs(2378));
    layer5_outputs(4939) <= (layer4_outputs(2027)) and (layer4_outputs(818));
    layer5_outputs(4940) <= layer4_outputs(2982);
    layer5_outputs(4941) <= not(layer4_outputs(3867));
    layer5_outputs(4942) <= (layer4_outputs(2962)) and not (layer4_outputs(2431));
    layer5_outputs(4943) <= not(layer4_outputs(2424));
    layer5_outputs(4944) <= not(layer4_outputs(1950));
    layer5_outputs(4945) <= (layer4_outputs(3729)) or (layer4_outputs(4301));
    layer5_outputs(4946) <= not(layer4_outputs(4081));
    layer5_outputs(4947) <= '1';
    layer5_outputs(4948) <= not((layer4_outputs(907)) or (layer4_outputs(728)));
    layer5_outputs(4949) <= (layer4_outputs(2982)) and not (layer4_outputs(814));
    layer5_outputs(4950) <= '0';
    layer5_outputs(4951) <= not(layer4_outputs(42));
    layer5_outputs(4952) <= layer4_outputs(3964);
    layer5_outputs(4953) <= layer4_outputs(2046);
    layer5_outputs(4954) <= not(layer4_outputs(4525));
    layer5_outputs(4955) <= (layer4_outputs(899)) and not (layer4_outputs(989));
    layer5_outputs(4956) <= not((layer4_outputs(3084)) or (layer4_outputs(83)));
    layer5_outputs(4957) <= layer4_outputs(4582);
    layer5_outputs(4958) <= not(layer4_outputs(928)) or (layer4_outputs(2570));
    layer5_outputs(4959) <= not(layer4_outputs(3184));
    layer5_outputs(4960) <= not(layer4_outputs(588));
    layer5_outputs(4961) <= (layer4_outputs(1782)) xor (layer4_outputs(1962));
    layer5_outputs(4962) <= not(layer4_outputs(3283));
    layer5_outputs(4963) <= layer4_outputs(547);
    layer5_outputs(4964) <= layer4_outputs(5085);
    layer5_outputs(4965) <= not(layer4_outputs(1933)) or (layer4_outputs(4142));
    layer5_outputs(4966) <= not(layer4_outputs(721));
    layer5_outputs(4967) <= not((layer4_outputs(3038)) or (layer4_outputs(902)));
    layer5_outputs(4968) <= (layer4_outputs(543)) and not (layer4_outputs(1027));
    layer5_outputs(4969) <= not((layer4_outputs(4407)) and (layer4_outputs(3643)));
    layer5_outputs(4970) <= not((layer4_outputs(1757)) xor (layer4_outputs(2975)));
    layer5_outputs(4971) <= '1';
    layer5_outputs(4972) <= not(layer4_outputs(798));
    layer5_outputs(4973) <= layer4_outputs(1268);
    layer5_outputs(4974) <= (layer4_outputs(547)) and (layer4_outputs(3229));
    layer5_outputs(4975) <= not(layer4_outputs(3707));
    layer5_outputs(4976) <= not((layer4_outputs(778)) xor (layer4_outputs(2441)));
    layer5_outputs(4977) <= layer4_outputs(2389);
    layer5_outputs(4978) <= not(layer4_outputs(4069)) or (layer4_outputs(4546));
    layer5_outputs(4979) <= not((layer4_outputs(4543)) and (layer4_outputs(4820)));
    layer5_outputs(4980) <= layer4_outputs(3831);
    layer5_outputs(4981) <= (layer4_outputs(521)) and not (layer4_outputs(803));
    layer5_outputs(4982) <= (layer4_outputs(3277)) and not (layer4_outputs(5075));
    layer5_outputs(4983) <= not(layer4_outputs(2635));
    layer5_outputs(4984) <= layer4_outputs(168);
    layer5_outputs(4985) <= layer4_outputs(4392);
    layer5_outputs(4986) <= layer4_outputs(1217);
    layer5_outputs(4987) <= not(layer4_outputs(2304));
    layer5_outputs(4988) <= (layer4_outputs(3984)) or (layer4_outputs(4662));
    layer5_outputs(4989) <= not(layer4_outputs(3709));
    layer5_outputs(4990) <= (layer4_outputs(4127)) and not (layer4_outputs(2819));
    layer5_outputs(4991) <= not(layer4_outputs(4427)) or (layer4_outputs(1276));
    layer5_outputs(4992) <= not((layer4_outputs(424)) or (layer4_outputs(3234)));
    layer5_outputs(4993) <= not((layer4_outputs(1730)) and (layer4_outputs(2690)));
    layer5_outputs(4994) <= not(layer4_outputs(4303));
    layer5_outputs(4995) <= not(layer4_outputs(893));
    layer5_outputs(4996) <= '1';
    layer5_outputs(4997) <= not(layer4_outputs(2627));
    layer5_outputs(4998) <= not((layer4_outputs(3919)) or (layer4_outputs(1168)));
    layer5_outputs(4999) <= not(layer4_outputs(1085)) or (layer4_outputs(217));
    layer5_outputs(5000) <= layer4_outputs(3608);
    layer5_outputs(5001) <= layer4_outputs(743);
    layer5_outputs(5002) <= layer4_outputs(4409);
    layer5_outputs(5003) <= (layer4_outputs(2849)) and (layer4_outputs(1872));
    layer5_outputs(5004) <= '0';
    layer5_outputs(5005) <= (layer4_outputs(2620)) and not (layer4_outputs(689));
    layer5_outputs(5006) <= (layer4_outputs(1202)) and not (layer4_outputs(1173));
    layer5_outputs(5007) <= (layer4_outputs(823)) or (layer4_outputs(2799));
    layer5_outputs(5008) <= layer4_outputs(4243);
    layer5_outputs(5009) <= not((layer4_outputs(401)) or (layer4_outputs(3839)));
    layer5_outputs(5010) <= not((layer4_outputs(2013)) or (layer4_outputs(445)));
    layer5_outputs(5011) <= layer4_outputs(2435);
    layer5_outputs(5012) <= layer4_outputs(1067);
    layer5_outputs(5013) <= (layer4_outputs(903)) and not (layer4_outputs(3360));
    layer5_outputs(5014) <= layer4_outputs(2004);
    layer5_outputs(5015) <= not(layer4_outputs(4537));
    layer5_outputs(5016) <= not(layer4_outputs(1024));
    layer5_outputs(5017) <= not(layer4_outputs(1106));
    layer5_outputs(5018) <= (layer4_outputs(4482)) and not (layer4_outputs(5010));
    layer5_outputs(5019) <= not(layer4_outputs(1614));
    layer5_outputs(5020) <= not(layer4_outputs(2160));
    layer5_outputs(5021) <= (layer4_outputs(1470)) or (layer4_outputs(2524));
    layer5_outputs(5022) <= (layer4_outputs(4989)) and not (layer4_outputs(3736));
    layer5_outputs(5023) <= '0';
    layer5_outputs(5024) <= not(layer4_outputs(393));
    layer5_outputs(5025) <= '1';
    layer5_outputs(5026) <= not(layer4_outputs(1786));
    layer5_outputs(5027) <= not(layer4_outputs(1473)) or (layer4_outputs(4987));
    layer5_outputs(5028) <= (layer4_outputs(3160)) xor (layer4_outputs(996));
    layer5_outputs(5029) <= not(layer4_outputs(628));
    layer5_outputs(5030) <= not(layer4_outputs(1302)) or (layer4_outputs(3582));
    layer5_outputs(5031) <= not((layer4_outputs(4878)) and (layer4_outputs(1853)));
    layer5_outputs(5032) <= not((layer4_outputs(1203)) or (layer4_outputs(4985)));
    layer5_outputs(5033) <= layer4_outputs(2309);
    layer5_outputs(5034) <= not(layer4_outputs(2149)) or (layer4_outputs(4710));
    layer5_outputs(5035) <= (layer4_outputs(3208)) xor (layer4_outputs(2759));
    layer5_outputs(5036) <= not(layer4_outputs(2642));
    layer5_outputs(5037) <= not(layer4_outputs(4860)) or (layer4_outputs(1469));
    layer5_outputs(5038) <= layer4_outputs(2877);
    layer5_outputs(5039) <= layer4_outputs(4439);
    layer5_outputs(5040) <= (layer4_outputs(3505)) and (layer4_outputs(3620));
    layer5_outputs(5041) <= (layer4_outputs(2861)) or (layer4_outputs(5103));
    layer5_outputs(5042) <= not(layer4_outputs(4525));
    layer5_outputs(5043) <= not(layer4_outputs(4673)) or (layer4_outputs(3998));
    layer5_outputs(5044) <= not((layer4_outputs(2909)) xor (layer4_outputs(2649)));
    layer5_outputs(5045) <= layer4_outputs(4227);
    layer5_outputs(5046) <= (layer4_outputs(402)) xor (layer4_outputs(4847));
    layer5_outputs(5047) <= not(layer4_outputs(2777));
    layer5_outputs(5048) <= not((layer4_outputs(1965)) or (layer4_outputs(1634)));
    layer5_outputs(5049) <= not(layer4_outputs(943));
    layer5_outputs(5050) <= (layer4_outputs(2931)) or (layer4_outputs(802));
    layer5_outputs(5051) <= not(layer4_outputs(1539));
    layer5_outputs(5052) <= not(layer4_outputs(3607)) or (layer4_outputs(3289));
    layer5_outputs(5053) <= not(layer4_outputs(9));
    layer5_outputs(5054) <= (layer4_outputs(4723)) and (layer4_outputs(4995));
    layer5_outputs(5055) <= layer4_outputs(4012);
    layer5_outputs(5056) <= not(layer4_outputs(1538)) or (layer4_outputs(440));
    layer5_outputs(5057) <= (layer4_outputs(4369)) and not (layer4_outputs(3849));
    layer5_outputs(5058) <= layer4_outputs(2392);
    layer5_outputs(5059) <= not(layer4_outputs(1004)) or (layer4_outputs(1744));
    layer5_outputs(5060) <= layer4_outputs(4601);
    layer5_outputs(5061) <= not((layer4_outputs(4066)) and (layer4_outputs(3747)));
    layer5_outputs(5062) <= not((layer4_outputs(2702)) or (layer4_outputs(4352)));
    layer5_outputs(5063) <= layer4_outputs(1939);
    layer5_outputs(5064) <= not(layer4_outputs(2184));
    layer5_outputs(5065) <= not(layer4_outputs(1102));
    layer5_outputs(5066) <= layer4_outputs(1161);
    layer5_outputs(5067) <= not(layer4_outputs(742)) or (layer4_outputs(1368));
    layer5_outputs(5068) <= (layer4_outputs(1199)) and not (layer4_outputs(3855));
    layer5_outputs(5069) <= not((layer4_outputs(2774)) or (layer4_outputs(3711)));
    layer5_outputs(5070) <= not((layer4_outputs(4515)) or (layer4_outputs(2381)));
    layer5_outputs(5071) <= not(layer4_outputs(1451));
    layer5_outputs(5072) <= (layer4_outputs(4522)) or (layer4_outputs(3192));
    layer5_outputs(5073) <= not((layer4_outputs(1585)) xor (layer4_outputs(4722)));
    layer5_outputs(5074) <= not((layer4_outputs(4701)) or (layer4_outputs(4128)));
    layer5_outputs(5075) <= not((layer4_outputs(1799)) and (layer4_outputs(2808)));
    layer5_outputs(5076) <= not((layer4_outputs(4291)) or (layer4_outputs(4982)));
    layer5_outputs(5077) <= layer4_outputs(1673);
    layer5_outputs(5078) <= not(layer4_outputs(557)) or (layer4_outputs(4844));
    layer5_outputs(5079) <= (layer4_outputs(3496)) and (layer4_outputs(3013));
    layer5_outputs(5080) <= not(layer4_outputs(1452));
    layer5_outputs(5081) <= (layer4_outputs(2937)) or (layer4_outputs(1104));
    layer5_outputs(5082) <= layer4_outputs(2562);
    layer5_outputs(5083) <= layer4_outputs(4993);
    layer5_outputs(5084) <= (layer4_outputs(865)) or (layer4_outputs(2062));
    layer5_outputs(5085) <= '1';
    layer5_outputs(5086) <= (layer4_outputs(3203)) and not (layer4_outputs(1074));
    layer5_outputs(5087) <= not((layer4_outputs(3533)) and (layer4_outputs(1513)));
    layer5_outputs(5088) <= not((layer4_outputs(4311)) xor (layer4_outputs(880)));
    layer5_outputs(5089) <= (layer4_outputs(451)) or (layer4_outputs(667));
    layer5_outputs(5090) <= not((layer4_outputs(968)) xor (layer4_outputs(1897)));
    layer5_outputs(5091) <= layer4_outputs(4076);
    layer5_outputs(5092) <= not((layer4_outputs(4314)) xor (layer4_outputs(4674)));
    layer5_outputs(5093) <= not(layer4_outputs(4673));
    layer5_outputs(5094) <= layer4_outputs(226);
    layer5_outputs(5095) <= layer4_outputs(3240);
    layer5_outputs(5096) <= not(layer4_outputs(5003));
    layer5_outputs(5097) <= layer4_outputs(695);
    layer5_outputs(5098) <= not(layer4_outputs(1088));
    layer5_outputs(5099) <= (layer4_outputs(5042)) or (layer4_outputs(1279));
    layer5_outputs(5100) <= not((layer4_outputs(2529)) and (layer4_outputs(3589)));
    layer5_outputs(5101) <= not(layer4_outputs(2391));
    layer5_outputs(5102) <= not(layer4_outputs(2763)) or (layer4_outputs(4841));
    layer5_outputs(5103) <= '1';
    layer5_outputs(5104) <= layer4_outputs(4923);
    layer5_outputs(5105) <= not((layer4_outputs(2726)) or (layer4_outputs(2752)));
    layer5_outputs(5106) <= not(layer4_outputs(4437));
    layer5_outputs(5107) <= not((layer4_outputs(1958)) and (layer4_outputs(578)));
    layer5_outputs(5108) <= layer4_outputs(4011);
    layer5_outputs(5109) <= not((layer4_outputs(4130)) xor (layer4_outputs(1886)));
    layer5_outputs(5110) <= (layer4_outputs(1115)) and not (layer4_outputs(4029));
    layer5_outputs(5111) <= (layer4_outputs(4727)) and not (layer4_outputs(4311));
    layer5_outputs(5112) <= not((layer4_outputs(409)) or (layer4_outputs(3499)));
    layer5_outputs(5113) <= (layer4_outputs(3107)) or (layer4_outputs(4957));
    layer5_outputs(5114) <= (layer4_outputs(2969)) xor (layer4_outputs(2801));
    layer5_outputs(5115) <= (layer4_outputs(4921)) or (layer4_outputs(4446));
    layer5_outputs(5116) <= not((layer4_outputs(405)) or (layer4_outputs(4766)));
    layer5_outputs(5117) <= layer4_outputs(3159);
    layer5_outputs(5118) <= not(layer4_outputs(4131));
    layer5_outputs(5119) <= not(layer4_outputs(424));
    layer6_outputs(0) <= (layer5_outputs(4942)) and not (layer5_outputs(1152));
    layer6_outputs(1) <= (layer5_outputs(3799)) and (layer5_outputs(1481));
    layer6_outputs(2) <= layer5_outputs(3218);
    layer6_outputs(3) <= not(layer5_outputs(2804));
    layer6_outputs(4) <= not(layer5_outputs(624));
    layer6_outputs(5) <= not(layer5_outputs(1447)) or (layer5_outputs(1009));
    layer6_outputs(6) <= (layer5_outputs(4815)) and not (layer5_outputs(219));
    layer6_outputs(7) <= layer5_outputs(2372);
    layer6_outputs(8) <= layer5_outputs(1192);
    layer6_outputs(9) <= layer5_outputs(4821);
    layer6_outputs(10) <= layer5_outputs(983);
    layer6_outputs(11) <= (layer5_outputs(1276)) xor (layer5_outputs(793));
    layer6_outputs(12) <= not(layer5_outputs(4420));
    layer6_outputs(13) <= layer5_outputs(3618);
    layer6_outputs(14) <= layer5_outputs(3047);
    layer6_outputs(15) <= not(layer5_outputs(2540));
    layer6_outputs(16) <= not((layer5_outputs(2456)) xor (layer5_outputs(1344)));
    layer6_outputs(17) <= not((layer5_outputs(2829)) and (layer5_outputs(4992)));
    layer6_outputs(18) <= layer5_outputs(859);
    layer6_outputs(19) <= (layer5_outputs(3837)) or (layer5_outputs(4480));
    layer6_outputs(20) <= not(layer5_outputs(5014));
    layer6_outputs(21) <= '0';
    layer6_outputs(22) <= not(layer5_outputs(3187));
    layer6_outputs(23) <= not(layer5_outputs(3458));
    layer6_outputs(24) <= not(layer5_outputs(466));
    layer6_outputs(25) <= layer5_outputs(3165);
    layer6_outputs(26) <= (layer5_outputs(2852)) and (layer5_outputs(87));
    layer6_outputs(27) <= layer5_outputs(3974);
    layer6_outputs(28) <= not(layer5_outputs(1457)) or (layer5_outputs(4185));
    layer6_outputs(29) <= not(layer5_outputs(4752));
    layer6_outputs(30) <= not(layer5_outputs(3722));
    layer6_outputs(31) <= not(layer5_outputs(1818));
    layer6_outputs(32) <= layer5_outputs(3679);
    layer6_outputs(33) <= layer5_outputs(1247);
    layer6_outputs(34) <= not(layer5_outputs(1642));
    layer6_outputs(35) <= not((layer5_outputs(2470)) xor (layer5_outputs(4970)));
    layer6_outputs(36) <= not(layer5_outputs(3547));
    layer6_outputs(37) <= (layer5_outputs(575)) xor (layer5_outputs(242));
    layer6_outputs(38) <= (layer5_outputs(1412)) and not (layer5_outputs(5048));
    layer6_outputs(39) <= not((layer5_outputs(2292)) or (layer5_outputs(3291)));
    layer6_outputs(40) <= not(layer5_outputs(926));
    layer6_outputs(41) <= layer5_outputs(4466);
    layer6_outputs(42) <= layer5_outputs(4184);
    layer6_outputs(43) <= '0';
    layer6_outputs(44) <= not(layer5_outputs(3891));
    layer6_outputs(45) <= layer5_outputs(194);
    layer6_outputs(46) <= (layer5_outputs(4738)) xor (layer5_outputs(4330));
    layer6_outputs(47) <= not(layer5_outputs(3303));
    layer6_outputs(48) <= layer5_outputs(42);
    layer6_outputs(49) <= not(layer5_outputs(3041));
    layer6_outputs(50) <= not((layer5_outputs(3968)) xor (layer5_outputs(4885)));
    layer6_outputs(51) <= not(layer5_outputs(4880));
    layer6_outputs(52) <= not((layer5_outputs(2369)) and (layer5_outputs(407)));
    layer6_outputs(53) <= (layer5_outputs(3755)) xor (layer5_outputs(2241));
    layer6_outputs(54) <= layer5_outputs(3247);
    layer6_outputs(55) <= not(layer5_outputs(1013)) or (layer5_outputs(3772));
    layer6_outputs(56) <= not((layer5_outputs(1496)) or (layer5_outputs(722)));
    layer6_outputs(57) <= not(layer5_outputs(3930));
    layer6_outputs(58) <= not(layer5_outputs(4111));
    layer6_outputs(59) <= layer5_outputs(4812);
    layer6_outputs(60) <= layer5_outputs(4703);
    layer6_outputs(61) <= layer5_outputs(1494);
    layer6_outputs(62) <= (layer5_outputs(1589)) and (layer5_outputs(1397));
    layer6_outputs(63) <= not(layer5_outputs(506)) or (layer5_outputs(1164));
    layer6_outputs(64) <= not(layer5_outputs(2637));
    layer6_outputs(65) <= layer5_outputs(732);
    layer6_outputs(66) <= (layer5_outputs(2111)) and not (layer5_outputs(342));
    layer6_outputs(67) <= not((layer5_outputs(1439)) and (layer5_outputs(3422)));
    layer6_outputs(68) <= '0';
    layer6_outputs(69) <= not((layer5_outputs(1220)) xor (layer5_outputs(4973)));
    layer6_outputs(70) <= (layer5_outputs(4396)) and (layer5_outputs(1094));
    layer6_outputs(71) <= not((layer5_outputs(1629)) xor (layer5_outputs(1492)));
    layer6_outputs(72) <= not(layer5_outputs(976));
    layer6_outputs(73) <= not(layer5_outputs(4394));
    layer6_outputs(74) <= not(layer5_outputs(3189));
    layer6_outputs(75) <= layer5_outputs(3565);
    layer6_outputs(76) <= not((layer5_outputs(1648)) xor (layer5_outputs(1616)));
    layer6_outputs(77) <= not(layer5_outputs(3252)) or (layer5_outputs(4178));
    layer6_outputs(78) <= not(layer5_outputs(3061));
    layer6_outputs(79) <= not(layer5_outputs(1203));
    layer6_outputs(80) <= layer5_outputs(1531);
    layer6_outputs(81) <= layer5_outputs(308);
    layer6_outputs(82) <= layer5_outputs(2866);
    layer6_outputs(83) <= not((layer5_outputs(4762)) or (layer5_outputs(1597)));
    layer6_outputs(84) <= not(layer5_outputs(2415));
    layer6_outputs(85) <= not((layer5_outputs(1687)) or (layer5_outputs(801)));
    layer6_outputs(86) <= layer5_outputs(1027);
    layer6_outputs(87) <= not(layer5_outputs(4486));
    layer6_outputs(88) <= not(layer5_outputs(4830));
    layer6_outputs(89) <= (layer5_outputs(1951)) xor (layer5_outputs(805));
    layer6_outputs(90) <= not(layer5_outputs(3269));
    layer6_outputs(91) <= not(layer5_outputs(4915));
    layer6_outputs(92) <= layer5_outputs(1566);
    layer6_outputs(93) <= layer5_outputs(1333);
    layer6_outputs(94) <= not(layer5_outputs(3414));
    layer6_outputs(95) <= '1';
    layer6_outputs(96) <= not(layer5_outputs(2644));
    layer6_outputs(97) <= layer5_outputs(4077);
    layer6_outputs(98) <= not((layer5_outputs(3340)) or (layer5_outputs(1609)));
    layer6_outputs(99) <= layer5_outputs(4524);
    layer6_outputs(100) <= layer5_outputs(3161);
    layer6_outputs(101) <= not(layer5_outputs(726));
    layer6_outputs(102) <= (layer5_outputs(1028)) or (layer5_outputs(1876));
    layer6_outputs(103) <= not(layer5_outputs(2643));
    layer6_outputs(104) <= layer5_outputs(4961);
    layer6_outputs(105) <= (layer5_outputs(3765)) or (layer5_outputs(1855));
    layer6_outputs(106) <= layer5_outputs(4623);
    layer6_outputs(107) <= not(layer5_outputs(732));
    layer6_outputs(108) <= not((layer5_outputs(837)) and (layer5_outputs(1278)));
    layer6_outputs(109) <= not((layer5_outputs(3356)) or (layer5_outputs(1612)));
    layer6_outputs(110) <= layer5_outputs(4329);
    layer6_outputs(111) <= (layer5_outputs(486)) and not (layer5_outputs(505));
    layer6_outputs(112) <= layer5_outputs(303);
    layer6_outputs(113) <= not((layer5_outputs(3575)) xor (layer5_outputs(798)));
    layer6_outputs(114) <= (layer5_outputs(2248)) and (layer5_outputs(4923));
    layer6_outputs(115) <= not(layer5_outputs(4872));
    layer6_outputs(116) <= (layer5_outputs(3808)) xor (layer5_outputs(1127));
    layer6_outputs(117) <= layer5_outputs(4730);
    layer6_outputs(118) <= not((layer5_outputs(1117)) and (layer5_outputs(1990)));
    layer6_outputs(119) <= layer5_outputs(2083);
    layer6_outputs(120) <= not((layer5_outputs(3593)) and (layer5_outputs(2644)));
    layer6_outputs(121) <= not(layer5_outputs(2565));
    layer6_outputs(122) <= (layer5_outputs(4725)) and not (layer5_outputs(5095));
    layer6_outputs(123) <= not(layer5_outputs(4169));
    layer6_outputs(124) <= (layer5_outputs(1585)) and not (layer5_outputs(2285));
    layer6_outputs(125) <= not(layer5_outputs(3595)) or (layer5_outputs(3029));
    layer6_outputs(126) <= not(layer5_outputs(1913));
    layer6_outputs(127) <= layer5_outputs(2230);
    layer6_outputs(128) <= not((layer5_outputs(2958)) xor (layer5_outputs(4364)));
    layer6_outputs(129) <= (layer5_outputs(3149)) and not (layer5_outputs(3546));
    layer6_outputs(130) <= not(layer5_outputs(2753));
    layer6_outputs(131) <= not((layer5_outputs(1115)) and (layer5_outputs(2886)));
    layer6_outputs(132) <= not((layer5_outputs(1432)) and (layer5_outputs(2738)));
    layer6_outputs(133) <= not(layer5_outputs(1780));
    layer6_outputs(134) <= (layer5_outputs(165)) and (layer5_outputs(2127));
    layer6_outputs(135) <= not(layer5_outputs(2550));
    layer6_outputs(136) <= layer5_outputs(4297);
    layer6_outputs(137) <= not(layer5_outputs(3773)) or (layer5_outputs(1958));
    layer6_outputs(138) <= not(layer5_outputs(4822));
    layer6_outputs(139) <= not(layer5_outputs(3911));
    layer6_outputs(140) <= (layer5_outputs(2501)) or (layer5_outputs(2144));
    layer6_outputs(141) <= layer5_outputs(398);
    layer6_outputs(142) <= (layer5_outputs(1478)) and not (layer5_outputs(1051));
    layer6_outputs(143) <= not(layer5_outputs(378));
    layer6_outputs(144) <= (layer5_outputs(1114)) and (layer5_outputs(3491));
    layer6_outputs(145) <= (layer5_outputs(1289)) and not (layer5_outputs(3923));
    layer6_outputs(146) <= (layer5_outputs(2776)) xor (layer5_outputs(324));
    layer6_outputs(147) <= (layer5_outputs(3009)) or (layer5_outputs(2745));
    layer6_outputs(148) <= not(layer5_outputs(2984));
    layer6_outputs(149) <= layer5_outputs(1197);
    layer6_outputs(150) <= not(layer5_outputs(4851));
    layer6_outputs(151) <= (layer5_outputs(82)) and not (layer5_outputs(1845));
    layer6_outputs(152) <= not(layer5_outputs(3024));
    layer6_outputs(153) <= (layer5_outputs(4426)) xor (layer5_outputs(2249));
    layer6_outputs(154) <= layer5_outputs(2020);
    layer6_outputs(155) <= not(layer5_outputs(3253));
    layer6_outputs(156) <= not(layer5_outputs(2294));
    layer6_outputs(157) <= layer5_outputs(189);
    layer6_outputs(158) <= not(layer5_outputs(5086)) or (layer5_outputs(4252));
    layer6_outputs(159) <= (layer5_outputs(1289)) xor (layer5_outputs(144));
    layer6_outputs(160) <= not(layer5_outputs(4624));
    layer6_outputs(161) <= (layer5_outputs(54)) and not (layer5_outputs(1296));
    layer6_outputs(162) <= (layer5_outputs(853)) xor (layer5_outputs(2642));
    layer6_outputs(163) <= not(layer5_outputs(2345));
    layer6_outputs(164) <= not(layer5_outputs(2457));
    layer6_outputs(165) <= not(layer5_outputs(886));
    layer6_outputs(166) <= (layer5_outputs(227)) and not (layer5_outputs(3102));
    layer6_outputs(167) <= layer5_outputs(4695);
    layer6_outputs(168) <= (layer5_outputs(3642)) xor (layer5_outputs(4427));
    layer6_outputs(169) <= not((layer5_outputs(4416)) and (layer5_outputs(4218)));
    layer6_outputs(170) <= layer5_outputs(5047);
    layer6_outputs(171) <= not((layer5_outputs(1377)) xor (layer5_outputs(752)));
    layer6_outputs(172) <= not(layer5_outputs(1562)) or (layer5_outputs(948));
    layer6_outputs(173) <= '1';
    layer6_outputs(174) <= layer5_outputs(3314);
    layer6_outputs(175) <= not(layer5_outputs(3183));
    layer6_outputs(176) <= not(layer5_outputs(88)) or (layer5_outputs(1803));
    layer6_outputs(177) <= not(layer5_outputs(4184));
    layer6_outputs(178) <= not(layer5_outputs(2246)) or (layer5_outputs(1724));
    layer6_outputs(179) <= layer5_outputs(1559);
    layer6_outputs(180) <= layer5_outputs(3474);
    layer6_outputs(181) <= not((layer5_outputs(643)) xor (layer5_outputs(2720)));
    layer6_outputs(182) <= layer5_outputs(3748);
    layer6_outputs(183) <= not(layer5_outputs(4629));
    layer6_outputs(184) <= (layer5_outputs(4806)) and not (layer5_outputs(211));
    layer6_outputs(185) <= not((layer5_outputs(3330)) and (layer5_outputs(423)));
    layer6_outputs(186) <= layer5_outputs(1314);
    layer6_outputs(187) <= layer5_outputs(4128);
    layer6_outputs(188) <= layer5_outputs(1687);
    layer6_outputs(189) <= layer5_outputs(312);
    layer6_outputs(190) <= not(layer5_outputs(3112));
    layer6_outputs(191) <= not(layer5_outputs(211));
    layer6_outputs(192) <= not((layer5_outputs(2160)) xor (layer5_outputs(411)));
    layer6_outputs(193) <= not(layer5_outputs(2126));
    layer6_outputs(194) <= not(layer5_outputs(4285));
    layer6_outputs(195) <= layer5_outputs(4240);
    layer6_outputs(196) <= not(layer5_outputs(4928));
    layer6_outputs(197) <= not(layer5_outputs(4123));
    layer6_outputs(198) <= not(layer5_outputs(232));
    layer6_outputs(199) <= layer5_outputs(1106);
    layer6_outputs(200) <= not(layer5_outputs(1488));
    layer6_outputs(201) <= (layer5_outputs(1588)) or (layer5_outputs(504));
    layer6_outputs(202) <= not(layer5_outputs(1665));
    layer6_outputs(203) <= not(layer5_outputs(2042));
    layer6_outputs(204) <= layer5_outputs(2571);
    layer6_outputs(205) <= (layer5_outputs(4406)) and not (layer5_outputs(2177));
    layer6_outputs(206) <= layer5_outputs(1836);
    layer6_outputs(207) <= (layer5_outputs(4713)) xor (layer5_outputs(1523));
    layer6_outputs(208) <= layer5_outputs(3346);
    layer6_outputs(209) <= (layer5_outputs(3255)) or (layer5_outputs(2618));
    layer6_outputs(210) <= (layer5_outputs(3056)) or (layer5_outputs(355));
    layer6_outputs(211) <= not(layer5_outputs(1693));
    layer6_outputs(212) <= layer5_outputs(1073);
    layer6_outputs(213) <= not(layer5_outputs(3475));
    layer6_outputs(214) <= not((layer5_outputs(4933)) xor (layer5_outputs(241)));
    layer6_outputs(215) <= layer5_outputs(2236);
    layer6_outputs(216) <= not(layer5_outputs(4875));
    layer6_outputs(217) <= layer5_outputs(4593);
    layer6_outputs(218) <= not(layer5_outputs(3347));
    layer6_outputs(219) <= not(layer5_outputs(4931));
    layer6_outputs(220) <= '1';
    layer6_outputs(221) <= not(layer5_outputs(3371));
    layer6_outputs(222) <= layer5_outputs(679);
    layer6_outputs(223) <= not(layer5_outputs(715));
    layer6_outputs(224) <= (layer5_outputs(4440)) xor (layer5_outputs(950));
    layer6_outputs(225) <= not(layer5_outputs(3274));
    layer6_outputs(226) <= not((layer5_outputs(2000)) xor (layer5_outputs(3326)));
    layer6_outputs(227) <= layer5_outputs(1226);
    layer6_outputs(228) <= layer5_outputs(3108);
    layer6_outputs(229) <= (layer5_outputs(782)) xor (layer5_outputs(250));
    layer6_outputs(230) <= not(layer5_outputs(4335)) or (layer5_outputs(5119));
    layer6_outputs(231) <= not((layer5_outputs(4070)) or (layer5_outputs(2987)));
    layer6_outputs(232) <= not(layer5_outputs(3031));
    layer6_outputs(233) <= not(layer5_outputs(3180));
    layer6_outputs(234) <= layer5_outputs(3767);
    layer6_outputs(235) <= not(layer5_outputs(2240));
    layer6_outputs(236) <= layer5_outputs(1828);
    layer6_outputs(237) <= (layer5_outputs(3056)) and (layer5_outputs(2952));
    layer6_outputs(238) <= layer5_outputs(3448);
    layer6_outputs(239) <= (layer5_outputs(1463)) xor (layer5_outputs(2327));
    layer6_outputs(240) <= not(layer5_outputs(4829));
    layer6_outputs(241) <= not(layer5_outputs(2742)) or (layer5_outputs(4849));
    layer6_outputs(242) <= not((layer5_outputs(4072)) and (layer5_outputs(3580)));
    layer6_outputs(243) <= not(layer5_outputs(1377));
    layer6_outputs(244) <= layer5_outputs(3179);
    layer6_outputs(245) <= not(layer5_outputs(3494));
    layer6_outputs(246) <= layer5_outputs(654);
    layer6_outputs(247) <= layer5_outputs(3313);
    layer6_outputs(248) <= not(layer5_outputs(4946));
    layer6_outputs(249) <= (layer5_outputs(2442)) xor (layer5_outputs(5025));
    layer6_outputs(250) <= not(layer5_outputs(4332));
    layer6_outputs(251) <= (layer5_outputs(1363)) and (layer5_outputs(4791));
    layer6_outputs(252) <= not((layer5_outputs(2638)) xor (layer5_outputs(4669)));
    layer6_outputs(253) <= not((layer5_outputs(2268)) or (layer5_outputs(3065)));
    layer6_outputs(254) <= layer5_outputs(1963);
    layer6_outputs(255) <= not(layer5_outputs(5063));
    layer6_outputs(256) <= not(layer5_outputs(3936));
    layer6_outputs(257) <= not(layer5_outputs(685));
    layer6_outputs(258) <= not(layer5_outputs(2601));
    layer6_outputs(259) <= not(layer5_outputs(966));
    layer6_outputs(260) <= not(layer5_outputs(397));
    layer6_outputs(261) <= not((layer5_outputs(59)) xor (layer5_outputs(2128)));
    layer6_outputs(262) <= (layer5_outputs(4741)) and not (layer5_outputs(42));
    layer6_outputs(263) <= layer5_outputs(2837);
    layer6_outputs(264) <= not((layer5_outputs(4643)) xor (layer5_outputs(2406)));
    layer6_outputs(265) <= not(layer5_outputs(874));
    layer6_outputs(266) <= not(layer5_outputs(4214)) or (layer5_outputs(3157));
    layer6_outputs(267) <= layer5_outputs(5077);
    layer6_outputs(268) <= not(layer5_outputs(4071));
    layer6_outputs(269) <= not(layer5_outputs(321));
    layer6_outputs(270) <= not(layer5_outputs(4420));
    layer6_outputs(271) <= (layer5_outputs(2681)) and not (layer5_outputs(2606));
    layer6_outputs(272) <= layer5_outputs(3496);
    layer6_outputs(273) <= layer5_outputs(3595);
    layer6_outputs(274) <= not(layer5_outputs(4155));
    layer6_outputs(275) <= (layer5_outputs(4038)) and not (layer5_outputs(3528));
    layer6_outputs(276) <= not(layer5_outputs(4172));
    layer6_outputs(277) <= not(layer5_outputs(1727));
    layer6_outputs(278) <= layer5_outputs(2867);
    layer6_outputs(279) <= not(layer5_outputs(2632));
    layer6_outputs(280) <= layer5_outputs(3831);
    layer6_outputs(281) <= (layer5_outputs(4479)) and not (layer5_outputs(4197));
    layer6_outputs(282) <= not(layer5_outputs(3427));
    layer6_outputs(283) <= layer5_outputs(2985);
    layer6_outputs(284) <= not(layer5_outputs(3168)) or (layer5_outputs(2843));
    layer6_outputs(285) <= (layer5_outputs(4012)) and (layer5_outputs(3215));
    layer6_outputs(286) <= layer5_outputs(1866);
    layer6_outputs(287) <= (layer5_outputs(2092)) xor (layer5_outputs(4963));
    layer6_outputs(288) <= layer5_outputs(3498);
    layer6_outputs(289) <= layer5_outputs(2490);
    layer6_outputs(290) <= not(layer5_outputs(4674));
    layer6_outputs(291) <= not((layer5_outputs(4711)) or (layer5_outputs(385)));
    layer6_outputs(292) <= layer5_outputs(1978);
    layer6_outputs(293) <= not(layer5_outputs(4108));
    layer6_outputs(294) <= (layer5_outputs(887)) and not (layer5_outputs(4544));
    layer6_outputs(295) <= layer5_outputs(2652);
    layer6_outputs(296) <= not((layer5_outputs(5058)) xor (layer5_outputs(4557)));
    layer6_outputs(297) <= not(layer5_outputs(2864));
    layer6_outputs(298) <= layer5_outputs(1713);
    layer6_outputs(299) <= not(layer5_outputs(2521));
    layer6_outputs(300) <= not(layer5_outputs(1753));
    layer6_outputs(301) <= layer5_outputs(187);
    layer6_outputs(302) <= not((layer5_outputs(1175)) xor (layer5_outputs(2509)));
    layer6_outputs(303) <= not(layer5_outputs(3279));
    layer6_outputs(304) <= (layer5_outputs(116)) xor (layer5_outputs(3733));
    layer6_outputs(305) <= not(layer5_outputs(2794));
    layer6_outputs(306) <= not(layer5_outputs(3665));
    layer6_outputs(307) <= (layer5_outputs(3054)) xor (layer5_outputs(3457));
    layer6_outputs(308) <= layer5_outputs(4038);
    layer6_outputs(309) <= not((layer5_outputs(653)) or (layer5_outputs(1406)));
    layer6_outputs(310) <= not((layer5_outputs(3125)) and (layer5_outputs(3718)));
    layer6_outputs(311) <= layer5_outputs(4070);
    layer6_outputs(312) <= layer5_outputs(2445);
    layer6_outputs(313) <= not(layer5_outputs(2143));
    layer6_outputs(314) <= not(layer5_outputs(2286));
    layer6_outputs(315) <= not(layer5_outputs(1211));
    layer6_outputs(316) <= (layer5_outputs(777)) and not (layer5_outputs(3620));
    layer6_outputs(317) <= layer5_outputs(130);
    layer6_outputs(318) <= layer5_outputs(708);
    layer6_outputs(319) <= layer5_outputs(2629);
    layer6_outputs(320) <= layer5_outputs(343);
    layer6_outputs(321) <= not((layer5_outputs(4075)) or (layer5_outputs(4796)));
    layer6_outputs(322) <= not(layer5_outputs(2670)) or (layer5_outputs(354));
    layer6_outputs(323) <= not((layer5_outputs(1597)) xor (layer5_outputs(3094)));
    layer6_outputs(324) <= not(layer5_outputs(2421)) or (layer5_outputs(1086));
    layer6_outputs(325) <= layer5_outputs(1816);
    layer6_outputs(326) <= layer5_outputs(4073);
    layer6_outputs(327) <= layer5_outputs(2819);
    layer6_outputs(328) <= not(layer5_outputs(3000));
    layer6_outputs(329) <= layer5_outputs(432);
    layer6_outputs(330) <= layer5_outputs(4652);
    layer6_outputs(331) <= layer5_outputs(3931);
    layer6_outputs(332) <= (layer5_outputs(4529)) and not (layer5_outputs(3073));
    layer6_outputs(333) <= (layer5_outputs(1180)) xor (layer5_outputs(5054));
    layer6_outputs(334) <= not(layer5_outputs(1290));
    layer6_outputs(335) <= layer5_outputs(230);
    layer6_outputs(336) <= not((layer5_outputs(2679)) or (layer5_outputs(2326)));
    layer6_outputs(337) <= layer5_outputs(3726);
    layer6_outputs(338) <= not((layer5_outputs(2399)) xor (layer5_outputs(3173)));
    layer6_outputs(339) <= '1';
    layer6_outputs(340) <= layer5_outputs(1331);
    layer6_outputs(341) <= not(layer5_outputs(1801));
    layer6_outputs(342) <= not(layer5_outputs(3814));
    layer6_outputs(343) <= layer5_outputs(33);
    layer6_outputs(344) <= layer5_outputs(2479);
    layer6_outputs(345) <= not((layer5_outputs(3440)) or (layer5_outputs(4784)));
    layer6_outputs(346) <= (layer5_outputs(1745)) xor (layer5_outputs(3922));
    layer6_outputs(347) <= (layer5_outputs(3179)) xor (layer5_outputs(3750));
    layer6_outputs(348) <= layer5_outputs(2784);
    layer6_outputs(349) <= (layer5_outputs(90)) xor (layer5_outputs(4036));
    layer6_outputs(350) <= layer5_outputs(4882);
    layer6_outputs(351) <= not(layer5_outputs(3611)) or (layer5_outputs(1942));
    layer6_outputs(352) <= not((layer5_outputs(1563)) and (layer5_outputs(132)));
    layer6_outputs(353) <= layer5_outputs(4016);
    layer6_outputs(354) <= layer5_outputs(5080);
    layer6_outputs(355) <= layer5_outputs(3907);
    layer6_outputs(356) <= (layer5_outputs(4637)) xor (layer5_outputs(4598));
    layer6_outputs(357) <= layer5_outputs(1989);
    layer6_outputs(358) <= not(layer5_outputs(4097)) or (layer5_outputs(1455));
    layer6_outputs(359) <= not(layer5_outputs(50));
    layer6_outputs(360) <= (layer5_outputs(173)) and not (layer5_outputs(345));
    layer6_outputs(361) <= layer5_outputs(4613);
    layer6_outputs(362) <= not(layer5_outputs(4571));
    layer6_outputs(363) <= not(layer5_outputs(3695)) or (layer5_outputs(4868));
    layer6_outputs(364) <= layer5_outputs(4442);
    layer6_outputs(365) <= (layer5_outputs(174)) xor (layer5_outputs(1400));
    layer6_outputs(366) <= layer5_outputs(4241);
    layer6_outputs(367) <= (layer5_outputs(1351)) and not (layer5_outputs(4688));
    layer6_outputs(368) <= layer5_outputs(1275);
    layer6_outputs(369) <= (layer5_outputs(2897)) xor (layer5_outputs(715));
    layer6_outputs(370) <= not(layer5_outputs(3965));
    layer6_outputs(371) <= not(layer5_outputs(4168));
    layer6_outputs(372) <= not((layer5_outputs(4576)) and (layer5_outputs(2046)));
    layer6_outputs(373) <= layer5_outputs(2127);
    layer6_outputs(374) <= not(layer5_outputs(5116));
    layer6_outputs(375) <= (layer5_outputs(557)) xor (layer5_outputs(4750));
    layer6_outputs(376) <= (layer5_outputs(1235)) and not (layer5_outputs(3318));
    layer6_outputs(377) <= layer5_outputs(2635);
    layer6_outputs(378) <= layer5_outputs(3646);
    layer6_outputs(379) <= not(layer5_outputs(3187));
    layer6_outputs(380) <= (layer5_outputs(2408)) and (layer5_outputs(2063));
    layer6_outputs(381) <= not(layer5_outputs(3745));
    layer6_outputs(382) <= layer5_outputs(4473);
    layer6_outputs(383) <= (layer5_outputs(4542)) and (layer5_outputs(2433));
    layer6_outputs(384) <= layer5_outputs(2658);
    layer6_outputs(385) <= not(layer5_outputs(2691)) or (layer5_outputs(2913));
    layer6_outputs(386) <= (layer5_outputs(3606)) xor (layer5_outputs(15));
    layer6_outputs(387) <= layer5_outputs(4207);
    layer6_outputs(388) <= (layer5_outputs(863)) and not (layer5_outputs(906));
    layer6_outputs(389) <= (layer5_outputs(417)) and (layer5_outputs(4452));
    layer6_outputs(390) <= layer5_outputs(54);
    layer6_outputs(391) <= not((layer5_outputs(1941)) or (layer5_outputs(2722)));
    layer6_outputs(392) <= (layer5_outputs(4902)) and (layer5_outputs(1918));
    layer6_outputs(393) <= not(layer5_outputs(3270));
    layer6_outputs(394) <= layer5_outputs(970);
    layer6_outputs(395) <= not(layer5_outputs(4766));
    layer6_outputs(396) <= not((layer5_outputs(2615)) xor (layer5_outputs(3144)));
    layer6_outputs(397) <= layer5_outputs(4147);
    layer6_outputs(398) <= (layer5_outputs(4386)) and not (layer5_outputs(1105));
    layer6_outputs(399) <= layer5_outputs(1308);
    layer6_outputs(400) <= (layer5_outputs(472)) xor (layer5_outputs(1353));
    layer6_outputs(401) <= not((layer5_outputs(2573)) or (layer5_outputs(18)));
    layer6_outputs(402) <= not(layer5_outputs(4663));
    layer6_outputs(403) <= layer5_outputs(4273);
    layer6_outputs(404) <= layer5_outputs(3523);
    layer6_outputs(405) <= layer5_outputs(680);
    layer6_outputs(406) <= not(layer5_outputs(1670));
    layer6_outputs(407) <= (layer5_outputs(1081)) xor (layer5_outputs(2999));
    layer6_outputs(408) <= not(layer5_outputs(4196));
    layer6_outputs(409) <= layer5_outputs(3875);
    layer6_outputs(410) <= (layer5_outputs(2302)) and not (layer5_outputs(2963));
    layer6_outputs(411) <= layer5_outputs(2828);
    layer6_outputs(412) <= layer5_outputs(4687);
    layer6_outputs(413) <= layer5_outputs(1506);
    layer6_outputs(414) <= layer5_outputs(957);
    layer6_outputs(415) <= (layer5_outputs(3873)) xor (layer5_outputs(3160));
    layer6_outputs(416) <= layer5_outputs(2034);
    layer6_outputs(417) <= layer5_outputs(2027);
    layer6_outputs(418) <= layer5_outputs(3359);
    layer6_outputs(419) <= not(layer5_outputs(865));
    layer6_outputs(420) <= layer5_outputs(488);
    layer6_outputs(421) <= not(layer5_outputs(2226));
    layer6_outputs(422) <= not(layer5_outputs(743));
    layer6_outputs(423) <= (layer5_outputs(549)) xor (layer5_outputs(4665));
    layer6_outputs(424) <= not((layer5_outputs(662)) or (layer5_outputs(3809)));
    layer6_outputs(425) <= (layer5_outputs(3679)) and not (layer5_outputs(4063));
    layer6_outputs(426) <= (layer5_outputs(1051)) or (layer5_outputs(287));
    layer6_outputs(427) <= not((layer5_outputs(2281)) xor (layer5_outputs(2224)));
    layer6_outputs(428) <= not(layer5_outputs(1110));
    layer6_outputs(429) <= not(layer5_outputs(3870));
    layer6_outputs(430) <= layer5_outputs(3079);
    layer6_outputs(431) <= not((layer5_outputs(4100)) xor (layer5_outputs(1320)));
    layer6_outputs(432) <= not(layer5_outputs(1756)) or (layer5_outputs(4167));
    layer6_outputs(433) <= not(layer5_outputs(929)) or (layer5_outputs(1303));
    layer6_outputs(434) <= layer5_outputs(2663);
    layer6_outputs(435) <= not(layer5_outputs(3506));
    layer6_outputs(436) <= '0';
    layer6_outputs(437) <= (layer5_outputs(4712)) xor (layer5_outputs(1404));
    layer6_outputs(438) <= layer5_outputs(1858);
    layer6_outputs(439) <= not((layer5_outputs(1322)) and (layer5_outputs(933)));
    layer6_outputs(440) <= not(layer5_outputs(4872));
    layer6_outputs(441) <= not(layer5_outputs(4487)) or (layer5_outputs(290));
    layer6_outputs(442) <= not((layer5_outputs(4288)) or (layer5_outputs(2374)));
    layer6_outputs(443) <= '1';
    layer6_outputs(444) <= layer5_outputs(2658);
    layer6_outputs(445) <= not(layer5_outputs(3787));
    layer6_outputs(446) <= not(layer5_outputs(283));
    layer6_outputs(447) <= layer5_outputs(4576);
    layer6_outputs(448) <= layer5_outputs(572);
    layer6_outputs(449) <= layer5_outputs(4828);
    layer6_outputs(450) <= not(layer5_outputs(2093));
    layer6_outputs(451) <= not(layer5_outputs(2185));
    layer6_outputs(452) <= layer5_outputs(3222);
    layer6_outputs(453) <= layer5_outputs(3364);
    layer6_outputs(454) <= layer5_outputs(339);
    layer6_outputs(455) <= layer5_outputs(1984);
    layer6_outputs(456) <= (layer5_outputs(3938)) or (layer5_outputs(4619));
    layer6_outputs(457) <= not(layer5_outputs(2494));
    layer6_outputs(458) <= not(layer5_outputs(1115));
    layer6_outputs(459) <= layer5_outputs(370);
    layer6_outputs(460) <= (layer5_outputs(835)) and (layer5_outputs(217));
    layer6_outputs(461) <= (layer5_outputs(3700)) xor (layer5_outputs(2949));
    layer6_outputs(462) <= layer5_outputs(4087);
    layer6_outputs(463) <= not((layer5_outputs(4999)) or (layer5_outputs(1151)));
    layer6_outputs(464) <= (layer5_outputs(3408)) and not (layer5_outputs(40));
    layer6_outputs(465) <= not(layer5_outputs(3764));
    layer6_outputs(466) <= not(layer5_outputs(2797));
    layer6_outputs(467) <= (layer5_outputs(3629)) and (layer5_outputs(232));
    layer6_outputs(468) <= layer5_outputs(274);
    layer6_outputs(469) <= layer5_outputs(3144);
    layer6_outputs(470) <= layer5_outputs(1324);
    layer6_outputs(471) <= (layer5_outputs(3540)) and not (layer5_outputs(2623));
    layer6_outputs(472) <= (layer5_outputs(562)) and not (layer5_outputs(898));
    layer6_outputs(473) <= not(layer5_outputs(1792));
    layer6_outputs(474) <= layer5_outputs(2324);
    layer6_outputs(475) <= not(layer5_outputs(4319));
    layer6_outputs(476) <= not(layer5_outputs(3395));
    layer6_outputs(477) <= not((layer5_outputs(3493)) xor (layer5_outputs(5035)));
    layer6_outputs(478) <= not(layer5_outputs(279));
    layer6_outputs(479) <= not(layer5_outputs(4250));
    layer6_outputs(480) <= not(layer5_outputs(3136));
    layer6_outputs(481) <= layer5_outputs(1341);
    layer6_outputs(482) <= (layer5_outputs(1801)) and not (layer5_outputs(4401));
    layer6_outputs(483) <= not(layer5_outputs(625));
    layer6_outputs(484) <= not(layer5_outputs(4286));
    layer6_outputs(485) <= not(layer5_outputs(960));
    layer6_outputs(486) <= layer5_outputs(2409);
    layer6_outputs(487) <= layer5_outputs(3230);
    layer6_outputs(488) <= not(layer5_outputs(4689)) or (layer5_outputs(1153));
    layer6_outputs(489) <= not((layer5_outputs(4765)) xor (layer5_outputs(4913)));
    layer6_outputs(490) <= not((layer5_outputs(127)) and (layer5_outputs(1070)));
    layer6_outputs(491) <= layer5_outputs(4112);
    layer6_outputs(492) <= (layer5_outputs(3942)) and not (layer5_outputs(1665));
    layer6_outputs(493) <= not(layer5_outputs(4200));
    layer6_outputs(494) <= (layer5_outputs(933)) and not (layer5_outputs(591));
    layer6_outputs(495) <= not(layer5_outputs(70)) or (layer5_outputs(2921));
    layer6_outputs(496) <= layer5_outputs(2708);
    layer6_outputs(497) <= not((layer5_outputs(2585)) xor (layer5_outputs(1441)));
    layer6_outputs(498) <= not(layer5_outputs(4935));
    layer6_outputs(499) <= not(layer5_outputs(4284));
    layer6_outputs(500) <= (layer5_outputs(2148)) xor (layer5_outputs(3209));
    layer6_outputs(501) <= not(layer5_outputs(43));
    layer6_outputs(502) <= layer5_outputs(2411);
    layer6_outputs(503) <= not(layer5_outputs(2220));
    layer6_outputs(504) <= layer5_outputs(265);
    layer6_outputs(505) <= not(layer5_outputs(1814));
    layer6_outputs(506) <= not((layer5_outputs(2649)) xor (layer5_outputs(740)));
    layer6_outputs(507) <= (layer5_outputs(3244)) xor (layer5_outputs(3789));
    layer6_outputs(508) <= not((layer5_outputs(3564)) xor (layer5_outputs(3900)));
    layer6_outputs(509) <= layer5_outputs(2994);
    layer6_outputs(510) <= not((layer5_outputs(1227)) xor (layer5_outputs(521)));
    layer6_outputs(511) <= not(layer5_outputs(1903));
    layer6_outputs(512) <= (layer5_outputs(675)) and not (layer5_outputs(4228));
    layer6_outputs(513) <= not(layer5_outputs(3399)) or (layer5_outputs(2493));
    layer6_outputs(514) <= layer5_outputs(719);
    layer6_outputs(515) <= layer5_outputs(2273);
    layer6_outputs(516) <= (layer5_outputs(2999)) and not (layer5_outputs(1721));
    layer6_outputs(517) <= (layer5_outputs(3590)) or (layer5_outputs(1929));
    layer6_outputs(518) <= not(layer5_outputs(213));
    layer6_outputs(519) <= '0';
    layer6_outputs(520) <= not(layer5_outputs(2794));
    layer6_outputs(521) <= (layer5_outputs(164)) and not (layer5_outputs(3811));
    layer6_outputs(522) <= (layer5_outputs(262)) and not (layer5_outputs(921));
    layer6_outputs(523) <= not(layer5_outputs(2544));
    layer6_outputs(524) <= not(layer5_outputs(3731));
    layer6_outputs(525) <= layer5_outputs(3660);
    layer6_outputs(526) <= (layer5_outputs(3632)) and not (layer5_outputs(805));
    layer6_outputs(527) <= (layer5_outputs(1786)) xor (layer5_outputs(1357));
    layer6_outputs(528) <= not(layer5_outputs(1126)) or (layer5_outputs(3469));
    layer6_outputs(529) <= layer5_outputs(3850);
    layer6_outputs(530) <= not(layer5_outputs(2183)) or (layer5_outputs(3914));
    layer6_outputs(531) <= layer5_outputs(2397);
    layer6_outputs(532) <= not((layer5_outputs(2367)) or (layer5_outputs(4633)));
    layer6_outputs(533) <= not((layer5_outputs(4411)) and (layer5_outputs(963)));
    layer6_outputs(534) <= (layer5_outputs(1443)) and not (layer5_outputs(3624));
    layer6_outputs(535) <= not(layer5_outputs(893));
    layer6_outputs(536) <= not(layer5_outputs(1542));
    layer6_outputs(537) <= not(layer5_outputs(2865));
    layer6_outputs(538) <= '1';
    layer6_outputs(539) <= not(layer5_outputs(1893));
    layer6_outputs(540) <= layer5_outputs(2475);
    layer6_outputs(541) <= layer5_outputs(2632);
    layer6_outputs(542) <= not((layer5_outputs(3112)) or (layer5_outputs(3139)));
    layer6_outputs(543) <= (layer5_outputs(3209)) and (layer5_outputs(5011));
    layer6_outputs(544) <= layer5_outputs(3736);
    layer6_outputs(545) <= not(layer5_outputs(2682));
    layer6_outputs(546) <= not(layer5_outputs(3588));
    layer6_outputs(547) <= (layer5_outputs(1936)) or (layer5_outputs(2477));
    layer6_outputs(548) <= (layer5_outputs(1740)) and (layer5_outputs(2366));
    layer6_outputs(549) <= (layer5_outputs(167)) xor (layer5_outputs(2880));
    layer6_outputs(550) <= layer5_outputs(876);
    layer6_outputs(551) <= layer5_outputs(4469);
    layer6_outputs(552) <= layer5_outputs(3531);
    layer6_outputs(553) <= layer5_outputs(4214);
    layer6_outputs(554) <= not(layer5_outputs(3692));
    layer6_outputs(555) <= not((layer5_outputs(169)) xor (layer5_outputs(1354)));
    layer6_outputs(556) <= not(layer5_outputs(4056));
    layer6_outputs(557) <= layer5_outputs(2694);
    layer6_outputs(558) <= not((layer5_outputs(1451)) and (layer5_outputs(2165)));
    layer6_outputs(559) <= (layer5_outputs(517)) xor (layer5_outputs(4132));
    layer6_outputs(560) <= not(layer5_outputs(4346));
    layer6_outputs(561) <= layer5_outputs(236);
    layer6_outputs(562) <= not(layer5_outputs(1997));
    layer6_outputs(563) <= (layer5_outputs(3288)) or (layer5_outputs(2790));
    layer6_outputs(564) <= not((layer5_outputs(2625)) xor (layer5_outputs(95)));
    layer6_outputs(565) <= layer5_outputs(2304);
    layer6_outputs(566) <= not(layer5_outputs(3301)) or (layer5_outputs(4425));
    layer6_outputs(567) <= layer5_outputs(1484);
    layer6_outputs(568) <= not((layer5_outputs(734)) or (layer5_outputs(983)));
    layer6_outputs(569) <= not(layer5_outputs(810));
    layer6_outputs(570) <= (layer5_outputs(1598)) xor (layer5_outputs(2907));
    layer6_outputs(571) <= layer5_outputs(1206);
    layer6_outputs(572) <= not(layer5_outputs(1882));
    layer6_outputs(573) <= layer5_outputs(4014);
    layer6_outputs(574) <= not(layer5_outputs(2781));
    layer6_outputs(575) <= layer5_outputs(1483);
    layer6_outputs(576) <= not(layer5_outputs(3015)) or (layer5_outputs(1695));
    layer6_outputs(577) <= layer5_outputs(420);
    layer6_outputs(578) <= (layer5_outputs(2961)) and not (layer5_outputs(2060));
    layer6_outputs(579) <= not((layer5_outputs(3971)) and (layer5_outputs(4985)));
    layer6_outputs(580) <= not(layer5_outputs(3378));
    layer6_outputs(581) <= not((layer5_outputs(4627)) xor (layer5_outputs(1230)));
    layer6_outputs(582) <= not(layer5_outputs(876));
    layer6_outputs(583) <= not(layer5_outputs(394));
    layer6_outputs(584) <= layer5_outputs(2529);
    layer6_outputs(585) <= not((layer5_outputs(2821)) xor (layer5_outputs(1646)));
    layer6_outputs(586) <= not(layer5_outputs(3529)) or (layer5_outputs(45));
    layer6_outputs(587) <= not(layer5_outputs(1169));
    layer6_outputs(588) <= not(layer5_outputs(757));
    layer6_outputs(589) <= not((layer5_outputs(4869)) and (layer5_outputs(2274)));
    layer6_outputs(590) <= not((layer5_outputs(261)) or (layer5_outputs(1277)));
    layer6_outputs(591) <= not(layer5_outputs(3608));
    layer6_outputs(592) <= layer5_outputs(3579);
    layer6_outputs(593) <= not(layer5_outputs(623));
    layer6_outputs(594) <= not(layer5_outputs(305));
    layer6_outputs(595) <= (layer5_outputs(2513)) xor (layer5_outputs(4771));
    layer6_outputs(596) <= layer5_outputs(4298);
    layer6_outputs(597) <= layer5_outputs(2004);
    layer6_outputs(598) <= not((layer5_outputs(1291)) and (layer5_outputs(1021)));
    layer6_outputs(599) <= not((layer5_outputs(3829)) xor (layer5_outputs(4130)));
    layer6_outputs(600) <= '0';
    layer6_outputs(601) <= layer5_outputs(1683);
    layer6_outputs(602) <= not(layer5_outputs(4393));
    layer6_outputs(603) <= (layer5_outputs(4133)) and not (layer5_outputs(1596));
    layer6_outputs(604) <= '1';
    layer6_outputs(605) <= layer5_outputs(934);
    layer6_outputs(606) <= (layer5_outputs(582)) xor (layer5_outputs(4548));
    layer6_outputs(607) <= not(layer5_outputs(3891));
    layer6_outputs(608) <= not((layer5_outputs(2434)) xor (layer5_outputs(1233)));
    layer6_outputs(609) <= not(layer5_outputs(1480)) or (layer5_outputs(270));
    layer6_outputs(610) <= (layer5_outputs(1207)) xor (layer5_outputs(1455));
    layer6_outputs(611) <= not(layer5_outputs(882)) or (layer5_outputs(5009));
    layer6_outputs(612) <= not(layer5_outputs(3169));
    layer6_outputs(613) <= (layer5_outputs(3413)) xor (layer5_outputs(3380));
    layer6_outputs(614) <= layer5_outputs(1666);
    layer6_outputs(615) <= layer5_outputs(2722);
    layer6_outputs(616) <= (layer5_outputs(4194)) and not (layer5_outputs(1824));
    layer6_outputs(617) <= not(layer5_outputs(3779));
    layer6_outputs(618) <= layer5_outputs(2106);
    layer6_outputs(619) <= not(layer5_outputs(2256));
    layer6_outputs(620) <= not(layer5_outputs(1500));
    layer6_outputs(621) <= (layer5_outputs(1816)) or (layer5_outputs(4960));
    layer6_outputs(622) <= not(layer5_outputs(1210));
    layer6_outputs(623) <= layer5_outputs(2528);
    layer6_outputs(624) <= layer5_outputs(3053);
    layer6_outputs(625) <= not((layer5_outputs(2963)) xor (layer5_outputs(1486)));
    layer6_outputs(626) <= not(layer5_outputs(1237)) or (layer5_outputs(2259));
    layer6_outputs(627) <= (layer5_outputs(1988)) or (layer5_outputs(5026));
    layer6_outputs(628) <= not(layer5_outputs(140)) or (layer5_outputs(1437));
    layer6_outputs(629) <= layer5_outputs(3631);
    layer6_outputs(630) <= layer5_outputs(3477);
    layer6_outputs(631) <= layer5_outputs(3694);
    layer6_outputs(632) <= not(layer5_outputs(474));
    layer6_outputs(633) <= not(layer5_outputs(3492));
    layer6_outputs(634) <= not((layer5_outputs(293)) xor (layer5_outputs(3439)));
    layer6_outputs(635) <= not(layer5_outputs(2112));
    layer6_outputs(636) <= not(layer5_outputs(3225));
    layer6_outputs(637) <= not(layer5_outputs(3996));
    layer6_outputs(638) <= (layer5_outputs(44)) and not (layer5_outputs(878));
    layer6_outputs(639) <= layer5_outputs(3703);
    layer6_outputs(640) <= layer5_outputs(3734);
    layer6_outputs(641) <= (layer5_outputs(3103)) or (layer5_outputs(3386));
    layer6_outputs(642) <= (layer5_outputs(2056)) and not (layer5_outputs(1902));
    layer6_outputs(643) <= (layer5_outputs(769)) and not (layer5_outputs(4422));
    layer6_outputs(644) <= (layer5_outputs(1219)) and not (layer5_outputs(4140));
    layer6_outputs(645) <= not(layer5_outputs(960));
    layer6_outputs(646) <= layer5_outputs(2702);
    layer6_outputs(647) <= not((layer5_outputs(4924)) xor (layer5_outputs(4668)));
    layer6_outputs(648) <= not(layer5_outputs(791));
    layer6_outputs(649) <= layer5_outputs(4201);
    layer6_outputs(650) <= not(layer5_outputs(1391));
    layer6_outputs(651) <= layer5_outputs(2678);
    layer6_outputs(652) <= (layer5_outputs(1286)) xor (layer5_outputs(139));
    layer6_outputs(653) <= layer5_outputs(795);
    layer6_outputs(654) <= not(layer5_outputs(3100)) or (layer5_outputs(2157));
    layer6_outputs(655) <= not((layer5_outputs(4255)) and (layer5_outputs(1454)));
    layer6_outputs(656) <= not(layer5_outputs(1806));
    layer6_outputs(657) <= not(layer5_outputs(2068));
    layer6_outputs(658) <= not((layer5_outputs(2618)) or (layer5_outputs(3174)));
    layer6_outputs(659) <= not(layer5_outputs(2271)) or (layer5_outputs(1511));
    layer6_outputs(660) <= (layer5_outputs(2131)) or (layer5_outputs(3761));
    layer6_outputs(661) <= not(layer5_outputs(737));
    layer6_outputs(662) <= '0';
    layer6_outputs(663) <= (layer5_outputs(2764)) and (layer5_outputs(1362));
    layer6_outputs(664) <= (layer5_outputs(943)) xor (layer5_outputs(2430));
    layer6_outputs(665) <= not(layer5_outputs(3314));
    layer6_outputs(666) <= (layer5_outputs(600)) and not (layer5_outputs(2336));
    layer6_outputs(667) <= '1';
    layer6_outputs(668) <= layer5_outputs(3657);
    layer6_outputs(669) <= not(layer5_outputs(815));
    layer6_outputs(670) <= not(layer5_outputs(4360)) or (layer5_outputs(3409));
    layer6_outputs(671) <= not(layer5_outputs(4948)) or (layer5_outputs(4699));
    layer6_outputs(672) <= not(layer5_outputs(3847));
    layer6_outputs(673) <= not(layer5_outputs(2185));
    layer6_outputs(674) <= (layer5_outputs(869)) and (layer5_outputs(2853));
    layer6_outputs(675) <= not(layer5_outputs(918)) or (layer5_outputs(3159));
    layer6_outputs(676) <= (layer5_outputs(88)) and (layer5_outputs(1609));
    layer6_outputs(677) <= not(layer5_outputs(1685)) or (layer5_outputs(1091));
    layer6_outputs(678) <= not(layer5_outputs(907));
    layer6_outputs(679) <= layer5_outputs(2838);
    layer6_outputs(680) <= (layer5_outputs(4797)) and not (layer5_outputs(1066));
    layer6_outputs(681) <= layer5_outputs(213);
    layer6_outputs(682) <= not(layer5_outputs(4313));
    layer6_outputs(683) <= not((layer5_outputs(482)) xor (layer5_outputs(3048)));
    layer6_outputs(684) <= not((layer5_outputs(2798)) xor (layer5_outputs(2858)));
    layer6_outputs(685) <= layer5_outputs(3567);
    layer6_outputs(686) <= (layer5_outputs(146)) and not (layer5_outputs(2052));
    layer6_outputs(687) <= layer5_outputs(4375);
    layer6_outputs(688) <= not(layer5_outputs(3137));
    layer6_outputs(689) <= layer5_outputs(3421);
    layer6_outputs(690) <= layer5_outputs(331);
    layer6_outputs(691) <= (layer5_outputs(4565)) and not (layer5_outputs(4422));
    layer6_outputs(692) <= layer5_outputs(4414);
    layer6_outputs(693) <= not(layer5_outputs(3141));
    layer6_outputs(694) <= layer5_outputs(472);
    layer6_outputs(695) <= not(layer5_outputs(601)) or (layer5_outputs(2616));
    layer6_outputs(696) <= (layer5_outputs(675)) or (layer5_outputs(4205));
    layer6_outputs(697) <= not((layer5_outputs(1973)) and (layer5_outputs(2986)));
    layer6_outputs(698) <= not(layer5_outputs(3011));
    layer6_outputs(699) <= not(layer5_outputs(365));
    layer6_outputs(700) <= (layer5_outputs(1655)) or (layer5_outputs(655));
    layer6_outputs(701) <= not((layer5_outputs(2307)) xor (layer5_outputs(4586)));
    layer6_outputs(702) <= not(layer5_outputs(3369));
    layer6_outputs(703) <= not((layer5_outputs(314)) and (layer5_outputs(1270)));
    layer6_outputs(704) <= not(layer5_outputs(1166));
    layer6_outputs(705) <= layer5_outputs(3289);
    layer6_outputs(706) <= not((layer5_outputs(2563)) and (layer5_outputs(2114)));
    layer6_outputs(707) <= layer5_outputs(4918);
    layer6_outputs(708) <= (layer5_outputs(4310)) and not (layer5_outputs(1337));
    layer6_outputs(709) <= (layer5_outputs(3961)) xor (layer5_outputs(2645));
    layer6_outputs(710) <= layer5_outputs(2318);
    layer6_outputs(711) <= not(layer5_outputs(2892));
    layer6_outputs(712) <= not((layer5_outputs(3640)) or (layer5_outputs(4472)));
    layer6_outputs(713) <= not(layer5_outputs(4658));
    layer6_outputs(714) <= not(layer5_outputs(481));
    layer6_outputs(715) <= not(layer5_outputs(4718));
    layer6_outputs(716) <= not(layer5_outputs(4590));
    layer6_outputs(717) <= not((layer5_outputs(193)) xor (layer5_outputs(4185)));
    layer6_outputs(718) <= not(layer5_outputs(3865));
    layer6_outputs(719) <= (layer5_outputs(2888)) and not (layer5_outputs(4894));
    layer6_outputs(720) <= (layer5_outputs(595)) and (layer5_outputs(3276));
    layer6_outputs(721) <= layer5_outputs(2926);
    layer6_outputs(722) <= not(layer5_outputs(438));
    layer6_outputs(723) <= layer5_outputs(2873);
    layer6_outputs(724) <= (layer5_outputs(1426)) or (layer5_outputs(690));
    layer6_outputs(725) <= layer5_outputs(3904);
    layer6_outputs(726) <= layer5_outputs(4612);
    layer6_outputs(727) <= (layer5_outputs(1097)) or (layer5_outputs(101));
    layer6_outputs(728) <= not((layer5_outputs(3403)) xor (layer5_outputs(1895)));
    layer6_outputs(729) <= not(layer5_outputs(1006)) or (layer5_outputs(4499));
    layer6_outputs(730) <= not((layer5_outputs(849)) and (layer5_outputs(1640)));
    layer6_outputs(731) <= not(layer5_outputs(3544));
    layer6_outputs(732) <= layer5_outputs(4888);
    layer6_outputs(733) <= not(layer5_outputs(3191));
    layer6_outputs(734) <= not(layer5_outputs(3470));
    layer6_outputs(735) <= not(layer5_outputs(835));
    layer6_outputs(736) <= layer5_outputs(4176);
    layer6_outputs(737) <= layer5_outputs(4107);
    layer6_outputs(738) <= not(layer5_outputs(1669));
    layer6_outputs(739) <= layer5_outputs(3805);
    layer6_outputs(740) <= (layer5_outputs(3572)) and not (layer5_outputs(4146));
    layer6_outputs(741) <= not(layer5_outputs(1158));
    layer6_outputs(742) <= not((layer5_outputs(4090)) or (layer5_outputs(4736)));
    layer6_outputs(743) <= (layer5_outputs(436)) or (layer5_outputs(4848));
    layer6_outputs(744) <= layer5_outputs(1154);
    layer6_outputs(745) <= not((layer5_outputs(524)) and (layer5_outputs(1835)));
    layer6_outputs(746) <= layer5_outputs(1519);
    layer6_outputs(747) <= not(layer5_outputs(4115));
    layer6_outputs(748) <= not(layer5_outputs(2066));
    layer6_outputs(749) <= (layer5_outputs(4121)) or (layer5_outputs(3245));
    layer6_outputs(750) <= (layer5_outputs(3051)) or (layer5_outputs(4910));
    layer6_outputs(751) <= (layer5_outputs(3027)) and not (layer5_outputs(1984));
    layer6_outputs(752) <= layer5_outputs(3962);
    layer6_outputs(753) <= not((layer5_outputs(3445)) xor (layer5_outputs(3597)));
    layer6_outputs(754) <= (layer5_outputs(2921)) and not (layer5_outputs(2222));
    layer6_outputs(755) <= not((layer5_outputs(3220)) and (layer5_outputs(3543)));
    layer6_outputs(756) <= not(layer5_outputs(5048)) or (layer5_outputs(1347));
    layer6_outputs(757) <= not(layer5_outputs(1651));
    layer6_outputs(758) <= layer5_outputs(4931);
    layer6_outputs(759) <= not(layer5_outputs(4405));
    layer6_outputs(760) <= layer5_outputs(545);
    layer6_outputs(761) <= not((layer5_outputs(1777)) xor (layer5_outputs(1321)));
    layer6_outputs(762) <= not(layer5_outputs(603));
    layer6_outputs(763) <= not((layer5_outputs(2705)) or (layer5_outputs(3878)));
    layer6_outputs(764) <= not((layer5_outputs(1165)) and (layer5_outputs(2541)));
    layer6_outputs(765) <= '1';
    layer6_outputs(766) <= (layer5_outputs(4697)) and not (layer5_outputs(2619));
    layer6_outputs(767) <= layer5_outputs(3301);
    layer6_outputs(768) <= layer5_outputs(4228);
    layer6_outputs(769) <= not(layer5_outputs(203));
    layer6_outputs(770) <= layer5_outputs(4790);
    layer6_outputs(771) <= (layer5_outputs(2889)) or (layer5_outputs(3013));
    layer6_outputs(772) <= (layer5_outputs(770)) or (layer5_outputs(3585));
    layer6_outputs(773) <= not((layer5_outputs(1297)) and (layer5_outputs(3473)));
    layer6_outputs(774) <= layer5_outputs(3035);
    layer6_outputs(775) <= not(layer5_outputs(4518));
    layer6_outputs(776) <= (layer5_outputs(1545)) or (layer5_outputs(1470));
    layer6_outputs(777) <= layer5_outputs(909);
    layer6_outputs(778) <= not(layer5_outputs(3915));
    layer6_outputs(779) <= layer5_outputs(3295);
    layer6_outputs(780) <= not(layer5_outputs(3640));
    layer6_outputs(781) <= not(layer5_outputs(1900)) or (layer5_outputs(2478));
    layer6_outputs(782) <= not(layer5_outputs(5008));
    layer6_outputs(783) <= not((layer5_outputs(1854)) and (layer5_outputs(3345)));
    layer6_outputs(784) <= layer5_outputs(1561);
    layer6_outputs(785) <= not((layer5_outputs(2211)) xor (layer5_outputs(2294)));
    layer6_outputs(786) <= not(layer5_outputs(2571));
    layer6_outputs(787) <= not((layer5_outputs(4859)) xor (layer5_outputs(2977)));
    layer6_outputs(788) <= layer5_outputs(1472);
    layer6_outputs(789) <= not(layer5_outputs(2910));
    layer6_outputs(790) <= not(layer5_outputs(2255));
    layer6_outputs(791) <= (layer5_outputs(1825)) and (layer5_outputs(2275));
    layer6_outputs(792) <= not(layer5_outputs(4763)) or (layer5_outputs(134));
    layer6_outputs(793) <= not((layer5_outputs(3801)) and (layer5_outputs(4636)));
    layer6_outputs(794) <= layer5_outputs(3061);
    layer6_outputs(795) <= layer5_outputs(3940);
    layer6_outputs(796) <= layer5_outputs(4502);
    layer6_outputs(797) <= layer5_outputs(3311);
    layer6_outputs(798) <= (layer5_outputs(1231)) or (layer5_outputs(4098));
    layer6_outputs(799) <= not(layer5_outputs(1299));
    layer6_outputs(800) <= not(layer5_outputs(1868));
    layer6_outputs(801) <= not(layer5_outputs(4377)) or (layer5_outputs(3083));
    layer6_outputs(802) <= not((layer5_outputs(3023)) xor (layer5_outputs(4204)));
    layer6_outputs(803) <= not(layer5_outputs(2962));
    layer6_outputs(804) <= not(layer5_outputs(5108));
    layer6_outputs(805) <= not(layer5_outputs(660));
    layer6_outputs(806) <= layer5_outputs(4127);
    layer6_outputs(807) <= layer5_outputs(3949);
    layer6_outputs(808) <= not((layer5_outputs(4806)) xor (layer5_outputs(4528)));
    layer6_outputs(809) <= not(layer5_outputs(163)) or (layer5_outputs(945));
    layer6_outputs(810) <= not((layer5_outputs(2228)) and (layer5_outputs(5055)));
    layer6_outputs(811) <= (layer5_outputs(1942)) and (layer5_outputs(1608));
    layer6_outputs(812) <= (layer5_outputs(4764)) and not (layer5_outputs(2231));
    layer6_outputs(813) <= layer5_outputs(2018);
    layer6_outputs(814) <= layer5_outputs(57);
    layer6_outputs(815) <= not(layer5_outputs(4777));
    layer6_outputs(816) <= not(layer5_outputs(1348));
    layer6_outputs(817) <= layer5_outputs(179);
    layer6_outputs(818) <= (layer5_outputs(5055)) and not (layer5_outputs(4484));
    layer6_outputs(819) <= not(layer5_outputs(3193));
    layer6_outputs(820) <= not(layer5_outputs(1326));
    layer6_outputs(821) <= '0';
    layer6_outputs(822) <= (layer5_outputs(4354)) or (layer5_outputs(2802));
    layer6_outputs(823) <= (layer5_outputs(1819)) or (layer5_outputs(1911));
    layer6_outputs(824) <= (layer5_outputs(4617)) and not (layer5_outputs(1724));
    layer6_outputs(825) <= layer5_outputs(313);
    layer6_outputs(826) <= layer5_outputs(3680);
    layer6_outputs(827) <= (layer5_outputs(1461)) and not (layer5_outputs(175));
    layer6_outputs(828) <= not(layer5_outputs(1307));
    layer6_outputs(829) <= layer5_outputs(776);
    layer6_outputs(830) <= not(layer5_outputs(3155));
    layer6_outputs(831) <= layer5_outputs(2016);
    layer6_outputs(832) <= not(layer5_outputs(4268));
    layer6_outputs(833) <= (layer5_outputs(1971)) xor (layer5_outputs(2719));
    layer6_outputs(834) <= layer5_outputs(4409);
    layer6_outputs(835) <= layer5_outputs(4240);
    layer6_outputs(836) <= not(layer5_outputs(613));
    layer6_outputs(837) <= (layer5_outputs(4451)) or (layer5_outputs(3509));
    layer6_outputs(838) <= not(layer5_outputs(3321)) or (layer5_outputs(1043));
    layer6_outputs(839) <= layer5_outputs(3268);
    layer6_outputs(840) <= not(layer5_outputs(996));
    layer6_outputs(841) <= not(layer5_outputs(1244));
    layer6_outputs(842) <= layer5_outputs(1279);
    layer6_outputs(843) <= layer5_outputs(1657);
    layer6_outputs(844) <= not(layer5_outputs(3800));
    layer6_outputs(845) <= not(layer5_outputs(2825));
    layer6_outputs(846) <= layer5_outputs(739);
    layer6_outputs(847) <= layer5_outputs(2427);
    layer6_outputs(848) <= not((layer5_outputs(4681)) or (layer5_outputs(4337)));
    layer6_outputs(849) <= layer5_outputs(813);
    layer6_outputs(850) <= not(layer5_outputs(3819)) or (layer5_outputs(1737));
    layer6_outputs(851) <= not(layer5_outputs(2551)) or (layer5_outputs(3476));
    layer6_outputs(852) <= (layer5_outputs(4666)) or (layer5_outputs(3533));
    layer6_outputs(853) <= not(layer5_outputs(4488));
    layer6_outputs(854) <= (layer5_outputs(2264)) or (layer5_outputs(159));
    layer6_outputs(855) <= layer5_outputs(4906);
    layer6_outputs(856) <= not(layer5_outputs(2701));
    layer6_outputs(857) <= not(layer5_outputs(2386)) or (layer5_outputs(3673));
    layer6_outputs(858) <= layer5_outputs(4079);
    layer6_outputs(859) <= not(layer5_outputs(3000));
    layer6_outputs(860) <= not(layer5_outputs(4494));
    layer6_outputs(861) <= layer5_outputs(5097);
    layer6_outputs(862) <= not((layer5_outputs(97)) or (layer5_outputs(3504)));
    layer6_outputs(863) <= not((layer5_outputs(2463)) and (layer5_outputs(3761)));
    layer6_outputs(864) <= (layer5_outputs(3258)) and not (layer5_outputs(3845));
    layer6_outputs(865) <= (layer5_outputs(3988)) and not (layer5_outputs(1802));
    layer6_outputs(866) <= not((layer5_outputs(2337)) xor (layer5_outputs(839)));
    layer6_outputs(867) <= not(layer5_outputs(3393));
    layer6_outputs(868) <= layer5_outputs(2110);
    layer6_outputs(869) <= not(layer5_outputs(1393));
    layer6_outputs(870) <= (layer5_outputs(5074)) and not (layer5_outputs(2612));
    layer6_outputs(871) <= not(layer5_outputs(2171));
    layer6_outputs(872) <= not((layer5_outputs(3513)) or (layer5_outputs(293)));
    layer6_outputs(873) <= (layer5_outputs(4169)) and (layer5_outputs(1154));
    layer6_outputs(874) <= not(layer5_outputs(3597)) or (layer5_outputs(1593));
    layer6_outputs(875) <= not(layer5_outputs(2729)) or (layer5_outputs(284));
    layer6_outputs(876) <= not((layer5_outputs(24)) and (layer5_outputs(2061)));
    layer6_outputs(877) <= layer5_outputs(4410);
    layer6_outputs(878) <= not(layer5_outputs(3970));
    layer6_outputs(879) <= not((layer5_outputs(1293)) xor (layer5_outputs(447)));
    layer6_outputs(880) <= (layer5_outputs(4983)) and not (layer5_outputs(3178));
    layer6_outputs(881) <= not(layer5_outputs(3481));
    layer6_outputs(882) <= not(layer5_outputs(4091));
    layer6_outputs(883) <= (layer5_outputs(1761)) and not (layer5_outputs(3456));
    layer6_outputs(884) <= not(layer5_outputs(1862));
    layer6_outputs(885) <= not(layer5_outputs(1495));
    layer6_outputs(886) <= not(layer5_outputs(2254)) or (layer5_outputs(3281));
    layer6_outputs(887) <= not((layer5_outputs(4986)) and (layer5_outputs(3362)));
    layer6_outputs(888) <= (layer5_outputs(4927)) xor (layer5_outputs(2507));
    layer6_outputs(889) <= not(layer5_outputs(499));
    layer6_outputs(890) <= not(layer5_outputs(4720));
    layer6_outputs(891) <= (layer5_outputs(1837)) xor (layer5_outputs(3545));
    layer6_outputs(892) <= layer5_outputs(2040);
    layer6_outputs(893) <= (layer5_outputs(608)) and not (layer5_outputs(4232));
    layer6_outputs(894) <= (layer5_outputs(4085)) and not (layer5_outputs(1068));
    layer6_outputs(895) <= layer5_outputs(5027);
    layer6_outputs(896) <= (layer5_outputs(1682)) xor (layer5_outputs(1982));
    layer6_outputs(897) <= (layer5_outputs(878)) and (layer5_outputs(2238));
    layer6_outputs(898) <= not((layer5_outputs(717)) xor (layer5_outputs(3811)));
    layer6_outputs(899) <= not((layer5_outputs(2586)) and (layer5_outputs(1956)));
    layer6_outputs(900) <= not(layer5_outputs(2330));
    layer6_outputs(901) <= (layer5_outputs(622)) and (layer5_outputs(421));
    layer6_outputs(902) <= not(layer5_outputs(1988)) or (layer5_outputs(4432));
    layer6_outputs(903) <= layer5_outputs(4737);
    layer6_outputs(904) <= (layer5_outputs(3625)) or (layer5_outputs(1487));
    layer6_outputs(905) <= (layer5_outputs(4119)) and not (layer5_outputs(4506));
    layer6_outputs(906) <= (layer5_outputs(3085)) and (layer5_outputs(4663));
    layer6_outputs(907) <= layer5_outputs(2068);
    layer6_outputs(908) <= not(layer5_outputs(5000)) or (layer5_outputs(2572));
    layer6_outputs(909) <= layer5_outputs(2540);
    layer6_outputs(910) <= (layer5_outputs(3792)) and (layer5_outputs(4494));
    layer6_outputs(911) <= layer5_outputs(704);
    layer6_outputs(912) <= not(layer5_outputs(4717));
    layer6_outputs(913) <= layer5_outputs(1726);
    layer6_outputs(914) <= not(layer5_outputs(1865));
    layer6_outputs(915) <= not(layer5_outputs(3552)) or (layer5_outputs(1768));
    layer6_outputs(916) <= (layer5_outputs(2186)) and (layer5_outputs(2626));
    layer6_outputs(917) <= layer5_outputs(3992);
    layer6_outputs(918) <= not(layer5_outputs(4159));
    layer6_outputs(919) <= not(layer5_outputs(4418));
    layer6_outputs(920) <= not(layer5_outputs(2249));
    layer6_outputs(921) <= not(layer5_outputs(350));
    layer6_outputs(922) <= not((layer5_outputs(4868)) and (layer5_outputs(3703)));
    layer6_outputs(923) <= not((layer5_outputs(2944)) or (layer5_outputs(5114)));
    layer6_outputs(924) <= (layer5_outputs(654)) and (layer5_outputs(910));
    layer6_outputs(925) <= (layer5_outputs(4721)) or (layer5_outputs(4788));
    layer6_outputs(926) <= layer5_outputs(1181);
    layer6_outputs(927) <= not(layer5_outputs(3899));
    layer6_outputs(928) <= not(layer5_outputs(5057));
    layer6_outputs(929) <= not(layer5_outputs(997));
    layer6_outputs(930) <= (layer5_outputs(3353)) or (layer5_outputs(1752));
    layer6_outputs(931) <= not(layer5_outputs(4108));
    layer6_outputs(932) <= not(layer5_outputs(437));
    layer6_outputs(933) <= layer5_outputs(3879);
    layer6_outputs(934) <= not(layer5_outputs(3622)) or (layer5_outputs(2154));
    layer6_outputs(935) <= layer5_outputs(2291);
    layer6_outputs(936) <= not(layer5_outputs(3152));
    layer6_outputs(937) <= layer5_outputs(2359);
    layer6_outputs(938) <= not((layer5_outputs(1574)) or (layer5_outputs(1044)));
    layer6_outputs(939) <= layer5_outputs(3280);
    layer6_outputs(940) <= (layer5_outputs(5030)) and not (layer5_outputs(413));
    layer6_outputs(941) <= not(layer5_outputs(1208)) or (layer5_outputs(126));
    layer6_outputs(942) <= layer5_outputs(3939);
    layer6_outputs(943) <= not((layer5_outputs(340)) or (layer5_outputs(1716)));
    layer6_outputs(944) <= layer5_outputs(2910);
    layer6_outputs(945) <= not(layer5_outputs(4381));
    layer6_outputs(946) <= (layer5_outputs(2095)) or (layer5_outputs(566));
    layer6_outputs(947) <= layer5_outputs(1204);
    layer6_outputs(948) <= (layer5_outputs(3452)) or (layer5_outputs(3735));
    layer6_outputs(949) <= layer5_outputs(1832);
    layer6_outputs(950) <= not(layer5_outputs(4585));
    layer6_outputs(951) <= not((layer5_outputs(705)) and (layer5_outputs(2089)));
    layer6_outputs(952) <= (layer5_outputs(1581)) and not (layer5_outputs(1203));
    layer6_outputs(953) <= layer5_outputs(3131);
    layer6_outputs(954) <= not(layer5_outputs(3825));
    layer6_outputs(955) <= not(layer5_outputs(1008));
    layer6_outputs(956) <= not((layer5_outputs(3930)) xor (layer5_outputs(4611)));
    layer6_outputs(957) <= not(layer5_outputs(2912));
    layer6_outputs(958) <= (layer5_outputs(2227)) or (layer5_outputs(2099));
    layer6_outputs(959) <= not(layer5_outputs(2688));
    layer6_outputs(960) <= (layer5_outputs(4103)) and (layer5_outputs(626));
    layer6_outputs(961) <= not((layer5_outputs(3086)) xor (layer5_outputs(3752)));
    layer6_outputs(962) <= not((layer5_outputs(3883)) xor (layer5_outputs(2929)));
    layer6_outputs(963) <= not(layer5_outputs(360));
    layer6_outputs(964) <= not(layer5_outputs(377));
    layer6_outputs(965) <= (layer5_outputs(459)) and (layer5_outputs(1697));
    layer6_outputs(966) <= not(layer5_outputs(3878));
    layer6_outputs(967) <= layer5_outputs(2454);
    layer6_outputs(968) <= not(layer5_outputs(459));
    layer6_outputs(969) <= layer5_outputs(4019);
    layer6_outputs(970) <= (layer5_outputs(4839)) and not (layer5_outputs(4230));
    layer6_outputs(971) <= (layer5_outputs(2537)) xor (layer5_outputs(4322));
    layer6_outputs(972) <= not((layer5_outputs(2479)) or (layer5_outputs(3046)));
    layer6_outputs(973) <= layer5_outputs(3359);
    layer6_outputs(974) <= not(layer5_outputs(1202));
    layer6_outputs(975) <= layer5_outputs(1084);
    layer6_outputs(976) <= layer5_outputs(3182);
    layer6_outputs(977) <= layer5_outputs(1155);
    layer6_outputs(978) <= layer5_outputs(4416);
    layer6_outputs(979) <= not(layer5_outputs(2775));
    layer6_outputs(980) <= (layer5_outputs(1527)) or (layer5_outputs(4715));
    layer6_outputs(981) <= not(layer5_outputs(1535)) or (layer5_outputs(4692));
    layer6_outputs(982) <= not((layer5_outputs(461)) xor (layer5_outputs(1509)));
    layer6_outputs(983) <= layer5_outputs(4278);
    layer6_outputs(984) <= not(layer5_outputs(5110)) or (layer5_outputs(3173));
    layer6_outputs(985) <= layer5_outputs(1847);
    layer6_outputs(986) <= not(layer5_outputs(3873)) or (layer5_outputs(2257));
    layer6_outputs(987) <= layer5_outputs(5049);
    layer6_outputs(988) <= (layer5_outputs(4170)) xor (layer5_outputs(3333));
    layer6_outputs(989) <= not(layer5_outputs(645));
    layer6_outputs(990) <= layer5_outputs(4608);
    layer6_outputs(991) <= not((layer5_outputs(961)) xor (layer5_outputs(4398)));
    layer6_outputs(992) <= not(layer5_outputs(4084));
    layer6_outputs(993) <= not(layer5_outputs(4532));
    layer6_outputs(994) <= (layer5_outputs(811)) and (layer5_outputs(913));
    layer6_outputs(995) <= layer5_outputs(3357);
    layer6_outputs(996) <= layer5_outputs(3404);
    layer6_outputs(997) <= not(layer5_outputs(3812));
    layer6_outputs(998) <= (layer5_outputs(2616)) xor (layer5_outputs(3080));
    layer6_outputs(999) <= layer5_outputs(2071);
    layer6_outputs(1000) <= not(layer5_outputs(971));
    layer6_outputs(1001) <= not(layer5_outputs(1588));
    layer6_outputs(1002) <= layer5_outputs(15);
    layer6_outputs(1003) <= (layer5_outputs(2972)) xor (layer5_outputs(1015));
    layer6_outputs(1004) <= layer5_outputs(3335);
    layer6_outputs(1005) <= not((layer5_outputs(3567)) or (layer5_outputs(3326)));
    layer6_outputs(1006) <= not((layer5_outputs(1695)) and (layer5_outputs(3883)));
    layer6_outputs(1007) <= (layer5_outputs(3835)) and not (layer5_outputs(5009));
    layer6_outputs(1008) <= layer5_outputs(3001);
    layer6_outputs(1009) <= not((layer5_outputs(4758)) or (layer5_outputs(1065)));
    layer6_outputs(1010) <= not(layer5_outputs(4779)) or (layer5_outputs(4823));
    layer6_outputs(1011) <= not((layer5_outputs(2038)) xor (layer5_outputs(2604)));
    layer6_outputs(1012) <= layer5_outputs(3067);
    layer6_outputs(1013) <= layer5_outputs(4579);
    layer6_outputs(1014) <= layer5_outputs(491);
    layer6_outputs(1015) <= layer5_outputs(110);
    layer6_outputs(1016) <= layer5_outputs(43);
    layer6_outputs(1017) <= layer5_outputs(1332);
    layer6_outputs(1018) <= not((layer5_outputs(4057)) or (layer5_outputs(1649)));
    layer6_outputs(1019) <= '1';
    layer6_outputs(1020) <= layer5_outputs(2555);
    layer6_outputs(1021) <= not((layer5_outputs(3020)) and (layer5_outputs(2115)));
    layer6_outputs(1022) <= not((layer5_outputs(2024)) xor (layer5_outputs(2650)));
    layer6_outputs(1023) <= not(layer5_outputs(4568)) or (layer5_outputs(3937));
    layer6_outputs(1024) <= not((layer5_outputs(171)) xor (layer5_outputs(862)));
    layer6_outputs(1025) <= layer5_outputs(4465);
    layer6_outputs(1026) <= not((layer5_outputs(5107)) or (layer5_outputs(1387)));
    layer6_outputs(1027) <= layer5_outputs(862);
    layer6_outputs(1028) <= not(layer5_outputs(2100));
    layer6_outputs(1029) <= not(layer5_outputs(2728));
    layer6_outputs(1030) <= not(layer5_outputs(3729));
    layer6_outputs(1031) <= layer5_outputs(79);
    layer6_outputs(1032) <= not(layer5_outputs(4455));
    layer6_outputs(1033) <= not(layer5_outputs(3947)) or (layer5_outputs(2130));
    layer6_outputs(1034) <= layer5_outputs(816);
    layer6_outputs(1035) <= (layer5_outputs(3986)) and not (layer5_outputs(2152));
    layer6_outputs(1036) <= not((layer5_outputs(3425)) xor (layer5_outputs(4609)));
    layer6_outputs(1037) <= not(layer5_outputs(2593));
    layer6_outputs(1038) <= not(layer5_outputs(4316));
    layer6_outputs(1039) <= layer5_outputs(4202);
    layer6_outputs(1040) <= not(layer5_outputs(1787));
    layer6_outputs(1041) <= layer5_outputs(4254);
    layer6_outputs(1042) <= (layer5_outputs(444)) and (layer5_outputs(4636));
    layer6_outputs(1043) <= (layer5_outputs(4583)) and not (layer5_outputs(609));
    layer6_outputs(1044) <= (layer5_outputs(604)) xor (layer5_outputs(4282));
    layer6_outputs(1045) <= layer5_outputs(2122);
    layer6_outputs(1046) <= not(layer5_outputs(2677));
    layer6_outputs(1047) <= (layer5_outputs(4171)) and not (layer5_outputs(286));
    layer6_outputs(1048) <= layer5_outputs(4354);
    layer6_outputs(1049) <= layer5_outputs(1153);
    layer6_outputs(1050) <= not(layer5_outputs(3165));
    layer6_outputs(1051) <= '0';
    layer6_outputs(1052) <= not(layer5_outputs(2515));
    layer6_outputs(1053) <= layer5_outputs(1875);
    layer6_outputs(1054) <= layer5_outputs(2198);
    layer6_outputs(1055) <= not(layer5_outputs(1384));
    layer6_outputs(1056) <= not(layer5_outputs(1351));
    layer6_outputs(1057) <= not((layer5_outputs(4201)) xor (layer5_outputs(2283)));
    layer6_outputs(1058) <= (layer5_outputs(1)) and not (layer5_outputs(2934));
    layer6_outputs(1059) <= not(layer5_outputs(1570));
    layer6_outputs(1060) <= not(layer5_outputs(51));
    layer6_outputs(1061) <= (layer5_outputs(2666)) and not (layer5_outputs(2077));
    layer6_outputs(1062) <= not((layer5_outputs(5076)) and (layer5_outputs(3981)));
    layer6_outputs(1063) <= layer5_outputs(242);
    layer6_outputs(1064) <= not(layer5_outputs(1463));
    layer6_outputs(1065) <= layer5_outputs(2419);
    layer6_outputs(1066) <= not(layer5_outputs(4618));
    layer6_outputs(1067) <= layer5_outputs(4827);
    layer6_outputs(1068) <= not(layer5_outputs(4344));
    layer6_outputs(1069) <= layer5_outputs(100);
    layer6_outputs(1070) <= (layer5_outputs(853)) and not (layer5_outputs(4734));
    layer6_outputs(1071) <= not(layer5_outputs(281));
    layer6_outputs(1072) <= not(layer5_outputs(3669));
    layer6_outputs(1073) <= (layer5_outputs(215)) or (layer5_outputs(4574));
    layer6_outputs(1074) <= (layer5_outputs(3568)) or (layer5_outputs(2208));
    layer6_outputs(1075) <= not(layer5_outputs(4740));
    layer6_outputs(1076) <= layer5_outputs(4626);
    layer6_outputs(1077) <= not((layer5_outputs(2459)) and (layer5_outputs(3759)));
    layer6_outputs(1078) <= (layer5_outputs(4932)) xor (layer5_outputs(32));
    layer6_outputs(1079) <= not((layer5_outputs(4220)) xor (layer5_outputs(1722)));
    layer6_outputs(1080) <= layer5_outputs(5063);
    layer6_outputs(1081) <= not(layer5_outputs(23)) or (layer5_outputs(4125));
    layer6_outputs(1082) <= not(layer5_outputs(616));
    layer6_outputs(1083) <= not(layer5_outputs(2894));
    layer6_outputs(1084) <= not(layer5_outputs(2001));
    layer6_outputs(1085) <= not((layer5_outputs(1793)) xor (layer5_outputs(2461)));
    layer6_outputs(1086) <= '0';
    layer6_outputs(1087) <= not((layer5_outputs(2402)) xor (layer5_outputs(2425)));
    layer6_outputs(1088) <= (layer5_outputs(3087)) and not (layer5_outputs(4604));
    layer6_outputs(1089) <= (layer5_outputs(3978)) and not (layer5_outputs(3718));
    layer6_outputs(1090) <= not(layer5_outputs(515));
    layer6_outputs(1091) <= layer5_outputs(201);
    layer6_outputs(1092) <= (layer5_outputs(3403)) and not (layer5_outputs(1042));
    layer6_outputs(1093) <= not(layer5_outputs(1706));
    layer6_outputs(1094) <= layer5_outputs(304);
    layer6_outputs(1095) <= not((layer5_outputs(4684)) xor (layer5_outputs(1268)));
    layer6_outputs(1096) <= (layer5_outputs(1101)) xor (layer5_outputs(2050));
    layer6_outputs(1097) <= not(layer5_outputs(4679)) or (layer5_outputs(2160));
    layer6_outputs(1098) <= layer5_outputs(561);
    layer6_outputs(1099) <= layer5_outputs(3600);
    layer6_outputs(1100) <= not((layer5_outputs(4010)) and (layer5_outputs(1140)));
    layer6_outputs(1101) <= (layer5_outputs(3340)) and not (layer5_outputs(1164));
    layer6_outputs(1102) <= not(layer5_outputs(4206));
    layer6_outputs(1103) <= (layer5_outputs(4783)) xor (layer5_outputs(3698));
    layer6_outputs(1104) <= layer5_outputs(593);
    layer6_outputs(1105) <= layer5_outputs(2409);
    layer6_outputs(1106) <= (layer5_outputs(4309)) and (layer5_outputs(2689));
    layer6_outputs(1107) <= not((layer5_outputs(445)) xor (layer5_outputs(4800)));
    layer6_outputs(1108) <= not(layer5_outputs(4138));
    layer6_outputs(1109) <= not((layer5_outputs(897)) and (layer5_outputs(1375)));
    layer6_outputs(1110) <= (layer5_outputs(4375)) and (layer5_outputs(4969));
    layer6_outputs(1111) <= (layer5_outputs(2395)) or (layer5_outputs(212));
    layer6_outputs(1112) <= layer5_outputs(239);
    layer6_outputs(1113) <= not(layer5_outputs(2600));
    layer6_outputs(1114) <= not(layer5_outputs(1476));
    layer6_outputs(1115) <= (layer5_outputs(2310)) xor (layer5_outputs(3312));
    layer6_outputs(1116) <= '0';
    layer6_outputs(1117) <= layer5_outputs(2411);
    layer6_outputs(1118) <= layer5_outputs(4711);
    layer6_outputs(1119) <= (layer5_outputs(1461)) and not (layer5_outputs(1549));
    layer6_outputs(1120) <= layer5_outputs(2554);
    layer6_outputs(1121) <= layer5_outputs(4766);
    layer6_outputs(1122) <= (layer5_outputs(4594)) or (layer5_outputs(2889));
    layer6_outputs(1123) <= not(layer5_outputs(976));
    layer6_outputs(1124) <= layer5_outputs(1960);
    layer6_outputs(1125) <= (layer5_outputs(3334)) xor (layer5_outputs(106));
    layer6_outputs(1126) <= layer5_outputs(3709);
    layer6_outputs(1127) <= (layer5_outputs(364)) and not (layer5_outputs(530));
    layer6_outputs(1128) <= layer5_outputs(1773);
    layer6_outputs(1129) <= (layer5_outputs(1410)) or (layer5_outputs(3169));
    layer6_outputs(1130) <= not((layer5_outputs(157)) or (layer5_outputs(485)));
    layer6_outputs(1131) <= layer5_outputs(2107);
    layer6_outputs(1132) <= not(layer5_outputs(1696));
    layer6_outputs(1133) <= layer5_outputs(3440);
    layer6_outputs(1134) <= (layer5_outputs(2611)) and (layer5_outputs(2517));
    layer6_outputs(1135) <= not((layer5_outputs(2284)) and (layer5_outputs(256)));
    layer6_outputs(1136) <= layer5_outputs(720);
    layer6_outputs(1137) <= layer5_outputs(1812);
    layer6_outputs(1138) <= '1';
    layer6_outputs(1139) <= not(layer5_outputs(2299));
    layer6_outputs(1140) <= not(layer5_outputs(1251));
    layer6_outputs(1141) <= not(layer5_outputs(1424));
    layer6_outputs(1142) <= not(layer5_outputs(1974));
    layer6_outputs(1143) <= layer5_outputs(1612);
    layer6_outputs(1144) <= not(layer5_outputs(5107));
    layer6_outputs(1145) <= not(layer5_outputs(1581));
    layer6_outputs(1146) <= layer5_outputs(294);
    layer6_outputs(1147) <= layer5_outputs(3827);
    layer6_outputs(1148) <= layer5_outputs(2084);
    layer6_outputs(1149) <= not(layer5_outputs(1066));
    layer6_outputs(1150) <= layer5_outputs(3245);
    layer6_outputs(1151) <= (layer5_outputs(1677)) or (layer5_outputs(2854));
    layer6_outputs(1152) <= not(layer5_outputs(1633));
    layer6_outputs(1153) <= not((layer5_outputs(1667)) or (layer5_outputs(5112)));
    layer6_outputs(1154) <= layer5_outputs(1586);
    layer6_outputs(1155) <= (layer5_outputs(1861)) and not (layer5_outputs(473));
    layer6_outputs(1156) <= not((layer5_outputs(946)) xor (layer5_outputs(1853)));
    layer6_outputs(1157) <= not(layer5_outputs(2756));
    layer6_outputs(1158) <= not(layer5_outputs(638)) or (layer5_outputs(4986));
    layer6_outputs(1159) <= not(layer5_outputs(1516)) or (layer5_outputs(1791));
    layer6_outputs(1160) <= not(layer5_outputs(3695)) or (layer5_outputs(4854));
    layer6_outputs(1161) <= not((layer5_outputs(3535)) xor (layer5_outputs(2851)));
    layer6_outputs(1162) <= '1';
    layer6_outputs(1163) <= layer5_outputs(4915);
    layer6_outputs(1164) <= not((layer5_outputs(1639)) or (layer5_outputs(1555)));
    layer6_outputs(1165) <= layer5_outputs(2052);
    layer6_outputs(1166) <= not((layer5_outputs(3132)) or (layer5_outputs(4000)));
    layer6_outputs(1167) <= layer5_outputs(2064);
    layer6_outputs(1168) <= not((layer5_outputs(2087)) or (layer5_outputs(4825)));
    layer6_outputs(1169) <= not((layer5_outputs(3411)) and (layer5_outputs(4222)));
    layer6_outputs(1170) <= not(layer5_outputs(4351));
    layer6_outputs(1171) <= not((layer5_outputs(4581)) xor (layer5_outputs(2634)));
    layer6_outputs(1172) <= not(layer5_outputs(910)) or (layer5_outputs(2334));
    layer6_outputs(1173) <= not((layer5_outputs(5023)) xor (layer5_outputs(3918)));
    layer6_outputs(1174) <= (layer5_outputs(3420)) and not (layer5_outputs(5014));
    layer6_outputs(1175) <= (layer5_outputs(1905)) or (layer5_outputs(2422));
    layer6_outputs(1176) <= not(layer5_outputs(725));
    layer6_outputs(1177) <= (layer5_outputs(673)) xor (layer5_outputs(4009));
    layer6_outputs(1178) <= not(layer5_outputs(5060));
    layer6_outputs(1179) <= not(layer5_outputs(4266));
    layer6_outputs(1180) <= not(layer5_outputs(745));
    layer6_outputs(1181) <= not((layer5_outputs(1605)) and (layer5_outputs(3383)));
    layer6_outputs(1182) <= (layer5_outputs(2321)) or (layer5_outputs(648));
    layer6_outputs(1183) <= layer5_outputs(4482);
    layer6_outputs(1184) <= not(layer5_outputs(3519));
    layer6_outputs(1185) <= not(layer5_outputs(495));
    layer6_outputs(1186) <= (layer5_outputs(4445)) or (layer5_outputs(3772));
    layer6_outputs(1187) <= not(layer5_outputs(3844)) or (layer5_outputs(4199));
    layer6_outputs(1188) <= not((layer5_outputs(4950)) and (layer5_outputs(2315)));
    layer6_outputs(1189) <= not(layer5_outputs(567));
    layer6_outputs(1190) <= not(layer5_outputs(1515)) or (layer5_outputs(4116));
    layer6_outputs(1191) <= layer5_outputs(2137);
    layer6_outputs(1192) <= (layer5_outputs(3089)) or (layer5_outputs(2120));
    layer6_outputs(1193) <= not(layer5_outputs(1031));
    layer6_outputs(1194) <= layer5_outputs(2957);
    layer6_outputs(1195) <= not((layer5_outputs(1826)) or (layer5_outputs(751)));
    layer6_outputs(1196) <= layer5_outputs(475);
    layer6_outputs(1197) <= not(layer5_outputs(5001));
    layer6_outputs(1198) <= layer5_outputs(266);
    layer6_outputs(1199) <= (layer5_outputs(4755)) xor (layer5_outputs(1817));
    layer6_outputs(1200) <= not((layer5_outputs(239)) xor (layer5_outputs(2933)));
    layer6_outputs(1201) <= not((layer5_outputs(798)) xor (layer5_outputs(3383)));
    layer6_outputs(1202) <= not((layer5_outputs(3414)) xor (layer5_outputs(2497)));
    layer6_outputs(1203) <= layer5_outputs(4714);
    layer6_outputs(1204) <= not(layer5_outputs(2098)) or (layer5_outputs(4662));
    layer6_outputs(1205) <= not(layer5_outputs(3751));
    layer6_outputs(1206) <= not(layer5_outputs(3579));
    layer6_outputs(1207) <= layer5_outputs(1851);
    layer6_outputs(1208) <= layer5_outputs(342);
    layer6_outputs(1209) <= (layer5_outputs(2301)) or (layer5_outputs(1248));
    layer6_outputs(1210) <= (layer5_outputs(782)) and (layer5_outputs(2763));
    layer6_outputs(1211) <= layer5_outputs(3696);
    layer6_outputs(1212) <= layer5_outputs(1441);
    layer6_outputs(1213) <= not(layer5_outputs(985));
    layer6_outputs(1214) <= not(layer5_outputs(2998));
    layer6_outputs(1215) <= not((layer5_outputs(317)) xor (layer5_outputs(1447)));
    layer6_outputs(1216) <= not(layer5_outputs(4846)) or (layer5_outputs(3858));
    layer6_outputs(1217) <= layer5_outputs(3802);
    layer6_outputs(1218) <= layer5_outputs(570);
    layer6_outputs(1219) <= not(layer5_outputs(320));
    layer6_outputs(1220) <= (layer5_outputs(4648)) or (layer5_outputs(901));
    layer6_outputs(1221) <= layer5_outputs(3298);
    layer6_outputs(1222) <= not(layer5_outputs(1730));
    layer6_outputs(1223) <= not(layer5_outputs(838));
    layer6_outputs(1224) <= (layer5_outputs(4125)) xor (layer5_outputs(2578));
    layer6_outputs(1225) <= not(layer5_outputs(81)) or (layer5_outputs(2996));
    layer6_outputs(1226) <= layer5_outputs(4087);
    layer6_outputs(1227) <= not((layer5_outputs(4412)) or (layer5_outputs(3905)));
    layer6_outputs(1228) <= (layer5_outputs(4513)) xor (layer5_outputs(1457));
    layer6_outputs(1229) <= not((layer5_outputs(4842)) xor (layer5_outputs(3910)));
    layer6_outputs(1230) <= not(layer5_outputs(541));
    layer6_outputs(1231) <= (layer5_outputs(3727)) and not (layer5_outputs(186));
    layer6_outputs(1232) <= layer5_outputs(3421);
    layer6_outputs(1233) <= not((layer5_outputs(3149)) xor (layer5_outputs(2369)));
    layer6_outputs(1234) <= not((layer5_outputs(3945)) xor (layer5_outputs(16)));
    layer6_outputs(1235) <= (layer5_outputs(3617)) and not (layer5_outputs(4449));
    layer6_outputs(1236) <= layer5_outputs(4994);
    layer6_outputs(1237) <= (layer5_outputs(1928)) xor (layer5_outputs(3467));
    layer6_outputs(1238) <= layer5_outputs(3577);
    layer6_outputs(1239) <= not((layer5_outputs(3990)) xor (layer5_outputs(3273)));
    layer6_outputs(1240) <= not(layer5_outputs(296));
    layer6_outputs(1241) <= (layer5_outputs(1857)) and (layer5_outputs(3505));
    layer6_outputs(1242) <= not(layer5_outputs(1914));
    layer6_outputs(1243) <= not(layer5_outputs(4953));
    layer6_outputs(1244) <= (layer5_outputs(1480)) and not (layer5_outputs(2199));
    layer6_outputs(1245) <= not(layer5_outputs(2541));
    layer6_outputs(1246) <= (layer5_outputs(3635)) xor (layer5_outputs(2450));
    layer6_outputs(1247) <= not((layer5_outputs(579)) and (layer5_outputs(2433)));
    layer6_outputs(1248) <= layer5_outputs(2008);
    layer6_outputs(1249) <= (layer5_outputs(1428)) xor (layer5_outputs(1037));
    layer6_outputs(1250) <= '1';
    layer6_outputs(1251) <= not((layer5_outputs(4939)) xor (layer5_outputs(4287)));
    layer6_outputs(1252) <= layer5_outputs(11);
    layer6_outputs(1253) <= layer5_outputs(1311);
    layer6_outputs(1254) <= not((layer5_outputs(4993)) and (layer5_outputs(2323)));
    layer6_outputs(1255) <= not(layer5_outputs(940));
    layer6_outputs(1256) <= not(layer5_outputs(4437));
    layer6_outputs(1257) <= layer5_outputs(4481);
    layer6_outputs(1258) <= not(layer5_outputs(3220)) or (layer5_outputs(2731));
    layer6_outputs(1259) <= (layer5_outputs(2595)) xor (layer5_outputs(3712));
    layer6_outputs(1260) <= layer5_outputs(2124);
    layer6_outputs(1261) <= layer5_outputs(1785);
    layer6_outputs(1262) <= not(layer5_outputs(1833));
    layer6_outputs(1263) <= layer5_outputs(110);
    layer6_outputs(1264) <= (layer5_outputs(4937)) xor (layer5_outputs(3768));
    layer6_outputs(1265) <= layer5_outputs(968);
    layer6_outputs(1266) <= not((layer5_outputs(3513)) or (layer5_outputs(2854)));
    layer6_outputs(1267) <= layer5_outputs(202);
    layer6_outputs(1268) <= layer5_outputs(1901);
    layer6_outputs(1269) <= not((layer5_outputs(1050)) or (layer5_outputs(4162)));
    layer6_outputs(1270) <= layer5_outputs(1620);
    layer6_outputs(1271) <= layer5_outputs(4069);
    layer6_outputs(1272) <= (layer5_outputs(508)) or (layer5_outputs(1225));
    layer6_outputs(1273) <= not(layer5_outputs(2867)) or (layer5_outputs(687));
    layer6_outputs(1274) <= not((layer5_outputs(4272)) and (layer5_outputs(907)));
    layer6_outputs(1275) <= layer5_outputs(1085);
    layer6_outputs(1276) <= not(layer5_outputs(3909)) or (layer5_outputs(828));
    layer6_outputs(1277) <= layer5_outputs(3285);
    layer6_outputs(1278) <= layer5_outputs(839);
    layer6_outputs(1279) <= layer5_outputs(2686);
    layer6_outputs(1280) <= layer5_outputs(1460);
    layer6_outputs(1281) <= layer5_outputs(3756);
    layer6_outputs(1282) <= layer5_outputs(1558);
    layer6_outputs(1283) <= (layer5_outputs(2094)) and not (layer5_outputs(1599));
    layer6_outputs(1284) <= (layer5_outputs(5042)) and not (layer5_outputs(3443));
    layer6_outputs(1285) <= not((layer5_outputs(448)) xor (layer5_outputs(544)));
    layer6_outputs(1286) <= (layer5_outputs(1944)) and not (layer5_outputs(4844));
    layer6_outputs(1287) <= not(layer5_outputs(5041)) or (layer5_outputs(1922));
    layer6_outputs(1288) <= not(layer5_outputs(2700));
    layer6_outputs(1289) <= not((layer5_outputs(731)) or (layer5_outputs(896)));
    layer6_outputs(1290) <= not(layer5_outputs(3100));
    layer6_outputs(1291) <= layer5_outputs(4183);
    layer6_outputs(1292) <= '1';
    layer6_outputs(1293) <= not(layer5_outputs(564));
    layer6_outputs(1294) <= not(layer5_outputs(3388));
    layer6_outputs(1295) <= layer5_outputs(1869);
    layer6_outputs(1296) <= (layer5_outputs(2991)) xor (layer5_outputs(1603));
    layer6_outputs(1297) <= layer5_outputs(4779);
    layer6_outputs(1298) <= not(layer5_outputs(2601));
    layer6_outputs(1299) <= layer5_outputs(3963);
    layer6_outputs(1300) <= (layer5_outputs(1136)) or (layer5_outputs(4554));
    layer6_outputs(1301) <= (layer5_outputs(1549)) or (layer5_outputs(83));
    layer6_outputs(1302) <= layer5_outputs(2820);
    layer6_outputs(1303) <= (layer5_outputs(819)) xor (layer5_outputs(3791));
    layer6_outputs(1304) <= layer5_outputs(3682);
    layer6_outputs(1305) <= not(layer5_outputs(1845));
    layer6_outputs(1306) <= (layer5_outputs(3135)) and not (layer5_outputs(2418));
    layer6_outputs(1307) <= not(layer5_outputs(2766));
    layer6_outputs(1308) <= layer5_outputs(3946);
    layer6_outputs(1309) <= not(layer5_outputs(2276));
    layer6_outputs(1310) <= not((layer5_outputs(658)) and (layer5_outputs(3944)));
    layer6_outputs(1311) <= layer5_outputs(4650);
    layer6_outputs(1312) <= layer5_outputs(3466);
    layer6_outputs(1313) <= not(layer5_outputs(4530));
    layer6_outputs(1314) <= not((layer5_outputs(4887)) and (layer5_outputs(4234)));
    layer6_outputs(1315) <= layer5_outputs(381);
    layer6_outputs(1316) <= not((layer5_outputs(4162)) xor (layer5_outputs(860)));
    layer6_outputs(1317) <= layer5_outputs(3024);
    layer6_outputs(1318) <= not(layer5_outputs(666));
    layer6_outputs(1319) <= not(layer5_outputs(4662)) or (layer5_outputs(2599));
    layer6_outputs(1320) <= not((layer5_outputs(4139)) xor (layer5_outputs(1954)));
    layer6_outputs(1321) <= not(layer5_outputs(1598));
    layer6_outputs(1322) <= not(layer5_outputs(4343));
    layer6_outputs(1323) <= not(layer5_outputs(1613)) or (layer5_outputs(1871));
    layer6_outputs(1324) <= (layer5_outputs(3893)) xor (layer5_outputs(2941));
    layer6_outputs(1325) <= layer5_outputs(2354);
    layer6_outputs(1326) <= not(layer5_outputs(1930));
    layer6_outputs(1327) <= (layer5_outputs(2264)) or (layer5_outputs(3134));
    layer6_outputs(1328) <= not(layer5_outputs(2606)) or (layer5_outputs(1661));
    layer6_outputs(1329) <= layer5_outputs(1910);
    layer6_outputs(1330) <= (layer5_outputs(4957)) and (layer5_outputs(4726));
    layer6_outputs(1331) <= not(layer5_outputs(4775)) or (layer5_outputs(2216));
    layer6_outputs(1332) <= layer5_outputs(4044);
    layer6_outputs(1333) <= not(layer5_outputs(4705));
    layer6_outputs(1334) <= not(layer5_outputs(1384)) or (layer5_outputs(3841));
    layer6_outputs(1335) <= not(layer5_outputs(3975)) or (layer5_outputs(3190));
    layer6_outputs(1336) <= not((layer5_outputs(3188)) xor (layer5_outputs(4661)));
    layer6_outputs(1337) <= layer5_outputs(1806);
    layer6_outputs(1338) <= not(layer5_outputs(676));
    layer6_outputs(1339) <= not(layer5_outputs(994));
    layer6_outputs(1340) <= layer5_outputs(2803);
    layer6_outputs(1341) <= not((layer5_outputs(3750)) xor (layer5_outputs(4275)));
    layer6_outputs(1342) <= (layer5_outputs(4457)) xor (layer5_outputs(4245));
    layer6_outputs(1343) <= layer5_outputs(3275);
    layer6_outputs(1344) <= not((layer5_outputs(2276)) xor (layer5_outputs(4769)));
    layer6_outputs(1345) <= (layer5_outputs(2960)) xor (layer5_outputs(2645));
    layer6_outputs(1346) <= '0';
    layer6_outputs(1347) <= layer5_outputs(1199);
    layer6_outputs(1348) <= not((layer5_outputs(2195)) xor (layer5_outputs(3807)));
    layer6_outputs(1349) <= not(layer5_outputs(2260));
    layer6_outputs(1350) <= not(layer5_outputs(2270));
    layer6_outputs(1351) <= layer5_outputs(881);
    layer6_outputs(1352) <= not(layer5_outputs(3495));
    layer6_outputs(1353) <= (layer5_outputs(200)) or (layer5_outputs(2955));
    layer6_outputs(1354) <= not(layer5_outputs(4333));
    layer6_outputs(1355) <= not(layer5_outputs(4761)) or (layer5_outputs(4680));
    layer6_outputs(1356) <= not((layer5_outputs(936)) and (layer5_outputs(428)));
    layer6_outputs(1357) <= (layer5_outputs(939)) xor (layer5_outputs(4439));
    layer6_outputs(1358) <= not(layer5_outputs(5111));
    layer6_outputs(1359) <= not((layer5_outputs(532)) xor (layer5_outputs(4601)));
    layer6_outputs(1360) <= (layer5_outputs(5082)) and not (layer5_outputs(3791));
    layer6_outputs(1361) <= not(layer5_outputs(3262));
    layer6_outputs(1362) <= (layer5_outputs(4945)) and not (layer5_outputs(2695));
    layer6_outputs(1363) <= not(layer5_outputs(3111));
    layer6_outputs(1364) <= not(layer5_outputs(1421)) or (layer5_outputs(2457));
    layer6_outputs(1365) <= not(layer5_outputs(1413));
    layer6_outputs(1366) <= not(layer5_outputs(2115));
    layer6_outputs(1367) <= (layer5_outputs(4429)) xor (layer5_outputs(5075));
    layer6_outputs(1368) <= layer5_outputs(2366);
    layer6_outputs(1369) <= not((layer5_outputs(2244)) and (layer5_outputs(1921)));
    layer6_outputs(1370) <= not((layer5_outputs(3133)) xor (layer5_outputs(2371)));
    layer6_outputs(1371) <= not(layer5_outputs(2231)) or (layer5_outputs(2788));
    layer6_outputs(1372) <= (layer5_outputs(656)) xor (layer5_outputs(1370));
    layer6_outputs(1373) <= not(layer5_outputs(5077));
    layer6_outputs(1374) <= layer5_outputs(3934);
    layer6_outputs(1375) <= (layer5_outputs(2271)) and (layer5_outputs(3426));
    layer6_outputs(1376) <= (layer5_outputs(471)) or (layer5_outputs(1023));
    layer6_outputs(1377) <= not(layer5_outputs(319));
    layer6_outputs(1378) <= not(layer5_outputs(781));
    layer6_outputs(1379) <= layer5_outputs(3097);
    layer6_outputs(1380) <= (layer5_outputs(3163)) or (layer5_outputs(286));
    layer6_outputs(1381) <= (layer5_outputs(3174)) or (layer5_outputs(1083));
    layer6_outputs(1382) <= not(layer5_outputs(4659));
    layer6_outputs(1383) <= layer5_outputs(1301);
    layer6_outputs(1384) <= (layer5_outputs(5069)) and not (layer5_outputs(3124));
    layer6_outputs(1385) <= not(layer5_outputs(2413));
    layer6_outputs(1386) <= layer5_outputs(343);
    layer6_outputs(1387) <= (layer5_outputs(584)) and (layer5_outputs(5015));
    layer6_outputs(1388) <= layer5_outputs(1823);
    layer6_outputs(1389) <= (layer5_outputs(3942)) and not (layer5_outputs(2918));
    layer6_outputs(1390) <= not(layer5_outputs(5003));
    layer6_outputs(1391) <= not(layer5_outputs(3001));
    layer6_outputs(1392) <= not(layer5_outputs(3511));
    layer6_outputs(1393) <= not(layer5_outputs(1206));
    layer6_outputs(1394) <= (layer5_outputs(3184)) xor (layer5_outputs(2661));
    layer6_outputs(1395) <= not((layer5_outputs(3979)) xor (layer5_outputs(2665)));
    layer6_outputs(1396) <= layer5_outputs(4261);
    layer6_outputs(1397) <= not((layer5_outputs(2784)) xor (layer5_outputs(4153)));
    layer6_outputs(1398) <= layer5_outputs(2217);
    layer6_outputs(1399) <= not(layer5_outputs(3982)) or (layer5_outputs(2289));
    layer6_outputs(1400) <= not(layer5_outputs(880));
    layer6_outputs(1401) <= layer5_outputs(2693);
    layer6_outputs(1402) <= not((layer5_outputs(2429)) xor (layer5_outputs(1601)));
    layer6_outputs(1403) <= '0';
    layer6_outputs(1404) <= not((layer5_outputs(2779)) and (layer5_outputs(37)));
    layer6_outputs(1405) <= (layer5_outputs(430)) xor (layer5_outputs(3070));
    layer6_outputs(1406) <= not(layer5_outputs(4053));
    layer6_outputs(1407) <= layer5_outputs(3551);
    layer6_outputs(1408) <= (layer5_outputs(1953)) and not (layer5_outputs(940));
    layer6_outputs(1409) <= not(layer5_outputs(836)) or (layer5_outputs(1390));
    layer6_outputs(1410) <= not(layer5_outputs(2062));
    layer6_outputs(1411) <= not(layer5_outputs(1551));
    layer6_outputs(1412) <= (layer5_outputs(652)) and not (layer5_outputs(1350));
    layer6_outputs(1413) <= not((layer5_outputs(269)) or (layer5_outputs(1252)));
    layer6_outputs(1414) <= (layer5_outputs(2956)) and not (layer5_outputs(3033));
    layer6_outputs(1415) <= not((layer5_outputs(1212)) and (layer5_outputs(4391)));
    layer6_outputs(1416) <= (layer5_outputs(2384)) or (layer5_outputs(5073));
    layer6_outputs(1417) <= (layer5_outputs(2075)) and not (layer5_outputs(4988));
    layer6_outputs(1418) <= (layer5_outputs(3318)) and (layer5_outputs(4110));
    layer6_outputs(1419) <= layer5_outputs(3415);
    layer6_outputs(1420) <= (layer5_outputs(4018)) xor (layer5_outputs(694));
    layer6_outputs(1421) <= not((layer5_outputs(4707)) xor (layer5_outputs(142)));
    layer6_outputs(1422) <= not(layer5_outputs(267));
    layer6_outputs(1423) <= not(layer5_outputs(3665));
    layer6_outputs(1424) <= not(layer5_outputs(3010));
    layer6_outputs(1425) <= layer5_outputs(4592);
    layer6_outputs(1426) <= '0';
    layer6_outputs(1427) <= (layer5_outputs(2526)) or (layer5_outputs(425));
    layer6_outputs(1428) <= (layer5_outputs(4503)) and not (layer5_outputs(1209));
    layer6_outputs(1429) <= (layer5_outputs(4407)) or (layer5_outputs(1678));
    layer6_outputs(1430) <= not(layer5_outputs(4246)) or (layer5_outputs(1075));
    layer6_outputs(1431) <= layer5_outputs(4695);
    layer6_outputs(1432) <= not(layer5_outputs(1366));
    layer6_outputs(1433) <= not((layer5_outputs(4066)) xor (layer5_outputs(2471)));
    layer6_outputs(1434) <= (layer5_outputs(4104)) and not (layer5_outputs(3520));
    layer6_outputs(1435) <= not(layer5_outputs(1241));
    layer6_outputs(1436) <= not((layer5_outputs(5051)) xor (layer5_outputs(1087)));
    layer6_outputs(1437) <= (layer5_outputs(1383)) xor (layer5_outputs(3561));
    layer6_outputs(1438) <= layer5_outputs(496);
    layer6_outputs(1439) <= layer5_outputs(1495);
    layer6_outputs(1440) <= not(layer5_outputs(1572));
    layer6_outputs(1441) <= '1';
    layer6_outputs(1442) <= layer5_outputs(2628);
    layer6_outputs(1443) <= not(layer5_outputs(1644));
    layer6_outputs(1444) <= not(layer5_outputs(175)) or (layer5_outputs(2807));
    layer6_outputs(1445) <= '0';
    layer6_outputs(1446) <= layer5_outputs(1201);
    layer6_outputs(1447) <= layer5_outputs(1414);
    layer6_outputs(1448) <= not(layer5_outputs(945)) or (layer5_outputs(1170));
    layer6_outputs(1449) <= not(layer5_outputs(990)) or (layer5_outputs(2350));
    layer6_outputs(1450) <= (layer5_outputs(3912)) and not (layer5_outputs(3538));
    layer6_outputs(1451) <= not(layer5_outputs(1770));
    layer6_outputs(1452) <= layer5_outputs(228);
    layer6_outputs(1453) <= not(layer5_outputs(3946));
    layer6_outputs(1454) <= not(layer5_outputs(1049));
    layer6_outputs(1455) <= not(layer5_outputs(2113)) or (layer5_outputs(4324));
    layer6_outputs(1456) <= not(layer5_outputs(696));
    layer6_outputs(1457) <= layer5_outputs(2574);
    layer6_outputs(1458) <= not((layer5_outputs(1311)) xor (layer5_outputs(335)));
    layer6_outputs(1459) <= layer5_outputs(5053);
    layer6_outputs(1460) <= '0';
    layer6_outputs(1461) <= layer5_outputs(1970);
    layer6_outputs(1462) <= not((layer5_outputs(982)) or (layer5_outputs(4267)));
    layer6_outputs(1463) <= not(layer5_outputs(4496));
    layer6_outputs(1464) <= not(layer5_outputs(1385));
    layer6_outputs(1465) <= not(layer5_outputs(3777)) or (layer5_outputs(1498));
    layer6_outputs(1466) <= not(layer5_outputs(4895));
    layer6_outputs(1467) <= layer5_outputs(1409);
    layer6_outputs(1468) <= not(layer5_outputs(3933));
    layer6_outputs(1469) <= not(layer5_outputs(1485));
    layer6_outputs(1470) <= not(layer5_outputs(3461)) or (layer5_outputs(2706));
    layer6_outputs(1471) <= layer5_outputs(558);
    layer6_outputs(1472) <= (layer5_outputs(3293)) and (layer5_outputs(2037));
    layer6_outputs(1473) <= (layer5_outputs(2844)) and (layer5_outputs(4122));
    layer6_outputs(1474) <= not(layer5_outputs(4803)) or (layer5_outputs(4655));
    layer6_outputs(1475) <= layer5_outputs(4941);
    layer6_outputs(1476) <= not(layer5_outputs(2694));
    layer6_outputs(1477) <= (layer5_outputs(1352)) and (layer5_outputs(646));
    layer6_outputs(1478) <= (layer5_outputs(3068)) xor (layer5_outputs(3651));
    layer6_outputs(1479) <= '1';
    layer6_outputs(1480) <= (layer5_outputs(4996)) xor (layer5_outputs(787));
    layer6_outputs(1481) <= layer5_outputs(1867);
    layer6_outputs(1482) <= not(layer5_outputs(3981));
    layer6_outputs(1483) <= not(layer5_outputs(4053));
    layer6_outputs(1484) <= layer5_outputs(5052);
    layer6_outputs(1485) <= layer5_outputs(4389);
    layer6_outputs(1486) <= (layer5_outputs(2859)) and (layer5_outputs(2012));
    layer6_outputs(1487) <= layer5_outputs(3053);
    layer6_outputs(1488) <= layer5_outputs(5034);
    layer6_outputs(1489) <= (layer5_outputs(376)) and (layer5_outputs(3976));
    layer6_outputs(1490) <= not((layer5_outputs(904)) xor (layer5_outputs(334)));
    layer6_outputs(1491) <= '1';
    layer6_outputs(1492) <= layer5_outputs(4632);
    layer6_outputs(1493) <= not(layer5_outputs(115)) or (layer5_outputs(4058));
    layer6_outputs(1494) <= layer5_outputs(612);
    layer6_outputs(1495) <= layer5_outputs(3482);
    layer6_outputs(1496) <= layer5_outputs(3036);
    layer6_outputs(1497) <= not((layer5_outputs(3232)) or (layer5_outputs(3307)));
    layer6_outputs(1498) <= layer5_outputs(1908);
    layer6_outputs(1499) <= (layer5_outputs(3759)) and (layer5_outputs(4657));
    layer6_outputs(1500) <= not(layer5_outputs(3737));
    layer6_outputs(1501) <= (layer5_outputs(5079)) and not (layer5_outputs(3971));
    layer6_outputs(1502) <= not(layer5_outputs(3114));
    layer6_outputs(1503) <= not(layer5_outputs(668)) or (layer5_outputs(4505));
    layer6_outputs(1504) <= not(layer5_outputs(1683));
    layer6_outputs(1505) <= (layer5_outputs(2891)) xor (layer5_outputs(1008));
    layer6_outputs(1506) <= layer5_outputs(4250);
    layer6_outputs(1507) <= layer5_outputs(3997);
    layer6_outputs(1508) <= not((layer5_outputs(2355)) and (layer5_outputs(4877)));
    layer6_outputs(1509) <= not((layer5_outputs(1797)) and (layer5_outputs(674)));
    layer6_outputs(1510) <= not(layer5_outputs(2984));
    layer6_outputs(1511) <= (layer5_outputs(4010)) or (layer5_outputs(561));
    layer6_outputs(1512) <= not(layer5_outputs(3479));
    layer6_outputs(1513) <= not(layer5_outputs(2711));
    layer6_outputs(1514) <= layer5_outputs(270);
    layer6_outputs(1515) <= (layer5_outputs(890)) and not (layer5_outputs(734));
    layer6_outputs(1516) <= (layer5_outputs(3297)) and (layer5_outputs(4178));
    layer6_outputs(1517) <= (layer5_outputs(3530)) and not (layer5_outputs(4621));
    layer6_outputs(1518) <= (layer5_outputs(3278)) xor (layer5_outputs(4370));
    layer6_outputs(1519) <= not(layer5_outputs(3313));
    layer6_outputs(1520) <= not(layer5_outputs(2823));
    layer6_outputs(1521) <= layer5_outputs(1558);
    layer6_outputs(1522) <= layer5_outputs(533);
    layer6_outputs(1523) <= not((layer5_outputs(2316)) or (layer5_outputs(669)));
    layer6_outputs(1524) <= not(layer5_outputs(3059));
    layer6_outputs(1525) <= layer5_outputs(3119);
    layer6_outputs(1526) <= not(layer5_outputs(3831));
    layer6_outputs(1527) <= layer5_outputs(2619);
    layer6_outputs(1528) <= not(layer5_outputs(2296));
    layer6_outputs(1529) <= not(layer5_outputs(190));
    layer6_outputs(1530) <= (layer5_outputs(893)) xor (layer5_outputs(246));
    layer6_outputs(1531) <= not(layer5_outputs(1277));
    layer6_outputs(1532) <= (layer5_outputs(3190)) xor (layer5_outputs(5006));
    layer6_outputs(1533) <= layer5_outputs(543);
    layer6_outputs(1534) <= (layer5_outputs(4374)) and (layer5_outputs(3553));
    layer6_outputs(1535) <= not(layer5_outputs(4300)) or (layer5_outputs(2376));
    layer6_outputs(1536) <= not(layer5_outputs(4602));
    layer6_outputs(1537) <= not(layer5_outputs(1654));
    layer6_outputs(1538) <= not((layer5_outputs(143)) and (layer5_outputs(3254)));
    layer6_outputs(1539) <= not(layer5_outputs(281));
    layer6_outputs(1540) <= not(layer5_outputs(3386));
    layer6_outputs(1541) <= not(layer5_outputs(2402));
    layer6_outputs(1542) <= (layer5_outputs(2662)) and not (layer5_outputs(2585));
    layer6_outputs(1543) <= layer5_outputs(4987);
    layer6_outputs(1544) <= layer5_outputs(3463);
    layer6_outputs(1545) <= layer5_outputs(1210);
    layer6_outputs(1546) <= (layer5_outputs(227)) and not (layer5_outputs(1855));
    layer6_outputs(1547) <= not(layer5_outputs(1926)) or (layer5_outputs(1403));
    layer6_outputs(1548) <= not((layer5_outputs(3317)) xor (layer5_outputs(1547)));
    layer6_outputs(1549) <= not(layer5_outputs(4347)) or (layer5_outputs(634));
    layer6_outputs(1550) <= not(layer5_outputs(2790));
    layer6_outputs(1551) <= (layer5_outputs(4687)) or (layer5_outputs(3401));
    layer6_outputs(1552) <= layer5_outputs(50);
    layer6_outputs(1553) <= (layer5_outputs(4698)) and (layer5_outputs(4930));
    layer6_outputs(1554) <= not(layer5_outputs(4613)) or (layer5_outputs(2597));
    layer6_outputs(1555) <= not((layer5_outputs(3636)) or (layer5_outputs(3277)));
    layer6_outputs(1556) <= not((layer5_outputs(909)) xor (layer5_outputs(631)));
    layer6_outputs(1557) <= not((layer5_outputs(3702)) xor (layer5_outputs(415)));
    layer6_outputs(1558) <= layer5_outputs(1174);
    layer6_outputs(1559) <= not(layer5_outputs(2817));
    layer6_outputs(1560) <= layer5_outputs(3863);
    layer6_outputs(1561) <= not((layer5_outputs(2145)) and (layer5_outputs(3536)));
    layer6_outputs(1562) <= layer5_outputs(2394);
    layer6_outputs(1563) <= layer5_outputs(4290);
    layer6_outputs(1564) <= not((layer5_outputs(4387)) and (layer5_outputs(2138)));
    layer6_outputs(1565) <= (layer5_outputs(4365)) xor (layer5_outputs(1119));
    layer6_outputs(1566) <= not(layer5_outputs(991)) or (layer5_outputs(2924));
    layer6_outputs(1567) <= not((layer5_outputs(3957)) xor (layer5_outputs(4874)));
    layer6_outputs(1568) <= (layer5_outputs(81)) and not (layer5_outputs(3447));
    layer6_outputs(1569) <= not((layer5_outputs(173)) xor (layer5_outputs(3231)));
    layer6_outputs(1570) <= (layer5_outputs(4239)) and (layer5_outputs(2340));
    layer6_outputs(1571) <= not(layer5_outputs(4811)) or (layer5_outputs(2226));
    layer6_outputs(1572) <= not(layer5_outputs(4977));
    layer6_outputs(1573) <= (layer5_outputs(1186)) and not (layer5_outputs(4624));
    layer6_outputs(1574) <= not(layer5_outputs(2792));
    layer6_outputs(1575) <= not(layer5_outputs(3381));
    layer6_outputs(1576) <= not((layer5_outputs(4792)) xor (layer5_outputs(4672)));
    layer6_outputs(1577) <= layer5_outputs(4351);
    layer6_outputs(1578) <= not((layer5_outputs(714)) xor (layer5_outputs(4040)));
    layer6_outputs(1579) <= not(layer5_outputs(3040));
    layer6_outputs(1580) <= not(layer5_outputs(1392));
    layer6_outputs(1581) <= not((layer5_outputs(2262)) xor (layer5_outputs(2221)));
    layer6_outputs(1582) <= (layer5_outputs(120)) xor (layer5_outputs(638));
    layer6_outputs(1583) <= layer5_outputs(2909);
    layer6_outputs(1584) <= not((layer5_outputs(4770)) xor (layer5_outputs(2958)));
    layer6_outputs(1585) <= not((layer5_outputs(665)) xor (layer5_outputs(1569)));
    layer6_outputs(1586) <= layer5_outputs(511);
    layer6_outputs(1587) <= not(layer5_outputs(1111));
    layer6_outputs(1588) <= (layer5_outputs(548)) and not (layer5_outputs(67));
    layer6_outputs(1589) <= (layer5_outputs(2056)) xor (layer5_outputs(1658));
    layer6_outputs(1590) <= layer5_outputs(3510);
    layer6_outputs(1591) <= not(layer5_outputs(1930));
    layer6_outputs(1592) <= not(layer5_outputs(2965));
    layer6_outputs(1593) <= '0';
    layer6_outputs(1594) <= not((layer5_outputs(1530)) and (layer5_outputs(4956)));
    layer6_outputs(1595) <= not(layer5_outputs(4625));
    layer6_outputs(1596) <= not((layer5_outputs(1583)) xor (layer5_outputs(1896)));
    layer6_outputs(1597) <= not(layer5_outputs(601));
    layer6_outputs(1598) <= not(layer5_outputs(1735)) or (layer5_outputs(2536));
    layer6_outputs(1599) <= (layer5_outputs(4212)) and (layer5_outputs(3741));
    layer6_outputs(1600) <= not((layer5_outputs(4467)) xor (layer5_outputs(3569)));
    layer6_outputs(1601) <= layer5_outputs(1681);
    layer6_outputs(1602) <= not(layer5_outputs(1789));
    layer6_outputs(1603) <= not(layer5_outputs(3526)) or (layer5_outputs(2139));
    layer6_outputs(1604) <= layer5_outputs(1395);
    layer6_outputs(1605) <= not(layer5_outputs(3022)) or (layer5_outputs(4131));
    layer6_outputs(1606) <= not((layer5_outputs(1701)) and (layer5_outputs(2351)));
    layer6_outputs(1607) <= layer5_outputs(3737);
    layer6_outputs(1608) <= not((layer5_outputs(3951)) xor (layer5_outputs(2335)));
    layer6_outputs(1609) <= not((layer5_outputs(3050)) xor (layer5_outputs(628)));
    layer6_outputs(1610) <= layer5_outputs(3861);
    layer6_outputs(1611) <= not(layer5_outputs(547));
    layer6_outputs(1612) <= not(layer5_outputs(4912));
    layer6_outputs(1613) <= not(layer5_outputs(1345));
    layer6_outputs(1614) <= (layer5_outputs(4427)) and (layer5_outputs(2639));
    layer6_outputs(1615) <= not((layer5_outputs(3166)) or (layer5_outputs(4834)));
    layer6_outputs(1616) <= not(layer5_outputs(137));
    layer6_outputs(1617) <= not((layer5_outputs(1875)) or (layer5_outputs(4383)));
    layer6_outputs(1618) <= not(layer5_outputs(1261));
    layer6_outputs(1619) <= not(layer5_outputs(2176));
    layer6_outputs(1620) <= not(layer5_outputs(3229));
    layer6_outputs(1621) <= not(layer5_outputs(2820));
    layer6_outputs(1622) <= (layer5_outputs(2403)) and not (layer5_outputs(218));
    layer6_outputs(1623) <= layer5_outputs(2047);
    layer6_outputs(1624) <= not(layer5_outputs(3860));
    layer6_outputs(1625) <= (layer5_outputs(262)) xor (layer5_outputs(3964));
    layer6_outputs(1626) <= (layer5_outputs(280)) xor (layer5_outputs(1462));
    layer6_outputs(1627) <= layer5_outputs(4224);
    layer6_outputs(1628) <= layer5_outputs(514);
    layer6_outputs(1629) <= layer5_outputs(4731);
    layer6_outputs(1630) <= not(layer5_outputs(4349));
    layer6_outputs(1631) <= (layer5_outputs(2034)) or (layer5_outputs(539));
    layer6_outputs(1632) <= not(layer5_outputs(1016)) or (layer5_outputs(2251));
    layer6_outputs(1633) <= layer5_outputs(754);
    layer6_outputs(1634) <= not(layer5_outputs(711));
    layer6_outputs(1635) <= (layer5_outputs(2659)) or (layer5_outputs(4061));
    layer6_outputs(1636) <= not((layer5_outputs(1535)) and (layer5_outputs(391)));
    layer6_outputs(1637) <= not(layer5_outputs(2757));
    layer6_outputs(1638) <= layer5_outputs(1045);
    layer6_outputs(1639) <= layer5_outputs(2696);
    layer6_outputs(1640) <= not((layer5_outputs(3925)) xor (layer5_outputs(2357)));
    layer6_outputs(1641) <= (layer5_outputs(558)) and not (layer5_outputs(493));
    layer6_outputs(1642) <= (layer5_outputs(1957)) xor (layer5_outputs(3410));
    layer6_outputs(1643) <= not(layer5_outputs(1985));
    layer6_outputs(1644) <= not((layer5_outputs(847)) and (layer5_outputs(334)));
    layer6_outputs(1645) <= layer5_outputs(363);
    layer6_outputs(1646) <= not(layer5_outputs(31));
    layer6_outputs(1647) <= layer5_outputs(5040);
    layer6_outputs(1648) <= not(layer5_outputs(648));
    layer6_outputs(1649) <= layer5_outputs(3123);
    layer6_outputs(1650) <= not((layer5_outputs(2974)) or (layer5_outputs(3632)));
    layer6_outputs(1651) <= not(layer5_outputs(2621));
    layer6_outputs(1652) <= layer5_outputs(1432);
    layer6_outputs(1653) <= not(layer5_outputs(869));
    layer6_outputs(1654) <= layer5_outputs(192);
    layer6_outputs(1655) <= not(layer5_outputs(2600));
    layer6_outputs(1656) <= not((layer5_outputs(1775)) xor (layer5_outputs(277)));
    layer6_outputs(1657) <= not(layer5_outputs(1512));
    layer6_outputs(1658) <= not(layer5_outputs(3366)) or (layer5_outputs(1188));
    layer6_outputs(1659) <= not(layer5_outputs(1071));
    layer6_outputs(1660) <= not(layer5_outputs(2779));
    layer6_outputs(1661) <= not(layer5_outputs(1482)) or (layer5_outputs(730));
    layer6_outputs(1662) <= not(layer5_outputs(4547)) or (layer5_outputs(2124));
    layer6_outputs(1663) <= not(layer5_outputs(4326));
    layer6_outputs(1664) <= layer5_outputs(2086);
    layer6_outputs(1665) <= (layer5_outputs(4574)) and (layer5_outputs(2567));
    layer6_outputs(1666) <= layer5_outputs(961);
    layer6_outputs(1667) <= layer5_outputs(3647);
    layer6_outputs(1668) <= (layer5_outputs(3207)) xor (layer5_outputs(4387));
    layer6_outputs(1669) <= (layer5_outputs(2304)) and not (layer5_outputs(465));
    layer6_outputs(1670) <= layer5_outputs(21);
    layer6_outputs(1671) <= (layer5_outputs(2414)) xor (layer5_outputs(1729));
    layer6_outputs(1672) <= not((layer5_outputs(2471)) and (layer5_outputs(4683)));
    layer6_outputs(1673) <= layer5_outputs(3944);
    layer6_outputs(1674) <= (layer5_outputs(114)) and not (layer5_outputs(3619));
    layer6_outputs(1675) <= not(layer5_outputs(649));
    layer6_outputs(1676) <= (layer5_outputs(2007)) and (layer5_outputs(3689));
    layer6_outputs(1677) <= not(layer5_outputs(1979));
    layer6_outputs(1678) <= (layer5_outputs(3697)) and not (layer5_outputs(4430));
    layer6_outputs(1679) <= (layer5_outputs(2538)) xor (layer5_outputs(574));
    layer6_outputs(1680) <= (layer5_outputs(1487)) xor (layer5_outputs(2435));
    layer6_outputs(1681) <= layer5_outputs(1867);
    layer6_outputs(1682) <= layer5_outputs(255);
    layer6_outputs(1683) <= not(layer5_outputs(808));
    layer6_outputs(1684) <= layer5_outputs(2778);
    layer6_outputs(1685) <= layer5_outputs(4413);
    layer6_outputs(1686) <= layer5_outputs(2424);
    layer6_outputs(1687) <= not(layer5_outputs(272));
    layer6_outputs(1688) <= not(layer5_outputs(3177));
    layer6_outputs(1689) <= not(layer5_outputs(1939));
    layer6_outputs(1690) <= not(layer5_outputs(562)) or (layer5_outputs(1641));
    layer6_outputs(1691) <= layer5_outputs(2132);
    layer6_outputs(1692) <= not(layer5_outputs(1759));
    layer6_outputs(1693) <= layer5_outputs(4879);
    layer6_outputs(1694) <= layer5_outputs(3271);
    layer6_outputs(1695) <= (layer5_outputs(2194)) and not (layer5_outputs(4747));
    layer6_outputs(1696) <= layer5_outputs(300);
    layer6_outputs(1697) <= not(layer5_outputs(1011));
    layer6_outputs(1698) <= not(layer5_outputs(2673));
    layer6_outputs(1699) <= layer5_outputs(4039);
    layer6_outputs(1700) <= not(layer5_outputs(4470));
    layer6_outputs(1701) <= not(layer5_outputs(2515));
    layer6_outputs(1702) <= (layer5_outputs(830)) or (layer5_outputs(1986));
    layer6_outputs(1703) <= '0';
    layer6_outputs(1704) <= (layer5_outputs(1213)) and (layer5_outputs(2584));
    layer6_outputs(1705) <= layer5_outputs(4850);
    layer6_outputs(1706) <= (layer5_outputs(1938)) xor (layer5_outputs(4259));
    layer6_outputs(1707) <= not((layer5_outputs(2162)) xor (layer5_outputs(4854)));
    layer6_outputs(1708) <= (layer5_outputs(2062)) and not (layer5_outputs(1751));
    layer6_outputs(1709) <= not(layer5_outputs(27));
    layer6_outputs(1710) <= not(layer5_outputs(2594));
    layer6_outputs(1711) <= (layer5_outputs(362)) or (layer5_outputs(109));
    layer6_outputs(1712) <= (layer5_outputs(2588)) and not (layer5_outputs(3741));
    layer6_outputs(1713) <= not(layer5_outputs(1013)) or (layer5_outputs(3603));
    layer6_outputs(1714) <= not(layer5_outputs(237));
    layer6_outputs(1715) <= layer5_outputs(3887);
    layer6_outputs(1716) <= not((layer5_outputs(1242)) or (layer5_outputs(1912)));
    layer6_outputs(1717) <= not(layer5_outputs(1396));
    layer6_outputs(1718) <= not(layer5_outputs(3832));
    layer6_outputs(1719) <= not(layer5_outputs(71));
    layer6_outputs(1720) <= layer5_outputs(3188);
    layer6_outputs(1721) <= '0';
    layer6_outputs(1722) <= not(layer5_outputs(4031)) or (layer5_outputs(4374));
    layer6_outputs(1723) <= not(layer5_outputs(1298));
    layer6_outputs(1724) <= (layer5_outputs(4062)) and not (layer5_outputs(534));
    layer6_outputs(1725) <= layer5_outputs(568);
    layer6_outputs(1726) <= layer5_outputs(499);
    layer6_outputs(1727) <= layer5_outputs(3794);
    layer6_outputs(1728) <= (layer5_outputs(199)) xor (layer5_outputs(3158));
    layer6_outputs(1729) <= layer5_outputs(4001);
    layer6_outputs(1730) <= (layer5_outputs(687)) and not (layer5_outputs(3705));
    layer6_outputs(1731) <= not(layer5_outputs(397));
    layer6_outputs(1732) <= not((layer5_outputs(619)) xor (layer5_outputs(2997)));
    layer6_outputs(1733) <= (layer5_outputs(4747)) and not (layer5_outputs(3822));
    layer6_outputs(1734) <= not((layer5_outputs(2216)) xor (layer5_outputs(3129)));
    layer6_outputs(1735) <= not((layer5_outputs(4093)) xor (layer5_outputs(1132)));
    layer6_outputs(1736) <= not((layer5_outputs(4350)) and (layer5_outputs(688)));
    layer6_outputs(1737) <= layer5_outputs(3242);
    layer6_outputs(1738) <= not((layer5_outputs(1486)) or (layer5_outputs(1034)));
    layer6_outputs(1739) <= layer5_outputs(4664);
    layer6_outputs(1740) <= layer5_outputs(1267);
    layer6_outputs(1741) <= layer5_outputs(296);
    layer6_outputs(1742) <= (layer5_outputs(2390)) and not (layer5_outputs(4949));
    layer6_outputs(1743) <= layer5_outputs(749);
    layer6_outputs(1744) <= not((layer5_outputs(4678)) xor (layer5_outputs(2717)));
    layer6_outputs(1745) <= not(layer5_outputs(2550));
    layer6_outputs(1746) <= not(layer5_outputs(855));
    layer6_outputs(1747) <= layer5_outputs(489);
    layer6_outputs(1748) <= not(layer5_outputs(288));
    layer6_outputs(1749) <= not(layer5_outputs(1172)) or (layer5_outputs(4720));
    layer6_outputs(1750) <= (layer5_outputs(2870)) and not (layer5_outputs(4372));
    layer6_outputs(1751) <= not(layer5_outputs(1098));
    layer6_outputs(1752) <= layer5_outputs(1822);
    layer6_outputs(1753) <= not((layer5_outputs(4233)) or (layer5_outputs(1741)));
    layer6_outputs(1754) <= not(layer5_outputs(2281));
    layer6_outputs(1755) <= not(layer5_outputs(2494));
    layer6_outputs(1756) <= (layer5_outputs(5033)) and not (layer5_outputs(3028));
    layer6_outputs(1757) <= not((layer5_outputs(2647)) xor (layer5_outputs(742)));
    layer6_outputs(1758) <= layer5_outputs(60);
    layer6_outputs(1759) <= (layer5_outputs(3601)) and not (layer5_outputs(1371));
    layer6_outputs(1760) <= not((layer5_outputs(456)) or (layer5_outputs(288)));
    layer6_outputs(1761) <= not(layer5_outputs(3767));
    layer6_outputs(1762) <= (layer5_outputs(4254)) and not (layer5_outputs(2987));
    layer6_outputs(1763) <= layer5_outputs(2030);
    layer6_outputs(1764) <= (layer5_outputs(3225)) xor (layer5_outputs(1382));
    layer6_outputs(1765) <= layer5_outputs(3538);
    layer6_outputs(1766) <= (layer5_outputs(1697)) and (layer5_outputs(2943));
    layer6_outputs(1767) <= not((layer5_outputs(268)) xor (layer5_outputs(1711)));
    layer6_outputs(1768) <= layer5_outputs(1851);
    layer6_outputs(1769) <= layer5_outputs(5037);
    layer6_outputs(1770) <= not(layer5_outputs(1456)) or (layer5_outputs(484));
    layer6_outputs(1771) <= not((layer5_outputs(323)) xor (layer5_outputs(204)));
    layer6_outputs(1772) <= not(layer5_outputs(2296));
    layer6_outputs(1773) <= not((layer5_outputs(2158)) xor (layer5_outputs(2467)));
    layer6_outputs(1774) <= layer5_outputs(5094);
    layer6_outputs(1775) <= not(layer5_outputs(3747));
    layer6_outputs(1776) <= not(layer5_outputs(4148)) or (layer5_outputs(5075));
    layer6_outputs(1777) <= not(layer5_outputs(4292));
    layer6_outputs(1778) <= layer5_outputs(2481);
    layer6_outputs(1779) <= not((layer5_outputs(1642)) xor (layer5_outputs(2009)));
    layer6_outputs(1780) <= (layer5_outputs(315)) and (layer5_outputs(927));
    layer6_outputs(1781) <= layer5_outputs(2032);
    layer6_outputs(1782) <= not((layer5_outputs(753)) and (layer5_outputs(2498)));
    layer6_outputs(1783) <= not((layer5_outputs(2850)) or (layer5_outputs(2250)));
    layer6_outputs(1784) <= layer5_outputs(911);
    layer6_outputs(1785) <= layer5_outputs(988);
    layer6_outputs(1786) <= (layer5_outputs(2051)) xor (layer5_outputs(2519));
    layer6_outputs(1787) <= layer5_outputs(191);
    layer6_outputs(1788) <= layer5_outputs(4483);
    layer6_outputs(1789) <= (layer5_outputs(1517)) and (layer5_outputs(4558));
    layer6_outputs(1790) <= not(layer5_outputs(4452));
    layer6_outputs(1791) <= not(layer5_outputs(3667));
    layer6_outputs(1792) <= not(layer5_outputs(1883));
    layer6_outputs(1793) <= not(layer5_outputs(3994));
    layer6_outputs(1794) <= layer5_outputs(2811);
    layer6_outputs(1795) <= not((layer5_outputs(4055)) or (layer5_outputs(1180)));
    layer6_outputs(1796) <= not(layer5_outputs(2136));
    layer6_outputs(1797) <= (layer5_outputs(5038)) xor (layer5_outputs(2552));
    layer6_outputs(1798) <= layer5_outputs(28);
    layer6_outputs(1799) <= layer5_outputs(965);
    layer6_outputs(1800) <= layer5_outputs(1571);
    layer6_outputs(1801) <= not((layer5_outputs(1582)) and (layer5_outputs(1552)));
    layer6_outputs(1802) <= (layer5_outputs(4448)) xor (layer5_outputs(3763));
    layer6_outputs(1803) <= not(layer5_outputs(1644));
    layer6_outputs(1804) <= layer5_outputs(4308);
    layer6_outputs(1805) <= not(layer5_outputs(3475)) or (layer5_outputs(3753));
    layer6_outputs(1806) <= not((layer5_outputs(1436)) or (layer5_outputs(1694)));
    layer6_outputs(1807) <= layer5_outputs(3246);
    layer6_outputs(1808) <= not(layer5_outputs(2770));
    layer6_outputs(1809) <= not(layer5_outputs(767));
    layer6_outputs(1810) <= (layer5_outputs(2667)) xor (layer5_outputs(392));
    layer6_outputs(1811) <= not(layer5_outputs(1396));
    layer6_outputs(1812) <= layer5_outputs(529);
    layer6_outputs(1813) <= not((layer5_outputs(3064)) xor (layer5_outputs(702)));
    layer6_outputs(1814) <= not(layer5_outputs(1442));
    layer6_outputs(1815) <= layer5_outputs(2031);
    layer6_outputs(1816) <= (layer5_outputs(2588)) and (layer5_outputs(531));
    layer6_outputs(1817) <= not(layer5_outputs(4985));
    layer6_outputs(1818) <= not((layer5_outputs(3566)) or (layer5_outputs(1992)));
    layer6_outputs(1819) <= not(layer5_outputs(4723));
    layer6_outputs(1820) <= not(layer5_outputs(322));
    layer6_outputs(1821) <= layer5_outputs(1334);
    layer6_outputs(1822) <= not((layer5_outputs(4145)) xor (layer5_outputs(4270)));
    layer6_outputs(1823) <= not(layer5_outputs(3354));
    layer6_outputs(1824) <= layer5_outputs(1074);
    layer6_outputs(1825) <= not(layer5_outputs(259)) or (layer5_outputs(2723));
    layer6_outputs(1826) <= not((layer5_outputs(694)) or (layer5_outputs(1038)));
    layer6_outputs(1827) <= not(layer5_outputs(2792));
    layer6_outputs(1828) <= layer5_outputs(1419);
    layer6_outputs(1829) <= (layer5_outputs(4944)) or (layer5_outputs(2156));
    layer6_outputs(1830) <= layer5_outputs(76);
    layer6_outputs(1831) <= layer5_outputs(1315);
    layer6_outputs(1832) <= (layer5_outputs(2653)) or (layer5_outputs(4485));
    layer6_outputs(1833) <= not((layer5_outputs(3303)) and (layer5_outputs(3136)));
    layer6_outputs(1834) <= not(layer5_outputs(1533));
    layer6_outputs(1835) <= (layer5_outputs(2416)) and not (layer5_outputs(5024));
    layer6_outputs(1836) <= (layer5_outputs(1757)) xor (layer5_outputs(2340));
    layer6_outputs(1837) <= '0';
    layer6_outputs(1838) <= not(layer5_outputs(2221));
    layer6_outputs(1839) <= (layer5_outputs(2703)) and not (layer5_outputs(4974));
    layer6_outputs(1840) <= layer5_outputs(1888);
    layer6_outputs(1841) <= not((layer5_outputs(1255)) and (layer5_outputs(2192)));
    layer6_outputs(1842) <= not(layer5_outputs(4727));
    layer6_outputs(1843) <= not(layer5_outputs(3324));
    layer6_outputs(1844) <= layer5_outputs(837);
    layer6_outputs(1845) <= (layer5_outputs(1274)) and (layer5_outputs(4933));
    layer6_outputs(1846) <= not((layer5_outputs(1769)) xor (layer5_outputs(1846)));
    layer6_outputs(1847) <= layer5_outputs(5038);
    layer6_outputs(1848) <= layer5_outputs(4413);
    layer6_outputs(1849) <= (layer5_outputs(4796)) xor (layer5_outputs(3287));
    layer6_outputs(1850) <= layer5_outputs(3082);
    layer6_outputs(1851) <= not(layer5_outputs(3294));
    layer6_outputs(1852) <= (layer5_outputs(1505)) and not (layer5_outputs(2859));
    layer6_outputs(1853) <= not(layer5_outputs(5072)) or (layer5_outputs(432));
    layer6_outputs(1854) <= not(layer5_outputs(4595)) or (layer5_outputs(3104));
    layer6_outputs(1855) <= layer5_outputs(4667);
    layer6_outputs(1856) <= not(layer5_outputs(4109)) or (layer5_outputs(5061));
    layer6_outputs(1857) <= layer5_outputs(2057);
    layer6_outputs(1858) <= layer5_outputs(3030);
    layer6_outputs(1859) <= layer5_outputs(1993);
    layer6_outputs(1860) <= layer5_outputs(1189);
    layer6_outputs(1861) <= not(layer5_outputs(2584));
    layer6_outputs(1862) <= (layer5_outputs(1453)) xor (layer5_outputs(4093));
    layer6_outputs(1863) <= not(layer5_outputs(3147));
    layer6_outputs(1864) <= not(layer5_outputs(1862));
    layer6_outputs(1865) <= (layer5_outputs(3569)) and (layer5_outputs(1325));
    layer6_outputs(1866) <= not(layer5_outputs(4028));
    layer6_outputs(1867) <= not(layer5_outputs(1310)) or (layer5_outputs(1330));
    layer6_outputs(1868) <= not(layer5_outputs(919));
    layer6_outputs(1869) <= layer5_outputs(758);
    layer6_outputs(1870) <= not(layer5_outputs(4799)) or (layer5_outputs(949));
    layer6_outputs(1871) <= (layer5_outputs(142)) and (layer5_outputs(1711));
    layer6_outputs(1872) <= not((layer5_outputs(4718)) xor (layer5_outputs(4916)));
    layer6_outputs(1873) <= (layer5_outputs(2074)) or (layer5_outputs(3237));
    layer6_outputs(1874) <= not((layer5_outputs(163)) xor (layer5_outputs(2474)));
    layer6_outputs(1875) <= layer5_outputs(2595);
    layer6_outputs(1876) <= layer5_outputs(5010);
    layer6_outputs(1877) <= not(layer5_outputs(667));
    layer6_outputs(1878) <= layer5_outputs(629);
    layer6_outputs(1879) <= not(layer5_outputs(2011));
    layer6_outputs(1880) <= not((layer5_outputs(4131)) or (layer5_outputs(4396)));
    layer6_outputs(1881) <= not((layer5_outputs(4151)) and (layer5_outputs(4749)));
    layer6_outputs(1882) <= not((layer5_outputs(352)) or (layer5_outputs(424)));
    layer6_outputs(1883) <= not(layer5_outputs(53));
    layer6_outputs(1884) <= not((layer5_outputs(4795)) and (layer5_outputs(2649)));
    layer6_outputs(1885) <= not(layer5_outputs(3743));
    layer6_outputs(1886) <= not(layer5_outputs(1314));
    layer6_outputs(1887) <= (layer5_outputs(2975)) and not (layer5_outputs(3894));
    layer6_outputs(1888) <= (layer5_outputs(2660)) and not (layer5_outputs(3205));
    layer6_outputs(1889) <= not(layer5_outputs(3323));
    layer6_outputs(1890) <= not(layer5_outputs(2003));
    layer6_outputs(1891) <= not((layer5_outputs(3973)) xor (layer5_outputs(3078)));
    layer6_outputs(1892) <= not(layer5_outputs(1191));
    layer6_outputs(1893) <= not(layer5_outputs(3116));
    layer6_outputs(1894) <= not(layer5_outputs(2530));
    layer6_outputs(1895) <= (layer5_outputs(3740)) xor (layer5_outputs(5084));
    layer6_outputs(1896) <= layer5_outputs(4997);
    layer6_outputs(1897) <= layer5_outputs(4908);
    layer6_outputs(1898) <= (layer5_outputs(969)) and not (layer5_outputs(103));
    layer6_outputs(1899) <= '1';
    layer6_outputs(1900) <= (layer5_outputs(5101)) and (layer5_outputs(3171));
    layer6_outputs(1901) <= layer5_outputs(1102);
    layer6_outputs(1902) <= layer5_outputs(4777);
    layer6_outputs(1903) <= layer5_outputs(2392);
    layer6_outputs(1904) <= not(layer5_outputs(4110));
    layer6_outputs(1905) <= (layer5_outputs(1290)) and not (layer5_outputs(4147));
    layer6_outputs(1906) <= not(layer5_outputs(663)) or (layer5_outputs(2948));
    layer6_outputs(1907) <= not((layer5_outputs(1266)) xor (layer5_outputs(4788)));
    layer6_outputs(1908) <= not(layer5_outputs(4380)) or (layer5_outputs(3439));
    layer6_outputs(1909) <= (layer5_outputs(1025)) and (layer5_outputs(1353));
    layer6_outputs(1910) <= layer5_outputs(1760);
    layer6_outputs(1911) <= '1';
    layer6_outputs(1912) <= layer5_outputs(2537);
    layer6_outputs(1913) <= (layer5_outputs(817)) xor (layer5_outputs(3643));
    layer6_outputs(1914) <= (layer5_outputs(1971)) xor (layer5_outputs(3537));
    layer6_outputs(1915) <= (layer5_outputs(2590)) or (layer5_outputs(3633));
    layer6_outputs(1916) <= not((layer5_outputs(1003)) xor (layer5_outputs(2300)));
    layer6_outputs(1917) <= (layer5_outputs(800)) xor (layer5_outputs(1923));
    layer6_outputs(1918) <= layer5_outputs(4149);
    layer6_outputs(1919) <= layer5_outputs(3487);
    layer6_outputs(1920) <= not((layer5_outputs(4969)) xor (layer5_outputs(1948)));
    layer6_outputs(1921) <= layer5_outputs(3974);
    layer6_outputs(1922) <= not(layer5_outputs(2260));
    layer6_outputs(1923) <= not(layer5_outputs(4433));
    layer6_outputs(1924) <= not((layer5_outputs(1222)) or (layer5_outputs(2564)));
    layer6_outputs(1925) <= not((layer5_outputs(1511)) xor (layer5_outputs(3910)));
    layer6_outputs(1926) <= not(layer5_outputs(4626));
    layer6_outputs(1927) <= not(layer5_outputs(2328));
    layer6_outputs(1928) <= not((layer5_outputs(536)) and (layer5_outputs(2568)));
    layer6_outputs(1929) <= layer5_outputs(292);
    layer6_outputs(1930) <= not(layer5_outputs(958)) or (layer5_outputs(2491));
    layer6_outputs(1931) <= (layer5_outputs(861)) or (layer5_outputs(563));
    layer6_outputs(1932) <= not(layer5_outputs(1616));
    layer6_outputs(1933) <= layer5_outputs(3424);
    layer6_outputs(1934) <= layer5_outputs(3246);
    layer6_outputs(1935) <= not((layer5_outputs(5088)) or (layer5_outputs(4257)));
    layer6_outputs(1936) <= layer5_outputs(4032);
    layer6_outputs(1937) <= not((layer5_outputs(765)) or (layer5_outputs(2657)));
    layer6_outputs(1938) <= layer5_outputs(2078);
    layer6_outputs(1939) <= not(layer5_outputs(5020)) or (layer5_outputs(4998));
    layer6_outputs(1940) <= not((layer5_outputs(1468)) or (layer5_outputs(4927)));
    layer6_outputs(1941) <= (layer5_outputs(4241)) and (layer5_outputs(3625));
    layer6_outputs(1942) <= layer5_outputs(26);
    layer6_outputs(1943) <= not(layer5_outputs(1763));
    layer6_outputs(1944) <= layer5_outputs(2313);
    layer6_outputs(1945) <= not(layer5_outputs(191)) or (layer5_outputs(1543));
    layer6_outputs(1946) <= layer5_outputs(1188);
    layer6_outputs(1947) <= layer5_outputs(503);
    layer6_outputs(1948) <= not(layer5_outputs(5059));
    layer6_outputs(1949) <= not(layer5_outputs(3686));
    layer6_outputs(1950) <= not(layer5_outputs(3508)) or (layer5_outputs(598));
    layer6_outputs(1951) <= (layer5_outputs(2430)) xor (layer5_outputs(3154));
    layer6_outputs(1952) <= not(layer5_outputs(2029));
    layer6_outputs(1953) <= not((layer5_outputs(4043)) and (layer5_outputs(3151)));
    layer6_outputs(1954) <= not(layer5_outputs(3073));
    layer6_outputs(1955) <= not((layer5_outputs(161)) or (layer5_outputs(234)));
    layer6_outputs(1956) <= not((layer5_outputs(4562)) xor (layer5_outputs(3233)));
    layer6_outputs(1957) <= not(layer5_outputs(4891)) or (layer5_outputs(3670));
    layer6_outputs(1958) <= not(layer5_outputs(2935));
    layer6_outputs(1959) <= layer5_outputs(4450);
    layer6_outputs(1960) <= (layer5_outputs(4121)) and (layer5_outputs(864));
    layer6_outputs(1961) <= (layer5_outputs(4795)) or (layer5_outputs(1493));
    layer6_outputs(1962) <= (layer5_outputs(1465)) xor (layer5_outputs(3195));
    layer6_outputs(1963) <= not(layer5_outputs(1807));
    layer6_outputs(1964) <= layer5_outputs(4801);
    layer6_outputs(1965) <= layer5_outputs(336);
    layer6_outputs(1966) <= not((layer5_outputs(2396)) and (layer5_outputs(761)));
    layer6_outputs(1967) <= not(layer5_outputs(306));
    layer6_outputs(1968) <= not(layer5_outputs(266));
    layer6_outputs(1969) <= not((layer5_outputs(2364)) or (layer5_outputs(3622)));
    layer6_outputs(1970) <= not(layer5_outputs(3596)) or (layer5_outputs(3332));
    layer6_outputs(1971) <= layer5_outputs(56);
    layer6_outputs(1972) <= not(layer5_outputs(2044));
    layer6_outputs(1973) <= layer5_outputs(2557);
    layer6_outputs(1974) <= not(layer5_outputs(4273));
    layer6_outputs(1975) <= layer5_outputs(4643);
    layer6_outputs(1976) <= layer5_outputs(1011);
    layer6_outputs(1977) <= not(layer5_outputs(1452));
    layer6_outputs(1978) <= not(layer5_outputs(4323)) or (layer5_outputs(4563));
    layer6_outputs(1979) <= (layer5_outputs(3049)) and not (layer5_outputs(2));
    layer6_outputs(1980) <= not(layer5_outputs(2695));
    layer6_outputs(1981) <= not(layer5_outputs(4355));
    layer6_outputs(1982) <= not(layer5_outputs(3117)) or (layer5_outputs(257));
    layer6_outputs(1983) <= layer5_outputs(3953);
    layer6_outputs(1984) <= not(layer5_outputs(3606));
    layer6_outputs(1985) <= (layer5_outputs(2006)) or (layer5_outputs(2718));
    layer6_outputs(1986) <= (layer5_outputs(419)) and not (layer5_outputs(4803));
    layer6_outputs(1987) <= not(layer5_outputs(3586)) or (layer5_outputs(1584));
    layer6_outputs(1988) <= not(layer5_outputs(2900));
    layer6_outputs(1989) <= not(layer5_outputs(4504));
    layer6_outputs(1990) <= not(layer5_outputs(758));
    layer6_outputs(1991) <= (layer5_outputs(3154)) and not (layer5_outputs(3466));
    layer6_outputs(1992) <= (layer5_outputs(2363)) and not (layer5_outputs(2990));
    layer6_outputs(1993) <= not((layer5_outputs(1175)) or (layer5_outputs(841)));
    layer6_outputs(1994) <= not((layer5_outputs(1389)) and (layer5_outputs(4813)));
    layer6_outputs(1995) <= layer5_outputs(1838);
    layer6_outputs(1996) <= layer5_outputs(4001);
    layer6_outputs(1997) <= layer5_outputs(2819);
    layer6_outputs(1998) <= layer5_outputs(4712);
    layer6_outputs(1999) <= not((layer5_outputs(2680)) xor (layer5_outputs(4336)));
    layer6_outputs(2000) <= layer5_outputs(4549);
    layer6_outputs(2001) <= (layer5_outputs(700)) and (layer5_outputs(4443));
    layer6_outputs(2002) <= (layer5_outputs(3331)) and (layer5_outputs(4531));
    layer6_outputs(2003) <= not(layer5_outputs(476)) or (layer5_outputs(3433));
    layer6_outputs(2004) <= not(layer5_outputs(2565));
    layer6_outputs(2005) <= not((layer5_outputs(3484)) or (layer5_outputs(2621)));
    layer6_outputs(2006) <= not(layer5_outputs(3141)) or (layer5_outputs(2960));
    layer6_outputs(2007) <= not(layer5_outputs(2904)) or (layer5_outputs(1562));
    layer6_outputs(2008) <= (layer5_outputs(4126)) and (layer5_outputs(1355));
    layer6_outputs(2009) <= not(layer5_outputs(3932));
    layer6_outputs(2010) <= not(layer5_outputs(4411));
    layer6_outputs(2011) <= not(layer5_outputs(2651));
    layer6_outputs(2012) <= (layer5_outputs(1001)) and not (layer5_outputs(1929));
    layer6_outputs(2013) <= layer5_outputs(337);
    layer6_outputs(2014) <= (layer5_outputs(253)) and not (layer5_outputs(3603));
    layer6_outputs(2015) <= (layer5_outputs(4390)) and not (layer5_outputs(685));
    layer6_outputs(2016) <= (layer5_outputs(2380)) and not (layer5_outputs(4978));
    layer6_outputs(2017) <= not(layer5_outputs(2029));
    layer6_outputs(2018) <= not(layer5_outputs(4599));
    layer6_outputs(2019) <= layer5_outputs(36);
    layer6_outputs(2020) <= not(layer5_outputs(5051));
    layer6_outputs(2021) <= not((layer5_outputs(727)) or (layer5_outputs(29)));
    layer6_outputs(2022) <= (layer5_outputs(1595)) and not (layer5_outputs(1200));
    layer6_outputs(2023) <= layer5_outputs(3987);
    layer6_outputs(2024) <= not(layer5_outputs(2182));
    layer6_outputs(2025) <= layer5_outputs(3732);
    layer6_outputs(2026) <= not((layer5_outputs(2405)) xor (layer5_outputs(1704)));
    layer6_outputs(2027) <= not(layer5_outputs(150));
    layer6_outputs(2028) <= not(layer5_outputs(2416)) or (layer5_outputs(4671));
    layer6_outputs(2029) <= not(layer5_outputs(3732));
    layer6_outputs(2030) <= not((layer5_outputs(2205)) and (layer5_outputs(3406)));
    layer6_outputs(2031) <= not((layer5_outputs(2507)) and (layer5_outputs(2942)));
    layer6_outputs(2032) <= layer5_outputs(4392);
    layer6_outputs(2033) <= layer5_outputs(3375);
    layer6_outputs(2034) <= (layer5_outputs(4577)) and not (layer5_outputs(4651));
    layer6_outputs(2035) <= not(layer5_outputs(1621));
    layer6_outputs(2036) <= (layer5_outputs(75)) xor (layer5_outputs(5056));
    layer6_outputs(2037) <= not(layer5_outputs(4961));
    layer6_outputs(2038) <= not((layer5_outputs(2652)) xor (layer5_outputs(2676)));
    layer6_outputs(2039) <= not(layer5_outputs(1749)) or (layer5_outputs(1765));
    layer6_outputs(2040) <= not((layer5_outputs(2927)) and (layer5_outputs(1684)));
    layer6_outputs(2041) <= layer5_outputs(2331);
    layer6_outputs(2042) <= not(layer5_outputs(2175));
    layer6_outputs(2043) <= (layer5_outputs(2926)) and (layer5_outputs(2646));
    layer6_outputs(2044) <= not(layer5_outputs(3213));
    layer6_outputs(2045) <= not(layer5_outputs(748));
    layer6_outputs(2046) <= layer5_outputs(260);
    layer6_outputs(2047) <= layer5_outputs(183);
    layer6_outputs(2048) <= not(layer5_outputs(658));
    layer6_outputs(2049) <= (layer5_outputs(677)) xor (layer5_outputs(2092));
    layer6_outputs(2050) <= not(layer5_outputs(3964));
    layer6_outputs(2051) <= layer5_outputs(4261);
    layer6_outputs(2052) <= layer5_outputs(22);
    layer6_outputs(2053) <= not((layer5_outputs(750)) xor (layer5_outputs(2630)));
    layer6_outputs(2054) <= (layer5_outputs(61)) and not (layer5_outputs(4009));
    layer6_outputs(2055) <= (layer5_outputs(2549)) xor (layer5_outputs(3054));
    layer6_outputs(2056) <= layer5_outputs(2696);
    layer6_outputs(2057) <= not(layer5_outputs(4867)) or (layer5_outputs(3228));
    layer6_outputs(2058) <= (layer5_outputs(3128)) and (layer5_outputs(1569));
    layer6_outputs(2059) <= not((layer5_outputs(4186)) xor (layer5_outputs(56)));
    layer6_outputs(2060) <= layer5_outputs(1074);
    layer6_outputs(2061) <= layer5_outputs(2359);
    layer6_outputs(2062) <= layer5_outputs(5027);
    layer6_outputs(2063) <= not(layer5_outputs(1550));
    layer6_outputs(2064) <= not(layer5_outputs(4832));
    layer6_outputs(2065) <= not(layer5_outputs(1417));
    layer6_outputs(2066) <= not(layer5_outputs(4082)) or (layer5_outputs(712));
    layer6_outputs(2067) <= layer5_outputs(3781);
    layer6_outputs(2068) <= (layer5_outputs(4277)) and not (layer5_outputs(3932));
    layer6_outputs(2069) <= not((layer5_outputs(655)) xor (layer5_outputs(4656)));
    layer6_outputs(2070) <= (layer5_outputs(3886)) xor (layer5_outputs(3305));
    layer6_outputs(2071) <= not(layer5_outputs(1610));
    layer6_outputs(2072) <= not((layer5_outputs(788)) xor (layer5_outputs(2473)));
    layer6_outputs(2073) <= (layer5_outputs(3859)) and not (layer5_outputs(4561));
    layer6_outputs(2074) <= layer5_outputs(1632);
    layer6_outputs(2075) <= layer5_outputs(1636);
    layer6_outputs(2076) <= not((layer5_outputs(2783)) and (layer5_outputs(1759)));
    layer6_outputs(2077) <= layer5_outputs(2461);
    layer6_outputs(2078) <= (layer5_outputs(0)) xor (layer5_outputs(851));
    layer6_outputs(2079) <= not((layer5_outputs(1846)) xor (layer5_outputs(65)));
    layer6_outputs(2080) <= layer5_outputs(1284);
    layer6_outputs(2081) <= not(layer5_outputs(4157));
    layer6_outputs(2082) <= not(layer5_outputs(4685));
    layer6_outputs(2083) <= layer5_outputs(5011);
    layer6_outputs(2084) <= layer5_outputs(565);
    layer6_outputs(2085) <= not(layer5_outputs(1963));
    layer6_outputs(2086) <= not((layer5_outputs(2762)) xor (layer5_outputs(3519)));
    layer6_outputs(2087) <= (layer5_outputs(2793)) and not (layer5_outputs(4865));
    layer6_outputs(2088) <= not((layer5_outputs(2462)) and (layer5_outputs(2816)));
    layer6_outputs(2089) <= (layer5_outputs(1159)) or (layer5_outputs(2675));
    layer6_outputs(2090) <= (layer5_outputs(2605)) xor (layer5_outputs(2499));
    layer6_outputs(2091) <= (layer5_outputs(3370)) and not (layer5_outputs(2342));
    layer6_outputs(2092) <= not((layer5_outputs(823)) and (layer5_outputs(2922)));
    layer6_outputs(2093) <= '1';
    layer6_outputs(2094) <= not(layer5_outputs(2134));
    layer6_outputs(2095) <= not(layer5_outputs(5007));
    layer6_outputs(2096) <= (layer5_outputs(1510)) or (layer5_outputs(465));
    layer6_outputs(2097) <= not((layer5_outputs(1368)) or (layer5_outputs(4836)));
    layer6_outputs(2098) <= not(layer5_outputs(128)) or (layer5_outputs(3437));
    layer6_outputs(2099) <= (layer5_outputs(143)) and (layer5_outputs(1249));
    layer6_outputs(2100) <= not(layer5_outputs(4719));
    layer6_outputs(2101) <= layer5_outputs(2534);
    layer6_outputs(2102) <= layer5_outputs(2313);
    layer6_outputs(2103) <= layer5_outputs(3613);
    layer6_outputs(2104) <= layer5_outputs(2176);
    layer6_outputs(2105) <= not((layer5_outputs(369)) or (layer5_outputs(779)));
    layer6_outputs(2106) <= layer5_outputs(276);
    layer6_outputs(2107) <= not(layer5_outputs(536));
    layer6_outputs(2108) <= layer5_outputs(3003);
    layer6_outputs(2109) <= (layer5_outputs(330)) xor (layer5_outputs(4306));
    layer6_outputs(2110) <= not(layer5_outputs(2758));
    layer6_outputs(2111) <= (layer5_outputs(1273)) and not (layer5_outputs(1220));
    layer6_outputs(2112) <= layer5_outputs(1952);
    layer6_outputs(2113) <= not(layer5_outputs(3681));
    layer6_outputs(2114) <= not(layer5_outputs(502));
    layer6_outputs(2115) <= layer5_outputs(2000);
    layer6_outputs(2116) <= layer5_outputs(5092);
    layer6_outputs(2117) <= not(layer5_outputs(1625));
    layer6_outputs(2118) <= (layer5_outputs(3215)) or (layer5_outputs(2558));
    layer6_outputs(2119) <= not((layer5_outputs(2361)) xor (layer5_outputs(3620)));
    layer6_outputs(2120) <= (layer5_outputs(2311)) and not (layer5_outputs(55));
    layer6_outputs(2121) <= not(layer5_outputs(2689));
    layer6_outputs(2122) <= (layer5_outputs(3641)) and (layer5_outputs(3906));
    layer6_outputs(2123) <= layer5_outputs(3366);
    layer6_outputs(2124) <= not(layer5_outputs(3692));
    layer6_outputs(2125) <= (layer5_outputs(4587)) and not (layer5_outputs(3996));
    layer6_outputs(2126) <= not(layer5_outputs(4192)) or (layer5_outputs(1887));
    layer6_outputs(2127) <= (layer5_outputs(2267)) and (layer5_outputs(4769));
    layer6_outputs(2128) <= not(layer5_outputs(3364));
    layer6_outputs(2129) <= (layer5_outputs(556)) xor (layer5_outputs(2676));
    layer6_outputs(2130) <= (layer5_outputs(904)) and (layer5_outputs(3745));
    layer6_outputs(2131) <= (layer5_outputs(2983)) xor (layer5_outputs(4609));
    layer6_outputs(2132) <= not((layer5_outputs(2344)) xor (layer5_outputs(595)));
    layer6_outputs(2133) <= not(layer5_outputs(231));
    layer6_outputs(2134) <= (layer5_outputs(2213)) xor (layer5_outputs(475));
    layer6_outputs(2135) <= not(layer5_outputs(4573)) or (layer5_outputs(3417));
    layer6_outputs(2136) <= layer5_outputs(2301);
    layer6_outputs(2137) <= not((layer5_outputs(1793)) xor (layer5_outputs(1946)));
    layer6_outputs(2138) <= not(layer5_outputs(4746));
    layer6_outputs(2139) <= layer5_outputs(1573);
    layer6_outputs(2140) <= layer5_outputs(2010);
    layer6_outputs(2141) <= not(layer5_outputs(1844));
    layer6_outputs(2142) <= '0';
    layer6_outputs(2143) <= not(layer5_outputs(348));
    layer6_outputs(2144) <= (layer5_outputs(2714)) and not (layer5_outputs(1053));
    layer6_outputs(2145) <= layer5_outputs(535);
    layer6_outputs(2146) <= not((layer5_outputs(3534)) xor (layer5_outputs(4702)));
    layer6_outputs(2147) <= layer5_outputs(3546);
    layer6_outputs(2148) <= not(layer5_outputs(3888));
    layer6_outputs(2149) <= not((layer5_outputs(546)) xor (layer5_outputs(3258)));
    layer6_outputs(2150) <= layer5_outputs(4313);
    layer6_outputs(2151) <= layer5_outputs(245);
    layer6_outputs(2152) <= layer5_outputs(1778);
    layer6_outputs(2153) <= not(layer5_outputs(1391));
    layer6_outputs(2154) <= (layer5_outputs(156)) and not (layer5_outputs(319));
    layer6_outputs(2155) <= not((layer5_outputs(427)) xor (layer5_outputs(4754)));
    layer6_outputs(2156) <= not(layer5_outputs(277)) or (layer5_outputs(3680));
    layer6_outputs(2157) <= not(layer5_outputs(2047));
    layer6_outputs(2158) <= not((layer5_outputs(1760)) and (layer5_outputs(4692)));
    layer6_outputs(2159) <= layer5_outputs(1280);
    layer6_outputs(2160) <= (layer5_outputs(3560)) xor (layer5_outputs(121));
    layer6_outputs(2161) <= layer5_outputs(2113);
    layer6_outputs(2162) <= (layer5_outputs(2213)) and not (layer5_outputs(3531));
    layer6_outputs(2163) <= not(layer5_outputs(1167));
    layer6_outputs(2164) <= layer5_outputs(2314);
    layer6_outputs(2165) <= (layer5_outputs(550)) and (layer5_outputs(1842));
    layer6_outputs(2166) <= not((layer5_outputs(1361)) or (layer5_outputs(246)));
    layer6_outputs(2167) <= not(layer5_outputs(2656));
    layer6_outputs(2168) <= (layer5_outputs(309)) and not (layer5_outputs(3384));
    layer6_outputs(2169) <= (layer5_outputs(4595)) and not (layer5_outputs(348));
    layer6_outputs(2170) <= (layer5_outputs(4224)) xor (layer5_outputs(3249));
    layer6_outputs(2171) <= not(layer5_outputs(2868));
    layer6_outputs(2172) <= not(layer5_outputs(3713));
    layer6_outputs(2173) <= not((layer5_outputs(2826)) and (layer5_outputs(1684)));
    layer6_outputs(2174) <= not((layer5_outputs(3456)) or (layer5_outputs(1385)));
    layer6_outputs(2175) <= not(layer5_outputs(2681));
    layer6_outputs(2176) <= (layer5_outputs(3517)) xor (layer5_outputs(2453));
    layer6_outputs(2177) <= (layer5_outputs(3512)) and not (layer5_outputs(5010));
    layer6_outputs(2178) <= not(layer5_outputs(2103));
    layer6_outputs(2179) <= '1';
    layer6_outputs(2180) <= layer5_outputs(2054);
    layer6_outputs(2181) <= not(layer5_outputs(4237));
    layer6_outputs(2182) <= not(layer5_outputs(849));
    layer6_outputs(2183) <= not(layer5_outputs(4061));
    layer6_outputs(2184) <= (layer5_outputs(71)) and not (layer5_outputs(444));
    layer6_outputs(2185) <= not((layer5_outputs(4956)) xor (layer5_outputs(1961)));
    layer6_outputs(2186) <= (layer5_outputs(3417)) and not (layer5_outputs(1010));
    layer6_outputs(2187) <= not(layer5_outputs(4978));
    layer6_outputs(2188) <= layer5_outputs(3763);
    layer6_outputs(2189) <= (layer5_outputs(2598)) and not (layer5_outputs(1719));
    layer6_outputs(2190) <= (layer5_outputs(3156)) and not (layer5_outputs(3711));
    layer6_outputs(2191) <= not(layer5_outputs(4811));
    layer6_outputs(2192) <= not((layer5_outputs(1431)) or (layer5_outputs(2648)));
    layer6_outputs(2193) <= not((layer5_outputs(3956)) xor (layer5_outputs(1741)));
    layer6_outputs(2194) <= layer5_outputs(4008);
    layer6_outputs(2195) <= not((layer5_outputs(3346)) and (layer5_outputs(1061)));
    layer6_outputs(2196) <= (layer5_outputs(3108)) xor (layer5_outputs(640));
    layer6_outputs(2197) <= (layer5_outputs(1871)) xor (layer5_outputs(3810));
    layer6_outputs(2198) <= not((layer5_outputs(726)) or (layer5_outputs(89)));
    layer6_outputs(2199) <= not(layer5_outputs(3328));
    layer6_outputs(2200) <= not((layer5_outputs(105)) or (layer5_outputs(2139)));
    layer6_outputs(2201) <= not(layer5_outputs(3002));
    layer6_outputs(2202) <= layer5_outputs(908);
    layer6_outputs(2203) <= not(layer5_outputs(4841));
    layer6_outputs(2204) <= (layer5_outputs(3973)) and not (layer5_outputs(4188));
    layer6_outputs(2205) <= layer5_outputs(4929);
    layer6_outputs(2206) <= not(layer5_outputs(719));
    layer6_outputs(2207) <= not(layer5_outputs(3111));
    layer6_outputs(2208) <= layer5_outputs(2462);
    layer6_outputs(2209) <= layer5_outputs(4836);
    layer6_outputs(2210) <= not(layer5_outputs(1196));
    layer6_outputs(2211) <= not((layer5_outputs(2858)) xor (layer5_outputs(1019)));
    layer6_outputs(2212) <= not(layer5_outputs(1693));
    layer6_outputs(2213) <= not((layer5_outputs(3239)) or (layer5_outputs(1999)));
    layer6_outputs(2214) <= layer5_outputs(3200);
    layer6_outputs(2215) <= layer5_outputs(2930);
    layer6_outputs(2216) <= (layer5_outputs(4405)) or (layer5_outputs(1424));
    layer6_outputs(2217) <= layer5_outputs(4158);
    layer6_outputs(2218) <= not((layer5_outputs(1618)) xor (layer5_outputs(1020)));
    layer6_outputs(2219) <= not((layer5_outputs(3449)) xor (layer5_outputs(301)));
    layer6_outputs(2220) <= (layer5_outputs(2996)) and not (layer5_outputs(1764));
    layer6_outputs(2221) <= not(layer5_outputs(5007));
    layer6_outputs(2222) <= (layer5_outputs(2881)) and (layer5_outputs(4696));
    layer6_outputs(2223) <= not(layer5_outputs(2750));
    layer6_outputs(2224) <= not(layer5_outputs(2946)) or (layer5_outputs(3784));
    layer6_outputs(2225) <= (layer5_outputs(1661)) and (layer5_outputs(3598));
    layer6_outputs(2226) <= not((layer5_outputs(2703)) or (layer5_outputs(1829)));
    layer6_outputs(2227) <= not(layer5_outputs(4438));
    layer6_outputs(2228) <= not(layer5_outputs(596));
    layer6_outputs(2229) <= not(layer5_outputs(3696));
    layer6_outputs(2230) <= not((layer5_outputs(4589)) and (layer5_outputs(952)));
    layer6_outputs(2231) <= not((layer5_outputs(2563)) xor (layer5_outputs(556)));
    layer6_outputs(2232) <= layer5_outputs(208);
    layer6_outputs(2233) <= not(layer5_outputs(512)) or (layer5_outputs(2173));
    layer6_outputs(2234) <= not(layer5_outputs(4658));
    layer6_outputs(2235) <= layer5_outputs(217);
    layer6_outputs(2236) <= not(layer5_outputs(4606));
    layer6_outputs(2237) <= not(layer5_outputs(2959));
    layer6_outputs(2238) <= not((layer5_outputs(3724)) and (layer5_outputs(3110)));
    layer6_outputs(2239) <= '0';
    layer6_outputs(2240) <= layer5_outputs(1295);
    layer6_outputs(2241) <= layer5_outputs(2824);
    layer6_outputs(2242) <= not((layer5_outputs(4525)) or (layer5_outputs(1738)));
    layer6_outputs(2243) <= layer5_outputs(3748);
    layer6_outputs(2244) <= not(layer5_outputs(2672));
    layer6_outputs(2245) <= (layer5_outputs(1853)) xor (layer5_outputs(4940));
    layer6_outputs(2246) <= '0';
    layer6_outputs(2247) <= (layer5_outputs(4701)) and (layer5_outputs(1057));
    layer6_outputs(2248) <= not(layer5_outputs(3068)) or (layer5_outputs(60));
    layer6_outputs(2249) <= (layer5_outputs(3474)) and not (layer5_outputs(4303));
    layer6_outputs(2250) <= not((layer5_outputs(1872)) or (layer5_outputs(4741)));
    layer6_outputs(2251) <= (layer5_outputs(2051)) and not (layer5_outputs(3052));
    layer6_outputs(2252) <= (layer5_outputs(2322)) and (layer5_outputs(73));
    layer6_outputs(2253) <= not(layer5_outputs(3221));
    layer6_outputs(2254) <= (layer5_outputs(1602)) and not (layer5_outputs(509));
    layer6_outputs(2255) <= layer5_outputs(3444);
    layer6_outputs(2256) <= (layer5_outputs(4681)) or (layer5_outputs(2872));
    layer6_outputs(2257) <= layer5_outputs(2980);
    layer6_outputs(2258) <= not(layer5_outputs(2091));
    layer6_outputs(2259) <= not(layer5_outputs(2210));
    layer6_outputs(2260) <= (layer5_outputs(6)) xor (layer5_outputs(1344));
    layer6_outputs(2261) <= not((layer5_outputs(4266)) or (layer5_outputs(4521)));
    layer6_outputs(2262) <= not(layer5_outputs(1090)) or (layer5_outputs(2341));
    layer6_outputs(2263) <= not(layer5_outputs(3143));
    layer6_outputs(2264) <= layer5_outputs(3575);
    layer6_outputs(2265) <= (layer5_outputs(2441)) xor (layer5_outputs(678));
    layer6_outputs(2266) <= not(layer5_outputs(1617));
    layer6_outputs(2267) <= layer5_outputs(602);
    layer6_outputs(2268) <= layer5_outputs(833);
    layer6_outputs(2269) <= (layer5_outputs(3507)) xor (layer5_outputs(688));
    layer6_outputs(2270) <= (layer5_outputs(1496)) or (layer5_outputs(2209));
    layer6_outputs(2271) <= not(layer5_outputs(747));
    layer6_outputs(2272) <= (layer5_outputs(477)) xor (layer5_outputs(2688));
    layer6_outputs(2273) <= layer5_outputs(3356);
    layer6_outputs(2274) <= layer5_outputs(3153);
    layer6_outputs(2275) <= not(layer5_outputs(4357)) or (layer5_outputs(1065));
    layer6_outputs(2276) <= layer5_outputs(2626);
    layer6_outputs(2277) <= layer5_outputs(1629);
    layer6_outputs(2278) <= (layer5_outputs(3183)) xor (layer5_outputs(3613));
    layer6_outputs(2279) <= layer5_outputs(4569);
    layer6_outputs(2280) <= not(layer5_outputs(3518));
    layer6_outputs(2281) <= '1';
    layer6_outputs(2282) <= layer5_outputs(3734);
    layer6_outputs(2283) <= layer5_outputs(2245);
    layer6_outputs(2284) <= (layer5_outputs(1361)) or (layer5_outputs(1779));
    layer6_outputs(2285) <= layer5_outputs(4890);
    layer6_outputs(2286) <= layer5_outputs(2520);
    layer6_outputs(2287) <= (layer5_outputs(4267)) and not (layer5_outputs(992));
    layer6_outputs(2288) <= not(layer5_outputs(380));
    layer6_outputs(2289) <= layer5_outputs(372);
    layer6_outputs(2290) <= not(layer5_outputs(580));
    layer6_outputs(2291) <= '1';
    layer6_outputs(2292) <= not(layer5_outputs(576));
    layer6_outputs(2293) <= (layer5_outputs(1128)) xor (layer5_outputs(2560));
    layer6_outputs(2294) <= layer5_outputs(1446);
    layer6_outputs(2295) <= (layer5_outputs(418)) and not (layer5_outputs(1137));
    layer6_outputs(2296) <= (layer5_outputs(2581)) and not (layer5_outputs(2104));
    layer6_outputs(2297) <= not(layer5_outputs(1913)) or (layer5_outputs(565));
    layer6_outputs(2298) <= (layer5_outputs(4060)) xor (layer5_outputs(2637));
    layer6_outputs(2299) <= layer5_outputs(1020);
    layer6_outputs(2300) <= layer5_outputs(2511);
    layer6_outputs(2301) <= layer5_outputs(1501);
    layer6_outputs(2302) <= not(layer5_outputs(1007));
    layer6_outputs(2303) <= (layer5_outputs(1653)) xor (layer5_outputs(2642));
    layer6_outputs(2304) <= layer5_outputs(3138);
    layer6_outputs(2305) <= not((layer5_outputs(4937)) and (layer5_outputs(4216)));
    layer6_outputs(2306) <= not(layer5_outputs(453));
    layer6_outputs(2307) <= layer5_outputs(3677);
    layer6_outputs(2308) <= not(layer5_outputs(2876)) or (layer5_outputs(1966));
    layer6_outputs(2309) <= not((layer5_outputs(1999)) or (layer5_outputs(2602)));
    layer6_outputs(2310) <= not((layer5_outputs(695)) xor (layer5_outputs(405)));
    layer6_outputs(2311) <= not(layer5_outputs(4270));
    layer6_outputs(2312) <= (layer5_outputs(267)) and not (layer5_outputs(3067));
    layer6_outputs(2313) <= (layer5_outputs(2943)) xor (layer5_outputs(1795));
    layer6_outputs(2314) <= layer5_outputs(1805);
    layer6_outputs(2315) <= layer5_outputs(4336);
    layer6_outputs(2316) <= (layer5_outputs(1398)) and (layer5_outputs(1707));
    layer6_outputs(2317) <= (layer5_outputs(1573)) and not (layer5_outputs(125));
    layer6_outputs(2318) <= layer5_outputs(1503);
    layer6_outputs(2319) <= not((layer5_outputs(3841)) xor (layer5_outputs(4728)));
    layer6_outputs(2320) <= not(layer5_outputs(2492)) or (layer5_outputs(3485));
    layer6_outputs(2321) <= (layer5_outputs(1916)) xor (layer5_outputs(5105));
    layer6_outputs(2322) <= not((layer5_outputs(956)) xor (layer5_outputs(1133)));
    layer6_outputs(2323) <= layer5_outputs(1560);
    layer6_outputs(2324) <= not((layer5_outputs(3564)) and (layer5_outputs(4974)));
    layer6_outputs(2325) <= layer5_outputs(2557);
    layer6_outputs(2326) <= layer5_outputs(540);
    layer6_outputs(2327) <= layer5_outputs(2153);
    layer6_outputs(2328) <= layer5_outputs(3895);
    layer6_outputs(2329) <= layer5_outputs(1994);
    layer6_outputs(2330) <= layer5_outputs(4129);
    layer6_outputs(2331) <= (layer5_outputs(3836)) or (layer5_outputs(4418));
    layer6_outputs(2332) <= not((layer5_outputs(439)) or (layer5_outputs(4575)));
    layer6_outputs(2333) <= layer5_outputs(4810);
    layer6_outputs(2334) <= not((layer5_outputs(4255)) and (layer5_outputs(3725)));
    layer6_outputs(2335) <= not(layer5_outputs(3336));
    layer6_outputs(2336) <= not(layer5_outputs(3343));
    layer6_outputs(2337) <= not((layer5_outputs(3963)) xor (layer5_outputs(2863)));
    layer6_outputs(2338) <= not((layer5_outputs(3007)) xor (layer5_outputs(4419)));
    layer6_outputs(2339) <= layer5_outputs(592);
    layer6_outputs(2340) <= not(layer5_outputs(2938));
    layer6_outputs(2341) <= layer5_outputs(4115);
    layer6_outputs(2342) <= not(layer5_outputs(1318));
    layer6_outputs(2343) <= not(layer5_outputs(2129));
    layer6_outputs(2344) <= layer5_outputs(4102);
    layer6_outputs(2345) <= layer5_outputs(3296);
    layer6_outputs(2346) <= (layer5_outputs(420)) and not (layer5_outputs(4260));
    layer6_outputs(2347) <= not(layer5_outputs(1204));
    layer6_outputs(2348) <= not(layer5_outputs(3370)) or (layer5_outputs(1903));
    layer6_outputs(2349) <= (layer5_outputs(814)) xor (layer5_outputs(1518));
    layer6_outputs(2350) <= not(layer5_outputs(1227));
    layer6_outputs(2351) <= (layer5_outputs(2675)) xor (layer5_outputs(698));
    layer6_outputs(2352) <= '1';
    layer6_outputs(2353) <= not(layer5_outputs(1946));
    layer6_outputs(2354) <= not(layer5_outputs(1482));
    layer6_outputs(2355) <= layer5_outputs(4139);
    layer6_outputs(2356) <= not(layer5_outputs(1166));
    layer6_outputs(2357) <= not(layer5_outputs(4641));
    layer6_outputs(2358) <= not((layer5_outputs(446)) or (layer5_outputs(4964)));
    layer6_outputs(2359) <= not(layer5_outputs(1124));
    layer6_outputs(2360) <= not(layer5_outputs(1532));
    layer6_outputs(2361) <= layer5_outputs(378);
    layer6_outputs(2362) <= not(layer5_outputs(2439));
    layer6_outputs(2363) <= (layer5_outputs(1262)) xor (layer5_outputs(4362));
    layer6_outputs(2364) <= layer5_outputs(1063);
    layer6_outputs(2365) <= not((layer5_outputs(1810)) xor (layer5_outputs(4382)));
    layer6_outputs(2366) <= layer5_outputs(624);
    layer6_outputs(2367) <= not(layer5_outputs(2841));
    layer6_outputs(2368) <= not(layer5_outputs(5021)) or (layer5_outputs(3354));
    layer6_outputs(2369) <= not((layer5_outputs(1147)) or (layer5_outputs(4293)));
    layer6_outputs(2370) <= not((layer5_outputs(2748)) or (layer5_outputs(2223)));
    layer6_outputs(2371) <= '0';
    layer6_outputs(2372) <= not(layer5_outputs(3157));
    layer6_outputs(2373) <= not(layer5_outputs(3105));
    layer6_outputs(2374) <= layer5_outputs(671);
    layer6_outputs(2375) <= not(layer5_outputs(3958));
    layer6_outputs(2376) <= '1';
    layer6_outputs(2377) <= layer5_outputs(4840);
    layer6_outputs(2378) <= not(layer5_outputs(1790)) or (layer5_outputs(3208));
    layer6_outputs(2379) <= layer5_outputs(4210);
    layer6_outputs(2380) <= layer5_outputs(368);
    layer6_outputs(2381) <= not(layer5_outputs(2229));
    layer6_outputs(2382) <= (layer5_outputs(493)) and not (layer5_outputs(4600));
    layer6_outputs(2383) <= not((layer5_outputs(2152)) xor (layer5_outputs(3345)));
    layer6_outputs(2384) <= layer5_outputs(5028);
    layer6_outputs(2385) <= not((layer5_outputs(3107)) xor (layer5_outputs(4776)));
    layer6_outputs(2386) <= not((layer5_outputs(4596)) and (layer5_outputs(1740)));
    layer6_outputs(2387) <= layer5_outputs(2828);
    layer6_outputs(2388) <= not(layer5_outputs(4362));
    layer6_outputs(2389) <= layer5_outputs(509);
    layer6_outputs(2390) <= layer5_outputs(3958);
    layer6_outputs(2391) <= (layer5_outputs(4269)) xor (layer5_outputs(4863));
    layer6_outputs(2392) <= layer5_outputs(2365);
    layer6_outputs(2393) <= (layer5_outputs(4364)) or (layer5_outputs(3355));
    layer6_outputs(2394) <= not(layer5_outputs(4545));
    layer6_outputs(2395) <= not((layer5_outputs(701)) xor (layer5_outputs(821)));
    layer6_outputs(2396) <= not((layer5_outputs(3105)) or (layer5_outputs(3863)));
    layer6_outputs(2397) <= not(layer5_outputs(2527)) or (layer5_outputs(4356));
    layer6_outputs(2398) <= not(layer5_outputs(761));
    layer6_outputs(2399) <= not(layer5_outputs(2175));
    layer6_outputs(2400) <= layer5_outputs(304);
    layer6_outputs(2401) <= not((layer5_outputs(2526)) xor (layer5_outputs(2525)));
    layer6_outputs(2402) <= (layer5_outputs(875)) xor (layer5_outputs(4845));
    layer6_outputs(2403) <= (layer5_outputs(2715)) and not (layer5_outputs(1776));
    layer6_outputs(2404) <= not(layer5_outputs(2631));
    layer6_outputs(2405) <= (layer5_outputs(2678)) and not (layer5_outputs(2346));
    layer6_outputs(2406) <= not(layer5_outputs(1663)) or (layer5_outputs(2916));
    layer6_outputs(2407) <= layer5_outputs(3331);
    layer6_outputs(2408) <= not(layer5_outputs(2460));
    layer6_outputs(2409) <= not(layer5_outputs(1707)) or (layer5_outputs(4682));
    layer6_outputs(2410) <= not(layer5_outputs(4730));
    layer6_outputs(2411) <= not((layer5_outputs(4526)) or (layer5_outputs(1038)));
    layer6_outputs(2412) <= (layer5_outputs(3322)) and not (layer5_outputs(1195));
    layer6_outputs(2413) <= layer5_outputs(799);
    layer6_outputs(2414) <= not(layer5_outputs(1727));
    layer6_outputs(2415) <= not((layer5_outputs(548)) or (layer5_outputs(1006)));
    layer6_outputs(2416) <= not((layer5_outputs(216)) or (layer5_outputs(1475)));
    layer6_outputs(2417) <= layer5_outputs(587);
    layer6_outputs(2418) <= (layer5_outputs(299)) xor (layer5_outputs(4150));
    layer6_outputs(2419) <= not(layer5_outputs(3511));
    layer6_outputs(2420) <= layer5_outputs(3527);
    layer6_outputs(2421) <= not(layer5_outputs(3098));
    layer6_outputs(2422) <= (layer5_outputs(225)) and not (layer5_outputs(4223));
    layer6_outputs(2423) <= not(layer5_outputs(1945));
    layer6_outputs(2424) <= not(layer5_outputs(1245)) or (layer5_outputs(1400));
    layer6_outputs(2425) <= not(layer5_outputs(112));
    layer6_outputs(2426) <= layer5_outputs(1582);
    layer6_outputs(2427) <= layer5_outputs(2087);
    layer6_outputs(2428) <= '0';
    layer6_outputs(2429) <= (layer5_outputs(220)) xor (layer5_outputs(30));
    layer6_outputs(2430) <= not((layer5_outputs(4884)) xor (layer5_outputs(4523)));
    layer6_outputs(2431) <= layer5_outputs(4744);
    layer6_outputs(2432) <= (layer5_outputs(3387)) and (layer5_outputs(307));
    layer6_outputs(2433) <= not(layer5_outputs(4754)) or (layer5_outputs(1754));
    layer6_outputs(2434) <= layer5_outputs(4882);
    layer6_outputs(2435) <= not((layer5_outputs(4947)) xor (layer5_outputs(2306)));
    layer6_outputs(2436) <= (layer5_outputs(365)) and not (layer5_outputs(4538));
    layer6_outputs(2437) <= not((layer5_outputs(3847)) or (layer5_outputs(2638)));
    layer6_outputs(2438) <= not(layer5_outputs(912));
    layer6_outputs(2439) <= layer5_outputs(3135);
    layer6_outputs(2440) <= not(layer5_outputs(3181));
    layer6_outputs(2441) <= layer5_outputs(1450);
    layer6_outputs(2442) <= not(layer5_outputs(2660)) or (layer5_outputs(3815));
    layer6_outputs(2443) <= not((layer5_outputs(3018)) or (layer5_outputs(255)));
    layer6_outputs(2444) <= not(layer5_outputs(3307));
    layer6_outputs(2445) <= not(layer5_outputs(4750));
    layer6_outputs(2446) <= (layer5_outputs(4571)) and (layer5_outputs(3539));
    layer6_outputs(2447) <= not(layer5_outputs(1528));
    layer6_outputs(2448) <= not(layer5_outputs(1433));
    layer6_outputs(2449) <= not(layer5_outputs(3300)) or (layer5_outputs(2915));
    layer6_outputs(2450) <= not(layer5_outputs(3042));
    layer6_outputs(2451) <= not(layer5_outputs(633)) or (layer5_outputs(3573));
    layer6_outputs(2452) <= (layer5_outputs(3818)) or (layer5_outputs(3962));
    layer6_outputs(2453) <= (layer5_outputs(353)) or (layer5_outputs(1733));
    layer6_outputs(2454) <= layer5_outputs(3310);
    layer6_outputs(2455) <= not(layer5_outputs(3462));
    layer6_outputs(2456) <= (layer5_outputs(4634)) xor (layer5_outputs(2905));
    layer6_outputs(2457) <= not(layer5_outputs(1781));
    layer6_outputs(2458) <= not((layer5_outputs(166)) or (layer5_outputs(4260)));
    layer6_outputs(2459) <= (layer5_outputs(2438)) and (layer5_outputs(4045));
    layer6_outputs(2460) <= not(layer5_outputs(469)) or (layer5_outputs(4182));
    layer6_outputs(2461) <= not(layer5_outputs(4032));
    layer6_outputs(2462) <= not(layer5_outputs(4661)) or (layer5_outputs(2533));
    layer6_outputs(2463) <= not(layer5_outputs(5106));
    layer6_outputs(2464) <= layer5_outputs(1894);
    layer6_outputs(2465) <= not(layer5_outputs(1868));
    layer6_outputs(2466) <= layer5_outputs(4907);
    layer6_outputs(2467) <= not(layer5_outputs(122));
    layer6_outputs(2468) <= (layer5_outputs(3342)) and not (layer5_outputs(1134));
    layer6_outputs(2469) <= not(layer5_outputs(2476));
    layer6_outputs(2470) <= not((layer5_outputs(5023)) and (layer5_outputs(2181)));
    layer6_outputs(2471) <= '0';
    layer6_outputs(2472) <= not(layer5_outputs(1993));
    layer6_outputs(2473) <= not(layer5_outputs(696)) or (layer5_outputs(3454));
    layer6_outputs(2474) <= (layer5_outputs(4310)) xor (layer5_outputs(3224));
    layer6_outputs(2475) <= layer5_outputs(902);
    layer6_outputs(2476) <= layer5_outputs(1232);
    layer6_outputs(2477) <= not(layer5_outputs(3688));
    layer6_outputs(2478) <= not(layer5_outputs(4389));
    layer6_outputs(2479) <= layer5_outputs(947);
    layer6_outputs(2480) <= layer5_outputs(4278);
    layer6_outputs(2481) <= (layer5_outputs(2319)) xor (layer5_outputs(665));
    layer6_outputs(2482) <= not(layer5_outputs(3159));
    layer6_outputs(2483) <= not(layer5_outputs(935));
    layer6_outputs(2484) <= (layer5_outputs(2871)) or (layer5_outputs(3540));
    layer6_outputs(2485) <= (layer5_outputs(2196)) xor (layer5_outputs(2614));
    layer6_outputs(2486) <= (layer5_outputs(4621)) and not (layer5_outputs(3542));
    layer6_outputs(2487) <= not(layer5_outputs(2312));
    layer6_outputs(2488) <= not((layer5_outputs(3786)) and (layer5_outputs(2475)));
    layer6_outputs(2489) <= layer5_outputs(429);
    layer6_outputs(2490) <= not(layer5_outputs(1381));
    layer6_outputs(2491) <= not(layer5_outputs(4861));
    layer6_outputs(2492) <= not(layer5_outputs(3170));
    layer6_outputs(2493) <= not(layer5_outputs(1934));
    layer6_outputs(2494) <= not(layer5_outputs(2598)) or (layer5_outputs(701));
    layer6_outputs(2495) <= not(layer5_outputs(385));
    layer6_outputs(2496) <= not(layer5_outputs(4549));
    layer6_outputs(2497) <= layer5_outputs(4884);
    layer6_outputs(2498) <= not(layer5_outputs(3648));
    layer6_outputs(2499) <= (layer5_outputs(1407)) and not (layer5_outputs(3324));
    layer6_outputs(2500) <= layer5_outputs(2990);
    layer6_outputs(2501) <= (layer5_outputs(2594)) and (layer5_outputs(3378));
    layer6_outputs(2502) <= layer5_outputs(1670);
    layer6_outputs(2503) <= layer5_outputs(2317);
    layer6_outputs(2504) <= (layer5_outputs(4066)) xor (layer5_outputs(2166));
    layer6_outputs(2505) <= layer5_outputs(3259);
    layer6_outputs(2506) <= (layer5_outputs(97)) or (layer5_outputs(182));
    layer6_outputs(2507) <= not(layer5_outputs(491));
    layer6_outputs(2508) <= (layer5_outputs(4098)) and not (layer5_outputs(3857));
    layer6_outputs(2509) <= not(layer5_outputs(3272));
    layer6_outputs(2510) <= not(layer5_outputs(3020)) or (layer5_outputs(604));
    layer6_outputs(2511) <= not(layer5_outputs(2362));
    layer6_outputs(2512) <= layer5_outputs(2579);
    layer6_outputs(2513) <= layer5_outputs(3739);
    layer6_outputs(2514) <= not(layer5_outputs(793));
    layer6_outputs(2515) <= (layer5_outputs(3627)) xor (layer5_outputs(480));
    layer6_outputs(2516) <= not((layer5_outputs(1925)) xor (layer5_outputs(1854)));
    layer6_outputs(2517) <= not(layer5_outputs(1737));
    layer6_outputs(2518) <= not(layer5_outputs(774)) or (layer5_outputs(3127));
    layer6_outputs(2519) <= '0';
    layer6_outputs(2520) <= (layer5_outputs(2966)) and not (layer5_outputs(3137));
    layer6_outputs(2521) <= (layer5_outputs(670)) xor (layer5_outputs(1215));
    layer6_outputs(2522) <= not(layer5_outputs(4368));
    layer6_outputs(2523) <= not(layer5_outputs(2863));
    layer6_outputs(2524) <= layer5_outputs(4853);
    layer6_outputs(2525) <= (layer5_outputs(2513)) and not (layer5_outputs(1173));
    layer6_outputs(2526) <= (layer5_outputs(3348)) and not (layer5_outputs(2520));
    layer6_outputs(2527) <= not(layer5_outputs(2671));
    layer6_outputs(2528) <= (layer5_outputs(4472)) and not (layer5_outputs(3742));
    layer6_outputs(2529) <= layer5_outputs(1755);
    layer6_outputs(2530) <= not(layer5_outputs(1699)) or (layer5_outputs(2975));
    layer6_outputs(2531) <= layer5_outputs(4155);
    layer6_outputs(2532) <= not(layer5_outputs(2964));
    layer6_outputs(2533) <= (layer5_outputs(3843)) xor (layer5_outputs(4871));
    layer6_outputs(2534) <= not(layer5_outputs(4026));
    layer6_outputs(2535) <= (layer5_outputs(3204)) and not (layer5_outputs(5067));
    layer6_outputs(2536) <= not(layer5_outputs(133));
    layer6_outputs(2537) <= (layer5_outputs(2813)) xor (layer5_outputs(258));
    layer6_outputs(2538) <= (layer5_outputs(3449)) xor (layer5_outputs(3204));
    layer6_outputs(2539) <= layer5_outputs(2070);
    layer6_outputs(2540) <= not(layer5_outputs(3395));
    layer6_outputs(2541) <= not(layer5_outputs(2802));
    layer6_outputs(2542) <= layer5_outputs(3453);
    layer6_outputs(2543) <= layer5_outputs(2036);
    layer6_outputs(2544) <= not(layer5_outputs(4091));
    layer6_outputs(2545) <= not(layer5_outputs(4855)) or (layer5_outputs(4229));
    layer6_outputs(2546) <= layer5_outputs(4821);
    layer6_outputs(2547) <= layer5_outputs(3933);
    layer6_outputs(2548) <= layer5_outputs(2657);
    layer6_outputs(2549) <= not(layer5_outputs(690));
    layer6_outputs(2550) <= (layer5_outputs(524)) and not (layer5_outputs(4164));
    layer6_outputs(2551) <= layer5_outputs(1416);
    layer6_outputs(2552) <= layer5_outputs(4049);
    layer6_outputs(2553) <= (layer5_outputs(4398)) and (layer5_outputs(4922));
    layer6_outputs(2554) <= not(layer5_outputs(674));
    layer6_outputs(2555) <= '1';
    layer6_outputs(2556) <= layer5_outputs(3091);
    layer6_outputs(2557) <= (layer5_outputs(3035)) or (layer5_outputs(2284));
    layer6_outputs(2558) <= (layer5_outputs(1207)) or (layer5_outputs(2932));
    layer6_outputs(2559) <= not((layer5_outputs(1703)) and (layer5_outputs(3321)));
    layer6_outputs(2560) <= not(layer5_outputs(1494)) or (layer5_outputs(3810));
    layer6_outputs(2561) <= not(layer5_outputs(75));
    layer6_outputs(2562) <= layer5_outputs(1241);
    layer6_outputs(2563) <= not(layer5_outputs(10));
    layer6_outputs(2564) <= (layer5_outputs(4560)) and (layer5_outputs(2012));
    layer6_outputs(2565) <= not((layer5_outputs(979)) and (layer5_outputs(977)));
    layer6_outputs(2566) <= layer5_outputs(4921);
    layer6_outputs(2567) <= not(layer5_outputs(1138));
    layer6_outputs(2568) <= layer5_outputs(356);
    layer6_outputs(2569) <= layer5_outputs(1505);
    layer6_outputs(2570) <= not(layer5_outputs(1472));
    layer6_outputs(2571) <= not(layer5_outputs(462));
    layer6_outputs(2572) <= layer5_outputs(4550);
    layer6_outputs(2573) <= layer5_outputs(1860);
    layer6_outputs(2574) <= (layer5_outputs(681)) xor (layer5_outputs(3754));
    layer6_outputs(2575) <= not(layer5_outputs(4440));
    layer6_outputs(2576) <= layer5_outputs(1821);
    layer6_outputs(2577) <= (layer5_outputs(3406)) xor (layer5_outputs(2624));
    layer6_outputs(2578) <= layer5_outputs(979);
    layer6_outputs(2579) <= layer5_outputs(4495);
    layer6_outputs(2580) <= (layer5_outputs(939)) and not (layer5_outputs(778));
    layer6_outputs(2581) <= layer5_outputs(1392);
    layer6_outputs(2582) <= not(layer5_outputs(1246));
    layer6_outputs(2583) <= not(layer5_outputs(2112));
    layer6_outputs(2584) <= not((layer5_outputs(4282)) and (layer5_outputs(2930)));
    layer6_outputs(2585) <= layer5_outputs(3377);
    layer6_outputs(2586) <= (layer5_outputs(1183)) and not (layer5_outputs(4474));
    layer6_outputs(2587) <= not(layer5_outputs(516));
    layer6_outputs(2588) <= (layer5_outputs(2053)) or (layer5_outputs(1055));
    layer6_outputs(2589) <= layer5_outputs(3783);
    layer6_outputs(2590) <= not(layer5_outputs(297)) or (layer5_outputs(4620));
    layer6_outputs(2591) <= (layer5_outputs(2554)) or (layer5_outputs(41));
    layer6_outputs(2592) <= layer5_outputs(2237);
    layer6_outputs(2593) <= layer5_outputs(4159);
    layer6_outputs(2594) <= not(layer5_outputs(1045));
    layer6_outputs(2595) <= not((layer5_outputs(4979)) or (layer5_outputs(2668)));
    layer6_outputs(2596) <= not((layer5_outputs(1113)) or (layer5_outputs(1675)));
    layer6_outputs(2597) <= not(layer5_outputs(1488));
    layer6_outputs(2598) <= layer5_outputs(1214);
    layer6_outputs(2599) <= not(layer5_outputs(4759)) or (layer5_outputs(4552));
    layer6_outputs(2600) <= layer5_outputs(400);
    layer6_outputs(2601) <= not(layer5_outputs(1253)) or (layer5_outputs(1019));
    layer6_outputs(2602) <= not(layer5_outputs(2266)) or (layer5_outputs(3175));
    layer6_outputs(2603) <= not(layer5_outputs(4457));
    layer6_outputs(2604) <= layer5_outputs(391);
    layer6_outputs(2605) <= not(layer5_outputs(4280));
    layer6_outputs(2606) <= not((layer5_outputs(848)) xor (layer5_outputs(636)));
    layer6_outputs(2607) <= not(layer5_outputs(1328));
    layer6_outputs(2608) <= not(layer5_outputs(4887));
    layer6_outputs(2609) <= layer5_outputs(4083);
    layer6_outputs(2610) <= (layer5_outputs(1668)) and not (layer5_outputs(764));
    layer6_outputs(2611) <= not(layer5_outputs(3107));
    layer6_outputs(2612) <= not(layer5_outputs(1150));
    layer6_outputs(2613) <= not((layer5_outputs(3058)) or (layer5_outputs(3717)));
    layer6_outputs(2614) <= layer5_outputs(4216);
    layer6_outputs(2615) <= (layer5_outputs(1850)) and (layer5_outputs(2169));
    layer6_outputs(2616) <= not(layer5_outputs(4991));
    layer6_outputs(2617) <= not(layer5_outputs(388));
    layer6_outputs(2618) <= not((layer5_outputs(2141)) or (layer5_outputs(1699)));
    layer6_outputs(2619) <= not(layer5_outputs(4600));
    layer6_outputs(2620) <= not(layer5_outputs(2793));
    layer6_outputs(2621) <= not((layer5_outputs(1912)) and (layer5_outputs(1367)));
    layer6_outputs(2622) <= layer5_outputs(4318);
    layer6_outputs(2623) <= not((layer5_outputs(2061)) xor (layer5_outputs(1114)));
    layer6_outputs(2624) <= not(layer5_outputs(1100));
    layer6_outputs(2625) <= not(layer5_outputs(1313));
    layer6_outputs(2626) <= (layer5_outputs(3079)) xor (layer5_outputs(4682));
    layer6_outputs(2627) <= layer5_outputs(4138);
    layer6_outputs(2628) <= '1';
    layer6_outputs(2629) <= not((layer5_outputs(1534)) or (layer5_outputs(2852)));
    layer6_outputs(2630) <= not(layer5_outputs(4025));
    layer6_outputs(2631) <= not((layer5_outputs(1464)) xor (layer5_outputs(1343)));
    layer6_outputs(2632) <= layer5_outputs(2162);
    layer6_outputs(2633) <= (layer5_outputs(2003)) and not (layer5_outputs(757));
    layer6_outputs(2634) <= not((layer5_outputs(1196)) xor (layer5_outputs(4798)));
    layer6_outputs(2635) <= not(layer5_outputs(4650)) or (layer5_outputs(1365));
    layer6_outputs(2636) <= layer5_outputs(697);
    layer6_outputs(2637) <= (layer5_outputs(4357)) xor (layer5_outputs(1977));
    layer6_outputs(2638) <= layer5_outputs(3272);
    layer6_outputs(2639) <= not(layer5_outputs(1675));
    layer6_outputs(2640) <= not(layer5_outputs(4130));
    layer6_outputs(2641) <= not(layer5_outputs(4127));
    layer6_outputs(2642) <= layer5_outputs(3738);
    layer6_outputs(2643) <= (layer5_outputs(2150)) and (layer5_outputs(3339));
    layer6_outputs(2644) <= (layer5_outputs(1176)) or (layer5_outputs(466));
    layer6_outputs(2645) <= (layer5_outputs(1994)) and not (layer5_outputs(284));
    layer6_outputs(2646) <= not(layer5_outputs(299));
    layer6_outputs(2647) <= (layer5_outputs(4967)) or (layer5_outputs(2320));
    layer6_outputs(2648) <= not(layer5_outputs(2553)) or (layer5_outputs(442));
    layer6_outputs(2649) <= (layer5_outputs(2093)) xor (layer5_outputs(3738));
    layer6_outputs(2650) <= layer5_outputs(249);
    layer6_outputs(2651) <= not(layer5_outputs(4081));
    layer6_outputs(2652) <= not(layer5_outputs(964));
    layer6_outputs(2653) <= '1';
    layer6_outputs(2654) <= (layer5_outputs(1620)) and not (layer5_outputs(1279));
    layer6_outputs(2655) <= not(layer5_outputs(3755));
    layer6_outputs(2656) <= not(layer5_outputs(1680));
    layer6_outputs(2657) <= layer5_outputs(3690);
    layer6_outputs(2658) <= not(layer5_outputs(1815));
    layer6_outputs(2659) <= layer5_outputs(4508);
    layer6_outputs(2660) <= not(layer5_outputs(2289));
    layer6_outputs(2661) <= layer5_outputs(3954);
    layer6_outputs(2662) <= not(layer5_outputs(1420)) or (layer5_outputs(2232));
    layer6_outputs(2663) <= (layer5_outputs(4199)) xor (layer5_outputs(3075));
    layer6_outputs(2664) <= layer5_outputs(522);
    layer6_outputs(2665) <= layer5_outputs(3251);
    layer6_outputs(2666) <= not((layer5_outputs(3662)) and (layer5_outputs(241)));
    layer6_outputs(2667) <= not(layer5_outputs(92));
    layer6_outputs(2668) <= not(layer5_outputs(2505));
    layer6_outputs(2669) <= layer5_outputs(3350);
    layer6_outputs(2670) <= not(layer5_outputs(3408)) or (layer5_outputs(4560));
    layer6_outputs(2671) <= (layer5_outputs(2725)) and (layer5_outputs(243));
    layer6_outputs(2672) <= not((layer5_outputs(487)) and (layer5_outputs(2458)));
    layer6_outputs(2673) <= not(layer5_outputs(4043)) or (layer5_outputs(4136));
    layer6_outputs(2674) <= (layer5_outputs(3126)) and not (layer5_outputs(2070));
    layer6_outputs(2675) <= layer5_outputs(372);
    layer6_outputs(2676) <= layer5_outputs(4748);
    layer6_outputs(2677) <= (layer5_outputs(2997)) and not (layer5_outputs(1765));
    layer6_outputs(2678) <= not((layer5_outputs(3798)) and (layer5_outputs(3249)));
    layer6_outputs(2679) <= layer5_outputs(1954);
    layer6_outputs(2680) <= not(layer5_outputs(234));
    layer6_outputs(2681) <= not(layer5_outputs(549)) or (layer5_outputs(3127));
    layer6_outputs(2682) <= layer5_outputs(602);
    layer6_outputs(2683) <= layer5_outputs(2142);
    layer6_outputs(2684) <= layer5_outputs(510);
    layer6_outputs(2685) <= not(layer5_outputs(3972));
    layer6_outputs(2686) <= not(layer5_outputs(4197));
    layer6_outputs(2687) <= not((layer5_outputs(2491)) or (layer5_outputs(946)));
    layer6_outputs(2688) <= layer5_outputs(2090);
    layer6_outputs(2689) <= layer5_outputs(1906);
    layer6_outputs(2690) <= (layer5_outputs(2178)) xor (layer5_outputs(631));
    layer6_outputs(2691) <= not(layer5_outputs(1540));
    layer6_outputs(2692) <= not(layer5_outputs(3925)) or (layer5_outputs(512));
    layer6_outputs(2693) <= not(layer5_outputs(3867));
    layer6_outputs(2694) <= (layer5_outputs(5001)) xor (layer5_outputs(871));
    layer6_outputs(2695) <= not((layer5_outputs(3840)) xor (layer5_outputs(1223)));
    layer6_outputs(2696) <= not((layer5_outputs(3450)) and (layer5_outputs(4541)));
    layer6_outputs(2697) <= not(layer5_outputs(4431));
    layer6_outputs(2698) <= not(layer5_outputs(2633));
    layer6_outputs(2699) <= not(layer5_outputs(4981));
    layer6_outputs(2700) <= not((layer5_outputs(2847)) and (layer5_outputs(4881)));
    layer6_outputs(2701) <= layer5_outputs(2857);
    layer6_outputs(2702) <= layer5_outputs(282);
    layer6_outputs(2703) <= not((layer5_outputs(5090)) xor (layer5_outputs(2640)));
    layer6_outputs(2704) <= not(layer5_outputs(5114));
    layer6_outputs(2705) <= not((layer5_outputs(1010)) xor (layer5_outputs(4736)));
    layer6_outputs(2706) <= not(layer5_outputs(2901));
    layer6_outputs(2707) <= layer5_outputs(5059);
    layer6_outputs(2708) <= layer5_outputs(899);
    layer6_outputs(2709) <= not(layer5_outputs(2395));
    layer6_outputs(2710) <= not(layer5_outputs(1292));
    layer6_outputs(2711) <= '0';
    layer6_outputs(2712) <= not(layer5_outputs(1323));
    layer6_outputs(2713) <= layer5_outputs(3486);
    layer6_outputs(2714) <= (layer5_outputs(855)) or (layer5_outputs(802));
    layer6_outputs(2715) <= not(layer5_outputs(4941));
    layer6_outputs(2716) <= not(layer5_outputs(443));
    layer6_outputs(2717) <= (layer5_outputs(4356)) and not (layer5_outputs(184));
    layer6_outputs(2718) <= layer5_outputs(3477);
    layer6_outputs(2719) <= layer5_outputs(4312);
    layer6_outputs(2720) <= (layer5_outputs(3070)) and not (layer5_outputs(2923));
    layer6_outputs(2721) <= not((layer5_outputs(1402)) xor (layer5_outputs(2225)));
    layer6_outputs(2722) <= not(layer5_outputs(2290));
    layer6_outputs(2723) <= (layer5_outputs(4426)) xor (layer5_outputs(3670));
    layer6_outputs(2724) <= (layer5_outputs(2215)) and not (layer5_outputs(4361));
    layer6_outputs(2725) <= not(layer5_outputs(1381));
    layer6_outputs(2726) <= layer5_outputs(2252);
    layer6_outputs(2727) <= layer5_outputs(2256);
    layer6_outputs(2728) <= not((layer5_outputs(151)) and (layer5_outputs(4567)));
    layer6_outputs(2729) <= layer5_outputs(742);
    layer6_outputs(2730) <= not(layer5_outputs(1864));
    layer6_outputs(2731) <= not((layer5_outputs(2523)) or (layer5_outputs(4156)));
    layer6_outputs(2732) <= layer5_outputs(1131);
    layer6_outputs(2733) <= layer5_outputs(4998);
    layer6_outputs(2734) <= not((layer5_outputs(4373)) and (layer5_outputs(4080)));
    layer6_outputs(2735) <= not(layer5_outputs(4539));
    layer6_outputs(2736) <= layer5_outputs(4094);
    layer6_outputs(2737) <= not(layer5_outputs(3999));
    layer6_outputs(2738) <= not((layer5_outputs(1069)) and (layer5_outputs(1405)));
    layer6_outputs(2739) <= not(layer5_outputs(178));
    layer6_outputs(2740) <= layer5_outputs(4629);
    layer6_outputs(2741) <= not(layer5_outputs(2890));
    layer6_outputs(2742) <= not(layer5_outputs(5118));
    layer6_outputs(2743) <= not((layer5_outputs(4477)) xor (layer5_outputs(3109)));
    layer6_outputs(2744) <= not(layer5_outputs(538)) or (layer5_outputs(1459));
    layer6_outputs(2745) <= not(layer5_outputs(2119)) or (layer5_outputs(5091));
    layer6_outputs(2746) <= not(layer5_outputs(1092));
    layer6_outputs(2747) <= (layer5_outputs(1018)) or (layer5_outputs(2860));
    layer6_outputs(2748) <= not(layer5_outputs(1171));
    layer6_outputs(2749) <= not(layer5_outputs(750)) or (layer5_outputs(3023));
    layer6_outputs(2750) <= not(layer5_outputs(2933));
    layer6_outputs(2751) <= (layer5_outputs(4793)) and (layer5_outputs(3970));
    layer6_outputs(2752) <= not(layer5_outputs(2538));
    layer6_outputs(2753) <= not(layer5_outputs(3549));
    layer6_outputs(2754) <= not(layer5_outputs(2465));
    layer6_outputs(2755) <= (layer5_outputs(2622)) and (layer5_outputs(889));
    layer6_outputs(2756) <= not(layer5_outputs(3803));
    layer6_outputs(2757) <= not((layer5_outputs(4096)) xor (layer5_outputs(2830)));
    layer6_outputs(2758) <= not(layer5_outputs(3836));
    layer6_outputs(2759) <= not(layer5_outputs(1537));
    layer6_outputs(2760) <= not((layer5_outputs(1811)) and (layer5_outputs(526)));
    layer6_outputs(2761) <= not((layer5_outputs(783)) and (layer5_outputs(3941)));
    layer6_outputs(2762) <= not(layer5_outputs(2039));
    layer6_outputs(2763) <= (layer5_outputs(2161)) and (layer5_outputs(3299));
    layer6_outputs(2764) <= '1';
    layer6_outputs(2765) <= not(layer5_outputs(4674)) or (layer5_outputs(3487));
    layer6_outputs(2766) <= layer5_outputs(1235);
    layer6_outputs(2767) <= layer5_outputs(4877);
    layer6_outputs(2768) <= not(layer5_outputs(980)) or (layer5_outputs(2522));
    layer6_outputs(2769) <= layer5_outputs(3604);
    layer6_outputs(2770) <= not((layer5_outputs(1247)) and (layer5_outputs(4860)));
    layer6_outputs(2771) <= layer5_outputs(5002);
    layer6_outputs(2772) <= layer5_outputs(3162);
    layer6_outputs(2773) <= not(layer5_outputs(4995)) or (layer5_outputs(2297));
    layer6_outputs(2774) <= layer5_outputs(3271);
    layer6_outputs(2775) <= not(layer5_outputs(327)) or (layer5_outputs(1794));
    layer6_outputs(2776) <= not(layer5_outputs(127));
    layer6_outputs(2777) <= (layer5_outputs(1310)) and not (layer5_outputs(918));
    layer6_outputs(2778) <= layer5_outputs(877);
    layer6_outputs(2779) <= (layer5_outputs(2625)) xor (layer5_outputs(3839));
    layer6_outputs(2780) <= (layer5_outputs(3419)) and not (layer5_outputs(2149));
    layer6_outputs(2781) <= (layer5_outputs(5066)) or (layer5_outputs(5074));
    layer6_outputs(2782) <= layer5_outputs(4857);
    layer6_outputs(2783) <= '1';
    layer6_outputs(2784) <= layer5_outputs(575);
    layer6_outputs(2785) <= not(layer5_outputs(4438));
    layer6_outputs(2786) <= not(layer5_outputs(1872));
    layer6_outputs(2787) <= not(layer5_outputs(3416));
    layer6_outputs(2788) <= not(layer5_outputs(4217));
    layer6_outputs(2789) <= not((layer5_outputs(2484)) xor (layer5_outputs(4546)));
    layer6_outputs(2790) <= not((layer5_outputs(285)) xor (layer5_outputs(2862)));
    layer6_outputs(2791) <= not((layer5_outputs(2274)) and (layer5_outputs(4705)));
    layer6_outputs(2792) <= not(layer5_outputs(2892)) or (layer5_outputs(86));
    layer6_outputs(2793) <= not(layer5_outputs(2432));
    layer6_outputs(2794) <= not(layer5_outputs(5086));
    layer6_outputs(2795) <= layer5_outputs(5037);
    layer6_outputs(2796) <= '0';
    layer6_outputs(2797) <= layer5_outputs(5118);
    layer6_outputs(2798) <= not(layer5_outputs(4316));
    layer6_outputs(2799) <= not((layer5_outputs(1032)) xor (layer5_outputs(2720)));
    layer6_outputs(2800) <= layer5_outputs(1238);
    layer6_outputs(2801) <= not(layer5_outputs(2880)) or (layer5_outputs(2414));
    layer6_outputs(2802) <= not(layer5_outputs(1577));
    layer6_outputs(2803) <= (layer5_outputs(5013)) and not (layer5_outputs(48));
    layer6_outputs(2804) <= layer5_outputs(4664);
    layer6_outputs(2805) <= not((layer5_outputs(2261)) or (layer5_outputs(2970)));
    layer6_outputs(2806) <= not(layer5_outputs(2693));
    layer6_outputs(2807) <= not((layer5_outputs(2545)) and (layer5_outputs(4137)));
    layer6_outputs(2808) <= (layer5_outputs(4256)) xor (layer5_outputs(494));
    layer6_outputs(2809) <= not(layer5_outputs(1553));
    layer6_outputs(2810) <= (layer5_outputs(3885)) and not (layer5_outputs(2500));
    layer6_outputs(2811) <= not(layer5_outputs(4668));
    layer6_outputs(2812) <= layer5_outputs(4461);
    layer6_outputs(2813) <= layer5_outputs(3839);
    layer6_outputs(2814) <= layer5_outputs(3242);
    layer6_outputs(2815) <= not((layer5_outputs(297)) xor (layer5_outputs(3798)));
    layer6_outputs(2816) <= layer5_outputs(1822);
    layer6_outputs(2817) <= layer5_outputs(4177);
    layer6_outputs(2818) <= not((layer5_outputs(2751)) xor (layer5_outputs(1915)));
    layer6_outputs(2819) <= layer5_outputs(5095);
    layer6_outputs(2820) <= layer5_outputs(3800);
    layer6_outputs(2821) <= not(layer5_outputs(1091)) or (layer5_outputs(795));
    layer6_outputs(2822) <= not((layer5_outputs(3315)) xor (layer5_outputs(2159)));
    layer6_outputs(2823) <= not(layer5_outputs(3704));
    layer6_outputs(2824) <= not(layer5_outputs(2769));
    layer6_outputs(2825) <= (layer5_outputs(2345)) xor (layer5_outputs(2740));
    layer6_outputs(2826) <= layer5_outputs(14);
    layer6_outputs(2827) <= layer5_outputs(3191);
    layer6_outputs(2828) <= not(layer5_outputs(2251)) or (layer5_outputs(3521));
    layer6_outputs(2829) <= (layer5_outputs(298)) xor (layer5_outputs(4760));
    layer6_outputs(2830) <= layer5_outputs(2542);
    layer6_outputs(2831) <= (layer5_outputs(4844)) xor (layer5_outputs(3497));
    layer6_outputs(2832) <= not(layer5_outputs(14));
    layer6_outputs(2833) <= layer5_outputs(5021);
    layer6_outputs(2834) <= (layer5_outputs(540)) xor (layer5_outputs(1260));
    layer6_outputs(2835) <= not(layer5_outputs(2147));
    layer6_outputs(2836) <= not(layer5_outputs(3541));
    layer6_outputs(2837) <= not(layer5_outputs(703));
    layer6_outputs(2838) <= not(layer5_outputs(881));
    layer6_outputs(2839) <= not(layer5_outputs(4510));
    layer6_outputs(2840) <= (layer5_outputs(4245)) xor (layer5_outputs(4906));
    layer6_outputs(2841) <= layer5_outputs(3337);
    layer6_outputs(2842) <= layer5_outputs(4193);
    layer6_outputs(2843) <= not((layer5_outputs(115)) xor (layer5_outputs(2777)));
    layer6_outputs(2844) <= not(layer5_outputs(2986));
    layer6_outputs(2845) <= layer5_outputs(3972);
    layer6_outputs(2846) <= (layer5_outputs(4723)) and not (layer5_outputs(3088));
    layer6_outputs(2847) <= layer5_outputs(3714);
    layer6_outputs(2848) <= layer5_outputs(2150);
    layer6_outputs(2849) <= not(layer5_outputs(1211));
    layer6_outputs(2850) <= layer5_outputs(3155);
    layer6_outputs(2851) <= not((layer5_outputs(2464)) and (layer5_outputs(3256)));
    layer6_outputs(2852) <= not(layer5_outputs(4522));
    layer6_outputs(2853) <= layer5_outputs(240);
    layer6_outputs(2854) <= layer5_outputs(214);
    layer6_outputs(2855) <= layer5_outputs(4377);
    layer6_outputs(2856) <= not((layer5_outputs(1613)) xor (layer5_outputs(1216)));
    layer6_outputs(2857) <= not(layer5_outputs(4119)) or (layer5_outputs(723));
    layer6_outputs(2858) <= (layer5_outputs(1417)) and not (layer5_outputs(4984));
    layer6_outputs(2859) <= layer5_outputs(3368);
    layer6_outputs(2860) <= layer5_outputs(4394);
    layer6_outputs(2861) <= layer5_outputs(1186);
    layer6_outputs(2862) <= layer5_outputs(4916);
    layer6_outputs(2863) <= not(layer5_outputs(2752));
    layer6_outputs(2864) <= not((layer5_outputs(1372)) xor (layer5_outputs(1120)));
    layer6_outputs(2865) <= not((layer5_outputs(2822)) and (layer5_outputs(571)));
    layer6_outputs(2866) <= not(layer5_outputs(4365));
    layer6_outputs(2867) <= layer5_outputs(2751);
    layer6_outputs(2868) <= not(layer5_outputs(4002));
    layer6_outputs(2869) <= (layer5_outputs(3808)) and not (layer5_outputs(84));
    layer6_outputs(2870) <= not(layer5_outputs(4444));
    layer6_outputs(2871) <= layer5_outputs(3830);
    layer6_outputs(2872) <= (layer5_outputs(2730)) and not (layer5_outputs(582));
    layer6_outputs(2873) <= not((layer5_outputs(1156)) or (layer5_outputs(9)));
    layer6_outputs(2874) <= layer5_outputs(4381);
    layer6_outputs(2875) <= '1';
    layer6_outputs(2876) <= (layer5_outputs(16)) and not (layer5_outputs(1194));
    layer6_outputs(2877) <= not((layer5_outputs(18)) xor (layer5_outputs(1481)));
    layer6_outputs(2878) <= not((layer5_outputs(3966)) xor (layer5_outputs(431)));
    layer6_outputs(2879) <= (layer5_outputs(3895)) and not (layer5_outputs(219));
    layer6_outputs(2880) <= layer5_outputs(4453);
    layer6_outputs(2881) <= not(layer5_outputs(2535));
    layer6_outputs(2882) <= '1';
    layer6_outputs(2883) <= layer5_outputs(4725);
    layer6_outputs(2884) <= (layer5_outputs(1747)) xor (layer5_outputs(3385));
    layer6_outputs(2885) <= layer5_outputs(2132);
    layer6_outputs(2886) <= not(layer5_outputs(3199));
    layer6_outputs(2887) <= (layer5_outputs(3072)) and (layer5_outputs(3379));
    layer6_outputs(2888) <= not(layer5_outputs(3927));
    layer6_outputs(2889) <= not(layer5_outputs(679));
    layer6_outputs(2890) <= not(layer5_outputs(1131)) or (layer5_outputs(518));
    layer6_outputs(2891) <= not((layer5_outputs(2510)) or (layer5_outputs(3268)));
    layer6_outputs(2892) <= not(layer5_outputs(3801)) or (layer5_outputs(1269));
    layer6_outputs(2893) <= layer5_outputs(1643);
    layer6_outputs(2894) <= not(layer5_outputs(3310));
    layer6_outputs(2895) <= not(layer5_outputs(455));
    layer6_outputs(2896) <= (layer5_outputs(4407)) xor (layer5_outputs(4300));
    layer6_outputs(2897) <= not(layer5_outputs(3357));
    layer6_outputs(2898) <= layer5_outputs(4740);
    layer6_outputs(2899) <= layer5_outputs(222);
    layer6_outputs(2900) <= (layer5_outputs(2914)) xor (layer5_outputs(3762));
    layer6_outputs(2901) <= layer5_outputs(168);
    layer6_outputs(2902) <= not(layer5_outputs(915));
    layer6_outputs(2903) <= layer5_outputs(4041);
    layer6_outputs(2904) <= not(layer5_outputs(737));
    layer6_outputs(2905) <= layer5_outputs(4638);
    layer6_outputs(2906) <= not(layer5_outputs(3869));
    layer6_outputs(2907) <= not(layer5_outputs(1442));
    layer6_outputs(2908) <= not((layer5_outputs(4516)) xor (layer5_outputs(1827)));
    layer6_outputs(2909) <= not(layer5_outputs(4433)) or (layer5_outputs(520));
    layer6_outputs(2910) <= (layer5_outputs(791)) and not (layer5_outputs(1570));
    layer6_outputs(2911) <= '1';
    layer6_outputs(2912) <= (layer5_outputs(3689)) and not (layer5_outputs(2909));
    layer6_outputs(2913) <= layer5_outputs(1144);
    layer6_outputs(2914) <= layer5_outputs(799);
    layer6_outputs(2915) <= not(layer5_outputs(4067));
    layer6_outputs(2916) <= layer5_outputs(3677);
    layer6_outputs(2917) <= not((layer5_outputs(1393)) and (layer5_outputs(4180)));
    layer6_outputs(2918) <= not((layer5_outputs(3367)) or (layer5_outputs(2840)));
    layer6_outputs(2919) <= layer5_outputs(3014);
    layer6_outputs(2920) <= (layer5_outputs(3350)) xor (layer5_outputs(1698));
    layer6_outputs(2921) <= not(layer5_outputs(2009));
    layer6_outputs(2922) <= (layer5_outputs(996)) and not (layer5_outputs(3011));
    layer6_outputs(2923) <= not((layer5_outputs(1184)) xor (layer5_outputs(2919)));
    layer6_outputs(2924) <= layer5_outputs(525);
    layer6_outputs(2925) <= not(layer5_outputs(1518));
    layer6_outputs(2926) <= (layer5_outputs(911)) and not (layer5_outputs(628));
    layer6_outputs(2927) <= layer5_outputs(3985);
    layer6_outputs(2928) <= not(layer5_outputs(1673));
    layer6_outputs(2929) <= layer5_outputs(3694);
    layer6_outputs(2930) <= (layer5_outputs(2443)) xor (layer5_outputs(3021));
    layer6_outputs(2931) <= layer5_outputs(158);
    layer6_outputs(2932) <= not(layer5_outputs(3397));
    layer6_outputs(2933) <= not(layer5_outputs(4948));
    layer6_outputs(2934) <= layer5_outputs(312);
    layer6_outputs(2935) <= (layer5_outputs(2873)) and (layer5_outputs(3816));
    layer6_outputs(2936) <= not(layer5_outputs(201));
    layer6_outputs(2937) <= not(layer5_outputs(3929));
    layer6_outputs(2938) <= not(layer5_outputs(4524));
    layer6_outputs(2939) <= layer5_outputs(955);
    layer6_outputs(2940) <= not((layer5_outputs(4951)) and (layer5_outputs(3948)));
    layer6_outputs(2941) <= not(layer5_outputs(1571));
    layer6_outputs(2942) <= (layer5_outputs(1449)) and (layer5_outputs(178));
    layer6_outputs(2943) <= not(layer5_outputs(4425));
    layer6_outputs(2944) <= layer5_outputs(4531);
    layer6_outputs(2945) <= not(layer5_outputs(4474));
    layer6_outputs(2946) <= not(layer5_outputs(764));
    layer6_outputs(2947) <= (layer5_outputs(2380)) and not (layer5_outputs(2324));
    layer6_outputs(2948) <= '1';
    layer6_outputs(2949) <= not(layer5_outputs(2883));
    layer6_outputs(2950) <= not((layer5_outputs(1236)) xor (layer5_outputs(4722)));
    layer6_outputs(2951) <= layer5_outputs(2935);
    layer6_outputs(2952) <= (layer5_outputs(2293)) or (layer5_outputs(1974));
    layer6_outputs(2953) <= not((layer5_outputs(589)) or (layer5_outputs(2168)));
    layer6_outputs(2954) <= (layer5_outputs(3172)) and not (layer5_outputs(1404));
    layer6_outputs(2955) <= (layer5_outputs(4424)) and (layer5_outputs(1419));
    layer6_outputs(2956) <= (layer5_outputs(3585)) xor (layer5_outputs(1546));
    layer6_outputs(2957) <= layer5_outputs(2230);
    layer6_outputs(2958) <= (layer5_outputs(2786)) xor (layer5_outputs(2138));
    layer6_outputs(2959) <= not(layer5_outputs(2738)) or (layer5_outputs(3244));
    layer6_outputs(2960) <= not(layer5_outputs(4866));
    layer6_outputs(2961) <= not(layer5_outputs(4337));
    layer6_outputs(2962) <= not(layer5_outputs(769));
    layer6_outputs(2963) <= (layer5_outputs(2207)) xor (layer5_outputs(864));
    layer6_outputs(2964) <= not((layer5_outputs(1728)) or (layer5_outputs(379)));
    layer6_outputs(2965) <= not(layer5_outputs(1792));
    layer6_outputs(2966) <= (layer5_outputs(1083)) and (layer5_outputs(5116));
    layer6_outputs(2967) <= not((layer5_outputs(4918)) and (layer5_outputs(1163)));
    layer6_outputs(2968) <= layer5_outputs(1224);
    layer6_outputs(2969) <= layer5_outputs(1);
    layer6_outputs(2970) <= not(layer5_outputs(2315));
    layer6_outputs(2971) <= layer5_outputs(4675);
    layer6_outputs(2972) <= not(layer5_outputs(2135));
    layer6_outputs(2973) <= not(layer5_outputs(4966));
    layer6_outputs(2974) <= not(layer5_outputs(2382));
    layer6_outputs(2975) <= (layer5_outputs(468)) xor (layer5_outputs(932));
    layer6_outputs(2976) <= layer5_outputs(4236);
    layer6_outputs(2977) <= not(layer5_outputs(442));
    layer6_outputs(2978) <= not(layer5_outputs(4168));
    layer6_outputs(2979) <= layer5_outputs(1427);
    layer6_outputs(2980) <= layer5_outputs(24);
    layer6_outputs(2981) <= not((layer5_outputs(3317)) xor (layer5_outputs(3)));
    layer6_outputs(2982) <= layer5_outputs(150);
    layer6_outputs(2983) <= layer5_outputs(2976);
    layer6_outputs(2984) <= not((layer5_outputs(3828)) or (layer5_outputs(1036)));
    layer6_outputs(2985) <= (layer5_outputs(4670)) and not (layer5_outputs(363));
    layer6_outputs(2986) <= layer5_outputs(4583);
    layer6_outputs(2987) <= not(layer5_outputs(2783));
    layer6_outputs(2988) <= not((layer5_outputs(4859)) xor (layer5_outputs(2205)));
    layer6_outputs(2989) <= not(layer5_outputs(3234));
    layer6_outputs(2990) <= not(layer5_outputs(248));
    layer6_outputs(2991) <= (layer5_outputs(2250)) and (layer5_outputs(373));
    layer6_outputs(2992) <= not(layer5_outputs(4058)) or (layer5_outputs(1698));
    layer6_outputs(2993) <= not((layer5_outputs(1389)) and (layer5_outputs(2188)));
    layer6_outputs(2994) <= not(layer5_outputs(5000));
    layer6_outputs(2995) <= layer5_outputs(2833);
    layer6_outputs(2996) <= layer5_outputs(3708);
    layer6_outputs(2997) <= not(layer5_outputs(1096));
    layer6_outputs(2998) <= (layer5_outputs(846)) xor (layer5_outputs(4728));
    layer6_outputs(2999) <= not((layer5_outputs(3084)) xor (layer5_outputs(2981)));
    layer6_outputs(3000) <= layer5_outputs(2805);
    layer6_outputs(3001) <= layer5_outputs(1111);
    layer6_outputs(3002) <= (layer5_outputs(2254)) and (layer5_outputs(3852));
    layer6_outputs(3003) <= (layer5_outputs(3138)) and (layer5_outputs(2255));
    layer6_outputs(3004) <= layer5_outputs(2458);
    layer6_outputs(3005) <= not(layer5_outputs(1414));
    layer6_outputs(3006) <= (layer5_outputs(3099)) xor (layer5_outputs(1794));
    layer6_outputs(3007) <= not(layer5_outputs(4780));
    layer6_outputs(3008) <= layer5_outputs(4564);
    layer6_outputs(3009) <= not(layer5_outputs(3252));
    layer6_outputs(3010) <= (layer5_outputs(3653)) and (layer5_outputs(3605));
    layer6_outputs(3011) <= not(layer5_outputs(2280)) or (layer5_outputs(1317));
    layer6_outputs(3012) <= layer5_outputs(4359);
    layer6_outputs(3013) <= (layer5_outputs(4822)) and (layer5_outputs(4286));
    layer6_outputs(3014) <= not(layer5_outputs(1578));
    layer6_outputs(3015) <= not(layer5_outputs(371));
    layer6_outputs(3016) <= layer5_outputs(2643);
    layer6_outputs(3017) <= layer5_outputs(3919);
    layer6_outputs(3018) <= (layer5_outputs(3514)) and not (layer5_outputs(4899));
    layer6_outputs(3019) <= not(layer5_outputs(3894));
    layer6_outputs(3020) <= not(layer5_outputs(1024));
    layer6_outputs(3021) <= layer5_outputs(4352);
    layer6_outputs(3022) <= (layer5_outputs(1513)) and not (layer5_outputs(4946));
    layer6_outputs(3023) <= not((layer5_outputs(476)) or (layer5_outputs(1600)));
    layer6_outputs(3024) <= layer5_outputs(1782);
    layer6_outputs(3025) <= not(layer5_outputs(12));
    layer6_outputs(3026) <= (layer5_outputs(4132)) or (layer5_outputs(728));
    layer6_outputs(3027) <= (layer5_outputs(4652)) and not (layer5_outputs(2095));
    layer6_outputs(3028) <= not((layer5_outputs(4021)) and (layer5_outputs(1189)));
    layer6_outputs(3029) <= not((layer5_outputs(3661)) and (layer5_outputs(3874)));
    layer6_outputs(3030) <= layer5_outputs(2519);
    layer6_outputs(3031) <= not(layer5_outputs(3868));
    layer6_outputs(3032) <= not(layer5_outputs(2387));
    layer6_outputs(3033) <= not(layer5_outputs(2699));
    layer6_outputs(3034) <= layer5_outputs(4669);
    layer6_outputs(3035) <= (layer5_outputs(4706)) and (layer5_outputs(2311));
    layer6_outputs(3036) <= (layer5_outputs(3758)) or (layer5_outputs(4275));
    layer6_outputs(3037) <= '1';
    layer6_outputs(3038) <= not((layer5_outputs(4380)) xor (layer5_outputs(3672)));
    layer6_outputs(3039) <= layer5_outputs(1788);
    layer6_outputs(3040) <= not(layer5_outputs(4428));
    layer6_outputs(3041) <= not(layer5_outputs(2744));
    layer6_outputs(3042) <= not((layer5_outputs(435)) and (layer5_outputs(3468)));
    layer6_outputs(3043) <= not((layer5_outputs(3523)) and (layer5_outputs(4331)));
    layer6_outputs(3044) <= (layer5_outputs(2840)) and (layer5_outputs(1732));
    layer6_outputs(3045) <= layer5_outputs(3533);
    layer6_outputs(3046) <= not(layer5_outputs(895)) or (layer5_outputs(2243));
    layer6_outputs(3047) <= (layer5_outputs(1135)) xor (layer5_outputs(480));
    layer6_outputs(3048) <= not(layer5_outputs(2309));
    layer6_outputs(3049) <= not(layer5_outputs(4078)) or (layer5_outputs(1585));
    layer6_outputs(3050) <= layer5_outputs(1955);
    layer6_outputs(3051) <= layer5_outputs(3043);
    layer6_outputs(3052) <= (layer5_outputs(2299)) xor (layer5_outputs(4605));
    layer6_outputs(3053) <= layer5_outputs(1657);
    layer6_outputs(3054) <= not(layer5_outputs(2917));
    layer6_outputs(3055) <= not((layer5_outputs(3797)) xor (layer5_outputs(1369)));
    layer6_outputs(3056) <= (layer5_outputs(4221)) and not (layer5_outputs(4983));
    layer6_outputs(3057) <= not(layer5_outputs(2542)) or (layer5_outputs(95));
    layer6_outputs(3058) <= layer5_outputs(3275);
    layer6_outputs(3059) <= not(layer5_outputs(923));
    layer6_outputs(3060) <= not(layer5_outputs(5112));
    layer6_outputs(3061) <= not(layer5_outputs(2295));
    layer6_outputs(3062) <= not(layer5_outputs(4244)) or (layer5_outputs(619));
    layer6_outputs(3063) <= not(layer5_outputs(4489)) or (layer5_outputs(328));
    layer6_outputs(3064) <= layer5_outputs(1068);
    layer6_outputs(3065) <= layer5_outputs(2123);
    layer6_outputs(3066) <= layer5_outputs(2842);
    layer6_outputs(3067) <= layer5_outputs(4209);
    layer6_outputs(3068) <= layer5_outputs(20);
    layer6_outputs(3069) <= layer5_outputs(3655);
    layer6_outputs(3070) <= layer5_outputs(903);
    layer6_outputs(3071) <= not((layer5_outputs(768)) xor (layer5_outputs(4454)));
    layer6_outputs(3072) <= layer5_outputs(2371);
    layer6_outputs(3073) <= (layer5_outputs(1373)) and not (layer5_outputs(4909));
    layer6_outputs(3074) <= (layer5_outputs(2067)) and (layer5_outputs(4594));
    layer6_outputs(3075) <= not(layer5_outputs(4673));
    layer6_outputs(3076) <= not(layer5_outputs(1884));
    layer6_outputs(3077) <= not(layer5_outputs(852));
    layer6_outputs(3078) <= not(layer5_outputs(1294));
    layer6_outputs(3079) <= not((layer5_outputs(1258)) xor (layer5_outputs(386)));
    layer6_outputs(3080) <= (layer5_outputs(3989)) and not (layer5_outputs(2640));
    layer6_outputs(3081) <= (layer5_outputs(4225)) xor (layer5_outputs(2766));
    layer6_outputs(3082) <= not(layer5_outputs(4678)) or (layer5_outputs(1107));
    layer6_outputs(3083) <= layer5_outputs(2883);
    layer6_outputs(3084) <= layer5_outputs(1125);
    layer6_outputs(3085) <= not(layer5_outputs(4021));
    layer6_outputs(3086) <= not((layer5_outputs(1282)) xor (layer5_outputs(4249)));
    layer6_outputs(3087) <= not((layer5_outputs(3311)) xor (layer5_outputs(4568)));
    layer6_outputs(3088) <= not((layer5_outputs(2367)) xor (layer5_outputs(3228)));
    layer6_outputs(3089) <= layer5_outputs(2848);
    layer6_outputs(3090) <= not(layer5_outputs(2733)) or (layer5_outputs(2882));
    layer6_outputs(3091) <= not(layer5_outputs(4497));
    layer6_outputs(3092) <= not(layer5_outputs(1347));
    layer6_outputs(3093) <= not(layer5_outputs(4828));
    layer6_outputs(3094) <= layer5_outputs(3447);
    layer6_outputs(3095) <= (layer5_outputs(1784)) xor (layer5_outputs(2436));
    layer6_outputs(3096) <= not(layer5_outputs(4901));
    layer6_outputs(3097) <= not(layer5_outputs(588));
    layer6_outputs(3098) <= not((layer5_outputs(5032)) or (layer5_outputs(3955)));
    layer6_outputs(3099) <= not(layer5_outputs(2141));
    layer6_outputs(3100) <= (layer5_outputs(4517)) xor (layer5_outputs(2144));
    layer6_outputs(3101) <= not((layer5_outputs(2161)) xor (layer5_outputs(181)));
    layer6_outputs(3102) <= (layer5_outputs(426)) and (layer5_outputs(1257));
    layer6_outputs(3103) <= (layer5_outputs(2404)) xor (layer5_outputs(3492));
    layer6_outputs(3104) <= (layer5_outputs(4088)) and (layer5_outputs(129));
    layer6_outputs(3105) <= layer5_outputs(2384);
    layer6_outputs(3106) <= not(layer5_outputs(1423));
    layer6_outputs(3107) <= not((layer5_outputs(3550)) xor (layer5_outputs(3092)));
    layer6_outputs(3108) <= not(layer5_outputs(3372));
    layer6_outputs(3109) <= not(layer5_outputs(1039)) or (layer5_outputs(1022));
    layer6_outputs(3110) <= not(layer5_outputs(1732)) or (layer5_outputs(2710));
    layer6_outputs(3111) <= layer5_outputs(4907);
    layer6_outputs(3112) <= layer5_outputs(645);
    layer6_outputs(3113) <= not(layer5_outputs(2220));
    layer6_outputs(3114) <= not(layer5_outputs(1117)) or (layer5_outputs(2441));
    layer6_outputs(3115) <= (layer5_outputs(4521)) xor (layer5_outputs(1221));
    layer6_outputs(3116) <= not(layer5_outputs(3803));
    layer6_outputs(3117) <= not(layer5_outputs(3851));
    layer6_outputs(3118) <= (layer5_outputs(1980)) and not (layer5_outputs(4290));
    layer6_outputs(3119) <= not((layer5_outputs(3210)) and (layer5_outputs(4829)));
    layer6_outputs(3120) <= layer5_outputs(2785);
    layer6_outputs(3121) <= layer5_outputs(337);
    layer6_outputs(3122) <= not(layer5_outputs(2982));
    layer6_outputs(3123) <= not((layer5_outputs(4226)) xor (layer5_outputs(1664)));
    layer6_outputs(3124) <= (layer5_outputs(4005)) and not (layer5_outputs(3957));
    layer6_outputs(3125) <= layer5_outputs(4582);
    layer6_outputs(3126) <= not(layer5_outputs(1345));
    layer6_outputs(3127) <= not(layer5_outputs(4198));
    layer6_outputs(3128) <= not(layer5_outputs(4460));
    layer6_outputs(3129) <= layer5_outputs(5050);
    layer6_outputs(3130) <= not(layer5_outputs(4960));
    layer6_outputs(3131) <= not(layer5_outputs(3866));
    layer6_outputs(3132) <= not((layer5_outputs(4492)) xor (layer5_outputs(3265)));
    layer6_outputs(3133) <= not(layer5_outputs(2426));
    layer6_outputs(3134) <= layer5_outputs(1493);
    layer6_outputs(3135) <= layer5_outputs(2978);
    layer6_outputs(3136) <= layer5_outputs(3465);
    layer6_outputs(3137) <= not((layer5_outputs(251)) or (layer5_outputs(1893)));
    layer6_outputs(3138) <= layer5_outputs(2190);
    layer6_outputs(3139) <= layer5_outputs(3955);
    layer6_outputs(3140) <= not(layer5_outputs(3796));
    layer6_outputs(3141) <= not((layer5_outputs(174)) or (layer5_outputs(1190)));
    layer6_outputs(3142) <= layer5_outputs(3820);
    layer6_outputs(3143) <= (layer5_outputs(4794)) xor (layer5_outputs(5117));
    layer6_outputs(3144) <= layer5_outputs(566);
    layer6_outputs(3145) <= layer5_outputs(2449);
    layer6_outputs(3146) <= not(layer5_outputs(2427));
    layer6_outputs(3147) <= (layer5_outputs(4708)) xor (layer5_outputs(1967));
    layer6_outputs(3148) <= not(layer5_outputs(4505));
    layer6_outputs(3149) <= not(layer5_outputs(4897));
    layer6_outputs(3150) <= (layer5_outputs(1859)) and not (layer5_outputs(3175));
    layer6_outputs(3151) <= not(layer5_outputs(4773));
    layer6_outputs(3152) <= not(layer5_outputs(2055));
    layer6_outputs(3153) <= layer5_outputs(2308);
    layer6_outputs(3154) <= (layer5_outputs(1935)) or (layer5_outputs(3602));
    layer6_outputs(3155) <= not(layer5_outputs(4330));
    layer6_outputs(3156) <= '0';
    layer6_outputs(3157) <= (layer5_outputs(3480)) xor (layer5_outputs(4181));
    layer6_outputs(3158) <= '1';
    layer6_outputs(3159) <= (layer5_outputs(1768)) and (layer5_outputs(2410));
    layer6_outputs(3160) <= layer5_outputs(4817);
    layer6_outputs(3161) <= not(layer5_outputs(2716));
    layer6_outputs(3162) <= (layer5_outputs(2704)) and not (layer5_outputs(1243));
    layer6_outputs(3163) <= (layer5_outputs(2364)) or (layer5_outputs(3874));
    layer6_outputs(3164) <= '1';
    layer6_outputs(3165) <= not(layer5_outputs(4312));
    layer6_outputs(3166) <= not(layer5_outputs(2312));
    layer6_outputs(3167) <= layer5_outputs(2808);
    layer6_outputs(3168) <= (layer5_outputs(1647)) or (layer5_outputs(1182));
    layer6_outputs(3169) <= not(layer5_outputs(3236));
    layer6_outputs(3170) <= layer5_outputs(1743);
    layer6_outputs(3171) <= not((layer5_outputs(2214)) and (layer5_outputs(618)));
    layer6_outputs(3172) <= not(layer5_outputs(3507)) or (layer5_outputs(3607));
    layer6_outputs(3173) <= (layer5_outputs(2807)) and (layer5_outputs(1168));
    layer6_outputs(3174) <= not(layer5_outputs(1388));
    layer6_outputs(3175) <= layer5_outputs(2682);
    layer6_outputs(3176) <= not(layer5_outputs(3211));
    layer6_outputs(3177) <= layer5_outputs(3057);
    layer6_outputs(3178) <= layer5_outputs(2994);
    layer6_outputs(3179) <= not((layer5_outputs(3062)) or (layer5_outputs(4421)));
    layer6_outputs(3180) <= layer5_outputs(2673);
    layer6_outputs(3181) <= not(layer5_outputs(4361));
    layer6_outputs(3182) <= not(layer5_outputs(325));
    layer6_outputs(3183) <= not(layer5_outputs(2759));
    layer6_outputs(3184) <= not(layer5_outputs(747)) or (layer5_outputs(4116));
    layer6_outputs(3185) <= (layer5_outputs(2671)) and (layer5_outputs(4434));
    layer6_outputs(3186) <= not((layer5_outputs(3701)) and (layer5_outputs(4642)));
    layer6_outputs(3187) <= not(layer5_outputs(4731));
    layer6_outputs(3188) <= layer5_outputs(2360);
    layer6_outputs(3189) <= (layer5_outputs(2372)) and not (layer5_outputs(3960));
    layer6_outputs(3190) <= (layer5_outputs(3852)) and not (layer5_outputs(1004));
    layer6_outputs(3191) <= not(layer5_outputs(2591));
    layer6_outputs(3192) <= layer5_outputs(4443);
    layer6_outputs(3193) <= layer5_outputs(574);
    layer6_outputs(3194) <= layer5_outputs(1736);
    layer6_outputs(3195) <= (layer5_outputs(4458)) and not (layer5_outputs(545));
    layer6_outputs(3196) <= not(layer5_outputs(3026));
    layer6_outputs(3197) <= not((layer5_outputs(4305)) and (layer5_outputs(82)));
    layer6_outputs(3198) <= (layer5_outputs(2864)) or (layer5_outputs(3713));
    layer6_outputs(3199) <= not(layer5_outputs(597));
    layer6_outputs(3200) <= not((layer5_outputs(2286)) xor (layer5_outputs(874)));
    layer6_outputs(3201) <= layer5_outputs(1395);
    layer6_outputs(3202) <= not(layer5_outputs(3795)) or (layer5_outputs(483));
    layer6_outputs(3203) <= not(layer5_outputs(1819)) or (layer5_outputs(4863));
    layer6_outputs(3204) <= layer5_outputs(599);
    layer6_outputs(3205) <= (layer5_outputs(1548)) and not (layer5_outputs(2352));
    layer6_outputs(3206) <= not(layer5_outputs(3140));
    layer6_outputs(3207) <= not(layer5_outputs(1014));
    layer6_outputs(3208) <= not(layer5_outputs(1833));
    layer6_outputs(3209) <= layer5_outputs(4528);
    layer6_outputs(3210) <= not(layer5_outputs(1778));
    layer6_outputs(3211) <= not((layer5_outputs(2022)) or (layer5_outputs(310)));
    layer6_outputs(3212) <= not(layer5_outputs(713));
    layer6_outputs(3213) <= not(layer5_outputs(1972));
    layer6_outputs(3214) <= not(layer5_outputs(3851));
    layer6_outputs(3215) <= layer5_outputs(4853);
    layer6_outputs(3216) <= not((layer5_outputs(357)) or (layer5_outputs(963)));
    layer6_outputs(3217) <= not(layer5_outputs(4835));
    layer6_outputs(3218) <= not(layer5_outputs(2836));
    layer6_outputs(3219) <= (layer5_outputs(4065)) and (layer5_outputs(615));
    layer6_outputs(3220) <= layer5_outputs(3316);
    layer6_outputs(3221) <= not(layer5_outputs(3482)) or (layer5_outputs(4555));
    layer6_outputs(3222) <= (layer5_outputs(843)) xor (layer5_outputs(477));
    layer6_outputs(3223) <= layer5_outputs(4645);
    layer6_outputs(3224) <= layer5_outputs(4856);
    layer6_outputs(3225) <= not(layer5_outputs(941));
    layer6_outputs(3226) <= not((layer5_outputs(2194)) and (layer5_outputs(8)));
    layer6_outputs(3227) <= not(layer5_outputs(2714));
    layer6_outputs(3228) <= (layer5_outputs(3349)) xor (layer5_outputs(4487));
    layer6_outputs(3229) <= layer5_outputs(3015);
    layer6_outputs(3230) <= (layer5_outputs(395)) xor (layer5_outputs(3197));
    layer6_outputs(3231) <= not(layer5_outputs(449));
    layer6_outputs(3232) <= (layer5_outputs(527)) xor (layer5_outputs(2024));
    layer6_outputs(3233) <= layer5_outputs(3194);
    layer6_outputs(3234) <= (layer5_outputs(4976)) and not (layer5_outputs(3415));
    layer6_outputs(3235) <= (layer5_outputs(206)) and not (layer5_outputs(2182));
    layer6_outputs(3236) <= not(layer5_outputs(2936));
    layer6_outputs(3237) <= not((layer5_outputs(1036)) and (layer5_outputs(3004)));
    layer6_outputs(3238) <= (layer5_outputs(4172)) and (layer5_outputs(891));
    layer6_outputs(3239) <= not(layer5_outputs(2961)) or (layer5_outputs(3428));
    layer6_outputs(3240) <= layer5_outputs(2349);
    layer6_outputs(3241) <= layer5_outputs(111);
    layer6_outputs(3242) <= layer5_outputs(3196);
    layer6_outputs(3243) <= not(layer5_outputs(1182));
    layer6_outputs(3244) <= not(layer5_outputs(2370)) or (layer5_outputs(3559));
    layer6_outputs(3245) <= not((layer5_outputs(44)) xor (layer5_outputs(1383)));
    layer6_outputs(3246) <= layer5_outputs(172);
    layer6_outputs(3247) <= (layer5_outputs(4326)) xor (layer5_outputs(3730));
    layer6_outputs(3248) <= not(layer5_outputs(3615));
    layer6_outputs(3249) <= (layer5_outputs(573)) and (layer5_outputs(2572));
    layer6_outputs(3250) <= not(layer5_outputs(3823));
    layer6_outputs(3251) <= layer5_outputs(590);
    layer6_outputs(3252) <= not(layer5_outputs(1922)) or (layer5_outputs(1989));
    layer6_outputs(3253) <= '0';
    layer6_outputs(3254) <= not((layer5_outputs(899)) xor (layer5_outputs(1748)));
    layer6_outputs(3255) <= layer5_outputs(1677);
    layer6_outputs(3256) <= layer5_outputs(349);
    layer6_outputs(3257) <= (layer5_outputs(302)) or (layer5_outputs(873));
    layer6_outputs(3258) <= (layer5_outputs(4566)) and (layer5_outputs(626));
    layer6_outputs(3259) <= not(layer5_outputs(382));
    layer6_outputs(3260) <= layer5_outputs(367);
    layer6_outputs(3261) <= not(layer5_outputs(3072));
    layer6_outputs(3262) <= (layer5_outputs(439)) and not (layer5_outputs(2377));
    layer6_outputs(3263) <= (layer5_outputs(1587)) and not (layer5_outputs(3630));
    layer6_outputs(3264) <= not((layer5_outputs(3158)) and (layer5_outputs(4923)));
    layer6_outputs(3265) <= (layer5_outputs(3943)) and (layer5_outputs(2218));
    layer6_outputs(3266) <= layer5_outputs(1710);
    layer6_outputs(3267) <= not(layer5_outputs(4079)) or (layer5_outputs(3896));
    layer6_outputs(3268) <= layer5_outputs(4739);
    layer6_outputs(3269) <= (layer5_outputs(2339)) and not (layer5_outputs(1717));
    layer6_outputs(3270) <= not(layer5_outputs(1348)) or (layer5_outputs(4683));
    layer6_outputs(3271) <= layer5_outputs(144);
    layer6_outputs(3272) <= not(layer5_outputs(906));
    layer6_outputs(3273) <= layer5_outputs(1641);
    layer6_outputs(3274) <= layer5_outputs(4484);
    layer6_outputs(3275) <= not(layer5_outputs(506));
    layer6_outputs(3276) <= (layer5_outputs(2390)) and not (layer5_outputs(2318));
    layer6_outputs(3277) <= layer5_outputs(4238);
    layer6_outputs(3278) <= not(layer5_outputs(3009));
    layer6_outputs(3279) <= layer5_outputs(457);
    layer6_outputs(3280) <= layer5_outputs(388);
    layer6_outputs(3281) <= layer5_outputs(2004);
    layer6_outputs(3282) <= not(layer5_outputs(1004)) or (layer5_outputs(3777));
    layer6_outputs(3283) <= layer5_outputs(1953);
    layer6_outputs(3284) <= layer5_outputs(4141);
    layer6_outputs(3285) <= layer5_outputs(1586);
    layer6_outputs(3286) <= not(layer5_outputs(1667)) or (layer5_outputs(4084));
    layer6_outputs(3287) <= (layer5_outputs(4493)) and not (layer5_outputs(4976));
    layer6_outputs(3288) <= not(layer5_outputs(4949));
    layer6_outputs(3289) <= not(layer5_outputs(2060));
    layer6_outputs(3290) <= not((layer5_outputs(927)) or (layer5_outputs(4886)));
    layer6_outputs(3291) <= not(layer5_outputs(1606)) or (layer5_outputs(320));
    layer6_outputs(3292) <= layer5_outputs(289);
    layer6_outputs(3293) <= not(layer5_outputs(2263));
    layer6_outputs(3294) <= not(layer5_outputs(4329));
    layer6_outputs(3295) <= not(layer5_outputs(3368));
    layer6_outputs(3296) <= layer5_outputs(629);
    layer6_outputs(3297) <= (layer5_outputs(87)) and not (layer5_outputs(692));
    layer6_outputs(3298) <= not(layer5_outputs(57));
    layer6_outputs(3299) <= (layer5_outputs(4191)) and (layer5_outputs(5003));
    layer6_outputs(3300) <= not(layer5_outputs(94));
    layer6_outputs(3301) <= (layer5_outputs(2002)) xor (layer5_outputs(585));
    layer6_outputs(3302) <= layer5_outputs(867);
    layer6_outputs(3303) <= not(layer5_outputs(2154));
    layer6_outputs(3304) <= layer5_outputs(4798);
    layer6_outputs(3305) <= (layer5_outputs(1688)) and not (layer5_outputs(3034));
    layer6_outputs(3306) <= (layer5_outputs(3749)) and (layer5_outputs(3016));
    layer6_outputs(3307) <= not(layer5_outputs(4615));
    layer6_outputs(3308) <= layer5_outputs(956);
    layer6_outputs(3309) <= not(layer5_outputs(4335));
    layer6_outputs(3310) <= layer5_outputs(552);
    layer6_outputs(3311) <= not(layer5_outputs(4596));
    layer6_outputs(3312) <= layer5_outputs(5099);
    layer6_outputs(3313) <= layer5_outputs(2718);
    layer6_outputs(3314) <= not(layer5_outputs(4935));
    layer6_outputs(3315) <= not(layer5_outputs(2440));
    layer6_outputs(3316) <= (layer5_outputs(1422)) xor (layer5_outputs(3558));
    layer6_outputs(3317) <= not(layer5_outputs(479));
    layer6_outputs(3318) <= '1';
    layer6_outputs(3319) <= not((layer5_outputs(2988)) xor (layer5_outputs(2391)));
    layer6_outputs(3320) <= not(layer5_outputs(2177));
    layer6_outputs(3321) <= not((layer5_outputs(4995)) xor (layer5_outputs(3855)));
    layer6_outputs(3322) <= (layer5_outputs(4230)) xor (layer5_outputs(2140));
    layer6_outputs(3323) <= not((layer5_outputs(2432)) or (layer5_outputs(3227)));
    layer6_outputs(3324) <= (layer5_outputs(641)) and not (layer5_outputs(1899));
    layer6_outputs(3325) <= layer5_outputs(1870);
    layer6_outputs(3326) <= not(layer5_outputs(3843)) or (layer5_outputs(3781));
    layer6_outputs(3327) <= not(layer5_outputs(205));
    layer6_outputs(3328) <= not(layer5_outputs(2831));
    layer6_outputs(3329) <= not(layer5_outputs(2662));
    layer6_outputs(3330) <= not(layer5_outputs(884));
    layer6_outputs(3331) <= layer5_outputs(2180);
    layer6_outputs(3332) <= layer5_outputs(3543);
    layer6_outputs(3333) <= not(layer5_outputs(1897));
    layer6_outputs(3334) <= layer5_outputs(4875);
    layer6_outputs(3335) <= not(layer5_outputs(873)) or (layer5_outputs(1676));
    layer6_outputs(3336) <= layer5_outputs(12);
    layer6_outputs(3337) <= layer5_outputs(3031);
    layer6_outputs(3338) <= layer5_outputs(1725);
    layer6_outputs(3339) <= not(layer5_outputs(1990));
    layer6_outputs(3340) <= not((layer5_outputs(1030)) xor (layer5_outputs(2589)));
    layer6_outputs(3341) <= layer5_outputs(384);
    layer6_outputs(3342) <= not(layer5_outputs(3950));
    layer6_outputs(3343) <= layer5_outputs(3473);
    layer6_outputs(3344) <= not((layer5_outputs(4693)) xor (layer5_outputs(682)));
    layer6_outputs(3345) <= not(layer5_outputs(3130));
    layer6_outputs(3346) <= not((layer5_outputs(4143)) or (layer5_outputs(2208)));
    layer6_outputs(3347) <= (layer5_outputs(1928)) or (layer5_outputs(1997));
    layer6_outputs(3348) <= (layer5_outputs(1451)) or (layer5_outputs(1026));
    layer6_outputs(3349) <= not(layer5_outputs(4006));
    layer6_outputs(3350) <= (layer5_outputs(2948)) or (layer5_outputs(4460));
    layer6_outputs(3351) <= not(layer5_outputs(1232));
    layer6_outputs(3352) <= layer5_outputs(2130);
    layer6_outputs(3353) <= not(layer5_outputs(2046));
    layer6_outputs(3354) <= not((layer5_outputs(2148)) xor (layer5_outputs(2198)));
    layer6_outputs(3355) <= not(layer5_outputs(3226)) or (layer5_outputs(4620));
    layer6_outputs(3356) <= layer5_outputs(4953);
    layer6_outputs(3357) <= '1';
    layer6_outputs(3358) <= layer5_outputs(3216);
    layer6_outputs(3359) <= (layer5_outputs(4186)) xor (layer5_outputs(3039));
    layer6_outputs(3360) <= layer5_outputs(1072);
    layer6_outputs(3361) <= layer5_outputs(612);
    layer6_outputs(3362) <= not(layer5_outputs(985));
    layer6_outputs(3363) <= not(layer5_outputs(4036)) or (layer5_outputs(2551));
    layer6_outputs(3364) <= not(layer5_outputs(230));
    layer6_outputs(3365) <= layer5_outputs(3309);
    layer6_outputs(3366) <= not(layer5_outputs(1144));
    layer6_outputs(3367) <= not(layer5_outputs(3608));
    layer6_outputs(3368) <= not(layer5_outputs(3098));
    layer6_outputs(3369) <= layer5_outputs(4485);
    layer6_outputs(3370) <= (layer5_outputs(2440)) and not (layer5_outputs(1975));
    layer6_outputs(3371) <= layer5_outputs(1713);
    layer6_outputs(3372) <= (layer5_outputs(3302)) and not (layer5_outputs(3017));
    layer6_outputs(3373) <= not(layer5_outputs(4022)) or (layer5_outputs(5046));
    layer6_outputs(3374) <= layer5_outputs(1839);
    layer6_outputs(3375) <= layer5_outputs(2973);
    layer6_outputs(3376) <= layer5_outputs(4047);
    layer6_outputs(3377) <= layer5_outputs(1917);
    layer6_outputs(3378) <= not(layer5_outputs(1231));
    layer6_outputs(3379) <= not((layer5_outputs(1360)) and (layer5_outputs(76)));
    layer6_outputs(3380) <= (layer5_outputs(2206)) xor (layer5_outputs(999));
    layer6_outputs(3381) <= not((layer5_outputs(1848)) xor (layer5_outputs(2887)));
    layer6_outputs(3382) <= not(layer5_outputs(276));
    layer6_outputs(3383) <= layer5_outputs(4507);
    layer6_outputs(3384) <= layer5_outputs(4841);
    layer6_outputs(3385) <= layer5_outputs(1671);
    layer6_outputs(3386) <= not(layer5_outputs(4219));
    layer6_outputs(3387) <= (layer5_outputs(3405)) and not (layer5_outputs(2266));
    layer6_outputs(3388) <= layer5_outputs(2771);
    layer6_outputs(3389) <= layer5_outputs(461);
    layer6_outputs(3390) <= not(layer5_outputs(3864));
    layer6_outputs(3391) <= (layer5_outputs(4901)) xor (layer5_outputs(1600));
    layer6_outputs(3392) <= (layer5_outputs(2370)) xor (layer5_outputs(1354));
    layer6_outputs(3393) <= not((layer5_outputs(841)) xor (layer5_outputs(2191)));
    layer6_outputs(3394) <= not(layer5_outputs(3880));
    layer6_outputs(3395) <= layer5_outputs(112);
    layer6_outputs(3396) <= not(layer5_outputs(3788));
    layer6_outputs(3397) <= (layer5_outputs(223)) or (layer5_outputs(1331));
    layer6_outputs(3398) <= (layer5_outputs(347)) and (layer5_outputs(775));
    layer6_outputs(3399) <= (layer5_outputs(756)) and (layer5_outputs(974));
    layer6_outputs(3400) <= not(layer5_outputs(1365));
    layer6_outputs(3401) <= not(layer5_outputs(1470));
    layer6_outputs(3402) <= not(layer5_outputs(4117));
    layer6_outputs(3403) <= not(layer5_outputs(2158));
    layer6_outputs(3404) <= (layer5_outputs(4846)) and (layer5_outputs(1338));
    layer6_outputs(3405) <= layer5_outputs(3997);
    layer6_outputs(3406) <= layer5_outputs(3101);
    layer6_outputs(3407) <= not(layer5_outputs(1269));
    layer6_outputs(3408) <= not(layer5_outputs(4054));
    layer6_outputs(3409) <= not(layer5_outputs(1305)) or (layer5_outputs(375));
    layer6_outputs(3410) <= (layer5_outputs(1342)) and not (layer5_outputs(3176));
    layer6_outputs(3411) <= not(layer5_outputs(2373));
    layer6_outputs(3412) <= not(layer5_outputs(3060));
    layer6_outputs(3413) <= not(layer5_outputs(30)) or (layer5_outputs(1714));
    layer6_outputs(3414) <= not((layer5_outputs(1239)) or (layer5_outputs(4534)));
    layer6_outputs(3415) <= not((layer5_outputs(1563)) xor (layer5_outputs(4231)));
    layer6_outputs(3416) <= not(layer5_outputs(4005)) or (layer5_outputs(3941));
    layer6_outputs(3417) <= layer5_outputs(2207);
    layer6_outputs(3418) <= not(layer5_outputs(4893)) or (layer5_outputs(4990));
    layer6_outputs(3419) <= not(layer5_outputs(107));
    layer6_outputs(3420) <= layer5_outputs(111);
    layer6_outputs(3421) <= not(layer5_outputs(3115)) or (layer5_outputs(2420));
    layer6_outputs(3422) <= not(layer5_outputs(1435));
    layer6_outputs(3423) <= (layer5_outputs(1002)) and not (layer5_outputs(3501));
    layer6_outputs(3424) <= not(layer5_outputs(4253)) or (layer5_outputs(3255));
    layer6_outputs(3425) <= not(layer5_outputs(4699));
    layer6_outputs(3426) <= '1';
    layer6_outputs(3427) <= layer5_outputs(316);
    layer6_outputs(3428) <= (layer5_outputs(3714)) and not (layer5_outputs(3724));
    layer6_outputs(3429) <= layer5_outputs(197);
    layer6_outputs(3430) <= (layer5_outputs(2903)) or (layer5_outputs(2775));
    layer6_outputs(3431) <= (layer5_outputs(3200)) or (layer5_outputs(3042));
    layer6_outputs(3432) <= not((layer5_outputs(3316)) or (layer5_outputs(1336)));
    layer6_outputs(3433) <= not(layer5_outputs(4551));
    layer6_outputs(3434) <= not(layer5_outputs(294));
    layer6_outputs(3435) <= not(layer5_outputs(2824));
    layer6_outputs(3436) <= not(layer5_outputs(2242));
    layer6_outputs(3437) <= not(layer5_outputs(3235)) or (layer5_outputs(147));
    layer6_outputs(3438) <= not(layer5_outputs(1932));
    layer6_outputs(3439) <= (layer5_outputs(22)) and not (layer5_outputs(1397));
    layer6_outputs(3440) <= not((layer5_outputs(4295)) and (layer5_outputs(3590)));
    layer6_outputs(3441) <= not(layer5_outputs(1406));
    layer6_outputs(3442) <= (layer5_outputs(3855)) and not (layer5_outputs(2901));
    layer6_outputs(3443) <= layer5_outputs(3956);
    layer6_outputs(3444) <= layer5_outputs(1317);
    layer6_outputs(3445) <= layer5_outputs(2920);
    layer6_outputs(3446) <= not(layer5_outputs(964));
    layer6_outputs(3447) <= not(layer5_outputs(4651));
    layer6_outputs(3448) <= not((layer5_outputs(331)) and (layer5_outputs(1445)));
    layer6_outputs(3449) <= not(layer5_outputs(1681));
    layer6_outputs(3450) <= not(layer5_outputs(4385));
    layer6_outputs(3451) <= not(layer5_outputs(2932));
    layer6_outputs(3452) <= not((layer5_outputs(1986)) and (layer5_outputs(4349)));
    layer6_outputs(3453) <= layer5_outputs(4926);
    layer6_outputs(3454) <= not((layer5_outputs(4843)) xor (layer5_outputs(1136)));
    layer6_outputs(3455) <= (layer5_outputs(3740)) and not (layer5_outputs(528));
    layer6_outputs(3456) <= layer5_outputs(668);
    layer6_outputs(3457) <= not(layer5_outputs(1564));
    layer6_outputs(3458) <= (layer5_outputs(3612)) or (layer5_outputs(460));
    layer6_outputs(3459) <= (layer5_outputs(366)) or (layer5_outputs(4611));
    layer6_outputs(3460) <= not(layer5_outputs(3185));
    layer6_outputs(3461) <= not((layer5_outputs(1980)) xor (layer5_outputs(4864)));
    layer6_outputs(3462) <= (layer5_outputs(1840)) xor (layer5_outputs(1096));
    layer6_outputs(3463) <= (layer5_outputs(3924)) xor (layer5_outputs(326));
    layer6_outputs(3464) <= layer5_outputs(2861);
    layer6_outputs(3465) <= (layer5_outputs(3612)) and not (layer5_outputs(2842));
    layer6_outputs(3466) <= (layer5_outputs(1538)) or (layer5_outputs(1540));
    layer6_outputs(3467) <= not(layer5_outputs(1579));
    layer6_outputs(3468) <= (layer5_outputs(3678)) and not (layer5_outputs(1437));
    layer6_outputs(3469) <= not(layer5_outputs(919));
    layer6_outputs(3470) <= layer5_outputs(2865);
    layer6_outputs(3471) <= not(layer5_outputs(3376));
    layer6_outputs(3472) <= not(layer5_outputs(4497)) or (layer5_outputs(4314));
    layer6_outputs(3473) <= layer5_outputs(2844);
    layer6_outputs(3474) <= not(layer5_outputs(1894));
    layer6_outputs(3475) <= layer5_outputs(2120);
    layer6_outputs(3476) <= not(layer5_outputs(301)) or (layer5_outputs(762));
    layer6_outputs(3477) <= not(layer5_outputs(3649)) or (layer5_outputs(2757));
    layer6_outputs(3478) <= layer5_outputs(2291);
    layer6_outputs(3479) <= not(layer5_outputs(4913));
    layer6_outputs(3480) <= (layer5_outputs(209)) and (layer5_outputs(2482));
    layer6_outputs(3481) <= layer5_outputs(1596);
    layer6_outputs(3482) <= not((layer5_outputs(2259)) or (layer5_outputs(1339)));
    layer6_outputs(3483) <= '1';
    layer6_outputs(3484) <= not((layer5_outputs(3893)) and (layer5_outputs(3335)));
    layer6_outputs(3485) <= layer5_outputs(2523);
    layer6_outputs(3486) <= not(layer5_outputs(704)) or (layer5_outputs(2322));
    layer6_outputs(3487) <= layer5_outputs(2728);
    layer6_outputs(3488) <= (layer5_outputs(1233)) xor (layer5_outputs(3592));
    layer6_outputs(3489) <= layer5_outputs(3360);
    layer6_outputs(3490) <= layer5_outputs(4065);
    layer6_outputs(3491) <= (layer5_outputs(3172)) xor (layer5_outputs(4077));
    layer6_outputs(3492) <= not(layer5_outputs(4737));
    layer6_outputs(3493) <= not(layer5_outputs(827)) or (layer5_outputs(953));
    layer6_outputs(3494) <= (layer5_outputs(3557)) xor (layer5_outputs(2952));
    layer6_outputs(3495) <= not(layer5_outputs(2919));
    layer6_outputs(3496) <= (layer5_outputs(1976)) xor (layer5_outputs(3025));
    layer6_outputs(3497) <= not(layer5_outputs(1866));
    layer6_outputs(3498) <= layer5_outputs(1270);
    layer6_outputs(3499) <= layer5_outputs(2899);
    layer6_outputs(3500) <= layer5_outputs(1088);
    layer6_outputs(3501) <= not(layer5_outputs(4885));
    layer6_outputs(3502) <= (layer5_outputs(2285)) and not (layer5_outputs(1565));
    layer6_outputs(3503) <= layer5_outputs(3888);
    layer6_outputs(3504) <= layer5_outputs(4049);
    layer6_outputs(3505) <= not(layer5_outputs(4153));
    layer6_outputs(3506) <= layer5_outputs(3667);
    layer6_outputs(3507) <= layer5_outputs(3243);
    layer6_outputs(3508) <= not((layer5_outputs(3502)) xor (layer5_outputs(4247)));
    layer6_outputs(3509) <= layer5_outputs(1513);
    layer6_outputs(3510) <= not(layer5_outputs(4696));
    layer6_outputs(3511) <= layer5_outputs(1652);
    layer6_outputs(3512) <= (layer5_outputs(139)) xor (layer5_outputs(2469));
    layer6_outputs(3513) <= not(layer5_outputs(5098));
    layer6_outputs(3514) <= not(layer5_outputs(2373));
    layer6_outputs(3515) <= layer5_outputs(2125);
    layer6_outputs(3516) <= not(layer5_outputs(3877));
    layer6_outputs(3517) <= not((layer5_outputs(3096)) xor (layer5_outputs(3621)));
    layer6_outputs(3518) <= not(layer5_outputs(4456)) or (layer5_outputs(104));
    layer6_outputs(3519) <= not(layer5_outputs(3775));
    layer6_outputs(3520) <= layer5_outputs(954);
    layer6_outputs(3521) <= layer5_outputs(434);
    layer6_outputs(3522) <= layer5_outputs(1386);
    layer6_outputs(3523) <= not((layer5_outputs(2306)) xor (layer5_outputs(316)));
    layer6_outputs(3524) <= layer5_outputs(720);
    layer6_outputs(3525) <= layer5_outputs(2580);
    layer6_outputs(3526) <= not(layer5_outputs(2884));
    layer6_outputs(3527) <= not(layer5_outputs(3347)) or (layer5_outputs(4195));
    layer6_outputs(3528) <= layer5_outputs(3945);
    layer6_outputs(3529) <= layer5_outputs(4359);
    layer6_outputs(3530) <= layer5_outputs(4020);
    layer6_outputs(3531) <= (layer5_outputs(398)) and (layer5_outputs(1002));
    layer6_outputs(3532) <= (layer5_outputs(751)) and (layer5_outputs(806));
    layer6_outputs(3533) <= layer5_outputs(2641);
    layer6_outputs(3534) <= not(layer5_outputs(3876));
    layer6_outputs(3535) <= (layer5_outputs(2006)) and not (layer5_outputs(2021));
    layer6_outputs(3536) <= not((layer5_outputs(678)) xor (layer5_outputs(1959)));
    layer6_outputs(3537) <= (layer5_outputs(3751)) and not (layer5_outputs(1379));
    layer6_outputs(3538) <= layer5_outputs(2804);
    layer6_outputs(3539) <= layer5_outputs(4686);
    layer6_outputs(3540) <= layer5_outputs(2953);
    layer6_outputs(3541) <= layer5_outputs(2547);
    layer6_outputs(3542) <= (layer5_outputs(5068)) xor (layer5_outputs(4376));
    layer6_outputs(3543) <= not(layer5_outputs(3110));
    layer6_outputs(3544) <= layer5_outputs(550);
    layer6_outputs(3545) <= layer5_outputs(4378);
    layer6_outputs(3546) <= not(layer5_outputs(4358));
    layer6_outputs(3547) <= not((layer5_outputs(2712)) or (layer5_outputs(4739)));
    layer6_outputs(3548) <= not((layer5_outputs(2496)) and (layer5_outputs(4654)));
    layer6_outputs(3549) <= not(layer5_outputs(4211));
    layer6_outputs(3550) <= layer5_outputs(5093);
    layer6_outputs(3551) <= layer5_outputs(4431);
    layer6_outputs(3552) <= not((layer5_outputs(1274)) xor (layer5_outputs(2451)));
    layer6_outputs(3553) <= (layer5_outputs(4510)) and not (layer5_outputs(74));
    layer6_outputs(3554) <= not(layer5_outputs(3656));
    layer6_outputs(3555) <= (layer5_outputs(4912)) or (layer5_outputs(3558));
    layer6_outputs(3556) <= layer5_outputs(3066);
    layer6_outputs(3557) <= not((layer5_outputs(3815)) or (layer5_outputs(2125)));
    layer6_outputs(3558) <= layer5_outputs(917);
    layer6_outputs(3559) <= layer5_outputs(2020);
    layer6_outputs(3560) <= not(layer5_outputs(3937));
    layer6_outputs(3561) <= not(layer5_outputs(4527));
    layer6_outputs(3562) <= '1';
    layer6_outputs(3563) <= not((layer5_outputs(488)) xor (layer5_outputs(2383)));
    layer6_outputs(3564) <= not((layer5_outputs(2078)) and (layer5_outputs(3231)));
    layer6_outputs(3565) <= not(layer5_outputs(1891)) or (layer5_outputs(718));
    layer6_outputs(3566) <= layer5_outputs(1237);
    layer6_outputs(3567) <= (layer5_outputs(3610)) or (layer5_outputs(117));
    layer6_outputs(3568) <= not(layer5_outputs(1192));
    layer6_outputs(3569) <= not(layer5_outputs(1639)) or (layer5_outputs(2075));
    layer6_outputs(3570) <= not(layer5_outputs(4727));
    layer6_outputs(3571) <= not(layer5_outputs(4908));
    layer6_outputs(3572) <= not((layer5_outputs(4536)) xor (layer5_outputs(3381)));
    layer6_outputs(3573) <= layer5_outputs(4390);
    layer6_outputs(3574) <= (layer5_outputs(4383)) or (layer5_outputs(2400));
    layer6_outputs(3575) <= not((layer5_outputs(3526)) or (layer5_outputs(3459)));
    layer6_outputs(3576) <= not(layer5_outputs(3693));
    layer6_outputs(3577) <= layer5_outputs(306);
    layer6_outputs(3578) <= not(layer5_outputs(3365));
    layer6_outputs(3579) <= layer5_outputs(228);
    layer6_outputs(3580) <= not(layer5_outputs(894));
    layer6_outputs(3581) <= (layer5_outputs(1217)) xor (layer5_outputs(4358));
    layer6_outputs(3582) <= (layer5_outputs(273)) and not (layer5_outputs(4196));
    layer6_outputs(3583) <= not(layer5_outputs(2633)) or (layer5_outputs(2991));
    layer6_outputs(3584) <= (layer5_outputs(1873)) xor (layer5_outputs(4307));
    layer6_outputs(3585) <= not((layer5_outputs(2439)) or (layer5_outputs(1194)));
    layer6_outputs(3586) <= not((layer5_outputs(4838)) or (layer5_outputs(4102)));
    layer6_outputs(3587) <= layer5_outputs(4553);
    layer6_outputs(3588) <= layer5_outputs(3868);
    layer6_outputs(3589) <= layer5_outputs(3101);
    layer6_outputs(3590) <= not((layer5_outputs(2583)) xor (layer5_outputs(4540)));
    layer6_outputs(3591) <= layer5_outputs(2917);
    layer6_outputs(3592) <= (layer5_outputs(1219)) xor (layer5_outputs(3502));
    layer6_outputs(3593) <= (layer5_outputs(2798)) xor (layer5_outputs(4133));
    layer6_outputs(3594) <= not((layer5_outputs(2137)) xor (layer5_outputs(597)));
    layer6_outputs(3595) <= not((layer5_outputs(1299)) xor (layer5_outputs(1878)));
    layer6_outputs(3596) <= '1';
    layer6_outputs(3597) <= layer5_outputs(2235);
    layer6_outputs(3598) <= layer5_outputs(1590);
    layer6_outputs(3599) <= (layer5_outputs(1359)) or (layer5_outputs(3609));
    layer6_outputs(3600) <= not((layer5_outputs(1174)) and (layer5_outputs(4694)));
    layer6_outputs(3601) <= not(layer5_outputs(504));
    layer6_outputs(3602) <= not((layer5_outputs(1222)) xor (layer5_outputs(2506)));
    layer6_outputs(3603) <= not(layer5_outputs(86));
    layer6_outputs(3604) <= not(layer5_outputs(2627));
    layer6_outputs(3605) <= (layer5_outputs(4880)) and (layer5_outputs(2382));
    layer6_outputs(3606) <= not((layer5_outputs(1171)) xor (layer5_outputs(2504)));
    layer6_outputs(3607) <= not(layer5_outputs(4314)) or (layer5_outputs(4500));
    layer6_outputs(3608) <= not(layer5_outputs(777));
    layer6_outputs(3609) <= (layer5_outputs(3010)) and (layer5_outputs(159));
    layer6_outputs(3610) <= (layer5_outputs(298)) and not (layer5_outputs(1580));
    layer6_outputs(3611) <= not((layer5_outputs(4925)) xor (layer5_outputs(3062)));
    layer6_outputs(3612) <= layer5_outputs(1718);
    layer6_outputs(3613) <= not((layer5_outputs(2743)) xor (layer5_outputs(2548)));
    layer6_outputs(3614) <= layer5_outputs(3064);
    layer6_outputs(3615) <= '1';
    layer6_outputs(3616) <= layer5_outputs(4449);
    layer6_outputs(3617) <= not(layer5_outputs(916));
    layer6_outputs(3618) <= (layer5_outputs(3881)) and (layer5_outputs(3294));
    layer6_outputs(3619) <= layer5_outputs(2022);
    layer6_outputs(3620) <= (layer5_outputs(3197)) and (layer5_outputs(113));
    layer6_outputs(3621) <= not((layer5_outputs(3032)) xor (layer5_outputs(1284)));
    layer6_outputs(3622) <= not(layer5_outputs(3797));
    layer6_outputs(3623) <= layer5_outputs(1924);
    layer6_outputs(3624) <= not(layer5_outputs(3915)) or (layer5_outputs(2044));
    layer6_outputs(3625) <= (layer5_outputs(1618)) xor (layer5_outputs(1595));
    layer6_outputs(3626) <= layer5_outputs(3443);
    layer6_outputs(3627) <= not(layer5_outputs(977)) or (layer5_outputs(969));
    layer6_outputs(3628) <= layer5_outputs(931);
    layer6_outputs(3629) <= layer5_outputs(79);
    layer6_outputs(3630) <= (layer5_outputs(3279)) or (layer5_outputs(1891));
    layer6_outputs(3631) <= (layer5_outputs(883)) or (layer5_outputs(5019));
    layer6_outputs(3632) <= (layer5_outputs(2234)) xor (layer5_outputs(4693));
    layer6_outputs(3633) <= not(layer5_outputs(3361)) or (layer5_outputs(4732));
    layer6_outputs(3634) <= (layer5_outputs(3793)) or (layer5_outputs(3427));
    layer6_outputs(3635) <= layer5_outputs(408);
    layer6_outputs(3636) <= not(layer5_outputs(4081));
    layer6_outputs(3637) <= layer5_outputs(1251);
    layer6_outputs(3638) <= (layer5_outputs(2437)) and (layer5_outputs(3537));
    layer6_outputs(3639) <= not(layer5_outputs(1663));
    layer6_outputs(3640) <= not(layer5_outputs(2191));
    layer6_outputs(3641) <= (layer5_outputs(3938)) or (layer5_outputs(417));
    layer6_outputs(3642) <= (layer5_outputs(3041)) and not (layer5_outputs(748));
    layer6_outputs(3643) <= (layer5_outputs(2752)) and (layer5_outputs(1433));
    layer6_outputs(3644) <= not(layer5_outputs(1774));
    layer6_outputs(3645) <= not((layer5_outputs(3593)) xor (layer5_outputs(2193)));
    layer6_outputs(3646) <= not(layer5_outputs(1674));
    layer6_outputs(3647) <= not(layer5_outputs(2888));
    layer6_outputs(3648) <= not(layer5_outputs(3216));
    layer6_outputs(3649) <= (layer5_outputs(2014)) xor (layer5_outputs(4896));
    layer6_outputs(3650) <= layer5_outputs(2155);
    layer6_outputs(3651) <= not((layer5_outputs(5087)) xor (layer5_outputs(3485)));
    layer6_outputs(3652) <= layer5_outputs(399);
    layer6_outputs(3653) <= layer5_outputs(1198);
    layer6_outputs(3654) <= layer5_outputs(3664);
    layer6_outputs(3655) <= (layer5_outputs(5065)) and (layer5_outputs(3503));
    layer6_outputs(3656) <= not(layer5_outputs(152));
    layer6_outputs(3657) <= not(layer5_outputs(4746)) or (layer5_outputs(2838));
    layer6_outputs(3658) <= not(layer5_outputs(83));
    layer6_outputs(3659) <= not((layer5_outputs(474)) and (layer5_outputs(792)));
    layer6_outputs(3660) <= not(layer5_outputs(1738));
    layer6_outputs(3661) <= not((layer5_outputs(1187)) or (layer5_outputs(3705)));
    layer6_outputs(3662) <= not(layer5_outputs(989));
    layer6_outputs(3663) <= layer5_outputs(3080);
    layer6_outputs(3664) <= not((layer5_outputs(1756)) or (layer5_outputs(3392)));
    layer6_outputs(3665) <= (layer5_outputs(275)) and not (layer5_outputs(436));
    layer6_outputs(3666) <= (layer5_outputs(3262)) xor (layer5_outputs(971));
    layer6_outputs(3667) <= (layer5_outputs(834)) and not (layer5_outputs(4982));
    layer6_outputs(3668) <= not((layer5_outputs(4437)) xor (layer5_outputs(3596)));
    layer6_outputs(3669) <= (layer5_outputs(2826)) and (layer5_outputs(4264));
    layer6_outputs(3670) <= not(layer5_outputs(1958));
    layer6_outputs(3671) <= (layer5_outputs(4512)) and not (layer5_outputs(2861));
    layer6_outputs(3672) <= (layer5_outputs(37)) or (layer5_outputs(4623));
    layer6_outputs(3673) <= layer5_outputs(2302);
    layer6_outputs(3674) <= (layer5_outputs(800)) and not (layer5_outputs(4593));
    layer6_outputs(3675) <= (layer5_outputs(3038)) or (layer5_outputs(272));
    layer6_outputs(3676) <= layer5_outputs(1079);
    layer6_outputs(3677) <= not(layer5_outputs(2209));
    layer6_outputs(3678) <= not(layer5_outputs(3491));
    layer6_outputs(3679) <= (layer5_outputs(3192)) xor (layer5_outputs(3792));
    layer6_outputs(3680) <= not(layer5_outputs(1473)) or (layer5_outputs(1313));
    layer6_outputs(3681) <= not(layer5_outputs(908)) or (layer5_outputs(886));
    layer6_outputs(3682) <= (layer5_outputs(2035)) xor (layer5_outputs(733));
    layer6_outputs(3683) <= not(layer5_outputs(1288));
    layer6_outputs(3684) <= (layer5_outputs(1450)) and not (layer5_outputs(573));
    layer6_outputs(3685) <= '0';
    layer6_outputs(3686) <= layer5_outputs(832);
    layer6_outputs(3687) <= not((layer5_outputs(4553)) and (layer5_outputs(4656)));
    layer6_outputs(3688) <= layer5_outputs(3826);
    layer6_outputs(3689) <= not(layer5_outputs(2452)) or (layer5_outputs(421));
    layer6_outputs(3690) <= '1';
    layer6_outputs(3691) <= (layer5_outputs(2665)) and not (layer5_outputs(2620));
    layer6_outputs(3692) <= '1';
    layer6_outputs(3693) <= layer5_outputs(130);
    layer6_outputs(3694) <= not(layer5_outputs(1753));
    layer6_outputs(3695) <= not(layer5_outputs(2307));
    layer6_outputs(3696) <= not((layer5_outputs(4436)) xor (layer5_outputs(1497)));
    layer6_outputs(3697) <= layer5_outputs(932);
    layer6_outputs(3698) <= layer5_outputs(587);
    layer6_outputs(3699) <= '1';
    layer6_outputs(3700) <= not(layer5_outputs(205)) or (layer5_outputs(2521));
    layer6_outputs(3701) <= not(layer5_outputs(1673));
    layer6_outputs(3702) <= not((layer5_outputs(807)) xor (layer5_outputs(93)));
    layer6_outputs(3703) <= not(layer5_outputs(3730));
    layer6_outputs(3704) <= layer5_outputs(2890);
    layer6_outputs(3705) <= (layer5_outputs(3594)) and (layer5_outputs(1089));
    layer6_outputs(3706) <= not(layer5_outputs(4400));
    layer6_outputs(3707) <= not((layer5_outputs(1536)) and (layer5_outputs(2898)));
    layer6_outputs(3708) <= not(layer5_outputs(2897)) or (layer5_outputs(3418));
    layer6_outputs(3709) <= layer5_outputs(2583);
    layer6_outputs(3710) <= not((layer5_outputs(4142)) xor (layer5_outputs(1739)));
    layer6_outputs(3711) <= not(layer5_outputs(1898));
    layer6_outputs(3712) <= not(layer5_outputs(318));
    layer6_outputs(3713) <= '1';
    layer6_outputs(3714) <= not(layer5_outputs(959));
    layer6_outputs(3715) <= not(layer5_outputs(4391));
    layer6_outputs(3716) <= not(layer5_outputs(1652));
    layer6_outputs(3717) <= (layer5_outputs(1529)) xor (layer5_outputs(1148));
    layer6_outputs(3718) <= not((layer5_outputs(221)) or (layer5_outputs(4921)));
    layer6_outputs(3719) <= not(layer5_outputs(2424));
    layer6_outputs(3720) <= (layer5_outputs(2444)) and not (layer5_outputs(2025));
    layer6_outputs(3721) <= layer5_outputs(3766);
    layer6_outputs(3722) <= (layer5_outputs(2080)) or (layer5_outputs(833));
    layer6_outputs(3723) <= not(layer5_outputs(1030));
    layer6_outputs(3724) <= not((layer5_outputs(3908)) xor (layer5_outputs(771)));
    layer6_outputs(3725) <= not(layer5_outputs(3574));
    layer6_outputs(3726) <= layer5_outputs(2497);
    layer6_outputs(3727) <= not(layer5_outputs(4733));
    layer6_outputs(3728) <= (layer5_outputs(3599)) or (layer5_outputs(698));
    layer6_outputs(3729) <= not(layer5_outputs(3012));
    layer6_outputs(3730) <= layer5_outputs(3418);
    layer6_outputs(3731) <= not(layer5_outputs(4400));
    layer6_outputs(3732) <= layer5_outputs(4729);
    layer6_outputs(3733) <= layer5_outputs(4017);
    layer6_outputs(3734) <= layer5_outputs(1112);
    layer6_outputs(3735) <= not(layer5_outputs(4507));
    layer6_outputs(3736) <= layer5_outputs(389);
    layer6_outputs(3737) <= not(layer5_outputs(449));
    layer6_outputs(3738) <= (layer5_outputs(4482)) and (layer5_outputs(4192));
    layer6_outputs(3739) <= not(layer5_outputs(1476));
    layer6_outputs(3740) <= (layer5_outputs(4291)) xor (layer5_outputs(4334));
    layer6_outputs(3741) <= not(layer5_outputs(4920)) or (layer5_outputs(3237));
    layer6_outputs(3742) <= layer5_outputs(3442);
    layer6_outputs(3743) <= not(layer5_outputs(1519));
    layer6_outputs(3744) <= not(layer5_outputs(3091));
    layer6_outputs(3745) <= layer5_outputs(2833);
    layer6_outputs(3746) <= not(layer5_outputs(2817));
    layer6_outputs(3747) <= layer5_outputs(1248);
    layer6_outputs(3748) <= not(layer5_outputs(3044)) or (layer5_outputs(4075));
    layer6_outputs(3749) <= (layer5_outputs(2721)) or (layer5_outputs(2455));
    layer6_outputs(3750) <= (layer5_outputs(1606)) xor (layer5_outputs(2048));
    layer6_outputs(3751) <= not(layer5_outputs(2244));
    layer6_outputs(3752) <= not(layer5_outputs(3666));
    layer6_outputs(3753) <= (layer5_outputs(3409)) and (layer5_outputs(2566));
    layer6_outputs(3754) <= layer5_outputs(4459);
    layer6_outputs(3755) <= (layer5_outputs(4535)) and (layer5_outputs(41));
    layer6_outputs(3756) <= layer5_outputs(994);
    layer6_outputs(3757) <= (layer5_outputs(4892)) xor (layer5_outputs(4502));
    layer6_outputs(3758) <= not(layer5_outputs(3871));
    layer6_outputs(3759) <= (layer5_outputs(1303)) xor (layer5_outputs(741));
    layer6_outputs(3760) <= not(layer5_outputs(215));
    layer6_outputs(3761) <= layer5_outputs(647);
    layer6_outputs(3762) <= (layer5_outputs(2512)) and (layer5_outputs(4248));
    layer6_outputs(3763) <= layer5_outputs(208);
    layer6_outputs(3764) <= layer5_outputs(68);
    layer6_outputs(3765) <= layer5_outputs(2493);
    layer6_outputs(3766) <= (layer5_outputs(1498)) xor (layer5_outputs(3084));
    layer6_outputs(3767) <= layer5_outputs(2450);
    layer6_outputs(3768) <= not((layer5_outputs(2032)) or (layer5_outputs(4523)));
    layer6_outputs(3769) <= not((layer5_outputs(3790)) xor (layer5_outputs(3565)));
    layer6_outputs(3770) <= (layer5_outputs(3674)) and not (layer5_outputs(2015));
    layer6_outputs(3771) <= not((layer5_outputs(749)) and (layer5_outputs(1093)));
    layer6_outputs(3772) <= not(layer5_outputs(2001));
    layer6_outputs(3773) <= (layer5_outputs(1440)) and not (layer5_outputs(1757));
    layer6_outputs(3774) <= (layer5_outputs(1947)) xor (layer5_outputs(3293));
    layer6_outputs(3775) <= not(layer5_outputs(4082)) or (layer5_outputs(2887));
    layer6_outputs(3776) <= layer5_outputs(349);
    layer6_outputs(3777) <= layer5_outputs(74);
    layer6_outputs(3778) <= layer5_outputs(1788);
    layer6_outputs(3779) <= layer5_outputs(371);
    layer6_outputs(3780) <= not((layer5_outputs(98)) xor (layer5_outputs(4622)));
    layer6_outputs(3781) <= not(layer5_outputs(3773));
    layer6_outputs(3782) <= not(layer5_outputs(937)) or (layer5_outputs(4170));
    layer6_outputs(3783) <= not(layer5_outputs(4508));
    layer6_outputs(3784) <= (layer5_outputs(4244)) and not (layer5_outputs(2147));
    layer6_outputs(3785) <= (layer5_outputs(2444)) xor (layer5_outputs(903));
    layer6_outputs(3786) <= not(layer5_outputs(2533));
    layer6_outputs(3787) <= (layer5_outputs(1440)) and (layer5_outputs(818));
    layer6_outputs(3788) <= (layer5_outputs(193)) xor (layer5_outputs(4903));
    layer6_outputs(3789) <= '1';
    layer6_outputs(3790) <= layer5_outputs(3676);
    layer6_outputs(3791) <= not(layer5_outputs(10)) or (layer5_outputs(3662));
    layer6_outputs(3792) <= not(layer5_outputs(4463));
    layer6_outputs(3793) <= not((layer5_outputs(1009)) or (layer5_outputs(2401)));
    layer6_outputs(3794) <= not(layer5_outputs(1863));
    layer6_outputs(3795) <= layer5_outputs(3132);
    layer6_outputs(3796) <= not(layer5_outputs(1662));
    layer6_outputs(3797) <= (layer5_outputs(218)) and not (layer5_outputs(1099));
    layer6_outputs(3798) <= not(layer5_outputs(2974));
    layer6_outputs(3799) <= not(layer5_outputs(2238));
    layer6_outputs(3800) <= not(layer5_outputs(4917));
    layer6_outputs(3801) <= not(layer5_outputs(3719));
    layer6_outputs(3802) <= not(layer5_outputs(3065));
    layer6_outputs(3803) <= layer5_outputs(263);
    layer6_outputs(3804) <= (layer5_outputs(210)) and (layer5_outputs(3704));
    layer6_outputs(3805) <= (layer5_outputs(3892)) xor (layer5_outputs(4090));
    layer6_outputs(3806) <= (layer5_outputs(4772)) and not (layer5_outputs(369));
    layer6_outputs(3807) <= (layer5_outputs(3916)) and (layer5_outputs(2378));
    layer6_outputs(3808) <= not(layer5_outputs(3500));
    layer6_outputs(3809) <= layer5_outputs(1374);
    layer6_outputs(3810) <= not(layer5_outputs(697));
    layer6_outputs(3811) <= layer5_outputs(3764);
    layer6_outputs(3812) <= layer5_outputs(3432);
    layer6_outputs(3813) <= (layer5_outputs(1746)) xor (layer5_outputs(3646));
    layer6_outputs(3814) <= not(layer5_outputs(3805));
    layer6_outputs(3815) <= not((layer5_outputs(4610)) or (layer5_outputs(3379)));
    layer6_outputs(3816) <= '1';
    layer6_outputs(3817) <= not(layer5_outputs(1626));
    layer6_outputs(3818) <= '1';
    layer6_outputs(3819) <= not(layer5_outputs(563));
    layer6_outputs(3820) <= not(layer5_outputs(2108)) or (layer5_outputs(4614));
    layer6_outputs(3821) <= layer5_outputs(4509);
    layer6_outputs(3822) <= not(layer5_outputs(2577)) or (layer5_outputs(4704));
    layer6_outputs(3823) <= '0';
    layer6_outputs(3824) <= not((layer5_outputs(1688)) or (layer5_outputs(4323)));
    layer6_outputs(3825) <= (layer5_outputs(1631)) or (layer5_outputs(2033));
    layer6_outputs(3826) <= not((layer5_outputs(2469)) xor (layer5_outputs(3435)));
    layer6_outputs(3827) <= not(layer5_outputs(3952)) or (layer5_outputs(1449));
    layer6_outputs(3828) <= layer5_outputs(350);
    layer6_outputs(3829) <= layer5_outputs(1106);
    layer6_outputs(3830) <= not(layer5_outputs(4589));
    layer6_outputs(3831) <= layer5_outputs(4790);
    layer6_outputs(3832) <= layer5_outputs(1123);
    layer6_outputs(3833) <= layer5_outputs(1322);
    layer6_outputs(3834) <= not(layer5_outputs(1205));
    layer6_outputs(3835) <= (layer5_outputs(1033)) and not (layer5_outputs(2202));
    layer6_outputs(3836) <= layer5_outputs(1873);
    layer6_outputs(3837) <= (layer5_outputs(1379)) and (layer5_outputs(3532));
    layer6_outputs(3838) <= (layer5_outputs(212)) or (layer5_outputs(3325));
    layer6_outputs(3839) <= not((layer5_outputs(1110)) or (layer5_outputs(712)));
    layer6_outputs(3840) <= not((layer5_outputs(2247)) xor (layer5_outputs(1159)));
    layer6_outputs(3841) <= not(layer5_outputs(3774));
    layer6_outputs(3842) <= not(layer5_outputs(2646));
    layer6_outputs(3843) <= layer5_outputs(4258);
    layer6_outputs(3844) <= not(layer5_outputs(4501));
    layer6_outputs(3845) <= not(layer5_outputs(1287));
    layer6_outputs(3846) <= (layer5_outputs(2773)) or (layer5_outputs(1744));
    layer6_outputs(3847) <= (layer5_outputs(1637)) xor (layer5_outputs(1937));
    layer6_outputs(3848) <= not(layer5_outputs(1134)) or (layer5_outputs(93));
    layer6_outputs(3849) <= not(layer5_outputs(4289)) or (layer5_outputs(4444));
    layer6_outputs(3850) <= layer5_outputs(2316);
    layer6_outputs(3851) <= not((layer5_outputs(1995)) or (layer5_outputs(5109)));
    layer6_outputs(3852) <= not((layer5_outputs(598)) and (layer5_outputs(3394)));
    layer6_outputs(3853) <= layer5_outputs(4003);
    layer6_outputs(3854) <= not(layer5_outputs(993));
    layer6_outputs(3855) <= (layer5_outputs(4852)) or (layer5_outputs(517));
    layer6_outputs(3856) <= not(layer5_outputs(4265));
    layer6_outputs(3857) <= (layer5_outputs(1983)) and (layer5_outputs(3824));
    layer6_outputs(3858) <= not((layer5_outputs(2334)) and (layer5_outputs(1469)));
    layer6_outputs(3859) <= not(layer5_outputs(4572)) or (layer5_outputs(4315));
    layer6_outputs(3860) <= not(layer5_outputs(32)) or (layer5_outputs(2156));
    layer6_outputs(3861) <= layer5_outputs(4506);
    layer6_outputs(3862) <= (layer5_outputs(4035)) and not (layer5_outputs(1720));
    layer6_outputs(3863) <= not(layer5_outputs(1388));
    layer6_outputs(3864) <= not(layer5_outputs(1821));
    layer6_outputs(3865) <= not(layer5_outputs(2531)) or (layer5_outputs(3167));
    layer6_outputs(3866) <= layer5_outputs(4529);
    layer6_outputs(3867) <= not(layer5_outputs(2667)) or (layer5_outputs(2472));
    layer6_outputs(3868) <= (layer5_outputs(553)) and not (layer5_outputs(2014));
    layer6_outputs(3869) <= not(layer5_outputs(4639)) or (layer5_outputs(3181));
    layer6_outputs(3870) <= (layer5_outputs(1747)) or (layer5_outputs(3544));
    layer6_outputs(3871) <= not(layer5_outputs(1686));
    layer6_outputs(3872) <= not((layer5_outputs(2059)) or (layer5_outputs(735)));
    layer6_outputs(3873) <= not(layer5_outputs(3306));
    layer6_outputs(3874) <= layer5_outputs(3305);
    layer6_outputs(3875) <= not(layer5_outputs(131));
    layer6_outputs(3876) <= '0';
    layer6_outputs(3877) <= (layer5_outputs(710)) xor (layer5_outputs(4782));
    layer6_outputs(3878) <= not(layer5_outputs(1625));
    layer6_outputs(3879) <= not(layer5_outputs(3762));
    layer6_outputs(3880) <= (layer5_outputs(3086)) and not (layer5_outputs(611));
    layer6_outputs(3881) <= layer5_outputs(3332);
    layer6_outputs(3882) <= layer5_outputs(4825);
    layer6_outputs(3883) <= not(layer5_outputs(5090));
    layer6_outputs(3884) <= not(layer5_outputs(4384)) or (layer5_outputs(4539));
    layer6_outputs(3885) <= not((layer5_outputs(3574)) or (layer5_outputs(1879)));
    layer6_outputs(3886) <= not((layer5_outputs(3429)) or (layer5_outputs(2995)));
    layer6_outputs(3887) <= not(layer5_outputs(3412));
    layer6_outputs(3888) <= (layer5_outputs(3253)) and not (layer5_outputs(4092));
    layer6_outputs(3889) <= not(layer5_outputs(670));
    layer6_outputs(3890) <= layer5_outputs(3599);
    layer6_outputs(3891) <= not(layer5_outputs(1327));
    layer6_outputs(3892) <= layer5_outputs(3266);
    layer6_outputs(3893) <= layer5_outputs(4763);
    layer6_outputs(3894) <= (layer5_outputs(501)) and (layer5_outputs(1886));
    layer6_outputs(3895) <= layer5_outputs(4114);
    layer6_outputs(3896) <= layer5_outputs(3451);
    layer6_outputs(3897) <= not(layer5_outputs(2410));
    layer6_outputs(3898) <= layer5_outputs(2431);
    layer6_outputs(3899) <= not((layer5_outputs(254)) xor (layer5_outputs(4256)));
    layer6_outputs(3900) <= layer5_outputs(4833);
    layer6_outputs(3901) <= layer5_outputs(3936);
    layer6_outputs(3902) <= layer5_outputs(3114);
    layer6_outputs(3903) <= '1';
    layer6_outputs(3904) <= layer5_outputs(1904);
    layer6_outputs(3905) <= not((layer5_outputs(3834)) or (layer5_outputs(403)));
    layer6_outputs(3906) <= not(layer5_outputs(2064)) or (layer5_outputs(2053));
    layer6_outputs(3907) <= not(layer5_outputs(4236));
    layer6_outputs(3908) <= not((layer5_outputs(3078)) and (layer5_outputs(1338)));
    layer6_outputs(3909) <= layer5_outputs(3706);
    layer6_outputs(3910) <= (layer5_outputs(392)) and (layer5_outputs(661));
    layer6_outputs(3911) <= layer5_outputs(2791);
    layer6_outputs(3912) <= (layer5_outputs(2488)) or (layer5_outputs(1774));
    layer6_outputs(3913) <= not(layer5_outputs(55));
    layer6_outputs(3914) <= (layer5_outputs(578)) and not (layer5_outputs(4441));
    layer6_outputs(3915) <= not((layer5_outputs(4977)) and (layer5_outputs(1611)));
    layer6_outputs(3916) <= layer5_outputs(2904);
    layer6_outputs(3917) <= not((layer5_outputs(360)) xor (layer5_outputs(2851)));
    layer6_outputs(3918) <= not(layer5_outputs(3436)) or (layer5_outputs(4074));
    layer6_outputs(3919) <= (layer5_outputs(1940)) xor (layer5_outputs(98));
    layer6_outputs(3920) <= layer5_outputs(2227);
    layer6_outputs(3921) <= layer5_outputs(453);
    layer6_outputs(3922) <= (layer5_outputs(1650)) and not (layer5_outputs(4612));
    layer6_outputs(3923) <= layer5_outputs(2413);
    layer6_outputs(3924) <= layer5_outputs(2534);
    layer6_outputs(3925) <= not(layer5_outputs(1122));
    layer6_outputs(3926) <= not(layer5_outputs(3582)) or (layer5_outputs(4382));
    layer6_outputs(3927) <= (layer5_outputs(2293)) or (layer5_outputs(1371));
    layer6_outputs(3928) <= not(layer5_outputs(2269));
    layer6_outputs(3929) <= not(layer5_outputs(172));
    layer6_outputs(3930) <= not(layer5_outputs(3987));
    layer6_outputs(3931) <= layer5_outputs(3218);
    layer6_outputs(3932) <= layer5_outputs(1097);
    layer6_outputs(3933) <= not((layer5_outputs(3736)) xor (layer5_outputs(2187)));
    layer6_outputs(3934) <= not((layer5_outputs(1783)) and (layer5_outputs(2989)));
    layer6_outputs(3935) <= (layer5_outputs(583)) and not (layer5_outputs(3168));
    layer6_outputs(3936) <= not(layer5_outputs(3032));
    layer6_outputs(3937) <= (layer5_outputs(4399)) and not (layer5_outputs(300));
    layer6_outputs(3938) <= not(layer5_outputs(4833));
    layer6_outputs(3939) <= not((layer5_outputs(332)) or (layer5_outputs(4429)));
    layer6_outputs(3940) <= not(layer5_outputs(3327)) or (layer5_outputs(3034));
    layer6_outputs(3941) <= not((layer5_outputs(4187)) and (layer5_outputs(100)));
    layer6_outputs(3942) <= not(layer5_outputs(3928));
    layer6_outputs(3943) <= layer5_outputs(189);
    layer6_outputs(3944) <= (layer5_outputs(851)) xor (layer5_outputs(2059));
    layer6_outputs(3945) <= not(layer5_outputs(2855));
    layer6_outputs(3946) <= (layer5_outputs(2279)) and (layer5_outputs(1950));
    layer6_outputs(3947) <= not(layer5_outputs(4542));
    layer6_outputs(3948) <= not((layer5_outputs(4117)) xor (layer5_outputs(256)));
    layer6_outputs(3949) <= (layer5_outputs(2453)) xor (layer5_outputs(3870));
    layer6_outputs(3950) <= layer5_outputs(552);
    layer6_outputs(3951) <= not((layer5_outputs(4903)) and (layer5_outputs(2348)));
    layer6_outputs(3952) <= (layer5_outputs(1507)) and not (layer5_outputs(2731));
    layer6_outputs(3953) <= not((layer5_outputs(2378)) or (layer5_outputs(4764)));
    layer6_outputs(3954) <= not((layer5_outputs(1666)) xor (layer5_outputs(4886)));
    layer6_outputs(3955) <= layer5_outputs(2135);
    layer6_outputs(3956) <= layer5_outputs(4870);
    layer6_outputs(3957) <= (layer5_outputs(311)) and (layer5_outputs(921));
    layer6_outputs(3958) <= not((layer5_outputs(404)) xor (layer5_outputs(5031)));
    layer6_outputs(3959) <= not(layer5_outputs(3410));
    layer6_outputs(3960) <= (layer5_outputs(755)) and not (layer5_outputs(185));
    layer6_outputs(3961) <= layer5_outputs(579);
    layer6_outputs(3962) <= not(layer5_outputs(4280));
    layer6_outputs(3963) <= not((layer5_outputs(1726)) and (layer5_outputs(860)));
    layer6_outputs(3964) <= layer5_outputs(2241);
    layer6_outputs(3965) <= layer5_outputs(1960);
    layer6_outputs(3966) <= not(layer5_outputs(2922));
    layer6_outputs(3967) <= layer5_outputs(2806);
    layer6_outputs(3968) <= layer5_outputs(85);
    layer6_outputs(3969) <= layer5_outputs(3563);
    layer6_outputs(3970) <= (layer5_outputs(523)) and (layer5_outputs(126));
    layer6_outputs(3971) <= (layer5_outputs(3659)) xor (layer5_outputs(3576));
    layer6_outputs(3972) <= layer5_outputs(3122);
    layer6_outputs(3973) <= layer5_outputs(1094);
    layer6_outputs(3974) <= layer5_outputs(2532);
    layer6_outputs(3975) <= '0';
    layer6_outputs(3976) <= layer5_outputs(5012);
    layer6_outputs(3977) <= not((layer5_outputs(4274)) and (layer5_outputs(2937)));
    layer6_outputs(3978) <= (layer5_outputs(2815)) xor (layer5_outputs(3768));
    layer6_outputs(3979) <= (layer5_outputs(5089)) xor (layer5_outputs(1422));
    layer6_outputs(3980) <= not(layer5_outputs(4533)) or (layer5_outputs(973));
    layer6_outputs(3981) <= not(layer5_outputs(394));
    layer6_outputs(3982) <= not(layer5_outputs(2498));
    layer6_outputs(3983) <= (layer5_outputs(570)) and not (layer5_outputs(2620));
    layer6_outputs(3984) <= layer5_outputs(4883);
    layer6_outputs(3985) <= not(layer5_outputs(4239));
    layer6_outputs(3986) <= not((layer5_outputs(2724)) or (layer5_outputs(5119)));
    layer6_outputs(3987) <= layer5_outputs(3260);
    layer6_outputs(3988) <= not(layer5_outputs(3500));
    layer6_outputs(3989) <= not(layer5_outputs(183));
    layer6_outputs(3990) <= not(layer5_outputs(497));
    layer6_outputs(3991) <= layer5_outputs(606);
    layer6_outputs(3992) <= (layer5_outputs(746)) xor (layer5_outputs(621));
    layer6_outputs(3993) <= layer5_outputs(1257);
    layer6_outputs(3994) <= not((layer5_outputs(4909)) and (layer5_outputs(981)));
    layer6_outputs(3995) <= not((layer5_outputs(3129)) xor (layer5_outputs(182)));
    layer6_outputs(3996) <= not(layer5_outputs(3698));
    layer6_outputs(3997) <= layer5_outputs(1213);
    layer6_outputs(3998) <= layer5_outputs(1446);
    layer6_outputs(3999) <= not(layer5_outputs(1195));
    layer6_outputs(4000) <= layer5_outputs(2217);
    layer6_outputs(4001) <= not(layer5_outputs(118));
    layer6_outputs(4002) <= '1';
    layer6_outputs(4003) <= not((layer5_outputs(4205)) or (layer5_outputs(3468)));
    layer6_outputs(4004) <= not((layer5_outputs(2771)) and (layer5_outputs(4154)));
    layer6_outputs(4005) <= not(layer5_outputs(4659));
    layer6_outputs(4006) <= '1';
    layer6_outputs(4007) <= (layer5_outputs(226)) or (layer5_outputs(3238));
    layer6_outputs(4008) <= layer5_outputs(4966);
    layer6_outputs(4009) <= layer5_outputs(2010);
    layer6_outputs(4010) <= (layer5_outputs(1939)) and not (layer5_outputs(1725));
    layer6_outputs(4011) <= (layer5_outputs(596)) and not (layer5_outputs(2058));
    layer6_outputs(4012) <= (layer5_outputs(1165)) and not (layer5_outputs(2399));
    layer6_outputs(4013) <= not(layer5_outputs(4536));
    layer6_outputs(4014) <= (layer5_outputs(2937)) xor (layer5_outputs(1575));
    layer6_outputs(4015) <= layer5_outputs(4716);
    layer6_outputs(4016) <= not(layer5_outputs(5018));
    layer6_outputs(4017) <= not(layer5_outputs(102));
    layer6_outputs(4018) <= not((layer5_outputs(4086)) xor (layer5_outputs(2038)));
    layer6_outputs(4019) <= not((layer5_outputs(424)) xor (layer5_outputs(2893)));
    layer6_outputs(4020) <= not(layer5_outputs(2973));
    layer6_outputs(4021) <= not(layer5_outputs(3557));
    layer6_outputs(4022) <= (layer5_outputs(3561)) and not (layer5_outputs(3441));
    layer6_outputs(4023) <= not(layer5_outputs(3563));
    layer6_outputs(4024) <= (layer5_outputs(1886)) and not (layer5_outputs(3691));
    layer6_outputs(4025) <= not((layer5_outputs(59)) and (layer5_outputs(1655)));
    layer6_outputs(4026) <= not(layer5_outputs(1800));
    layer6_outputs(4027) <= (layer5_outputs(4786)) and (layer5_outputs(165));
    layer6_outputs(4028) <= not(layer5_outputs(5113)) or (layer5_outputs(2741));
    layer6_outputs(4029) <= layer5_outputs(3984);
    layer6_outputs(4030) <= layer5_outputs(383);
    layer6_outputs(4031) <= (layer5_outputs(2627)) and not (layer5_outputs(1254));
    layer6_outputs(4032) <= (layer5_outputs(3645)) xor (layer5_outputs(3264));
    layer6_outputs(4033) <= not(layer5_outputs(3746)) or (layer5_outputs(2745));
    layer6_outputs(4034) <= not((layer5_outputs(243)) xor (layer5_outputs(2685)));
    layer6_outputs(4035) <= layer5_outputs(368);
    layer6_outputs(4036) <= not(layer5_outputs(2612)) or (layer5_outputs(866));
    layer6_outputs(4037) <= layer5_outputs(2098);
    layer6_outputs(4038) <= (layer5_outputs(135)) xor (layer5_outputs(4042));
    layer6_outputs(4039) <= not(layer5_outputs(1271));
    layer6_outputs(4040) <= layer5_outputs(3045);
    layer6_outputs(4041) <= layer5_outputs(4862);
    layer6_outputs(4042) <= (layer5_outputs(1679)) or (layer5_outputs(2971));
    layer6_outputs(4043) <= not(layer5_outputs(2546));
    layer6_outputs(4044) <= not((layer5_outputs(3856)) or (layer5_outputs(4388)));
    layer6_outputs(4045) <= not(layer5_outputs(2834)) or (layer5_outputs(4625));
    layer6_outputs(4046) <= not(layer5_outputs(1940));
    layer6_outputs(4047) <= (layer5_outputs(1084)) and not (layer5_outputs(4013));
    layer6_outputs(4048) <= not(layer5_outputs(248));
    layer6_outputs(4049) <= (layer5_outputs(2733)) or (layer5_outputs(3782));
    layer6_outputs(4050) <= not((layer5_outputs(1653)) or (layer5_outputs(4925)));
    layer6_outputs(4051) <= (layer5_outputs(177)) and not (layer5_outputs(2388));
    layer6_outputs(4052) <= '1';
    layer6_outputs(4053) <= layer5_outputs(1515);
    layer6_outputs(4054) <= not(layer5_outputs(2946));
    layer6_outputs(4055) <= not(layer5_outputs(3003));
    layer6_outputs(4056) <= layer5_outputs(3134);
    layer6_outputs(4057) <= not(layer5_outputs(4064));
    layer6_outputs(4058) <= not(layer5_outputs(3899));
    layer6_outputs(4059) <= (layer5_outputs(351)) and not (layer5_outputs(1787));
    layer6_outputs(4060) <= (layer5_outputs(357)) xor (layer5_outputs(707));
    layer6_outputs(4061) <= not(layer5_outputs(865));
    layer6_outputs(4062) <= not(layer5_outputs(3770));
    layer6_outputs(4063) <= not(layer5_outputs(3758));
    layer6_outputs(4064) <= layer5_outputs(577);
    layer6_outputs(4065) <= (layer5_outputs(498)) xor (layer5_outputs(4321));
    layer6_outputs(4066) <= not((layer5_outputs(3030)) or (layer5_outputs(1272)));
    layer6_outputs(4067) <= (layer5_outputs(303)) and not (layer5_outputs(2655));
    layer6_outputs(4068) <= not((layer5_outputs(3917)) xor (layer5_outputs(4830)));
    layer6_outputs(4069) <= not(layer5_outputs(3568)) or (layer5_outputs(3257));
    layer6_outputs(4070) <= layer5_outputs(1146);
    layer6_outputs(4071) <= not(layer5_outputs(2765));
    layer6_outputs(4072) <= (layer5_outputs(710)) and (layer5_outputs(1477));
    layer6_outputs(4073) <= not(layer5_outputs(2803));
    layer6_outputs(4074) <= layer5_outputs(2886);
    layer6_outputs(4075) <= layer5_outputs(1307);
    layer6_outputs(4076) <= not((layer5_outputs(529)) or (layer5_outputs(4910)));
    layer6_outputs(4077) <= (layer5_outputs(4156)) or (layer5_outputs(2114));
    layer6_outputs(4078) <= not(layer5_outputs(186));
    layer6_outputs(4079) <= not((layer5_outputs(3556)) or (layer5_outputs(2478)));
    layer6_outputs(4080) <= layer5_outputs(4501);
    layer6_outputs(4081) <= not(layer5_outputs(2257));
    layer6_outputs(4082) <= not((layer5_outputs(197)) or (layer5_outputs(3660)));
    layer6_outputs(4083) <= (layer5_outputs(1209)) and not (layer5_outputs(5108));
    layer6_outputs(4084) <= not(layer5_outputs(4975));
    layer6_outputs(4085) <= not(layer5_outputs(1368));
    layer6_outputs(4086) <= not((layer5_outputs(615)) or (layer5_outputs(3583)));
    layer6_outputs(4087) <= not(layer5_outputs(4639));
    layer6_outputs(4088) <= (layer5_outputs(4667)) and not (layer5_outputs(1380));
    layer6_outputs(4089) <= not(layer5_outputs(640));
    layer6_outputs(4090) <= layer5_outputs(4936);
    layer6_outputs(4091) <= (layer5_outputs(105)) xor (layer5_outputs(1420));
    layer6_outputs(4092) <= not(layer5_outputs(3069));
    layer6_outputs(4093) <= not((layer5_outputs(1504)) xor (layer5_outputs(4304)));
    layer6_outputs(4094) <= not((layer5_outputs(1064)) or (layer5_outputs(2173)));
    layer6_outputs(4095) <= not(layer5_outputs(2247));
    layer6_outputs(4096) <= (layer5_outputs(820)) or (layer5_outputs(344));
    layer6_outputs(4097) <= not((layer5_outputs(850)) xor (layer5_outputs(4415)));
    layer6_outputs(4098) <= not((layer5_outputs(4059)) xor (layer5_outputs(632)));
    layer6_outputs(4099) <= (layer5_outputs(4981)) or (layer5_outputs(390));
    layer6_outputs(4100) <= not(layer5_outputs(3232)) or (layer5_outputs(1706));
    layer6_outputs(4101) <= not(layer5_outputs(2489));
    layer6_outputs(4102) <= not((layer5_outputs(4789)) or (layer5_outputs(4120)));
    layer6_outputs(4103) <= layer5_outputs(1320);
    layer6_outputs(4104) <= not(layer5_outputs(3328));
    layer6_outputs(4105) <= not((layer5_outputs(203)) and (layer5_outputs(1041)));
    layer6_outputs(4106) <= not(layer5_outputs(4028));
    layer6_outputs(4107) <= not(layer5_outputs(3940)) or (layer5_outputs(1197));
    layer6_outputs(4108) <= layer5_outputs(4176);
    layer6_outputs(4109) <= (layer5_outputs(4493)) and not (layer5_outputs(207));
    layer6_outputs(4110) <= layer5_outputs(192);
    layer6_outputs(4111) <= layer5_outputs(362);
    layer6_outputs(4112) <= not(layer5_outputs(2810));
    layer6_outputs(4113) <= not(layer5_outputs(4129));
    layer6_outputs(4114) <= layer5_outputs(0);
    layer6_outputs(4115) <= layer5_outputs(3959);
    layer6_outputs(4116) <= layer5_outputs(3802);
    layer6_outputs(4117) <= (layer5_outputs(1243)) and not (layer5_outputs(2853));
    layer6_outputs(4118) <= layer5_outputs(1634);
    layer6_outputs(4119) <= not((layer5_outputs(1490)) xor (layer5_outputs(664)));
    layer6_outputs(4120) <= layer5_outputs(5012);
    layer6_outputs(4121) <= layer5_outputs(2035);
    layer6_outputs(4122) <= not(layer5_outputs(2613));
    layer6_outputs(4123) <= layer5_outputs(4208);
    layer6_outputs(4124) <= layer5_outputs(1158);
    layer6_outputs(4125) <= not(layer5_outputs(3572));
    layer6_outputs(4126) <= layer5_outputs(3992);
    layer6_outputs(4127) <= not((layer5_outputs(4480)) xor (layer5_outputs(1265)));
    layer6_outputs(4128) <= not((layer5_outputs(2501)) xor (layer5_outputs(2428)));
    layer6_outputs(4129) <= layer5_outputs(2746);
    layer6_outputs(4130) <= (layer5_outputs(470)) and not (layer5_outputs(383));
    layer6_outputs(4131) <= layer5_outputs(1734);
    layer6_outputs(4132) <= not((layer5_outputs(3813)) and (layer5_outputs(3837)));
    layer6_outputs(4133) <= not(layer5_outputs(149));
    layer6_outputs(4134) <= not((layer5_outputs(1054)) or (layer5_outputs(374)));
    layer6_outputs(4135) <= not((layer5_outputs(2243)) xor (layer5_outputs(2055)));
    layer6_outputs(4136) <= not(layer5_outputs(888));
    layer6_outputs(4137) <= not(layer5_outputs(4262)) or (layer5_outputs(4287));
    layer6_outputs(4138) <= layer5_outputs(3929);
    layer6_outputs(4139) <= layer5_outputs(3991);
    layer6_outputs(4140) <= layer5_outputs(3710);
    layer6_outputs(4141) <= not(layer5_outputs(4932)) or (layer5_outputs(2393));
    layer6_outputs(4142) <= not((layer5_outputs(617)) or (layer5_outputs(4962)));
    layer6_outputs(4143) <= not(layer5_outputs(990));
    layer6_outputs(4144) <= not(layer5_outputs(4544));
    layer6_outputs(4145) <= (layer5_outputs(1376)) xor (layer5_outputs(2754));
    layer6_outputs(4146) <= (layer5_outputs(4143)) and not (layer5_outputs(2776));
    layer6_outputs(4147) <= layer5_outputs(936);
    layer6_outputs(4148) <= not((layer5_outputs(4514)) or (layer5_outputs(2172)));
    layer6_outputs(4149) <= layer5_outputs(3582);
    layer6_outputs(4150) <= not(layer5_outputs(2535));
    layer6_outputs(4151) <= layer5_outputs(3967);
    layer6_outputs(4152) <= not((layer5_outputs(4151)) xor (layer5_outputs(1500)));
    layer6_outputs(4153) <= not(layer5_outputs(1686));
    layer6_outputs(4154) <= not(layer5_outputs(4491));
    layer6_outputs(4155) <= not(layer5_outputs(4972));
    layer6_outputs(4156) <= not(layer5_outputs(1340));
    layer6_outputs(4157) <= not(layer5_outputs(1510));
    layer6_outputs(4158) <= layer5_outputs(965);
    layer6_outputs(4159) <= not(layer5_outputs(5052));
    layer6_outputs(4160) <= layer5_outputs(4644);
    layer6_outputs(4161) <= layer5_outputs(1042);
    layer6_outputs(4162) <= not((layer5_outputs(4473)) xor (layer5_outputs(1991)));
    layer6_outputs(4163) <= layer5_outputs(653);
    layer6_outputs(4164) <= not(layer5_outputs(4660));
    layer6_outputs(4165) <= not(layer5_outputs(3081));
    layer6_outputs(4166) <= not(layer5_outputs(937));
    layer6_outputs(4167) <= not(layer5_outputs(2710));
    layer6_outputs(4168) <= layer5_outputs(4573);
    layer6_outputs(4169) <= layer5_outputs(641);
    layer6_outputs(4170) <= (layer5_outputs(3820)) xor (layer5_outputs(3578));
    layer6_outputs(4171) <= not(layer5_outputs(2386));
    layer6_outputs(4172) <= not(layer5_outputs(3775));
    layer6_outputs(4173) <= layer5_outputs(753);
    layer6_outputs(4174) <= layer5_outputs(1327);
    layer6_outputs(4175) <= layer5_outputs(4069);
    layer6_outputs(4176) <= not((layer5_outputs(957)) or (layer5_outputs(3638)));
    layer6_outputs(4177) <= (layer5_outputs(3889)) or (layer5_outputs(1669));
    layer6_outputs(4178) <= not(layer5_outputs(4934));
    layer6_outputs(4179) <= not(layer5_outputs(4445)) or (layer5_outputs(1772));
    layer6_outputs(4180) <= layer5_outputs(2126);
    layer6_outputs(4181) <= not(layer5_outputs(3429));
    layer6_outputs(4182) <= not(layer5_outputs(735));
    layer6_outputs(4183) <= '0';
    layer6_outputs(4184) <= layer5_outputs(1607);
    layer6_outputs(4185) <= not((layer5_outputs(2683)) or (layer5_outputs(651)));
    layer6_outputs(4186) <= not((layer5_outputs(2456)) xor (layer5_outputs(3550)));
    layer6_outputs(4187) <= layer5_outputs(924);
    layer6_outputs(4188) <= layer5_outputs(2602);
    layer6_outputs(4189) <= not(layer5_outputs(591));
    layer6_outputs(4190) <= (layer5_outputs(2610)) and not (layer5_outputs(634));
    layer6_outputs(4191) <= not(layer5_outputs(1127)) or (layer5_outputs(4112));
    layer6_outputs(4192) <= not((layer5_outputs(4341)) and (layer5_outputs(2344)));
    layer6_outputs(4193) <= not(layer5_outputs(1943));
    layer6_outputs(4194) <= not(layer5_outputs(1000));
    layer6_outputs(4195) <= layer5_outputs(3442);
    layer6_outputs(4196) <= not(layer5_outputs(3036));
    layer6_outputs(4197) <= layer5_outputs(4714);
    layer6_outputs(4198) <= (layer5_outputs(3077)) and (layer5_outputs(3337));
    layer6_outputs(4199) <= not(layer5_outputs(4781));
    layer6_outputs(4200) <= '1';
    layer6_outputs(4201) <= (layer5_outputs(1905)) and not (layer5_outputs(4992));
    layer6_outputs(4202) <= (layer5_outputs(2091)) or (layer5_outputs(1426));
    layer6_outputs(4203) <= (layer5_outputs(109)) or (layer5_outputs(4852));
    layer6_outputs(4204) <= layer5_outputs(830);
    layer6_outputs(4205) <= '1';
    layer6_outputs(4206) <= layer5_outputs(1835);
    layer6_outputs(4207) <= not(layer5_outputs(3648));
    layer6_outputs(4208) <= not(layer5_outputs(4104)) or (layer5_outputs(4392));
    layer6_outputs(4209) <= (layer5_outputs(321)) and not (layer5_outputs(1469));
    layer6_outputs(4210) <= not(layer5_outputs(333));
    layer6_outputs(4211) <= not(layer5_outputs(206));
    layer6_outputs(4212) <= (layer5_outputs(1017)) xor (layer5_outputs(1402));
    layer6_outputs(4213) <= not(layer5_outputs(1138));
    layer6_outputs(4214) <= layer5_outputs(3864);
    layer6_outputs(4215) <= not(layer5_outputs(164)) or (layer5_outputs(457));
    layer6_outputs(4216) <= not(layer5_outputs(3176)) or (layer5_outputs(1162));
    layer6_outputs(4217) <= layer5_outputs(1287);
    layer6_outputs(4218) <= not((layer5_outputs(1340)) xor (layer5_outputs(4979)));
    layer6_outputs(4219) <= (layer5_outputs(4105)) and not (layer5_outputs(4893));
    layer6_outputs(4220) <= layer5_outputs(1462);
    layer6_outputs(4221) <= (layer5_outputs(2814)) and (layer5_outputs(639));
    layer6_outputs(4222) <= layer5_outputs(3039);
    layer6_outputs(4223) <= (layer5_outputs(96)) xor (layer5_outputs(402));
    layer6_outputs(4224) <= layer5_outputs(3471);
    layer6_outputs(4225) <= (layer5_outputs(1659)) xor (layer5_outputs(659));
    layer6_outputs(4226) <= not(layer5_outputs(393));
    layer6_outputs(4227) <= (layer5_outputs(323)) xor (layer5_outputs(3284));
    layer6_outputs(4228) <= layer5_outputs(4831);
    layer6_outputs(4229) <= not((layer5_outputs(1300)) xor (layer5_outputs(2882)));
    layer6_outputs(4230) <= not(layer5_outputs(973));
    layer6_outputs(4231) <= not((layer5_outputs(752)) xor (layer5_outputs(3823)));
    layer6_outputs(4232) <= not((layer5_outputs(1527)) xor (layer5_outputs(1777)));
    layer6_outputs(4233) <= layer5_outputs(235);
    layer6_outputs(4234) <= layer5_outputs(4952);
    layer6_outputs(4235) <= (layer5_outputs(4113)) or (layer5_outputs(4306));
    layer6_outputs(4236) <= not(layer5_outputs(827)) or (layer5_outputs(4321));
    layer6_outputs(4237) <= layer5_outputs(3495);
    layer6_outputs(4238) <= not(layer5_outputs(4211));
    layer6_outputs(4239) <= not(layer5_outputs(4943));
    layer6_outputs(4240) <= layer5_outputs(374);
    layer6_outputs(4241) <= layer5_outputs(305);
    layer6_outputs(4242) <= not((layer5_outputs(2916)) and (layer5_outputs(263)));
    layer6_outputs(4243) <= not((layer5_outputs(2415)) xor (layer5_outputs(2228)));
    layer6_outputs(4244) <= (layer5_outputs(5111)) and not (layer5_outputs(2421));
    layer6_outputs(4245) <= not((layer5_outputs(1026)) or (layer5_outputs(2097)));
    layer6_outputs(4246) <= not((layer5_outputs(4242)) xor (layer5_outputs(2088)));
    layer6_outputs(4247) <= not(layer5_outputs(4865));
    layer6_outputs(4248) <= (layer5_outputs(2969)) and not (layer5_outputs(4051));
    layer6_outputs(4249) <= layer5_outputs(4823);
    layer6_outputs(4250) <= (layer5_outputs(4742)) xor (layer5_outputs(1660));
    layer6_outputs(4251) <= not(layer5_outputs(649));
    layer6_outputs(4252) <= not((layer5_outputs(807)) xor (layer5_outputs(2391)));
    layer6_outputs(4253) <= not((layer5_outputs(3524)) xor (layer5_outputs(691)));
    layer6_outputs(4254) <= not(layer5_outputs(3240));
    layer6_outputs(4255) <= (layer5_outputs(2907)) or (layer5_outputs(633));
    layer6_outputs(4256) <= (layer5_outputs(4964)) xor (layer5_outputs(2067));
    layer6_outputs(4257) <= (layer5_outputs(2273)) and not (layer5_outputs(2966));
    layer6_outputs(4258) <= not(layer5_outputs(441));
    layer6_outputs(4259) <= not(layer5_outputs(1814));
    layer6_outputs(4260) <= (layer5_outputs(5064)) xor (layer5_outputs(713));
    layer6_outputs(4261) <= not(layer5_outputs(4238));
    layer6_outputs(4262) <= not(layer5_outputs(4498)) or (layer5_outputs(1460));
    layer6_outputs(4263) <= layer5_outputs(3164);
    layer6_outputs(4264) <= not(layer5_outputs(1945));
    layer6_outputs(4265) <= layer5_outputs(3687);
    layer6_outputs(4266) <= not(layer5_outputs(1564));
    layer6_outputs(4267) <= (layer5_outputs(3229)) xor (layer5_outputs(2744));
    layer6_outputs(4268) <= layer5_outputs(3683);
    layer6_outputs(4269) <= not((layer5_outputs(136)) xor (layer5_outputs(4826)));
    layer6_outputs(4270) <= (layer5_outputs(2069)) xor (layer5_outputs(4786));
    layer6_outputs(4271) <= layer5_outputs(1668);
    layer6_outputs(4272) <= layer5_outputs(1544);
    layer6_outputs(4273) <= (layer5_outputs(4223)) xor (layer5_outputs(1783));
    layer6_outputs(4274) <= not(layer5_outputs(1146));
    layer6_outputs(4275) <= layer5_outputs(448);
    layer6_outputs(4276) <= layer5_outputs(410);
    layer6_outputs(4277) <= not(layer5_outputs(663));
    layer6_outputs(4278) <= not((layer5_outputs(2179)) xor (layer5_outputs(1077)));
    layer6_outputs(4279) <= not(layer5_outputs(4285));
    layer6_outputs(4280) <= (layer5_outputs(1252)) xor (layer5_outputs(4897));
    layer6_outputs(4281) <= not(layer5_outputs(1062));
    layer6_outputs(4282) <= (layer5_outputs(4149)) xor (layer5_outputs(844));
    layer6_outputs(4283) <= layer5_outputs(820);
    layer6_outputs(4284) <= layer5_outputs(2305);
    layer6_outputs(4285) <= '1';
    layer6_outputs(4286) <= not(layer5_outputs(2881));
    layer6_outputs(4287) <= not(layer5_outputs(1592));
    layer6_outputs(4288) <= not((layer5_outputs(724)) xor (layer5_outputs(606)));
    layer6_outputs(4289) <= not(layer5_outputs(1076));
    layer6_outputs(4290) <= (layer5_outputs(221)) xor (layer5_outputs(47));
    layer6_outputs(4291) <= layer5_outputs(2749);
    layer6_outputs(4292) <= (layer5_outputs(883)) and not (layer5_outputs(2769));
    layer6_outputs(4293) <= not((layer5_outputs(1078)) or (layer5_outputs(271)));
    layer6_outputs(4294) <= (layer5_outputs(852)) and not (layer5_outputs(2954));
    layer6_outputs(4295) <= not(layer5_outputs(1088)) or (layer5_outputs(1378));
    layer6_outputs(4296) <= layer5_outputs(2982);
    layer6_outputs(4297) <= not((layer5_outputs(1607)) or (layer5_outputs(48)));
    layer6_outputs(4298) <= layer5_outputs(2388);
    layer6_outputs(4299) <= not(layer5_outputs(2834)) or (layer5_outputs(3261));
    layer6_outputs(4300) <= not(layer5_outputs(3012));
    layer6_outputs(4301) <= (layer5_outputs(4988)) and (layer5_outputs(2896));
    layer6_outputs(4302) <= (layer5_outputs(2748)) or (layer5_outputs(4399));
    layer6_outputs(4303) <= not((layer5_outputs(4890)) and (layer5_outputs(2482)));
    layer6_outputs(4304) <= not(layer5_outputs(2614)) or (layer5_outputs(5061));
    layer6_outputs(4305) <= not(layer5_outputs(5087));
    layer6_outputs(4306) <= (layer5_outputs(2090)) or (layer5_outputs(4602));
    layer6_outputs(4307) <= layer5_outputs(767);
    layer6_outputs(4308) <= (layer5_outputs(3515)) and not (layer5_outputs(1181));
    layer6_outputs(4309) <= not(layer5_outputs(3090));
    layer6_outputs(4310) <= not((layer5_outputs(555)) or (layer5_outputs(2050)));
    layer6_outputs(4311) <= not(layer5_outputs(3898));
    layer6_outputs(4312) <= not((layer5_outputs(779)) xor (layer5_outputs(1723)));
    layer6_outputs(4313) <= (layer5_outputs(3995)) xor (layer5_outputs(4345));
    layer6_outputs(4314) <= (layer5_outputs(152)) and (layer5_outputs(4334));
    layer6_outputs(4315) <= layer5_outputs(4106);
    layer6_outputs(4316) <= not(layer5_outputs(808));
    layer6_outputs(4317) <= '1';
    layer6_outputs(4318) <= (layer5_outputs(3329)) and (layer5_outputs(2668));
    layer6_outputs(4319) <= not(layer5_outputs(2855));
    layer6_outputs(4320) <= not(layer5_outputs(3822));
    layer6_outputs(4321) <= layer5_outputs(738);
    layer6_outputs(4322) <= layer5_outputs(3604);
    layer6_outputs(4323) <= layer5_outputs(167);
    layer6_outputs(4324) <= layer5_outputs(3353);
    layer6_outputs(4325) <= not((layer5_outputs(2502)) xor (layer5_outputs(2447)));
    layer6_outputs(4326) <= (layer5_outputs(4164)) and not (layer5_outputs(4017));
    layer6_outputs(4327) <= not(layer5_outputs(3369));
    layer6_outputs(4328) <= not(layer5_outputs(3795));
    layer6_outputs(4329) <= not((layer5_outputs(3993)) xor (layer5_outputs(2117)));
    layer6_outputs(4330) <= layer5_outputs(285);
    layer6_outputs(4331) <= layer5_outputs(4423);
    layer6_outputs(4332) <= not((layer5_outputs(3401)) or (layer5_outputs(4200)));
    layer6_outputs(4333) <= not(layer5_outputs(882));
    layer6_outputs(4334) <= not(layer5_outputs(2028));
    layer6_outputs(4335) <= layer5_outputs(3697);
    layer6_outputs(4336) <= layer5_outputs(822);
    layer6_outputs(4337) <= layer5_outputs(2089);
    layer6_outputs(4338) <= not(layer5_outputs(471)) or (layer5_outputs(1552));
    layer6_outputs(4339) <= not(layer5_outputs(4688));
    layer6_outputs(4340) <= (layer5_outputs(2502)) and not (layer5_outputs(609));
    layer6_outputs(4341) <= layer5_outputs(872);
    layer6_outputs(4342) <= not(layer5_outputs(3494));
    layer6_outputs(4343) <= not(layer5_outputs(1346));
    layer6_outputs(4344) <= not(layer5_outputs(478));
    layer6_outputs(4345) <= layer5_outputs(1191);
    layer6_outputs(4346) <= not(layer5_outputs(2812)) or (layer5_outputs(4412));
    layer6_outputs(4347) <= not(layer5_outputs(3816)) or (layer5_outputs(2980));
    layer6_outputs(4348) <= not(layer5_outputs(2845));
    layer6_outputs(4349) <= not(layer5_outputs(559));
    layer6_outputs(4350) <= not(layer5_outputs(1466));
    layer6_outputs(4351) <= not(layer5_outputs(4213));
    layer6_outputs(4352) <= (layer5_outputs(2385)) and not (layer5_outputs(766));
    layer6_outputs(4353) <= layer5_outputs(5070);
    layer6_outputs(4354) <= (layer5_outputs(1844)) or (layer5_outputs(3186));
    layer6_outputs(4355) <= layer5_outputs(1121);
    layer6_outputs(4356) <= not(layer5_outputs(1539));
    layer6_outputs(4357) <= not(layer5_outputs(2348));
    layer6_outputs(4358) <= not(layer5_outputs(3889));
    layer6_outputs(4359) <= not((layer5_outputs(962)) xor (layer5_outputs(3652)));
    layer6_outputs(4360) <= (layer5_outputs(5106)) and not (layer5_outputs(560));
    layer6_outputs(4361) <= (layer5_outputs(4193)) and not (layer5_outputs(1941));
    layer6_outputs(4362) <= (layer5_outputs(275)) or (layer5_outputs(551));
    layer6_outputs(4363) <= layer5_outputs(5);
    layer6_outputs(4364) <= layer5_outputs(834);
    layer6_outputs(4365) <= not(layer5_outputs(2446));
    layer6_outputs(4366) <= not(layer5_outputs(832));
    layer6_outputs(4367) <= layer5_outputs(711);
    layer6_outputs(4368) <= not(layer5_outputs(560));
    layer6_outputs(4369) <= not(layer5_outputs(513));
    layer6_outputs(4370) <= not(layer5_outputs(1889));
    layer6_outputs(4371) <= not((layer5_outputs(1645)) or (layer5_outputs(4088)));
    layer6_outputs(4372) <= not((layer5_outputs(2806)) and (layer5_outputs(4902)));
    layer6_outputs(4373) <= not((layer5_outputs(422)) and (layer5_outputs(4068)));
    layer6_outputs(4374) <= layer5_outputs(944);
    layer6_outputs(4375) <= not(layer5_outputs(2684));
    layer6_outputs(4376) <= not((layer5_outputs(2377)) xor (layer5_outputs(2811)));
    layer6_outputs(4377) <= not(layer5_outputs(2641)) or (layer5_outputs(1823));
    layer6_outputs(4378) <= layer5_outputs(324);
    layer6_outputs(4379) <= layer5_outputs(4591);
    layer6_outputs(4380) <= layer5_outputs(4037);
    layer6_outputs(4381) <= not(layer5_outputs(2422));
    layer6_outputs(4382) <= not(layer5_outputs(3444)) or (layer5_outputs(1526));
    layer6_outputs(4383) <= not(layer5_outputs(3657));
    layer6_outputs(4384) <= not(layer5_outputs(1643));
    layer6_outputs(4385) <= (layer5_outputs(593)) and not (layer5_outputs(2782));
    layer6_outputs(4386) <= not((layer5_outputs(393)) and (layer5_outputs(526)));
    layer6_outputs(4387) <= not((layer5_outputs(4027)) and (layer5_outputs(1156)));
    layer6_outputs(4388) <= layer5_outputs(4866);
    layer6_outputs(4389) <= not(layer5_outputs(2690));
    layer6_outputs(4390) <= (layer5_outputs(1874)) xor (layer5_outputs(387));
    layer6_outputs(4391) <= not((layer5_outputs(250)) xor (layer5_outputs(2780)));
    layer6_outputs(4392) <= not((layer5_outputs(5088)) xor (layer5_outputs(3426)));
    layer6_outputs(4393) <= not(layer5_outputs(341)) or (layer5_outputs(840));
    layer6_outputs(4394) <= not(layer5_outputs(3360)) or (layer5_outputs(437));
    layer6_outputs(4395) <= (layer5_outputs(4784)) xor (layer5_outputs(1130));
    layer6_outputs(4396) <= not(layer5_outputs(3150)) or (layer5_outputs(3002));
    layer6_outputs(4397) <= (layer5_outputs(825)) and (layer5_outputs(2604));
    layer6_outputs(4398) <= not(layer5_outputs(4753));
    layer6_outputs(4399) <= not(layer5_outputs(1399));
    layer6_outputs(4400) <= layer5_outputs(928);
    layer6_outputs(4401) <= not(layer5_outputs(1561));
    layer6_outputs(4402) <= not(layer5_outputs(3145)) or (layer5_outputs(2661));
    layer6_outputs(4403) <= layer5_outputs(3006);
    layer6_outputs(4404) <= layer5_outputs(196);
    layer6_outputs(4405) <= (layer5_outputs(3351)) and (layer5_outputs(2049));
    layer6_outputs(4406) <= not((layer5_outputs(3430)) and (layer5_outputs(3796)));
    layer6_outputs(4407) <= layer5_outputs(4580);
    layer6_outputs(4408) <= (layer5_outputs(2732)) xor (layer5_outputs(35));
    layer6_outputs(4409) <= not(layer5_outputs(4442));
    layer6_outputs(4410) <= not((layer5_outputs(2133)) xor (layer5_outputs(607)));
    layer6_outputs(4411) <= (layer5_outputs(515)) or (layer5_outputs(3419));
    layer6_outputs(4412) <= '0';
    layer6_outputs(4413) <= layer5_outputs(497);
    layer6_outputs(4414) <= not((layer5_outputs(3616)) or (layer5_outputs(3425)));
    layer6_outputs(4415) <= (layer5_outputs(1843)) and not (layer5_outputs(2690));
    layer6_outputs(4416) <= layer5_outputs(1329);
    layer6_outputs(4417) <= not(layer5_outputs(2026));
    layer6_outputs(4418) <= not(layer5_outputs(1779)) or (layer5_outputs(4475));
    layer6_outputs(4419) <= not(layer5_outputs(146));
    layer6_outputs(4420) <= (layer5_outputs(3058)) and not (layer5_outputs(3862));
    layer6_outputs(4421) <= layer5_outputs(3113);
    layer6_outputs(4422) <= layer5_outputs(4283);
    layer6_outputs(4423) <= layer5_outputs(4124);
    layer6_outputs(4424) <= layer5_outputs(4537);
    layer6_outputs(4425) <= not(layer5_outputs(2847));
    layer6_outputs(4426) <= '0';
    layer6_outputs(4427) <= (layer5_outputs(1638)) and not (layer5_outputs(406));
    layer6_outputs(4428) <= not((layer5_outputs(3774)) or (layer5_outputs(4052)));
    layer6_outputs(4429) <= not(layer5_outputs(2684)) or (layer5_outputs(1434));
    layer6_outputs(4430) <= (layer5_outputs(3690)) xor (layer5_outputs(962));
    layer6_outputs(4431) <= not(layer5_outputs(3322)) or (layer5_outputs(537));
    layer6_outputs(4432) <= not(layer5_outputs(3094));
    layer6_outputs(4433) <= layer5_outputs(2116);
    layer6_outputs(4434) <= '0';
    layer6_outputs(4435) <= not((layer5_outputs(532)) or (layer5_outputs(1430)));
    layer6_outputs(4436) <= layer5_outputs(4922);
    layer6_outputs(4437) <= not(layer5_outputs(3498));
    layer6_outputs(4438) <= (layer5_outputs(4072)) or (layer5_outputs(667));
    layer6_outputs(4439) <= not(layer5_outputs(4479));
    layer6_outputs(4440) <= (layer5_outputs(4980)) and (layer5_outputs(1580));
    layer6_outputs(4441) <= layer5_outputs(2753);
    layer6_outputs(4442) <= not((layer5_outputs(3501)) or (layer5_outputs(1246)));
    layer6_outputs(4443) <= (layer5_outputs(3226)) and (layer5_outputs(2483));
    layer6_outputs(4444) <= not(layer5_outputs(3450));
    layer6_outputs(4445) <= layer5_outputs(3259);
    layer6_outputs(4446) <= (layer5_outputs(1234)) and not (layer5_outputs(4490));
    layer6_outputs(4447) <= not(layer5_outputs(402));
    layer6_outputs(4448) <= layer5_outputs(1885);
    layer6_outputs(4449) <= layer5_outputs(470);
    layer6_outputs(4450) <= not((layer5_outputs(2979)) and (layer5_outputs(5028)));
    layer6_outputs(4451) <= (layer5_outputs(2713)) and (layer5_outputs(1998));
    layer6_outputs(4452) <= layer5_outputs(1553);
    layer6_outputs(4453) <= not(layer5_outputs(4107));
    layer6_outputs(4454) <= layer5_outputs(692);
    layer6_outputs(4455) <= (layer5_outputs(3746)) and not (layer5_outputs(725));
    layer6_outputs(4456) <= not(layer5_outputs(4870)) or (layer5_outputs(4004));
    layer6_outputs(4457) <= (layer5_outputs(1082)) xor (layer5_outputs(4800));
    layer6_outputs(4458) <= (layer5_outputs(1415)) xor (layer5_outputs(4183));
    layer6_outputs(4459) <= (layer5_outputs(714)) and not (layer5_outputs(2288));
    layer6_outputs(4460) <= not(layer5_outputs(1190)) or (layer5_outputs(1022));
    layer6_outputs(4461) <= not(layer5_outputs(5093));
    layer6_outputs(4462) <= layer5_outputs(3969);
    layer6_outputs(4463) <= layer5_outputs(2071);
    layer6_outputs(4464) <= (layer5_outputs(5005)) and not (layer5_outputs(2404));
    layer6_outputs(4465) <= not((layer5_outputs(2270)) and (layer5_outputs(427)));
    layer6_outputs(4466) <= not(layer5_outputs(3725));
    layer6_outputs(4467) <= not(layer5_outputs(3652));
    layer6_outputs(4468) <= not(layer5_outputs(2746));
    layer6_outputs(4469) <= (layer5_outputs(603)) xor (layer5_outputs(4095));
    layer6_outputs(4470) <= not((layer5_outputs(4141)) and (layer5_outputs(1333)));
    layer6_outputs(4471) <= not(layer5_outputs(2108));
    layer6_outputs(4472) <= layer5_outputs(616);
    layer6_outputs(4473) <= not((layer5_outputs(3559)) xor (layer5_outputs(3327)));
    layer6_outputs(4474) <= layer5_outputs(116);
    layer6_outputs(4475) <= (layer5_outputs(1283)) xor (layer5_outputs(2082));
    layer6_outputs(4476) <= layer5_outputs(2236);
    layer6_outputs(4477) <= layer5_outputs(1916);
    layer6_outputs(4478) <= (layer5_outputs(467)) and not (layer5_outputs(481));
    layer6_outputs(4479) <= not((layer5_outputs(4311)) and (layer5_outputs(4352)));
    layer6_outputs(4480) <= not(layer5_outputs(897));
    layer6_outputs(4481) <= not((layer5_outputs(2145)) xor (layer5_outputs(1456)));
    layer6_outputs(4482) <= not(layer5_outputs(4732));
    layer6_outputs(4483) <= not((layer5_outputs(3935)) xor (layer5_outputs(1910)));
    layer6_outputs(4484) <= (layer5_outputs(17)) and not (layer5_outputs(3729));
    layer6_outputs(4485) <= not(layer5_outputs(3389));
    layer6_outputs(4486) <= not(layer5_outputs(2397));
    layer6_outputs(4487) <= layer5_outputs(2528);
    layer6_outputs(4488) <= not((layer5_outputs(4067)) and (layer5_outputs(58)));
    layer6_outputs(4489) <= not((layer5_outputs(1927)) xor (layer5_outputs(3509)));
    layer6_outputs(4490) <= layer5_outputs(1584);
    layer6_outputs(4491) <= not(layer5_outputs(92)) or (layer5_outputs(1283));
    layer6_outputs(4492) <= layer5_outputs(2168);
    layer6_outputs(4493) <= not((layer5_outputs(5043)) xor (layer5_outputs(1003)));
    layer6_outputs(4494) <= layer5_outputs(771);
    layer6_outputs(4495) <= layer5_outputs(3469);
    layer6_outputs(4496) <= (layer5_outputs(3261)) or (layer5_outputs(929));
    layer6_outputs(4497) <= not((layer5_outputs(482)) xor (layer5_outputs(4315)));
    layer6_outputs(4498) <= not(layer5_outputs(4234));
    layer6_outputs(4499) <= not(layer5_outputs(53)) or (layer5_outputs(4675));
    layer6_outputs(4500) <= layer5_outputs(4543);
    layer6_outputs(4501) <= not(layer5_outputs(1635)) or (layer5_outputs(1514));
    layer6_outputs(4502) <= (layer5_outputs(567)) and (layer5_outputs(5));
    layer6_outputs(4503) <= not(layer5_outputs(1755));
    layer6_outputs(4504) <= not(layer5_outputs(154));
    layer6_outputs(4505) <= layer5_outputs(3645);
    layer6_outputs(4506) <= not(layer5_outputs(1477));
    layer6_outputs(4507) <= not(layer5_outputs(4370));
    layer6_outputs(4508) <= (layer5_outputs(3377)) or (layer5_outputs(4832));
    layer6_outputs(4509) <= (layer5_outputs(3769)) or (layer5_outputs(2328));
    layer6_outputs(4510) <= layer5_outputs(1120);
    layer6_outputs(4511) <= not(layer5_outputs(2830));
    layer6_outputs(4512) <= not(layer5_outputs(3090));
    layer6_outputs(4513) <= not(layer5_outputs(3806));
    layer6_outputs(4514) <= not((layer5_outputs(2337)) xor (layer5_outputs(2575)));
    layer6_outputs(4515) <= not(layer5_outputs(249));
    layer6_outputs(4516) <= (layer5_outputs(605)) and not (layer5_outputs(413));
    layer6_outputs(4517) <= not(layer5_outputs(3306));
    layer6_outputs(4518) <= layer5_outputs(4655);
    layer6_outputs(4519) <= (layer5_outputs(1703)) xor (layer5_outputs(3223));
    layer6_outputs(4520) <= not(layer5_outputs(4083)) or (layer5_outputs(1541));
    layer6_outputs(4521) <= not(layer5_outputs(4166));
    layer6_outputs(4522) <= layer5_outputs(1508);
    layer6_outputs(4523) <= (layer5_outputs(913)) xor (layer5_outputs(4048));
    layer6_outputs(4524) <= not(layer5_outputs(2192));
    layer6_outputs(4525) <= not(layer5_outputs(871)) or (layer5_outputs(1095));
    layer6_outputs(4526) <= not(layer5_outputs(4878));
    layer6_outputs(4527) <= not(layer5_outputs(2715));
    layer6_outputs(4528) <= layer5_outputs(3715);
    layer6_outputs(4529) <= (layer5_outputs(2300)) or (layer5_outputs(4450));
    layer6_outputs(4530) <= not(layer5_outputs(401));
    layer6_outputs(4531) <= not((layer5_outputs(1128)) xor (layer5_outputs(3016)));
    layer6_outputs(4532) <= layer5_outputs(2105);
    layer6_outputs(4533) <= not(layer5_outputs(3562));
    layer6_outputs(4534) <= not(layer5_outputs(702));
    layer6_outputs(4535) <= not(layer5_outputs(4561));
    layer6_outputs(4536) <= not(layer5_outputs(3720)) or (layer5_outputs(809));
    layer6_outputs(4537) <= (layer5_outputs(4019)) xor (layer5_outputs(3180));
    layer6_outputs(4538) <= not((layer5_outputs(2934)) or (layer5_outputs(3087)));
    layer6_outputs(4539) <= layer5_outputs(4954);
    layer6_outputs(4540) <= not(layer5_outputs(884));
    layer6_outputs(4541) <= not((layer5_outputs(4686)) or (layer5_outputs(1637)));
    layer6_outputs(4542) <= not(layer5_outputs(2287));
    layer6_outputs(4543) <= layer5_outputs(905);
    layer6_outputs(4544) <= layer5_outputs(3708);
    layer6_outputs(4545) <= (layer5_outputs(2875)) xor (layer5_outputs(2872));
    layer6_outputs(4546) <= layer5_outputs(500);
    layer6_outputs(4547) <= (layer5_outputs(3118)) or (layer5_outputs(4503));
    layer6_outputs(4548) <= not((layer5_outputs(49)) or (layer5_outputs(1587)));
    layer6_outputs(4549) <= layer5_outputs(1970);
    layer6_outputs(4550) <= '1';
    layer6_outputs(4551) <= not(layer5_outputs(868)) or (layer5_outputs(3081));
    layer6_outputs(4552) <= layer5_outputs(4495);
    layer6_outputs(4553) <= not((layer5_outputs(838)) xor (layer5_outputs(4635)));
    layer6_outputs(4554) <= (layer5_outputs(3771)) and not (layer5_outputs(2272));
    layer6_outputs(4555) <= layer5_outputs(2480);
    layer6_outputs(4556) <= not(layer5_outputs(4051));
    layer6_outputs(4557) <= (layer5_outputs(2522)) and (layer5_outputs(3669));
    layer6_outputs(4558) <= not(layer5_outputs(4105));
    layer6_outputs(4559) <= not((layer5_outputs(5032)) xor (layer5_outputs(155)));
    layer6_outputs(4560) <= (layer5_outputs(3142)) xor (layer5_outputs(4973));
    layer6_outputs(4561) <= not(layer5_outputs(34));
    layer6_outputs(4562) <= not(layer5_outputs(4475));
    layer6_outputs(4563) <= not(layer5_outputs(2711));
    layer6_outputs(4564) <= not((layer5_outputs(3651)) xor (layer5_outputs(4434)));
    layer6_outputs(4565) <= layer5_outputs(1979);
    layer6_outputs(4566) <= not((layer5_outputs(3998)) and (layer5_outputs(4831)));
    layer6_outputs(4567) <= (layer5_outputs(1764)) or (layer5_outputs(1611));
    layer6_outputs(4568) <= not((layer5_outputs(1258)) and (layer5_outputs(1746)));
    layer6_outputs(4569) <= layer5_outputs(4000);
    layer6_outputs(4570) <= not(layer5_outputs(636)) or (layer5_outputs(5034));
    layer6_outputs(4571) <= layer5_outputs(2472);
    layer6_outputs(4572) <= not(layer5_outputs(1565));
    layer6_outputs(4573) <= not(layer5_outputs(3445));
    layer6_outputs(4574) <= not(layer5_outputs(1479));
    layer6_outputs(4575) <= not((layer5_outputs(3102)) xor (layer5_outputs(635)));
    layer6_outputs(4576) <= (layer5_outputs(3588)) and not (layer5_outputs(721));
    layer6_outputs(4577) <= (layer5_outputs(1073)) or (layer5_outputs(155));
    layer6_outputs(4578) <= (layer5_outputs(3876)) and (layer5_outputs(4938));
    layer6_outputs(4579) <= layer5_outputs(429);
    layer6_outputs(4580) <= layer5_outputs(1416);
    layer6_outputs(4581) <= '1';
    layer6_outputs(4582) <= not((layer5_outputs(2816)) or (layer5_outputs(1551)));
    layer6_outputs(4583) <= (layer5_outputs(69)) and not (layer5_outputs(3607));
    layer6_outputs(4584) <= '1';
    layer6_outputs(4585) <= not(layer5_outputs(5015));
    layer6_outputs(4586) <= not((layer5_outputs(4015)) and (layer5_outputs(5040)));
    layer6_outputs(4587) <= (layer5_outputs(1622)) and (layer5_outputs(3238));
    layer6_outputs(4588) <= (layer5_outputs(1734)) and not (layer5_outputs(3130));
    layer6_outputs(4589) <= not((layer5_outputs(1275)) and (layer5_outputs(2636)));
    layer6_outputs(4590) <= layer5_outputs(4603);
    layer6_outputs(4591) <= not(layer5_outputs(1955));
    layer6_outputs(4592) <= (layer5_outputs(149)) and not (layer5_outputs(401));
    layer6_outputs(4593) <= not(layer5_outputs(537)) or (layer5_outputs(2073));
    layer6_outputs(4594) <= '1';
    layer6_outputs(4595) <= (layer5_outputs(2891)) and (layer5_outputs(1102));
    layer6_outputs(4596) <= not((layer5_outputs(210)) or (layer5_outputs(5060)));
    layer6_outputs(4597) <= layer5_outputs(377);
    layer6_outputs(4598) <= not(layer5_outputs(2109));
    layer6_outputs(4599) <= not(layer5_outputs(3116));
    layer6_outputs(4600) <= layer5_outputs(4520);
    layer6_outputs(4601) <= layer5_outputs(4637);
    layer6_outputs(4602) <= layer5_outputs(1452);
    layer6_outputs(4603) <= layer5_outputs(2199);
    layer6_outputs(4604) <= layer5_outputs(4118);
    layer6_outputs(4605) <= layer5_outputs(2906);
    layer6_outputs(4606) <= not((layer5_outputs(2911)) xor (layer5_outputs(2545)));
    layer6_outputs(4607) <= not(layer5_outputs(1961)) or (layer5_outputs(4638));
    layer6_outputs(4608) <= not((layer5_outputs(3133)) xor (layer5_outputs(3817)));
    layer6_outputs(4609) <= not((layer5_outputs(2782)) xor (layer5_outputs(4366)));
    layer6_outputs(4610) <= not((layer5_outputs(2809)) or (layer5_outputs(2713)));
    layer6_outputs(4611) <= (layer5_outputs(458)) and not (layer5_outputs(2560));
    layer6_outputs(4612) <= not(layer5_outputs(180));
    layer6_outputs(4613) <= layer5_outputs(4046);
    layer6_outputs(4614) <= not(layer5_outputs(4180)) or (layer5_outputs(4463));
    layer6_outputs(4615) <= not(layer5_outputs(1202)) or (layer5_outputs(3019));
    layer6_outputs(4616) <= not((layer5_outputs(485)) xor (layer5_outputs(5018)));
    layer6_outputs(4617) <= not((layer5_outputs(1069)) xor (layer5_outputs(627)));
    layer6_outputs(4618) <= not(layer5_outputs(931));
    layer6_outputs(4619) <= not(layer5_outputs(1981));
    layer6_outputs(4620) <= not(layer5_outputs(1321));
    layer6_outputs(4621) <= layer5_outputs(3451);
    layer6_outputs(4622) <= not(layer5_outputs(1624));
    layer6_outputs(4623) <= layer5_outputs(507);
    layer6_outputs(4624) <= layer5_outputs(1983);
    layer6_outputs(4625) <= '0';
    layer6_outputs(4626) <= not(layer5_outputs(3288));
    layer6_outputs(4627) <= not((layer5_outputs(914)) and (layer5_outputs(118)));
    layer6_outputs(4628) <= layer5_outputs(244);
    layer6_outputs(4629) <= not(layer5_outputs(3728));
    layer6_outputs(4630) <= not((layer5_outputs(2837)) and (layer5_outputs(3374)));
    layer6_outputs(4631) <= layer5_outputs(2785);
    layer6_outputs(4632) <= (layer5_outputs(2832)) xor (layer5_outputs(2774));
    layer6_outputs(4633) <= layer5_outputs(3026);
    layer6_outputs(4634) <= not(layer5_outputs(781)) or (layer5_outputs(5065));
    layer6_outputs(4635) <= not(layer5_outputs(4819));
    layer6_outputs(4636) <= (layer5_outputs(238)) and not (layer5_outputs(689));
    layer6_outputs(4637) <= not((layer5_outputs(1594)) xor (layer5_outputs(3390)));
    layer6_outputs(4638) <= layer5_outputs(2536);
    layer6_outputs(4639) <= not(layer5_outputs(3743));
    layer6_outputs(4640) <= (layer5_outputs(3716)) or (layer5_outputs(2374));
    layer6_outputs(4641) <= not(layer5_outputs(1176));
    layer6_outputs(4642) <= not((layer5_outputs(3361)) or (layer5_outputs(4415)));
    layer6_outputs(4643) <= (layer5_outputs(1909)) and (layer5_outputs(4395));
    layer6_outputs(4644) <= not(layer5_outputs(3223)) or (layer5_outputs(5091));
    layer6_outputs(4645) <= not((layer5_outputs(2701)) or (layer5_outputs(3437)));
    layer6_outputs(4646) <= layer5_outputs(1896);
    layer6_outputs(4647) <= (layer5_outputs(4896)) xor (layer5_outputs(3008));
    layer6_outputs(4648) <= layer5_outputs(729);
    layer6_outputs(4649) <= layer5_outputs(3858);
    layer6_outputs(4650) <= not((layer5_outputs(2787)) xor (layer5_outputs(1459)));
    layer6_outputs(4651) <= (layer5_outputs(3668)) xor (layer5_outputs(5022));
    layer6_outputs(4652) <= not(layer5_outputs(4408));
    layer6_outputs(4653) <= not((layer5_outputs(5100)) or (layer5_outputs(3988)));
    layer6_outputs(4654) <= (layer5_outputs(672)) xor (layer5_outputs(4303));
    layer6_outputs(4655) <= (layer5_outputs(610)) xor (layer5_outputs(4748));
    layer6_outputs(4656) <= not(layer5_outputs(353));
    layer6_outputs(4657) <= layer5_outputs(2278);
    layer6_outputs(4658) <= (layer5_outputs(2336)) and not (layer5_outputs(5102));
    layer6_outputs(4659) <= '1';
    layer6_outputs(4660) <= (layer5_outputs(786)) and not (layer5_outputs(2486));
    layer6_outputs(4661) <= not(layer5_outputs(1356));
    layer6_outputs(4662) <= layer5_outputs(4816);
    layer6_outputs(4663) <= (layer5_outputs(38)) and (layer5_outputs(2110));
    layer6_outputs(4664) <= not((layer5_outputs(2939)) xor (layer5_outputs(2579)));
    layer6_outputs(4665) <= (layer5_outputs(1892)) xor (layer5_outputs(3402));
    layer6_outputs(4666) <= (layer5_outputs(1996)) and not (layer5_outputs(2936));
    layer6_outputs(4667) <= not(layer5_outputs(559));
    layer6_outputs(4668) <= not(layer5_outputs(3479));
    layer6_outputs(4669) <= layer5_outputs(1632);
    layer6_outputs(4670) <= not((layer5_outputs(1329)) xor (layer5_outputs(2829)));
    layer6_outputs(4671) <= (layer5_outputs(405)) and (layer5_outputs(2846));
    layer6_outputs(4672) <= not(layer5_outputs(887)) or (layer5_outputs(3517));
    layer6_outputs(4673) <= layer5_outputs(700);
    layer6_outputs(4674) <= not(layer5_outputs(2011)) or (layer5_outputs(2972));
    layer6_outputs(4675) <= (layer5_outputs(4004)) and not (layer5_outputs(3423));
    layer6_outputs(4676) <= not(layer5_outputs(2240));
    layer6_outputs(4677) <= not(layer5_outputs(1268));
    layer6_outputs(4678) <= layer5_outputs(915);
    layer6_outputs(4679) <= not(layer5_outputs(600));
    layer6_outputs(4680) <= (layer5_outputs(978)) or (layer5_outputs(2692));
    layer6_outputs(4681) <= (layer5_outputs(4233)) and not (layer5_outputs(3628));
    layer6_outputs(4682) <= layer5_outputs(1240);
    layer6_outputs(4683) <= layer5_outputs(2556);
    layer6_outputs(4684) <= (layer5_outputs(982)) and not (layer5_outputs(2346));
    layer6_outputs(4685) <= (layer5_outputs(2405)) and (layer5_outputs(2419));
    layer6_outputs(4686) <= not(layer5_outputs(2879));
    layer6_outputs(4687) <= not(layer5_outputs(207)) or (layer5_outputs(676));
    layer6_outputs(4688) <= not(layer5_outputs(914));
    layer6_outputs(4689) <= (layer5_outputs(1752)) xor (layer5_outputs(4632));
    layer6_outputs(4690) <= layer5_outputs(236);
    layer6_outputs(4691) <= not((layer5_outputs(3436)) xor (layer5_outputs(2985)));
    layer6_outputs(4692) <= layer5_outputs(1771);
    layer6_outputs(4693) <= not(layer5_outputs(1890));
    layer6_outputs(4694) <= layer5_outputs(1411);
    layer6_outputs(4695) <= not((layer5_outputs(930)) or (layer5_outputs(3520)));
    layer6_outputs(4696) <= (layer5_outputs(543)) xor (layer5_outputs(3728));
    layer6_outputs(4697) <= not((layer5_outputs(1751)) xor (layer5_outputs(4327)));
    layer6_outputs(4698) <= layer5_outputs(2224);
    layer6_outputs(4699) <= (layer5_outputs(1521)) and not (layer5_outputs(3113));
    layer6_outputs(4700) <= layer5_outputs(168);
    layer6_outputs(4701) <= not((layer5_outputs(2977)) xor (layer5_outputs(2465)));
    layer6_outputs(4702) <= not((layer5_outputs(1113)) or (layer5_outputs(2358)));
    layer6_outputs(4703) <= not(layer5_outputs(80));
    layer6_outputs(4704) <= (layer5_outputs(759)) xor (layer5_outputs(2288));
    layer6_outputs(4705) <= not((layer5_outputs(4857)) or (layer5_outputs(5025)));
    layer6_outputs(4706) <= layer5_outputs(1502);
    layer6_outputs(4707) <= not(layer5_outputs(153)) or (layer5_outputs(4512));
    layer6_outputs(4708) <= not(layer5_outputs(3904)) or (layer5_outputs(2269));
    layer6_outputs(4709) <= not((layer5_outputs(2953)) and (layer5_outputs(4708)));
    layer6_outputs(4710) <= layer5_outputs(1349);
    layer6_outputs(4711) <= (layer5_outputs(2615)) and not (layer5_outputs(3486));
    layer6_outputs(4712) <= (layer5_outputs(430)) xor (layer5_outputs(1889));
    layer6_outputs(4713) <= layer5_outputs(1533);
    layer6_outputs(4714) <= not((layer5_outputs(867)) or (layer5_outputs(1623)));
    layer6_outputs(4715) <= (layer5_outputs(2835)) and not (layer5_outputs(1919));
    layer6_outputs(4716) <= not(layer5_outputs(3203)) or (layer5_outputs(2159));
    layer6_outputs(4717) <= not(layer5_outputs(3074));
    layer6_outputs(4718) <= not((layer5_outputs(2552)) or (layer5_outputs(494)));
    layer6_outputs(4719) <= layer5_outputs(1754);
    layer6_outputs(4720) <= layer5_outputs(1901);
    layer6_outputs(4721) <= not((layer5_outputs(3643)) or (layer5_outputs(651)));
    layer6_outputs(4722) <= not(layer5_outputs(313));
    layer6_outputs(4723) <= not(layer5_outputs(1758));
    layer6_outputs(4724) <= not(layer5_outputs(4071)) or (layer5_outputs(464));
    layer6_outputs(4725) <= not(layer5_outputs(3471));
    layer6_outputs(4726) <= not((layer5_outputs(2008)) or (layer5_outputs(487)));
    layer6_outputs(4727) <= layer5_outputs(72);
    layer6_outputs(4728) <= not(layer5_outputs(3536));
    layer6_outputs(4729) <= not((layer5_outputs(866)) or (layer5_outputs(1429)));
    layer6_outputs(4730) <= not((layer5_outputs(2893)) or (layer5_outputs(2073)));
    layer6_outputs(4731) <= (layer5_outputs(2559)) xor (layer5_outputs(3711));
    layer6_outputs(4732) <= layer5_outputs(3623);
    layer6_outputs(4733) <= not(layer5_outputs(3739));
    layer6_outputs(4734) <= not(layer5_outputs(4993));
    layer6_outputs(4735) <= (layer5_outputs(3051)) and (layer5_outputs(2655));
    layer6_outputs(4736) <= not(layer5_outputs(2759));
    layer6_outputs(4737) <= layer5_outputs(3542);
    layer6_outputs(4738) <= not((layer5_outputs(784)) xor (layer5_outputs(1071)));
    layer6_outputs(4739) <= not(layer5_outputs(3875)) or (layer5_outputs(3809));
    layer6_outputs(4740) <= not((layer5_outputs(4834)) or (layer5_outputs(4518)));
    layer6_outputs(4741) <= layer5_outputs(539);
    layer6_outputs(4742) <= layer5_outputs(4092);
    layer6_outputs(4743) <= layer5_outputs(1430);
    layer6_outputs(4744) <= not(layer5_outputs(3029));
    layer6_outputs(4745) <= not(layer5_outputs(4753));
    layer6_outputs(4746) <= not((layer5_outputs(972)) xor (layer5_outputs(1214)));
    layer6_outputs(4747) <= layer5_outputs(2212);
    layer6_outputs(4748) <= not(layer5_outputs(4936)) or (layer5_outputs(2122));
    layer6_outputs(4749) <= not((layer5_outputs(3037)) xor (layer5_outputs(2171)));
    layer6_outputs(4750) <= (layer5_outputs(4955)) and not (layer5_outputs(1579));
    layer6_outputs(4751) <= not(layer5_outputs(1408));
    layer6_outputs(4752) <= not(layer5_outputs(845));
    layer6_outputs(4753) <= not(layer5_outputs(2449));
    layer6_outputs(4754) <= not(layer5_outputs(4671));
    layer6_outputs(4755) <= not(layer5_outputs(2884)) or (layer5_outputs(821));
    layer6_outputs(4756) <= not((layer5_outputs(1221)) xor (layer5_outputs(3432)));
    layer6_outputs(4757) <= not(layer5_outputs(2489));
    layer6_outputs(4758) <= not(layer5_outputs(1547));
    layer6_outputs(4759) <= layer5_outputs(1557);
    layer6_outputs(4760) <= layer5_outputs(1319);
    layer6_outputs(4761) <= not(layer5_outputs(3424));
    layer6_outputs(4762) <= not(layer5_outputs(4050));
    layer6_outputs(4763) <= layer5_outputs(3256);
    layer6_outputs(4764) <= '1';
    layer6_outputs(4765) <= (layer5_outputs(1151)) and (layer5_outputs(220));
    layer6_outputs(4766) <= layer5_outputs(967);
    layer6_outputs(4767) <= not(layer5_outputs(1898));
    layer6_outputs(4768) <= layer5_outputs(831);
    layer6_outputs(4769) <= not((layer5_outputs(3512)) or (layer5_outputs(519)));
    layer6_outputs(4770) <= layer5_outputs(4556);
    layer6_outputs(4771) <= not(layer5_outputs(5042));
    layer6_outputs(4772) <= (layer5_outputs(160)) and (layer5_outputs(5066));
    layer6_outputs(4773) <= not(layer5_outputs(2755));
    layer6_outputs(4774) <= layer5_outputs(1758);
    layer6_outputs(4775) <= not(layer5_outputs(3813));
    layer6_outputs(4776) <= not((layer5_outputs(4476)) xor (layer5_outputs(2875)));
    layer6_outputs(4777) <= layer5_outputs(5036);
    layer6_outputs(4778) <= layer5_outputs(4259);
    layer6_outputs(4779) <= not(layer5_outputs(3388));
    layer6_outputs(4780) <= layer5_outputs(3177);
    layer6_outputs(4781) <= not(layer5_outputs(2210)) or (layer5_outputs(468));
    layer6_outputs(4782) <= not((layer5_outputs(1715)) xor (layer5_outputs(4430)));
    layer6_outputs(4783) <= not(layer5_outputs(3025));
    layer6_outputs(4784) <= not(layer5_outputs(2989));
    layer6_outputs(4785) <= layer5_outputs(3208);
    layer6_outputs(4786) <= layer5_outputs(4395);
    layer6_outputs(4787) <= layer5_outputs(709);
    layer6_outputs(4788) <= not((layer5_outputs(705)) xor (layer5_outputs(1483)));
    layer6_outputs(4789) <= layer5_outputs(356);
    layer6_outputs(4790) <= not((layer5_outputs(2709)) or (layer5_outputs(525)));
    layer6_outputs(4791) <= (layer5_outputs(2821)) xor (layer5_outputs(1884));
    layer6_outputs(4792) <= layer5_outputs(2874);
    layer6_outputs(4793) <= (layer5_outputs(2253)) and not (layer5_outputs(2094));
    layer6_outputs(4794) <= not(layer5_outputs(4120)) or (layer5_outputs(3458));
    layer6_outputs(4795) <= layer5_outputs(4163);
    layer6_outputs(4796) <= layer5_outputs(2508);
    layer6_outputs(4797) <= layer5_outputs(1861);
    layer6_outputs(4798) <= (layer5_outputs(1572)) and not (layer5_outputs(3614));
    layer6_outputs(4799) <= (layer5_outputs(664)) xor (layer5_outputs(3457));
    layer6_outputs(4800) <= (layer5_outputs(2403)) xor (layer5_outputs(290));
    layer6_outputs(4801) <= layer5_outputs(3295);
    layer6_outputs(4802) <= '1';
    layer6_outputs(4803) <= (layer5_outputs(4943)) xor (layer5_outputs(2368));
    layer6_outputs(4804) <= layer5_outputs(2516);
    layer6_outputs(4805) <= not(layer5_outputs(4332));
    layer6_outputs(4806) <= (layer5_outputs(2452)) xor (layer5_outputs(2805));
    layer6_outputs(4807) <= layer5_outputs(1032);
    layer6_outputs(4808) <= not(layer5_outputs(3203)) or (layer5_outputs(1689));
    layer6_outputs(4809) <= (layer5_outputs(2735)) xor (layer5_outputs(4898));
    layer6_outputs(4810) <= not(layer5_outputs(1244));
    layer6_outputs(4811) <= layer5_outputs(4161);
    layer6_outputs(4812) <= not(layer5_outputs(4327)) or (layer5_outputs(859));
    layer6_outputs(4813) <= not((layer5_outputs(2193)) xor (layer5_outputs(2225)));
    layer6_outputs(4814) <= (layer5_outputs(1601)) and not (layer5_outputs(2028));
    layer6_outputs(4815) <= layer5_outputs(2741);
    layer6_outputs(4816) <= (layer5_outputs(754)) and not (layer5_outputs(5036));
    layer6_outputs(4817) <= (layer5_outputs(4989)) or (layer5_outputs(4630));
    layer6_outputs(4818) <= layer5_outputs(4229);
    layer6_outputs(4819) <= (layer5_outputs(3570)) or (layer5_outputs(3394));
    layer6_outputs(4820) <= not(layer5_outputs(3976));
    layer6_outputs(4821) <= not(layer5_outputs(3247));
    layer6_outputs(4822) <= not(layer5_outputs(1293)) or (layer5_outputs(1070));
    layer6_outputs(4823) <= not(layer5_outputs(2755));
    layer6_outputs(4824) <= layer5_outputs(119);
    layer6_outputs(4825) <= not(layer5_outputs(3292));
    layer6_outputs(4826) <= '0';
    layer6_outputs(4827) <= (layer5_outputs(2648)) and not (layer5_outputs(3095));
    layer6_outputs(4828) <= (layer5_outputs(1729)) and (layer5_outputs(4402));
    layer6_outputs(4829) <= (layer5_outputs(252)) or (layer5_outputs(3266));
    layer6_outputs(4830) <= layer5_outputs(825);
    layer6_outputs(4831) <= layer5_outputs(2672);
    layer6_outputs(4832) <= layer5_outputs(1485);
    layer6_outputs(4833) <= not(layer5_outputs(133));
    layer6_outputs(4834) <= not(layer5_outputs(3986));
    layer6_outputs(4835) <= not((layer5_outputs(4227)) xor (layer5_outputs(3686)));
    layer6_outputs(4836) <= (layer5_outputs(3842)) and (layer5_outputs(1923));
    layer6_outputs(4837) <= layer5_outputs(1260);
    layer6_outputs(4838) <= (layer5_outputs(454)) xor (layer5_outputs(4023));
    layer6_outputs(4839) <= not(layer5_outputs(478));
    layer6_outputs(4840) <= (layer5_outputs(1576)) and not (layer5_outputs(78));
    layer6_outputs(4841) <= not((layer5_outputs(4778)) xor (layer5_outputs(2186)));
    layer6_outputs(4842) <= not(layer5_outputs(1319));
    layer6_outputs(4843) <= layer5_outputs(1046);
    layer6_outputs(4844) <= layer5_outputs(728);
    layer6_outputs(4845) <= (layer5_outputs(520)) or (layer5_outputs(2630));
    layer6_outputs(4846) <= not(layer5_outputs(4541));
    layer6_outputs(4847) <= layer5_outputs(4758);
    layer6_outputs(4848) <= layer5_outputs(2758);
    layer6_outputs(4849) <= not((layer5_outputs(3991)) xor (layer5_outputs(434)));
    layer6_outputs(4850) <= layer5_outputs(1623);
    layer6_outputs(4851) <= (layer5_outputs(4980)) xor (layer5_outputs(2096));
    layer6_outputs(4852) <= not(layer5_outputs(840)) or (layer5_outputs(4308));
    layer6_outputs(4853) <= not((layer5_outputs(5043)) or (layer5_outputs(4297)));
    layer6_outputs(4854) <= not(layer5_outputs(3844));
    layer6_outputs(4855) <= (layer5_outputs(3534)) and not (layer5_outputs(1934));
    layer6_outputs(4856) <= layer5_outputs(2949);
    layer6_outputs(4857) <= not(layer5_outputs(2768));
    layer6_outputs(4858) <= not(layer5_outputs(2437));
    layer6_outputs(4859) <= not(layer5_outputs(3480));
    layer6_outputs(4860) <= (layer5_outputs(5096)) xor (layer5_outputs(1622));
    layer6_outputs(4861) <= not(layer5_outputs(3085));
    layer6_outputs(4862) <= (layer5_outputs(2350)) xor (layer5_outputs(4837));
    layer6_outputs(4863) <= not(layer5_outputs(2463));
    layer6_outputs(4864) <= (layer5_outputs(2206)) and not (layer5_outputs(1271));
    layer6_outputs(4865) <= (layer5_outputs(4294)) or (layer5_outputs(3671));
    layer6_outputs(4866) <= not((layer5_outputs(3308)) and (layer5_outputs(4439)));
    layer6_outputs(4867) <= layer5_outputs(2607);
    layer6_outputs(4868) <= not(layer5_outputs(80));
    layer6_outputs(4869) <= layer5_outputs(2016);
    layer6_outputs(4870) <= not(layer5_outputs(4006));
    layer6_outputs(4871) <= not((layer5_outputs(3897)) and (layer5_outputs(4376)));
    layer6_outputs(4872) <= not((layer5_outputs(1297)) xor (layer5_outputs(120)));
    layer6_outputs(4873) <= (layer5_outputs(3799)) and not (layer5_outputs(344));
    layer6_outputs(4874) <= layer5_outputs(4781);
    layer6_outputs(4875) <= layer5_outputs(4860);
    layer6_outputs(4876) <= not(layer5_outputs(5101));
    layer6_outputs(4877) <= layer5_outputs(2219);
    layer6_outputs(4878) <= not(layer5_outputs(4217)) or (layer5_outputs(3286));
    layer6_outputs(4879) <= not(layer5_outputs(2801));
    layer6_outputs(4880) <= (layer5_outputs(3914)) and (layer5_outputs(1951));
    layer6_outputs(4881) <= (layer5_outputs(3454)) or (layer5_outputs(2664));
    layer6_outputs(4882) <= not(layer5_outputs(1140));
    layer6_outputs(4883) <= layer5_outputs(3441);
    layer6_outputs(4884) <= (layer5_outputs(4054)) and not (layer5_outputs(1583));
    layer6_outputs(4885) <= not((layer5_outputs(621)) xor (layer5_outputs(4572)));
    layer6_outputs(4886) <= not(layer5_outputs(3685)) or (layer5_outputs(4243));
    layer6_outputs(4887) <= not(layer5_outputs(2418));
    layer6_outputs(4888) <= (layer5_outputs(4585)) and (layer5_outputs(858));
    layer6_outputs(4889) <= (layer5_outputs(1431)) and not (layer5_outputs(1489));
    layer6_outputs(4890) <= (layer5_outputs(452)) and not (layer5_outputs(2697));
    layer6_outputs(4891) <= (layer5_outputs(1177)) xor (layer5_outputs(3911));
    layer6_outputs(4892) <= not(layer5_outputs(1149)) or (layer5_outputs(1090));
    layer6_outputs(4893) <= not(layer5_outputs(1770));
    layer6_outputs(4894) <= layer5_outputs(3027);
    layer6_outputs(4895) <= layer5_outputs(3270);
    layer6_outputs(4896) <= not(layer5_outputs(3343));
    layer6_outputs(4897) <= layer5_outputs(4628);
    layer6_outputs(4898) <= not((layer5_outputs(3387)) xor (layer5_outputs(890)));
    layer6_outputs(4899) <= (layer5_outputs(1394)) or (layer5_outputs(382));
    layer6_outputs(4900) <= layer5_outputs(4208);
    layer6_outputs(4901) <= not((layer5_outputs(1484)) or (layer5_outputs(1100)));
    layer6_outputs(4902) <= not((layer5_outputs(1847)) xor (layer5_outputs(422)));
    layer6_outputs(4903) <= layer5_outputs(2603);
    layer6_outputs(4904) <= not(layer5_outputs(1050));
    layer6_outputs(4905) <= not(layer5_outputs(4646));
    layer6_outputs(4906) <= not((layer5_outputs(1093)) and (layer5_outputs(77)));
    layer6_outputs(4907) <= not((layer5_outputs(1692)) or (layer5_outputs(622)));
    layer6_outputs(4908) <= not(layer5_outputs(4235));
    layer6_outputs(4909) <= layer5_outputs(1060);
    layer6_outputs(4910) <= not(layer5_outputs(3075));
    layer6_outputs(4911) <= not(layer5_outputs(922));
    layer6_outputs(4912) <= not(layer5_outputs(1316));
    layer6_outputs(4913) <= not((layer5_outputs(3319)) or (layer5_outputs(3202)));
    layer6_outputs(4914) <= not(layer5_outputs(4768)) or (layer5_outputs(824));
    layer6_outputs(4915) <= not(layer5_outputs(3398));
    layer6_outputs(4916) <= not(layer5_outputs(4851));
    layer6_outputs(4917) <= not(layer5_outputs(1408)) or (layer5_outputs(3953));
    layer6_outputs(4918) <= layer5_outputs(1769);
    layer6_outputs(4919) <= not(layer5_outputs(2347));
    layer6_outputs(4920) <= layer5_outputs(414);
    layer6_outputs(4921) <= not(layer5_outputs(3234));
    layer6_outputs(4922) <= layer5_outputs(4034);
    layer6_outputs(4923) <= layer5_outputs(5024);
    layer6_outputs(4924) <= layer5_outputs(4003);
    layer6_outputs(4925) <= not(layer5_outputs(1078));
    layer6_outputs(4926) <= layer5_outputs(3463);
    layer6_outputs(4927) <= (layer5_outputs(4855)) and (layer5_outputs(4554));
    layer6_outputs(4928) <= not(layer5_outputs(1119));
    layer6_outputs(4929) <= (layer5_outputs(4562)) and (layer5_outputs(502));
    layer6_outputs(4930) <= layer5_outputs(4989);
    layer6_outputs(4931) <= not(layer5_outputs(326));
    layer6_outputs(4932) <= layer5_outputs(3283);
    layer6_outputs(4933) <= (layer5_outputs(483)) xor (layer5_outputs(1103));
    layer6_outputs(4934) <= not(layer5_outputs(3103));
    layer6_outputs(4935) <= not(layer5_outputs(2686));
    layer6_outputs(4936) <= layer5_outputs(2639);
    layer6_outputs(4937) <= layer5_outputs(4749);
    layer6_outputs(4938) <= (layer5_outputs(1557)) and not (layer5_outputs(2750));
    layer6_outputs(4939) <= layer5_outputs(1813);
    layer6_outputs(4940) <= not(layer5_outputs(999));
    layer6_outputs(4941) <= (layer5_outputs(3118)) and (layer5_outputs(4774));
    layer6_outputs(4942) <= not((layer5_outputs(4269)) xor (layer5_outputs(5080)));
    layer6_outputs(4943) <= not((layer5_outputs(4879)) xor (layer5_outputs(4344)));
    layer6_outputs(4944) <= layer5_outputs(1328);
    layer6_outputs(4945) <= (layer5_outputs(4984)) and not (layer5_outputs(4525));
    layer6_outputs(4946) <= not(layer5_outputs(3752));
    layer6_outputs(4947) <= layer5_outputs(1185);
    layer6_outputs(4948) <= '1';
    layer6_outputs(4949) <= not((layer5_outputs(4253)) and (layer5_outputs(2445)));
    layer6_outputs(4950) <= not(layer5_outputs(1992));
    layer6_outputs(4951) <= layer5_outputs(1802);
    layer6_outputs(4952) <= not((layer5_outputs(1878)) and (layer5_outputs(1614)));
    layer6_outputs(4953) <= not((layer5_outputs(3119)) and (layer5_outputs(1544)));
    layer6_outputs(4954) <= not((layer5_outputs(2233)) xor (layer5_outputs(1369)));
    layer6_outputs(4955) <= not(layer5_outputs(464)) or (layer5_outputs(2079));
    layer6_outputs(4956) <= not(layer5_outputs(25));
    layer6_outputs(4957) <= not(layer5_outputs(418));
    layer6_outputs(4958) <= layer5_outputs(1938);
    layer6_outputs(4959) <= (layer5_outputs(1355)) and (layer5_outputs(1249));
    layer6_outputs(4960) <= (layer5_outputs(5056)) or (layer5_outputs(1173));
    layer6_outputs(4961) <= layer5_outputs(4835);
    layer6_outputs(4962) <= layer5_outputs(4670);
    layer6_outputs(4963) <= not(layer5_outputs(3983)) or (layer5_outputs(4938));
    layer6_outputs(4964) <= not(layer5_outputs(2506));
    layer6_outputs(4965) <= (layer5_outputs(2054)) and (layer5_outputs(1471));
    layer6_outputs(4966) <= (layer5_outputs(1796)) or (layer5_outputs(4894));
    layer6_outputs(4967) <= (layer5_outputs(774)) and not (layer5_outputs(4451));
    layer6_outputs(4968) <= not(layer5_outputs(226)) or (layer5_outputs(4195));
    layer6_outputs(4969) <= (layer5_outputs(1326)) or (layer5_outputs(3260));
    layer6_outputs(4970) <= layer5_outputs(935);
    layer6_outputs(4971) <= (layer5_outputs(2797)) and not (layer5_outputs(4301));
    layer6_outputs(4972) <= not(layer5_outputs(7));
    layer6_outputs(4973) <= not((layer5_outputs(3920)) and (layer5_outputs(4045)));
    layer6_outputs(4974) <= (layer5_outputs(2303)) and (layer5_outputs(495));
    layer6_outputs(4975) <= not(layer5_outputs(3722));
    layer6_outputs(4976) <= '1';
    layer6_outputs(4977) <= layer5_outputs(3594);
    layer6_outputs(4978) <= not((layer5_outputs(2203)) xor (layer5_outputs(717)));
    layer6_outputs(4979) <= (layer5_outputs(2455)) xor (layer5_outputs(2772));
    layer6_outputs(4980) <= not(layer5_outputs(145));
    layer6_outputs(4981) <= layer5_outputs(2573);
    layer6_outputs(4982) <= not(layer5_outputs(2609));
    layer6_outputs(4983) <= (layer5_outputs(2401)) xor (layer5_outputs(3397));
    layer6_outputs(4984) <= not(layer5_outputs(1238));
    layer6_outputs(4985) <= layer5_outputs(854);
    layer6_outputs(4986) <= (layer5_outputs(1359)) and not (layer5_outputs(2007));
    layer6_outputs(4987) <= not(layer5_outputs(2546));
    layer6_outputs(4988) <= layer5_outputs(1316);
    layer6_outputs(4989) <= not((layer5_outputs(2979)) and (layer5_outputs(2031)));
    layer6_outputs(4990) <= not(layer5_outputs(1018));
    layer6_outputs(4991) <= '1';
    layer6_outputs(4992) <= not((layer5_outputs(4251)) and (layer5_outputs(1742)));
    layer6_outputs(4993) <= not(layer5_outputs(431));
    layer6_outputs(4994) <= layer5_outputs(1935);
    layer6_outputs(4995) <= (layer5_outputs(4606)) and not (layer5_outputs(4755));
    layer6_outputs(4996) <= '0';
    layer6_outputs(4997) <= not((layer5_outputs(2582)) and (layer5_outputs(1956)));
    layer6_outputs(4998) <= layer5_outputs(4235);
    layer6_outputs(4999) <= layer5_outputs(4911);
    layer6_outputs(5000) <= not(layer5_outputs(3212));
    layer6_outputs(5001) <= (layer5_outputs(1876)) and not (layer5_outputs(2335));
    layer6_outputs(5002) <= not(layer5_outputs(409));
    layer6_outputs(5003) <= (layer5_outputs(352)) and (layer5_outputs(492));
    layer6_outputs(5004) <= (layer5_outputs(4944)) xor (layer5_outputs(4179));
    layer6_outputs(5005) <= layer5_outputs(1696);
    layer6_outputs(5006) <= not((layer5_outputs(1109)) and (layer5_outputs(4601)));
    layer6_outputs(5007) <= not((layer5_outputs(1972)) or (layer5_outputs(2202)));
    layer6_outputs(5008) <= layer5_outputs(564);
    layer6_outputs(5009) <= (layer5_outputs(4031)) or (layer5_outputs(156));
    layer6_outputs(5010) <= not(layer5_outputs(901));
    layer6_outputs(5011) <= (layer5_outputs(3219)) and not (layer5_outputs(4074));
    layer6_outputs(5012) <= layer5_outputs(4453);
    layer6_outputs(5013) <= not(layer5_outputs(3476));
    layer6_outputs(5014) <= not(layer5_outputs(2539));
    layer6_outputs(5015) <= not(layer5_outputs(4089));
    layer6_outputs(5016) <= layer5_outputs(3923);
    layer6_outputs(5017) <= not(layer5_outputs(3296)) or (layer5_outputs(4324));
    layer6_outputs(5018) <= not(layer5_outputs(3642));
    layer6_outputs(5019) <= layer5_outputs(2272);
    layer6_outputs(5020) <= not(layer5_outputs(2460)) or (layer5_outputs(4289));
    layer6_outputs(5021) <= layer5_outputs(802);
    layer6_outputs(5022) <= '0';
    layer6_outputs(5023) <= not((layer5_outputs(5039)) xor (layer5_outputs(36)));
    layer6_outputs(5024) <= not(layer5_outputs(4881));
    layer6_outputs(5025) <= not(layer5_outputs(4722));
    layer6_outputs(5026) <= layer5_outputs(69);
    layer6_outputs(5027) <= (layer5_outputs(1545)) xor (layer5_outputs(4068));
    layer6_outputs(5028) <= not(layer5_outputs(224));
    layer6_outputs(5029) <= (layer5_outputs(3243)) and (layer5_outputs(3644));
    layer6_outputs(5030) <= (layer5_outputs(1761)) or (layer5_outputs(730));
    layer6_outputs(5031) <= (layer5_outputs(1072)) xor (layer5_outputs(1474));
    layer6_outputs(5032) <= (layer5_outputs(2412)) or (layer5_outputs(817));
    layer6_outputs(5033) <= not((layer5_outputs(2942)) xor (layer5_outputs(1907)));
    layer6_outputs(5034) <= layer5_outputs(4640);
    layer6_outputs(5035) <= not(layer5_outputs(1809));
    layer6_outputs(5036) <= not((layer5_outputs(5050)) and (layer5_outputs(3683)));
    layer6_outputs(5037) <= not(layer5_outputs(355));
    layer6_outputs(5038) <= not(layer5_outputs(4114)) or (layer5_outputs(3006));
    layer6_outputs(5039) <= (layer5_outputs(1161)) and not (layer5_outputs(3076));
    layer6_outputs(5040) <= not((layer5_outputs(4738)) and (layer5_outputs(26)));
    layer6_outputs(5041) <= (layer5_outputs(1375)) or (layer5_outputs(1139));
    layer6_outputs(5042) <= not(layer5_outputs(3887));
    layer6_outputs(5043) <= (layer5_outputs(3827)) or (layer5_outputs(1985));
    layer6_outputs(5044) <= layer5_outputs(2962);
    layer6_outputs(5045) <= (layer5_outputs(3699)) and not (layer5_outputs(302));
    layer6_outputs(5046) <= not(layer5_outputs(3282)) or (layer5_outputs(2074));
    layer6_outputs(5047) <= layer5_outputs(998);
    layer6_outputs(5048) <= (layer5_outputs(1259)) and not (layer5_outputs(4519));
    layer6_outputs(5049) <= not(layer5_outputs(3339)) or (layer5_outputs(1987));
    layer6_outputs(5050) <= (layer5_outputs(3221)) xor (layer5_outputs(2435));
    layer6_outputs(5051) <= not(layer5_outputs(1304));
    layer6_outputs(5052) <= not((layer5_outputs(1664)) xor (layer5_outputs(1798)));
    layer6_outputs(5053) <= not((layer5_outputs(2878)) xor (layer5_outputs(4145)));
    layer6_outputs(5054) <= not(layer5_outputs(4191));
    layer6_outputs(5055) <= not(layer5_outputs(4540));
    layer6_outputs(5056) <= not(layer5_outputs(3684));
    layer6_outputs(5057) <= not(layer5_outputs(794));
    layer6_outputs(5058) <= layer5_outputs(617);
    layer6_outputs(5059) <= layer5_outputs(2166);
    layer6_outputs(5060) <= not(layer5_outputs(2420));
    layer6_outputs(5061) <= not(layer5_outputs(4610));
    layer6_outputs(5062) <= not(layer5_outputs(2518)) or (layer5_outputs(2800));
    layer6_outputs(5063) <= layer5_outputs(4645);
    layer6_outputs(5064) <= layer5_outputs(500);
    layer6_outputs(5065) <= layer5_outputs(1315);
    layer6_outputs(5066) <= (layer5_outputs(2058)) and (layer5_outputs(2485));
    layer6_outputs(5067) <= layer5_outputs(2818);
    layer6_outputs(5068) <= not(layer5_outputs(3919));
    layer6_outputs(5069) <= not(layer5_outputs(1978)) or (layer5_outputs(3977));
    layer6_outputs(5070) <= not((layer5_outputs(190)) and (layer5_outputs(1401)));
    layer6_outputs(5071) <= (layer5_outputs(2768)) xor (layer5_outputs(3998));
    layer6_outputs(5072) <= (layer5_outputs(2129)) and (layer5_outputs(137));
    layer6_outputs(5073) <= layer5_outputs(1633);
    layer6_outputs(5074) <= (layer5_outputs(3074)) or (layer5_outputs(2204));
    layer6_outputs(5075) <= layer5_outputs(3975);
    layer6_outputs(5076) <= layer5_outputs(2488);
    layer6_outputs(5077) <= '1';
    layer6_outputs(5078) <= not(layer5_outputs(1374));
    layer6_outputs(5079) <= not(layer5_outputs(2516));
    layer6_outputs(5080) <= not((layer5_outputs(1829)) or (layer5_outputs(4516)));
    layer6_outputs(5081) <= not((layer5_outputs(1145)) xor (layer5_outputs(975)));
    layer6_outputs(5082) <= not((layer5_outputs(4221)) and (layer5_outputs(4135)));
    layer6_outputs(5083) <= (layer5_outputs(4034)) xor (layer5_outputs(4530));
    layer6_outputs(5084) <= not(layer5_outputs(2659));
    layer6_outputs(5085) <= layer5_outputs(870);
    layer6_outputs(5086) <= '1';
    layer6_outputs(5087) <= not((layer5_outputs(783)) and (layer5_outputs(4570)));
    layer6_outputs(5088) <= not(layer5_outputs(2635));
    layer6_outputs(5089) <= layer5_outputs(2477);
    layer6_outputs(5090) <= (layer5_outputs(4641)) or (layer5_outputs(3372));
    layer6_outputs(5091) <= layer5_outputs(2292);
    layer6_outputs(5092) <= not(layer5_outputs(4685));
    layer6_outputs(5093) <= layer5_outputs(2265);
    layer6_outputs(5094) <= not((layer5_outputs(1057)) and (layer5_outputs(684)));
    layer6_outputs(5095) <= layer5_outputs(1991);
    layer6_outputs(5096) <= layer5_outputs(824);
    layer6_outputs(5097) <= not(layer5_outputs(3464)) or (layer5_outputs(4690));
    layer6_outputs(5098) <= (layer5_outputs(2018)) and not (layer5_outputs(3004));
    layer6_outputs(5099) <= layer5_outputs(39);
    layer6_outputs(5100) <= (layer5_outputs(2664)) xor (layer5_outputs(2181));
    layer6_outputs(5101) <= layer5_outputs(5096);
    layer6_outputs(5102) <= (layer5_outputs(3860)) and not (layer5_outputs(4967));
    layer6_outputs(5103) <= not(layer5_outputs(1849)) or (layer5_outputs(2042));
    layer6_outputs(5104) <= layer5_outputs(4743);
    layer6_outputs(5105) <= layer5_outputs(756);
    layer6_outputs(5106) <= layer5_outputs(4567);
    layer6_outputs(5107) <= not(layer5_outputs(768));
    layer6_outputs(5108) <= layer5_outputs(3459);
    layer6_outputs(5109) <= (layer5_outputs(3488)) and not (layer5_outputs(1909));
    layer6_outputs(5110) <= layer5_outputs(3610);
    layer6_outputs(5111) <= layer5_outputs(2057);
    layer6_outputs(5112) <= not((layer5_outputs(1016)) or (layer5_outputs(282)));
    layer6_outputs(5113) <= layer5_outputs(1785);
    layer6_outputs(5114) <= not((layer5_outputs(672)) or (layer5_outputs(451)));
    layer6_outputs(5115) <= not((layer5_outputs(3407)) or (layer5_outputs(1337)));
    layer6_outputs(5116) <= not(layer5_outputs(1242));
    layer6_outputs(5117) <= not(layer5_outputs(423));
    layer6_outputs(5118) <= layer5_outputs(2574);
    layer6_outputs(5119) <= not(layer5_outputs(4888)) or (layer5_outputs(1614));
    outputs(0) <= layer6_outputs(3511);
    outputs(1) <= not(layer6_outputs(3515));
    outputs(2) <= not(layer6_outputs(2080));
    outputs(3) <= layer6_outputs(1052);
    outputs(4) <= not((layer6_outputs(4166)) xor (layer6_outputs(2482)));
    outputs(5) <= layer6_outputs(1959);
    outputs(6) <= layer6_outputs(2283);
    outputs(7) <= layer6_outputs(2879);
    outputs(8) <= layer6_outputs(2048);
    outputs(9) <= layer6_outputs(1898);
    outputs(10) <= layer6_outputs(2642);
    outputs(11) <= layer6_outputs(4969);
    outputs(12) <= not(layer6_outputs(4848));
    outputs(13) <= not(layer6_outputs(3977));
    outputs(14) <= not(layer6_outputs(3646));
    outputs(15) <= layer6_outputs(5117);
    outputs(16) <= layer6_outputs(1120);
    outputs(17) <= layer6_outputs(1128);
    outputs(18) <= not((layer6_outputs(2326)) xor (layer6_outputs(1746)));
    outputs(19) <= not(layer6_outputs(1197));
    outputs(20) <= layer6_outputs(4433);
    outputs(21) <= not(layer6_outputs(1496));
    outputs(22) <= (layer6_outputs(5062)) and (layer6_outputs(739));
    outputs(23) <= layer6_outputs(4502);
    outputs(24) <= not(layer6_outputs(1148));
    outputs(25) <= not(layer6_outputs(1928)) or (layer6_outputs(3762));
    outputs(26) <= not(layer6_outputs(896));
    outputs(27) <= layer6_outputs(1679);
    outputs(28) <= not((layer6_outputs(1943)) xor (layer6_outputs(2895)));
    outputs(29) <= not(layer6_outputs(260));
    outputs(30) <= not((layer6_outputs(5078)) xor (layer6_outputs(2078)));
    outputs(31) <= layer6_outputs(3766);
    outputs(32) <= not((layer6_outputs(4600)) and (layer6_outputs(2771)));
    outputs(33) <= (layer6_outputs(3212)) xor (layer6_outputs(2328));
    outputs(34) <= not((layer6_outputs(3635)) xor (layer6_outputs(1046)));
    outputs(35) <= (layer6_outputs(4216)) and not (layer6_outputs(644));
    outputs(36) <= layer6_outputs(423);
    outputs(37) <= not((layer6_outputs(2939)) or (layer6_outputs(3646)));
    outputs(38) <= (layer6_outputs(3254)) xor (layer6_outputs(2436));
    outputs(39) <= not(layer6_outputs(4858));
    outputs(40) <= not(layer6_outputs(3524));
    outputs(41) <= (layer6_outputs(285)) xor (layer6_outputs(2856));
    outputs(42) <= (layer6_outputs(672)) or (layer6_outputs(1194));
    outputs(43) <= not(layer6_outputs(3411));
    outputs(44) <= not(layer6_outputs(4916));
    outputs(45) <= not(layer6_outputs(1584));
    outputs(46) <= layer6_outputs(1918);
    outputs(47) <= layer6_outputs(1429);
    outputs(48) <= not((layer6_outputs(2539)) xor (layer6_outputs(577)));
    outputs(49) <= not(layer6_outputs(293));
    outputs(50) <= not((layer6_outputs(387)) or (layer6_outputs(5060)));
    outputs(51) <= not(layer6_outputs(3591));
    outputs(52) <= not(layer6_outputs(4017));
    outputs(53) <= layer6_outputs(947);
    outputs(54) <= not(layer6_outputs(524));
    outputs(55) <= not((layer6_outputs(1436)) or (layer6_outputs(2730)));
    outputs(56) <= layer6_outputs(3452);
    outputs(57) <= layer6_outputs(1552);
    outputs(58) <= not(layer6_outputs(3317));
    outputs(59) <= not(layer6_outputs(1054));
    outputs(60) <= not((layer6_outputs(2990)) or (layer6_outputs(2309)));
    outputs(61) <= not(layer6_outputs(3571));
    outputs(62) <= layer6_outputs(726);
    outputs(63) <= (layer6_outputs(4044)) xor (layer6_outputs(602));
    outputs(64) <= layer6_outputs(3587);
    outputs(65) <= (layer6_outputs(59)) xor (layer6_outputs(133));
    outputs(66) <= layer6_outputs(1576);
    outputs(67) <= not(layer6_outputs(252));
    outputs(68) <= layer6_outputs(3495);
    outputs(69) <= not(layer6_outputs(4676));
    outputs(70) <= not(layer6_outputs(1438));
    outputs(71) <= not((layer6_outputs(2803)) xor (layer6_outputs(3315)));
    outputs(72) <= not(layer6_outputs(3450));
    outputs(73) <= not(layer6_outputs(4641));
    outputs(74) <= layer6_outputs(4971);
    outputs(75) <= layer6_outputs(3007);
    outputs(76) <= layer6_outputs(4150);
    outputs(77) <= layer6_outputs(4416);
    outputs(78) <= not(layer6_outputs(641));
    outputs(79) <= layer6_outputs(5093);
    outputs(80) <= not(layer6_outputs(4144));
    outputs(81) <= not(layer6_outputs(2963));
    outputs(82) <= not((layer6_outputs(4552)) xor (layer6_outputs(1674)));
    outputs(83) <= not(layer6_outputs(4336));
    outputs(84) <= (layer6_outputs(3868)) xor (layer6_outputs(324));
    outputs(85) <= layer6_outputs(4571);
    outputs(86) <= layer6_outputs(1359);
    outputs(87) <= not(layer6_outputs(1518));
    outputs(88) <= layer6_outputs(4140);
    outputs(89) <= layer6_outputs(4139);
    outputs(90) <= not(layer6_outputs(2236));
    outputs(91) <= not((layer6_outputs(4857)) xor (layer6_outputs(4333)));
    outputs(92) <= not((layer6_outputs(3754)) and (layer6_outputs(1187)));
    outputs(93) <= layer6_outputs(1221);
    outputs(94) <= layer6_outputs(4294);
    outputs(95) <= not(layer6_outputs(3155));
    outputs(96) <= not((layer6_outputs(1354)) xor (layer6_outputs(974)));
    outputs(97) <= not(layer6_outputs(3861));
    outputs(98) <= layer6_outputs(325);
    outputs(99) <= not(layer6_outputs(817));
    outputs(100) <= not((layer6_outputs(2560)) and (layer6_outputs(1381)));
    outputs(101) <= not((layer6_outputs(2920)) xor (layer6_outputs(4846)));
    outputs(102) <= layer6_outputs(2319);
    outputs(103) <= not(layer6_outputs(4296));
    outputs(104) <= layer6_outputs(3432);
    outputs(105) <= (layer6_outputs(3816)) and (layer6_outputs(3201));
    outputs(106) <= layer6_outputs(4895);
    outputs(107) <= not(layer6_outputs(1495));
    outputs(108) <= layer6_outputs(2878);
    outputs(109) <= not(layer6_outputs(630));
    outputs(110) <= not((layer6_outputs(2639)) xor (layer6_outputs(4620)));
    outputs(111) <= layer6_outputs(3808);
    outputs(112) <= (layer6_outputs(664)) and not (layer6_outputs(4620));
    outputs(113) <= not(layer6_outputs(239));
    outputs(114) <= not(layer6_outputs(1448));
    outputs(115) <= (layer6_outputs(2016)) xor (layer6_outputs(4055));
    outputs(116) <= layer6_outputs(1940);
    outputs(117) <= (layer6_outputs(4888)) and not (layer6_outputs(1665));
    outputs(118) <= not(layer6_outputs(443)) or (layer6_outputs(567));
    outputs(119) <= not(layer6_outputs(1331)) or (layer6_outputs(2421));
    outputs(120) <= not(layer6_outputs(3723));
    outputs(121) <= not(layer6_outputs(1300));
    outputs(122) <= layer6_outputs(4190);
    outputs(123) <= layer6_outputs(3626);
    outputs(124) <= not(layer6_outputs(89));
    outputs(125) <= not(layer6_outputs(3827));
    outputs(126) <= layer6_outputs(2881);
    outputs(127) <= (layer6_outputs(3546)) xor (layer6_outputs(557));
    outputs(128) <= not((layer6_outputs(4010)) or (layer6_outputs(2059)));
    outputs(129) <= (layer6_outputs(1807)) xor (layer6_outputs(4557));
    outputs(130) <= (layer6_outputs(2474)) xor (layer6_outputs(364));
    outputs(131) <= (layer6_outputs(2613)) and not (layer6_outputs(4094));
    outputs(132) <= (layer6_outputs(4759)) xor (layer6_outputs(264));
    outputs(133) <= layer6_outputs(1701);
    outputs(134) <= not(layer6_outputs(78));
    outputs(135) <= not(layer6_outputs(4869));
    outputs(136) <= layer6_outputs(360);
    outputs(137) <= not((layer6_outputs(4455)) xor (layer6_outputs(4035)));
    outputs(138) <= layer6_outputs(2844);
    outputs(139) <= (layer6_outputs(2026)) or (layer6_outputs(811));
    outputs(140) <= layer6_outputs(1526);
    outputs(141) <= not((layer6_outputs(2995)) xor (layer6_outputs(4843)));
    outputs(142) <= (layer6_outputs(3359)) or (layer6_outputs(686));
    outputs(143) <= layer6_outputs(1090);
    outputs(144) <= not(layer6_outputs(4804));
    outputs(145) <= (layer6_outputs(1560)) xor (layer6_outputs(821));
    outputs(146) <= not(layer6_outputs(4842));
    outputs(147) <= not(layer6_outputs(4030));
    outputs(148) <= (layer6_outputs(241)) xor (layer6_outputs(4768));
    outputs(149) <= layer6_outputs(130);
    outputs(150) <= layer6_outputs(7);
    outputs(151) <= not(layer6_outputs(2787));
    outputs(152) <= not(layer6_outputs(3349));
    outputs(153) <= layer6_outputs(3406);
    outputs(154) <= not(layer6_outputs(946));
    outputs(155) <= (layer6_outputs(3)) xor (layer6_outputs(1067));
    outputs(156) <= not(layer6_outputs(4037));
    outputs(157) <= not(layer6_outputs(4858));
    outputs(158) <= layer6_outputs(1748);
    outputs(159) <= (layer6_outputs(1447)) and (layer6_outputs(2914));
    outputs(160) <= layer6_outputs(2633);
    outputs(161) <= not(layer6_outputs(1931));
    outputs(162) <= (layer6_outputs(2157)) xor (layer6_outputs(1013));
    outputs(163) <= layer6_outputs(4323);
    outputs(164) <= not((layer6_outputs(1397)) or (layer6_outputs(4319)));
    outputs(165) <= not(layer6_outputs(168));
    outputs(166) <= not((layer6_outputs(1866)) xor (layer6_outputs(2299)));
    outputs(167) <= not((layer6_outputs(4997)) xor (layer6_outputs(895)));
    outputs(168) <= (layer6_outputs(49)) and not (layer6_outputs(1548));
    outputs(169) <= not((layer6_outputs(3796)) or (layer6_outputs(998)));
    outputs(170) <= layer6_outputs(3053);
    outputs(171) <= not(layer6_outputs(4131));
    outputs(172) <= layer6_outputs(3550);
    outputs(173) <= (layer6_outputs(3244)) xor (layer6_outputs(1691));
    outputs(174) <= not(layer6_outputs(4573));
    outputs(175) <= not((layer6_outputs(246)) or (layer6_outputs(515)));
    outputs(176) <= (layer6_outputs(4974)) xor (layer6_outputs(218));
    outputs(177) <= not(layer6_outputs(1068));
    outputs(178) <= layer6_outputs(1317);
    outputs(179) <= (layer6_outputs(4932)) xor (layer6_outputs(539));
    outputs(180) <= layer6_outputs(1926);
    outputs(181) <= not(layer6_outputs(5013));
    outputs(182) <= not((layer6_outputs(4899)) and (layer6_outputs(4802)));
    outputs(183) <= layer6_outputs(4849);
    outputs(184) <= (layer6_outputs(5021)) xor (layer6_outputs(1143));
    outputs(185) <= layer6_outputs(1170);
    outputs(186) <= layer6_outputs(4418);
    outputs(187) <= not((layer6_outputs(700)) and (layer6_outputs(4845)));
    outputs(188) <= not((layer6_outputs(2705)) and (layer6_outputs(3583)));
    outputs(189) <= not(layer6_outputs(1643));
    outputs(190) <= not(layer6_outputs(2060));
    outputs(191) <= not(layer6_outputs(4279));
    outputs(192) <= not(layer6_outputs(1198));
    outputs(193) <= not((layer6_outputs(839)) xor (layer6_outputs(178)));
    outputs(194) <= not(layer6_outputs(2676));
    outputs(195) <= not(layer6_outputs(966));
    outputs(196) <= not(layer6_outputs(4310));
    outputs(197) <= layer6_outputs(1814);
    outputs(198) <= layer6_outputs(4743);
    outputs(199) <= layer6_outputs(5101);
    outputs(200) <= not(layer6_outputs(2992));
    outputs(201) <= not(layer6_outputs(4496));
    outputs(202) <= (layer6_outputs(4159)) xor (layer6_outputs(1116));
    outputs(203) <= not(layer6_outputs(1970));
    outputs(204) <= layer6_outputs(5042);
    outputs(205) <= (layer6_outputs(3681)) xor (layer6_outputs(1125));
    outputs(206) <= not((layer6_outputs(3440)) xor (layer6_outputs(3737)));
    outputs(207) <= not(layer6_outputs(3957));
    outputs(208) <= not((layer6_outputs(3760)) xor (layer6_outputs(984)));
    outputs(209) <= not(layer6_outputs(3351));
    outputs(210) <= layer6_outputs(1468);
    outputs(211) <= not((layer6_outputs(642)) or (layer6_outputs(1362)));
    outputs(212) <= not((layer6_outputs(5048)) or (layer6_outputs(4490)));
    outputs(213) <= not(layer6_outputs(2541));
    outputs(214) <= not(layer6_outputs(2248));
    outputs(215) <= not((layer6_outputs(855)) and (layer6_outputs(3719)));
    outputs(216) <= (layer6_outputs(2123)) and not (layer6_outputs(357));
    outputs(217) <= layer6_outputs(2532);
    outputs(218) <= layer6_outputs(2023);
    outputs(219) <= layer6_outputs(2643);
    outputs(220) <= not(layer6_outputs(3945));
    outputs(221) <= (layer6_outputs(215)) xor (layer6_outputs(1602));
    outputs(222) <= not((layer6_outputs(2588)) xor (layer6_outputs(1543)));
    outputs(223) <= not(layer6_outputs(85));
    outputs(224) <= layer6_outputs(590);
    outputs(225) <= layer6_outputs(1177);
    outputs(226) <= not(layer6_outputs(1484));
    outputs(227) <= not((layer6_outputs(3399)) xor (layer6_outputs(78)));
    outputs(228) <= not(layer6_outputs(1637));
    outputs(229) <= layer6_outputs(1128);
    outputs(230) <= layer6_outputs(144);
    outputs(231) <= not(layer6_outputs(1752));
    outputs(232) <= not(layer6_outputs(4894));
    outputs(233) <= (layer6_outputs(1676)) xor (layer6_outputs(2361));
    outputs(234) <= not(layer6_outputs(3494));
    outputs(235) <= layer6_outputs(4785);
    outputs(236) <= not(layer6_outputs(2902));
    outputs(237) <= not(layer6_outputs(3633));
    outputs(238) <= layer6_outputs(3843);
    outputs(239) <= not(layer6_outputs(4096));
    outputs(240) <= not(layer6_outputs(2030));
    outputs(241) <= not(layer6_outputs(4475));
    outputs(242) <= not(layer6_outputs(1206));
    outputs(243) <= (layer6_outputs(1631)) and not (layer6_outputs(2994));
    outputs(244) <= layer6_outputs(2082);
    outputs(245) <= (layer6_outputs(2564)) xor (layer6_outputs(893));
    outputs(246) <= layer6_outputs(3617);
    outputs(247) <= layer6_outputs(4184);
    outputs(248) <= layer6_outputs(51);
    outputs(249) <= layer6_outputs(256);
    outputs(250) <= not(layer6_outputs(4917));
    outputs(251) <= (layer6_outputs(1465)) xor (layer6_outputs(1842));
    outputs(252) <= not(layer6_outputs(3360));
    outputs(253) <= not(layer6_outputs(3936));
    outputs(254) <= (layer6_outputs(879)) and not (layer6_outputs(2688));
    outputs(255) <= not((layer6_outputs(4192)) xor (layer6_outputs(2085)));
    outputs(256) <= not(layer6_outputs(315));
    outputs(257) <= not(layer6_outputs(682));
    outputs(258) <= layer6_outputs(3862);
    outputs(259) <= not((layer6_outputs(2798)) xor (layer6_outputs(1304)));
    outputs(260) <= not(layer6_outputs(2575));
    outputs(261) <= not(layer6_outputs(1352));
    outputs(262) <= not((layer6_outputs(4893)) and (layer6_outputs(4373)));
    outputs(263) <= layer6_outputs(2965);
    outputs(264) <= not(layer6_outputs(4963));
    outputs(265) <= (layer6_outputs(3994)) xor (layer6_outputs(4661));
    outputs(266) <= not(layer6_outputs(2597));
    outputs(267) <= layer6_outputs(1356);
    outputs(268) <= not((layer6_outputs(628)) xor (layer6_outputs(765)));
    outputs(269) <= layer6_outputs(18);
    outputs(270) <= not(layer6_outputs(1098));
    outputs(271) <= (layer6_outputs(3037)) xor (layer6_outputs(1104));
    outputs(272) <= (layer6_outputs(214)) and not (layer6_outputs(4338));
    outputs(273) <= not((layer6_outputs(4381)) xor (layer6_outputs(439)));
    outputs(274) <= layer6_outputs(2874);
    outputs(275) <= not(layer6_outputs(1745));
    outputs(276) <= not(layer6_outputs(2128));
    outputs(277) <= not((layer6_outputs(4385)) or (layer6_outputs(2201)));
    outputs(278) <= not(layer6_outputs(3252));
    outputs(279) <= layer6_outputs(299);
    outputs(280) <= not(layer6_outputs(4833));
    outputs(281) <= not(layer6_outputs(1558));
    outputs(282) <= (layer6_outputs(2340)) and (layer6_outputs(498));
    outputs(283) <= not((layer6_outputs(1247)) xor (layer6_outputs(5055)));
    outputs(284) <= layer6_outputs(1309);
    outputs(285) <= layer6_outputs(1896);
    outputs(286) <= not(layer6_outputs(1886));
    outputs(287) <= layer6_outputs(2450);
    outputs(288) <= (layer6_outputs(172)) xor (layer6_outputs(1060));
    outputs(289) <= layer6_outputs(1167);
    outputs(290) <= layer6_outputs(41);
    outputs(291) <= not((layer6_outputs(1971)) xor (layer6_outputs(2523)));
    outputs(292) <= not((layer6_outputs(3600)) and (layer6_outputs(2849)));
    outputs(293) <= not((layer6_outputs(2737)) xor (layer6_outputs(4704)));
    outputs(294) <= not(layer6_outputs(4689));
    outputs(295) <= not(layer6_outputs(210));
    outputs(296) <= layer6_outputs(592);
    outputs(297) <= (layer6_outputs(3801)) and (layer6_outputs(433));
    outputs(298) <= (layer6_outputs(949)) or (layer6_outputs(4062));
    outputs(299) <= not(layer6_outputs(4867)) or (layer6_outputs(3106));
    outputs(300) <= layer6_outputs(3597);
    outputs(301) <= (layer6_outputs(985)) xor (layer6_outputs(68));
    outputs(302) <= layer6_outputs(2813);
    outputs(303) <= not((layer6_outputs(2704)) xor (layer6_outputs(1600)));
    outputs(304) <= (layer6_outputs(29)) and not (layer6_outputs(2189));
    outputs(305) <= (layer6_outputs(4662)) and not (layer6_outputs(4816));
    outputs(306) <= layer6_outputs(4126);
    outputs(307) <= not(layer6_outputs(595));
    outputs(308) <= layer6_outputs(3325);
    outputs(309) <= not(layer6_outputs(2999));
    outputs(310) <= layer6_outputs(199);
    outputs(311) <= not(layer6_outputs(1707));
    outputs(312) <= layer6_outputs(952);
    outputs(313) <= not(layer6_outputs(220)) or (layer6_outputs(4301));
    outputs(314) <= (layer6_outputs(3817)) and not (layer6_outputs(4641));
    outputs(315) <= not(layer6_outputs(1786));
    outputs(316) <= (layer6_outputs(2153)) xor (layer6_outputs(4549));
    outputs(317) <= not(layer6_outputs(868));
    outputs(318) <= layer6_outputs(444);
    outputs(319) <= layer6_outputs(4442);
    outputs(320) <= layer6_outputs(3983);
    outputs(321) <= not((layer6_outputs(4410)) xor (layer6_outputs(4997)));
    outputs(322) <= not((layer6_outputs(4520)) xor (layer6_outputs(3740)));
    outputs(323) <= (layer6_outputs(1929)) xor (layer6_outputs(5008));
    outputs(324) <= not(layer6_outputs(511));
    outputs(325) <= layer6_outputs(714);
    outputs(326) <= not(layer6_outputs(141));
    outputs(327) <= (layer6_outputs(3711)) or (layer6_outputs(3787));
    outputs(328) <= not(layer6_outputs(3973));
    outputs(329) <= layer6_outputs(4700);
    outputs(330) <= not(layer6_outputs(1463));
    outputs(331) <= layer6_outputs(3829);
    outputs(332) <= not(layer6_outputs(4228));
    outputs(333) <= not(layer6_outputs(4817));
    outputs(334) <= (layer6_outputs(4358)) xor (layer6_outputs(1492));
    outputs(335) <= (layer6_outputs(3129)) and (layer6_outputs(4074));
    outputs(336) <= layer6_outputs(2587);
    outputs(337) <= layer6_outputs(3290);
    outputs(338) <= layer6_outputs(3582);
    outputs(339) <= not(layer6_outputs(2697));
    outputs(340) <= layer6_outputs(3589);
    outputs(341) <= not(layer6_outputs(4341));
    outputs(342) <= layer6_outputs(2390);
    outputs(343) <= not(layer6_outputs(2684));
    outputs(344) <= layer6_outputs(738);
    outputs(345) <= layer6_outputs(4669);
    outputs(346) <= layer6_outputs(1685);
    outputs(347) <= not(layer6_outputs(690));
    outputs(348) <= layer6_outputs(746);
    outputs(349) <= not(layer6_outputs(4451));
    outputs(350) <= not(layer6_outputs(4107)) or (layer6_outputs(283));
    outputs(351) <= not(layer6_outputs(284)) or (layer6_outputs(4203));
    outputs(352) <= (layer6_outputs(5072)) xor (layer6_outputs(2977));
    outputs(353) <= layer6_outputs(4944);
    outputs(354) <= layer6_outputs(2084);
    outputs(355) <= (layer6_outputs(177)) and not (layer6_outputs(1434));
    outputs(356) <= not(layer6_outputs(3572));
    outputs(357) <= not(layer6_outputs(2529));
    outputs(358) <= not((layer6_outputs(4622)) or (layer6_outputs(1710)));
    outputs(359) <= not(layer6_outputs(3082)) or (layer6_outputs(4486));
    outputs(360) <= layer6_outputs(843);
    outputs(361) <= (layer6_outputs(3736)) xor (layer6_outputs(2912));
    outputs(362) <= layer6_outputs(4090);
    outputs(363) <= not(layer6_outputs(2343));
    outputs(364) <= layer6_outputs(2166);
    outputs(365) <= layer6_outputs(1390);
    outputs(366) <= not((layer6_outputs(1020)) xor (layer6_outputs(2586)));
    outputs(367) <= not((layer6_outputs(3678)) xor (layer6_outputs(1417)));
    outputs(368) <= not(layer6_outputs(266));
    outputs(369) <= layer6_outputs(4482);
    outputs(370) <= layer6_outputs(3819);
    outputs(371) <= layer6_outputs(4696);
    outputs(372) <= not((layer6_outputs(4272)) xor (layer6_outputs(4316)));
    outputs(373) <= layer6_outputs(2530);
    outputs(374) <= layer6_outputs(120);
    outputs(375) <= layer6_outputs(1819);
    outputs(376) <= layer6_outputs(564);
    outputs(377) <= layer6_outputs(1601);
    outputs(378) <= not(layer6_outputs(649));
    outputs(379) <= layer6_outputs(4518);
    outputs(380) <= not((layer6_outputs(2985)) xor (layer6_outputs(2636)));
    outputs(381) <= not(layer6_outputs(573));
    outputs(382) <= not(layer6_outputs(4815));
    outputs(383) <= not((layer6_outputs(2122)) xor (layer6_outputs(3208)));
    outputs(384) <= (layer6_outputs(1533)) xor (layer6_outputs(1324));
    outputs(385) <= not(layer6_outputs(317));
    outputs(386) <= not(layer6_outputs(2250));
    outputs(387) <= not(layer6_outputs(1203));
    outputs(388) <= layer6_outputs(4729);
    outputs(389) <= not((layer6_outputs(802)) xor (layer6_outputs(715)));
    outputs(390) <= (layer6_outputs(3194)) xor (layer6_outputs(4632));
    outputs(391) <= not((layer6_outputs(2600)) xor (layer6_outputs(2397)));
    outputs(392) <= not(layer6_outputs(2121));
    outputs(393) <= not(layer6_outputs(1993));
    outputs(394) <= not(layer6_outputs(2837));
    outputs(395) <= not(layer6_outputs(1594)) or (layer6_outputs(2184));
    outputs(396) <= not(layer6_outputs(5050));
    outputs(397) <= not(layer6_outputs(1470));
    outputs(398) <= layer6_outputs(3543);
    outputs(399) <= (layer6_outputs(3421)) and (layer6_outputs(3314));
    outputs(400) <= not(layer6_outputs(4100));
    outputs(401) <= not((layer6_outputs(2257)) or (layer6_outputs(5084)));
    outputs(402) <= (layer6_outputs(1153)) xor (layer6_outputs(4432));
    outputs(403) <= layer6_outputs(1859);
    outputs(404) <= (layer6_outputs(829)) and not (layer6_outputs(903));
    outputs(405) <= (layer6_outputs(1761)) xor (layer6_outputs(5081));
    outputs(406) <= layer6_outputs(1446);
    outputs(407) <= layer6_outputs(4970);
    outputs(408) <= not((layer6_outputs(3476)) and (layer6_outputs(4465)));
    outputs(409) <= not(layer6_outputs(1572));
    outputs(410) <= (layer6_outputs(2286)) or (layer6_outputs(4538));
    outputs(411) <= layer6_outputs(4294);
    outputs(412) <= (layer6_outputs(2030)) xor (layer6_outputs(598));
    outputs(413) <= layer6_outputs(1959);
    outputs(414) <= (layer6_outputs(63)) xor (layer6_outputs(2945));
    outputs(415) <= not((layer6_outputs(3153)) xor (layer6_outputs(1550)));
    outputs(416) <= not(layer6_outputs(3929));
    outputs(417) <= not(layer6_outputs(776));
    outputs(418) <= not(layer6_outputs(1551));
    outputs(419) <= not((layer6_outputs(2823)) xor (layer6_outputs(5021)));
    outputs(420) <= not((layer6_outputs(4892)) xor (layer6_outputs(1094)));
    outputs(421) <= not(layer6_outputs(1508));
    outputs(422) <= not(layer6_outputs(915)) or (layer6_outputs(4522));
    outputs(423) <= (layer6_outputs(3236)) xor (layer6_outputs(394));
    outputs(424) <= not(layer6_outputs(3441));
    outputs(425) <= not(layer6_outputs(561));
    outputs(426) <= not(layer6_outputs(2725));
    outputs(427) <= not((layer6_outputs(2183)) or (layer6_outputs(2236)));
    outputs(428) <= (layer6_outputs(3459)) and (layer6_outputs(112));
    outputs(429) <= not(layer6_outputs(2663));
    outputs(430) <= not(layer6_outputs(2712));
    outputs(431) <= not(layer6_outputs(4355));
    outputs(432) <= layer6_outputs(4666);
    outputs(433) <= (layer6_outputs(4012)) xor (layer6_outputs(5074));
    outputs(434) <= layer6_outputs(1962);
    outputs(435) <= (layer6_outputs(2631)) and not (layer6_outputs(2403));
    outputs(436) <= not(layer6_outputs(2147));
    outputs(437) <= not((layer6_outputs(393)) or (layer6_outputs(4824)));
    outputs(438) <= not((layer6_outputs(1536)) xor (layer6_outputs(938)));
    outputs(439) <= (layer6_outputs(2455)) and (layer6_outputs(1552));
    outputs(440) <= not((layer6_outputs(3792)) or (layer6_outputs(2293)));
    outputs(441) <= (layer6_outputs(2978)) or (layer6_outputs(3149));
    outputs(442) <= not(layer6_outputs(2867));
    outputs(443) <= (layer6_outputs(719)) xor (layer6_outputs(2572));
    outputs(444) <= layer6_outputs(290);
    outputs(445) <= not(layer6_outputs(4650));
    outputs(446) <= (layer6_outputs(4820)) xor (layer6_outputs(1919));
    outputs(447) <= layer6_outputs(4403);
    outputs(448) <= layer6_outputs(2151);
    outputs(449) <= layer6_outputs(3234);
    outputs(450) <= not(layer6_outputs(916));
    outputs(451) <= (layer6_outputs(2271)) or (layer6_outputs(3557));
    outputs(452) <= not(layer6_outputs(1240));
    outputs(453) <= not(layer6_outputs(2107));
    outputs(454) <= layer6_outputs(2378);
    outputs(455) <= layer6_outputs(461);
    outputs(456) <= not(layer6_outputs(581));
    outputs(457) <= layer6_outputs(3573);
    outputs(458) <= not((layer6_outputs(3454)) xor (layer6_outputs(3309)));
    outputs(459) <= not(layer6_outputs(3109));
    outputs(460) <= layer6_outputs(1133);
    outputs(461) <= layer6_outputs(3581);
    outputs(462) <= not(layer6_outputs(3688));
    outputs(463) <= layer6_outputs(4325);
    outputs(464) <= layer6_outputs(4599);
    outputs(465) <= not(layer6_outputs(3898));
    outputs(466) <= layer6_outputs(3705);
    outputs(467) <= not((layer6_outputs(2801)) xor (layer6_outputs(384)));
    outputs(468) <= not((layer6_outputs(2649)) or (layer6_outputs(3539)));
    outputs(469) <= not(layer6_outputs(3788));
    outputs(470) <= not((layer6_outputs(3276)) xor (layer6_outputs(3762)));
    outputs(471) <= layer6_outputs(51);
    outputs(472) <= layer6_outputs(4087);
    outputs(473) <= not(layer6_outputs(3279));
    outputs(474) <= layer6_outputs(2651);
    outputs(475) <= not(layer6_outputs(4122));
    outputs(476) <= not(layer6_outputs(3951));
    outputs(477) <= layer6_outputs(1956);
    outputs(478) <= layer6_outputs(1560);
    outputs(479) <= (layer6_outputs(2474)) xor (layer6_outputs(458));
    outputs(480) <= layer6_outputs(98);
    outputs(481) <= (layer6_outputs(925)) xor (layer6_outputs(1154));
    outputs(482) <= layer6_outputs(421);
    outputs(483) <= layer6_outputs(4479);
    outputs(484) <= layer6_outputs(3448);
    outputs(485) <= layer6_outputs(2898);
    outputs(486) <= layer6_outputs(353);
    outputs(487) <= not(layer6_outputs(3701));
    outputs(488) <= layer6_outputs(2282);
    outputs(489) <= (layer6_outputs(4034)) or (layer6_outputs(1888));
    outputs(490) <= not(layer6_outputs(552));
    outputs(491) <= (layer6_outputs(3250)) xor (layer6_outputs(1899));
    outputs(492) <= layer6_outputs(1732);
    outputs(493) <= layer6_outputs(5089);
    outputs(494) <= not(layer6_outputs(4717)) or (layer6_outputs(4582));
    outputs(495) <= not(layer6_outputs(3072));
    outputs(496) <= not((layer6_outputs(4237)) xor (layer6_outputs(1746)));
    outputs(497) <= not(layer6_outputs(4804));
    outputs(498) <= not(layer6_outputs(3001));
    outputs(499) <= not((layer6_outputs(1050)) xor (layer6_outputs(3919)));
    outputs(500) <= not((layer6_outputs(1766)) or (layer6_outputs(4524)));
    outputs(501) <= layer6_outputs(389);
    outputs(502) <= not((layer6_outputs(587)) xor (layer6_outputs(4232)));
    outputs(503) <= not(layer6_outputs(4904));
    outputs(504) <= layer6_outputs(3045);
    outputs(505) <= not(layer6_outputs(1696));
    outputs(506) <= not(layer6_outputs(2517));
    outputs(507) <= not(layer6_outputs(4222));
    outputs(508) <= (layer6_outputs(191)) and not (layer6_outputs(3200));
    outputs(509) <= not((layer6_outputs(1242)) or (layer6_outputs(3917)));
    outputs(510) <= (layer6_outputs(3266)) xor (layer6_outputs(499));
    outputs(511) <= not(layer6_outputs(931));
    outputs(512) <= layer6_outputs(2581);
    outputs(513) <= layer6_outputs(907);
    outputs(514) <= not(layer6_outputs(1207));
    outputs(515) <= not((layer6_outputs(1510)) xor (layer6_outputs(4762)));
    outputs(516) <= not(layer6_outputs(1716)) or (layer6_outputs(742));
    outputs(517) <= not((layer6_outputs(62)) or (layer6_outputs(1535)));
    outputs(518) <= (layer6_outputs(2725)) and not (layer6_outputs(513));
    outputs(519) <= layer6_outputs(2702);
    outputs(520) <= layer6_outputs(2652);
    outputs(521) <= not(layer6_outputs(4132));
    outputs(522) <= layer6_outputs(2683);
    outputs(523) <= layer6_outputs(1299);
    outputs(524) <= not((layer6_outputs(3433)) or (layer6_outputs(1579)));
    outputs(525) <= not(layer6_outputs(4074));
    outputs(526) <= not(layer6_outputs(361));
    outputs(527) <= (layer6_outputs(3868)) and not (layer6_outputs(2097));
    outputs(528) <= not(layer6_outputs(4861));
    outputs(529) <= (layer6_outputs(4989)) xor (layer6_outputs(4467));
    outputs(530) <= not(layer6_outputs(1905));
    outputs(531) <= (layer6_outputs(1174)) and (layer6_outputs(545));
    outputs(532) <= not(layer6_outputs(2799));
    outputs(533) <= layer6_outputs(3094);
    outputs(534) <= not(layer6_outputs(4118));
    outputs(535) <= layer6_outputs(294);
    outputs(536) <= not(layer6_outputs(4042));
    outputs(537) <= layer6_outputs(518);
    outputs(538) <= layer6_outputs(2755);
    outputs(539) <= (layer6_outputs(4777)) xor (layer6_outputs(3836));
    outputs(540) <= not((layer6_outputs(2002)) or (layer6_outputs(4382)));
    outputs(541) <= not((layer6_outputs(68)) or (layer6_outputs(1855)));
    outputs(542) <= not(layer6_outputs(3083));
    outputs(543) <= (layer6_outputs(4023)) and not (layer6_outputs(4121));
    outputs(544) <= not(layer6_outputs(2692));
    outputs(545) <= not((layer6_outputs(2630)) xor (layer6_outputs(4567)));
    outputs(546) <= not(layer6_outputs(2930));
    outputs(547) <= not((layer6_outputs(3330)) and (layer6_outputs(4103)));
    outputs(548) <= not(layer6_outputs(2386));
    outputs(549) <= layer6_outputs(4592);
    outputs(550) <= layer6_outputs(1340);
    outputs(551) <= layer6_outputs(1230);
    outputs(552) <= layer6_outputs(713);
    outputs(553) <= not(layer6_outputs(1165));
    outputs(554) <= not(layer6_outputs(35));
    outputs(555) <= layer6_outputs(4154);
    outputs(556) <= layer6_outputs(70);
    outputs(557) <= layer6_outputs(1497);
    outputs(558) <= layer6_outputs(4431);
    outputs(559) <= (layer6_outputs(4316)) or (layer6_outputs(4768));
    outputs(560) <= layer6_outputs(3908);
    outputs(561) <= not(layer6_outputs(2081));
    outputs(562) <= not(layer6_outputs(1658));
    outputs(563) <= layer6_outputs(606);
    outputs(564) <= (layer6_outputs(846)) xor (layer6_outputs(2602));
    outputs(565) <= not(layer6_outputs(4775));
    outputs(566) <= (layer6_outputs(1302)) and (layer6_outputs(782));
    outputs(567) <= (layer6_outputs(3980)) and not (layer6_outputs(1861));
    outputs(568) <= layer6_outputs(219);
    outputs(569) <= not(layer6_outputs(1818));
    outputs(570) <= (layer6_outputs(4698)) and (layer6_outputs(1512));
    outputs(571) <= (layer6_outputs(3926)) and not (layer6_outputs(1545));
    outputs(572) <= layer6_outputs(9);
    outputs(573) <= layer6_outputs(1071);
    outputs(574) <= not(layer6_outputs(1041));
    outputs(575) <= not(layer6_outputs(3359));
    outputs(576) <= layer6_outputs(304);
    outputs(577) <= (layer6_outputs(932)) and (layer6_outputs(4344));
    outputs(578) <= not(layer6_outputs(1275));
    outputs(579) <= not(layer6_outputs(3783));
    outputs(580) <= not(layer6_outputs(2713));
    outputs(581) <= not(layer6_outputs(1675));
    outputs(582) <= not(layer6_outputs(2955));
    outputs(583) <= not(layer6_outputs(3721));
    outputs(584) <= not(layer6_outputs(517));
    outputs(585) <= not(layer6_outputs(2056)) or (layer6_outputs(4798));
    outputs(586) <= layer6_outputs(64);
    outputs(587) <= not((layer6_outputs(1567)) or (layer6_outputs(1011)));
    outputs(588) <= not(layer6_outputs(4470)) or (layer6_outputs(988));
    outputs(589) <= not((layer6_outputs(1479)) xor (layer6_outputs(3209)));
    outputs(590) <= not(layer6_outputs(3525));
    outputs(591) <= layer6_outputs(2251);
    outputs(592) <= layer6_outputs(3060);
    outputs(593) <= layer6_outputs(3049);
    outputs(594) <= layer6_outputs(4805);
    outputs(595) <= not(layer6_outputs(2983));
    outputs(596) <= not(layer6_outputs(4737));
    outputs(597) <= not(layer6_outputs(1064));
    outputs(598) <= (layer6_outputs(2576)) and (layer6_outputs(887));
    outputs(599) <= layer6_outputs(4972);
    outputs(600) <= layer6_outputs(4651);
    outputs(601) <= (layer6_outputs(906)) and (layer6_outputs(3382));
    outputs(602) <= (layer6_outputs(2556)) and not (layer6_outputs(3298));
    outputs(603) <= layer6_outputs(836);
    outputs(604) <= not(layer6_outputs(4950));
    outputs(605) <= not(layer6_outputs(4417));
    outputs(606) <= not(layer6_outputs(1736));
    outputs(607) <= not(layer6_outputs(4734));
    outputs(608) <= layer6_outputs(4272);
    outputs(609) <= (layer6_outputs(313)) and not (layer6_outputs(4348));
    outputs(610) <= layer6_outputs(1914);
    outputs(611) <= (layer6_outputs(2306)) and not (layer6_outputs(3930));
    outputs(612) <= not(layer6_outputs(4044));
    outputs(613) <= (layer6_outputs(1019)) and not (layer6_outputs(52));
    outputs(614) <= not(layer6_outputs(3608));
    outputs(615) <= not(layer6_outputs(4534));
    outputs(616) <= not(layer6_outputs(3308));
    outputs(617) <= not((layer6_outputs(1116)) xor (layer6_outputs(1921)));
    outputs(618) <= not(layer6_outputs(2850));
    outputs(619) <= layer6_outputs(2103);
    outputs(620) <= not(layer6_outputs(1631)) or (layer6_outputs(3949));
    outputs(621) <= not(layer6_outputs(3620));
    outputs(622) <= not(layer6_outputs(289));
    outputs(623) <= (layer6_outputs(3078)) and not (layer6_outputs(2664));
    outputs(624) <= not(layer6_outputs(657));
    outputs(625) <= not(layer6_outputs(3867));
    outputs(626) <= layer6_outputs(3666);
    outputs(627) <= not(layer6_outputs(4364));
    outputs(628) <= (layer6_outputs(3630)) xor (layer6_outputs(4368));
    outputs(629) <= (layer6_outputs(2892)) and not (layer6_outputs(3796));
    outputs(630) <= not(layer6_outputs(180));
    outputs(631) <= layer6_outputs(1232);
    outputs(632) <= layer6_outputs(631);
    outputs(633) <= not(layer6_outputs(2582));
    outputs(634) <= not(layer6_outputs(1975));
    outputs(635) <= not(layer6_outputs(1141));
    outputs(636) <= not(layer6_outputs(4160));
    outputs(637) <= not(layer6_outputs(4498)) or (layer6_outputs(3375));
    outputs(638) <= not(layer6_outputs(4444));
    outputs(639) <= layer6_outputs(4526);
    outputs(640) <= layer6_outputs(1772);
    outputs(641) <= (layer6_outputs(3430)) and (layer6_outputs(2949));
    outputs(642) <= not(layer6_outputs(528));
    outputs(643) <= not(layer6_outputs(2120));
    outputs(644) <= not(layer6_outputs(1056)) or (layer6_outputs(865));
    outputs(645) <= layer6_outputs(2777);
    outputs(646) <= layer6_outputs(2312);
    outputs(647) <= layer6_outputs(3535);
    outputs(648) <= not(layer6_outputs(4284));
    outputs(649) <= layer6_outputs(4854);
    outputs(650) <= (layer6_outputs(4501)) and not (layer6_outputs(2700));
    outputs(651) <= (layer6_outputs(868)) and (layer6_outputs(3331));
    outputs(652) <= not(layer6_outputs(3422));
    outputs(653) <= (layer6_outputs(4089)) and (layer6_outputs(3486));
    outputs(654) <= not((layer6_outputs(5043)) and (layer6_outputs(4605)));
    outputs(655) <= (layer6_outputs(4841)) xor (layer6_outputs(2196));
    outputs(656) <= layer6_outputs(1182);
    outputs(657) <= not((layer6_outputs(2)) xor (layer6_outputs(3112)));
    outputs(658) <= (layer6_outputs(2473)) and (layer6_outputs(1983));
    outputs(659) <= layer6_outputs(648);
    outputs(660) <= not((layer6_outputs(3038)) xor (layer6_outputs(2068)));
    outputs(661) <= (layer6_outputs(183)) and not (layer6_outputs(1724));
    outputs(662) <= layer6_outputs(4791);
    outputs(663) <= not(layer6_outputs(2453)) or (layer6_outputs(1473));
    outputs(664) <= layer6_outputs(2852);
    outputs(665) <= not(layer6_outputs(4208));
    outputs(666) <= (layer6_outputs(215)) and not (layer6_outputs(5061));
    outputs(667) <= not(layer6_outputs(4494));
    outputs(668) <= not(layer6_outputs(1946));
    outputs(669) <= (layer6_outputs(5065)) and not (layer6_outputs(4736));
    outputs(670) <= layer6_outputs(3049);
    outputs(671) <= (layer6_outputs(1284)) and not (layer6_outputs(3386));
    outputs(672) <= not(layer6_outputs(3051));
    outputs(673) <= layer6_outputs(249);
    outputs(674) <= not((layer6_outputs(2448)) or (layer6_outputs(3306)));
    outputs(675) <= not(layer6_outputs(268)) or (layer6_outputs(870));
    outputs(676) <= (layer6_outputs(2035)) xor (layer6_outputs(2003));
    outputs(677) <= layer6_outputs(4839);
    outputs(678) <= not(layer6_outputs(1681));
    outputs(679) <= not(layer6_outputs(4900));
    outputs(680) <= layer6_outputs(3974);
    outputs(681) <= (layer6_outputs(1345)) and (layer6_outputs(1832));
    outputs(682) <= layer6_outputs(1654);
    outputs(683) <= (layer6_outputs(1617)) and (layer6_outputs(3772));
    outputs(684) <= not(layer6_outputs(1321));
    outputs(685) <= not(layer6_outputs(3657));
    outputs(686) <= not((layer6_outputs(3132)) and (layer6_outputs(201)));
    outputs(687) <= layer6_outputs(4667);
    outputs(688) <= not((layer6_outputs(669)) xor (layer6_outputs(3462)));
    outputs(689) <= (layer6_outputs(708)) xor (layer6_outputs(2366));
    outputs(690) <= (layer6_outputs(1145)) and (layer6_outputs(1750));
    outputs(691) <= not(layer6_outputs(2599));
    outputs(692) <= not(layer6_outputs(1293));
    outputs(693) <= layer6_outputs(2703);
    outputs(694) <= not(layer6_outputs(5095));
    outputs(695) <= not(layer6_outputs(3775));
    outputs(696) <= layer6_outputs(4172);
    outputs(697) <= layer6_outputs(4435);
    outputs(698) <= (layer6_outputs(4512)) and not (layer6_outputs(2751));
    outputs(699) <= not(layer6_outputs(2208));
    outputs(700) <= not(layer6_outputs(441));
    outputs(701) <= (layer6_outputs(1315)) and (layer6_outputs(4355));
    outputs(702) <= not(layer6_outputs(1204));
    outputs(703) <= (layer6_outputs(2371)) xor (layer6_outputs(4690));
    outputs(704) <= (layer6_outputs(4437)) xor (layer6_outputs(4529));
    outputs(705) <= not(layer6_outputs(883));
    outputs(706) <= not(layer6_outputs(3786));
    outputs(707) <= layer6_outputs(3219);
    outputs(708) <= not(layer6_outputs(1211));
    outputs(709) <= not(layer6_outputs(255));
    outputs(710) <= not(layer6_outputs(310));
    outputs(711) <= (layer6_outputs(3582)) xor (layer6_outputs(403));
    outputs(712) <= layer6_outputs(4638);
    outputs(713) <= not(layer6_outputs(4259));
    outputs(714) <= layer6_outputs(357);
    outputs(715) <= not((layer6_outputs(108)) xor (layer6_outputs(2213)));
    outputs(716) <= layer6_outputs(5000);
    outputs(717) <= layer6_outputs(4590);
    outputs(718) <= layer6_outputs(963);
    outputs(719) <= layer6_outputs(2593);
    outputs(720) <= layer6_outputs(3252);
    outputs(721) <= (layer6_outputs(1969)) and not (layer6_outputs(3602));
    outputs(722) <= not(layer6_outputs(1409));
    outputs(723) <= (layer6_outputs(4732)) xor (layer6_outputs(3938));
    outputs(724) <= not(layer6_outputs(2808));
    outputs(725) <= not(layer6_outputs(3501));
    outputs(726) <= not(layer6_outputs(1540));
    outputs(727) <= layer6_outputs(4853);
    outputs(728) <= not(layer6_outputs(2524));
    outputs(729) <= not((layer6_outputs(1459)) xor (layer6_outputs(531)));
    outputs(730) <= (layer6_outputs(1978)) xor (layer6_outputs(4925));
    outputs(731) <= layer6_outputs(2935);
    outputs(732) <= (layer6_outputs(2669)) and not (layer6_outputs(3584));
    outputs(733) <= (layer6_outputs(4120)) and (layer6_outputs(1153));
    outputs(734) <= not(layer6_outputs(2720));
    outputs(735) <= layer6_outputs(4563);
    outputs(736) <= not(layer6_outputs(4247));
    outputs(737) <= (layer6_outputs(2887)) and not (layer6_outputs(2032));
    outputs(738) <= (layer6_outputs(1172)) and not (layer6_outputs(5038));
    outputs(739) <= layer6_outputs(2546);
    outputs(740) <= (layer6_outputs(3090)) and not (layer6_outputs(3638));
    outputs(741) <= layer6_outputs(4596);
    outputs(742) <= (layer6_outputs(450)) and not (layer6_outputs(401));
    outputs(743) <= not((layer6_outputs(350)) xor (layer6_outputs(3253)));
    outputs(744) <= not((layer6_outputs(4403)) or (layer6_outputs(4484)));
    outputs(745) <= (layer6_outputs(2218)) and not (layer6_outputs(1273));
    outputs(746) <= not(layer6_outputs(1623));
    outputs(747) <= not((layer6_outputs(2863)) xor (layer6_outputs(3232)));
    outputs(748) <= not(layer6_outputs(2791));
    outputs(749) <= not(layer6_outputs(2791));
    outputs(750) <= layer6_outputs(1796);
    outputs(751) <= not((layer6_outputs(854)) xor (layer6_outputs(951)));
    outputs(752) <= (layer6_outputs(265)) or (layer6_outputs(3293));
    outputs(753) <= layer6_outputs(2691);
    outputs(754) <= layer6_outputs(3598);
    outputs(755) <= (layer6_outputs(4917)) and not (layer6_outputs(4297));
    outputs(756) <= not((layer6_outputs(3610)) xor (layer6_outputs(4113)));
    outputs(757) <= not(layer6_outputs(5116));
    outputs(758) <= (layer6_outputs(1311)) and not (layer6_outputs(4986));
    outputs(759) <= layer6_outputs(5118);
    outputs(760) <= (layer6_outputs(4590)) and not (layer6_outputs(1505));
    outputs(761) <= (layer6_outputs(1425)) and not (layer6_outputs(3025));
    outputs(762) <= (layer6_outputs(744)) xor (layer6_outputs(2409));
    outputs(763) <= layer6_outputs(2389);
    outputs(764) <= not((layer6_outputs(2197)) xor (layer6_outputs(205)));
    outputs(765) <= (layer6_outputs(2780)) and (layer6_outputs(3763));
    outputs(766) <= not(layer6_outputs(3281)) or (layer6_outputs(2065));
    outputs(767) <= not(layer6_outputs(4375));
    outputs(768) <= (layer6_outputs(2154)) or (layer6_outputs(1388));
    outputs(769) <= not(layer6_outputs(2206));
    outputs(770) <= (layer6_outputs(4008)) and (layer6_outputs(1469));
    outputs(771) <= not(layer6_outputs(129));
    outputs(772) <= layer6_outputs(3974);
    outputs(773) <= (layer6_outputs(3481)) and (layer6_outputs(2147));
    outputs(774) <= not(layer6_outputs(3015));
    outputs(775) <= not((layer6_outputs(1288)) xor (layer6_outputs(291)));
    outputs(776) <= layer6_outputs(1901);
    outputs(777) <= layer6_outputs(3151);
    outputs(778) <= layer6_outputs(4027);
    outputs(779) <= not(layer6_outputs(372));
    outputs(780) <= (layer6_outputs(3426)) and not (layer6_outputs(605));
    outputs(781) <= not(layer6_outputs(1179));
    outputs(782) <= layer6_outputs(4101);
    outputs(783) <= not((layer6_outputs(1276)) or (layer6_outputs(2138)));
    outputs(784) <= not(layer6_outputs(310));
    outputs(785) <= not(layer6_outputs(5105));
    outputs(786) <= (layer6_outputs(179)) xor (layer6_outputs(2726));
    outputs(787) <= not(layer6_outputs(3389));
    outputs(788) <= layer6_outputs(1602);
    outputs(789) <= layer6_outputs(3028);
    outputs(790) <= not(layer6_outputs(4214));
    outputs(791) <= not((layer6_outputs(2028)) xor (layer6_outputs(2840)));
    outputs(792) <= layer6_outputs(2826);
    outputs(793) <= not(layer6_outputs(4914));
    outputs(794) <= (layer6_outputs(3848)) xor (layer6_outputs(1825));
    outputs(795) <= (layer6_outputs(1030)) xor (layer6_outputs(757));
    outputs(796) <= layer6_outputs(3556);
    outputs(797) <= (layer6_outputs(533)) and not (layer6_outputs(2886));
    outputs(798) <= not((layer6_outputs(2111)) xor (layer6_outputs(1897)));
    outputs(799) <= not((layer6_outputs(4180)) or (layer6_outputs(3536)));
    outputs(800) <= not(layer6_outputs(4603));
    outputs(801) <= not(layer6_outputs(2066));
    outputs(802) <= layer6_outputs(2343);
    outputs(803) <= not(layer6_outputs(3952));
    outputs(804) <= layer6_outputs(149);
    outputs(805) <= not((layer6_outputs(1873)) xor (layer6_outputs(4832)));
    outputs(806) <= not((layer6_outputs(679)) or (layer6_outputs(3024)));
    outputs(807) <= layer6_outputs(4901);
    outputs(808) <= layer6_outputs(643);
    outputs(809) <= layer6_outputs(4489);
    outputs(810) <= not(layer6_outputs(4745));
    outputs(811) <= layer6_outputs(58);
    outputs(812) <= (layer6_outputs(4564)) xor (layer6_outputs(287));
    outputs(813) <= not((layer6_outputs(340)) or (layer6_outputs(3017)));
    outputs(814) <= layer6_outputs(2687);
    outputs(815) <= (layer6_outputs(4219)) xor (layer6_outputs(2918));
    outputs(816) <= not(layer6_outputs(4903));
    outputs(817) <= (layer6_outputs(4597)) xor (layer6_outputs(119));
    outputs(818) <= not((layer6_outputs(3265)) xor (layer6_outputs(541)));
    outputs(819) <= layer6_outputs(1904);
    outputs(820) <= not(layer6_outputs(2808));
    outputs(821) <= (layer6_outputs(4438)) and not (layer6_outputs(2434));
    outputs(822) <= not(layer6_outputs(427));
    outputs(823) <= not(layer6_outputs(4359));
    outputs(824) <= layer6_outputs(1202);
    outputs(825) <= (layer6_outputs(3125)) xor (layer6_outputs(2911));
    outputs(826) <= layer6_outputs(1504);
    outputs(827) <= not((layer6_outputs(3311)) xor (layer6_outputs(2630)));
    outputs(828) <= layer6_outputs(2355);
    outputs(829) <= layer6_outputs(3268);
    outputs(830) <= not((layer6_outputs(614)) or (layer6_outputs(1386)));
    outputs(831) <= (layer6_outputs(4867)) and (layer6_outputs(410));
    outputs(832) <= layer6_outputs(1164);
    outputs(833) <= (layer6_outputs(4011)) or (layer6_outputs(3150));
    outputs(834) <= (layer6_outputs(2444)) and not (layer6_outputs(3447));
    outputs(835) <= not(layer6_outputs(2945));
    outputs(836) <= not(layer6_outputs(2552));
    outputs(837) <= (layer6_outputs(4241)) xor (layer6_outputs(2267));
    outputs(838) <= (layer6_outputs(2646)) and (layer6_outputs(2365));
    outputs(839) <= (layer6_outputs(4314)) and (layer6_outputs(638));
    outputs(840) <= layer6_outputs(3077);
    outputs(841) <= layer6_outputs(5001);
    outputs(842) <= not(layer6_outputs(4681));
    outputs(843) <= not(layer6_outputs(697));
    outputs(844) <= layer6_outputs(2606);
    outputs(845) <= not(layer6_outputs(3114));
    outputs(846) <= layer6_outputs(4453);
    outputs(847) <= not((layer6_outputs(4720)) xor (layer6_outputs(2869)));
    outputs(848) <= layer6_outputs(1286);
    outputs(849) <= not((layer6_outputs(1211)) or (layer6_outputs(1783)));
    outputs(850) <= (layer6_outputs(1870)) xor (layer6_outputs(2533));
    outputs(851) <= layer6_outputs(1451);
    outputs(852) <= layer6_outputs(535);
    outputs(853) <= (layer6_outputs(2571)) xor (layer6_outputs(804));
    outputs(854) <= not((layer6_outputs(4980)) xor (layer6_outputs(369)));
    outputs(855) <= layer6_outputs(4517);
    outputs(856) <= layer6_outputs(3970);
    outputs(857) <= not(layer6_outputs(2542));
    outputs(858) <= layer6_outputs(3336);
    outputs(859) <= layer6_outputs(2706);
    outputs(860) <= layer6_outputs(2411);
    outputs(861) <= layer6_outputs(1079);
    outputs(862) <= layer6_outputs(2894);
    outputs(863) <= layer6_outputs(2137);
    outputs(864) <= not(layer6_outputs(2981));
    outputs(865) <= not((layer6_outputs(1450)) and (layer6_outputs(2489)));
    outputs(866) <= not(layer6_outputs(440));
    outputs(867) <= not(layer6_outputs(180));
    outputs(868) <= (layer6_outputs(349)) and not (layer6_outputs(3650));
    outputs(869) <= not((layer6_outputs(1115)) xor (layer6_outputs(3122)));
    outputs(870) <= layer6_outputs(4036);
    outputs(871) <= not((layer6_outputs(4182)) xor (layer6_outputs(1888)));
    outputs(872) <= not((layer6_outputs(2838)) or (layer6_outputs(100)));
    outputs(873) <= not((layer6_outputs(1208)) xor (layer6_outputs(4257)));
    outputs(874) <= layer6_outputs(2889);
    outputs(875) <= not((layer6_outputs(69)) xor (layer6_outputs(2667)));
    outputs(876) <= (layer6_outputs(2233)) and not (layer6_outputs(1272));
    outputs(877) <= (layer6_outputs(2461)) xor (layer6_outputs(2247));
    outputs(878) <= (layer6_outputs(1892)) xor (layer6_outputs(3134));
    outputs(879) <= layer6_outputs(1375);
    outputs(880) <= layer6_outputs(442);
    outputs(881) <= not(layer6_outputs(2761));
    outputs(882) <= (layer6_outputs(2926)) and not (layer6_outputs(3551));
    outputs(883) <= (layer6_outputs(1272)) xor (layer6_outputs(4947));
    outputs(884) <= (layer6_outputs(1784)) and not (layer6_outputs(1418));
    outputs(885) <= not((layer6_outputs(3384)) or (layer6_outputs(2172)));
    outputs(886) <= not(layer6_outputs(2857));
    outputs(887) <= (layer6_outputs(4776)) and (layer6_outputs(4159));
    outputs(888) <= (layer6_outputs(60)) and (layer6_outputs(971));
    outputs(889) <= not(layer6_outputs(298));
    outputs(890) <= not(layer6_outputs(5104));
    outputs(891) <= not(layer6_outputs(1794));
    outputs(892) <= (layer6_outputs(3649)) xor (layer6_outputs(3454));
    outputs(893) <= layer6_outputs(3277);
    outputs(894) <= not(layer6_outputs(2795));
    outputs(895) <= (layer6_outputs(2095)) xor (layer6_outputs(3569));
    outputs(896) <= (layer6_outputs(2919)) and not (layer6_outputs(661));
    outputs(897) <= layer6_outputs(3921);
    outputs(898) <= not(layer6_outputs(858));
    outputs(899) <= (layer6_outputs(4099)) and (layer6_outputs(5113));
    outputs(900) <= layer6_outputs(3092);
    outputs(901) <= not(layer6_outputs(610));
    outputs(902) <= not(layer6_outputs(1256));
    outputs(903) <= not(layer6_outputs(993));
    outputs(904) <= not(layer6_outputs(449));
    outputs(905) <= not(layer6_outputs(1800));
    outputs(906) <= (layer6_outputs(5036)) and not (layer6_outputs(4769));
    outputs(907) <= (layer6_outputs(2490)) and not (layer6_outputs(3419));
    outputs(908) <= (layer6_outputs(4922)) xor (layer6_outputs(4593));
    outputs(909) <= not((layer6_outputs(901)) xor (layer6_outputs(5050)));
    outputs(910) <= not(layer6_outputs(1298));
    outputs(911) <= layer6_outputs(32);
    outputs(912) <= not((layer6_outputs(4379)) xor (layer6_outputs(914)));
    outputs(913) <= layer6_outputs(3840);
    outputs(914) <= not(layer6_outputs(4673));
    outputs(915) <= (layer6_outputs(3552)) and not (layer6_outputs(4926));
    outputs(916) <= '0';
    outputs(917) <= not(layer6_outputs(624));
    outputs(918) <= not(layer6_outputs(1075)) or (layer6_outputs(3664));
    outputs(919) <= not(layer6_outputs(210));
    outputs(920) <= not((layer6_outputs(5016)) or (layer6_outputs(2827)));
    outputs(921) <= not(layer6_outputs(2278));
    outputs(922) <= (layer6_outputs(1271)) and not (layer6_outputs(101));
    outputs(923) <= layer6_outputs(81);
    outputs(924) <= not((layer6_outputs(4886)) or (layer6_outputs(2484)));
    outputs(925) <= not(layer6_outputs(4187));
    outputs(926) <= not(layer6_outputs(1180));
    outputs(927) <= not((layer6_outputs(1928)) and (layer6_outputs(5119)));
    outputs(928) <= not(layer6_outputs(1846));
    outputs(929) <= layer6_outputs(1244);
    outputs(930) <= layer6_outputs(2505);
    outputs(931) <= (layer6_outputs(649)) and (layer6_outputs(45));
    outputs(932) <= (layer6_outputs(1431)) and not (layer6_outputs(762));
    outputs(933) <= layer6_outputs(3984);
    outputs(934) <= not(layer6_outputs(599));
    outputs(935) <= not(layer6_outputs(4581)) or (layer6_outputs(1248));
    outputs(936) <= (layer6_outputs(365)) and (layer6_outputs(1994));
    outputs(937) <= not((layer6_outputs(4879)) xor (layer6_outputs(4979)));
    outputs(938) <= not(layer6_outputs(1475));
    outputs(939) <= not((layer6_outputs(3956)) xor (layer6_outputs(4787)));
    outputs(940) <= (layer6_outputs(2159)) xor (layer6_outputs(1337));
    outputs(941) <= layer6_outputs(4249);
    outputs(942) <= not(layer6_outputs(2393)) or (layer6_outputs(2432));
    outputs(943) <= not(layer6_outputs(2275));
    outputs(944) <= layer6_outputs(2553);
    outputs(945) <= not((layer6_outputs(4908)) xor (layer6_outputs(3682)));
    outputs(946) <= (layer6_outputs(1111)) and (layer6_outputs(5040));
    outputs(947) <= layer6_outputs(2414);
    outputs(948) <= layer6_outputs(3888);
    outputs(949) <= (layer6_outputs(1009)) and not (layer6_outputs(3931));
    outputs(950) <= layer6_outputs(4595);
    outputs(951) <= not(layer6_outputs(4150));
    outputs(952) <= (layer6_outputs(1013)) xor (layer6_outputs(4945));
    outputs(953) <= not(layer6_outputs(1874));
    outputs(954) <= layer6_outputs(4114);
    outputs(955) <= not((layer6_outputs(1948)) xor (layer6_outputs(3399)));
    outputs(956) <= layer6_outputs(3803);
    outputs(957) <= (layer6_outputs(4885)) and not (layer6_outputs(4123));
    outputs(958) <= layer6_outputs(1079);
    outputs(959) <= layer6_outputs(2748);
    outputs(960) <= not(layer6_outputs(314));
    outputs(961) <= not(layer6_outputs(2784));
    outputs(962) <= layer6_outputs(1332);
    outputs(963) <= not(layer6_outputs(2798));
    outputs(964) <= layer6_outputs(563);
    outputs(965) <= not(layer6_outputs(2354));
    outputs(966) <= layer6_outputs(1529);
    outputs(967) <= (layer6_outputs(655)) and not (layer6_outputs(3345));
    outputs(968) <= layer6_outputs(3427);
    outputs(969) <= layer6_outputs(1127);
    outputs(970) <= layer6_outputs(3966);
    outputs(971) <= layer6_outputs(4191);
    outputs(972) <= not(layer6_outputs(115));
    outputs(973) <= not((layer6_outputs(2011)) xor (layer6_outputs(1026)));
    outputs(974) <= layer6_outputs(827);
    outputs(975) <= layer6_outputs(1497);
    outputs(976) <= (layer6_outputs(2885)) and (layer6_outputs(3637));
    outputs(977) <= layer6_outputs(2180);
    outputs(978) <= (layer6_outputs(1357)) xor (layer6_outputs(1958));
    outputs(979) <= not(layer6_outputs(2657));
    outputs(980) <= (layer6_outputs(1605)) xor (layer6_outputs(931));
    outputs(981) <= not(layer6_outputs(955));
    outputs(982) <= layer6_outputs(4078);
    outputs(983) <= layer6_outputs(2422);
    outputs(984) <= not(layer6_outputs(1997));
    outputs(985) <= layer6_outputs(335);
    outputs(986) <= not(layer6_outputs(2113));
    outputs(987) <= not(layer6_outputs(3550));
    outputs(988) <= not(layer6_outputs(4627));
    outputs(989) <= layer6_outputs(267);
    outputs(990) <= (layer6_outputs(5011)) and (layer6_outputs(3469));
    outputs(991) <= not(layer6_outputs(147));
    outputs(992) <= not(layer6_outputs(2765));
    outputs(993) <= not(layer6_outputs(4834));
    outputs(994) <= not(layer6_outputs(2768));
    outputs(995) <= not(layer6_outputs(3864));
    outputs(996) <= (layer6_outputs(1880)) xor (layer6_outputs(2416));
    outputs(997) <= not(layer6_outputs(1503));
    outputs(998) <= layer6_outputs(2559);
    outputs(999) <= layer6_outputs(2498);
    outputs(1000) <= not(layer6_outputs(2479));
    outputs(1001) <= layer6_outputs(2445);
    outputs(1002) <= layer6_outputs(2273);
    outputs(1003) <= (layer6_outputs(4138)) xor (layer6_outputs(4179));
    outputs(1004) <= not(layer6_outputs(1052));
    outputs(1005) <= layer6_outputs(2458);
    outputs(1006) <= (layer6_outputs(3279)) and not (layer6_outputs(3423));
    outputs(1007) <= layer6_outputs(872);
    outputs(1008) <= layer6_outputs(2486);
    outputs(1009) <= (layer6_outputs(3554)) xor (layer6_outputs(1330));
    outputs(1010) <= (layer6_outputs(2013)) and (layer6_outputs(2453));
    outputs(1011) <= (layer6_outputs(289)) xor (layer6_outputs(339));
    outputs(1012) <= not(layer6_outputs(740));
    outputs(1013) <= not((layer6_outputs(2186)) xor (layer6_outputs(1756)));
    outputs(1014) <= not((layer6_outputs(1461)) xor (layer6_outputs(927)));
    outputs(1015) <= (layer6_outputs(949)) and not (layer6_outputs(2436));
    outputs(1016) <= not(layer6_outputs(2656));
    outputs(1017) <= not(layer6_outputs(1936));
    outputs(1018) <= not(layer6_outputs(502));
    outputs(1019) <= (layer6_outputs(1985)) and not (layer6_outputs(308));
    outputs(1020) <= layer6_outputs(4642);
    outputs(1021) <= layer6_outputs(376);
    outputs(1022) <= layer6_outputs(4475);
    outputs(1023) <= (layer6_outputs(2611)) xor (layer6_outputs(3895));
    outputs(1024) <= not(layer6_outputs(4016)) or (layer6_outputs(4517));
    outputs(1025) <= not(layer6_outputs(4217));
    outputs(1026) <= not((layer6_outputs(740)) or (layer6_outputs(656)));
    outputs(1027) <= not(layer6_outputs(857));
    outputs(1028) <= not(layer6_outputs(4469));
    outputs(1029) <= not(layer6_outputs(622));
    outputs(1030) <= not(layer6_outputs(1352));
    outputs(1031) <= layer6_outputs(1252);
    outputs(1032) <= not(layer6_outputs(3800));
    outputs(1033) <= layer6_outputs(3912);
    outputs(1034) <= layer6_outputs(282);
    outputs(1035) <= layer6_outputs(1344);
    outputs(1036) <= not(layer6_outputs(1737));
    outputs(1037) <= not(layer6_outputs(2249));
    outputs(1038) <= not(layer6_outputs(3291));
    outputs(1039) <= not(layer6_outputs(3508));
    outputs(1040) <= layer6_outputs(3222);
    outputs(1041) <= not(layer6_outputs(2116));
    outputs(1042) <= not((layer6_outputs(3232)) and (layer6_outputs(1963)));
    outputs(1043) <= not(layer6_outputs(653)) or (layer6_outputs(2950));
    outputs(1044) <= layer6_outputs(4993);
    outputs(1045) <= layer6_outputs(4598);
    outputs(1046) <= layer6_outputs(881);
    outputs(1047) <= not(layer6_outputs(3435));
    outputs(1048) <= layer6_outputs(3025);
    outputs(1049) <= (layer6_outputs(1341)) xor (layer6_outputs(24));
    outputs(1050) <= (layer6_outputs(4906)) and not (layer6_outputs(1313));
    outputs(1051) <= layer6_outputs(3362);
    outputs(1052) <= not(layer6_outputs(3711)) or (layer6_outputs(3292));
    outputs(1053) <= not(layer6_outputs(3918));
    outputs(1054) <= not(layer6_outputs(2198));
    outputs(1055) <= layer6_outputs(503);
    outputs(1056) <= not((layer6_outputs(1911)) xor (layer6_outputs(2793)));
    outputs(1057) <= not(layer6_outputs(1007));
    outputs(1058) <= not(layer6_outputs(1564));
    outputs(1059) <= layer6_outputs(2481);
    outputs(1060) <= not(layer6_outputs(2604));
    outputs(1061) <= layer6_outputs(1290);
    outputs(1062) <= not(layer6_outputs(413));
    outputs(1063) <= not((layer6_outputs(1663)) and (layer6_outputs(4199)));
    outputs(1064) <= not(layer6_outputs(618));
    outputs(1065) <= layer6_outputs(402);
    outputs(1066) <= not(layer6_outputs(3842));
    outputs(1067) <= (layer6_outputs(2142)) xor (layer6_outputs(387));
    outputs(1068) <= layer6_outputs(396);
    outputs(1069) <= (layer6_outputs(4941)) xor (layer6_outputs(4583));
    outputs(1070) <= layer6_outputs(2296);
    outputs(1071) <= layer6_outputs(2962);
    outputs(1072) <= layer6_outputs(1692);
    outputs(1073) <= layer6_outputs(762);
    outputs(1074) <= not(layer6_outputs(710));
    outputs(1075) <= not(layer6_outputs(3420));
    outputs(1076) <= not(layer6_outputs(2));
    outputs(1077) <= not(layer6_outputs(2667));
    outputs(1078) <= (layer6_outputs(4007)) and not (layer6_outputs(948));
    outputs(1079) <= not(layer6_outputs(845));
    outputs(1080) <= (layer6_outputs(3207)) or (layer6_outputs(4559));
    outputs(1081) <= layer6_outputs(4274);
    outputs(1082) <= layer6_outputs(5095);
    outputs(1083) <= layer6_outputs(4503);
    outputs(1084) <= not((layer6_outputs(3047)) xor (layer6_outputs(824)));
    outputs(1085) <= not(layer6_outputs(572));
    outputs(1086) <= not(layer6_outputs(1527));
    outputs(1087) <= not((layer6_outputs(4100)) xor (layer6_outputs(4795)));
    outputs(1088) <= (layer6_outputs(2215)) and not (layer6_outputs(3704));
    outputs(1089) <= (layer6_outputs(4486)) xor (layer6_outputs(1594));
    outputs(1090) <= not(layer6_outputs(3909));
    outputs(1091) <= layer6_outputs(4165);
    outputs(1092) <= layer6_outputs(3478);
    outputs(1093) <= not(layer6_outputs(5083)) or (layer6_outputs(3701));
    outputs(1094) <= layer6_outputs(104);
    outputs(1095) <= not(layer6_outputs(4870));
    outputs(1096) <= layer6_outputs(2674);
    outputs(1097) <= (layer6_outputs(3226)) and not (layer6_outputs(3118));
    outputs(1098) <= not(layer6_outputs(4460));
    outputs(1099) <= not((layer6_outputs(314)) xor (layer6_outputs(897)));
    outputs(1100) <= layer6_outputs(360);
    outputs(1101) <= (layer6_outputs(169)) and not (layer6_outputs(4926));
    outputs(1102) <= not(layer6_outputs(106));
    outputs(1103) <= not(layer6_outputs(1645));
    outputs(1104) <= not(layer6_outputs(416));
    outputs(1105) <= layer6_outputs(1616);
    outputs(1106) <= layer6_outputs(5042);
    outputs(1107) <= (layer6_outputs(2828)) and not (layer6_outputs(2120));
    outputs(1108) <= not(layer6_outputs(558));
    outputs(1109) <= (layer6_outputs(2523)) and not (layer6_outputs(835));
    outputs(1110) <= not(layer6_outputs(1639)) or (layer6_outputs(2674));
    outputs(1111) <= not(layer6_outputs(2922));
    outputs(1112) <= layer6_outputs(2408);
    outputs(1113) <= layer6_outputs(3482);
    outputs(1114) <= (layer6_outputs(2785)) and not (layer6_outputs(3671));
    outputs(1115) <= layer6_outputs(4911);
    outputs(1116) <= layer6_outputs(2004);
    outputs(1117) <= layer6_outputs(2300);
    outputs(1118) <= (layer6_outputs(1115)) xor (layer6_outputs(3887));
    outputs(1119) <= layer6_outputs(2655);
    outputs(1120) <= not(layer6_outputs(494));
    outputs(1121) <= layer6_outputs(365);
    outputs(1122) <= layer6_outputs(2306);
    outputs(1123) <= (layer6_outputs(2313)) xor (layer6_outputs(2316));
    outputs(1124) <= not(layer6_outputs(2742));
    outputs(1125) <= layer6_outputs(4015);
    outputs(1126) <= not((layer6_outputs(3079)) xor (layer6_outputs(3009)));
    outputs(1127) <= (layer6_outputs(1929)) and (layer6_outputs(92));
    outputs(1128) <= not(layer6_outputs(158)) or (layer6_outputs(2720));
    outputs(1129) <= not(layer6_outputs(2998));
    outputs(1130) <= not(layer6_outputs(4232));
    outputs(1131) <= layer6_outputs(4515);
    outputs(1132) <= layer6_outputs(4298);
    outputs(1133) <= layer6_outputs(4416);
    outputs(1134) <= layer6_outputs(320);
    outputs(1135) <= not((layer6_outputs(3097)) or (layer6_outputs(559)));
    outputs(1136) <= not(layer6_outputs(479));
    outputs(1137) <= not((layer6_outputs(25)) xor (layer6_outputs(2864)));
    outputs(1138) <= layer6_outputs(979);
    outputs(1139) <= not(layer6_outputs(3497));
    outputs(1140) <= layer6_outputs(4095);
    outputs(1141) <= (layer6_outputs(4525)) and (layer6_outputs(696));
    outputs(1142) <= not(layer6_outputs(959));
    outputs(1143) <= (layer6_outputs(2096)) or (layer6_outputs(674));
    outputs(1144) <= layer6_outputs(2029);
    outputs(1145) <= not(layer6_outputs(1142));
    outputs(1146) <= layer6_outputs(3892);
    outputs(1147) <= not(layer6_outputs(4430));
    outputs(1148) <= not(layer6_outputs(1472));
    outputs(1149) <= layer6_outputs(3276);
    outputs(1150) <= (layer6_outputs(1109)) and not (layer6_outputs(4934));
    outputs(1151) <= not((layer6_outputs(2446)) and (layer6_outputs(3350)));
    outputs(1152) <= not(layer6_outputs(3430)) or (layer6_outputs(1957));
    outputs(1153) <= not(layer6_outputs(493));
    outputs(1154) <= layer6_outputs(2775);
    outputs(1155) <= (layer6_outputs(1955)) or (layer6_outputs(1799));
    outputs(1156) <= layer6_outputs(246);
    outputs(1157) <= layer6_outputs(2848);
    outputs(1158) <= not(layer6_outputs(390)) or (layer6_outputs(1918));
    outputs(1159) <= not(layer6_outputs(3638));
    outputs(1160) <= not((layer6_outputs(2642)) xor (layer6_outputs(361)));
    outputs(1161) <= not(layer6_outputs(2579));
    outputs(1162) <= (layer6_outputs(2503)) xor (layer6_outputs(2472));
    outputs(1163) <= (layer6_outputs(1151)) xor (layer6_outputs(4821));
    outputs(1164) <= layer6_outputs(2745);
    outputs(1165) <= layer6_outputs(1613);
    outputs(1166) <= layer6_outputs(3741);
    outputs(1167) <= not((layer6_outputs(820)) or (layer6_outputs(3824)));
    outputs(1168) <= not(layer6_outputs(1687));
    outputs(1169) <= not(layer6_outputs(773));
    outputs(1170) <= not((layer6_outputs(1611)) or (layer6_outputs(823)));
    outputs(1171) <= layer6_outputs(3122);
    outputs(1172) <= (layer6_outputs(3100)) and not (layer6_outputs(1715));
    outputs(1173) <= not(layer6_outputs(1701));
    outputs(1174) <= not(layer6_outputs(1623));
    outputs(1175) <= layer6_outputs(1813);
    outputs(1176) <= layer6_outputs(86);
    outputs(1177) <= not(layer6_outputs(2395));
    outputs(1178) <= layer6_outputs(2811);
    outputs(1179) <= not(layer6_outputs(4123));
    outputs(1180) <= not((layer6_outputs(5078)) or (layer6_outputs(4771)));
    outputs(1181) <= layer6_outputs(4292);
    outputs(1182) <= layer6_outputs(3512);
    outputs(1183) <= not(layer6_outputs(4364));
    outputs(1184) <= layer6_outputs(1082);
    outputs(1185) <= (layer6_outputs(2467)) and not (layer6_outputs(794));
    outputs(1186) <= (layer6_outputs(1903)) xor (layer6_outputs(3019));
    outputs(1187) <= layer6_outputs(3830);
    outputs(1188) <= layer6_outputs(2307);
    outputs(1189) <= (layer6_outputs(3198)) and not (layer6_outputs(4923));
    outputs(1190) <= not(layer6_outputs(4155));
    outputs(1191) <= layer6_outputs(502);
    outputs(1192) <= (layer6_outputs(1540)) xor (layer6_outputs(1570));
    outputs(1193) <= (layer6_outputs(2749)) and not (layer6_outputs(1402));
    outputs(1194) <= layer6_outputs(4942);
    outputs(1195) <= not((layer6_outputs(3756)) or (layer6_outputs(336)));
    outputs(1196) <= not(layer6_outputs(2426));
    outputs(1197) <= not(layer6_outputs(411));
    outputs(1198) <= not(layer6_outputs(3933));
    outputs(1199) <= not(layer6_outputs(995));
    outputs(1200) <= not((layer6_outputs(3492)) xor (layer6_outputs(3253)));
    outputs(1201) <= not((layer6_outputs(4277)) xor (layer6_outputs(3690)));
    outputs(1202) <= (layer6_outputs(3348)) and (layer6_outputs(3368));
    outputs(1203) <= layer6_outputs(1152);
    outputs(1204) <= not(layer6_outputs(647));
    outputs(1205) <= layer6_outputs(1375);
    outputs(1206) <= layer6_outputs(1706);
    outputs(1207) <= not((layer6_outputs(4551)) and (layer6_outputs(1544)));
    outputs(1208) <= (layer6_outputs(4372)) xor (layer6_outputs(2483));
    outputs(1209) <= (layer6_outputs(3467)) and not (layer6_outputs(3665));
    outputs(1210) <= (layer6_outputs(415)) and not (layer6_outputs(4588));
    outputs(1211) <= not((layer6_outputs(2886)) xor (layer6_outputs(102)));
    outputs(1212) <= not(layer6_outputs(2392));
    outputs(1213) <= layer6_outputs(895);
    outputs(1214) <= layer6_outputs(1659);
    outputs(1215) <= not((layer6_outputs(46)) and (layer6_outputs(586)));
    outputs(1216) <= (layer6_outputs(1849)) xor (layer6_outputs(2199));
    outputs(1217) <= not((layer6_outputs(323)) and (layer6_outputs(2391)));
    outputs(1218) <= not((layer6_outputs(404)) and (layer6_outputs(1086)));
    outputs(1219) <= not(layer6_outputs(3055));
    outputs(1220) <= not(layer6_outputs(3060));
    outputs(1221) <= layer6_outputs(4714);
    outputs(1222) <= not(layer6_outputs(1484));
    outputs(1223) <= not(layer6_outputs(2567));
    outputs(1224) <= not(layer6_outputs(2007));
    outputs(1225) <= (layer6_outputs(1690)) xor (layer6_outputs(2368));
    outputs(1226) <= not(layer6_outputs(3517));
    outputs(1227) <= not(layer6_outputs(1927));
    outputs(1228) <= layer6_outputs(522);
    outputs(1229) <= not(layer6_outputs(452));
    outputs(1230) <= layer6_outputs(3175);
    outputs(1231) <= not(layer6_outputs(1878));
    outputs(1232) <= layer6_outputs(94);
    outputs(1233) <= not(layer6_outputs(3725));
    outputs(1234) <= not(layer6_outputs(944));
    outputs(1235) <= (layer6_outputs(3739)) or (layer6_outputs(3768));
    outputs(1236) <= layer6_outputs(4548);
    outputs(1237) <= not(layer6_outputs(4129));
    outputs(1238) <= (layer6_outputs(825)) or (layer6_outputs(4528));
    outputs(1239) <= layer6_outputs(3070);
    outputs(1240) <= layer6_outputs(2202);
    outputs(1241) <= layer6_outputs(3310);
    outputs(1242) <= not(layer6_outputs(1439));
    outputs(1243) <= layer6_outputs(2738);
    outputs(1244) <= not(layer6_outputs(3744));
    outputs(1245) <= layer6_outputs(3748);
    outputs(1246) <= layer6_outputs(933);
    outputs(1247) <= not((layer6_outputs(136)) xor (layer6_outputs(753)));
    outputs(1248) <= layer6_outputs(1306);
    outputs(1249) <= layer6_outputs(3783);
    outputs(1250) <= not(layer6_outputs(2172));
    outputs(1251) <= (layer6_outputs(2917)) xor (layer6_outputs(4593));
    outputs(1252) <= not((layer6_outputs(4301)) or (layer6_outputs(2805)));
    outputs(1253) <= (layer6_outputs(1317)) xor (layer6_outputs(2187));
    outputs(1254) <= not(layer6_outputs(1199));
    outputs(1255) <= (layer6_outputs(1214)) xor (layer6_outputs(1041));
    outputs(1256) <= not(layer6_outputs(412));
    outputs(1257) <= not(layer6_outputs(1922)) or (layer6_outputs(3670));
    outputs(1258) <= not((layer6_outputs(1759)) xor (layer6_outputs(2297)));
    outputs(1259) <= (layer6_outputs(2287)) xor (layer6_outputs(4422));
    outputs(1260) <= layer6_outputs(4829);
    outputs(1261) <= layer6_outputs(2620);
    outputs(1262) <= layer6_outputs(249);
    outputs(1263) <= layer6_outputs(3980);
    outputs(1264) <= not(layer6_outputs(630));
    outputs(1265) <= layer6_outputs(233);
    outputs(1266) <= not((layer6_outputs(1018)) xor (layer6_outputs(157)));
    outputs(1267) <= not((layer6_outputs(671)) xor (layer6_outputs(1088)));
    outputs(1268) <= not(layer6_outputs(3942));
    outputs(1269) <= layer6_outputs(4516);
    outputs(1270) <= layer6_outputs(3712);
    outputs(1271) <= not(layer6_outputs(1210));
    outputs(1272) <= layer6_outputs(1924);
    outputs(1273) <= not(layer6_outputs(3716));
    outputs(1274) <= (layer6_outputs(2687)) or (layer6_outputs(1181));
    outputs(1275) <= not(layer6_outputs(4043));
    outputs(1276) <= not(layer6_outputs(1661));
    outputs(1277) <= layer6_outputs(1742);
    outputs(1278) <= not(layer6_outputs(4794));
    outputs(1279) <= (layer6_outputs(4227)) xor (layer6_outputs(4084));
    outputs(1280) <= not(layer6_outputs(2646));
    outputs(1281) <= layer6_outputs(2699);
    outputs(1282) <= (layer6_outputs(2861)) xor (layer6_outputs(4083));
    outputs(1283) <= not(layer6_outputs(1021));
    outputs(1284) <= not((layer6_outputs(5032)) xor (layer6_outputs(2245)));
    outputs(1285) <= not(layer6_outputs(3606));
    outputs(1286) <= layer6_outputs(4032);
    outputs(1287) <= not(layer6_outputs(3811));
    outputs(1288) <= layer6_outputs(539);
    outputs(1289) <= not((layer6_outputs(3040)) xor (layer6_outputs(145)));
    outputs(1290) <= not(layer6_outputs(5090));
    outputs(1291) <= not(layer6_outputs(1097));
    outputs(1292) <= not((layer6_outputs(4954)) xor (layer6_outputs(4808)));
    outputs(1293) <= not((layer6_outputs(4207)) and (layer6_outputs(3792)));
    outputs(1294) <= layer6_outputs(3916);
    outputs(1295) <= not((layer6_outputs(3099)) and (layer6_outputs(3651)));
    outputs(1296) <= not((layer6_outputs(3237)) and (layer6_outputs(1389)));
    outputs(1297) <= (layer6_outputs(5032)) xor (layer6_outputs(4583));
    outputs(1298) <= layer6_outputs(4614);
    outputs(1299) <= not(layer6_outputs(871));
    outputs(1300) <= layer6_outputs(2739);
    outputs(1301) <= (layer6_outputs(279)) xor (layer6_outputs(3085));
    outputs(1302) <= layer6_outputs(3089);
    outputs(1303) <= not(layer6_outputs(2330));
    outputs(1304) <= (layer6_outputs(1380)) xor (layer6_outputs(3529));
    outputs(1305) <= not(layer6_outputs(491));
    outputs(1306) <= not(layer6_outputs(3335));
    outputs(1307) <= layer6_outputs(2329);
    outputs(1308) <= not(layer6_outputs(1723));
    outputs(1309) <= layer6_outputs(2307);
    outputs(1310) <= layer6_outputs(3999);
    outputs(1311) <= not(layer6_outputs(738)) or (layer6_outputs(2213));
    outputs(1312) <= not(layer6_outputs(4987));
    outputs(1313) <= not(layer6_outputs(3204));
    outputs(1314) <= layer6_outputs(1278);
    outputs(1315) <= not(layer6_outputs(55));
    outputs(1316) <= layer6_outputs(1883);
    outputs(1317) <= layer6_outputs(216);
    outputs(1318) <= layer6_outputs(4324);
    outputs(1319) <= layer6_outputs(204);
    outputs(1320) <= not(layer6_outputs(2609));
    outputs(1321) <= not(layer6_outputs(1097));
    outputs(1322) <= layer6_outputs(3182);
    outputs(1323) <= not(layer6_outputs(4186));
    outputs(1324) <= layer6_outputs(1476);
    outputs(1325) <= not((layer6_outputs(4907)) and (layer6_outputs(4687)));
    outputs(1326) <= layer6_outputs(4894);
    outputs(1327) <= not(layer6_outputs(3347));
    outputs(1328) <= layer6_outputs(2497);
    outputs(1329) <= not(layer6_outputs(446));
    outputs(1330) <= not(layer6_outputs(321));
    outputs(1331) <= not(layer6_outputs(3167));
    outputs(1332) <= not(layer6_outputs(2561));
    outputs(1333) <= not(layer6_outputs(4022));
    outputs(1334) <= (layer6_outputs(1457)) or (layer6_outputs(2985));
    outputs(1335) <= layer6_outputs(1862);
    outputs(1336) <= layer6_outputs(4813);
    outputs(1337) <= (layer6_outputs(3371)) and not (layer6_outputs(5072));
    outputs(1338) <= layer6_outputs(4353);
    outputs(1339) <= layer6_outputs(3087);
    outputs(1340) <= not(layer6_outputs(2626));
    outputs(1341) <= not(layer6_outputs(737));
    outputs(1342) <= layer6_outputs(800);
    outputs(1343) <= not(layer6_outputs(2426));
    outputs(1344) <= not((layer6_outputs(3799)) xor (layer6_outputs(4554)));
    outputs(1345) <= layer6_outputs(1258);
    outputs(1346) <= layer6_outputs(4277);
    outputs(1347) <= (layer6_outputs(1802)) xor (layer6_outputs(2584));
    outputs(1348) <= layer6_outputs(3853);
    outputs(1349) <= (layer6_outputs(846)) xor (layer6_outputs(3195));
    outputs(1350) <= not(layer6_outputs(2651));
    outputs(1351) <= not(layer6_outputs(960));
    outputs(1352) <= not((layer6_outputs(2322)) xor (layer6_outputs(3110)));
    outputs(1353) <= not(layer6_outputs(10));
    outputs(1354) <= not(layer6_outputs(782)) or (layer6_outputs(4695));
    outputs(1355) <= not(layer6_outputs(1227));
    outputs(1356) <= not(layer6_outputs(1513));
    outputs(1357) <= not(layer6_outputs(2053)) or (layer6_outputs(3691));
    outputs(1358) <= not(layer6_outputs(4283));
    outputs(1359) <= (layer6_outputs(2190)) xor (layer6_outputs(3549));
    outputs(1360) <= layer6_outputs(1893);
    outputs(1361) <= not(layer6_outputs(3065));
    outputs(1362) <= (layer6_outputs(3342)) and not (layer6_outputs(3338));
    outputs(1363) <= not((layer6_outputs(2400)) or (layer6_outputs(2207)));
    outputs(1364) <= layer6_outputs(940);
    outputs(1365) <= not(layer6_outputs(2569)) or (layer6_outputs(2175));
    outputs(1366) <= not(layer6_outputs(4803)) or (layer6_outputs(3911));
    outputs(1367) <= not(layer6_outputs(3030));
    outputs(1368) <= (layer6_outputs(4441)) and (layer6_outputs(3695));
    outputs(1369) <= layer6_outputs(3120);
    outputs(1370) <= not(layer6_outputs(1845));
    outputs(1371) <= layer6_outputs(4515);
    outputs(1372) <= (layer6_outputs(2480)) or (layer6_outputs(1975));
    outputs(1373) <= not(layer6_outputs(272));
    outputs(1374) <= (layer6_outputs(1377)) and (layer6_outputs(3271));
    outputs(1375) <= layer6_outputs(4883);
    outputs(1376) <= not(layer6_outputs(4020));
    outputs(1377) <= not(layer6_outputs(2814)) or (layer6_outputs(97));
    outputs(1378) <= not(layer6_outputs(323));
    outputs(1379) <= (layer6_outputs(1514)) and not (layer6_outputs(2702));
    outputs(1380) <= not(layer6_outputs(583));
    outputs(1381) <= (layer6_outputs(1459)) and (layer6_outputs(840));
    outputs(1382) <= not(layer6_outputs(2920));
    outputs(1383) <= not(layer6_outputs(3477));
    outputs(1384) <= layer6_outputs(1068);
    outputs(1385) <= not((layer6_outputs(157)) and (layer6_outputs(1831)));
    outputs(1386) <= layer6_outputs(445);
    outputs(1387) <= not((layer6_outputs(1748)) xor (layer6_outputs(3433)));
    outputs(1388) <= not((layer6_outputs(2718)) or (layer6_outputs(3071)));
    outputs(1389) <= layer6_outputs(4204);
    outputs(1390) <= not(layer6_outputs(1843));
    outputs(1391) <= not(layer6_outputs(330));
    outputs(1392) <= (layer6_outputs(2709)) and (layer6_outputs(4591));
    outputs(1393) <= not(layer6_outputs(5030));
    outputs(1394) <= not(layer6_outputs(5106));
    outputs(1395) <= (layer6_outputs(2560)) and not (layer6_outputs(4485));
    outputs(1396) <= layer6_outputs(3017);
    outputs(1397) <= not(layer6_outputs(4758));
    outputs(1398) <= layer6_outputs(1822);
    outputs(1399) <= not(layer6_outputs(1251));
    outputs(1400) <= (layer6_outputs(2617)) or (layer6_outputs(254));
    outputs(1401) <= layer6_outputs(3809);
    outputs(1402) <= not((layer6_outputs(4115)) and (layer6_outputs(174)));
    outputs(1403) <= layer6_outputs(1343);
    outputs(1404) <= layer6_outputs(1743);
    outputs(1405) <= layer6_outputs(3556);
    outputs(1406) <= not(layer6_outputs(1360));
    outputs(1407) <= not(layer6_outputs(2782));
    outputs(1408) <= not(layer6_outputs(2443));
    outputs(1409) <= not(layer6_outputs(4504));
    outputs(1410) <= not(layer6_outputs(1984));
    outputs(1411) <= layer6_outputs(2872);
    outputs(1412) <= layer6_outputs(4958);
    outputs(1413) <= not(layer6_outputs(3280));
    outputs(1414) <= (layer6_outputs(3294)) xor (layer6_outputs(1930));
    outputs(1415) <= not(layer6_outputs(4368));
    outputs(1416) <= layer6_outputs(4151);
    outputs(1417) <= not((layer6_outputs(2401)) xor (layer6_outputs(864)));
    outputs(1418) <= (layer6_outputs(255)) xor (layer6_outputs(2788));
    outputs(1419) <= not(layer6_outputs(4936));
    outputs(1420) <= layer6_outputs(725);
    outputs(1421) <= not((layer6_outputs(2316)) or (layer6_outputs(1704)));
    outputs(1422) <= not((layer6_outputs(4914)) and (layer6_outputs(3725)));
    outputs(1423) <= layer6_outputs(2289);
    outputs(1424) <= layer6_outputs(2891);
    outputs(1425) <= not(layer6_outputs(2035));
    outputs(1426) <= not(layer6_outputs(2769));
    outputs(1427) <= layer6_outputs(3028);
    outputs(1428) <= not(layer6_outputs(1559));
    outputs(1429) <= layer6_outputs(1968);
    outputs(1430) <= not(layer6_outputs(1069));
    outputs(1431) <= not(layer6_outputs(22));
    outputs(1432) <= layer6_outputs(2708);
    outputs(1433) <= (layer6_outputs(85)) and not (layer6_outputs(4295));
    outputs(1434) <= layer6_outputs(3026);
    outputs(1435) <= not((layer6_outputs(3702)) or (layer6_outputs(2276)));
    outputs(1436) <= not(layer6_outputs(325));
    outputs(1437) <= layer6_outputs(3500);
    outputs(1438) <= not(layer6_outputs(2368));
    outputs(1439) <= (layer6_outputs(3305)) and not (layer6_outputs(379));
    outputs(1440) <= not((layer6_outputs(2830)) xor (layer6_outputs(302)));
    outputs(1441) <= not(layer6_outputs(3119));
    outputs(1442) <= not(layer6_outputs(3031)) or (layer6_outputs(2358));
    outputs(1443) <= layer6_outputs(79);
    outputs(1444) <= not(layer6_outputs(509));
    outputs(1445) <= not(layer6_outputs(2083)) or (layer6_outputs(386));
    outputs(1446) <= layer6_outputs(2912);
    outputs(1447) <= (layer6_outputs(3920)) or (layer6_outputs(797));
    outputs(1448) <= not(layer6_outputs(876)) or (layer6_outputs(251));
    outputs(1449) <= not(layer6_outputs(1138)) or (layer6_outputs(257));
    outputs(1450) <= layer6_outputs(3203);
    outputs(1451) <= not((layer6_outputs(2601)) xor (layer6_outputs(2495)));
    outputs(1452) <= (layer6_outputs(1339)) or (layer6_outputs(4941));
    outputs(1453) <= (layer6_outputs(1038)) and (layer6_outputs(3270));
    outputs(1454) <= layer6_outputs(4081);
    outputs(1455) <= layer6_outputs(312);
    outputs(1456) <= not(layer6_outputs(155));
    outputs(1457) <= (layer6_outputs(2357)) or (layer6_outputs(5112));
    outputs(1458) <= not(layer6_outputs(3160));
    outputs(1459) <= layer6_outputs(4221);
    outputs(1460) <= layer6_outputs(2776);
    outputs(1461) <= not((layer6_outputs(1502)) xor (layer6_outputs(4954)));
    outputs(1462) <= layer6_outputs(3375);
    outputs(1463) <= layer6_outputs(345);
    outputs(1464) <= layer6_outputs(1612);
    outputs(1465) <= not(layer6_outputs(493));
    outputs(1466) <= layer6_outputs(729);
    outputs(1467) <= not(layer6_outputs(948));
    outputs(1468) <= not((layer6_outputs(2011)) xor (layer6_outputs(3139)));
    outputs(1469) <= not(layer6_outputs(4241));
    outputs(1470) <= (layer6_outputs(3135)) xor (layer6_outputs(352));
    outputs(1471) <= not(layer6_outputs(1016));
    outputs(1472) <= not(layer6_outputs(454));
    outputs(1473) <= not(layer6_outputs(3001));
    outputs(1474) <= (layer6_outputs(5119)) and not (layer6_outputs(1168));
    outputs(1475) <= not(layer6_outputs(4154));
    outputs(1476) <= not(layer6_outputs(1633)) or (layer6_outputs(4365));
    outputs(1477) <= layer6_outputs(963);
    outputs(1478) <= layer6_outputs(4832);
    outputs(1479) <= not(layer6_outputs(4059));
    outputs(1480) <= layer6_outputs(4740);
    outputs(1481) <= not(layer6_outputs(3672));
    outputs(1482) <= not(layer6_outputs(1126));
    outputs(1483) <= layer6_outputs(607);
    outputs(1484) <= layer6_outputs(1412);
    outputs(1485) <= layer6_outputs(3199);
    outputs(1486) <= (layer6_outputs(2230)) and not (layer6_outputs(2688));
    outputs(1487) <= layer6_outputs(2140);
    outputs(1488) <= not(layer6_outputs(3324));
    outputs(1489) <= not(layer6_outputs(3944));
    outputs(1490) <= layer6_outputs(84);
    outputs(1491) <= (layer6_outputs(222)) or (layer6_outputs(2321));
    outputs(1492) <= not(layer6_outputs(3714));
    outputs(1493) <= layer6_outputs(16);
    outputs(1494) <= not((layer6_outputs(3337)) or (layer6_outputs(2590)));
    outputs(1495) <= layer6_outputs(1558);
    outputs(1496) <= layer6_outputs(595);
    outputs(1497) <= layer6_outputs(4818);
    outputs(1498) <= layer6_outputs(2250);
    outputs(1499) <= not((layer6_outputs(4474)) and (layer6_outputs(4824)));
    outputs(1500) <= layer6_outputs(233);
    outputs(1501) <= (layer6_outputs(391)) xor (layer6_outputs(2760));
    outputs(1502) <= not(layer6_outputs(3887));
    outputs(1503) <= not(layer6_outputs(813));
    outputs(1504) <= not(layer6_outputs(3460));
    outputs(1505) <= layer6_outputs(1042);
    outputs(1506) <= layer6_outputs(1024);
    outputs(1507) <= not((layer6_outputs(3005)) and (layer6_outputs(2650)));
    outputs(1508) <= not((layer6_outputs(4230)) xor (layer6_outputs(1513)));
    outputs(1509) <= layer6_outputs(260);
    outputs(1510) <= layer6_outputs(2719);
    outputs(1511) <= layer6_outputs(3272);
    outputs(1512) <= not((layer6_outputs(3795)) and (layer6_outputs(3566)));
    outputs(1513) <= (layer6_outputs(574)) or (layer6_outputs(4920));
    outputs(1514) <= not(layer6_outputs(4173));
    outputs(1515) <= not(layer6_outputs(4328));
    outputs(1516) <= (layer6_outputs(1586)) xor (layer6_outputs(3250));
    outputs(1517) <= not((layer6_outputs(3658)) or (layer6_outputs(3516)));
    outputs(1518) <= (layer6_outputs(3519)) xor (layer6_outputs(1287));
    outputs(1519) <= not(layer6_outputs(4308));
    outputs(1520) <= layer6_outputs(3932);
    outputs(1521) <= not((layer6_outputs(2142)) xor (layer6_outputs(421)));
    outputs(1522) <= (layer6_outputs(2652)) and not (layer6_outputs(826));
    outputs(1523) <= layer6_outputs(2872);
    outputs(1524) <= (layer6_outputs(162)) xor (layer6_outputs(88));
    outputs(1525) <= layer6_outputs(3901);
    outputs(1526) <= not(layer6_outputs(2859));
    outputs(1527) <= layer6_outputs(181);
    outputs(1528) <= not(layer6_outputs(2727));
    outputs(1529) <= not(layer6_outputs(3115));
    outputs(1530) <= (layer6_outputs(56)) and not (layer6_outputs(1270));
    outputs(1531) <= layer6_outputs(3859);
    outputs(1532) <= layer6_outputs(4063);
    outputs(1533) <= (layer6_outputs(163)) and not (layer6_outputs(3570));
    outputs(1534) <= layer6_outputs(1913);
    outputs(1535) <= (layer6_outputs(274)) xor (layer6_outputs(4147));
    outputs(1536) <= layer6_outputs(2388);
    outputs(1537) <= not(layer6_outputs(2557)) or (layer6_outputs(3156));
    outputs(1538) <= (layer6_outputs(2046)) or (layer6_outputs(1715));
    outputs(1539) <= layer6_outputs(1963);
    outputs(1540) <= not(layer6_outputs(1161));
    outputs(1541) <= not(layer6_outputs(3795));
    outputs(1542) <= not(layer6_outputs(1112));
    outputs(1543) <= not(layer6_outputs(3160));
    outputs(1544) <= layer6_outputs(2257);
    outputs(1545) <= not(layer6_outputs(3378)) or (layer6_outputs(2862));
    outputs(1546) <= layer6_outputs(2613);
    outputs(1547) <= not(layer6_outputs(3519));
    outputs(1548) <= not(layer6_outputs(1017));
    outputs(1549) <= (layer6_outputs(2376)) xor (layer6_outputs(4490));
    outputs(1550) <= not(layer6_outputs(1432));
    outputs(1551) <= not(layer6_outputs(3969));
    outputs(1552) <= layer6_outputs(144);
    outputs(1553) <= (layer6_outputs(2697)) xor (layer6_outputs(3243));
    outputs(1554) <= not(layer6_outputs(4107));
    outputs(1555) <= layer6_outputs(2826);
    outputs(1556) <= layer6_outputs(2869);
    outputs(1557) <= layer6_outputs(4384);
    outputs(1558) <= (layer6_outputs(768)) xor (layer6_outputs(4408));
    outputs(1559) <= layer6_outputs(732);
    outputs(1560) <= not(layer6_outputs(3503));
    outputs(1561) <= not(layer6_outputs(2734));
    outputs(1562) <= not(layer6_outputs(490));
    outputs(1563) <= (layer6_outputs(1365)) xor (layer6_outputs(1799));
    outputs(1564) <= (layer6_outputs(2240)) and (layer6_outputs(2314));
    outputs(1565) <= not(layer6_outputs(2350));
    outputs(1566) <= not((layer6_outputs(1765)) xor (layer6_outputs(136)));
    outputs(1567) <= not((layer6_outputs(2106)) or (layer6_outputs(1043)));
    outputs(1568) <= not(layer6_outputs(919));
    outputs(1569) <= not(layer6_outputs(1451));
    outputs(1570) <= (layer6_outputs(2308)) and (layer6_outputs(1564));
    outputs(1571) <= layer6_outputs(5045);
    outputs(1572) <= layer6_outputs(2283);
    outputs(1573) <= not((layer6_outputs(2645)) xor (layer6_outputs(778)));
    outputs(1574) <= layer6_outputs(3568);
    outputs(1575) <= not(layer6_outputs(141));
    outputs(1576) <= layer6_outputs(1519);
    outputs(1577) <= not((layer6_outputs(406)) xor (layer6_outputs(4710)));
    outputs(1578) <= not((layer6_outputs(4465)) xor (layer6_outputs(4507)));
    outputs(1579) <= not(layer6_outputs(4349));
    outputs(1580) <= not((layer6_outputs(3913)) xor (layer6_outputs(909)));
    outputs(1581) <= layer6_outputs(122);
    outputs(1582) <= not(layer6_outputs(793));
    outputs(1583) <= layer6_outputs(3065);
    outputs(1584) <= not((layer6_outputs(3531)) xor (layer6_outputs(3703)));
    outputs(1585) <= not(layer6_outputs(3264));
    outputs(1586) <= layer6_outputs(2735);
    outputs(1587) <= not((layer6_outputs(234)) or (layer6_outputs(4904)));
    outputs(1588) <= layer6_outputs(4749);
    outputs(1589) <= not(layer6_outputs(966)) or (layer6_outputs(1305));
    outputs(1590) <= layer6_outputs(4162);
    outputs(1591) <= not(layer6_outputs(2212));
    outputs(1592) <= not(layer6_outputs(3407));
    outputs(1593) <= layer6_outputs(2139);
    outputs(1594) <= not(layer6_outputs(29));
    outputs(1595) <= not(layer6_outputs(2614));
    outputs(1596) <= not(layer6_outputs(3652));
    outputs(1597) <= not(layer6_outputs(2088));
    outputs(1598) <= not(layer6_outputs(4506));
    outputs(1599) <= layer6_outputs(2182);
    outputs(1600) <= layer6_outputs(890);
    outputs(1601) <= not((layer6_outputs(1074)) xor (layer6_outputs(3441)));
    outputs(1602) <= not(layer6_outputs(1860));
    outputs(1603) <= (layer6_outputs(4045)) xor (layer6_outputs(390));
    outputs(1604) <= (layer6_outputs(2293)) and not (layer6_outputs(2633));
    outputs(1605) <= layer6_outputs(2121);
    outputs(1606) <= not(layer6_outputs(2451));
    outputs(1607) <= layer6_outputs(4546);
    outputs(1608) <= not((layer6_outputs(1008)) and (layer6_outputs(112)));
    outputs(1609) <= (layer6_outputs(870)) xor (layer6_outputs(3836));
    outputs(1610) <= (layer6_outputs(2310)) and (layer6_outputs(87));
    outputs(1611) <= layer6_outputs(399);
    outputs(1612) <= not(layer6_outputs(1003));
    outputs(1613) <= layer6_outputs(1580);
    outputs(1614) <= not((layer6_outputs(372)) xor (layer6_outputs(4337)));
    outputs(1615) <= (layer6_outputs(3733)) and (layer6_outputs(1291));
    outputs(1616) <= (layer6_outputs(4531)) and (layer6_outputs(5017));
    outputs(1617) <= not(layer6_outputs(641)) or (layer6_outputs(3199));
    outputs(1618) <= (layer6_outputs(105)) and not (layer6_outputs(4113));
    outputs(1619) <= not(layer6_outputs(1227));
    outputs(1620) <= not(layer6_outputs(123));
    outputs(1621) <= not(layer6_outputs(2476));
    outputs(1622) <= (layer6_outputs(1890)) and not (layer6_outputs(3313));
    outputs(1623) <= (layer6_outputs(4923)) and (layer6_outputs(3164));
    outputs(1624) <= layer6_outputs(5051);
    outputs(1625) <= layer6_outputs(87);
    outputs(1626) <= not(layer6_outputs(841));
    outputs(1627) <= (layer6_outputs(3427)) xor (layer6_outputs(3453));
    outputs(1628) <= not(layer6_outputs(2194));
    outputs(1629) <= layer6_outputs(2136);
    outputs(1630) <= not(layer6_outputs(437));
    outputs(1631) <= layer6_outputs(4831);
    outputs(1632) <= not(layer6_outputs(1941));
    outputs(1633) <= layer6_outputs(988);
    outputs(1634) <= layer6_outputs(1627);
    outputs(1635) <= not(layer6_outputs(1358));
    outputs(1636) <= (layer6_outputs(187)) and (layer6_outputs(3287));
    outputs(1637) <= not(layer6_outputs(968));
    outputs(1638) <= not(layer6_outputs(927));
    outputs(1639) <= (layer6_outputs(3864)) and not (layer6_outputs(1751));
    outputs(1640) <= layer6_outputs(2208);
    outputs(1641) <= layer6_outputs(2542);
    outputs(1642) <= not((layer6_outputs(1744)) xor (layer6_outputs(1899)));
    outputs(1643) <= not(layer6_outputs(3941));
    outputs(1644) <= layer6_outputs(3922);
    outputs(1645) <= not(layer6_outputs(5012));
    outputs(1646) <= not(layer6_outputs(748));
    outputs(1647) <= not(layer6_outputs(1626));
    outputs(1648) <= not((layer6_outputs(1374)) xor (layer6_outputs(4028)));
    outputs(1649) <= layer6_outputs(962);
    outputs(1650) <= layer6_outputs(1028);
    outputs(1651) <= layer6_outputs(5070);
    outputs(1652) <= (layer6_outputs(268)) xor (layer6_outputs(3137));
    outputs(1653) <= (layer6_outputs(271)) and not (layer6_outputs(702));
    outputs(1654) <= layer6_outputs(2888);
    outputs(1655) <= not(layer6_outputs(4366));
    outputs(1656) <= (layer6_outputs(3119)) xor (layer6_outputs(1803));
    outputs(1657) <= layer6_outputs(4683);
    outputs(1658) <= (layer6_outputs(3506)) xor (layer6_outputs(4217));
    outputs(1659) <= (layer6_outputs(2578)) and not (layer6_outputs(104));
    outputs(1660) <= not(layer6_outputs(934));
    outputs(1661) <= not((layer6_outputs(1936)) xor (layer6_outputs(2749)));
    outputs(1662) <= (layer6_outputs(3613)) and not (layer6_outputs(160));
    outputs(1663) <= not((layer6_outputs(780)) xor (layer6_outputs(3812)));
    outputs(1664) <= layer6_outputs(2742);
    outputs(1665) <= not((layer6_outputs(2284)) xor (layer6_outputs(3909)));
    outputs(1666) <= layer6_outputs(4740);
    outputs(1667) <= layer6_outputs(1867);
    outputs(1668) <= (layer6_outputs(4369)) xor (layer6_outputs(2055));
    outputs(1669) <= not((layer6_outputs(1969)) or (layer6_outputs(1763)));
    outputs(1670) <= (layer6_outputs(1712)) xor (layer6_outputs(1789));
    outputs(1671) <= layer6_outputs(3548);
    outputs(1672) <= not(layer6_outputs(3093));
    outputs(1673) <= (layer6_outputs(3233)) and (layer6_outputs(636));
    outputs(1674) <= not(layer6_outputs(651));
    outputs(1675) <= (layer6_outputs(2640)) xor (layer6_outputs(2750));
    outputs(1676) <= not(layer6_outputs(1583));
    outputs(1677) <= layer6_outputs(750);
    outputs(1678) <= not(layer6_outputs(4436));
    outputs(1679) <= not(layer6_outputs(1922));
    outputs(1680) <= not((layer6_outputs(3982)) or (layer6_outputs(2879)));
    outputs(1681) <= layer6_outputs(2508);
    outputs(1682) <= (layer6_outputs(4346)) xor (layer6_outputs(1667));
    outputs(1683) <= not(layer6_outputs(3033));
    outputs(1684) <= not((layer6_outputs(3747)) xor (layer6_outputs(4731)));
    outputs(1685) <= not((layer6_outputs(1092)) xor (layer6_outputs(1757)));
    outputs(1686) <= layer6_outputs(1166);
    outputs(1687) <= layer6_outputs(546);
    outputs(1688) <= layer6_outputs(568);
    outputs(1689) <= not(layer6_outputs(1881));
    outputs(1690) <= (layer6_outputs(1724)) or (layer6_outputs(4877));
    outputs(1691) <= layer6_outputs(2897);
    outputs(1692) <= (layer6_outputs(91)) xor (layer6_outputs(1089));
    outputs(1693) <= layer6_outputs(975);
    outputs(1694) <= (layer6_outputs(1251)) xor (layer6_outputs(496));
    outputs(1695) <= not(layer6_outputs(571));
    outputs(1696) <= not(layer6_outputs(1339));
    outputs(1697) <= not((layer6_outputs(2040)) xor (layer6_outputs(2931)));
    outputs(1698) <= layer6_outputs(2607);
    outputs(1699) <= (layer6_outputs(4989)) and not (layer6_outputs(1014));
    outputs(1700) <= layer6_outputs(3162);
    outputs(1701) <= not(layer6_outputs(950));
    outputs(1702) <= not((layer6_outputs(495)) xor (layer6_outputs(3700)));
    outputs(1703) <= layer6_outputs(1578);
    outputs(1704) <= layer6_outputs(1986);
    outputs(1705) <= (layer6_outputs(923)) or (layer6_outputs(267));
    outputs(1706) <= not(layer6_outputs(3098));
    outputs(1707) <= layer6_outputs(2817);
    outputs(1708) <= not(layer6_outputs(3579));
    outputs(1709) <= not(layer6_outputs(4818));
    outputs(1710) <= layer6_outputs(1025);
    outputs(1711) <= not(layer6_outputs(1449));
    outputs(1712) <= not(layer6_outputs(4617));
    outputs(1713) <= layer6_outputs(3548);
    outputs(1714) <= not(layer6_outputs(2904));
    outputs(1715) <= layer6_outputs(4791);
    outputs(1716) <= layer6_outputs(3622);
    outputs(1717) <= (layer6_outputs(1849)) xor (layer6_outputs(4014));
    outputs(1718) <= layer6_outputs(2858);
    outputs(1719) <= layer6_outputs(3566);
    outputs(1720) <= not((layer6_outputs(3661)) xor (layer6_outputs(4741)));
    outputs(1721) <= layer6_outputs(2425);
    outputs(1722) <= (layer6_outputs(2087)) and not (layer6_outputs(94));
    outputs(1723) <= (layer6_outputs(3934)) and not (layer6_outputs(4975));
    outputs(1724) <= (layer6_outputs(1658)) and (layer6_outputs(3699));
    outputs(1725) <= not(layer6_outputs(394));
    outputs(1726) <= layer6_outputs(2566);
    outputs(1727) <= layer6_outputs(4244);
    outputs(1728) <= (layer6_outputs(2514)) and not (layer6_outputs(1883));
    outputs(1729) <= (layer6_outputs(4073)) and not (layer6_outputs(867));
    outputs(1730) <= not((layer6_outputs(1295)) xor (layer6_outputs(5054)));
    outputs(1731) <= not((layer6_outputs(928)) xor (layer6_outputs(1598)));
    outputs(1732) <= not(layer6_outputs(2455)) or (layer6_outputs(4247));
    outputs(1733) <= (layer6_outputs(2419)) and not (layer6_outputs(100));
    outputs(1734) <= (layer6_outputs(4023)) and (layer6_outputs(589));
    outputs(1735) <= not(layer6_outputs(547));
    outputs(1736) <= not(layer6_outputs(4575));
    outputs(1737) <= layer6_outputs(3358);
    outputs(1738) <= not(layer6_outputs(4068));
    outputs(1739) <= layer6_outputs(4153);
    outputs(1740) <= not(layer6_outputs(4172));
    outputs(1741) <= layer6_outputs(3015);
    outputs(1742) <= layer6_outputs(429);
    outputs(1743) <= (layer6_outputs(2054)) xor (layer6_outputs(2370));
    outputs(1744) <= (layer6_outputs(2322)) or (layer6_outputs(4012));
    outputs(1745) <= not((layer6_outputs(4696)) or (layer6_outputs(237)));
    outputs(1746) <= layer6_outputs(3249);
    outputs(1747) <= not(layer6_outputs(4896));
    outputs(1748) <= not(layer6_outputs(4764)) or (layer6_outputs(1179));
    outputs(1749) <= not(layer6_outputs(4532));
    outputs(1750) <= layer6_outputs(2583);
    outputs(1751) <= (layer6_outputs(1943)) and (layer6_outputs(4800));
    outputs(1752) <= (layer6_outputs(2203)) xor (layer6_outputs(2762));
    outputs(1753) <= layer6_outputs(1453);
    outputs(1754) <= layer6_outputs(1950);
    outputs(1755) <= layer6_outputs(859);
    outputs(1756) <= not(layer6_outputs(3730));
    outputs(1757) <= not(layer6_outputs(2047));
    outputs(1758) <= layer6_outputs(4690);
    outputs(1759) <= layer6_outputs(809);
    outputs(1760) <= (layer6_outputs(4742)) xor (layer6_outputs(3659));
    outputs(1761) <= layer6_outputs(668);
    outputs(1762) <= not(layer6_outputs(469));
    outputs(1763) <= (layer6_outputs(970)) xor (layer6_outputs(4686));
    outputs(1764) <= not(layer6_outputs(1548));
    outputs(1765) <= layer6_outputs(176);
    outputs(1766) <= (layer6_outputs(3055)) and (layer6_outputs(5024));
    outputs(1767) <= layer6_outputs(4491);
    outputs(1768) <= not(layer6_outputs(2554));
    outputs(1769) <= layer6_outputs(1624);
    outputs(1770) <= layer6_outputs(2732);
    outputs(1771) <= not(layer6_outputs(3844));
    outputs(1772) <= not(layer6_outputs(759));
    outputs(1773) <= layer6_outputs(402);
    outputs(1774) <= not(layer6_outputs(4371));
    outputs(1775) <= not(layer6_outputs(4540));
    outputs(1776) <= not((layer6_outputs(4615)) xor (layer6_outputs(204)));
    outputs(1777) <= layer6_outputs(256);
    outputs(1778) <= (layer6_outputs(2009)) xor (layer6_outputs(2757));
    outputs(1779) <= not(layer6_outputs(437)) or (layer6_outputs(4079));
    outputs(1780) <= not(layer6_outputs(3954));
    outputs(1781) <= layer6_outputs(3790);
    outputs(1782) <= layer6_outputs(969);
    outputs(1783) <= not((layer6_outputs(3296)) and (layer6_outputs(2381)));
    outputs(1784) <= not(layer6_outputs(956));
    outputs(1785) <= layer6_outputs(1816);
    outputs(1786) <= not(layer6_outputs(363));
    outputs(1787) <= not(layer6_outputs(1333));
    outputs(1788) <= not(layer6_outputs(2626));
    outputs(1789) <= layer6_outputs(905);
    outputs(1790) <= layer6_outputs(4307);
    outputs(1791) <= (layer6_outputs(1169)) and (layer6_outputs(2963));
    outputs(1792) <= not(layer6_outputs(706)) or (layer6_outputs(1136));
    outputs(1793) <= layer6_outputs(1935);
    outputs(1794) <= not((layer6_outputs(4967)) xor (layer6_outputs(3242)));
    outputs(1795) <= (layer6_outputs(197)) xor (layer6_outputs(3086));
    outputs(1796) <= not(layer6_outputs(489));
    outputs(1797) <= not(layer6_outputs(1579));
    outputs(1798) <= not(layer6_outputs(2420));
    outputs(1799) <= layer6_outputs(2910);
    outputs(1800) <= not(layer6_outputs(3724));
    outputs(1801) <= layer6_outputs(882);
    outputs(1802) <= layer6_outputs(669);
    outputs(1803) <= layer6_outputs(3074);
    outputs(1804) <= (layer6_outputs(332)) xor (layer6_outputs(2853));
    outputs(1805) <= not(layer6_outputs(3987));
    outputs(1806) <= not(layer6_outputs(2108));
    outputs(1807) <= not(layer6_outputs(638));
    outputs(1808) <= not(layer6_outputs(490));
    outputs(1809) <= (layer6_outputs(2015)) or (layer6_outputs(4571));
    outputs(1810) <= not(layer6_outputs(2092));
    outputs(1811) <= layer6_outputs(962);
    outputs(1812) <= layer6_outputs(4883);
    outputs(1813) <= layer6_outputs(3283);
    outputs(1814) <= not(layer6_outputs(280));
    outputs(1815) <= layer6_outputs(5112);
    outputs(1816) <= layer6_outputs(3765);
    outputs(1817) <= (layer6_outputs(5011)) or (layer6_outputs(712));
    outputs(1818) <= not(layer6_outputs(2350));
    outputs(1819) <= layer6_outputs(2585);
    outputs(1820) <= layer6_outputs(2379);
    outputs(1821) <= (layer6_outputs(3271)) and (layer6_outputs(1566));
    outputs(1822) <= (layer6_outputs(3284)) and (layer6_outputs(4377));
    outputs(1823) <= layer6_outputs(3558);
    outputs(1824) <= not(layer6_outputs(910));
    outputs(1825) <= layer6_outputs(1792);
    outputs(1826) <= not(layer6_outputs(4564));
    outputs(1827) <= (layer6_outputs(1287)) and (layer6_outputs(3756));
    outputs(1828) <= not(layer6_outputs(3177));
    outputs(1829) <= (layer6_outputs(629)) and not (layer6_outputs(3220));
    outputs(1830) <= not(layer6_outputs(2207));
    outputs(1831) <= not((layer6_outputs(4577)) xor (layer6_outputs(3686)));
    outputs(1832) <= not(layer6_outputs(1382));
    outputs(1833) <= not(layer6_outputs(2373));
    outputs(1834) <= (layer6_outputs(1330)) xor (layer6_outputs(2634));
    outputs(1835) <= layer6_outputs(5060);
    outputs(1836) <= layer6_outputs(1430);
    outputs(1837) <= not(layer6_outputs(645));
    outputs(1838) <= not(layer6_outputs(4409));
    outputs(1839) <= not(layer6_outputs(4397));
    outputs(1840) <= layer6_outputs(4157);
    outputs(1841) <= layer6_outputs(2219);
    outputs(1842) <= layer6_outputs(3885);
    outputs(1843) <= not(layer6_outputs(2672)) or (layer6_outputs(1685));
    outputs(1844) <= not((layer6_outputs(3639)) xor (layer6_outputs(33)));
    outputs(1845) <= layer6_outputs(3178);
    outputs(1846) <= not(layer6_outputs(597));
    outputs(1847) <= layer6_outputs(1391);
    outputs(1848) <= not(layer6_outputs(2660));
    outputs(1849) <= not(layer6_outputs(1449));
    outputs(1850) <= layer6_outputs(477);
    outputs(1851) <= not(layer6_outputs(3591)) or (layer6_outputs(4315));
    outputs(1852) <= layer6_outputs(3094);
    outputs(1853) <= not((layer6_outputs(1025)) xor (layer6_outputs(4659)));
    outputs(1854) <= layer6_outputs(1515);
    outputs(1855) <= layer6_outputs(1572);
    outputs(1856) <= not((layer6_outputs(1901)) or (layer6_outputs(2691)));
    outputs(1857) <= (layer6_outputs(3364)) xor (layer6_outputs(2804));
    outputs(1858) <= not(layer6_outputs(5015));
    outputs(1859) <= not(layer6_outputs(2781));
    outputs(1860) <= not((layer6_outputs(3827)) and (layer6_outputs(3579)));
    outputs(1861) <= not(layer6_outputs(4440)) or (layer6_outputs(4208));
    outputs(1862) <= (layer6_outputs(193)) xor (layer6_outputs(1937));
    outputs(1863) <= (layer6_outputs(4584)) xor (layer6_outputs(3264));
    outputs(1864) <= layer6_outputs(2610);
    outputs(1865) <= not(layer6_outputs(2412));
    outputs(1866) <= not(layer6_outputs(259));
    outputs(1867) <= not(layer6_outputs(1782));
    outputs(1868) <= (layer6_outputs(4918)) or (layer6_outputs(4193));
    outputs(1869) <= layer6_outputs(1347);
    outputs(1870) <= not(layer6_outputs(3693)) or (layer6_outputs(4092));
    outputs(1871) <= layer6_outputs(3557);
    outputs(1872) <= (layer6_outputs(2509)) xor (layer6_outputs(1978));
    outputs(1873) <= not(layer6_outputs(3168));
    outputs(1874) <= (layer6_outputs(4398)) and not (layer6_outputs(5039));
    outputs(1875) <= not(layer6_outputs(3652));
    outputs(1876) <= not(layer6_outputs(904));
    outputs(1877) <= layer6_outputs(5027);
    outputs(1878) <= layer6_outputs(2261);
    outputs(1879) <= (layer6_outputs(2823)) xor (layer6_outputs(3612));
    outputs(1880) <= not(layer6_outputs(4511));
    outputs(1881) <= not((layer6_outputs(3460)) xor (layer6_outputs(2525)));
    outputs(1882) <= layer6_outputs(709);
    outputs(1883) <= layer6_outputs(73);
    outputs(1884) <= (layer6_outputs(3692)) and not (layer6_outputs(5018));
    outputs(1885) <= layer6_outputs(3327);
    outputs(1886) <= layer6_outputs(3670);
    outputs(1887) <= layer6_outputs(4391);
    outputs(1888) <= (layer6_outputs(4588)) and not (layer6_outputs(2855));
    outputs(1889) <= (layer6_outputs(2976)) and not (layer6_outputs(1490));
    outputs(1890) <= layer6_outputs(635);
    outputs(1891) <= layer6_outputs(4513);
    outputs(1892) <= layer6_outputs(3595);
    outputs(1893) <= not((layer6_outputs(5094)) xor (layer6_outputs(4872)));
    outputs(1894) <= layer6_outputs(1714);
    outputs(1895) <= (layer6_outputs(1848)) or (layer6_outputs(2766));
    outputs(1896) <= layer6_outputs(4611);
    outputs(1897) <= layer6_outputs(663);
    outputs(1898) <= layer6_outputs(684);
    outputs(1899) <= layer6_outputs(511);
    outputs(1900) <= not(layer6_outputs(2249));
    outputs(1901) <= layer6_outputs(633);
    outputs(1902) <= (layer6_outputs(4632)) xor (layer6_outputs(4146));
    outputs(1903) <= layer6_outputs(4887);
    outputs(1904) <= not(layer6_outputs(2659));
    outputs(1905) <= layer6_outputs(4512);
    outputs(1906) <= layer6_outputs(945);
    outputs(1907) <= layer6_outputs(2716);
    outputs(1908) <= layer6_outputs(1787);
    outputs(1909) <= not(layer6_outputs(4040));
    outputs(1910) <= not(layer6_outputs(451));
    outputs(1911) <= not(layer6_outputs(1856));
    outputs(1912) <= layer6_outputs(4477);
    outputs(1913) <= layer6_outputs(977);
    outputs(1914) <= not((layer6_outputs(1923)) and (layer6_outputs(3778)));
    outputs(1915) <= layer6_outputs(894);
    outputs(1916) <= layer6_outputs(1332);
    outputs(1917) <= (layer6_outputs(1976)) and not (layer6_outputs(4959));
    outputs(1918) <= not(layer6_outputs(2398));
    outputs(1919) <= not(layer6_outputs(557));
    outputs(1920) <= not(layer6_outputs(4163));
    outputs(1921) <= not(layer6_outputs(4093));
    outputs(1922) <= not((layer6_outputs(3937)) or (layer6_outputs(4920)));
    outputs(1923) <= layer6_outputs(34);
    outputs(1924) <= (layer6_outputs(73)) and (layer6_outputs(2621));
    outputs(1925) <= not(layer6_outputs(1299));
    outputs(1926) <= not(layer6_outputs(459));
    outputs(1927) <= (layer6_outputs(4912)) xor (layer6_outputs(3098));
    outputs(1928) <= not(layer6_outputs(3198));
    outputs(1929) <= not((layer6_outputs(2612)) and (layer6_outputs(4968)));
    outputs(1930) <= not(layer6_outputs(2581));
    outputs(1931) <= not(layer6_outputs(515));
    outputs(1932) <= layer6_outputs(4507);
    outputs(1933) <= (layer6_outputs(1734)) or (layer6_outputs(4803));
    outputs(1934) <= layer6_outputs(2478);
    outputs(1935) <= layer6_outputs(2708);
    outputs(1936) <= not(layer6_outputs(3130));
    outputs(1937) <= (layer6_outputs(3352)) or (layer6_outputs(1284));
    outputs(1938) <= not(layer6_outputs(4956));
    outputs(1939) <= not(layer6_outputs(3960));
    outputs(1940) <= layer6_outputs(3607);
    outputs(1941) <= layer6_outputs(3087);
    outputs(1942) <= layer6_outputs(3409);
    outputs(1943) <= (layer6_outputs(694)) and not (layer6_outputs(901));
    outputs(1944) <= (layer6_outputs(4581)) and (layer6_outputs(4187));
    outputs(1945) <= not(layer6_outputs(182));
    outputs(1946) <= (layer6_outputs(1186)) xor (layer6_outputs(3186));
    outputs(1947) <= (layer6_outputs(1829)) and not (layer6_outputs(4838));
    outputs(1948) <= (layer6_outputs(2166)) xor (layer6_outputs(3166));
    outputs(1949) <= (layer6_outputs(2370)) or (layer6_outputs(5004));
    outputs(1950) <= layer6_outputs(1624);
    outputs(1951) <= not(layer6_outputs(593));
    outputs(1952) <= not(layer6_outputs(1427));
    outputs(1953) <= layer6_outputs(5057);
    outputs(1954) <= layer6_outputs(2305);
    outputs(1955) <= not(layer6_outputs(140));
    outputs(1956) <= (layer6_outputs(2090)) and not (layer6_outputs(3823));
    outputs(1957) <= layer6_outputs(850);
    outputs(1958) <= not((layer6_outputs(3176)) xor (layer6_outputs(4058)));
    outputs(1959) <= not(layer6_outputs(1893));
    outputs(1960) <= (layer6_outputs(1921)) and not (layer6_outputs(2206));
    outputs(1961) <= layer6_outputs(1391);
    outputs(1962) <= (layer6_outputs(2054)) or (layer6_outputs(3302));
    outputs(1963) <= layer6_outputs(1747);
    outputs(1964) <= layer6_outputs(4270);
    outputs(1965) <= not(layer6_outputs(125));
    outputs(1966) <= layer6_outputs(2165);
    outputs(1967) <= layer6_outputs(839);
    outputs(1968) <= layer6_outputs(1734);
    outputs(1969) <= not((layer6_outputs(2563)) xor (layer6_outputs(3067)));
    outputs(1970) <= not(layer6_outputs(1060)) or (layer6_outputs(4981));
    outputs(1971) <= not(layer6_outputs(657));
    outputs(1972) <= not(layer6_outputs(4939)) or (layer6_outputs(4493));
    outputs(1973) <= not(layer6_outputs(1191));
    outputs(1974) <= not((layer6_outputs(2432)) or (layer6_outputs(4909)));
    outputs(1975) <= layer6_outputs(653);
    outputs(1976) <= layer6_outputs(565);
    outputs(1977) <= not(layer6_outputs(661));
    outputs(1978) <= not(layer6_outputs(178));
    outputs(1979) <= not(layer6_outputs(585));
    outputs(1980) <= layer6_outputs(3790);
    outputs(1981) <= layer6_outputs(1866);
    outputs(1982) <= not((layer6_outputs(3329)) xor (layer6_outputs(1224)));
    outputs(1983) <= (layer6_outputs(1703)) xor (layer6_outputs(474));
    outputs(1984) <= not(layer6_outputs(4280));
    outputs(1985) <= not(layer6_outputs(2994));
    outputs(1986) <= layer6_outputs(2959);
    outputs(1987) <= not(layer6_outputs(1531));
    outputs(1988) <= not(layer6_outputs(1040));
    outputs(1989) <= layer6_outputs(909);
    outputs(1990) <= layer6_outputs(4348);
    outputs(1991) <= not(layer6_outputs(330));
    outputs(1992) <= not(layer6_outputs(1098));
    outputs(1993) <= layer6_outputs(699);
    outputs(1994) <= (layer6_outputs(4069)) xor (layer6_outputs(4680));
    outputs(1995) <= not(layer6_outputs(3134));
    outputs(1996) <= layer6_outputs(151);
    outputs(1997) <= layer6_outputs(4811);
    outputs(1998) <= (layer6_outputs(1587)) xor (layer6_outputs(1447));
    outputs(1999) <= not(layer6_outputs(4949));
    outputs(2000) <= not(layer6_outputs(4409));
    outputs(2001) <= not((layer6_outputs(727)) or (layer6_outputs(1387)));
    outputs(2002) <= (layer6_outputs(416)) and (layer6_outputs(1742));
    outputs(2003) <= not(layer6_outputs(1006));
    outputs(2004) <= layer6_outputs(4921);
    outputs(2005) <= (layer6_outputs(5023)) xor (layer6_outputs(1887));
    outputs(2006) <= layer6_outputs(1133);
    outputs(2007) <= layer6_outputs(4549);
    outputs(2008) <= not(layer6_outputs(2786));
    outputs(2009) <= not(layer6_outputs(4623));
    outputs(2010) <= not(layer6_outputs(1132));
    outputs(2011) <= layer6_outputs(3805);
    outputs(2012) <= layer6_outputs(2896);
    outputs(2013) <= not(layer6_outputs(3969));
    outputs(2014) <= layer6_outputs(1314);
    outputs(2015) <= layer6_outputs(4539);
    outputs(2016) <= (layer6_outputs(5105)) and not (layer6_outputs(3872));
    outputs(2017) <= layer6_outputs(3030);
    outputs(2018) <= layer6_outputs(1378);
    outputs(2019) <= layer6_outputs(3162);
    outputs(2020) <= layer6_outputs(27);
    outputs(2021) <= not(layer6_outputs(959));
    outputs(2022) <= not(layer6_outputs(2349));
    outputs(2023) <= not(layer6_outputs(3774));
    outputs(2024) <= not((layer6_outputs(4933)) xor (layer6_outputs(3043)));
    outputs(2025) <= not(layer6_outputs(1390));
    outputs(2026) <= layer6_outputs(1279);
    outputs(2027) <= layer6_outputs(4248);
    outputs(2028) <= layer6_outputs(1869);
    outputs(2029) <= (layer6_outputs(4417)) and not (layer6_outputs(2369));
    outputs(2030) <= layer6_outputs(4331);
    outputs(2031) <= (layer6_outputs(627)) and (layer6_outputs(4598));
    outputs(2032) <= not(layer6_outputs(4774));
    outputs(2033) <= not(layer6_outputs(1573));
    outputs(2034) <= layer6_outputs(4424);
    outputs(2035) <= not((layer6_outputs(219)) or (layer6_outputs(4057)));
    outputs(2036) <= not(layer6_outputs(727));
    outputs(2037) <= (layer6_outputs(4542)) xor (layer6_outputs(4189));
    outputs(2038) <= not((layer6_outputs(80)) or (layer6_outputs(4331)));
    outputs(2039) <= not((layer6_outputs(4352)) xor (layer6_outputs(1162)));
    outputs(2040) <= layer6_outputs(2989);
    outputs(2041) <= not(layer6_outputs(1308));
    outputs(2042) <= (layer6_outputs(1931)) or (layer6_outputs(3141));
    outputs(2043) <= not((layer6_outputs(2905)) or (layer6_outputs(3553)));
    outputs(2044) <= not(layer6_outputs(264));
    outputs(2045) <= not((layer6_outputs(2878)) xor (layer6_outputs(2186)));
    outputs(2046) <= not(layer6_outputs(2996));
    outputs(2047) <= layer6_outputs(4835);
    outputs(2048) <= layer6_outputs(1201);
    outputs(2049) <= not((layer6_outputs(3930)) xor (layer6_outputs(2090)));
    outputs(2050) <= layer6_outputs(2908);
    outputs(2051) <= not(layer6_outputs(4644));
    outputs(2052) <= layer6_outputs(3879);
    outputs(2053) <= not(layer6_outputs(221));
    outputs(2054) <= layer6_outputs(4563);
    outputs(2055) <= not(layer6_outputs(1461));
    outputs(2056) <= (layer6_outputs(1420)) xor (layer6_outputs(1184));
    outputs(2057) <= not((layer6_outputs(3262)) xor (layer6_outputs(2526)));
    outputs(2058) <= not(layer6_outputs(1777));
    outputs(2059) <= not((layer6_outputs(2258)) or (layer6_outputs(121)));
    outputs(2060) <= (layer6_outputs(698)) and not (layer6_outputs(2289));
    outputs(2061) <= layer6_outputs(4682);
    outputs(2062) <= not((layer6_outputs(4911)) xor (layer6_outputs(704)));
    outputs(2063) <= layer6_outputs(1428);
    outputs(2064) <= (layer6_outputs(3006)) xor (layer6_outputs(4725));
    outputs(2065) <= not(layer6_outputs(2664));
    outputs(2066) <= not(layer6_outputs(847));
    outputs(2067) <= not(layer6_outputs(2231));
    outputs(2068) <= layer6_outputs(3411);
    outputs(2069) <= not(layer6_outputs(2824));
    outputs(2070) <= not((layer6_outputs(2463)) and (layer6_outputs(3906)));
    outputs(2071) <= layer6_outputs(5039);
    outputs(2072) <= not(layer6_outputs(647));
    outputs(2073) <= layer6_outputs(3994);
    outputs(2074) <= layer6_outputs(1110);
    outputs(2075) <= not((layer6_outputs(3035)) xor (layer6_outputs(2398)));
    outputs(2076) <= not(layer6_outputs(2719));
    outputs(2077) <= not(layer6_outputs(5041));
    outputs(2078) <= layer6_outputs(3933);
    outputs(2079) <= not(layer6_outputs(4168));
    outputs(2080) <= not(layer6_outputs(2614));
    outputs(2081) <= not(layer6_outputs(4888));
    outputs(2082) <= layer6_outputs(2547);
    outputs(2083) <= not(layer6_outputs(755));
    outputs(2084) <= not(layer6_outputs(3363)) or (layer6_outputs(1749));
    outputs(2085) <= not(layer6_outputs(2033));
    outputs(2086) <= not(layer6_outputs(2834));
    outputs(2087) <= layer6_outputs(440);
    outputs(2088) <= not((layer6_outputs(2154)) xor (layer6_outputs(1047)));
    outputs(2089) <= layer6_outputs(1349);
    outputs(2090) <= not((layer6_outputs(4709)) and (layer6_outputs(232)));
    outputs(2091) <= layer6_outputs(2353);
    outputs(2092) <= layer6_outputs(211);
    outputs(2093) <= not((layer6_outputs(2067)) or (layer6_outputs(3875)));
    outputs(2094) <= layer6_outputs(4633);
    outputs(2095) <= layer6_outputs(3491);
    outputs(2096) <= layer6_outputs(974);
    outputs(2097) <= not(layer6_outputs(5044));
    outputs(2098) <= not(layer6_outputs(4938));
    outputs(2099) <= not(layer6_outputs(3554));
    outputs(2100) <= not(layer6_outputs(3584));
    outputs(2101) <= (layer6_outputs(3918)) and not (layer6_outputs(779));
    outputs(2102) <= not(layer6_outputs(3401));
    outputs(2103) <= layer6_outputs(4243);
    outputs(2104) <= layer6_outputs(1740);
    outputs(2105) <= not(layer6_outputs(1265));
    outputs(2106) <= layer6_outputs(2740);
    outputs(2107) <= not(layer6_outputs(203));
    outputs(2108) <= (layer6_outputs(3436)) xor (layer6_outputs(4120));
    outputs(2109) <= not(layer6_outputs(2129));
    outputs(2110) <= not(layer6_outputs(964));
    outputs(2111) <= not(layer6_outputs(383));
    outputs(2112) <= not(layer6_outputs(3139));
    outputs(2113) <= (layer6_outputs(1371)) xor (layer6_outputs(1895));
    outputs(2114) <= not(layer6_outputs(4866));
    outputs(2115) <= layer6_outputs(20);
    outputs(2116) <= not(layer6_outputs(3829));
    outputs(2117) <= layer6_outputs(3555);
    outputs(2118) <= layer6_outputs(3715);
    outputs(2119) <= (layer6_outputs(4722)) and not (layer6_outputs(3742));
    outputs(2120) <= (layer6_outputs(4595)) xor (layer6_outputs(455));
    outputs(2121) <= layer6_outputs(3708);
    outputs(2122) <= not(layer6_outputs(4021));
    outputs(2123) <= not(layer6_outputs(1023));
    outputs(2124) <= not(layer6_outputs(3749));
    outputs(2125) <= layer6_outputs(1649);
    outputs(2126) <= not(layer6_outputs(2058));
    outputs(2127) <= not(layer6_outputs(4700));
    outputs(2128) <= (layer6_outputs(660)) xor (layer6_outputs(812));
    outputs(2129) <= layer6_outputs(2268);
    outputs(2130) <= not(layer6_outputs(276));
    outputs(2131) <= layer6_outputs(4428);
    outputs(2132) <= not(layer6_outputs(3123));
    outputs(2133) <= not((layer6_outputs(2485)) xor (layer6_outputs(3537)));
    outputs(2134) <= layer6_outputs(1000);
    outputs(2135) <= (layer6_outputs(1808)) xor (layer6_outputs(4521));
    outputs(2136) <= layer6_outputs(1852);
    outputs(2137) <= (layer6_outputs(2875)) xor (layer6_outputs(3295));
    outputs(2138) <= (layer6_outputs(3353)) xor (layer6_outputs(1249));
    outputs(2139) <= not(layer6_outputs(350));
    outputs(2140) <= (layer6_outputs(3692)) and (layer6_outputs(4860));
    outputs(2141) <= not(layer6_outputs(3789)) or (layer6_outputs(3608));
    outputs(2142) <= layer6_outputs(4873);
    outputs(2143) <= not(layer6_outputs(297));
    outputs(2144) <= layer6_outputs(2929);
    outputs(2145) <= not(layer6_outputs(684));
    outputs(2146) <= (layer6_outputs(593)) xor (layer6_outputs(4133));
    outputs(2147) <= not(layer6_outputs(420));
    outputs(2148) <= layer6_outputs(1665);
    outputs(2149) <= layer6_outputs(417);
    outputs(2150) <= not(layer6_outputs(4344));
    outputs(2151) <= layer6_outputs(4558);
    outputs(2152) <= (layer6_outputs(3623)) and not (layer6_outputs(807));
    outputs(2153) <= not(layer6_outputs(221));
    outputs(2154) <= not((layer6_outputs(407)) or (layer6_outputs(1306)));
    outputs(2155) <= layer6_outputs(3217);
    outputs(2156) <= not(layer6_outputs(3229)) or (layer6_outputs(1247));
    outputs(2157) <= not((layer6_outputs(36)) xor (layer6_outputs(3724)));
    outputs(2158) <= not(layer6_outputs(1562));
    outputs(2159) <= not(layer6_outputs(711));
    outputs(2160) <= not(layer6_outputs(4946));
    outputs(2161) <= (layer6_outputs(965)) xor (layer6_outputs(2043));
    outputs(2162) <= not(layer6_outputs(2285));
    outputs(2163) <= layer6_outputs(3563);
    outputs(2164) <= not(layer6_outputs(2079));
    outputs(2165) <= not(layer6_outputs(3625)) or (layer6_outputs(4789));
    outputs(2166) <= not((layer6_outputs(719)) or (layer6_outputs(3432)));
    outputs(2167) <= not(layer6_outputs(3062));
    outputs(2168) <= layer6_outputs(2007);
    outputs(2169) <= (layer6_outputs(1593)) or (layer6_outputs(4476));
    outputs(2170) <= layer6_outputs(2677);
    outputs(2171) <= not((layer6_outputs(4839)) xor (layer6_outputs(3866)));
    outputs(2172) <= not(layer6_outputs(767));
    outputs(2173) <= layer6_outputs(3236);
    outputs(2174) <= not(layer6_outputs(4829)) or (layer6_outputs(3684));
    outputs(2175) <= not((layer6_outputs(1844)) xor (layer6_outputs(519)));
    outputs(2176) <= not(layer6_outputs(5009));
    outputs(2177) <= layer6_outputs(340);
    outputs(2178) <= not(layer6_outputs(3470));
    outputs(2179) <= layer6_outputs(3455);
    outputs(2180) <= not(layer6_outputs(2973));
    outputs(2181) <= (layer6_outputs(980)) and (layer6_outputs(152));
    outputs(2182) <= not((layer6_outputs(1462)) or (layer6_outputs(1942)));
    outputs(2183) <= not(layer6_outputs(473));
    outputs(2184) <= not(layer6_outputs(4634));
    outputs(2185) <= not(layer6_outputs(3567)) or (layer6_outputs(449));
    outputs(2186) <= not(layer6_outputs(2413));
    outputs(2187) <= not(layer6_outputs(2385));
    outputs(2188) <= (layer6_outputs(5035)) and not (layer6_outputs(1992));
    outputs(2189) <= not(layer6_outputs(3401));
    outputs(2190) <= layer6_outputs(4067);
    outputs(2191) <= layer6_outputs(2789);
    outputs(2192) <= not(layer6_outputs(3859));
    outputs(2193) <= not(layer6_outputs(4626));
    outputs(2194) <= not(layer6_outputs(1907));
    outputs(2195) <= not((layer6_outputs(4306)) xor (layer6_outputs(418)));
    outputs(2196) <= not(layer6_outputs(480));
    outputs(2197) <= not(layer6_outputs(1191));
    outputs(2198) <= not((layer6_outputs(1260)) or (layer6_outputs(2733)));
    outputs(2199) <= layer6_outputs(578);
    outputs(2200) <= not((layer6_outputs(4064)) xor (layer6_outputs(1626)));
    outputs(2201) <= layer6_outputs(802);
    outputs(2202) <= layer6_outputs(1454);
    outputs(2203) <= layer6_outputs(248);
    outputs(2204) <= layer6_outputs(4827);
    outputs(2205) <= layer6_outputs(1551);
    outputs(2206) <= (layer6_outputs(853)) and not (layer6_outputs(1506));
    outputs(2207) <= (layer6_outputs(3697)) and not (layer6_outputs(758));
    outputs(2208) <= layer6_outputs(4771);
    outputs(2209) <= layer6_outputs(3540);
    outputs(2210) <= not((layer6_outputs(217)) xor (layer6_outputs(1078)));
    outputs(2211) <= not(layer6_outputs(359));
    outputs(2212) <= layer6_outputs(687);
    outputs(2213) <= not(layer6_outputs(4400));
    outputs(2214) <= (layer6_outputs(2001)) and (layer6_outputs(4978));
    outputs(2215) <= not(layer6_outputs(1720));
    outputs(2216) <= not(layer6_outputs(1409));
    outputs(2217) <= not(layer6_outputs(3499));
    outputs(2218) <= not(layer6_outputs(2767)) or (layer6_outputs(424));
    outputs(2219) <= not(layer6_outputs(4466));
    outputs(2220) <= layer6_outputs(659);
    outputs(2221) <= not(layer6_outputs(1193));
    outputs(2222) <= (layer6_outputs(300)) and not (layer6_outputs(1210));
    outputs(2223) <= layer6_outputs(1667);
    outputs(2224) <= layer6_outputs(4828);
    outputs(2225) <= not((layer6_outputs(5)) xor (layer6_outputs(1581)));
    outputs(2226) <= not(layer6_outputs(4324));
    outputs(2227) <= layer6_outputs(668);
    outputs(2228) <= (layer6_outputs(3856)) and not (layer6_outputs(3547));
    outputs(2229) <= layer6_outputs(4051);
    outputs(2230) <= layer6_outputs(2715);
    outputs(2231) <= not((layer6_outputs(849)) xor (layer6_outputs(1934)));
    outputs(2232) <= not(layer6_outputs(3284));
    outputs(2233) <= not(layer6_outputs(5044));
    outputs(2234) <= (layer6_outputs(2677)) xor (layer6_outputs(721));
    outputs(2235) <= layer6_outputs(2929);
    outputs(2236) <= (layer6_outputs(4961)) xor (layer6_outputs(1798));
    outputs(2237) <= layer6_outputs(5005);
    outputs(2238) <= not(layer6_outputs(939)) or (layer6_outputs(4330));
    outputs(2239) <= layer6_outputs(3461);
    outputs(2240) <= (layer6_outputs(3929)) xor (layer6_outputs(4415));
    outputs(2241) <= (layer6_outputs(4783)) xor (layer6_outputs(3365));
    outputs(2242) <= layer6_outputs(1925);
    outputs(2243) <= not((layer6_outputs(3488)) or (layer6_outputs(4370)));
    outputs(2244) <= layer6_outputs(1423);
    outputs(2245) <= not(layer6_outputs(5002));
    outputs(2246) <= (layer6_outputs(4717)) xor (layer6_outputs(1426));
    outputs(2247) <= (layer6_outputs(113)) and not (layer6_outputs(3422));
    outputs(2248) <= not(layer6_outputs(1219));
    outputs(2249) <= not((layer6_outputs(286)) or (layer6_outputs(4541)));
    outputs(2250) <= (layer6_outputs(2102)) or (layer6_outputs(2595));
    outputs(2251) <= not(layer6_outputs(3107));
    outputs(2252) <= layer6_outputs(1455);
    outputs(2253) <= not(layer6_outputs(2402));
    outputs(2254) <= (layer6_outputs(2797)) xor (layer6_outputs(4206));
    outputs(2255) <= not(layer6_outputs(4330));
    outputs(2256) <= not(layer6_outputs(3631));
    outputs(2257) <= layer6_outputs(4645);
    outputs(2258) <= layer6_outputs(4051);
    outputs(2259) <= layer6_outputs(2659);
    outputs(2260) <= not(layer6_outputs(4382));
    outputs(2261) <= not(layer6_outputs(528));
    outputs(2262) <= (layer6_outputs(934)) xor (layer6_outputs(4567));
    outputs(2263) <= not(layer6_outputs(1301));
    outputs(2264) <= not(layer6_outputs(692));
    outputs(2265) <= layer6_outputs(2536);
    outputs(2266) <= not(layer6_outputs(3369));
    outputs(2267) <= not(layer6_outputs(343));
    outputs(2268) <= not(layer6_outputs(2294));
    outputs(2269) <= not(layer6_outputs(3299));
    outputs(2270) <= not(layer6_outputs(3686));
    outputs(2271) <= layer6_outputs(2934);
    outputs(2272) <= not(layer6_outputs(1952));
    outputs(2273) <= layer6_outputs(1048);
    outputs(2274) <= not(layer6_outputs(4759));
    outputs(2275) <= not((layer6_outputs(2700)) xor (layer6_outputs(4747)));
    outputs(2276) <= layer6_outputs(1733);
    outputs(2277) <= layer6_outputs(2475);
    outputs(2278) <= not(layer6_outputs(3705));
    outputs(2279) <= layer6_outputs(2567);
    outputs(2280) <= not((layer6_outputs(398)) xor (layer6_outputs(482)));
    outputs(2281) <= (layer6_outputs(3302)) or (layer6_outputs(4915));
    outputs(2282) <= not(layer6_outputs(1697));
    outputs(2283) <= not((layer6_outputs(677)) and (layer6_outputs(2123)));
    outputs(2284) <= not(layer6_outputs(2298));
    outputs(2285) <= not(layer6_outputs(1468));
    outputs(2286) <= (layer6_outputs(4014)) xor (layer6_outputs(1215));
    outputs(2287) <= not(layer6_outputs(4221));
    outputs(2288) <= not((layer6_outputs(4184)) and (layer6_outputs(5082)));
    outputs(2289) <= layer6_outputs(2592);
    outputs(2290) <= not(layer6_outputs(2175));
    outputs(2291) <= layer6_outputs(2593);
    outputs(2292) <= not((layer6_outputs(3626)) or (layer6_outputs(476)));
    outputs(2293) <= layer6_outputs(5068);
    outputs(2294) <= not(layer6_outputs(2380));
    outputs(2295) <= layer6_outputs(1642);
    outputs(2296) <= layer6_outputs(2977);
    outputs(2297) <= not(layer6_outputs(1939));
    outputs(2298) <= not(layer6_outputs(154));
    outputs(2299) <= not(layer6_outputs(127));
    outputs(2300) <= layer6_outputs(3902);
    outputs(2301) <= (layer6_outputs(137)) and not (layer6_outputs(723));
    outputs(2302) <= not((layer6_outputs(2882)) xor (layer6_outputs(2500)));
    outputs(2303) <= layer6_outputs(1648);
    outputs(2304) <= not((layer6_outputs(689)) and (layer6_outputs(2089)));
    outputs(2305) <= layer6_outputs(1976);
    outputs(2306) <= not(layer6_outputs(1031));
    outputs(2307) <= not(layer6_outputs(4495));
    outputs(2308) <= layer6_outputs(3668);
    outputs(2309) <= not(layer6_outputs(3273));
    outputs(2310) <= not(layer6_outputs(44));
    outputs(2311) <= not(layer6_outputs(4237));
    outputs(2312) <= not(layer6_outputs(397));
    outputs(2313) <= not(layer6_outputs(4162));
    outputs(2314) <= layer6_outputs(4223);
    outputs(2315) <= layer6_outputs(3209);
    outputs(2316) <= not((layer6_outputs(987)) or (layer6_outputs(4452)));
    outputs(2317) <= layer6_outputs(2000);
    outputs(2318) <= not(layer6_outputs(3355)) or (layer6_outputs(3889));
    outputs(2319) <= (layer6_outputs(2491)) and not (layer6_outputs(4851));
    outputs(2320) <= not(layer6_outputs(4414));
    outputs(2321) <= not(layer6_outputs(1378));
    outputs(2322) <= not(layer6_outputs(4276));
    outputs(2323) <= layer6_outputs(4001);
    outputs(2324) <= not(layer6_outputs(2431));
    outputs(2325) <= layer6_outputs(4998);
    outputs(2326) <= layer6_outputs(850);
    outputs(2327) <= (layer6_outputs(2377)) xor (layer6_outputs(1556));
    outputs(2328) <= layer6_outputs(2295);
    outputs(2329) <= not(layer6_outputs(3924));
    outputs(2330) <= (layer6_outputs(2042)) or (layer6_outputs(1546));
    outputs(2331) <= (layer6_outputs(2112)) xor (layer6_outputs(5076));
    outputs(2332) <= not((layer6_outputs(3108)) xor (layer6_outputs(3071)));
    outputs(2333) <= not((layer6_outputs(3627)) xor (layer6_outputs(4677)));
    outputs(2334) <= not(layer6_outputs(2925));
    outputs(2335) <= layer6_outputs(4349);
    outputs(2336) <= not((layer6_outputs(2972)) xor (layer6_outputs(742)));
    outputs(2337) <= not(layer6_outputs(2524));
    outputs(2338) <= (layer6_outputs(5062)) xor (layer6_outputs(3466));
    outputs(2339) <= not(layer6_outputs(1093));
    outputs(2340) <= layer6_outputs(2344);
    outputs(2341) <= layer6_outputs(1842);
    outputs(2342) <= not(layer6_outputs(4218));
    outputs(2343) <= layer6_outputs(2586);
    outputs(2344) <= not(layer6_outputs(1243));
    outputs(2345) <= layer6_outputs(5106);
    outputs(2346) <= layer6_outputs(3993);
    outputs(2347) <= not(layer6_outputs(4952)) or (layer6_outputs(1555));
    outputs(2348) <= not(layer6_outputs(1933));
    outputs(2349) <= not(layer6_outputs(2334)) or (layer6_outputs(3648));
    outputs(2350) <= layer6_outputs(3251);
    outputs(2351) <= not(layer6_outputs(4984));
    outputs(2352) <= not(layer6_outputs(592));
    outputs(2353) <= not(layer6_outputs(4773));
    outputs(2354) <= layer6_outputs(3238);
    outputs(2355) <= not(layer6_outputs(1731));
    outputs(2356) <= not((layer6_outputs(1356)) xor (layer6_outputs(1417)));
    outputs(2357) <= layer6_outputs(3997);
    outputs(2358) <= not(layer6_outputs(3507));
    outputs(2359) <= not((layer6_outputs(2970)) or (layer6_outputs(3312)));
    outputs(2360) <= not(layer6_outputs(4927));
    outputs(2361) <= not(layer6_outputs(3163));
    outputs(2362) <= not(layer6_outputs(4812));
    outputs(2363) <= layer6_outputs(3103);
    outputs(2364) <= not((layer6_outputs(4235)) and (layer6_outputs(2970)));
    outputs(2365) <= (layer6_outputs(2492)) xor (layer6_outputs(277));
    outputs(2366) <= (layer6_outputs(3821)) xor (layer6_outputs(2407));
    outputs(2367) <= layer6_outputs(434);
    outputs(2368) <= (layer6_outputs(1313)) and not (layer6_outputs(3675));
    outputs(2369) <= layer6_outputs(1);
    outputs(2370) <= layer6_outputs(4236);
    outputs(2371) <= not(layer6_outputs(430));
    outputs(2372) <= not((layer6_outputs(819)) or (layer6_outputs(609)));
    outputs(2373) <= (layer6_outputs(3559)) xor (layer6_outputs(4749));
    outputs(2374) <= not((layer6_outputs(3418)) xor (layer6_outputs(1436)));
    outputs(2375) <= layer6_outputs(518);
    outputs(2376) <= not(layer6_outputs(615));
    outputs(2377) <= (layer6_outputs(2950)) or (layer6_outputs(4756));
    outputs(2378) <= not((layer6_outputs(2042)) xor (layer6_outputs(973)));
    outputs(2379) <= not((layer6_outputs(5034)) xor (layer6_outputs(4408)));
    outputs(2380) <= layer6_outputs(3648);
    outputs(2381) <= not(layer6_outputs(1376));
    outputs(2382) <= not(layer6_outputs(354));
    outputs(2383) <= not(layer6_outputs(2388));
    outputs(2384) <= layer6_outputs(4774);
    outputs(2385) <= layer6_outputs(2263);
    outputs(2386) <= not(layer6_outputs(2216));
    outputs(2387) <= (layer6_outputs(4334)) xor (layer6_outputs(519));
    outputs(2388) <= layer6_outputs(4935);
    outputs(2389) <= not((layer6_outputs(1823)) or (layer6_outputs(1996)));
    outputs(2390) <= layer6_outputs(24);
    outputs(2391) <= layer6_outputs(3360);
    outputs(2392) <= layer6_outputs(986);
    outputs(2393) <= not(layer6_outputs(1833));
    outputs(2394) <= not((layer6_outputs(292)) xor (layer6_outputs(2160)));
    outputs(2395) <= layer6_outputs(2217);
    outputs(2396) <= (layer6_outputs(3178)) and (layer6_outputs(4545));
    outputs(2397) <= not(layer6_outputs(2082));
    outputs(2398) <= layer6_outputs(4072);
    outputs(2399) <= not(layer6_outputs(3733));
    outputs(2400) <= (layer6_outputs(4018)) and not (layer6_outputs(4760));
    outputs(2401) <= not((layer6_outputs(131)) or (layer6_outputs(2065)));
    outputs(2402) <= not(layer6_outputs(2310)) or (layer6_outputs(3044));
    outputs(2403) <= not(layer6_outputs(1310));
    outputs(2404) <= not(layer6_outputs(3950));
    outputs(2405) <= not(layer6_outputs(3576)) or (layer6_outputs(4809));
    outputs(2406) <= layer6_outputs(3335);
    outputs(2407) <= not(layer6_outputs(3014));
    outputs(2408) <= (layer6_outputs(3170)) and (layer6_outputs(107));
    outputs(2409) <= not(layer6_outputs(4264));
    outputs(2410) <= not((layer6_outputs(3320)) xor (layer6_outputs(1555)));
    outputs(2411) <= not(layer6_outputs(1257));
    outputs(2412) <= not(layer6_outputs(3064));
    outputs(2413) <= not(layer6_outputs(999));
    outputs(2414) <= (layer6_outputs(1089)) xor (layer6_outputs(3116));
    outputs(2415) <= not(layer6_outputs(4983));
    outputs(2416) <= layer6_outputs(1845);
    outputs(2417) <= not(layer6_outputs(4444));
    outputs(2418) <= not((layer6_outputs(2492)) or (layer6_outputs(463)));
    outputs(2419) <= not(layer6_outputs(978));
    outputs(2420) <= not(layer6_outputs(1514));
    outputs(2421) <= layer6_outputs(4682);
    outputs(2422) <= layer6_outputs(1049);
    outputs(2423) <= layer6_outputs(1140);
    outputs(2424) <= layer6_outputs(318);
    outputs(2425) <= not(layer6_outputs(2699));
    outputs(2426) <= not((layer6_outputs(2993)) xor (layer6_outputs(3740)));
    outputs(2427) <= (layer6_outputs(446)) and not (layer6_outputs(4351));
    outputs(2428) <= not(layer6_outputs(4744));
    outputs(2429) <= not(layer6_outputs(3854));
    outputs(2430) <= layer6_outputs(1642);
    outputs(2431) <= layer6_outputs(844);
    outputs(2432) <= not(layer6_outputs(2109));
    outputs(2433) <= not(layer6_outputs(3246));
    outputs(2434) <= not((layer6_outputs(554)) xor (layer6_outputs(4411)));
    outputs(2435) <= layer6_outputs(1308);
    outputs(2436) <= not(layer6_outputs(4565));
    outputs(2437) <= not(layer6_outputs(1072));
    outputs(2438) <= (layer6_outputs(3549)) xor (layer6_outputs(3991));
    outputs(2439) <= (layer6_outputs(3951)) and (layer6_outputs(2511));
    outputs(2440) <= layer6_outputs(3680);
    outputs(2441) <= not(layer6_outputs(4295));
    outputs(2442) <= not(layer6_outputs(4298));
    outputs(2443) <= not(layer6_outputs(3825));
    outputs(2444) <= not((layer6_outputs(2783)) and (layer6_outputs(4721)));
    outputs(2445) <= not((layer6_outputs(891)) xor (layer6_outputs(4363)));
    outputs(2446) <= layer6_outputs(2499);
    outputs(2447) <= not(layer6_outputs(2914));
    outputs(2448) <= layer6_outputs(3834);
    outputs(2449) <= not(layer6_outputs(3008));
    outputs(2450) <= layer6_outputs(4726);
    outputs(2451) <= layer6_outputs(3197);
    outputs(2452) <= layer6_outputs(3988);
    outputs(2453) <= layer6_outputs(64);
    outputs(2454) <= layer6_outputs(4741);
    outputs(2455) <= layer6_outputs(1333);
    outputs(2456) <= layer6_outputs(3831);
    outputs(2457) <= not(layer6_outputs(4879));
    outputs(2458) <= layer6_outputs(3636);
    outputs(2459) <= layer6_outputs(4008);
    outputs(2460) <= not(layer6_outputs(270));
    outputs(2461) <= layer6_outputs(2218);
    outputs(2462) <= layer6_outputs(189);
    outputs(2463) <= not((layer6_outputs(536)) and (layer6_outputs(3237)));
    outputs(2464) <= layer6_outputs(3773);
    outputs(2465) <= not(layer6_outputs(1422));
    outputs(2466) <= (layer6_outputs(2072)) or (layer6_outputs(1991));
    outputs(2467) <= not(layer6_outputs(408)) or (layer6_outputs(2187));
    outputs(2468) <= layer6_outputs(4487);
    outputs(2469) <= layer6_outputs(4652);
    outputs(2470) <= not(layer6_outputs(4164));
    outputs(2471) <= layer6_outputs(613);
    outputs(2472) <= not(layer6_outputs(2395));
    outputs(2473) <= not(layer6_outputs(4066));
    outputs(2474) <= not(layer6_outputs(1559));
    outputs(2475) <= layer6_outputs(2059);
    outputs(2476) <= layer6_outputs(2005);
    outputs(2477) <= layer6_outputs(3217);
    outputs(2478) <= (layer6_outputs(3230)) and not (layer6_outputs(2034));
    outputs(2479) <= layer6_outputs(4772);
    outputs(2480) <= layer6_outputs(3907);
    outputs(2481) <= not(layer6_outputs(3578));
    outputs(2482) <= not(layer6_outputs(1444));
    outputs(2483) <= layer6_outputs(2442);
    outputs(2484) <= not(layer6_outputs(4181));
    outputs(2485) <= not((layer6_outputs(4291)) xor (layer6_outputs(1051)));
    outputs(2486) <= (layer6_outputs(4139)) xor (layer6_outputs(488));
    outputs(2487) <= layer6_outputs(2944);
    outputs(2488) <= (layer6_outputs(2410)) and not (layer6_outputs(2496));
    outputs(2489) <= not(layer6_outputs(663));
    outputs(2490) <= layer6_outputs(4560);
    outputs(2491) <= (layer6_outputs(998)) and (layer6_outputs(1972));
    outputs(2492) <= (layer6_outputs(1045)) and (layer6_outputs(4825));
    outputs(2493) <= not((layer6_outputs(3698)) and (layer6_outputs(3821)));
    outputs(2494) <= not(layer6_outputs(1217));
    outputs(2495) <= (layer6_outputs(3698)) and (layer6_outputs(4761));
    outputs(2496) <= not(layer6_outputs(2976));
    outputs(2497) <= layer6_outputs(759);
    outputs(2498) <= layer6_outputs(3750);
    outputs(2499) <= (layer6_outputs(2367)) and (layer6_outputs(899));
    outputs(2500) <= not((layer6_outputs(1250)) xor (layer6_outputs(2362)));
    outputs(2501) <= layer6_outputs(3737);
    outputs(2502) <= layer6_outputs(5033);
    outputs(2503) <= not(layer6_outputs(3525));
    outputs(2504) <= layer6_outputs(405);
    outputs(2505) <= not(layer6_outputs(654));
    outputs(2506) <= layer6_outputs(3176);
    outputs(2507) <= (layer6_outputs(2230)) and not (layer6_outputs(483));
    outputs(2508) <= layer6_outputs(3633);
    outputs(2509) <= (layer6_outputs(3565)) and (layer6_outputs(1835));
    outputs(2510) <= not((layer6_outputs(726)) xor (layer6_outputs(1346)));
    outputs(2511) <= (layer6_outputs(1297)) xor (layer6_outputs(3002));
    outputs(2512) <= layer6_outputs(1646);
    outputs(2513) <= layer6_outputs(250);
    outputs(2514) <= not(layer6_outputs(1684));
    outputs(2515) <= layer6_outputs(2183);
    outputs(2516) <= not(layer6_outputs(1820));
    outputs(2517) <= not(layer6_outputs(540));
    outputs(2518) <= not(layer6_outputs(944));
    outputs(2519) <= layer6_outputs(4821);
    outputs(2520) <= layer6_outputs(4166);
    outputs(2521) <= not(layer6_outputs(2709));
    outputs(2522) <= (layer6_outputs(3763)) or (layer6_outputs(3267));
    outputs(2523) <= layer6_outputs(11);
    outputs(2524) <= not(layer6_outputs(992));
    outputs(2525) <= not(layer6_outputs(1778));
    outputs(2526) <= layer6_outputs(537);
    outputs(2527) <= not(layer6_outputs(3721));
    outputs(2528) <= not((layer6_outputs(5000)) xor (layer6_outputs(1841)));
    outputs(2529) <= layer6_outputs(4578);
    outputs(2530) <= layer6_outputs(2224);
    outputs(2531) <= not((layer6_outputs(3699)) xor (layer6_outputs(1550)));
    outputs(2532) <= layer6_outputs(4689);
    outputs(2533) <= not(layer6_outputs(3117));
    outputs(2534) <= (layer6_outputs(4755)) and not (layer6_outputs(1093));
    outputs(2535) <= not(layer6_outputs(4061));
    outputs(2536) <= not(layer6_outputs(1910));
    outputs(2537) <= layer6_outputs(3235);
    outputs(2538) <= layer6_outputs(1495);
    outputs(2539) <= layer6_outputs(1604);
    outputs(2540) <= (layer6_outputs(5063)) xor (layer6_outputs(3213));
    outputs(2541) <= layer6_outputs(4855);
    outputs(2542) <= (layer6_outputs(733)) xor (layer6_outputs(4285));
    outputs(2543) <= not(layer6_outputs(799));
    outputs(2544) <= not(layer6_outputs(2481)) or (layer6_outputs(3285));
    outputs(2545) <= not(layer6_outputs(2576));
    outputs(2546) <= layer6_outputs(1045);
    outputs(2547) <= layer6_outputs(4360);
    outputs(2548) <= not(layer6_outputs(2896)) or (layer6_outputs(2915));
    outputs(2549) <= (layer6_outputs(3002)) xor (layer6_outputs(1012));
    outputs(2550) <= not(layer6_outputs(4556));
    outputs(2551) <= layer6_outputs(639);
    outputs(2552) <= not((layer6_outputs(3961)) xor (layer6_outputs(3621)));
    outputs(2553) <= (layer6_outputs(3958)) and (layer6_outputs(4253));
    outputs(2554) <= layer6_outputs(2237);
    outputs(2555) <= not(layer6_outputs(3221));
    outputs(2556) <= not(layer6_outputs(1213));
    outputs(2557) <= not(layer6_outputs(775));
    outputs(2558) <= layer6_outputs(4461);
    outputs(2559) <= not((layer6_outputs(2812)) and (layer6_outputs(4025)));
    outputs(2560) <= layer6_outputs(2051);
    outputs(2561) <= not((layer6_outputs(2520)) xor (layer6_outputs(1105)));
    outputs(2562) <= layer6_outputs(3634);
    outputs(2563) <= not(layer6_outputs(2786));
    outputs(2564) <= (layer6_outputs(652)) and not (layer6_outputs(5055));
    outputs(2565) <= not(layer6_outputs(2545));
    outputs(2566) <= not((layer6_outputs(2583)) xor (layer6_outputs(2679)));
    outputs(2567) <= not(layer6_outputs(3542));
    outputs(2568) <= layer6_outputs(2386);
    outputs(2569) <= layer6_outputs(2973);
    outputs(2570) <= layer6_outputs(2668);
    outputs(2571) <= not(layer6_outputs(2194));
    outputs(2572) <= (layer6_outputs(5075)) and (layer6_outputs(2452));
    outputs(2573) <= not((layer6_outputs(1038)) and (layer6_outputs(2986)));
    outputs(2574) <= not((layer6_outputs(4848)) and (layer6_outputs(561)));
    outputs(2575) <= (layer6_outputs(856)) xor (layer6_outputs(2555));
    outputs(2576) <= layer6_outputs(4611);
    outputs(2577) <= layer6_outputs(1130);
    outputs(2578) <= not((layer6_outputs(2115)) xor (layer6_outputs(3374)));
    outputs(2579) <= layer6_outputs(1729);
    outputs(2580) <= not((layer6_outputs(226)) xor (layer6_outputs(1686)));
    outputs(2581) <= layer6_outputs(1329);
    outputs(2582) <= not(layer6_outputs(3193));
    outputs(2583) <= layer6_outputs(1584);
    outputs(2584) <= layer6_outputs(4436);
    outputs(2585) <= not(layer6_outputs(4354));
    outputs(2586) <= (layer6_outputs(5035)) xor (layer6_outputs(418));
    outputs(2587) <= not((layer6_outputs(1868)) xor (layer6_outputs(2046)));
    outputs(2588) <= not(layer6_outputs(3165)) or (layer6_outputs(3946));
    outputs(2589) <= layer6_outputs(4155);
    outputs(2590) <= not(layer6_outputs(425));
    outputs(2591) <= not(layer6_outputs(4423));
    outputs(2592) <= (layer6_outputs(4718)) and not (layer6_outputs(3509));
    outputs(2593) <= layer6_outputs(2899);
    outputs(2594) <= layer6_outputs(1669);
    outputs(2595) <= not(layer6_outputs(2344));
    outputs(2596) <= layer6_outputs(2569);
    outputs(2597) <= layer6_outputs(3044);
    outputs(2598) <= not(layer6_outputs(3780));
    outputs(2599) <= layer6_outputs(3115);
    outputs(2600) <= not(layer6_outputs(2063));
    outputs(2601) <= not(layer6_outputs(3947));
    outputs(2602) <= not(layer6_outputs(982));
    outputs(2603) <= not(layer6_outputs(1318));
    outputs(2604) <= not(layer6_outputs(2372));
    outputs(2605) <= not(layer6_outputs(322));
    outputs(2606) <= layer6_outputs(4060);
    outputs(2607) <= layer6_outputs(2330);
    outputs(2608) <= layer6_outputs(884);
    outputs(2609) <= (layer6_outputs(1080)) xor (layer6_outputs(1242));
    outputs(2610) <= layer6_outputs(2269);
    outputs(2611) <= layer6_outputs(1132);
    outputs(2612) <= not(layer6_outputs(2215));
    outputs(2613) <= not(layer6_outputs(2375)) or (layer6_outputs(530));
    outputs(2614) <= (layer6_outputs(946)) xor (layer6_outputs(4035));
    outputs(2615) <= layer6_outputs(2551);
    outputs(2616) <= layer6_outputs(2634);
    outputs(2617) <= layer6_outputs(5071);
    outputs(2618) <= layer6_outputs(1053);
    outputs(2619) <= (layer6_outputs(3514)) xor (layer6_outputs(4283));
    outputs(2620) <= layer6_outputs(3301);
    outputs(2621) <= (layer6_outputs(646)) xor (layer6_outputs(3048));
    outputs(2622) <= (layer6_outputs(4006)) xor (layer6_outputs(3873));
    outputs(2623) <= layer6_outputs(1003);
    outputs(2624) <= layer6_outputs(1450);
    outputs(2625) <= not(layer6_outputs(4215));
    outputs(2626) <= not(layer6_outputs(454));
    outputs(2627) <= layer6_outputs(4949);
    outputs(2628) <= not(layer6_outputs(2341));
    outputs(2629) <= not((layer6_outputs(3568)) xor (layer6_outputs(301)));
    outputs(2630) <= not(layer6_outputs(5049));
    outputs(2631) <= not(layer6_outputs(4290));
    outputs(2632) <= not(layer6_outputs(4091));
    outputs(2633) <= not(layer6_outputs(460));
    outputs(2634) <= layer6_outputs(2597);
    outputs(2635) <= not(layer6_outputs(1964));
    outputs(2636) <= layer6_outputs(3629);
    outputs(2637) <= not(layer6_outputs(2479));
    outputs(2638) <= layer6_outputs(2480);
    outputs(2639) <= layer6_outputs(3173);
    outputs(2640) <= not((layer6_outputs(4692)) xor (layer6_outputs(1312)));
    outputs(2641) <= layer6_outputs(3041);
    outputs(2642) <= layer6_outputs(4049);
    outputs(2643) <= not(layer6_outputs(3272));
    outputs(2644) <= not((layer6_outputs(1437)) or (layer6_outputs(4034)));
    outputs(2645) <= not(layer6_outputs(2747)) or (layer6_outputs(4039));
    outputs(2646) <= not((layer6_outputs(1773)) xor (layer6_outputs(640)));
    outputs(2647) <= not((layer6_outputs(2069)) xor (layer6_outputs(2023)));
    outputs(2648) <= not(layer6_outputs(3269));
    outputs(2649) <= (layer6_outputs(1104)) xor (layer6_outputs(3537));
    outputs(2650) <= not(layer6_outputs(942));
    outputs(2651) <= layer6_outputs(2304);
    outputs(2652) <= (layer6_outputs(2296)) or (layer6_outputs(1271));
    outputs(2653) <= not(layer6_outputs(3997));
    outputs(2654) <= not((layer6_outputs(1948)) or (layer6_outputs(2278)));
    outputs(2655) <= not(layer6_outputs(1159)) or (layer6_outputs(1154));
    outputs(2656) <= layer6_outputs(4082);
    outputs(2657) <= layer6_outputs(3304);
    outputs(2658) <= (layer6_outputs(5)) xor (layer6_outputs(3429));
    outputs(2659) <= layer6_outputs(3145);
    outputs(2660) <= (layer6_outputs(690)) and not (layer6_outputs(1192));
    outputs(2661) <= (layer6_outputs(4175)) and (layer6_outputs(3562));
    outputs(2662) <= not(layer6_outputs(2076));
    outputs(2663) <= not((layer6_outputs(2338)) xor (layer6_outputs(1991)));
    outputs(2664) <= (layer6_outputs(1402)) xor (layer6_outputs(3321));
    outputs(2665) <= not(layer6_outputs(3392));
    outputs(2666) <= not((layer6_outputs(3581)) xor (layer6_outputs(1563)));
    outputs(2667) <= not(layer6_outputs(1438));
    outputs(2668) <= not(layer6_outputs(52));
    outputs(2669) <= layer6_outputs(4540);
    outputs(2670) <= layer6_outputs(3679);
    outputs(2671) <= not(layer6_outputs(3822));
    outputs(2672) <= (layer6_outputs(3366)) xor (layer6_outputs(1995));
    outputs(2673) <= (layer6_outputs(720)) and not (layer6_outputs(4770));
    outputs(2674) <= not(layer6_outputs(1207));
    outputs(2675) <= (layer6_outputs(1532)) or (layer6_outputs(116));
    outputs(2676) <= (layer6_outputs(1142)) xor (layer6_outputs(4161));
    outputs(2677) <= (layer6_outputs(4585)) or (layer6_outputs(2631));
    outputs(2678) <= not(layer6_outputs(1095));
    outputs(2679) <= layer6_outputs(2662);
    outputs(2680) <= not((layer6_outputs(2916)) or (layer6_outputs(2268)));
    outputs(2681) <= (layer6_outputs(3509)) xor (layer6_outputs(2531));
    outputs(2682) <= not(layer6_outputs(1912));
    outputs(2683) <= not((layer6_outputs(512)) xor (layer6_outputs(509)));
    outputs(2684) <= layer6_outputs(2327);
    outputs(2685) <= layer6_outputs(1996);
    outputs(2686) <= layer6_outputs(1031);
    outputs(2687) <= not(layer6_outputs(2290)) or (layer6_outputs(83));
    outputs(2688) <= layer6_outputs(4635);
    outputs(2689) <= not((layer6_outputs(4300)) xor (layer6_outputs(4675)));
    outputs(2690) <= layer6_outputs(2618);
    outputs(2691) <= not(layer6_outputs(4075));
    outputs(2692) <= (layer6_outputs(1823)) and (layer6_outputs(359));
    outputs(2693) <= not((layer6_outputs(5065)) xor (layer6_outputs(921)));
    outputs(2694) <= layer6_outputs(1366);
    outputs(2695) <= layer6_outputs(4110);
    outputs(2696) <= not(layer6_outputs(188));
    outputs(2697) <= layer6_outputs(2064);
    outputs(2698) <= not((layer6_outputs(632)) xor (layer6_outputs(484)));
    outputs(2699) <= not(layer6_outputs(2545));
    outputs(2700) <= not((layer6_outputs(2124)) xor (layer6_outputs(3019)));
    outputs(2701) <= layer6_outputs(4243);
    outputs(2702) <= (layer6_outputs(1827)) xor (layer6_outputs(1987));
    outputs(2703) <= (layer6_outputs(2790)) and not (layer6_outputs(1367));
    outputs(2704) <= not(layer6_outputs(4394));
    outputs(2705) <= not((layer6_outputs(3084)) xor (layer6_outputs(341)));
    outputs(2706) <= layer6_outputs(3273);
    outputs(2707) <= layer6_outputs(3765);
    outputs(2708) <= layer6_outputs(1717);
    outputs(2709) <= not(layer6_outputs(1314));
    outputs(2710) <= layer6_outputs(936);
    outputs(2711) <= not(layer6_outputs(799));
    outputs(2712) <= not((layer6_outputs(2156)) and (layer6_outputs(3142)));
    outputs(2713) <= (layer6_outputs(2706)) and not (layer6_outputs(3910));
    outputs(2714) <= not(layer6_outputs(715));
    outputs(2715) <= not(layer6_outputs(2451));
    outputs(2716) <= layer6_outputs(2018);
    outputs(2717) <= (layer6_outputs(2596)) xor (layer6_outputs(4207));
    outputs(2718) <= layer6_outputs(2660);
    outputs(2719) <= (layer6_outputs(337)) xor (layer6_outputs(225));
    outputs(2720) <= layer6_outputs(131);
    outputs(2721) <= not(layer6_outputs(1617));
    outputs(2722) <= not((layer6_outputs(3982)) xor (layer6_outputs(1782)));
    outputs(2723) <= layer6_outputs(3221);
    outputs(2724) <= not(layer6_outputs(5108));
    outputs(2725) <= not(layer6_outputs(82));
    outputs(2726) <= layer6_outputs(3481);
    outputs(2727) <= not(layer6_outputs(3267));
    outputs(2728) <= (layer6_outputs(2538)) xor (layer6_outputs(3848));
    outputs(2729) <= layer6_outputs(711);
    outputs(2730) <= (layer6_outputs(809)) and (layer6_outputs(8));
    outputs(2731) <= (layer6_outputs(1312)) xor (layer6_outputs(3669));
    outputs(2732) <= not(layer6_outputs(1267));
    outputs(2733) <= not(layer6_outputs(4285)) or (layer6_outputs(866));
    outputs(2734) <= layer6_outputs(3530);
    outputs(2735) <= (layer6_outputs(3676)) and not (layer6_outputs(1735));
    outputs(2736) <= not(layer6_outputs(3390));
    outputs(2737) <= layer6_outputs(1595);
    outputs(2738) <= not(layer6_outputs(2754));
    outputs(2739) <= not(layer6_outputs(1861));
    outputs(2740) <= not((layer6_outputs(4141)) and (layer6_outputs(4046)));
    outputs(2741) <= layer6_outputs(2482);
    outputs(2742) <= layer6_outputs(4950);
    outputs(2743) <= layer6_outputs(1160);
    outputs(2744) <= not((layer6_outputs(2259)) and (layer6_outputs(576)));
    outputs(2745) <= not((layer6_outputs(2430)) xor (layer6_outputs(3990)));
    outputs(2746) <= (layer6_outputs(3696)) xor (layer6_outputs(2185));
    outputs(2747) <= (layer6_outputs(2654)) xor (layer6_outputs(5092));
    outputs(2748) <= not(layer6_outputs(2623));
    outputs(2749) <= not(layer6_outputs(4471));
    outputs(2750) <= not(layer6_outputs(4738));
    outputs(2751) <= (layer6_outputs(3039)) xor (layer6_outputs(1582));
    outputs(2752) <= not(layer6_outputs(3490));
    outputs(2753) <= (layer6_outputs(3645)) xor (layer6_outputs(3007));
    outputs(2754) <= not(layer6_outputs(1886));
    outputs(2755) <= not((layer6_outputs(3456)) xor (layer6_outputs(382)));
    outputs(2756) <= layer6_outputs(3095);
    outputs(2757) <= not(layer6_outputs(333));
    outputs(2758) <= not(layer6_outputs(2809));
    outputs(2759) <= not(layer6_outputs(1625));
    outputs(2760) <= layer6_outputs(1535);
    outputs(2761) <= layer6_outputs(3574);
    outputs(2762) <= not(layer6_outputs(3415)) or (layer6_outputs(4048));
    outputs(2763) <= not(layer6_outputs(4468));
    outputs(2764) <= not(layer6_outputs(2399));
    outputs(2765) <= (layer6_outputs(3845)) and not (layer6_outputs(811));
    outputs(2766) <= not(layer6_outputs(2163));
    outputs(2767) <= layer6_outputs(3544);
    outputs(2768) <= (layer6_outputs(4420)) or (layer6_outputs(2169));
    outputs(2769) <= (layer6_outputs(4665)) xor (layer6_outputs(4415));
    outputs(2770) <= (layer6_outputs(717)) xor (layer6_outputs(3526));
    outputs(2771) <= (layer6_outputs(3943)) and (layer6_outputs(3830));
    outputs(2772) <= not((layer6_outputs(1755)) xor (layer6_outputs(2592)));
    outputs(2773) <= not(layer6_outputs(838));
    outputs(2774) <= not(layer6_outputs(1637));
    outputs(2775) <= layer6_outputs(2513);
    outputs(2776) <= (layer6_outputs(3806)) or (layer6_outputs(1073));
    outputs(2777) <= layer6_outputs(2490);
    outputs(2778) <= not(layer6_outputs(479));
    outputs(2779) <= not(layer6_outputs(3227)) or (layer6_outputs(2165));
    outputs(2780) <= (layer6_outputs(2842)) xor (layer6_outputs(4072));
    outputs(2781) <= (layer6_outputs(2757)) xor (layer6_outputs(487));
    outputs(2782) <= layer6_outputs(5101);
    outputs(2783) <= not(layer6_outputs(1443));
    outputs(2784) <= not(layer6_outputs(993));
    outputs(2785) <= (layer6_outputs(752)) or (layer6_outputs(4786));
    outputs(2786) <= (layer6_outputs(1395)) xor (layer6_outputs(2127));
    outputs(2787) <= (layer6_outputs(4708)) xor (layer6_outputs(1790));
    outputs(2788) <= layer6_outputs(3053);
    outputs(2789) <= (layer6_outputs(700)) xor (layer6_outputs(457));
    outputs(2790) <= not((layer6_outputs(2754)) or (layer6_outputs(2493)));
    outputs(2791) <= layer6_outputs(4251);
    outputs(2792) <= layer6_outputs(2180);
    outputs(2793) <= not(layer6_outputs(928));
    outputs(2794) <= not(layer6_outputs(3589));
    outputs(2795) <= not((layer6_outputs(2913)) and (layer6_outputs(4170)));
    outputs(2796) <= not(layer6_outputs(3193));
    outputs(2797) <= not(layer6_outputs(3941));
    outputs(2798) <= not(layer6_outputs(852));
    outputs(2799) <= (layer6_outputs(1596)) xor (layer6_outputs(4231));
    outputs(2800) <= (layer6_outputs(1640)) xor (layer6_outputs(4505));
    outputs(2801) <= not(layer6_outputs(1337));
    outputs(2802) <= (layer6_outputs(4506)) xor (layer6_outputs(4672));
    outputs(2803) <= not((layer6_outputs(937)) xor (layer6_outputs(4780)));
    outputs(2804) <= layer6_outputs(3247);
    outputs(2805) <= layer6_outputs(4706);
    outputs(2806) <= layer6_outputs(3315);
    outputs(2807) <= not((layer6_outputs(3101)) xor (layer6_outputs(332)));
    outputs(2808) <= layer6_outputs(4322);
    outputs(2809) <= not(layer6_outputs(3890));
    outputs(2810) <= '1';
    outputs(2811) <= not(layer6_outputs(1406));
    outputs(2812) <= not(layer6_outputs(920));
    outputs(2813) <= not((layer6_outputs(4092)) xor (layer6_outputs(2498)));
    outputs(2814) <= not((layer6_outputs(327)) xor (layer6_outputs(38)));
    outputs(2815) <= not((layer6_outputs(2714)) xor (layer6_outputs(2081)));
    outputs(2816) <= not((layer6_outputs(605)) xor (layer6_outputs(3410)));
    outputs(2817) <= not(layer6_outputs(833));
    outputs(2818) <= not(layer6_outputs(4339));
    outputs(2819) <= layer6_outputs(4060);
    outputs(2820) <= not(layer6_outputs(525));
    outputs(2821) <= (layer6_outputs(3379)) xor (layer6_outputs(1163));
    outputs(2822) <= (layer6_outputs(4413)) xor (layer6_outputs(2141));
    outputs(2823) <= (layer6_outputs(3336)) xor (layer6_outputs(1225));
    outputs(2824) <= layer6_outputs(184);
    outputs(2825) <= layer6_outputs(3405);
    outputs(2826) <= not(layer6_outputs(169));
    outputs(2827) <= not(layer6_outputs(2126));
    outputs(2828) <= not(layer6_outputs(456));
    outputs(2829) <= (layer6_outputs(634)) xor (layer6_outputs(1226));
    outputs(2830) <= layer6_outputs(5046);
    outputs(2831) <= not(layer6_outputs(4209));
    outputs(2832) <= not(layer6_outputs(4392));
    outputs(2833) <= (layer6_outputs(2680)) or (layer6_outputs(562));
    outputs(2834) <= (layer6_outputs(3243)) and not (layer6_outputs(348));
    outputs(2835) <= not(layer6_outputs(3342));
    outputs(2836) <= (layer6_outputs(3468)) xor (layer6_outputs(1063));
    outputs(2837) <= (layer6_outputs(326)) xor (layer6_outputs(3468));
    outputs(2838) <= not(layer6_outputs(2987));
    outputs(2839) <= not((layer6_outputs(4602)) xor (layer6_outputs(58)));
    outputs(2840) <= (layer6_outputs(5009)) and not (layer6_outputs(156));
    outputs(2841) <= not(layer6_outputs(2094)) or (layer6_outputs(3860));
    outputs(2842) <= not(layer6_outputs(3356));
    outputs(2843) <= not(layer6_outputs(3239));
    outputs(2844) <= layer6_outputs(2021);
    outputs(2845) <= layer6_outputs(2825);
    outputs(2846) <= not(layer6_outputs(2643));
    outputs(2847) <= (layer6_outputs(207)) xor (layer6_outputs(358));
    outputs(2848) <= not(layer6_outputs(1768));
    outputs(2849) <= not((layer6_outputs(650)) xor (layer6_outputs(1135)));
    outputs(2850) <= layer6_outputs(3594);
    outputs(2851) <= not(layer6_outputs(4670));
    outputs(2852) <= layer6_outputs(4519);
    outputs(2853) <= (layer6_outputs(1854)) and (layer6_outputs(2783));
    outputs(2854) <= not(layer6_outputs(2529)) or (layer6_outputs(3367));
    outputs(2855) <= not(layer6_outputs(1269));
    outputs(2856) <= not(layer6_outputs(1430));
    outputs(2857) <= not((layer6_outputs(3717)) xor (layer6_outputs(4205)));
    outputs(2858) <= layer6_outputs(4847);
    outputs(2859) <= not(layer6_outputs(3259));
    outputs(2860) <= layer6_outputs(2255);
    outputs(2861) <= layer6_outputs(534);
    outputs(2862) <= layer6_outputs(1190);
    outputs(2863) <= not(layer6_outputs(4001));
    outputs(2864) <= layer6_outputs(2951);
    outputs(2865) <= not(layer6_outputs(4195));
    outputs(2866) <= not((layer6_outputs(1858)) xor (layer6_outputs(2118)));
    outputs(2867) <= (layer6_outputs(833)) xor (layer6_outputs(4052));
    outputs(2868) <= not(layer6_outputs(808));
    outputs(2869) <= (layer6_outputs(3599)) and not (layer6_outputs(4143));
    outputs(2870) <= layer6_outputs(2772);
    outputs(2871) <= (layer6_outputs(981)) xor (layer6_outputs(3225));
    outputs(2872) <= not(layer6_outputs(699));
    outputs(2873) <= not(layer6_outputs(2238));
    outputs(2874) <= layer6_outputs(3400);
    outputs(2875) <= not(layer6_outputs(3616));
    outputs(2876) <= not(layer6_outputs(4287));
    outputs(2877) <= not(layer6_outputs(1768));
    outputs(2878) <= not(layer6_outputs(254));
    outputs(2879) <= layer6_outputs(5037);
    outputs(2880) <= layer6_outputs(4073);
    outputs(2881) <= not(layer6_outputs(1268));
    outputs(2882) <= not(layer6_outputs(3222));
    outputs(2883) <= layer6_outputs(1507);
    outputs(2884) <= not(layer6_outputs(4799));
    outputs(2885) <= not(layer6_outputs(3862));
    outputs(2886) <= layer6_outputs(3577);
    outputs(2887) <= layer6_outputs(2689);
    outputs(2888) <= not((layer6_outputs(2021)) xor (layer6_outputs(3690)));
    outputs(2889) <= layer6_outputs(744);
    outputs(2890) <= layer6_outputs(4173);
    outputs(2891) <= not(layer6_outputs(2088));
    outputs(2892) <= not(layer6_outputs(2070));
    outputs(2893) <= not((layer6_outputs(2243)) or (layer6_outputs(2259)));
    outputs(2894) <= (layer6_outputs(3505)) and not (layer6_outputs(624));
    outputs(2895) <= layer6_outputs(1373);
    outputs(2896) <= layer6_outputs(3127);
    outputs(2897) <= not(layer6_outputs(4391));
    outputs(2898) <= (layer6_outputs(4726)) or (layer6_outputs(1821));
    outputs(2899) <= layer6_outputs(498);
    outputs(2900) <= (layer6_outputs(2596)) and (layer6_outputs(3218));
    outputs(2901) <= not((layer6_outputs(4730)) xor (layer6_outputs(1296)));
    outputs(2902) <= not(layer6_outputs(1753));
    outputs(2903) <= layer6_outputs(1672);
    outputs(2904) <= not((layer6_outputs(4325)) or (layer6_outputs(4924)));
    outputs(2905) <= not(layer6_outputs(57));
    outputs(2906) <= (layer6_outputs(3344)) or (layer6_outputs(2671));
    outputs(2907) <= not((layer6_outputs(1077)) xor (layer6_outputs(275)));
    outputs(2908) <= layer6_outputs(240);
    outputs(2909) <= (layer6_outputs(2925)) xor (layer6_outputs(344));
    outputs(2910) <= not(layer6_outputs(687));
    outputs(2911) <= not(layer6_outputs(3728));
    outputs(2912) <= not((layer6_outputs(2324)) xor (layer6_outputs(1195)));
    outputs(2913) <= layer6_outputs(1541);
    outputs(2914) <= layer6_outputs(1203);
    outputs(2915) <= (layer6_outputs(3601)) xor (layer6_outputs(3310));
    outputs(2916) <= layer6_outputs(620);
    outputs(2917) <= (layer6_outputs(1310)) and not (layer6_outputs(4996));
    outputs(2918) <= not(layer6_outputs(1474));
    outputs(2919) <= not(layer6_outputs(626));
    outputs(2920) <= (layer6_outputs(1135)) xor (layer6_outputs(407));
    outputs(2921) <= not(layer6_outputs(138));
    outputs(2922) <= (layer6_outputs(133)) xor (layer6_outputs(4745));
    outputs(2923) <= not(layer6_outputs(4810));
    outputs(2924) <= not(layer6_outputs(2066));
    outputs(2925) <= layer6_outputs(4458);
    outputs(2926) <= not(layer6_outputs(3058));
    outputs(2927) <= (layer6_outputs(3575)) xor (layer6_outputs(1882));
    outputs(2928) <= (layer6_outputs(2535)) xor (layer6_outputs(4668));
    outputs(2929) <= not((layer6_outputs(2485)) xor (layer6_outputs(1533)));
    outputs(2930) <= (layer6_outputs(4171)) xor (layer6_outputs(1464));
    outputs(2931) <= layer6_outputs(4);
    outputs(2932) <= not(layer6_outputs(4784));
    outputs(2933) <= layer6_outputs(3655);
    outputs(2934) <= layer6_outputs(2162);
    outputs(2935) <= layer6_outputs(569);
    outputs(2936) <= not(layer6_outputs(86));
    outputs(2937) <= layer6_outputs(1442);
    outputs(2938) <= not((layer6_outputs(924)) xor (layer6_outputs(496)));
    outputs(2939) <= not(layer6_outputs(3266));
    outputs(2940) <= layer6_outputs(1680);
    outputs(2941) <= (layer6_outputs(620)) and not (layer6_outputs(4533));
    outputs(2942) <= not(layer6_outputs(1443));
    outputs(2943) <= not(layer6_outputs(4090));
    outputs(2944) <= layer6_outputs(4785);
    outputs(2945) <= layer6_outputs(2885);
    outputs(2946) <= layer6_outputs(4032);
    outputs(2947) <= not(layer6_outputs(1145));
    outputs(2948) <= not(layer6_outputs(514));
    outputs(2949) <= layer6_outputs(3117);
    outputs(2950) <= layer6_outputs(2406);
    outputs(2951) <= not(layer6_outputs(3935)) or (layer6_outputs(1336));
    outputs(2952) <= not(layer6_outputs(3240));
    outputs(2953) <= not(layer6_outputs(4943));
    outputs(2954) <= not(layer6_outputs(4425));
    outputs(2955) <= layer6_outputs(4840);
    outputs(2956) <= not(layer6_outputs(3869));
    outputs(2957) <= not(layer6_outputs(474)) or (layer6_outputs(288));
    outputs(2958) <= not(layer6_outputs(2815)) or (layer6_outputs(2574));
    outputs(2959) <= not(layer6_outputs(4887));
    outputs(2960) <= not(layer6_outputs(1062)) or (layer6_outputs(650));
    outputs(2961) <= not(layer6_outputs(1942));
    outputs(2962) <= layer6_outputs(1828);
    outputs(2963) <= not(layer6_outputs(4488));
    outputs(2964) <= layer6_outputs(4031);
    outputs(2965) <= layer6_outputs(3304);
    outputs(2966) <= (layer6_outputs(1791)) and not (layer6_outputs(4610));
    outputs(2967) <= layer6_outputs(146);
    outputs(2968) <= (layer6_outputs(1138)) xor (layer6_outputs(229));
    outputs(2969) <= layer6_outputs(4875);
    outputs(2970) <= not((layer6_outputs(4004)) xor (layer6_outputs(990)));
    outputs(2971) <= not(layer6_outputs(3869));
    outputs(2972) <= not(layer6_outputs(4627));
    outputs(2973) <= not(layer6_outputs(4459)) or (layer6_outputs(3372));
    outputs(2974) <= (layer6_outputs(2915)) xor (layer6_outputs(3489));
    outputs(2975) <= not(layer6_outputs(2137));
    outputs(2976) <= (layer6_outputs(3580)) and (layer6_outputs(1124));
    outputs(2977) <= (layer6_outputs(311)) xor (layer6_outputs(1705));
    outputs(2978) <= not((layer6_outputs(1222)) xor (layer6_outputs(4267)));
    outputs(2979) <= not((layer6_outputs(4488)) xor (layer6_outputs(4126)));
    outputs(2980) <= layer6_outputs(4844);
    outputs(2981) <= not(layer6_outputs(1971)) or (layer6_outputs(4965));
    outputs(2982) <= layer6_outputs(4176);
    outputs(2983) <= not(layer6_outputs(281)) or (layer6_outputs(65));
    outputs(2984) <= not(layer6_outputs(2028));
    outputs(2985) <= not(layer6_outputs(1491)) or (layer6_outputs(3895));
    outputs(2986) <= not((layer6_outputs(4414)) xor (layer6_outputs(4787)));
    outputs(2987) <= not(layer6_outputs(3908));
    outputs(2988) <= not(layer6_outputs(1646));
    outputs(2989) <= not((layer6_outputs(1400)) xor (layer6_outputs(140)));
    outputs(2990) <= layer6_outputs(4332);
    outputs(2991) <= not(layer6_outputs(1693));
    outputs(2992) <= layer6_outputs(1113);
    outputs(2993) <= not(layer6_outputs(3416));
    outputs(2994) <= not(layer6_outputs(3042));
    outputs(2995) <= layer6_outputs(4754);
    outputs(2996) <= (layer6_outputs(3173)) or (layer6_outputs(3904));
    outputs(2997) <= layer6_outputs(2589);
    outputs(2998) <= not((layer6_outputs(1606)) and (layer6_outputs(3076)));
    outputs(2999) <= layer6_outputs(1553);
    outputs(3000) <= layer6_outputs(186);
    outputs(3001) <= not(layer6_outputs(1660));
    outputs(3002) <= layer6_outputs(2544);
    outputs(3003) <= (layer6_outputs(951)) xor (layer6_outputs(2063));
    outputs(3004) <= not(layer6_outputs(877));
    outputs(3005) <= not(layer6_outputs(1958));
    outputs(3006) <= not((layer6_outputs(3011)) xor (layer6_outputs(1627)));
    outputs(3007) <= layer6_outputs(747);
    outputs(3008) <= not((layer6_outputs(1930)) xor (layer6_outputs(903)));
    outputs(3009) <= layer6_outputs(3130);
    outputs(3010) <= not(layer6_outputs(3371));
    outputs(3011) <= not((layer6_outputs(1523)) xor (layer6_outputs(3927)));
    outputs(3012) <= layer6_outputs(4859);
    outputs(3013) <= not(layer6_outputs(720)) or (layer6_outputs(969));
    outputs(3014) <= not((layer6_outputs(2544)) xor (layer6_outputs(3564)));
    outputs(3015) <= (layer6_outputs(3404)) or (layer6_outputs(1166));
    outputs(3016) <= layer6_outputs(656);
    outputs(3017) <= not(layer6_outputs(3195));
    outputs(3018) <= not((layer6_outputs(1298)) xor (layer6_outputs(2374)));
    outputs(3019) <= layer6_outputs(3603);
    outputs(3020) <= layer6_outputs(2618);
    outputs(3021) <= not((layer6_outputs(1188)) xor (layer6_outputs(4987)));
    outputs(3022) <= not((layer6_outputs(3189)) xor (layer6_outputs(3297)));
    outputs(3023) <= not(layer6_outputs(1947));
    outputs(3024) <= not((layer6_outputs(2475)) or (layer6_outputs(3245)));
    outputs(3025) <= layer6_outputs(4902);
    outputs(3026) <= (layer6_outputs(53)) xor (layer6_outputs(2328));
    outputs(3027) <= layer6_outputs(167);
    outputs(3028) <= not(layer6_outputs(3857));
    outputs(3029) <= not(layer6_outputs(2140));
    outputs(3030) <= not(layer6_outputs(4648)) or (layer6_outputs(0));
    outputs(3031) <= not(layer6_outputs(958));
    outputs(3032) <= not(layer6_outputs(3263));
    outputs(3033) <= layer6_outputs(2373);
    outputs(3034) <= (layer6_outputs(2027)) xor (layer6_outputs(3188));
    outputs(3035) <= not(layer6_outputs(57));
    outputs(3036) <= not(layer6_outputs(3620));
    outputs(3037) <= not((layer6_outputs(4721)) xor (layer6_outputs(4065)));
    outputs(3038) <= layer6_outputs(4524);
    outputs(3039) <= layer6_outputs(3743);
    outputs(3040) <= not(layer6_outputs(584));
    outputs(3041) <= (layer6_outputs(2562)) and (layer6_outputs(1196));
    outputs(3042) <= layer6_outputs(2794);
    outputs(3043) <= not((layer6_outputs(1563)) and (layer6_outputs(3280)));
    outputs(3044) <= layer6_outputs(2921);
    outputs(3045) <= not((layer6_outputs(2247)) xor (layer6_outputs(2800)));
    outputs(3046) <= (layer6_outputs(1754)) and (layer6_outputs(3658));
    outputs(3047) <= not((layer6_outputs(4198)) xor (layer6_outputs(4639)));
    outputs(3048) <= layer6_outputs(3837);
    outputs(3049) <= layer6_outputs(778);
    outputs(3050) <= not(layer6_outputs(614));
    outputs(3051) <= not(layer6_outputs(2488));
    outputs(3052) <= layer6_outputs(155);
    outputs(3053) <= (layer6_outputs(3)) xor (layer6_outputs(5037));
    outputs(3054) <= not((layer6_outputs(385)) xor (layer6_outputs(4846)));
    outputs(3055) <= layer6_outputs(3261);
    outputs(3056) <= (layer6_outputs(47)) and not (layer6_outputs(1189));
    outputs(3057) <= layer6_outputs(3438);
    outputs(3058) <= layer6_outputs(1764);
    outputs(3059) <= not(layer6_outputs(349));
    outputs(3060) <= not(layer6_outputs(1492));
    outputs(3061) <= not(layer6_outputs(4042));
    outputs(3062) <= not((layer6_outputs(3184)) xor (layer6_outputs(1818)));
    outputs(3063) <= not(layer6_outputs(1850)) or (layer6_outputs(1738));
    outputs(3064) <= not(layer6_outputs(2072));
    outputs(3065) <= not(layer6_outputs(3618));
    outputs(3066) <= (layer6_outputs(4233)) xor (layer6_outputs(296));
    outputs(3067) <= (layer6_outputs(2911)) and (layer6_outputs(1984));
    outputs(3068) <= not(layer6_outputs(251));
    outputs(3069) <= layer6_outputs(3931);
    outputs(3070) <= not(layer6_outputs(3154));
    outputs(3071) <= (layer6_outputs(4456)) and (layer6_outputs(2666));
    outputs(3072) <= not(layer6_outputs(1477));
    outputs(3073) <= not((layer6_outputs(281)) xor (layer6_outputs(3285)));
    outputs(3074) <= layer6_outputs(3890);
    outputs(3075) <= not((layer6_outputs(159)) or (layer6_outputs(1229)));
    outputs(3076) <= layer6_outputs(3238);
    outputs(3077) <= not(layer6_outputs(1474));
    outputs(3078) <= not(layer6_outputs(1999));
    outputs(3079) <= (layer6_outputs(2352)) xor (layer6_outputs(3018));
    outputs(3080) <= not(layer6_outputs(4393)) or (layer6_outputs(5058));
    outputs(3081) <= not(layer6_outputs(932));
    outputs(3082) <= not((layer6_outputs(4088)) xor (layer6_outputs(2657)));
    outputs(3083) <= not(layer6_outputs(2077)) or (layer6_outputs(2085));
    outputs(3084) <= (layer6_outputs(1147)) xor (layer6_outputs(2975));
    outputs(3085) <= not(layer6_outputs(1178));
    outputs(3086) <= (layer6_outputs(3343)) and not (layer6_outputs(3111));
    outputs(3087) <= not(layer6_outputs(2787));
    outputs(3088) <= layer6_outputs(673);
    outputs(3089) <= not(layer6_outputs(486));
    outputs(3090) <= not(layer6_outputs(771));
    outputs(3091) <= (layer6_outputs(1664)) or (layer6_outputs(5118));
    outputs(3092) <= not(layer6_outputs(766));
    outputs(3093) <= layer6_outputs(2463);
    outputs(3094) <= not(layer6_outputs(2341));
    outputs(3095) <= not(layer6_outputs(629));
    outputs(3096) <= not(layer6_outputs(1879));
    outputs(3097) <= (layer6_outputs(4094)) xor (layer6_outputs(4156));
    outputs(3098) <= (layer6_outputs(3564)) xor (layer6_outputs(2589));
    outputs(3099) <= not(layer6_outputs(2635));
    outputs(3100) <= not(layer6_outputs(1691));
    outputs(3101) <= (layer6_outputs(4953)) xor (layer6_outputs(480));
    outputs(3102) <= (layer6_outputs(1509)) and not (layer6_outputs(170));
    outputs(3103) <= layer6_outputs(3408);
    outputs(3104) <= (layer6_outputs(4719)) and not (layer6_outputs(2585));
    outputs(3105) <= layer6_outputs(788);
    outputs(3106) <= (layer6_outputs(4550)) xor (layer6_outputs(12));
    outputs(3107) <= (layer6_outputs(388)) xor (layer6_outputs(67));
    outputs(3108) <= not((layer6_outputs(1359)) xor (layer6_outputs(4284)));
    outputs(3109) <= not(layer6_outputs(4931));
    outputs(3110) <= (layer6_outputs(2489)) and not (layer6_outputs(4288));
    outputs(3111) <= layer6_outputs(619);
    outputs(3112) <= layer6_outputs(639);
    outputs(3113) <= layer6_outputs(4868);
    outputs(3114) <= not((layer6_outputs(4531)) xor (layer6_outputs(1657)));
    outputs(3115) <= layer6_outputs(3321);
    outputs(3116) <= layer6_outputs(211);
    outputs(3117) <= not((layer6_outputs(3710)) xor (layer6_outputs(3615)));
    outputs(3118) <= layer6_outputs(16);
    outputs(3119) <= not(layer6_outputs(3487));
    outputs(3120) <= layer6_outputs(968);
    outputs(3121) <= not(layer6_outputs(2622));
    outputs(3122) <= layer6_outputs(4149);
    outputs(3123) <= layer6_outputs(4321);
    outputs(3124) <= layer6_outputs(366);
    outputs(3125) <= not(layer6_outputs(1084));
    outputs(3126) <= layer6_outputs(4706);
    outputs(3127) <= layer6_outputs(1217);
    outputs(3128) <= layer6_outputs(4897);
    outputs(3129) <= layer6_outputs(1802);
    outputs(3130) <= not(layer6_outputs(109));
    outputs(3131) <= (layer6_outputs(4445)) and (layer6_outputs(4452));
    outputs(3132) <= layer6_outputs(2901);
    outputs(3133) <= (layer6_outputs(4431)) and not (layer6_outputs(813));
    outputs(3134) <= not(layer6_outputs(3849));
    outputs(3135) <= layer6_outputs(4234);
    outputs(3136) <= not(layer6_outputs(3609));
    outputs(3137) <= not(layer6_outputs(4299));
    outputs(3138) <= layer6_outputs(2301);
    outputs(3139) <= layer6_outputs(5107);
    outputs(3140) <= layer6_outputs(1434);
    outputs(3141) <= not(layer6_outputs(918));
    outputs(3142) <= not(layer6_outputs(1219));
    outputs(3143) <= not(layer6_outputs(1198));
    outputs(3144) <= not(layer6_outputs(4000));
    outputs(3145) <= not(layer6_outputs(1401));
    outputs(3146) <= (layer6_outputs(2690)) xor (layer6_outputs(2565));
    outputs(3147) <= (layer6_outputs(3880)) and not (layer6_outputs(4464));
    outputs(3148) <= not(layer6_outputs(3032));
    outputs(3149) <= layer6_outputs(5111);
    outputs(3150) <= layer6_outputs(769);
    outputs(3151) <= not(layer6_outputs(1657));
    outputs(3152) <= not(layer6_outputs(4473));
    outputs(3153) <= not(layer6_outputs(1954));
    outputs(3154) <= layer6_outputs(4733);
    outputs(3155) <= not(layer6_outputs(3452));
    outputs(3156) <= (layer6_outputs(2305)) xor (layer6_outputs(3707));
    outputs(3157) <= not(layer6_outputs(2295));
    outputs(3158) <= layer6_outputs(3959);
    outputs(3159) <= not(layer6_outputs(5103));
    outputs(3160) <= not(layer6_outputs(2189));
    outputs(3161) <= (layer6_outputs(3211)) and not (layer6_outputs(1797));
    outputs(3162) <= (layer6_outputs(2026)) and not (layer6_outputs(4167));
    outputs(3163) <= not(layer6_outputs(4421));
    outputs(3164) <= layer6_outputs(2609);
    outputs(3165) <= (layer6_outputs(5026)) and (layer6_outputs(4723));
    outputs(3166) <= not(layer6_outputs(756));
    outputs(3167) <= not(layer6_outputs(4082));
    outputs(3168) <= not(layer6_outputs(3641));
    outputs(3169) <= not((layer6_outputs(419)) or (layer6_outputs(1351)));
    outputs(3170) <= not(layer6_outputs(409));
    outputs(3171) <= not(layer6_outputs(885));
    outputs(3172) <= layer6_outputs(1718);
    outputs(3173) <= layer6_outputs(2947);
    outputs(3174) <= layer6_outputs(2543);
    outputs(3175) <= layer6_outputs(2159);
    outputs(3176) <= not(layer6_outputs(1575));
    outputs(3177) <= (layer6_outputs(1852)) and not (layer6_outputs(3517));
    outputs(3178) <= (layer6_outputs(1857)) and not (layer6_outputs(2198));
    outputs(3179) <= not((layer6_outputs(4229)) xor (layer6_outputs(3270)));
    outputs(3180) <= not((layer6_outputs(4033)) xor (layer6_outputs(3912)));
    outputs(3181) <= layer6_outputs(1633);
    outputs(3182) <= not(layer6_outputs(2835));
    outputs(3183) <= layer6_outputs(4546);
    outputs(3184) <= not((layer6_outputs(271)) xor (layer6_outputs(566)));
    outputs(3185) <= not(layer6_outputs(1362));
    outputs(3186) <= not(layer6_outputs(2846));
    outputs(3187) <= not(layer6_outputs(3863));
    outputs(3188) <= not(layer6_outputs(2055));
    outputs(3189) <= layer6_outputs(4024);
    outputs(3190) <= layer6_outputs(3662);
    outputs(3191) <= not(layer6_outputs(2188));
    outputs(3192) <= not((layer6_outputs(874)) and (layer6_outputs(315)));
    outputs(3193) <= layer6_outputs(814);
    outputs(3194) <= not(layer6_outputs(2502));
    outputs(3195) <= not(layer6_outputs(1340));
    outputs(3196) <= layer6_outputs(5099);
    outputs(3197) <= (layer6_outputs(3776)) xor (layer6_outputs(465));
    outputs(3198) <= not(layer6_outputs(3619));
    outputs(3199) <= layer6_outputs(1779);
    outputs(3200) <= not(layer6_outputs(3127));
    outputs(3201) <= not((layer6_outputs(1149)) or (layer6_outputs(3196)));
    outputs(3202) <= layer6_outputs(1007);
    outputs(3203) <= (layer6_outputs(2171)) and not (layer6_outputs(4793));
    outputs(3204) <= not((layer6_outputs(4109)) or (layer6_outputs(3781)));
    outputs(3205) <= layer6_outputs(4825);
    outputs(3206) <= layer6_outputs(692);
    outputs(3207) <= not(layer6_outputs(5075)) or (layer6_outputs(4163));
    outputs(3208) <= not(layer6_outputs(303));
    outputs(3209) <= (layer6_outputs(1590)) and (layer6_outputs(2275));
    outputs(3210) <= (layer6_outputs(3397)) and not (layer6_outputs(3121));
    outputs(3211) <= not(layer6_outputs(2464));
    outputs(3212) <= (layer6_outputs(4805)) and (layer6_outputs(3136));
    outputs(3213) <= (layer6_outputs(4988)) and not (layer6_outputs(3261));
    outputs(3214) <= layer6_outputs(1200);
    outputs(3215) <= layer6_outputs(277);
    outputs(3216) <= layer6_outputs(3152);
    outputs(3217) <= layer6_outputs(3100);
    outputs(3218) <= not(layer6_outputs(683));
    outputs(3219) <= layer6_outputs(999);
    outputs(3220) <= not((layer6_outputs(1325)) xor (layer6_outputs(2820)));
    outputs(3221) <= not(layer6_outputs(1370));
    outputs(3222) <= not(layer6_outputs(4757));
    outputs(3223) <= not((layer6_outputs(4179)) and (layer6_outputs(4937)));
    outputs(3224) <= not(layer6_outputs(4275));
    outputs(3225) <= layer6_outputs(240);
    outputs(3226) <= (layer6_outputs(4016)) xor (layer6_outputs(1144));
    outputs(3227) <= (layer6_outputs(1583)) and (layer6_outputs(4556));
    outputs(3228) <= not(layer6_outputs(258));
    outputs(3229) <= layer6_outputs(4988);
    outputs(3230) <= layer6_outputs(2534);
    outputs(3231) <= layer6_outputs(2302);
    outputs(3232) <= not(layer6_outputs(228));
    outputs(3233) <= layer6_outputs(2665);
    outputs(3234) <= (layer6_outputs(943)) xor (layer6_outputs(865));
    outputs(3235) <= not(layer6_outputs(1630));
    outputs(3236) <= layer6_outputs(3586);
    outputs(3237) <= layer6_outputs(982);
    outputs(3238) <= not(layer6_outputs(5053));
    outputs(3239) <= not(layer6_outputs(2375));
    outputs(3240) <= not(layer6_outputs(2701));
    outputs(3241) <= (layer6_outputs(3900)) xor (layer6_outputs(2477));
    outputs(3242) <= not(layer6_outputs(1199));
    outputs(3243) <= not(layer6_outputs(4025));
    outputs(3244) <= not(layer6_outputs(2205));
    outputs(3245) <= (layer6_outputs(113)) xor (layer6_outputs(2378));
    outputs(3246) <= layer6_outputs(3580);
    outputs(3247) <= layer6_outputs(3503);
    outputs(3248) <= layer6_outputs(1966);
    outputs(3249) <= not(layer6_outputs(4469));
    outputs(3250) <= layer6_outputs(2173);
    outputs(3251) <= not(layer6_outputs(3364));
    outputs(3252) <= layer6_outputs(1358);
    outputs(3253) <= layer6_outputs(2817);
    outputs(3254) <= (layer6_outputs(2124)) xor (layer6_outputs(2242));
    outputs(3255) <= not((layer6_outputs(343)) and (layer6_outputs(3233)));
    outputs(3256) <= not(layer6_outputs(4491));
    outputs(3257) <= not(layer6_outputs(585));
    outputs(3258) <= (layer6_outputs(2312)) and not (layer6_outputs(3165));
    outputs(3259) <= layer6_outputs(2600);
    outputs(3260) <= not((layer6_outputs(1770)) xor (layer6_outputs(2942)));
    outputs(3261) <= not(layer6_outputs(572));
    outputs(3262) <= layer6_outputs(1619);
    outputs(3263) <= layer6_outputs(3040);
    outputs(3264) <= not(layer6_outputs(55));
    outputs(3265) <= layer6_outputs(447);
    outputs(3266) <= not((layer6_outputs(1440)) xor (layer6_outputs(115)));
    outputs(3267) <= (layer6_outputs(3562)) and (layer6_outputs(1124));
    outputs(3268) <= layer6_outputs(3845);
    outputs(3269) <= not((layer6_outputs(367)) xor (layer6_outputs(2866)));
    outputs(3270) <= (layer6_outputs(4761)) or (layer6_outputs(3655));
    outputs(3271) <= (layer6_outputs(4572)) xor (layer6_outputs(801));
    outputs(3272) <= layer6_outputs(1989);
    outputs(3273) <= layer6_outputs(4080);
    outputs(3274) <= (layer6_outputs(4650)) xor (layer6_outputs(1033));
    outputs(3275) <= layer6_outputs(4732);
    outputs(3276) <= layer6_outputs(426);
    outputs(3277) <= not((layer6_outputs(2948)) xor (layer6_outputs(1864)));
    outputs(3278) <= layer6_outputs(4640);
    outputs(3279) <= layer6_outputs(1711);
    outputs(3280) <= layer6_outputs(4565);
    outputs(3281) <= not(layer6_outputs(1059));
    outputs(3282) <= not((layer6_outputs(3989)) xor (layer6_outputs(4750)));
    outputs(3283) <= not(layer6_outputs(4131));
    outputs(3284) <= layer6_outputs(3126);
    outputs(3285) <= not((layer6_outputs(4602)) xor (layer6_outputs(3709)));
    outputs(3286) <= layer6_outputs(4878);
    outputs(3287) <= layer6_outputs(4977);
    outputs(3288) <= layer6_outputs(2058);
    outputs(3289) <= layer6_outputs(4681);
    outputs(3290) <= layer6_outputs(1488);
    outputs(3291) <= not(layer6_outputs(2809));
    outputs(3292) <= layer6_outputs(4111);
    outputs(3293) <= not(layer6_outputs(4609));
    outputs(3294) <= layer6_outputs(80);
    outputs(3295) <= not(layer6_outputs(4422));
    outputs(3296) <= layer6_outputs(4599);
    outputs(3297) <= (layer6_outputs(843)) and not (layer6_outputs(2969));
    outputs(3298) <= not(layer6_outputs(2922));
    outputs(3299) <= not(layer6_outputs(4861));
    outputs(3300) <= not(layer6_outputs(3688));
    outputs(3301) <= not(layer6_outputs(3782));
    outputs(3302) <= layer6_outputs(3340);
    outputs(3303) <= (layer6_outputs(4250)) xor (layer6_outputs(471));
    outputs(3304) <= layer6_outputs(4897);
    outputs(3305) <= layer6_outputs(4366);
    outputs(3306) <= layer6_outputs(3693);
    outputs(3307) <= not(layer6_outputs(2205));
    outputs(3308) <= layer6_outputs(4739);
    outputs(3309) <= layer6_outputs(4383);
    outputs(3310) <= (layer6_outputs(2779)) and not (layer6_outputs(1986));
    outputs(3311) <= layer6_outputs(1604);
    outputs(3312) <= layer6_outputs(4111);
    outputs(3313) <= layer6_outputs(4882);
    outputs(3314) <= layer6_outputs(4404);
    outputs(3315) <= not(layer6_outputs(4258));
    outputs(3316) <= not(layer6_outputs(3128));
    outputs(3317) <= not(layer6_outputs(2998));
    outputs(3318) <= layer6_outputs(2661);
    outputs(3319) <= layer6_outputs(764);
    outputs(3320) <= (layer6_outputs(1889)) xor (layer6_outputs(790));
    outputs(3321) <= not((layer6_outputs(4601)) xor (layer6_outputs(760)));
    outputs(3322) <= not((layer6_outputs(3009)) and (layer6_outputs(4376)));
    outputs(3323) <= (layer6_outputs(3541)) xor (layer6_outputs(2582));
    outputs(3324) <= layer6_outputs(2020);
    outputs(3325) <= layer6_outputs(4908);
    outputs(3326) <= not(layer6_outputs(922));
    outputs(3327) <= (layer6_outputs(458)) and not (layer6_outputs(2649));
    outputs(3328) <= not(layer6_outputs(3538));
    outputs(3329) <= not((layer6_outputs(5063)) xor (layer6_outputs(1764)));
    outputs(3330) <= layer6_outputs(1868);
    outputs(3331) <= (layer6_outputs(4251)) and (layer6_outputs(3458));
    outputs(3332) <= layer6_outputs(3485);
    outputs(3333) <= not(layer6_outputs(682));
    outputs(3334) <= (layer6_outputs(3417)) and not (layer6_outputs(2730));
    outputs(3335) <= layer6_outputs(4367);
    outputs(3336) <= not(layer6_outputs(4722));
    outputs(3337) <= layer6_outputs(3474);
    outputs(3338) <= layer6_outputs(952);
    outputs(3339) <= not(layer6_outputs(2644));
    outputs(3340) <= not(layer6_outputs(2331));
    outputs(3341) <= not(layer6_outputs(1205));
    outputs(3342) <= (layer6_outputs(3322)) xor (layer6_outputs(2521));
    outputs(3343) <= not(layer6_outputs(1322));
    outputs(3344) <= layer6_outputs(1010);
    outputs(3345) <= layer6_outputs(2422);
    outputs(3346) <= not(layer6_outputs(3409)) or (layer6_outputs(3210));
    outputs(3347) <= not(layer6_outputs(2841));
    outputs(3348) <= (layer6_outputs(4220)) and (layer6_outputs(3471));
    outputs(3349) <= layer6_outputs(3443);
    outputs(3350) <= layer6_outputs(4279);
    outputs(3351) <= not(layer6_outputs(2562));
    outputs(3352) <= not(layer6_outputs(907));
    outputs(3353) <= not(layer6_outputs(1832));
    outputs(3354) <= not(layer6_outputs(2862));
    outputs(3355) <= layer6_outputs(124);
    outputs(3356) <= layer6_outputs(2001);
    outputs(3357) <= layer6_outputs(631);
    outputs(3358) <= layer6_outputs(4440);
    outputs(3359) <= layer6_outputs(2641);
    outputs(3360) <= not(layer6_outputs(2759));
    outputs(3361) <= not(layer6_outputs(122));
    outputs(3362) <= not(layer6_outputs(3215));
    outputs(3363) <= not(layer6_outputs(2570));
    outputs(3364) <= layer6_outputs(347);
    outputs(3365) <= layer6_outputs(3940);
    outputs(3366) <= not(layer6_outputs(137)) or (layer6_outputs(1941));
    outputs(3367) <= not(layer6_outputs(781));
    outputs(3368) <= not((layer6_outputs(3910)) or (layer6_outputs(3814)));
    outputs(3369) <= layer6_outputs(3916);
    outputs(3370) <= not(layer6_outputs(60));
    outputs(3371) <= not((layer6_outputs(1780)) and (layer6_outputs(3902)));
    outputs(3372) <= not(layer6_outputs(2946)) or (layer6_outputs(3901));
    outputs(3373) <= not(layer6_outputs(3147));
    outputs(3374) <= (layer6_outputs(5079)) and not (layer6_outputs(2068));
    outputs(3375) <= layer6_outputs(3752);
    outputs(3376) <= not((layer6_outputs(5115)) xor (layer6_outputs(2363)));
    outputs(3377) <= layer6_outputs(578);
    outputs(3378) <= not(layer6_outputs(786));
    outputs(3379) <= not(layer6_outputs(2957));
    outputs(3380) <= not(layer6_outputs(2057));
    outputs(3381) <= layer6_outputs(1898);
    outputs(3382) <= layer6_outputs(3003);
    outputs(3383) <= layer6_outputs(1431);
    outputs(3384) <= not((layer6_outputs(579)) and (layer6_outputs(3077)));
    outputs(3385) <= not(layer6_outputs(725));
    outputs(3386) <= not(layer6_outputs(2933));
    outputs(3387) <= layer6_outputs(722);
    outputs(3388) <= layer6_outputs(1793);
    outputs(3389) <= (layer6_outputs(3259)) and not (layer6_outputs(2174));
    outputs(3390) <= not(layer6_outputs(1649));
    outputs(3391) <= not(layer6_outputs(322));
    outputs(3392) <= (layer6_outputs(770)) and not (layer6_outputs(3146));
    outputs(3393) <= layer6_outputs(465);
    outputs(3394) <= not(layer6_outputs(2938));
    outputs(3395) <= layer6_outputs(3511);
    outputs(3396) <= (layer6_outputs(2765)) and not (layer6_outputs(1512));
    outputs(3397) <= layer6_outputs(75);
    outputs(3398) <= layer6_outputs(3068);
    outputs(3399) <= not(layer6_outputs(1979));
    outputs(3400) <= not((layer6_outputs(3587)) xor (layer6_outputs(1498)));
    outputs(3401) <= not(layer6_outputs(2989));
    outputs(3402) <= not(layer6_outputs(4374));
    outputs(3403) <= layer6_outputs(4876);
    outputs(3404) <= not(layer6_outputs(2148));
    outputs(3405) <= layer6_outputs(571);
    outputs(3406) <= layer6_outputs(1029);
    outputs(3407) <= (layer6_outputs(2097)) xor (layer6_outputs(436));
    outputs(3408) <= layer6_outputs(3477);
    outputs(3409) <= layer6_outputs(4834);
    outputs(3410) <= (layer6_outputs(2270)) and not (layer6_outputs(776));
    outputs(3411) <= not(layer6_outputs(1910));
    outputs(3412) <= (layer6_outputs(1264)) and not (layer6_outputs(4124));
    outputs(3413) <= not(layer6_outputs(1077));
    outputs(3414) <= (layer6_outputs(2412)) xor (layer6_outputs(428));
    outputs(3415) <= (layer6_outputs(1621)) and (layer6_outputs(2773));
    outputs(3416) <= (layer6_outputs(1302)) xor (layer6_outputs(3750));
    outputs(3417) <= not(layer6_outputs(4527));
    outputs(3418) <= not(layer6_outputs(3333));
    outputs(3419) <= not((layer6_outputs(2616)) xor (layer6_outputs(4261)));
    outputs(3420) <= not(layer6_outputs(431));
    outputs(3421) <= not(layer6_outputs(2336));
    outputs(3422) <= layer6_outputs(1505);
    outputs(3423) <= not(layer6_outputs(3451)) or (layer6_outputs(1727));
    outputs(3424) <= not(layer6_outputs(4753));
    outputs(3425) <= not(layer6_outputs(2334));
    outputs(3426) <= not(layer6_outputs(559));
    outputs(3427) <= (layer6_outputs(3408)) and not (layer6_outputs(3720));
    outputs(3428) <= layer6_outputs(3197);
    outputs(3429) <= layer6_outputs(1094);
    outputs(3430) <= not(layer6_outputs(558)) or (layer6_outputs(3685));
    outputs(3431) <= layer6_outputs(3597);
    outputs(3432) <= not(layer6_outputs(1990));
    outputs(3433) <= not((layer6_outputs(4587)) or (layer6_outputs(3492)));
    outputs(3434) <= (layer6_outputs(688)) xor (layer6_outputs(2528));
    outputs(3435) <= layer6_outputs(3735);
    outputs(3436) <= not(layer6_outputs(2363));
    outputs(3437) <= not(layer6_outputs(4138));
    outputs(3438) <= not(layer6_outputs(4973));
    outputs(3439) <= (layer6_outputs(1591)) and not (layer6_outputs(4238));
    outputs(3440) <= not(layer6_outputs(2961));
    outputs(3441) <= not((layer6_outputs(4036)) or (layer6_outputs(4575)));
    outputs(3442) <= layer6_outputs(3368);
    outputs(3443) <= layer6_outputs(1702);
    outputs(3444) <= not(layer6_outputs(92));
    outputs(3445) <= not(layer6_outputs(1114));
    outputs(3446) <= not(layer6_outputs(2152));
    outputs(3447) <= not(layer6_outputs(4872));
    outputs(3448) <= not(layer6_outputs(2961));
    outputs(3449) <= not(layer6_outputs(4276)) or (layer6_outputs(4500));
    outputs(3450) <= (layer6_outputs(3660)) or (layer6_outputs(114));
    outputs(3451) <= layer6_outputs(1905);
    outputs(3452) <= not(layer6_outputs(1678)) or (layer6_outputs(1810));
    outputs(3453) <= not(layer6_outputs(231));
    outputs(3454) <= layer6_outputs(4263);
    outputs(3455) <= layer6_outputs(4970);
    outputs(3456) <= not((layer6_outputs(3328)) or (layer6_outputs(4121)));
    outputs(3457) <= not(layer6_outputs(2234));
    outputs(3458) <= layer6_outputs(1791);
    outputs(3459) <= layer6_outputs(1896);
    outputs(3460) <= layer6_outputs(3149);
    outputs(3461) <= layer6_outputs(584);
    outputs(3462) <= not((layer6_outputs(3674)) or (layer6_outputs(1392)));
    outputs(3463) <= not(layer6_outputs(806));
    outputs(3464) <= not(layer6_outputs(1728)) or (layer6_outputs(2277));
    outputs(3465) <= not(layer6_outputs(427));
    outputs(3466) <= not(layer6_outputs(4466));
    outputs(3467) <= not(layer6_outputs(2892));
    outputs(3468) <= layer6_outputs(2605);
    outputs(3469) <= layer6_outputs(3169);
    outputs(3470) <= not(layer6_outputs(1415));
    outputs(3471) <= not(layer6_outputs(4801));
    outputs(3472) <= not(layer6_outputs(4449));
    outputs(3473) <= layer6_outputs(3126);
    outputs(3474) <= not(layer6_outputs(676));
    outputs(3475) <= not((layer6_outputs(2900)) or (layer6_outputs(2437)));
    outputs(3476) <= layer6_outputs(1774);
    outputs(3477) <= layer6_outputs(2968);
    outputs(3478) <= layer6_outputs(4981);
    outputs(3479) <= layer6_outputs(741);
    outputs(3480) <= layer6_outputs(3687);
    outputs(3481) <= (layer6_outputs(4618)) and not (layer6_outputs(2014));
    outputs(3482) <= layer6_outputs(3937);
    outputs(3483) <= layer6_outputs(822);
    outputs(3484) <= layer6_outputs(3154);
    outputs(3485) <= (layer6_outputs(989)) and (layer6_outputs(4442));
    outputs(3486) <= not((layer6_outputs(1316)) xor (layer6_outputs(4820)));
    outputs(3487) <= layer6_outputs(4239);
    outputs(3488) <= not(layer6_outputs(3374));
    outputs(3489) <= not(layer6_outputs(2992));
    outputs(3490) <= layer6_outputs(2265);
    outputs(3491) <= (layer6_outputs(2110)) and not (layer6_outputs(3389));
    outputs(3492) <= layer6_outputs(1146);
    outputs(3493) <= layer6_outputs(3731);
    outputs(3494) <= not(layer6_outputs(795));
    outputs(3495) <= layer6_outputs(769);
    outputs(3496) <= layer6_outputs(2423);
    outputs(3497) <= not(layer6_outputs(1998));
    outputs(3498) <= not(layer6_outputs(3061));
    outputs(3499) <= not(layer6_outputs(1797));
    outputs(3500) <= layer6_outputs(1565);
    outputs(3501) <= layer6_outputs(1944);
    outputs(3502) <= layer6_outputs(1951);
    outputs(3503) <= (layer6_outputs(84)) and (layer6_outputs(4328));
    outputs(3504) <= not(layer6_outputs(1109));
    outputs(3505) <= (layer6_outputs(1121)) and not (layer6_outputs(681));
    outputs(3506) <= not(layer6_outputs(908)) or (layer6_outputs(2887));
    outputs(3507) <= not(layer6_outputs(3046));
    outputs(3508) <= not(layer6_outputs(149));
    outputs(3509) <= layer6_outputs(1494);
    outputs(3510) <= not((layer6_outputs(3561)) xor (layer6_outputs(795)));
    outputs(3511) <= not(layer6_outputs(4720));
    outputs(3512) <= layer6_outputs(4703);
    outputs(3513) <= layer6_outputs(3771);
    outputs(3514) <= not((layer6_outputs(4788)) xor (layer6_outputs(3036)));
    outputs(3515) <= not((layer6_outputs(4910)) xor (layer6_outputs(83)));
    outputs(3516) <= not(layer6_outputs(4769));
    outputs(3517) <= layer6_outputs(4729);
    outputs(3518) <= layer6_outputs(2226);
    outputs(3519) <= layer6_outputs(5029);
    outputs(3520) <= not(layer6_outputs(2792));
    outputs(3521) <= not(layer6_outputs(3704));
    outputs(3522) <= not(layer6_outputs(3501));
    outputs(3523) <= not(layer6_outputs(3992));
    outputs(3524) <= layer6_outputs(1015);
    outputs(3525) <= layer6_outputs(688);
    outputs(3526) <= (layer6_outputs(123)) xor (layer6_outputs(4636));
    outputs(3527) <= (layer6_outputs(2401)) xor (layer6_outputs(1039));
    outputs(3528) <= not(layer6_outputs(1953)) or (layer6_outputs(374));
    outputs(3529) <= not(layer6_outputs(871));
    outputs(3530) <= not(layer6_outputs(3772)) or (layer6_outputs(2117));
    outputs(3531) <= not(layer6_outputs(2696));
    outputs(3532) <= (layer6_outputs(1509)) and not (layer6_outputs(3196));
    outputs(3533) <= not(layer6_outputs(2418));
    outputs(3534) <= layer6_outputs(5057);
    outputs(3535) <= layer6_outputs(610);
    outputs(3536) <= not(layer6_outputs(1632)) or (layer6_outputs(2568));
    outputs(3537) <= not(layer6_outputs(12));
    outputs(3538) <= not((layer6_outputs(2037)) or (layer6_outputs(1574)));
    outputs(3539) <= layer6_outputs(3471);
    outputs(3540) <= not(layer6_outputs(101));
    outputs(3541) <= layer6_outputs(4213);
    outputs(3542) <= layer6_outputs(961);
    outputs(3543) <= layer6_outputs(3391);
    outputs(3544) <= not(layer6_outputs(1351));
    outputs(3545) <= not((layer6_outputs(3588)) xor (layer6_outputs(2433)));
    outputs(3546) <= (layer6_outputs(5070)) and (layer6_outputs(840));
    outputs(3547) <= not(layer6_outputs(1059));
    outputs(3548) <= not(layer6_outputs(2234));
    outputs(3549) <= layer6_outputs(2880);
    outputs(3550) <= not(layer6_outputs(3607));
    outputs(3551) <= not(layer6_outputs(1183));
    outputs(3552) <= (layer6_outputs(3685)) xor (layer6_outputs(1258));
    outputs(3553) <= layer6_outputs(3378);
    outputs(3554) <= not(layer6_outputs(3356));
    outputs(3555) <= not(layer6_outputs(4374));
    outputs(3556) <= not(layer6_outputs(1999));
    outputs(3557) <= layer6_outputs(4471);
    outputs(3558) <= not(layer6_outputs(541));
    outputs(3559) <= not(layer6_outputs(2351));
    outputs(3560) <= not(layer6_outputs(23));
    outputs(3561) <= not(layer6_outputs(1277));
    outputs(3562) <= layer6_outputs(1110);
    outputs(3563) <= not((layer6_outputs(27)) and (layer6_outputs(2771)));
    outputs(3564) <= layer6_outputs(796);
    outputs(3565) <= not(layer6_outputs(1737));
    outputs(3566) <= layer6_outputs(763);
    outputs(3567) <= not(layer6_outputs(2139));
    outputs(3568) <= (layer6_outputs(2102)) xor (layer6_outputs(2252));
    outputs(3569) <= layer6_outputs(1131);
    outputs(3570) <= layer6_outputs(613);
    outputs(3571) <= not(layer6_outputs(77));
    outputs(3572) <= not(layer6_outputs(2163));
    outputs(3573) <= layer6_outputs(232);
    outputs(3574) <= layer6_outputs(79);
    outputs(3575) <= not(layer6_outputs(296));
    outputs(3576) <= layer6_outputs(4314);
    outputs(3577) <= layer6_outputs(4319);
    outputs(3578) <= not(layer6_outputs(3434));
    outputs(3579) <= not((layer6_outputs(1033)) xor (layer6_outputs(485)));
    outputs(3580) <= layer6_outputs(4788);
    outputs(3581) <= (layer6_outputs(3753)) xor (layer6_outputs(2958));
    outputs(3582) <= layer6_outputs(4511);
    outputs(3583) <= not(layer6_outputs(891));
    outputs(3584) <= not(layer6_outputs(3377));
    outputs(3585) <= '1';
    outputs(3586) <= layer6_outputs(1173);
    outputs(3587) <= layer6_outputs(1240);
    outputs(3588) <= layer6_outputs(2800);
    outputs(3589) <= not((layer6_outputs(2225)) or (layer6_outputs(701)));
    outputs(3590) <= not(layer6_outputs(3959));
    outputs(3591) <= (layer6_outputs(2518)) and not (layer6_outputs(1522));
    outputs(3592) <= not(layer6_outputs(4984));
    outputs(3593) <= layer6_outputs(3911);
    outputs(3594) <= layer6_outputs(1176);
    outputs(3595) <= not(layer6_outputs(1170));
    outputs(3596) <= not(layer6_outputs(1076));
    outputs(3597) <= not(layer6_outputs(627)) or (layer6_outputs(1824));
    outputs(3598) <= layer6_outputs(1983);
    outputs(3599) <= layer6_outputs(276);
    outputs(3600) <= (layer6_outputs(356)) xor (layer6_outputs(2083));
    outputs(3601) <= not((layer6_outputs(2027)) or (layer6_outputs(4171)));
    outputs(3602) <= layer6_outputs(4985);
    outputs(3603) <= layer6_outputs(3635);
    outputs(3604) <= not(layer6_outputs(2540));
    outputs(3605) <= not((layer6_outputs(391)) or (layer6_outputs(3524)));
    outputs(3606) <= not(layer6_outputs(1848));
    outputs(3607) <= not((layer6_outputs(780)) xor (layer6_outputs(2428)));
    outputs(3608) <= layer6_outputs(2681);
    outputs(3609) <= layer6_outputs(3987);
    outputs(3610) <= layer6_outputs(4510);
    outputs(3611) <= not(layer6_outputs(3536));
    outputs(3612) <= (layer6_outputs(3414)) xor (layer6_outputs(3677));
    outputs(3613) <= not(layer6_outputs(926));
    outputs(3614) <= not(layer6_outputs(1834));
    outputs(3615) <= not(layer6_outputs(3169));
    outputs(3616) <= layer6_outputs(4589);
    outputs(3617) <= (layer6_outputs(97)) and (layer6_outputs(4007));
    outputs(3618) <= layer6_outputs(3311);
    outputs(3619) <= layer6_outputs(309);
    outputs(3620) <= layer6_outputs(1222);
    outputs(3621) <= not((layer6_outputs(71)) xor (layer6_outputs(4013)));
    outputs(3622) <= layer6_outputs(1692);
    outputs(3623) <= not(layer6_outputs(4054));
    outputs(3624) <= not(layer6_outputs(4443));
    outputs(3625) <= not(layer6_outputs(67)) or (layer6_outputs(1176));
    outputs(3626) <= layer6_outputs(5068);
    outputs(3627) <= not(layer6_outputs(3513));
    outputs(3628) <= not((layer6_outputs(703)) xor (layer6_outputs(3106)));
    outputs(3629) <= not(layer6_outputs(3743));
    outputs(3630) <= (layer6_outputs(632)) and not (layer6_outputs(3706));
    outputs(3631) <= not((layer6_outputs(3141)) xor (layer6_outputs(4108)));
    outputs(3632) <= not(layer6_outputs(3245));
    outputs(3633) <= layer6_outputs(3891);
    outputs(3634) <= layer6_outputs(3953);
    outputs(3635) <= layer6_outputs(375);
    outputs(3636) <= layer6_outputs(2143);
    outputs(3637) <= not(layer6_outputs(1405));
    outputs(3638) <= not(layer6_outputs(269));
    outputs(3639) <= not((layer6_outputs(184)) xor (layer6_outputs(2881)));
    outputs(3640) <= not(layer6_outputs(1476));
    outputs(3641) <= not((layer6_outputs(3948)) xor (layer6_outputs(4461)));
    outputs(3642) <= layer6_outputs(4493);
    outputs(3643) <= not(layer6_outputs(2763));
    outputs(3644) <= (layer6_outputs(2606)) and not (layer6_outputs(1245));
    outputs(3645) <= (layer6_outputs(2039)) xor (layer6_outputs(4458));
    outputs(3646) <= layer6_outputs(4763);
    outputs(3647) <= layer6_outputs(4088);
    outputs(3648) <= not(layer6_outputs(1238));
    outputs(3649) <= layer6_outputs(1528);
    outputs(3650) <= not(layer6_outputs(1078));
    outputs(3651) <= (layer6_outputs(3785)) and (layer6_outputs(1547));
    outputs(3652) <= (layer6_outputs(4869)) xor (layer6_outputs(1919));
    outputs(3653) <= (layer6_outputs(2693)) xor (layer6_outputs(2191));
    outputs(3654) <= (layer6_outputs(435)) xor (layer6_outputs(4129));
    outputs(3655) <= layer6_outputs(4242);
    outputs(3656) <= not(layer6_outputs(4895));
    outputs(3657) <= layer6_outputs(4425);
    outputs(3658) <= not(layer6_outputs(4673));
    outputs(3659) <= not((layer6_outputs(4492)) and (layer6_outputs(510)));
    outputs(3660) <= layer6_outputs(4935);
    outputs(3661) <= layer6_outputs(1370);
    outputs(3662) <= layer6_outputs(1393);
    outputs(3663) <= (layer6_outputs(696)) and (layer6_outputs(2918));
    outputs(3664) <= layer6_outputs(2834);
    outputs(3665) <= (layer6_outputs(4203)) xor (layer6_outputs(2456));
    outputs(3666) <= layer6_outputs(2942);
    outputs(3667) <= layer6_outputs(3804);
    outputs(3668) <= not(layer6_outputs(2133));
    outputs(3669) <= layer6_outputs(3609);
    outputs(3670) <= layer6_outputs(4843);
    outputs(3671) <= not(layer6_outputs(4504));
    outputs(3672) <= (layer6_outputs(2168)) or (layer6_outputs(1414));
    outputs(3673) <= layer6_outputs(832);
    outputs(3674) <= not(layer6_outputs(2648));
    outputs(3675) <= not(layer6_outputs(4755)) or (layer6_outputs(478));
    outputs(3676) <= layer6_outputs(3142);
    outputs(3677) <= (layer6_outputs(2052)) xor (layer6_outputs(4716));
    outputs(3678) <= not((layer6_outputs(659)) xor (layer6_outputs(1727)));
    outputs(3679) <= not(layer6_outputs(4900));
    outputs(3680) <= not(layer6_outputs(4174));
    outputs(3681) <= not(layer6_outputs(1814));
    outputs(3682) <= (layer6_outputs(3865)) and (layer6_outputs(1034));
    outputs(3683) <= not((layer6_outputs(3963)) xor (layer6_outputs(3694)));
    outputs(3684) <= (layer6_outputs(816)) and not (layer6_outputs(4450));
    outputs(3685) <= not((layer6_outputs(4141)) xor (layer6_outputs(2866)));
    outputs(3686) <= layer6_outputs(1865);
    outputs(3687) <= not((layer6_outputs(1335)) and (layer6_outputs(286)));
    outputs(3688) <= layer6_outputs(1879);
    outputs(3689) <= (layer6_outputs(1887)) xor (layer6_outputs(1561));
    outputs(3690) <= not(layer6_outputs(3886));
    outputs(3691) <= not(layer6_outputs(189));
    outputs(3692) <= not(layer6_outputs(4463));
    outputs(3693) <= layer6_outputs(455);
    outputs(3694) <= not(layer6_outputs(1364));
    outputs(3695) <= not((layer6_outputs(4538)) xor (layer6_outputs(3449)));
    outputs(3696) <= layer6_outputs(4281);
    outputs(3697) <= (layer6_outputs(3445)) xor (layer6_outputs(916));
    outputs(3698) <= (layer6_outputs(3357)) and (layer6_outputs(2129));
    outputs(3699) <= (layer6_outputs(2266)) xor (layer6_outputs(426));
    outputs(3700) <= layer6_outputs(1771);
    outputs(3701) <= not(layer6_outputs(2149)) or (layer6_outputs(3975));
    outputs(3702) <= layer6_outputs(3333);
    outputs(3703) <= not(layer6_outputs(3841));
    outputs(3704) <= (layer6_outputs(4657)) and not (layer6_outputs(195));
    outputs(3705) <= (layer6_outputs(1619)) xor (layer6_outputs(324));
    outputs(3706) <= layer6_outputs(2926);
    outputs(3707) <= not(layer6_outputs(1788));
    outputs(3708) <= not(layer6_outputs(2302));
    outputs(3709) <= not(layer6_outputs(3971));
    outputs(3710) <= layer6_outputs(924);
    outputs(3711) <= layer6_outputs(3809);
    outputs(3712) <= not(layer6_outputs(3757));
    outputs(3713) <= not((layer6_outputs(2575)) or (layer6_outputs(2095)));
    outputs(3714) <= layer6_outputs(5052);
    outputs(3715) <= not(layer6_outputs(3914));
    outputs(3716) <= layer6_outputs(3425);
    outputs(3717) <= layer6_outputs(4096);
    outputs(3718) <= not((layer6_outputs(4693)) xor (layer6_outputs(162)));
    outputs(3719) <= not(layer6_outputs(2986));
    outputs(3720) <= not((layer6_outputs(1143)) xor (layer6_outputs(4878)));
    outputs(3721) <= not(layer6_outputs(2505));
    outputs(3722) <= not((layer6_outputs(3885)) xor (layer6_outputs(2105)));
    outputs(3723) <= layer6_outputs(2169);
    outputs(3724) <= not(layer6_outputs(4966)) or (layer6_outputs(1876));
    outputs(3725) <= not(layer6_outputs(1867));
    outputs(3726) <= not(layer6_outputs(4865));
    outputs(3727) <= layer6_outputs(3642);
    outputs(3728) <= layer6_outputs(567);
    outputs(3729) <= not(layer6_outputs(295));
    outputs(3730) <= not(layer6_outputs(3675));
    outputs(3731) <= not(layer6_outputs(3976));
    outputs(3732) <= (layer6_outputs(1383)) xor (layer6_outputs(1878));
    outputs(3733) <= not(layer6_outputs(3668));
    outputs(3734) <= not((layer6_outputs(3274)) and (layer6_outputs(4329)));
    outputs(3735) <= (layer6_outputs(3784)) or (layer6_outputs(470));
    outputs(3736) <= (layer6_outputs(3892)) xor (layer6_outputs(3628));
    outputs(3737) <= (layer6_outputs(3459)) and (layer6_outputs(2431));
    outputs(3738) <= not(layer6_outputs(1300));
    outputs(3739) <= layer6_outputs(2164);
    outputs(3740) <= not((layer6_outputs(1496)) xor (layer6_outputs(1697)));
    outputs(3741) <= not((layer6_outputs(3634)) and (layer6_outputs(2425)));
    outputs(3742) <= not((layer6_outputs(4003)) xor (layer6_outputs(2579)));
    outputs(3743) <= not((layer6_outputs(3299)) xor (layer6_outputs(1441)));
    outputs(3744) <= not(layer6_outputs(2406));
    outputs(3745) <= not(layer6_outputs(1106));
    outputs(3746) <= layer6_outputs(2515);
    outputs(3747) <= not(layer6_outputs(1621));
    outputs(3748) <= not(layer6_outputs(37));
    outputs(3749) <= layer6_outputs(2731);
    outputs(3750) <= not(layer6_outputs(5041));
    outputs(3751) <= (layer6_outputs(4373)) xor (layer6_outputs(1263));
    outputs(3752) <= not((layer6_outputs(2486)) xor (layer6_outputs(4378)));
    outputs(3753) <= not(layer6_outputs(1726));
    outputs(3754) <= layer6_outputs(3917);
    outputs(3755) <= (layer6_outputs(2456)) and not (layer6_outputs(4757));
    outputs(3756) <= (layer6_outputs(4537)) xor (layer6_outputs(4541));
    outputs(3757) <= not((layer6_outputs(2686)) xor (layer6_outputs(718)));
    outputs(3758) <= layer6_outputs(309);
    outputs(3759) <= not(layer6_outputs(3867));
    outputs(3760) <= (layer6_outputs(4944)) and not (layer6_outputs(1010));
    outputs(3761) <= layer6_outputs(2134);
    outputs(3762) <= layer6_outputs(292);
    outputs(3763) <= layer6_outputs(3678);
    outputs(3764) <= layer6_outputs(3388);
    outputs(3765) <= not((layer6_outputs(2937)) or (layer6_outputs(785)));
    outputs(3766) <= layer6_outputs(4746);
    outputs(3767) <= not((layer6_outputs(972)) xor (layer6_outputs(685)));
    outputs(3768) <= layer6_outputs(5073);
    outputs(3769) <= layer6_outputs(3656);
    outputs(3770) <= layer6_outputs(757);
    outputs(3771) <= not(layer6_outputs(4739));
    outputs(3772) <= not(layer6_outputs(4372));
    outputs(3773) <= layer6_outputs(1453);
    outputs(3774) <= not((layer6_outputs(4994)) xor (layer6_outputs(4658)));
    outputs(3775) <= layer6_outputs(3999);
    outputs(3776) <= not((layer6_outputs(75)) xor (layer6_outputs(262)));
    outputs(3777) <= layer6_outputs(3323);
    outputs(3778) <= not(layer6_outputs(4927));
    outputs(3779) <= layer6_outputs(3241);
    outputs(3780) <= layer6_outputs(1087);
    outputs(3781) <= (layer6_outputs(3182)) and not (layer6_outputs(2864));
    outputs(3782) <= (layer6_outputs(4180)) and not (layer6_outputs(1517));
    outputs(3783) <= (layer6_outputs(2983)) xor (layer6_outputs(5045));
    outputs(3784) <= not(layer6_outputs(1553));
    outputs(3785) <= '0';
    outputs(3786) <= not((layer6_outputs(4245)) xor (layer6_outputs(1664)));
    outputs(3787) <= not(layer6_outputs(2547));
    outputs(3788) <= layer6_outputs(4145);
    outputs(3789) <= not(layer6_outputs(2959));
    outputs(3790) <= not(layer6_outputs(689));
    outputs(3791) <= not((layer6_outputs(3522)) or (layer6_outputs(1397)));
    outputs(3792) <= layer6_outputs(1836);
    outputs(3793) <= layer6_outputs(683);
    outputs(3794) <= not((layer6_outputs(3697)) xor (layer6_outputs(2758)));
    outputs(3795) <= not((layer6_outputs(2415)) xor (layer6_outputs(4097)));
    outputs(3796) <= not(layer6_outputs(411));
    outputs(3797) <= not(layer6_outputs(3239));
    outputs(3798) <= not(layer6_outputs(2675));
    outputs(3799) <= not((layer6_outputs(3215)) xor (layer6_outputs(1566)));
    outputs(3800) <= not(layer6_outputs(2768));
    outputs(3801) <= layer6_outputs(2108);
    outputs(3802) <= (layer6_outputs(4701)) and (layer6_outputs(4449));
    outputs(3803) <= not(layer6_outputs(2049));
    outputs(3804) <= not(layer6_outputs(2476));
    outputs(3805) <= layer6_outputs(3425);
    outputs(3806) <= not(layer6_outputs(4249));
    outputs(3807) <= not(layer6_outputs(835));
    outputs(3808) <= layer6_outputs(2104);
    outputs(3809) <= (layer6_outputs(164)) and (layer6_outputs(3865));
    outputs(3810) <= (layer6_outputs(4390)) and not (layer6_outputs(1384));
    outputs(3811) <= layer6_outputs(4312);
    outputs(3812) <= not((layer6_outputs(4728)) xor (layer6_outputs(2956)));
    outputs(3813) <= not(layer6_outputs(3962));
    outputs(3814) <= (layer6_outputs(3494)) xor (layer6_outputs(3718));
    outputs(3815) <= not(layer6_outputs(1654));
    outputs(3816) <= layer6_outputs(717);
    outputs(3817) <= layer6_outputs(4472);
    outputs(3818) <= layer6_outputs(202);
    outputs(3819) <= not(layer6_outputs(2574));
    outputs(3820) <= not(layer6_outputs(2348));
    outputs(3821) <= not((layer6_outputs(3590)) xor (layer6_outputs(4693)));
    outputs(3822) <= not(layer6_outputs(2591));
    outputs(3823) <= layer6_outputs(166);
    outputs(3824) <= layer6_outputs(393);
    outputs(3825) <= layer6_outputs(4943);
    outputs(3826) <= not(layer6_outputs(429));
    outputs(3827) <= not(layer6_outputs(2337)) or (layer6_outputs(2471));
    outputs(3828) <= not(layer6_outputs(3016)) or (layer6_outputs(3412));
    outputs(3829) <= not(layer6_outputs(3571));
    outputs(3830) <= layer6_outputs(2971);
    outputs(3831) <= not(layer6_outputs(2413));
    outputs(3832) <= not(layer6_outputs(1682));
    outputs(3833) <= not(layer6_outputs(106));
    outputs(3834) <= layer6_outputs(327);
    outputs(3835) <= not(layer6_outputs(1218));
    outputs(3836) <= layer6_outputs(1412);
    outputs(3837) <= (layer6_outputs(216)) and not (layer6_outputs(1508));
    outputs(3838) <= not((layer6_outputs(4462)) xor (layer6_outputs(1294)));
    outputs(3839) <= layer6_outputs(3558);
    outputs(3840) <= layer6_outputs(2917);
    outputs(3841) <= (layer6_outputs(798)) xor (layer6_outputs(4645));
    outputs(3842) <= (layer6_outputs(4993)) or (layer6_outputs(1882));
    outputs(3843) <= not(layer6_outputs(2909));
    outputs(3844) <= (layer6_outputs(174)) xor (layer6_outputs(5115));
    outputs(3845) <= layer6_outputs(4040);
    outputs(3846) <= not(layer6_outputs(2126));
    outputs(3847) <= not(layer6_outputs(896));
    outputs(3848) <= (layer6_outputs(698)) and not (layer6_outputs(596));
    outputs(3849) <= not(layer6_outputs(2420));
    outputs(3850) <= not((layer6_outputs(234)) xor (layer6_outputs(1515)));
    outputs(3851) <= not(layer6_outputs(4135));
    outputs(3852) <= layer6_outputs(3457);
    outputs(3853) <= not(layer6_outputs(4015));
    outputs(3854) <= not((layer6_outputs(4213)) xor (layer6_outputs(2075)));
    outputs(3855) <= not((layer6_outputs(2838)) xor (layer6_outputs(4613)));
    outputs(3856) <= layer6_outputs(1743);
    outputs(3857) <= not(layer6_outputs(4345));
    outputs(3858) <= not(layer6_outputs(4110));
    outputs(3859) <= not(layer6_outputs(2038));
    outputs(3860) <= not((layer6_outputs(1585)) xor (layer6_outputs(2441)));
    outputs(3861) <= layer6_outputs(3785);
    outputs(3862) <= not(layer6_outputs(1405));
    outputs(3863) <= (layer6_outputs(2069)) xor (layer6_outputs(2580));
    outputs(3864) <= not(layer6_outputs(2909));
    outputs(3865) <= not(layer6_outputs(4580));
    outputs(3866) <= layer6_outputs(4487);
    outputs(3867) <= layer6_outputs(1268);
    outputs(3868) <= (layer6_outputs(3164)) and not (layer6_outputs(5080));
    outputs(3869) <= not((layer6_outputs(4224)) xor (layer6_outputs(1895)));
    outputs(3870) <= layer6_outputs(4435);
    outputs(3871) <= layer6_outputs(2772);
    outputs(3872) <= layer6_outputs(188);
    outputs(3873) <= layer6_outputs(3275);
    outputs(3874) <= layer6_outputs(42);
    outputs(3875) <= (layer6_outputs(1235)) or (layer6_outputs(4333));
    outputs(3876) <= not((layer6_outputs(2263)) or (layer6_outputs(1216)));
    outputs(3877) <= layer6_outputs(4071);
    outputs(3878) <= not(layer6_outputs(5064));
    outputs(3879) <= not(layer6_outputs(4708));
    outputs(3880) <= layer6_outputs(4257);
    outputs(3881) <= layer6_outputs(1733);
    outputs(3882) <= layer6_outputs(2561);
    outputs(3883) <= not(layer6_outputs(3769));
    outputs(3884) <= not(layer6_outputs(2894)) or (layer6_outputs(910));
    outputs(3885) <= layer6_outputs(2460);
    outputs(3886) <= not((layer6_outputs(3292)) or (layer6_outputs(1599)));
    outputs(3887) <= not(layer6_outputs(1396));
    outputs(3888) <= not((layer6_outputs(2031)) xor (layer6_outputs(1054)));
    outputs(3889) <= not(layer6_outputs(3362));
    outputs(3890) <= not((layer6_outputs(1246)) xor (layer6_outputs(1422)));
    outputs(3891) <= layer6_outputs(0);
    outputs(3892) <= layer6_outputs(3479);
    outputs(3893) <= not((layer6_outputs(1801)) xor (layer6_outputs(2822)));
    outputs(3894) <= not((layer6_outputs(2846)) xor (layer6_outputs(368)));
    outputs(3895) <= layer6_outputs(1401);
    outputs(3896) <= (layer6_outputs(2689)) xor (layer6_outputs(1766));
    outputs(3897) <= layer6_outputs(4375);
    outputs(3898) <= (layer6_outputs(1319)) xor (layer6_outputs(4983));
    outputs(3899) <= not(layer6_outputs(1193));
    outputs(3900) <= layer6_outputs(832);
    outputs(3901) <= not(layer6_outputs(2171));
    outputs(3902) <= layer6_outputs(2358);
    outputs(3903) <= not((layer6_outputs(1781)) xor (layer6_outputs(549)));
    outputs(3904) <= layer6_outputs(940);
    outputs(3905) <= not((layer6_outputs(4278)) xor (layer6_outputs(2726)));
    outputs(3906) <= not(layer6_outputs(4118));
    outputs(3907) <= (layer6_outputs(3852)) and not (layer6_outputs(4893));
    outputs(3908) <= layer6_outputs(2602);
    outputs(3909) <= not(layer6_outputs(1172));
    outputs(3910) <= (layer6_outputs(4405)) and not (layer6_outputs(4070));
    outputs(3911) <= not((layer6_outputs(1684)) xor (layer6_outputs(3823)));
    outputs(3912) <= not((layer6_outputs(2928)) xor (layer6_outputs(1334)));
    outputs(3913) <= not(layer6_outputs(1100));
    outputs(3914) <= not((layer6_outputs(1000)) xor (layer6_outputs(4702)));
    outputs(3915) <= not(layer6_outputs(1071));
    outputs(3916) <= (layer6_outputs(4837)) xor (layer6_outputs(4568));
    outputs(3917) <= not(layer6_outputs(1345));
    outputs(3918) <= not((layer6_outputs(2548)) or (layer6_outputs(2371)));
    outputs(3919) <= not(layer6_outputs(961));
    outputs(3920) <= not(layer6_outputs(4555));
    outputs(3921) <= (layer6_outputs(102)) and not (layer6_outputs(1413));
    outputs(3922) <= not(layer6_outputs(1494));
    outputs(3923) <= layer6_outputs(3611);
    outputs(3924) <= layer6_outputs(837);
    outputs(3925) <= (layer6_outputs(543)) xor (layer6_outputs(3669));
    outputs(3926) <= layer6_outputs(2790);
    outputs(3927) <= layer6_outputs(1507);
    outputs(3928) <= (layer6_outputs(3810)) and (layer6_outputs(3874));
    outputs(3929) <= (layer6_outputs(2057)) and not (layer6_outputs(2684));
    outputs(3930) <= not((layer6_outputs(2584)) xor (layer6_outputs(2177)));
    outputs(3931) <= layer6_outputs(1650);
    outputs(3932) <= not((layer6_outputs(2173)) xor (layer6_outputs(4778)));
    outputs(3933) <= not((layer6_outputs(1655)) xor (layer6_outputs(371)));
    outputs(3934) <= not(layer6_outputs(4177));
    outputs(3935) <= not(layer6_outputs(4463));
    outputs(3936) <= not(layer6_outputs(1029));
    outputs(3937) <= layer6_outputs(4478);
    outputs(3938) <= layer6_outputs(3738);
    outputs(3939) <= not((layer6_outputs(3625)) xor (layer6_outputs(3846)));
    outputs(3940) <= not((layer6_outputs(1019)) xor (layer6_outputs(512)));
    outputs(3941) <= not(layer6_outputs(4081));
    outputs(3942) <= (layer6_outputs(3303)) and not (layer6_outputs(5026));
    outputs(3943) <= (layer6_outputs(1997)) and not (layer6_outputs(3897));
    outputs(3944) <= layer6_outputs(258);
    outputs(3945) <= not((layer6_outputs(2975)) xor (layer6_outputs(4561)));
    outputs(3946) <= layer6_outputs(2694);
    outputs(3947) <= not(layer6_outputs(737));
    outputs(3948) <= layer6_outputs(3952);
    outputs(3949) <= (layer6_outputs(1671)) and not (layer6_outputs(196));
    outputs(3950) <= layer6_outputs(3480);
    outputs(3951) <= layer6_outputs(3654);
    outputs(3952) <= layer6_outputs(3637);
    outputs(3953) <= layer6_outputs(424);
    outputs(3954) <= not(layer6_outputs(2520));
    outputs(3955) <= not(layer6_outputs(3027));
    outputs(3956) <= layer6_outputs(3694);
    outputs(3957) <= layer6_outputs(2402);
    outputs(3958) <= not(layer6_outputs(3192));
    outputs(3959) <= layer6_outputs(2848);
    outputs(3960) <= (layer6_outputs(4727)) and not (layer6_outputs(3102));
    outputs(3961) <= not((layer6_outputs(3104)) xor (layer6_outputs(2736)));
    outputs(3962) <= not(layer6_outputs(4267));
    outputs(3963) <= not(layer6_outputs(261));
    outputs(3964) <= layer6_outputs(1903);
    outputs(3965) <= (layer6_outputs(283)) xor (layer6_outputs(1699));
    outputs(3966) <= layer6_outputs(4655);
    outputs(3967) <= layer6_outputs(4146);
    outputs(3968) <= (layer6_outputs(1736)) xor (layer6_outputs(3518));
    outputs(3969) <= layer6_outputs(2793);
    outputs(3970) <= not(layer6_outputs(2850));
    outputs(3971) <= not(layer6_outputs(1223));
    outputs(3972) <= (layer6_outputs(565)) and not (layer6_outputs(3083));
    outputs(3973) <= not(layer6_outputs(3630));
    outputs(3974) <= layer6_outputs(4178);
    outputs(3975) <= not(layer6_outputs(2029));
    outputs(3976) <= (layer6_outputs(1399)) xor (layer6_outputs(4270));
    outputs(3977) <= layer6_outputs(364);
    outputs(3978) <= layer6_outputs(4075);
    outputs(3979) <= (layer6_outputs(3719)) xor (layer6_outputs(2842));
    outputs(3980) <= not(layer6_outputs(3629));
    outputs(3981) <= not(layer6_outputs(1016));
    outputs(3982) <= layer6_outputs(1805);
    outputs(3983) <= (layer6_outputs(5074)) and not (layer6_outputs(3334));
    outputs(3984) <= layer6_outputs(231);
    outputs(3985) <= not(layer6_outputs(2410));
    outputs(3986) <= not(layer6_outputs(2354));
    outputs(3987) <= not(layer6_outputs(1158)) or (layer6_outputs(734));
    outputs(3988) <= layer6_outputs(1035);
    outputs(3989) <= not((layer6_outputs(4646)) or (layer6_outputs(770)));
    outputs(3990) <= (layer6_outputs(4255)) and not (layer6_outputs(2119));
    outputs(3991) <= layer6_outputs(2025);
    outputs(3992) <= not(layer6_outputs(702));
    outputs(3993) <= layer6_outputs(2682);
    outputs(3994) <= not(layer6_outputs(1530));
    outputs(3995) <= (layer6_outputs(436)) xor (layer6_outputs(3159));
    outputs(3996) <= not((layer6_outputs(4053)) xor (layer6_outputs(5005)));
    outputs(3997) <= layer6_outputs(4561);
    outputs(3998) <= not(layer6_outputs(3735));
    outputs(3999) <= layer6_outputs(412);
    outputs(4000) <= layer6_outputs(4342);
    outputs(4001) <= not(layer6_outputs(2348));
    outputs(4002) <= layer6_outputs(397);
    outputs(4003) <= not((layer6_outputs(1158)) and (layer6_outputs(3526)));
    outputs(4004) <= layer6_outputs(1772);
    outputs(4005) <= (layer6_outputs(3297)) xor (layer6_outputs(4037));
    outputs(4006) <= not(layer6_outputs(520));
    outputs(4007) <= (layer6_outputs(4648)) and not (layer6_outputs(285));
    outputs(4008) <= not(layer6_outputs(1541));
    outputs(4009) <= not(layer6_outputs(4021));
    outputs(4010) <= (layer6_outputs(4399)) and not (layer6_outputs(4336));
    outputs(4011) <= not((layer6_outputs(749)) and (layer6_outputs(4719)));
    outputs(4012) <= (layer6_outputs(362)) or (layer6_outputs(3753));
    outputs(4013) <= not(layer6_outputs(1591)) or (layer6_outputs(4688));
    outputs(4014) <= not(layer6_outputs(2990));
    outputs(4015) <= not(layer6_outputs(4327));
    outputs(4016) <= (layer6_outputs(4296)) and not (layer6_outputs(4445));
    outputs(4017) <= (layer6_outputs(117)) xor (layer6_outputs(3380));
    outputs(4018) <= not(layer6_outputs(1946));
    outputs(4019) <= layer6_outputs(1574);
    outputs(4020) <= not(layer6_outputs(2440));
    outputs(4021) <= not(layer6_outputs(3923));
    outputs(4022) <= layer6_outputs(611);
    outputs(4023) <= not(layer6_outputs(3860)) or (layer6_outputs(316));
    outputs(4024) <= not((layer6_outputs(1655)) xor (layer6_outputs(3720)));
    outputs(4025) <= not((layer6_outputs(3882)) xor (layer6_outputs(1529)));
    outputs(4026) <= not(layer6_outputs(814));
    outputs(4027) <= not(layer6_outputs(1212));
    outputs(4028) <= layer6_outputs(2512);
    outputs(4029) <= not(layer6_outputs(1055));
    outputs(4030) <= not(layer6_outputs(1950));
    outputs(4031) <= not((layer6_outputs(2948)) xor (layer6_outputs(2336)));
    outputs(4032) <= not((layer6_outputs(193)) or (layer6_outputs(153)));
    outputs(4033) <= layer6_outputs(3981);
    outputs(4034) <= layer6_outputs(1483);
    outputs(4035) <= layer6_outputs(1469);
    outputs(4036) <= not((layer6_outputs(4354)) xor (layer6_outputs(438)));
    outputs(4037) <= layer6_outputs(3712);
    outputs(4038) <= not(layer6_outputs(3940));
    outputs(4039) <= (layer6_outputs(1426)) and (layer6_outputs(705));
    outputs(4040) <= (layer6_outputs(2923)) and (layer6_outputs(1117));
    outputs(4041) <= layer6_outputs(2954);
    outputs(4042) <= (layer6_outputs(3170)) and (layer6_outputs(2670));
    outputs(4043) <= (layer6_outputs(4892)) xor (layer6_outputs(1710));
    outputs(4044) <= not((layer6_outputs(805)) xor (layer6_outputs(3379)));
    outputs(4045) <= layer6_outputs(4931);
    outputs(4046) <= not(layer6_outputs(1808));
    outputs(4047) <= not(layer6_outputs(3283));
    outputs(4048) <= layer6_outputs(388);
    outputs(4049) <= layer6_outputs(3857);
    outputs(4050) <= layer6_outputs(3888);
    outputs(4051) <= layer6_outputs(2132);
    outputs(4052) <= not((layer6_outputs(194)) or (layer6_outputs(554)));
    outputs(4053) <= layer6_outputs(238);
    outputs(4054) <= not((layer6_outputs(2349)) or (layer6_outputs(1517)));
    outputs(4055) <= not(layer6_outputs(3473)) or (layer6_outputs(96));
    outputs(4056) <= layer6_outputs(681);
    outputs(4057) <= (layer6_outputs(4866)) and (layer6_outputs(4360));
    outputs(4058) <= not(layer6_outputs(4264));
    outputs(4059) <= layer6_outputs(4291);
    outputs(4060) <= not(layer6_outputs(1053));
    outputs(4061) <= layer6_outputs(2211);
    outputs(4062) <= layer6_outputs(2721);
    outputs(4063) <= layer6_outputs(4616);
    outputs(4064) <= not(layer6_outputs(4570));
    outputs(4065) <= not(layer6_outputs(984));
    outputs(4066) <= layer6_outputs(3851);
    outputs(4067) <= (layer6_outputs(1835)) xor (layer6_outputs(995));
    outputs(4068) <= layer6_outputs(3739);
    outputs(4069) <= (layer6_outputs(2694)) and not (layer6_outputs(3474));
    outputs(4070) <= (layer6_outputs(1914)) xor (layer6_outputs(5018));
    outputs(4071) <= not(layer6_outputs(2491));
    outputs(4072) <= (layer6_outputs(5024)) and not (layer6_outputs(1140));
    outputs(4073) <= not((layer6_outputs(2590)) xor (layer6_outputs(3258)));
    outputs(4074) <= (layer6_outputs(2533)) xor (layer6_outputs(4909));
    outputs(4075) <= not(layer6_outputs(1582));
    outputs(4076) <= not(layer6_outputs(1635));
    outputs(4077) <= (layer6_outputs(1897)) and not (layer6_outputs(2517));
    outputs(4078) <= (layer6_outputs(1954)) and not (layer6_outputs(2893));
    outputs(4079) <= not(layer6_outputs(4214));
    outputs(4080) <= not(layer6_outputs(2032));
    outputs(4081) <= layer6_outputs(1869);
    outputs(4082) <= not((layer6_outputs(3366)) xor (layer6_outputs(1775)));
    outputs(4083) <= layer6_outputs(1650);
    outputs(4084) <= (layer6_outputs(218)) and not (layer6_outputs(828));
    outputs(4085) <= not(layer6_outputs(2494));
    outputs(4086) <= layer6_outputs(4109);
    outputs(4087) <= not(layer6_outputs(1487));
    outputs(4088) <= not((layer6_outputs(2243)) xor (layer6_outputs(4683)));
    outputs(4089) <= not(layer6_outputs(2256));
    outputs(4090) <= layer6_outputs(2752);
    outputs(4091) <= layer6_outputs(4196);
    outputs(4092) <= layer6_outputs(93);
    outputs(4093) <= not(layer6_outputs(2941));
    outputs(4094) <= not(layer6_outputs(306));
    outputs(4095) <= not(layer6_outputs(4503));
    outputs(4096) <= not((layer6_outputs(623)) and (layer6_outputs(1075)));
    outputs(4097) <= (layer6_outputs(4502)) and not (layer6_outputs(2162));
    outputs(4098) <= layer6_outputs(3404);
    outputs(4099) <= layer6_outputs(3113);
    outputs(4100) <= not((layer6_outputs(2335)) xor (layer6_outputs(3745)));
    outputs(4101) <= layer6_outputs(384);
    outputs(4102) <= layer6_outputs(2557);
    outputs(4103) <= not(layer6_outputs(2196)) or (layer6_outputs(1981));
    outputs(4104) <= (layer6_outputs(4585)) xor (layer6_outputs(4220));
    outputs(4105) <= not((layer6_outputs(2261)) xor (layer6_outputs(1074)));
    outputs(4106) <= not(layer6_outputs(82));
    outputs(4107) <= not(layer6_outputs(3161));
    outputs(4108) <= layer6_outputs(5085);
    outputs(4109) <= not(layer6_outputs(1027));
    outputs(4110) <= (layer6_outputs(1101)) xor (layer6_outputs(1180));
    outputs(4111) <= not(layer6_outputs(4031));
    outputs(4112) <= not(layer6_outputs(5015));
    outputs(4113) <= not(layer6_outputs(4930)) or (layer6_outputs(484));
    outputs(4114) <= not(layer6_outputs(431));
    outputs(4115) <= not(layer6_outputs(1651));
    outputs(4116) <= layer6_outputs(4357);
    outputs(4117) <= not((layer6_outputs(2680)) xor (layer6_outputs(5113)));
    outputs(4118) <= not(layer6_outputs(4712));
    outputs(4119) <= layer6_outputs(732);
    outputs(4120) <= layer6_outputs(5031);
    outputs(4121) <= not((layer6_outputs(4675)) xor (layer6_outputs(1485)));
    outputs(4122) <= layer6_outputs(4864);
    outputs(4123) <= not(layer6_outputs(1859));
    outputs(4124) <= layer6_outputs(955);
    outputs(4125) <= not((layer6_outputs(3671)) or (layer6_outputs(755)));
    outputs(4126) <= not((layer6_outputs(2865)) xor (layer6_outputs(3000)));
    outputs(4127) <= not((layer6_outputs(2549)) xor (layer6_outputs(4798)));
    outputs(4128) <= not(layer6_outputs(3328)) or (layer6_outputs(1750));
    outputs(4129) <= layer6_outputs(826);
    outputs(4130) <= not(layer6_outputs(3376));
    outputs(4131) <= (layer6_outputs(1846)) xor (layer6_outputs(4268));
    outputs(4132) <= layer6_outputs(3932);
    outputs(4133) <= not(layer6_outputs(4383));
    outputs(4134) <= (layer6_outputs(1675)) xor (layer6_outputs(342));
    outputs(4135) <= layer6_outputs(889);
    outputs(4136) <= (layer6_outputs(2761)) and (layer6_outputs(766));
    outputs(4137) <= layer6_outputs(3088);
    outputs(4138) <= not((layer6_outputs(4083)) xor (layer6_outputs(1263)));
    outputs(4139) <= layer6_outputs(3603);
    outputs(4140) <= layer6_outputs(4921);
    outputs(4141) <= (layer6_outputs(2931)) xor (layer6_outputs(1187));
    outputs(4142) <= (layer6_outputs(574)) xor (layer6_outputs(3793));
    outputs(4143) <= (layer6_outputs(869)) xor (layer6_outputs(1274));
    outputs(4144) <= not(layer6_outputs(2179)) or (layer6_outputs(5102));
    outputs(4145) <= not(layer6_outputs(2532));
    outputs(4146) <= layer6_outputs(3643);
    outputs(4147) <= layer6_outputs(930);
    outputs(4148) <= not(layer6_outputs(2438));
    outputs(4149) <= not(layer6_outputs(2789));
    outputs(4150) <= not(layer6_outputs(1155));
    outputs(4151) <= (layer6_outputs(4242)) and not (layer6_outputs(2467));
    outputs(4152) <= (layer6_outputs(4702)) or (layer6_outputs(4233));
    outputs(4153) <= (layer6_outputs(4995)) xor (layer6_outputs(487));
    outputs(4154) <= layer6_outputs(3420);
    outputs(4155) <= layer6_outputs(473);
    outputs(4156) <= not(layer6_outputs(4670)) or (layer6_outputs(4144));
    outputs(4157) <= layer6_outputs(2502);
    outputs(4158) <= (layer6_outputs(4226)) xor (layer6_outputs(3394));
    outputs(4159) <= not(layer6_outputs(4514));
    outputs(4160) <= not(layer6_outputs(4697)) or (layer6_outputs(1793));
    outputs(4161) <= not((layer6_outputs(694)) xor (layer6_outputs(3497)));
    outputs(4162) <= not(layer6_outputs(4392));
    outputs(4163) <= (layer6_outputs(1209)) and not (layer6_outputs(3123));
    outputs(4164) <= not((layer6_outputs(730)) xor (layer6_outputs(3012)));
    outputs(4165) <= layer6_outputs(434);
    outputs(4166) <= not(layer6_outputs(76));
    outputs(4167) <= layer6_outputs(2200);
    outputs(4168) <= (layer6_outputs(3188)) or (layer6_outputs(2262));
    outputs(4169) <= not(layer6_outputs(2804));
    outputs(4170) <= layer6_outputs(39);
    outputs(4171) <= layer6_outputs(779);
    outputs(4172) <= not((layer6_outputs(4871)) xor (layer6_outputs(1106)));
    outputs(4173) <= not(layer6_outputs(2908));
    outputs(4174) <= (layer6_outputs(637)) xor (layer6_outputs(4845));
    outputs(4175) <= not(layer6_outputs(2488));
    outputs(4176) <= not((layer6_outputs(1262)) and (layer6_outputs(2439)));
    outputs(4177) <= not((layer6_outputs(160)) xor (layer6_outputs(2361)));
    outputs(4178) <= (layer6_outputs(1320)) or (layer6_outputs(3815));
    outputs(4179) <= not((layer6_outputs(3758)) xor (layer6_outputs(4966)));
    outputs(4180) <= (layer6_outputs(1795)) xor (layer6_outputs(3353));
    outputs(4181) <= (layer6_outputs(273)) xor (layer6_outputs(2098));
    outputs(4182) <= layer6_outputs(1834);
    outputs(4183) <= layer6_outputs(1282);
    outputs(4184) <= layer6_outputs(3552);
    outputs(4185) <= (layer6_outputs(4991)) xor (layer6_outputs(1683));
    outputs(4186) <= not(layer6_outputs(2074));
    outputs(4187) <= layer6_outputs(2570);
    outputs(4188) <= layer6_outputs(2735);
    outputs(4189) <= not((layer6_outputs(3417)) or (layer6_outputs(4937)));
    outputs(4190) <= not(layer6_outputs(46)) or (layer6_outputs(4047));
    outputs(4191) <= not((layer6_outputs(3513)) xor (layer6_outputs(4925)));
    outputs(4192) <= layer6_outputs(1993);
    outputs(4193) <= not(layer6_outputs(4525));
    outputs(4194) <= not((layer6_outputs(4020)) xor (layer6_outputs(4889)));
    outputs(4195) <= layer6_outputs(4901);
    outputs(4196) <= layer6_outputs(45);
    outputs(4197) <= (layer6_outputs(1408)) and not (layer6_outputs(2777));
    outputs(4198) <= (layer6_outputs(1072)) xor (layer6_outputs(652));
    outputs(4199) <= (layer6_outputs(143)) xor (layer6_outputs(2729));
    outputs(4200) <= layer6_outputs(3775);
    outputs(4201) <= not(layer6_outputs(4823)) or (layer6_outputs(3067));
    outputs(4202) <= not(layer6_outputs(1739));
    outputs(4203) <= layer6_outputs(3305);
    outputs(4204) <= (layer6_outputs(1778)) xor (layer6_outputs(873));
    outputs(4205) <= not(layer6_outputs(4799));
    outputs(4206) <= (layer6_outputs(1221)) xor (layer6_outputs(1248));
    outputs(4207) <= layer6_outputs(3546);
    outputs(4208) <= layer6_outputs(1669);
    outputs(4209) <= not((layer6_outputs(2078)) xor (layer6_outputs(4751)));
    outputs(4210) <= not((layer6_outputs(1119)) or (layer6_outputs(3013)));
    outputs(4211) <= not(layer6_outputs(4969));
    outputs(4212) <= (layer6_outputs(1123)) xor (layer6_outputs(5097));
    outputs(4213) <= (layer6_outputs(3419)) xor (layer6_outputs(798));
    outputs(4214) <= (layer6_outputs(3288)) and not (layer6_outputs(8));
    outputs(4215) <= layer6_outputs(3032);
    outputs(4216) <= not((layer6_outputs(2921)) xor (layer6_outputs(3355)));
    outputs(4217) <= (layer6_outputs(856)) and (layer6_outputs(2907));
    outputs(4218) <= (layer6_outputs(3412)) xor (layer6_outputs(2890));
    outputs(4219) <= not(layer6_outputs(2573));
    outputs(4220) <= layer6_outputs(253);
    outputs(4221) <= layer6_outputs(1274);
    outputs(4222) <= not(layer6_outputs(1839));
    outputs(4223) <= not((layer6_outputs(4828)) xor (layer6_outputs(367)));
    outputs(4224) <= not(layer6_outputs(2091));
    outputs(4225) <= not((layer6_outputs(785)) xor (layer6_outputs(5006)));
    outputs(4226) <= not(layer6_outputs(506));
    outputs(4227) <= not((layer6_outputs(2833)) xor (layer6_outputs(4397)));
    outputs(4228) <= not((layer6_outputs(2131)) and (layer6_outputs(1614)));
    outputs(4229) <= layer6_outputs(4429);
    outputs(4230) <= (layer6_outputs(4145)) xor (layer6_outputs(3487));
    outputs(4231) <= layer6_outputs(1259);
    outputs(4232) <= layer6_outputs(818);
    outputs(4233) <= not(layer6_outputs(4617));
    outputs(4234) <= not(layer6_outputs(194));
    outputs(4235) <= not((layer6_outputs(3096)) and (layer6_outputs(3132)));
    outputs(4236) <= not((layer6_outputs(2774)) xor (layer6_outputs(4117)));
    outputs(4237) <= not(layer6_outputs(3540));
    outputs(4238) <= not(layer6_outputs(3369));
    outputs(4239) <= not(layer6_outputs(5108));
    outputs(4240) <= not((layer6_outputs(1159)) and (layer6_outputs(618)));
    outputs(4241) <= not((layer6_outputs(634)) and (layer6_outputs(2228)));
    outputs(4242) <= (layer6_outputs(4211)) and not (layer6_outputs(996));
    outputs(4243) <= not(layer6_outputs(1342));
    outputs(4244) <= not(layer6_outputs(1002));
    outputs(4245) <= layer6_outputs(4300);
    outputs(4246) <= not(layer6_outputs(1004));
    outputs(4247) <= layer6_outputs(4335);
    outputs(4248) <= (layer6_outputs(805)) xor (layer6_outputs(1168));
    outputs(4249) <= layer6_outputs(2086);
    outputs(4250) <= layer6_outputs(3575);
    outputs(4251) <= layer6_outputs(819);
    outputs(4252) <= (layer6_outputs(3466)) and (layer6_outputs(1851));
    outputs(4253) <= layer6_outputs(4898);
    outputs(4254) <= not(layer6_outputs(1926));
    outputs(4255) <= layer6_outputs(3334);
    outputs(4256) <= layer6_outputs(2324);
    outputs(4257) <= (layer6_outputs(4357)) and not (layer6_outputs(3313));
    outputs(4258) <= (layer6_outputs(4133)) xor (layer6_outputs(1012));
    outputs(4259) <= not(layer6_outputs(3442));
    outputs(4260) <= (layer6_outputs(4418)) and not (layer6_outputs(885));
    outputs(4261) <= not((layer6_outputs(2930)) and (layer6_outputs(1081)));
    outputs(4262) <= not(layer6_outputs(2683));
    outputs(4263) <= (layer6_outputs(353)) or (layer6_outputs(1336));
    outputs(4264) <= layer6_outputs(3093);
    outputs(4265) <= not(layer6_outputs(3624)) or (layer6_outputs(2913));
    outputs(4266) <= not(layer6_outputs(3831));
    outputs(4267) <= not(layer6_outputs(124));
    outputs(4268) <= not(layer6_outputs(1961));
    outputs(4269) <= layer6_outputs(4733);
    outputs(4270) <= (layer6_outputs(1767)) xor (layer6_outputs(208));
    outputs(4271) <= layer6_outputs(3832);
    outputs(4272) <= layer6_outputs(4709);
    outputs(4273) <= not(layer6_outputs(1129));
    outputs(4274) <= not(layer6_outputs(4684));
    outputs(4275) <= layer6_outputs(3407);
    outputs(4276) <= not(layer6_outputs(4811)) or (layer6_outputs(2603));
    outputs(4277) <= layer6_outputs(2347);
    outputs(4278) <= not(layer6_outputs(5012));
    outputs(4279) <= not(layer6_outputs(2381)) or (layer6_outputs(1421));
    outputs(4280) <= layer6_outputs(4691);
    outputs(4281) <= layer6_outputs(320);
    outputs(4282) <= (layer6_outputs(5010)) xor (layer6_outputs(2193));
    outputs(4283) <= not(layer6_outputs(3515));
    outputs(4284) <= layer6_outputs(2454);
    outputs(4285) <= (layer6_outputs(4513)) xor (layer6_outputs(640));
    outputs(4286) <= not((layer6_outputs(784)) xor (layer6_outputs(3248)));
    outputs(4287) <= (layer6_outputs(3729)) and (layer6_outputs(4618));
    outputs(4288) <= not(layer6_outputs(3863));
    outputs(4289) <= layer6_outputs(1328);
    outputs(4290) <= layer6_outputs(1021);
    outputs(4291) <= not((layer6_outputs(346)) xor (layer6_outputs(3278)));
    outputs(4292) <= not(layer6_outputs(3327));
    outputs(4293) <= not((layer6_outputs(2514)) xor (layer6_outputs(3808)));
    outputs(4294) <= layer6_outputs(2762);
    outputs(4295) <= layer6_outputs(942);
    outputs(4296) <= not((layer6_outputs(3738)) or (layer6_outputs(4668)));
    outputs(4297) <= layer6_outputs(3708);
    outputs(4298) <= layer6_outputs(1756);
    outputs(4299) <= (layer6_outputs(1539)) xor (layer6_outputs(3616));
    outputs(4300) <= not(layer6_outputs(4038));
    outputs(4301) <= layer6_outputs(3965);
    outputs(4302) <= layer6_outputs(3839);
    outputs(4303) <= (layer6_outputs(1844)) xor (layer6_outputs(2794));
    outputs(4304) <= layer6_outputs(1796);
    outputs(4305) <= (layer6_outputs(1732)) xor (layer6_outputs(4790));
    outputs(4306) <= layer6_outputs(4050);
    outputs(4307) <= layer6_outputs(2632);
    outputs(4308) <= layer6_outputs(2493);
    outputs(4309) <= not(layer6_outputs(4130));
    outputs(4310) <= not(layer6_outputs(1668));
    outputs(4311) <= not(layer6_outputs(4663));
    outputs(4312) <= layer6_outputs(3354);
    outputs(4313) <= (layer6_outputs(414)) xor (layer6_outputs(1482));
    outputs(4314) <= not(layer6_outputs(2000));
    outputs(4315) <= not((layer6_outputs(3383)) xor (layer6_outputs(3110)));
    outputs(4316) <= (layer6_outputs(3984)) xor (layer6_outputs(4245));
    outputs(4317) <= layer6_outputs(4210);
    outputs(4318) <= layer6_outputs(469);
    outputs(4319) <= not((layer6_outputs(3202)) and (layer6_outputs(4532)));
    outputs(4320) <= not(layer6_outputs(4152));
    outputs(4321) <= not(layer6_outputs(622));
    outputs(4322) <= layer6_outputs(4122);
    outputs(4323) <= (layer6_outputs(2984)) xor (layer6_outputs(4091));
    outputs(4324) <= not(layer6_outputs(601)) or (layer6_outputs(1006));
    outputs(4325) <= not(layer6_outputs(2157));
    outputs(4326) <= not(layer6_outputs(1643));
    outputs(4327) <= not(layer6_outputs(527));
    outputs(4328) <= layer6_outputs(1442);
    outputs(4329) <= not(layer6_outputs(644));
    outputs(4330) <= (layer6_outputs(1915)) and not (layer6_outputs(2114));
    outputs(4331) <= layer6_outputs(888);
    outputs(4332) <= not(layer6_outputs(4468));
    outputs(4333) <= (layer6_outputs(4991)) xor (layer6_outputs(2182));
    outputs(4334) <= not(layer6_outputs(4244));
    outputs(4335) <= not((layer6_outputs(30)) xor (layer6_outputs(3131)));
    outputs(4336) <= layer6_outputs(4451);
    outputs(4337) <= layer6_outputs(130);
    outputs(4338) <= layer6_outputs(294);
    outputs(4339) <= (layer6_outputs(842)) xor (layer6_outputs(3367));
    outputs(4340) <= not(layer6_outputs(1017));
    outputs(4341) <= layer6_outputs(4582);
    outputs(4342) <= layer6_outputs(1020);
    outputs(4343) <= layer6_outputs(1713);
    outputs(4344) <= layer6_outputs(678);
    outputs(4345) <= layer6_outputs(259);
    outputs(4346) <= not(layer6_outputs(3129));
    outputs(4347) <= layer6_outputs(4527);
    outputs(4348) <= layer6_outputs(1202);
    outputs(4349) <= layer6_outputs(1278);
    outputs(4350) <= not((layer6_outputs(4059)) xor (layer6_outputs(476)));
    outputs(4351) <= not(layer6_outputs(1726));
    outputs(4352) <= layer6_outputs(526);
    outputs(4353) <= layer6_outputs(2443);
    outputs(4354) <= layer6_outputs(3861);
    outputs(4355) <= not(layer6_outputs(4558));
    outputs(4356) <= not((layer6_outputs(1334)) and (layer6_outputs(191)));
    outputs(4357) <= not(layer6_outputs(445)) or (layer6_outputs(3075));
    outputs(4358) <= not(layer6_outputs(2827));
    outputs(4359) <= layer6_outputs(2728);
    outputs(4360) <= layer6_outputs(2980);
    outputs(4361) <= layer6_outputs(4188);
    outputs(4362) <= (layer6_outputs(2510)) and not (layer6_outputs(2130));
    outputs(4363) <= not(layer6_outputs(288));
    outputs(4364) <= (layer6_outputs(863)) and (layer6_outputs(4882));
    outputs(4365) <= (layer6_outputs(783)) xor (layer6_outputs(4099));
    outputs(4366) <= not(layer6_outputs(5111));
    outputs(4367) <= (layer6_outputs(1521)) or (layer6_outputs(3436));
    outputs(4368) <= not(layer6_outputs(3673));
    outputs(4369) <= layer6_outputs(4781);
    outputs(4370) <= (layer6_outputs(548)) xor (layer6_outputs(1543));
    outputs(4371) <= layer6_outputs(3512);
    outputs(4372) <= (layer6_outputs(2466)) xor (layer6_outputs(2444));
    outputs(4373) <= layer6_outputs(1122);
    outputs(4374) <= (layer6_outputs(2258)) xor (layer6_outputs(187));
    outputs(4375) <= (layer6_outputs(2518)) xor (layer6_outputs(3798));
    outputs(4376) <= layer6_outputs(4460);
    outputs(4377) <= not(layer6_outputs(1456));
    outputs(4378) <= layer6_outputs(2907);
    outputs(4379) <= layer6_outputs(750);
    outputs(4380) <= not((layer6_outputs(2286)) xor (layer6_outputs(2468)));
    outputs(4381) <= not(layer6_outputs(4773));
    outputs(4382) <= not(layer6_outputs(1873)) or (layer6_outputs(4679));
    outputs(4383) <= not((layer6_outputs(5098)) xor (layer6_outputs(4760)));
    outputs(4384) <= not(layer6_outputs(4530));
    outputs(4385) <= layer6_outputs(851);
    outputs(4386) <= (layer6_outputs(2507)) xor (layer6_outputs(2953));
    outputs(4387) <= '1';
    outputs(4388) <= (layer6_outputs(529)) xor (layer6_outputs(1830));
    outputs(4389) <= not(layer6_outputs(1705));
    outputs(4390) <= layer6_outputs(2510);
    outputs(4391) <= not(layer6_outputs(4370));
    outputs(4392) <= (layer6_outputs(5020)) and (layer6_outputs(3769));
    outputs(4393) <= (layer6_outputs(4289)) xor (layer6_outputs(2661));
    outputs(4394) <= not(layer6_outputs(2174));
    outputs(4395) <= not(layer6_outputs(3894));
    outputs(4396) <= layer6_outputs(841);
    outputs(4397) <= (layer6_outputs(2167)) xor (layer6_outputs(3166));
    outputs(4398) <= layer6_outputs(790);
    outputs(4399) <= not(layer6_outputs(3602));
    outputs(4400) <= (layer6_outputs(1634)) and not (layer6_outputs(4196));
    outputs(4401) <= layer6_outputs(2311);
    outputs(4402) <= not(layer6_outputs(2946));
    outputs(4403) <= not(layer6_outputs(4742));
    outputs(4404) <= layer6_outputs(4315);
    outputs(4405) <= layer6_outputs(2501);
    outputs(4406) <= layer6_outputs(3592);
    outputs(4407) <= (layer6_outputs(3091)) xor (layer6_outputs(1249));
    outputs(4408) <= layer6_outputs(4013);
    outputs(4409) <= layer6_outputs(3380);
    outputs(4410) <= not((layer6_outputs(1216)) and (layer6_outputs(2775)));
    outputs(4411) <= layer6_outputs(2300);
    outputs(4412) <= not(layer6_outputs(2148));
    outputs(4413) <= not(layer6_outputs(3641));
    outputs(4414) <= (layer6_outputs(3426)) and not (layer6_outputs(72));
    outputs(4415) <= layer6_outputs(2351);
    outputs(4416) <= not(layer6_outputs(148));
    outputs(4417) <= layer6_outputs(150);
    outputs(4418) <= layer6_outputs(491);
    outputs(4419) <= layer6_outputs(3746);
    outputs(4420) <= layer6_outputs(1148);
    outputs(4421) <= not(layer6_outputs(3478));
    outputs(4422) <= layer6_outputs(328);
    outputs(4423) <= (layer6_outputs(2739)) or (layer6_outputs(3080));
    outputs(4424) <= layer6_outputs(2100);
    outputs(4425) <= (layer6_outputs(2971)) xor (layer6_outputs(4002));
    outputs(4426) <= not((layer6_outputs(4119)) xor (layer6_outputs(161)));
    outputs(4427) <= not((layer6_outputs(3213)) and (layer6_outputs(838)));
    outputs(4428) <= not((layer6_outputs(4226)) xor (layer6_outputs(1238)));
    outputs(4429) <= not((layer6_outputs(326)) or (layer6_outputs(3382)));
    outputs(4430) <= layer6_outputs(1382);
    outputs(4431) <= (layer6_outputs(4347)) xor (layer6_outputs(2470));
    outputs(4432) <= not((layer6_outputs(1891)) xor (layer6_outputs(3461)));
    outputs(4433) <= (layer6_outputs(1810)) xor (layer6_outputs(4960));
    outputs(4434) <= (layer6_outputs(2067)) and not (layer6_outputs(4423));
    outputs(4435) <= not(layer6_outputs(4837));
    outputs(4436) <= (layer6_outputs(4508)) xor (layer6_outputs(2851));
    outputs(4437) <= layer6_outputs(4450);
    outputs(4438) <= not(layer6_outputs(2566));
    outputs(4439) <= layer6_outputs(2870);
    outputs(4440) <= (layer6_outputs(432)) xor (layer6_outputs(1641));
    outputs(4441) <= layer6_outputs(5043);
    outputs(4442) <= (layer6_outputs(351)) xor (layer6_outputs(3813));
    outputs(4443) <= not(layer6_outputs(3345));
    outputs(4444) <= not((layer6_outputs(2675)) xor (layer6_outputs(1173)));
    outputs(4445) <= not(layer6_outputs(380));
    outputs(4446) <= layer6_outputs(4077);
    outputs(4447) <= not((layer6_outputs(3893)) xor (layer6_outputs(4130)));
    outputs(4448) <= layer6_outputs(2387);
    outputs(4449) <= layer6_outputs(4246);
    outputs(4450) <= not((layer6_outputs(3102)) or (layer6_outputs(3612)));
    outputs(4451) <= (layer6_outputs(520)) and (layer6_outputs(5020));
    outputs(4452) <= not(layer6_outputs(2452));
    outputs(4453) <= not(layer6_outputs(2774));
    outputs(4454) <= not((layer6_outputs(2024)) and (layer6_outputs(4478)));
    outputs(4455) <= not(layer6_outputs(2260));
    outputs(4456) <= layer6_outputs(531);
    outputs(4457) <= (layer6_outputs(2937)) xor (layer6_outputs(2718));
    outputs(4458) <= not(layer6_outputs(2384));
    outputs(4459) <= (layer6_outputs(1321)) and not (layer6_outputs(2462));
    outputs(4460) <= (layer6_outputs(3822)) and not (layer6_outputs(3495));
    outputs(4461) <= not(layer6_outputs(2012));
    outputs(4462) <= not(layer6_outputs(2434));
    outputs(4463) <= not((layer6_outputs(4674)) xor (layer6_outputs(4685)));
    outputs(4464) <= layer6_outputs(804);
    outputs(4465) <= layer6_outputs(2527);
    outputs(4466) <= not(layer6_outputs(1364));
    outputs(4467) <= not(layer6_outputs(1613));
    outputs(4468) <= not((layer6_outputs(4544)) xor (layer6_outputs(4560)));
    outputs(4469) <= layer6_outputs(3314);
    outputs(4470) <= layer6_outputs(2061);
    outputs(4471) <= layer6_outputs(114);
    outputs(4472) <= not(layer6_outputs(751));
    outputs(4473) <= not(layer6_outputs(4266));
    outputs(4474) <= not(layer6_outputs(2409)) or (layer6_outputs(4815));
    outputs(4475) <= layer6_outputs(4951);
    outputs(4476) <= layer6_outputs(2244);
    outputs(4477) <= (layer6_outputs(3988)) and not (layer6_outputs(4455));
    outputs(4478) <= not((layer6_outputs(3200)) xor (layer6_outputs(3883)));
    outputs(4479) <= not(layer6_outputs(2947));
    outputs(4480) <= not(layer6_outputs(3679));
    outputs(4481) <= not(layer6_outputs(2131));
    outputs(4482) <= not((layer6_outputs(1288)) xor (layer6_outputs(2170)));
    outputs(4483) <= not((layer6_outputs(3406)) and (layer6_outputs(2686)));
    outputs(4484) <= not(layer6_outputs(4699));
    outputs(4485) <= layer6_outputs(307);
    outputs(4486) <= not(layer6_outputs(4367));
    outputs(4487) <= not(layer6_outputs(4400)) or (layer6_outputs(603));
    outputs(4488) <= layer6_outputs(3672);
    outputs(4489) <= not(layer6_outputs(2565));
    outputs(4490) <= layer6_outputs(2429);
    outputs(4491) <= layer6_outputs(177);
    outputs(4492) <= (layer6_outputs(583)) or (layer6_outputs(1504));
    outputs(4493) <= not(layer6_outputs(3880));
    outputs(4494) <= (layer6_outputs(4844)) xor (layer6_outputs(1917));
    outputs(4495) <= not((layer6_outputs(1228)) xor (layer6_outputs(4982)));
    outputs(4496) <= layer6_outputs(1806);
    outputs(4497) <= layer6_outputs(606);
    outputs(4498) <= (layer6_outputs(590)) xor (layer6_outputs(3464));
    outputs(4499) <= (layer6_outputs(831)) and not (layer6_outputs(2232));
    outputs(4500) <= not(layer6_outputs(2442)) or (layer6_outputs(2014));
    outputs(4501) <= not(layer6_outputs(4165));
    outputs(4502) <= not(layer6_outputs(103));
    outputs(4503) <= (layer6_outputs(4494)) and not (layer6_outputs(3021));
    outputs(4504) <= layer6_outputs(4017);
    outputs(4505) <= layer6_outputs(4994);
    outputs(4506) <= (layer6_outputs(3578)) and not (layer6_outputs(53));
    outputs(4507) <= (layer6_outputs(481)) and not (layer6_outputs(827));
    outputs(4508) <= not((layer6_outputs(1374)) xor (layer6_outputs(7)));
    outputs(4509) <= (layer6_outputs(2821)) xor (layer6_outputs(3174));
    outputs(4510) <= not(layer6_outputs(181));
    outputs(4511) <= (layer6_outputs(1022)) xor (layer6_outputs(608));
    outputs(4512) <= (layer6_outputs(2372)) xor (layer6_outputs(3842));
    outputs(4513) <= not(layer6_outputs(2227));
    outputs(4514) <= layer6_outputs(209);
    outputs(4515) <= layer6_outputs(1076);
    outputs(4516) <= not(layer6_outputs(2110));
    outputs(4517) <= not(layer6_outputs(2483));
    outputs(4518) <= not(layer6_outputs(226));
    outputs(4519) <= layer6_outputs(2450);
    outputs(4520) <= not(layer6_outputs(4216)) or (layer6_outputs(1567));
    outputs(4521) <= not((layer6_outputs(2214)) xor (layer6_outputs(1215)));
    outputs(4522) <= layer6_outputs(5102);
    outputs(4523) <= not(layer6_outputs(2448));
    outputs(4524) <= not((layer6_outputs(1565)) xor (layer6_outputs(2130)));
    outputs(4525) <= layer6_outputs(820);
    outputs(4526) <= (layer6_outputs(2629)) xor (layer6_outputs(2988));
    outputs(4527) <= not(layer6_outputs(3744));
    outputs(4528) <= not(layer6_outputs(4876));
    outputs(4529) <= (layer6_outputs(3946)) xor (layer6_outputs(4806));
    outputs(4530) <= not((layer6_outputs(676)) xor (layer6_outputs(3289)));
    outputs(4531) <= layer6_outputs(3231);
    outputs(4532) <= not((layer6_outputs(957)) and (layer6_outputs(2233)));
    outputs(4533) <= not(layer6_outputs(3061));
    outputs(4534) <= layer6_outputs(3210);
    outputs(4535) <= layer6_outputs(4303);
    outputs(4536) <= layer6_outputs(2017);
    outputs(4537) <= (layer6_outputs(1023)) xor (layer6_outputs(2241));
    outputs(4538) <= layer6_outputs(789);
    outputs(4539) <= not((layer6_outputs(5091)) xor (layer6_outputs(2405)));
    outputs(4540) <= layer6_outputs(4830);
    outputs(4541) <= not(layer6_outputs(1855));
    outputs(4542) <= not(layer6_outputs(4635)) or (layer6_outputs(3463));
    outputs(4543) <= not((layer6_outputs(611)) and (layer6_outputs(1)));
    outputs(4544) <= layer6_outputs(1475);
    outputs(4545) <= layer6_outputs(2578);
    outputs(4546) <= not(layer6_outputs(2932));
    outputs(4547) <= not(layer6_outputs(2012));
    outputs(4548) <= layer6_outputs(2119);
    outputs(4549) <= not(layer6_outputs(2276));
    outputs(4550) <= (layer6_outputs(4619)) xor (layer6_outputs(5091));
    outputs(4551) <= not(layer6_outputs(1326));
    outputs(4552) <= not((layer6_outputs(920)) xor (layer6_outputs(375)));
    outputs(4553) <= not(layer6_outputs(1811));
    outputs(4554) <= not((layer6_outputs(2993)) and (layer6_outputs(2982)));
    outputs(4555) <= layer6_outputs(2036);
    outputs(4556) <= (layer6_outputs(448)) xor (layer6_outputs(1678));
    outputs(4557) <= not(layer6_outputs(2509));
    outputs(4558) <= not(layer6_outputs(2152));
    outputs(4559) <= not(layer6_outputs(4707));
    outputs(4560) <= (layer6_outputs(3163)) and not (layer6_outputs(43));
    outputs(4561) <= layer6_outputs(505);
    outputs(4562) <= layer6_outputs(192);
    outputs(4563) <= layer6_outputs(5087);
    outputs(4564) <= (layer6_outputs(908)) and (layer6_outputs(150));
    outputs(4565) <= not(layer6_outputs(1651));
    outputs(4566) <= not(layer6_outputs(4831));
    outputs(4567) <= not(layer6_outputs(3121));
    outputs(4568) <= not((layer6_outputs(4361)) or (layer6_outputs(2366)));
    outputs(4569) <= not((layer6_outputs(3754)) xor (layer6_outputs(2045)));
    outputs(4570) <= not(layer6_outputs(736));
    outputs(4571) <= layer6_outputs(4114);
    outputs(4572) <= layer6_outputs(4371);
    outputs(4573) <= layer6_outputs(4106);
    outputs(4574) <= (layer6_outputs(1169)) and (layer6_outputs(2653));
    outputs(4575) <= not(layer6_outputs(4076));
    outputs(4576) <= (layer6_outputs(2729)) xor (layer6_outputs(3826));
    outputs(4577) <= (layer6_outputs(1331)) and not (layer6_outputs(1605));
    outputs(4578) <= not((layer6_outputs(1261)) or (layer6_outputs(2863)));
    outputs(4579) <= layer6_outputs(4864);
    outputs(4580) <= not(layer6_outputs(4501));
    outputs(4581) <= layer6_outputs(2640);
    outputs(4582) <= layer6_outputs(3393);
    outputs(4583) <= not(layer6_outputs(2038));
    outputs(4584) <= layer6_outputs(2898);
    outputs(4585) <= (layer6_outputs(540)) xor (layer6_outputs(978));
    outputs(4586) <= not(layer6_outputs(753));
    outputs(4587) <= layer6_outputs(2996);
    outputs(4588) <= layer6_outputs(4084);
    outputs(4589) <= layer6_outputs(2435);
    outputs(4590) <= layer6_outputs(2224);
    outputs(4591) <= not(layer6_outputs(731));
    outputs(4592) <= not((layer6_outputs(2891)) xor (layer6_outputs(3961)));
    outputs(4593) <= not(layer6_outputs(3405));
    outputs(4594) <= not((layer6_outputs(4175)) and (layer6_outputs(2495)));
    outputs(4595) <= not((layer6_outputs(1693)) and (layer6_outputs(1327)));
    outputs(4596) <= not((layer6_outputs(2329)) xor (layer6_outputs(2428)));
    outputs(4597) <= not((layer6_outputs(156)) and (layer6_outputs(3381)));
    outputs(4598) <= (layer6_outputs(4104)) xor (layer6_outputs(3143));
    outputs(4599) <= not(layer6_outputs(1057));
    outputs(4600) <= layer6_outputs(4467);
    outputs(4601) <= not(layer6_outputs(2573));
    outputs(4602) <= not(layer6_outputs(3451));
    outputs(4603) <= not(layer6_outputs(344));
    outputs(4604) <= not(layer6_outputs(4153));
    outputs(4605) <= not(layer6_outputs(4713));
    outputs(4606) <= not(layer6_outputs(3919));
    outputs(4607) <= not((layer6_outputs(2390)) xor (layer6_outputs(743)));
    outputs(4608) <= not(layer6_outputs(3185));
    outputs(4609) <= layer6_outputs(3223);
    outputs(4610) <= not(layer6_outputs(4482));
    outputs(4611) <= not(layer6_outputs(4005));
    outputs(4612) <= not((layer6_outputs(2979)) xor (layer6_outputs(1573)));
    outputs(4613) <= not(layer6_outputs(2048));
    outputs(4614) <= not(layer6_outputs(3534));
    outputs(4615) <= not(layer6_outputs(4055));
    outputs(4616) <= not(layer6_outputs(739));
    outputs(4617) <= layer6_outputs(1632);
    outputs(4618) <= not((layer6_outputs(1652)) xor (layer6_outputs(2756)));
    outputs(4619) <= not((layer6_outputs(4470)) xor (layer6_outputs(2319)));
    outputs(4620) <= (layer6_outputs(432)) and not (layer6_outputs(4698));
    outputs(4621) <= layer6_outputs(2568);
    outputs(4622) <= not(layer6_outputs(3068));
    outputs(4623) <= layer6_outputs(4961);
    outputs(4624) <= layer6_outputs(654);
    outputs(4625) <= (layer6_outputs(2462)) and (layer6_outputs(1639));
    outputs(4626) <= not(layer6_outputs(4971));
    outputs(4627) <= not(layer6_outputs(2605));
    outputs(4628) <= (layer6_outputs(3137)) xor (layer6_outputs(3789));
    outputs(4629) <= layer6_outputs(3155);
    outputs(4630) <= (layer6_outputs(4790)) xor (layer6_outputs(4688));
    outputs(4631) <= layer6_outputs(3039);
    outputs(4632) <= not((layer6_outputs(718)) xor (layer6_outputs(1837)));
    outputs(4633) <= not(layer6_outputs(3563));
    outputs(4634) <= not((layer6_outputs(4608)) xor (layer6_outputs(1230)));
    outputs(4635) <= not((layer6_outputs(2277)) xor (layer6_outputs(1571)));
    outputs(4636) <= not(layer6_outputs(163));
    outputs(4637) <= not(layer6_outputs(939));
    outputs(4638) <= layer6_outputs(4101);
    outputs(4639) <= layer6_outputs(2610);
    outputs(4640) <= not((layer6_outputs(3059)) xor (layer6_outputs(2220)));
    outputs(4641) <= not((layer6_outputs(3624)) xor (layer6_outputs(1205)));
    outputs(4642) <= (layer6_outputs(1368)) or (layer6_outputs(1473));
    outputs(4643) <= not(layer6_outputs(1433));
    outputs(4644) <= layer6_outputs(3618);
    outputs(4645) <= layer6_outputs(4784);
    outputs(4646) <= not(layer6_outputs(3621));
    outputs(4647) <= not(layer6_outputs(2540));
    outputs(4648) <= not(layer6_outputs(3326)) or (layer6_outputs(3205));
    outputs(4649) <= layer6_outputs(4710);
    outputs(4650) <= (layer6_outputs(2073)) and not (layer6_outputs(822));
    outputs(4651) <= not(layer6_outputs(550));
    outputs(4652) <= (layer6_outputs(1662)) and (layer6_outputs(1719));
    outputs(4653) <= not(layer6_outputs(612));
    outputs(4654) <= not(layer6_outputs(2522));
    outputs(4655) <= not(layer6_outputs(5031));
    outputs(4656) <= layer6_outputs(4651);
    outputs(4657) <= not(layer6_outputs(563));
    outputs(4658) <= (layer6_outputs(3499)) and not (layer6_outputs(2997));
    outputs(4659) <= not(layer6_outputs(4453));
    outputs(4660) <= layer6_outputs(1126);
    outputs(4661) <= layer6_outputs(4552);
    outputs(4662) <= not(layer6_outputs(4640));
    outputs(4663) <= layer6_outputs(1638);
    outputs(4664) <= not(layer6_outputs(2874));
    outputs(4665) <= not(layer6_outputs(4782));
    outputs(4666) <= (layer6_outputs(5116)) or (layer6_outputs(1865));
    outputs(4667) <= (layer6_outputs(313)) and not (layer6_outputs(2741));
    outputs(4668) <= not(layer6_outputs(3703));
    outputs(4669) <= not((layer6_outputs(175)) xor (layer6_outputs(845)));
    outputs(4670) <= layer6_outputs(4157);
    outputs(4671) <= not(layer6_outputs(564));
    outputs(4672) <= (layer6_outputs(5067)) xor (layer6_outputs(1812));
    outputs(4673) <= not(layer6_outputs(3595));
    outputs(4674) <= not(layer6_outputs(2962));
    outputs(4675) <= (layer6_outputs(1408)) xor (layer6_outputs(464));
    outputs(4676) <= layer6_outputs(1125);
    outputs(4677) <= layer6_outputs(4870);
    outputs(4678) <= layer6_outputs(4535);
    outputs(4679) <= not(layer6_outputs(5088));
    outputs(4680) <= not((layer6_outputs(4976)) xor (layer6_outputs(3957)));
    outputs(4681) <= not((layer6_outputs(2356)) xor (layer6_outputs(3458)));
    outputs(4682) <= layer6_outputs(466);
    outputs(4683) <= (layer6_outputs(442)) xor (layer6_outputs(1387));
    outputs(4684) <= not((layer6_outputs(2513)) xor (layer6_outputs(333)));
    outputs(4685) <= not((layer6_outputs(2195)) xor (layer6_outputs(679)));
    outputs(4686) <= not((layer6_outputs(853)) or (layer6_outputs(1291)));
    outputs(4687) <= layer6_outputs(2752);
    outputs(4688) <= layer6_outputs(3235);
    outputs(4689) <= layer6_outputs(1415);
    outputs(4690) <= layer6_outputs(4191);
    outputs(4691) <= not(layer6_outputs(5038));
    outputs(4692) <= not((layer6_outputs(4427)) xor (layer6_outputs(4194)));
    outputs(4693) <= not(layer6_outputs(132));
    outputs(4694) <= not(layer6_outputs(2465));
    outputs(4695) <= layer6_outputs(291);
    outputs(4696) <= not(layer6_outputs(1599));
    outputs(4697) <= layer6_outputs(1083);
    outputs(4698) <= not(layer6_outputs(203));
    outputs(4699) <= layer6_outputs(3619);
    outputs(4700) <= (layer6_outputs(2385)) xor (layer6_outputs(4801));
    outputs(4701) <= layer6_outputs(1762);
    outputs(4702) <= not(layer6_outputs(588));
    outputs(4703) <= layer6_outputs(4472);
    outputs(4704) <= (layer6_outputs(2389)) and not (layer6_outputs(4426));
    outputs(4705) <= layer6_outputs(5003);
    outputs(4706) <= not(layer6_outputs(13));
    outputs(4707) <= not(layer6_outputs(4862));
    outputs(4708) <= not(layer6_outputs(3559));
    outputs(4709) <= not(layer6_outputs(3086));
    outputs(4710) <= layer6_outputs(3023);
    outputs(4711) <= (layer6_outputs(675)) xor (layer6_outputs(1118));
    outputs(4712) <= layer6_outputs(2008);
    outputs(4713) <= layer6_outputs(4622);
    outputs(4714) <= not(layer6_outputs(4024));
    outputs(4715) <= (layer6_outputs(3080)) and not (layer6_outputs(4464));
    outputs(4716) <= not(layer6_outputs(1338));
    outputs(4717) <= layer6_outputs(890);
    outputs(4718) <= (layer6_outputs(2112)) xor (layer6_outputs(3660));
    outputs(4719) <= (layer6_outputs(4510)) and not (layer6_outputs(4777));
    outputs(4720) <= not((layer6_outputs(3990)) and (layer6_outputs(514)));
    outputs(4721) <= not(layer6_outputs(2223));
    outputs(4722) <= layer6_outputs(2181);
    outputs(4723) <= not((layer6_outputs(665)) xor (layer6_outputs(4134)));
    outputs(4724) <= layer6_outputs(4377);
    outputs(4725) <= layer6_outputs(2853);
    outputs(4726) <= not((layer6_outputs(1528)) xor (layer6_outputs(4802)));
    outputs(4727) <= (layer6_outputs(1156)) xor (layer6_outputs(3650));
    outputs(4728) <= (layer6_outputs(408)) and not (layer6_outputs(2285));
    outputs(4729) <= not((layer6_outputs(1538)) xor (layer6_outputs(284)));
    outputs(4730) <= layer6_outputs(960);
    outputs(4731) <= layer6_outputs(2778);
    outputs(4732) <= layer6_outputs(4261);
    outputs(4733) <= layer6_outputs(3148);
    outputs(4734) <= (layer6_outputs(1162)) xor (layer6_outputs(3983));
    outputs(4735) <= layer6_outputs(900);
    outputs(4736) <= not(layer6_outputs(4302));
    outputs(4737) <= layer6_outputs(3278);
    outputs(4738) <= not(layer6_outputs(3057));
    outputs(4739) <= layer6_outputs(2499);
    outputs(4740) <= (layer6_outputs(135)) xor (layer6_outputs(4229));
    outputs(4741) <= not(layer6_outputs(926));
    outputs(4742) <= (layer6_outputs(848)) and not (layer6_outputs(3212));
    outputs(4743) <= (layer6_outputs(395)) and not (layer6_outputs(4623));
    outputs(4744) <= (layer6_outputs(4271)) and not (layer6_outputs(3605));
    outputs(4745) <= not(layer6_outputs(1044));
    outputs(4746) <= (layer6_outputs(4086)) xor (layer6_outputs(3645));
    outputs(4747) <= layer6_outputs(238);
    outputs(4748) <= layer6_outputs(774);
    outputs(4749) <= layer6_outputs(1406);
    outputs(4750) <= (layer6_outputs(2318)) and not (layer6_outputs(2668));
    outputs(4751) <= not((layer6_outputs(2745)) or (layer6_outputs(4225)));
    outputs(4752) <= not(layer6_outputs(3962));
    outputs(4753) <= not(layer6_outputs(2320));
    outputs(4754) <= not(layer6_outputs(1354));
    outputs(4755) <= layer6_outputs(395);
    outputs(4756) <= (layer6_outputs(5051)) and not (layer6_outputs(3456));
    outputs(4757) <= not((layer6_outputs(930)) xor (layer6_outputs(3346)));
    outputs(4758) <= not(layer6_outputs(1967));
    outputs(4759) <= (layer6_outputs(3063)) xor (layer6_outputs(3161));
    outputs(4760) <= not(layer6_outputs(1064));
    outputs(4761) <= not(layer6_outputs(2272));
    outputs(4762) <= layer6_outputs(243);
    outputs(4763) <= not(layer6_outputs(1213));
    outputs(4764) <= layer6_outputs(4854);
    outputs(4765) <= layer6_outputs(1201);
    outputs(4766) <= not(layer6_outputs(3090)) or (layer6_outputs(2508));
    outputs(4767) <= layer6_outputs(3905);
    outputs(4768) <= layer6_outputs(4703);
    outputs(4769) <= not(layer6_outputs(3569));
    outputs(4770) <= not(layer6_outputs(562));
    outputs(4771) <= not(layer6_outputs(3125)) or (layer6_outputs(2136));
    outputs(4772) <= not(layer6_outputs(3185));
    outputs(4773) <= layer6_outputs(1965);
    outputs(4774) <= (layer6_outputs(1673)) and (layer6_outputs(1872));
    outputs(4775) <= not(layer6_outputs(1111));
    outputs(4776) <= not(layer6_outputs(2494));
    outputs(4777) <= not(layer6_outputs(4568));
    outputs(4778) <= not((layer6_outputs(2637)) xor (layer6_outputs(1603)));
    outputs(4779) <= not(layer6_outputs(167));
    outputs(4780) <= (layer6_outputs(2594)) xor (layer6_outputs(2228));
    outputs(4781) <= layer6_outputs(4407);
    outputs(4782) <= not((layer6_outputs(3214)) or (layer6_outputs(4735)));
    outputs(4783) <= (layer6_outputs(4089)) and not (layer6_outputs(1091));
    outputs(4784) <= not((layer6_outputs(775)) or (layer6_outputs(5117)));
    outputs(4785) <= (layer6_outputs(4543)) xor (layer6_outputs(4915));
    outputs(4786) <= (layer6_outputs(3877)) and (layer6_outputs(1980));
    outputs(4787) <= layer6_outputs(623);
    outputs(4788) <= layer6_outputs(2650);
    outputs(4789) <= layer6_outputs(2954);
    outputs(4790) <= layer6_outputs(4230);
    outputs(4791) <= not(layer6_outputs(672));
    outputs(4792) <= not(layer6_outputs(3647));
    outputs(4793) <= not((layer6_outputs(3465)) xor (layer6_outputs(810)));
    outputs(4794) <= layer6_outputs(3604);
    outputs(4795) <= layer6_outputs(146);
    outputs(4796) <= not(layer6_outputs(1435));
    outputs(4797) <= (layer6_outputs(1277)) and not (layer6_outputs(5022));
    outputs(4798) <= layer6_outputs(2644);
    outputs(4799) <= layer6_outputs(2346);
    outputs(4800) <= layer6_outputs(1972);
    outputs(4801) <= not(layer6_outputs(381));
    outputs(4802) <= (layer6_outputs(886)) xor (layer6_outputs(1951));
    outputs(4803) <= layer6_outputs(356);
    outputs(4804) <= layer6_outputs(2025);
    outputs(4805) <= not(layer6_outputs(2256));
    outputs(4806) <= not(layer6_outputs(3177));
    outputs(4807) <= layer6_outputs(2073);
    outputs(4808) <= (layer6_outputs(1569)) and not (layer6_outputs(6));
    outputs(4809) <= not(layer6_outputs(3520));
    outputs(4810) <= (layer6_outputs(1348)) xor (layer6_outputs(685));
    outputs(4811) <= layer6_outputs(503);
    outputs(4812) <= layer6_outputs(3788);
    outputs(4813) <= (layer6_outputs(2365)) and not (layer6_outputs(3189));
    outputs(4814) <= layer6_outputs(1367);
    outputs(4815) <= not((layer6_outputs(4764)) and (layer6_outputs(1913)));
    outputs(4816) <= not((layer6_outputs(2380)) and (layer6_outputs(3152)));
    outputs(4817) <= not(layer6_outputs(1923));
    outputs(4818) <= layer6_outputs(4273);
    outputs(4819) <= layer6_outputs(3034);
    outputs(4820) <= not(layer6_outputs(1781));
    outputs(4821) <= layer6_outputs(2792);
    outputs(4822) <= not((layer6_outputs(2279)) xor (layer6_outputs(2943)));
    outputs(4823) <= layer6_outputs(1618);
    outputs(4824) <= layer6_outputs(3538);
    outputs(4825) <= (layer6_outputs(1644)) xor (layer6_outputs(4647));
    outputs(4826) <= not(layer6_outputs(731));
    outputs(4827) <= not(layer6_outputs(1024));
    outputs(4828) <= not(layer6_outputs(2883));
    outputs(4829) <= layer6_outputs(2339);
    outputs(4830) <= (layer6_outputs(4178)) and (layer6_outputs(615));
    outputs(4831) <= layer6_outputs(1032);
    outputs(4832) <= not(layer6_outputs(3338));
    outputs(4833) <= (layer6_outputs(223)) xor (layer6_outputs(1804));
    outputs(4834) <= not(layer6_outputs(3993));
    outputs(4835) <= layer6_outputs(1084);
    outputs(4836) <= not((layer6_outputs(1682)) or (layer6_outputs(3642)));
    outputs(4837) <= layer6_outputs(1596);
    outputs(4838) <= not((layer6_outputs(4174)) or (layer6_outputs(803)));
    outputs(4839) <= (layer6_outputs(1155)) xor (layer6_outputs(3386));
    outputs(4840) <= not((layer6_outputs(2807)) xor (layer6_outputs(4390)));
    outputs(4841) <= not(layer6_outputs(2624)) or (layer6_outputs(4907));
    outputs(4842) <= layer6_outputs(2982);
    outputs(4843) <= (layer6_outputs(1107)) and not (layer6_outputs(3807));
    outputs(4844) <= layer6_outputs(4164);
    outputs(4845) <= not(layer6_outputs(3192)) or (layer6_outputs(862));
    outputs(4846) <= not((layer6_outputs(2266)) xor (layer6_outputs(4637)));
    outputs(4847) <= not(layer6_outputs(976));
    outputs(4848) <= not((layer6_outputs(4105)) or (layer6_outputs(3010)));
    outputs(4849) <= not((layer6_outputs(1644)) xor (layer6_outputs(5033)));
    outputs(4850) <= layer6_outputs(1900);
    outputs(4851) <= not((layer6_outputs(1161)) xor (layer6_outputs(3528)));
    outputs(4852) <= layer6_outputs(882);
    outputs(4853) <= not(layer6_outputs(917));
    outputs(4854) <= not(layer6_outputs(3541));
    outputs(4855) <= (layer6_outputs(2538)) xor (layer6_outputs(2222));
    outputs(4856) <= layer6_outputs(4407);
    outputs(4857) <= not((layer6_outputs(5079)) or (layer6_outputs(796)));
    outputs(4858) <= not((layer6_outputs(1717)) and (layer6_outputs(4456)));
    outputs(4859) <= (layer6_outputs(2477)) or (layer6_outputs(3674));
    outputs(4860) <= not(layer6_outputs(3295));
    outputs(4861) <= not(layer6_outputs(4939));
    outputs(4862) <= not(layer6_outputs(4519));
    outputs(4863) <= (layer6_outputs(42)) and not (layer6_outputs(791));
    outputs(4864) <= (layer6_outputs(1323)) xor (layer6_outputs(3469));
    outputs(4865) <= layer6_outputs(4912);
    outputs(4866) <= layer6_outputs(3950);
    outputs(4867) <= not((layer6_outputs(1235)) xor (layer6_outputs(3120)));
    outputs(4868) <= layer6_outputs(159);
    outputs(4869) <= not((layer6_outputs(2856)) xor (layer6_outputs(2939)));
    outputs(4870) <= (layer6_outputs(1472)) and not (layer6_outputs(1806));
    outputs(4871) <= not(layer6_outputs(1355));
    outputs(4872) <= not(layer6_outputs(4754));
    outputs(4873) <= layer6_outputs(3023);
    outputs(4874) <= layer6_outputs(1083);
    outputs(4875) <= not(layer6_outputs(1327));
    outputs(4876) <= not(layer6_outputs(1595)) or (layer6_outputs(2696));
    outputs(4877) <= layer6_outputs(5098);
    outputs(4878) <= layer6_outputs(858);
    outputs(4879) <= layer6_outputs(1839);
    outputs(4880) <= layer6_outputs(417);
    outputs(4881) <= not((layer6_outputs(911)) xor (layer6_outputs(2653)));
    outputs(4882) <= not(layer6_outputs(1488));
    outputs(4883) <= layer6_outputs(3673);
    outputs(4884) <= (layer6_outputs(3183)) and not (layer6_outputs(72));
    outputs(4885) <= not(layer6_outputs(1344));
    outputs(4886) <= layer6_outputs(4322);
    outputs(4887) <= not(layer6_outputs(4158)) or (layer6_outputs(3964));
    outputs(4888) <= (layer6_outputs(4202)) xor (layer6_outputs(3928));
    outputs(4889) <= not((layer6_outputs(5022)) or (layer6_outputs(887)));
    outputs(4890) <= not(layer6_outputs(3097));
    outputs(4891) <= (layer6_outputs(977)) xor (layer6_outputs(3881));
    outputs(4892) <= not((layer6_outputs(884)) xor (layer6_outputs(501)));
    outputs(4893) <= (layer6_outputs(4228)) and not (layer6_outputs(2241));
    outputs(4894) <= not(layer6_outputs(4847));
    outputs(4895) <= not(layer6_outputs(4079));
    outputs(4896) <= (layer6_outputs(1122)) and (layer6_outputs(3527));
    outputs(4897) <= (layer6_outputs(230)) xor (layer6_outputs(3748));
    outputs(4898) <= (layer6_outputs(3447)) and not (layer6_outputs(825));
    outputs(4899) <= (layer6_outputs(2203)) xor (layer6_outputs(3764));
    outputs(4900) <= not(layer6_outputs(4957));
    outputs(4901) <= not(layer6_outputs(1597));
    outputs(4902) <= not(layer6_outputs(651));
    outputs(4903) <= layer6_outputs(3777);
    outputs(4904) <= not(layer6_outputs(208));
    outputs(4905) <= not(layer6_outputs(4248));
    outputs(4906) <= (layer6_outputs(1304)) and not (layer6_outputs(31));
    outputs(4907) <= layer6_outputs(4341);
    outputs(4908) <= not(layer6_outputs(4347));
    outputs(4909) <= layer6_outputs(2867);
    outputs(4910) <= layer6_outputs(304);
    outputs(4911) <= not((layer6_outputs(2747)) xor (layer6_outputs(1393)));
    outputs(4912) <= (layer6_outputs(4263)) xor (layer6_outputs(4235));
    outputs(4913) <= layer6_outputs(4039);
    outputs(4914) <= not(layer6_outputs(2320));
    outputs(4915) <= (layer6_outputs(5007)) xor (layer6_outputs(3677));
    outputs(4916) <= layer6_outputs(2056);
    outputs(4917) <= not(layer6_outputs(2831)) or (layer6_outputs(3787));
    outputs(4918) <= (layer6_outputs(3022)) or (layer6_outputs(1588));
    outputs(4919) <= not(layer6_outputs(741));
    outputs(4920) <= (layer6_outputs(2101)) and (layer6_outputs(158));
    outputs(4921) <= not((layer6_outputs(2857)) xor (layer6_outputs(4200)));
    outputs(4922) <= not(layer6_outputs(1478));
    outputs(4923) <= not((layer6_outputs(1730)) or (layer6_outputs(1747)));
    outputs(4924) <= not(layer6_outputs(5040));
    outputs(4925) <= (layer6_outputs(4457)) xor (layer6_outputs(3617));
    outputs(4926) <= layer6_outputs(4473);
    outputs(4927) <= (layer6_outputs(4630)) and (layer6_outputs(2013));
    outputs(4928) <= layer6_outputs(786);
    outputs(4929) <= layer6_outputs(3717);
    outputs(4930) <= (layer6_outputs(1373)) and not (layer6_outputs(5093));
    outputs(4931) <= layer6_outputs(3347);
    outputs(4932) <= (layer6_outputs(3393)) and not (layer6_outputs(3998));
    outputs(4933) <= (layer6_outputs(525)) and not (layer6_outputs(337));
    outputs(4934) <= layer6_outputs(3489);
    outputs(4935) <= (layer6_outputs(877)) xor (layer6_outputs(466));
    outputs(4936) <= layer6_outputs(4800);
    outputs(4937) <= not((layer6_outputs(1259)) xor (layer6_outputs(4443)));
    outputs(4938) <= not(layer6_outputs(847));
    outputs(4939) <= not((layer6_outputs(1051)) xor (layer6_outputs(4149)));
    outputs(4940) <= not(layer6_outputs(591));
    outputs(4941) <= layer6_outputs(414);
    outputs(4942) <= not(layer6_outputs(4514));
    outputs(4943) <= (layer6_outputs(972)) or (layer6_outputs(425));
    outputs(4944) <= layer6_outputs(900);
    outputs(4945) <= (layer6_outputs(3187)) and not (layer6_outputs(3179));
    outputs(4946) <= not(layer6_outputs(186));
    outputs(4947) <= layer6_outputs(4851);
    outputs(4948) <= not(layer6_outputs(3431)) or (layer6_outputs(4676));
    outputs(4949) <= layer6_outputs(4624);
    outputs(4950) <= layer6_outputs(2355);
    outputs(4951) <= (layer6_outputs(2676)) and (layer6_outputs(892));
    outputs(4952) <= not(layer6_outputs(4621));
    outputs(4953) <= layer6_outputs(3644);
    outputs(4954) <= (layer6_outputs(3855)) and (layer6_outputs(4498));
    outputs(4955) <= layer6_outputs(3506);
    outputs(4956) <= not(layer6_outputs(1722));
    outputs(4957) <= layer6_outputs(1189);
    outputs(4958) <= (layer6_outputs(4873)) and not (layer6_outputs(2317));
    outputs(4959) <= not((layer6_outputs(5066)) xor (layer6_outputs(1539)));
    outputs(4960) <= not((layer6_outputs(2103)) or (layer6_outputs(2273)));
    outputs(4961) <= layer6_outputs(1194);
    outputs(4962) <= not(layer6_outputs(1702));
    outputs(4963) <= layer6_outputs(2109);
    outputs(4964) <= (layer6_outputs(4271)) and not (layer6_outputs(1372));
    outputs(4965) <= not(layer6_outputs(3361)) or (layer6_outputs(1876));
    outputs(4966) <= not(layer6_outputs(553));
    outputs(4967) <= layer6_outputs(4530);
    outputs(4968) <= not(layer6_outputs(2297)) or (layer6_outputs(3814));
    outputs(4969) <= not((layer6_outputs(983)) or (layer6_outputs(2064)));
    outputs(4970) <= not(layer6_outputs(3547));
    outputs(4971) <= not(layer6_outputs(2548));
    outputs(4972) <= not(layer6_outputs(3639));
    outputs(4973) <= layer6_outputs(3802);
    outputs(4974) <= not(layer6_outputs(4181));
    outputs(4975) <= (layer6_outputs(3020)) or (layer6_outputs(2635));
    outputs(4976) <= (layer6_outputs(4070)) and not (layer6_outputs(3807));
    outputs(4977) <= not(layer6_outputs(4903));
    outputs(4978) <= layer6_outputs(911);
    outputs(4979) <= layer6_outputs(5008);
    outputs(4980) <= not((layer6_outputs(2816)) xor (layer6_outputs(3884)));
    outputs(4981) <= layer6_outputs(3073);
    outputs(4982) <= not(layer6_outputs(866));
    outputs(4983) <= not((layer6_outputs(4137)) xor (layer6_outputs(4671)));
    outputs(4984) <= not(layer6_outputs(747));
    outputs(4985) <= (layer6_outputs(3172)) xor (layer6_outputs(2678));
    outputs(4986) <= layer6_outputs(1677);
    outputs(4987) <= (layer6_outputs(1575)) and (layer6_outputs(3514));
    outputs(4988) <= not((layer6_outputs(3045)) xor (layer6_outputs(1197)));
    outputs(4989) <= layer6_outputs(2841);
    outputs(4990) <= not(layer6_outputs(2619));
    outputs(4991) <= not((layer6_outputs(1546)) xor (layer6_outputs(4577)));
    outputs(4992) <= not(layer6_outputs(1236));
    outputs(4993) <= not((layer6_outputs(2469)) or (layer6_outputs(3810)));
    outputs(4994) <= (layer6_outputs(1480)) xor (layer6_outputs(2991));
    outputs(4995) <= not(layer6_outputs(2860));
    outputs(4996) <= layer6_outputs(2821);
    outputs(4997) <= not((layer6_outputs(2758)) or (layer6_outputs(119)));
    outputs(4998) <= not(layer6_outputs(2317));
    outputs(4999) <= layer6_outputs(883);
    outputs(5000) <= (layer6_outputs(3926)) and not (layer6_outputs(1577));
    outputs(5001) <= not(layer6_outputs(3004));
    outputs(5002) <= layer6_outputs(2248);
    outputs(5003) <= (layer6_outputs(3167)) and not (layer6_outputs(2469));
    outputs(5004) <= layer6_outputs(2813);
    outputs(5005) <= layer6_outputs(32);
    outputs(5006) <= not((layer6_outputs(1776)) xor (layer6_outputs(4275)));
    outputs(5007) <= (layer6_outputs(4182)) xor (layer6_outputs(1101));
    outputs(5008) <= not(layer6_outputs(3896));
    outputs(5009) <= (layer6_outputs(2698)) xor (layer6_outputs(3331));
    outputs(5010) <= not(layer6_outputs(695));
    outputs(5011) <= layer6_outputs(1900);
    outputs(5012) <= layer6_outputs(4305);
    outputs(5013) <= (layer6_outputs(2847)) xor (layer6_outputs(4932));
    outputs(5014) <= layer6_outputs(3453);
    outputs(5015) <= not((layer6_outputs(4046)) or (layer6_outputs(1977)));
    outputs(5016) <= layer6_outputs(1117);
    outputs(5017) <= (layer6_outputs(2932)) xor (layer6_outputs(954));
    outputs(5018) <= not(layer6_outputs(1456));
    outputs(5019) <= not((layer6_outputs(4985)) xor (layer6_outputs(3898)));
    outputs(5020) <= not(layer6_outputs(1519));
    outputs(5021) <= (layer6_outputs(1150)) xor (layer6_outputs(2209));
    outputs(5022) <= layer6_outputs(1723);
    outputs(5023) <= layer6_outputs(3745);
    outputs(5024) <= layer6_outputs(1049);
    outputs(5025) <= (layer6_outputs(1441)) xor (layer6_outputs(551));
    outputs(5026) <= layer6_outputs(3111);
    outputs(5027) <= (layer6_outputs(1783)) xor (layer6_outputs(3416));
    outputs(5028) <= layer6_outputs(1836);
    outputs(5029) <= layer6_outputs(678);
    outputs(5030) <= layer6_outputs(1704);
    outputs(5031) <= not(layer6_outputs(612));
    outputs(5032) <= not(layer6_outputs(1670));
    outputs(5033) <= layer6_outputs(15);
    outputs(5034) <= (layer6_outputs(2736)) xor (layer6_outputs(1831));
    outputs(5035) <= not(layer6_outputs(658));
    outputs(5036) <= not(layer6_outputs(3316));
    outputs(5037) <= not(layer6_outputs(2558));
    outputs(5038) <= not(layer6_outputs(1853));
    outputs(5039) <= layer6_outputs(1389);
    outputs(5040) <= (layer6_outputs(3561)) or (layer6_outputs(4318));
    outputs(5041) <= layer6_outputs(3606);
    outputs(5042) <= not(layer6_outputs(3752));
    outputs(5043) <= not(layer6_outputs(1236));
    outputs(5044) <= not(layer6_outputs(736));
    outputs(5045) <= not((layer6_outputs(4621)) xor (layer6_outputs(1208)));
    outputs(5046) <= not(layer6_outputs(1881));
    outputs(5047) <= layer6_outputs(334);
    outputs(5048) <= not((layer6_outputs(4946)) xor (layer6_outputs(2229)));
    outputs(5049) <= not(layer6_outputs(2006));
    outputs(5050) <= (layer6_outputs(4282)) and not (layer6_outputs(2265));
    outputs(5051) <= not(layer6_outputs(2290));
    outputs(5052) <= layer6_outputs(1608);
    outputs(5053) <= not((layer6_outputs(212)) xor (layer6_outputs(4553)));
    outputs(5054) <= layer6_outputs(2117);
    outputs(5055) <= (layer6_outputs(377)) and not (layer6_outputs(3702));
    outputs(5056) <= layer6_outputs(1731);
    outputs(5057) <= (layer6_outputs(1614)) or (layer6_outputs(2607));
    outputs(5058) <= (layer6_outputs(2773)) and not (layer6_outputs(4523));
    outputs(5059) <= not(layer6_outputs(4476));
    outputs(5060) <= (layer6_outputs(500)) xor (layer6_outputs(1403));
    outputs(5061) <= layer6_outputs(4419);
    outputs(5062) <= layer6_outputs(815);
    outputs(5063) <= not(layer6_outputs(3444));
    outputs(5064) <= not(layer6_outputs(126));
    outputs(5065) <= layer6_outputs(3891);
    outputs(5066) <= layer6_outputs(3732);
    outputs(5067) <= layer6_outputs(1112);
    outputs(5068) <= (layer6_outputs(2382)) xor (layer6_outputs(2164));
    outputs(5069) <= not(layer6_outputs(3786));
    outputs(5070) <= layer6_outputs(1762);
    outputs(5071) <= (layer6_outputs(3224)) and (layer6_outputs(3358));
    outputs(5072) <= (layer6_outputs(4335)) and (layer6_outputs(2666));
    outputs(5073) <= not((layer6_outputs(4269)) xor (layer6_outputs(1350)));
    outputs(5074) <= not(layer6_outputs(355));
    outputs(5075) <= layer6_outputs(4860);
    outputs(5076) <= not((layer6_outputs(589)) and (layer6_outputs(200)));
    outputs(5077) <= not(layer6_outputs(1556));
    outputs(5078) <= (layer6_outputs(3128)) and not (layer6_outputs(4351));
    outputs(5079) <= (layer6_outputs(2384)) xor (layer6_outputs(3588));
    outputs(5080) <= layer6_outputs(3622);
    outputs(5081) <= layer6_outputs(3636);
    outputs(5082) <= not(layer6_outputs(619));
    outputs(5083) <= layer6_outputs(3254);
    outputs(5084) <= layer6_outputs(869);
    outputs(5085) <= (layer6_outputs(3884)) and (layer6_outputs(3870));
    outputs(5086) <= not(layer6_outputs(1423));
    outputs(5087) <= not(layer6_outputs(4438));
    outputs(5088) <= layer6_outputs(3435);
    outputs(5089) <= (layer6_outputs(4664)) and not (layer6_outputs(1982));
    outputs(5090) <= not(layer6_outputs(2601)) or (layer6_outputs(4258));
    outputs(5091) <= not((layer6_outputs(517)) or (layer6_outputs(542)));
    outputs(5092) <= (layer6_outputs(4576)) xor (layer6_outputs(2711));
    outputs(5093) <= not(layer6_outputs(1906));
    outputs(5094) <= not((layer6_outputs(3551)) or (layer6_outputs(1542)));
    outputs(5095) <= not(layer6_outputs(2098));
    outputs(5096) <= layer6_outputs(2663);
    outputs(5097) <= not((layer6_outputs(1557)) xor (layer6_outputs(4281)));
    outputs(5098) <= layer6_outputs(3774);
    outputs(5099) <= layer6_outputs(1171);
    outputs(5100) <= not(layer6_outputs(3281)) or (layer6_outputs(3339));
    outputs(5101) <= layer6_outputs(1877);
    outputs(5102) <= not(layer6_outputs(5107));
    outputs(5103) <= not(layer6_outputs(1616));
    outputs(5104) <= (layer6_outputs(278)) xor (layer6_outputs(4212));
    outputs(5105) <= not(layer6_outputs(4652));
    outputs(5106) <= layer6_outputs(2024);
    outputs(5107) <= not((layer6_outputs(4193)) xor (layer6_outputs(2871)));
    outputs(5108) <= not(layer6_outputs(4499));
    outputs(5109) <= layer6_outputs(4405);
    outputs(5110) <= not(layer6_outputs(4579));
    outputs(5111) <= not(layer6_outputs(2345));
    outputs(5112) <= layer6_outputs(2264);
    outputs(5113) <= not((layer6_outputs(4967)) or (layer6_outputs(658)));
    outputs(5114) <= (layer6_outputs(2769)) and not (layer6_outputs(3330));
    outputs(5115) <= (layer6_outputs(655)) and (layer6_outputs(783));
    outputs(5116) <= layer6_outputs(4303);
    outputs(5117) <= (layer6_outputs(2107)) and not (layer6_outputs(2309));
    outputs(5118) <= (layer6_outputs(2052)) xor (layer6_outputs(1175));
    outputs(5119) <= not(layer6_outputs(812));

end Behavioral;
