library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);
    signal layer1_outputs : std_logic_vector(10239 downto 0);
    signal layer2_outputs : std_logic_vector(10239 downto 0);
    signal layer3_outputs : std_logic_vector(10239 downto 0);
    signal layer4_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= (inputs(167)) and not (inputs(118));
    layer0_outputs(1) <= inputs(188);
    layer0_outputs(2) <= not(inputs(168)) or (inputs(117));
    layer0_outputs(3) <= (inputs(84)) or (inputs(103));
    layer0_outputs(4) <= (inputs(206)) xor (inputs(175));
    layer0_outputs(5) <= not((inputs(119)) xor (inputs(56)));
    layer0_outputs(6) <= not((inputs(122)) and (inputs(172)));
    layer0_outputs(7) <= not(inputs(15)) or (inputs(24));
    layer0_outputs(8) <= inputs(101);
    layer0_outputs(9) <= inputs(171);
    layer0_outputs(10) <= not((inputs(185)) or (inputs(136)));
    layer0_outputs(11) <= (inputs(187)) and not (inputs(22));
    layer0_outputs(12) <= (inputs(205)) xor (inputs(28));
    layer0_outputs(13) <= not((inputs(154)) and (inputs(80)));
    layer0_outputs(14) <= not(inputs(81)) or (inputs(127));
    layer0_outputs(15) <= (inputs(83)) and not (inputs(32));
    layer0_outputs(16) <= (inputs(92)) xor (inputs(38));
    layer0_outputs(17) <= (inputs(208)) and not (inputs(200));
    layer0_outputs(18) <= not((inputs(171)) or (inputs(162)));
    layer0_outputs(19) <= not((inputs(105)) xor (inputs(223)));
    layer0_outputs(20) <= '0';
    layer0_outputs(21) <= (inputs(174)) xor (inputs(201));
    layer0_outputs(22) <= not(inputs(186));
    layer0_outputs(23) <= inputs(129);
    layer0_outputs(24) <= (inputs(95)) xor (inputs(162));
    layer0_outputs(25) <= (inputs(229)) or (inputs(101));
    layer0_outputs(26) <= not(inputs(245)) or (inputs(10));
    layer0_outputs(27) <= not((inputs(37)) xor (inputs(69)));
    layer0_outputs(28) <= not((inputs(216)) or (inputs(177)));
    layer0_outputs(29) <= not((inputs(20)) and (inputs(208)));
    layer0_outputs(30) <= not((inputs(87)) or (inputs(15)));
    layer0_outputs(31) <= (inputs(95)) and not (inputs(250));
    layer0_outputs(32) <= not(inputs(103));
    layer0_outputs(33) <= (inputs(198)) and not (inputs(94));
    layer0_outputs(34) <= inputs(209);
    layer0_outputs(35) <= not(inputs(250)) or (inputs(35));
    layer0_outputs(36) <= (inputs(85)) and (inputs(251));
    layer0_outputs(37) <= not(inputs(203));
    layer0_outputs(38) <= inputs(14);
    layer0_outputs(39) <= (inputs(144)) or (inputs(53));
    layer0_outputs(40) <= not((inputs(73)) or (inputs(163)));
    layer0_outputs(41) <= (inputs(195)) xor (inputs(69));
    layer0_outputs(42) <= (inputs(101)) and not (inputs(51));
    layer0_outputs(43) <= inputs(214);
    layer0_outputs(44) <= (inputs(109)) or (inputs(143));
    layer0_outputs(45) <= '1';
    layer0_outputs(46) <= (inputs(68)) or (inputs(185));
    layer0_outputs(47) <= (inputs(114)) and not (inputs(252));
    layer0_outputs(48) <= not((inputs(90)) or (inputs(74)));
    layer0_outputs(49) <= inputs(152);
    layer0_outputs(50) <= not((inputs(187)) or (inputs(140)));
    layer0_outputs(51) <= (inputs(70)) or (inputs(35));
    layer0_outputs(52) <= inputs(166);
    layer0_outputs(53) <= (inputs(119)) or (inputs(120));
    layer0_outputs(54) <= not(inputs(45)) or (inputs(202));
    layer0_outputs(55) <= (inputs(144)) and not (inputs(146));
    layer0_outputs(56) <= (inputs(249)) and not (inputs(244));
    layer0_outputs(57) <= (inputs(233)) or (inputs(23));
    layer0_outputs(58) <= not(inputs(188));
    layer0_outputs(59) <= not((inputs(9)) or (inputs(121)));
    layer0_outputs(60) <= (inputs(132)) and not (inputs(246));
    layer0_outputs(61) <= inputs(195);
    layer0_outputs(62) <= inputs(66);
    layer0_outputs(63) <= not((inputs(98)) or (inputs(231)));
    layer0_outputs(64) <= not((inputs(59)) or (inputs(116)));
    layer0_outputs(65) <= inputs(124);
    layer0_outputs(66) <= (inputs(43)) and not (inputs(39));
    layer0_outputs(67) <= not(inputs(184)) or (inputs(213));
    layer0_outputs(68) <= inputs(201);
    layer0_outputs(69) <= (inputs(198)) and (inputs(99));
    layer0_outputs(70) <= inputs(61);
    layer0_outputs(71) <= not((inputs(152)) xor (inputs(144)));
    layer0_outputs(72) <= inputs(72);
    layer0_outputs(73) <= not(inputs(131)) or (inputs(76));
    layer0_outputs(74) <= '0';
    layer0_outputs(75) <= (inputs(77)) xor (inputs(217));
    layer0_outputs(76) <= '0';
    layer0_outputs(77) <= not(inputs(112)) or (inputs(184));
    layer0_outputs(78) <= not((inputs(77)) or (inputs(91)));
    layer0_outputs(79) <= '0';
    layer0_outputs(80) <= not((inputs(159)) or (inputs(106)));
    layer0_outputs(81) <= inputs(161);
    layer0_outputs(82) <= inputs(152);
    layer0_outputs(83) <= not((inputs(70)) and (inputs(40)));
    layer0_outputs(84) <= not((inputs(103)) or (inputs(126)));
    layer0_outputs(85) <= not(inputs(37));
    layer0_outputs(86) <= not(inputs(194)) or (inputs(183));
    layer0_outputs(87) <= not((inputs(232)) xor (inputs(252)));
    layer0_outputs(88) <= '0';
    layer0_outputs(89) <= (inputs(85)) and not (inputs(245));
    layer0_outputs(90) <= (inputs(37)) or (inputs(71));
    layer0_outputs(91) <= inputs(86);
    layer0_outputs(92) <= (inputs(28)) and (inputs(172));
    layer0_outputs(93) <= not(inputs(110));
    layer0_outputs(94) <= (inputs(125)) and not (inputs(71));
    layer0_outputs(95) <= inputs(230);
    layer0_outputs(96) <= not(inputs(84));
    layer0_outputs(97) <= (inputs(182)) and not (inputs(211));
    layer0_outputs(98) <= (inputs(220)) or (inputs(54));
    layer0_outputs(99) <= not(inputs(226));
    layer0_outputs(100) <= not(inputs(185)) or (inputs(200));
    layer0_outputs(101) <= not((inputs(238)) or (inputs(26)));
    layer0_outputs(102) <= not((inputs(55)) and (inputs(215)));
    layer0_outputs(103) <= not((inputs(94)) or (inputs(238)));
    layer0_outputs(104) <= (inputs(201)) and not (inputs(62));
    layer0_outputs(105) <= (inputs(156)) xor (inputs(19));
    layer0_outputs(106) <= not(inputs(118)) or (inputs(52));
    layer0_outputs(107) <= not(inputs(4));
    layer0_outputs(108) <= not((inputs(187)) or (inputs(252)));
    layer0_outputs(109) <= '0';
    layer0_outputs(110) <= not((inputs(136)) or (inputs(121)));
    layer0_outputs(111) <= not(inputs(129)) or (inputs(80));
    layer0_outputs(112) <= '0';
    layer0_outputs(113) <= not(inputs(25)) or (inputs(172));
    layer0_outputs(114) <= not(inputs(54));
    layer0_outputs(115) <= (inputs(103)) and not (inputs(188));
    layer0_outputs(116) <= inputs(1);
    layer0_outputs(117) <= not(inputs(122)) or (inputs(20));
    layer0_outputs(118) <= not(inputs(83)) or (inputs(115));
    layer0_outputs(119) <= not((inputs(56)) or (inputs(181)));
    layer0_outputs(120) <= (inputs(136)) or (inputs(26));
    layer0_outputs(121) <= (inputs(235)) and (inputs(236));
    layer0_outputs(122) <= '1';
    layer0_outputs(123) <= not(inputs(110));
    layer0_outputs(124) <= not(inputs(140));
    layer0_outputs(125) <= not(inputs(191));
    layer0_outputs(126) <= '1';
    layer0_outputs(127) <= not((inputs(197)) and (inputs(219)));
    layer0_outputs(128) <= (inputs(87)) and not (inputs(37));
    layer0_outputs(129) <= inputs(214);
    layer0_outputs(130) <= not((inputs(205)) xor (inputs(219)));
    layer0_outputs(131) <= not(inputs(99)) or (inputs(29));
    layer0_outputs(132) <= not(inputs(95));
    layer0_outputs(133) <= '0';
    layer0_outputs(134) <= not((inputs(89)) or (inputs(233)));
    layer0_outputs(135) <= not((inputs(44)) or (inputs(6)));
    layer0_outputs(136) <= (inputs(135)) and not (inputs(98));
    layer0_outputs(137) <= not((inputs(19)) and (inputs(103)));
    layer0_outputs(138) <= not(inputs(224));
    layer0_outputs(139) <= not(inputs(171));
    layer0_outputs(140) <= not(inputs(112)) or (inputs(185));
    layer0_outputs(141) <= (inputs(74)) or (inputs(245));
    layer0_outputs(142) <= (inputs(58)) or (inputs(42));
    layer0_outputs(143) <= (inputs(130)) and not (inputs(179));
    layer0_outputs(144) <= not(inputs(131));
    layer0_outputs(145) <= (inputs(213)) xor (inputs(149));
    layer0_outputs(146) <= (inputs(75)) and (inputs(216));
    layer0_outputs(147) <= not(inputs(240)) or (inputs(249));
    layer0_outputs(148) <= inputs(124);
    layer0_outputs(149) <= (inputs(255)) and not (inputs(25));
    layer0_outputs(150) <= inputs(43);
    layer0_outputs(151) <= '0';
    layer0_outputs(152) <= (inputs(68)) and (inputs(43));
    layer0_outputs(153) <= not((inputs(181)) xor (inputs(24)));
    layer0_outputs(154) <= (inputs(245)) or (inputs(130));
    layer0_outputs(155) <= (inputs(131)) or (inputs(192));
    layer0_outputs(156) <= (inputs(139)) and not (inputs(132));
    layer0_outputs(157) <= inputs(124);
    layer0_outputs(158) <= not(inputs(102));
    layer0_outputs(159) <= '1';
    layer0_outputs(160) <= inputs(245);
    layer0_outputs(161) <= (inputs(75)) and not (inputs(100));
    layer0_outputs(162) <= '0';
    layer0_outputs(163) <= not((inputs(4)) and (inputs(218)));
    layer0_outputs(164) <= (inputs(22)) and not (inputs(155));
    layer0_outputs(165) <= not(inputs(184)) or (inputs(62));
    layer0_outputs(166) <= not((inputs(28)) or (inputs(98)));
    layer0_outputs(167) <= (inputs(167)) or (inputs(148));
    layer0_outputs(168) <= inputs(24);
    layer0_outputs(169) <= (inputs(12)) xor (inputs(49));
    layer0_outputs(170) <= '0';
    layer0_outputs(171) <= inputs(133);
    layer0_outputs(172) <= inputs(115);
    layer0_outputs(173) <= (inputs(112)) and not (inputs(213));
    layer0_outputs(174) <= not((inputs(229)) or (inputs(103)));
    layer0_outputs(175) <= inputs(40);
    layer0_outputs(176) <= (inputs(243)) and not (inputs(41));
    layer0_outputs(177) <= (inputs(184)) xor (inputs(88));
    layer0_outputs(178) <= (inputs(7)) or (inputs(219));
    layer0_outputs(179) <= not(inputs(182)) or (inputs(23));
    layer0_outputs(180) <= not((inputs(137)) or (inputs(90)));
    layer0_outputs(181) <= '1';
    layer0_outputs(182) <= (inputs(95)) and not (inputs(99));
    layer0_outputs(183) <= (inputs(16)) xor (inputs(161));
    layer0_outputs(184) <= (inputs(215)) xor (inputs(89));
    layer0_outputs(185) <= (inputs(124)) xor (inputs(252));
    layer0_outputs(186) <= not(inputs(110)) or (inputs(31));
    layer0_outputs(187) <= (inputs(12)) xor (inputs(100));
    layer0_outputs(188) <= not((inputs(5)) and (inputs(83)));
    layer0_outputs(189) <= inputs(52);
    layer0_outputs(190) <= not((inputs(255)) or (inputs(44)));
    layer0_outputs(191) <= not((inputs(233)) or (inputs(52)));
    layer0_outputs(192) <= not(inputs(135));
    layer0_outputs(193) <= inputs(122);
    layer0_outputs(194) <= not(inputs(103));
    layer0_outputs(195) <= (inputs(180)) and not (inputs(33));
    layer0_outputs(196) <= not((inputs(192)) xor (inputs(190)));
    layer0_outputs(197) <= inputs(21);
    layer0_outputs(198) <= not(inputs(139));
    layer0_outputs(199) <= (inputs(237)) or (inputs(117));
    layer0_outputs(200) <= (inputs(127)) and (inputs(228));
    layer0_outputs(201) <= not(inputs(180)) or (inputs(182));
    layer0_outputs(202) <= (inputs(233)) xor (inputs(229));
    layer0_outputs(203) <= '1';
    layer0_outputs(204) <= not(inputs(214));
    layer0_outputs(205) <= (inputs(227)) and not (inputs(90));
    layer0_outputs(206) <= (inputs(93)) and not (inputs(97));
    layer0_outputs(207) <= not((inputs(177)) or (inputs(136)));
    layer0_outputs(208) <= '0';
    layer0_outputs(209) <= inputs(69);
    layer0_outputs(210) <= not((inputs(29)) or (inputs(105)));
    layer0_outputs(211) <= '0';
    layer0_outputs(212) <= (inputs(122)) and not (inputs(253));
    layer0_outputs(213) <= '1';
    layer0_outputs(214) <= (inputs(228)) and (inputs(236));
    layer0_outputs(215) <= not(inputs(114)) or (inputs(222));
    layer0_outputs(216) <= not(inputs(218)) or (inputs(131));
    layer0_outputs(217) <= (inputs(213)) and (inputs(13));
    layer0_outputs(218) <= '0';
    layer0_outputs(219) <= not(inputs(152));
    layer0_outputs(220) <= not(inputs(153));
    layer0_outputs(221) <= (inputs(182)) and not (inputs(62));
    layer0_outputs(222) <= inputs(88);
    layer0_outputs(223) <= (inputs(115)) and (inputs(232));
    layer0_outputs(224) <= not((inputs(97)) or (inputs(226)));
    layer0_outputs(225) <= not(inputs(200)) or (inputs(117));
    layer0_outputs(226) <= not((inputs(138)) or (inputs(42)));
    layer0_outputs(227) <= (inputs(1)) and (inputs(49));
    layer0_outputs(228) <= '0';
    layer0_outputs(229) <= (inputs(152)) and not (inputs(235));
    layer0_outputs(230) <= not((inputs(118)) or (inputs(217)));
    layer0_outputs(231) <= not((inputs(94)) or (inputs(163)));
    layer0_outputs(232) <= not(inputs(138));
    layer0_outputs(233) <= '1';
    layer0_outputs(234) <= (inputs(105)) and (inputs(98));
    layer0_outputs(235) <= not((inputs(28)) xor (inputs(165)));
    layer0_outputs(236) <= inputs(229);
    layer0_outputs(237) <= (inputs(79)) and not (inputs(63));
    layer0_outputs(238) <= (inputs(137)) and not (inputs(43));
    layer0_outputs(239) <= '1';
    layer0_outputs(240) <= (inputs(208)) and not (inputs(58));
    layer0_outputs(241) <= not(inputs(171)) or (inputs(224));
    layer0_outputs(242) <= not(inputs(133));
    layer0_outputs(243) <= not(inputs(228));
    layer0_outputs(244) <= '1';
    layer0_outputs(245) <= inputs(109);
    layer0_outputs(246) <= inputs(6);
    layer0_outputs(247) <= (inputs(36)) and not (inputs(84));
    layer0_outputs(248) <= not(inputs(98)) or (inputs(240));
    layer0_outputs(249) <= not(inputs(38));
    layer0_outputs(250) <= not(inputs(15));
    layer0_outputs(251) <= not((inputs(237)) and (inputs(48)));
    layer0_outputs(252) <= '1';
    layer0_outputs(253) <= inputs(251);
    layer0_outputs(254) <= (inputs(242)) xor (inputs(182));
    layer0_outputs(255) <= (inputs(40)) xor (inputs(13));
    layer0_outputs(256) <= '0';
    layer0_outputs(257) <= (inputs(153)) xor (inputs(3));
    layer0_outputs(258) <= '1';
    layer0_outputs(259) <= inputs(116);
    layer0_outputs(260) <= inputs(111);
    layer0_outputs(261) <= '1';
    layer0_outputs(262) <= '1';
    layer0_outputs(263) <= (inputs(246)) or (inputs(103));
    layer0_outputs(264) <= inputs(217);
    layer0_outputs(265) <= inputs(188);
    layer0_outputs(266) <= (inputs(19)) and not (inputs(60));
    layer0_outputs(267) <= not((inputs(36)) or (inputs(25)));
    layer0_outputs(268) <= (inputs(123)) and not (inputs(111));
    layer0_outputs(269) <= not(inputs(91)) or (inputs(11));
    layer0_outputs(270) <= not(inputs(251)) or (inputs(181));
    layer0_outputs(271) <= inputs(1);
    layer0_outputs(272) <= (inputs(3)) or (inputs(217));
    layer0_outputs(273) <= not(inputs(139)) or (inputs(253));
    layer0_outputs(274) <= not(inputs(77));
    layer0_outputs(275) <= (inputs(201)) or (inputs(168));
    layer0_outputs(276) <= not(inputs(134)) or (inputs(146));
    layer0_outputs(277) <= (inputs(109)) and not (inputs(206));
    layer0_outputs(278) <= (inputs(248)) and (inputs(133));
    layer0_outputs(279) <= (inputs(7)) or (inputs(164));
    layer0_outputs(280) <= (inputs(150)) and not (inputs(217));
    layer0_outputs(281) <= inputs(161);
    layer0_outputs(282) <= (inputs(214)) or (inputs(20));
    layer0_outputs(283) <= (inputs(5)) xor (inputs(206));
    layer0_outputs(284) <= not((inputs(168)) xor (inputs(222)));
    layer0_outputs(285) <= (inputs(244)) or (inputs(184));
    layer0_outputs(286) <= not(inputs(19));
    layer0_outputs(287) <= inputs(181);
    layer0_outputs(288) <= '1';
    layer0_outputs(289) <= (inputs(156)) or (inputs(10));
    layer0_outputs(290) <= not(inputs(122));
    layer0_outputs(291) <= inputs(161);
    layer0_outputs(292) <= (inputs(104)) xor (inputs(104));
    layer0_outputs(293) <= not(inputs(126));
    layer0_outputs(294) <= (inputs(73)) or (inputs(46));
    layer0_outputs(295) <= (inputs(104)) and not (inputs(134));
    layer0_outputs(296) <= not((inputs(197)) and (inputs(42)));
    layer0_outputs(297) <= not(inputs(82)) or (inputs(50));
    layer0_outputs(298) <= not(inputs(112));
    layer0_outputs(299) <= not(inputs(119));
    layer0_outputs(300) <= '1';
    layer0_outputs(301) <= not((inputs(89)) or (inputs(146)));
    layer0_outputs(302) <= not((inputs(23)) xor (inputs(203)));
    layer0_outputs(303) <= (inputs(119)) and not (inputs(194));
    layer0_outputs(304) <= not(inputs(147));
    layer0_outputs(305) <= not(inputs(245));
    layer0_outputs(306) <= not(inputs(79));
    layer0_outputs(307) <= inputs(125);
    layer0_outputs(308) <= not(inputs(202));
    layer0_outputs(309) <= not(inputs(40));
    layer0_outputs(310) <= inputs(136);
    layer0_outputs(311) <= '1';
    layer0_outputs(312) <= inputs(42);
    layer0_outputs(313) <= not(inputs(212)) or (inputs(6));
    layer0_outputs(314) <= not(inputs(110));
    layer0_outputs(315) <= not((inputs(115)) or (inputs(121)));
    layer0_outputs(316) <= '1';
    layer0_outputs(317) <= inputs(137);
    layer0_outputs(318) <= inputs(14);
    layer0_outputs(319) <= '0';
    layer0_outputs(320) <= not(inputs(189));
    layer0_outputs(321) <= not(inputs(135));
    layer0_outputs(322) <= not(inputs(27)) or (inputs(244));
    layer0_outputs(323) <= not((inputs(205)) or (inputs(128)));
    layer0_outputs(324) <= (inputs(254)) or (inputs(16));
    layer0_outputs(325) <= not(inputs(140));
    layer0_outputs(326) <= not((inputs(50)) xor (inputs(93)));
    layer0_outputs(327) <= inputs(72);
    layer0_outputs(328) <= inputs(209);
    layer0_outputs(329) <= not(inputs(176)) or (inputs(94));
    layer0_outputs(330) <= not(inputs(21)) or (inputs(133));
    layer0_outputs(331) <= (inputs(171)) or (inputs(39));
    layer0_outputs(332) <= inputs(131);
    layer0_outputs(333) <= (inputs(122)) and not (inputs(110));
    layer0_outputs(334) <= inputs(91);
    layer0_outputs(335) <= not((inputs(205)) xor (inputs(196)));
    layer0_outputs(336) <= (inputs(31)) or (inputs(143));
    layer0_outputs(337) <= not((inputs(252)) and (inputs(121)));
    layer0_outputs(338) <= not((inputs(225)) xor (inputs(43)));
    layer0_outputs(339) <= (inputs(1)) xor (inputs(186));
    layer0_outputs(340) <= not((inputs(90)) or (inputs(205)));
    layer0_outputs(341) <= (inputs(90)) or (inputs(173));
    layer0_outputs(342) <= (inputs(97)) or (inputs(120));
    layer0_outputs(343) <= (inputs(205)) and not (inputs(245));
    layer0_outputs(344) <= not(inputs(206));
    layer0_outputs(345) <= not(inputs(216)) or (inputs(32));
    layer0_outputs(346) <= not((inputs(114)) or (inputs(73)));
    layer0_outputs(347) <= not((inputs(193)) xor (inputs(101)));
    layer0_outputs(348) <= (inputs(241)) and (inputs(191));
    layer0_outputs(349) <= not(inputs(226));
    layer0_outputs(350) <= (inputs(204)) and not (inputs(240));
    layer0_outputs(351) <= (inputs(27)) and not (inputs(246));
    layer0_outputs(352) <= not(inputs(97));
    layer0_outputs(353) <= (inputs(52)) and (inputs(251));
    layer0_outputs(354) <= (inputs(233)) xor (inputs(252));
    layer0_outputs(355) <= (inputs(107)) and not (inputs(178));
    layer0_outputs(356) <= not((inputs(113)) xor (inputs(197)));
    layer0_outputs(357) <= not(inputs(11)) or (inputs(67));
    layer0_outputs(358) <= not(inputs(63)) or (inputs(51));
    layer0_outputs(359) <= not((inputs(219)) xor (inputs(216)));
    layer0_outputs(360) <= not(inputs(140)) or (inputs(67));
    layer0_outputs(361) <= not(inputs(160));
    layer0_outputs(362) <= inputs(148);
    layer0_outputs(363) <= not((inputs(55)) or (inputs(118)));
    layer0_outputs(364) <= not((inputs(35)) or (inputs(115)));
    layer0_outputs(365) <= not((inputs(245)) xor (inputs(193)));
    layer0_outputs(366) <= (inputs(137)) or (inputs(173));
    layer0_outputs(367) <= not(inputs(136));
    layer0_outputs(368) <= (inputs(150)) or (inputs(133));
    layer0_outputs(369) <= '1';
    layer0_outputs(370) <= (inputs(87)) and not (inputs(192));
    layer0_outputs(371) <= not((inputs(20)) xor (inputs(136)));
    layer0_outputs(372) <= not((inputs(247)) or (inputs(99)));
    layer0_outputs(373) <= (inputs(78)) or (inputs(118));
    layer0_outputs(374) <= (inputs(244)) or (inputs(32));
    layer0_outputs(375) <= not((inputs(248)) or (inputs(197)));
    layer0_outputs(376) <= not(inputs(253));
    layer0_outputs(377) <= not((inputs(241)) or (inputs(110)));
    layer0_outputs(378) <= not(inputs(82));
    layer0_outputs(379) <= inputs(100);
    layer0_outputs(380) <= not((inputs(207)) xor (inputs(23)));
    layer0_outputs(381) <= '1';
    layer0_outputs(382) <= not(inputs(209)) or (inputs(33));
    layer0_outputs(383) <= (inputs(214)) and not (inputs(127));
    layer0_outputs(384) <= not((inputs(188)) or (inputs(54)));
    layer0_outputs(385) <= (inputs(41)) xor (inputs(16));
    layer0_outputs(386) <= not(inputs(52));
    layer0_outputs(387) <= (inputs(254)) and not (inputs(83));
    layer0_outputs(388) <= not((inputs(93)) or (inputs(65)));
    layer0_outputs(389) <= not(inputs(129));
    layer0_outputs(390) <= not(inputs(120));
    layer0_outputs(391) <= (inputs(94)) xor (inputs(250));
    layer0_outputs(392) <= inputs(161);
    layer0_outputs(393) <= not((inputs(215)) or (inputs(236)));
    layer0_outputs(394) <= '1';
    layer0_outputs(395) <= not(inputs(28));
    layer0_outputs(396) <= not((inputs(159)) xor (inputs(185)));
    layer0_outputs(397) <= (inputs(72)) and not (inputs(31));
    layer0_outputs(398) <= (inputs(150)) and not (inputs(48));
    layer0_outputs(399) <= inputs(217);
    layer0_outputs(400) <= '0';
    layer0_outputs(401) <= not(inputs(230));
    layer0_outputs(402) <= not((inputs(244)) xor (inputs(27)));
    layer0_outputs(403) <= inputs(189);
    layer0_outputs(404) <= not(inputs(73));
    layer0_outputs(405) <= not(inputs(120));
    layer0_outputs(406) <= not(inputs(249)) or (inputs(202));
    layer0_outputs(407) <= not(inputs(223));
    layer0_outputs(408) <= not((inputs(6)) xor (inputs(41)));
    layer0_outputs(409) <= (inputs(209)) xor (inputs(182));
    layer0_outputs(410) <= not(inputs(123));
    layer0_outputs(411) <= inputs(74);
    layer0_outputs(412) <= not(inputs(40));
    layer0_outputs(413) <= not(inputs(120));
    layer0_outputs(414) <= not((inputs(173)) xor (inputs(219)));
    layer0_outputs(415) <= (inputs(148)) or (inputs(33));
    layer0_outputs(416) <= not(inputs(132)) or (inputs(40));
    layer0_outputs(417) <= not(inputs(172)) or (inputs(142));
    layer0_outputs(418) <= inputs(139);
    layer0_outputs(419) <= not((inputs(35)) or (inputs(149)));
    layer0_outputs(420) <= inputs(144);
    layer0_outputs(421) <= not((inputs(135)) or (inputs(138)));
    layer0_outputs(422) <= not((inputs(194)) or (inputs(203)));
    layer0_outputs(423) <= not((inputs(186)) or (inputs(39)));
    layer0_outputs(424) <= not(inputs(91));
    layer0_outputs(425) <= inputs(129);
    layer0_outputs(426) <= not(inputs(5)) or (inputs(11));
    layer0_outputs(427) <= not(inputs(38)) or (inputs(191));
    layer0_outputs(428) <= not((inputs(35)) xor (inputs(222)));
    layer0_outputs(429) <= inputs(255);
    layer0_outputs(430) <= '0';
    layer0_outputs(431) <= not(inputs(220)) or (inputs(77));
    layer0_outputs(432) <= not(inputs(4)) or (inputs(81));
    layer0_outputs(433) <= not((inputs(103)) xor (inputs(224)));
    layer0_outputs(434) <= not(inputs(163));
    layer0_outputs(435) <= (inputs(253)) xor (inputs(69));
    layer0_outputs(436) <= (inputs(133)) and not (inputs(182));
    layer0_outputs(437) <= not((inputs(233)) or (inputs(234)));
    layer0_outputs(438) <= not((inputs(112)) xor (inputs(58)));
    layer0_outputs(439) <= (inputs(13)) or (inputs(12));
    layer0_outputs(440) <= '0';
    layer0_outputs(441) <= not((inputs(209)) or (inputs(154)));
    layer0_outputs(442) <= (inputs(56)) or (inputs(171));
    layer0_outputs(443) <= not((inputs(34)) or (inputs(56)));
    layer0_outputs(444) <= inputs(183);
    layer0_outputs(445) <= not((inputs(188)) xor (inputs(87)));
    layer0_outputs(446) <= not(inputs(214)) or (inputs(183));
    layer0_outputs(447) <= not((inputs(202)) or (inputs(226)));
    layer0_outputs(448) <= (inputs(126)) and not (inputs(12));
    layer0_outputs(449) <= '0';
    layer0_outputs(450) <= (inputs(74)) xor (inputs(59));
    layer0_outputs(451) <= (inputs(175)) xor (inputs(211));
    layer0_outputs(452) <= inputs(60);
    layer0_outputs(453) <= (inputs(203)) and not (inputs(10));
    layer0_outputs(454) <= not(inputs(113));
    layer0_outputs(455) <= not((inputs(46)) or (inputs(114)));
    layer0_outputs(456) <= not((inputs(33)) or (inputs(221)));
    layer0_outputs(457) <= (inputs(243)) xor (inputs(185));
    layer0_outputs(458) <= not((inputs(178)) and (inputs(211)));
    layer0_outputs(459) <= not((inputs(157)) and (inputs(41)));
    layer0_outputs(460) <= '0';
    layer0_outputs(461) <= (inputs(123)) and not (inputs(90));
    layer0_outputs(462) <= (inputs(13)) and not (inputs(9));
    layer0_outputs(463) <= not((inputs(181)) xor (inputs(255)));
    layer0_outputs(464) <= not((inputs(212)) xor (inputs(34)));
    layer0_outputs(465) <= not(inputs(45));
    layer0_outputs(466) <= '0';
    layer0_outputs(467) <= '1';
    layer0_outputs(468) <= inputs(25);
    layer0_outputs(469) <= not(inputs(237));
    layer0_outputs(470) <= (inputs(53)) and not (inputs(8));
    layer0_outputs(471) <= (inputs(220)) and not (inputs(54));
    layer0_outputs(472) <= (inputs(110)) and not (inputs(47));
    layer0_outputs(473) <= not(inputs(151));
    layer0_outputs(474) <= not(inputs(74));
    layer0_outputs(475) <= not(inputs(124));
    layer0_outputs(476) <= not(inputs(87)) or (inputs(191));
    layer0_outputs(477) <= '0';
    layer0_outputs(478) <= inputs(106);
    layer0_outputs(479) <= not(inputs(16));
    layer0_outputs(480) <= not(inputs(120));
    layer0_outputs(481) <= not((inputs(151)) or (inputs(158)));
    layer0_outputs(482) <= (inputs(86)) and not (inputs(191));
    layer0_outputs(483) <= inputs(218);
    layer0_outputs(484) <= (inputs(121)) and not (inputs(1));
    layer0_outputs(485) <= not(inputs(192)) or (inputs(154));
    layer0_outputs(486) <= inputs(215);
    layer0_outputs(487) <= (inputs(21)) xor (inputs(117));
    layer0_outputs(488) <= not(inputs(162)) or (inputs(29));
    layer0_outputs(489) <= not((inputs(7)) or (inputs(173)));
    layer0_outputs(490) <= '1';
    layer0_outputs(491) <= (inputs(120)) and (inputs(67));
    layer0_outputs(492) <= '0';
    layer0_outputs(493) <= (inputs(237)) xor (inputs(117));
    layer0_outputs(494) <= not((inputs(243)) or (inputs(132)));
    layer0_outputs(495) <= not((inputs(240)) or (inputs(74)));
    layer0_outputs(496) <= inputs(199);
    layer0_outputs(497) <= inputs(117);
    layer0_outputs(498) <= not(inputs(71)) or (inputs(253));
    layer0_outputs(499) <= '1';
    layer0_outputs(500) <= inputs(78);
    layer0_outputs(501) <= '1';
    layer0_outputs(502) <= '1';
    layer0_outputs(503) <= not((inputs(61)) or (inputs(49)));
    layer0_outputs(504) <= '1';
    layer0_outputs(505) <= '1';
    layer0_outputs(506) <= not(inputs(51)) or (inputs(99));
    layer0_outputs(507) <= not(inputs(51));
    layer0_outputs(508) <= not((inputs(212)) and (inputs(170)));
    layer0_outputs(509) <= inputs(61);
    layer0_outputs(510) <= not((inputs(68)) or (inputs(92)));
    layer0_outputs(511) <= not(inputs(75));
    layer0_outputs(512) <= not(inputs(120));
    layer0_outputs(513) <= not(inputs(183)) or (inputs(89));
    layer0_outputs(514) <= not(inputs(23)) or (inputs(61));
    layer0_outputs(515) <= (inputs(178)) and not (inputs(46));
    layer0_outputs(516) <= inputs(218);
    layer0_outputs(517) <= (inputs(222)) or (inputs(224));
    layer0_outputs(518) <= (inputs(13)) or (inputs(5));
    layer0_outputs(519) <= inputs(28);
    layer0_outputs(520) <= not(inputs(163));
    layer0_outputs(521) <= not(inputs(93)) or (inputs(71));
    layer0_outputs(522) <= (inputs(207)) and not (inputs(139));
    layer0_outputs(523) <= (inputs(229)) or (inputs(102));
    layer0_outputs(524) <= inputs(197);
    layer0_outputs(525) <= not((inputs(75)) and (inputs(73)));
    layer0_outputs(526) <= (inputs(213)) and not (inputs(68));
    layer0_outputs(527) <= '0';
    layer0_outputs(528) <= not((inputs(168)) or (inputs(106)));
    layer0_outputs(529) <= (inputs(69)) and not (inputs(170));
    layer0_outputs(530) <= not(inputs(145));
    layer0_outputs(531) <= not(inputs(84));
    layer0_outputs(532) <= not((inputs(140)) xor (inputs(200)));
    layer0_outputs(533) <= (inputs(26)) xor (inputs(118));
    layer0_outputs(534) <= inputs(118);
    layer0_outputs(535) <= '1';
    layer0_outputs(536) <= not((inputs(205)) xor (inputs(59)));
    layer0_outputs(537) <= not(inputs(29));
    layer0_outputs(538) <= not((inputs(83)) or (inputs(116)));
    layer0_outputs(539) <= (inputs(183)) and not (inputs(47));
    layer0_outputs(540) <= not((inputs(23)) and (inputs(13)));
    layer0_outputs(541) <= not(inputs(136));
    layer0_outputs(542) <= inputs(132);
    layer0_outputs(543) <= not(inputs(69)) or (inputs(197));
    layer0_outputs(544) <= not((inputs(36)) and (inputs(70)));
    layer0_outputs(545) <= not(inputs(163)) or (inputs(38));
    layer0_outputs(546) <= not(inputs(15));
    layer0_outputs(547) <= not((inputs(65)) xor (inputs(7)));
    layer0_outputs(548) <= (inputs(123)) xor (inputs(75));
    layer0_outputs(549) <= not(inputs(50));
    layer0_outputs(550) <= inputs(151);
    layer0_outputs(551) <= not((inputs(23)) or (inputs(112)));
    layer0_outputs(552) <= (inputs(201)) xor (inputs(143));
    layer0_outputs(553) <= '1';
    layer0_outputs(554) <= (inputs(221)) or (inputs(120));
    layer0_outputs(555) <= not(inputs(243)) or (inputs(14));
    layer0_outputs(556) <= not(inputs(122)) or (inputs(22));
    layer0_outputs(557) <= not(inputs(39)) or (inputs(98));
    layer0_outputs(558) <= not((inputs(65)) and (inputs(188)));
    layer0_outputs(559) <= not(inputs(144)) or (inputs(186));
    layer0_outputs(560) <= (inputs(39)) or (inputs(174));
    layer0_outputs(561) <= (inputs(107)) and not (inputs(226));
    layer0_outputs(562) <= (inputs(30)) xor (inputs(57));
    layer0_outputs(563) <= (inputs(14)) and not (inputs(118));
    layer0_outputs(564) <= not((inputs(138)) or (inputs(233)));
    layer0_outputs(565) <= not((inputs(79)) xor (inputs(15)));
    layer0_outputs(566) <= (inputs(147)) or (inputs(9));
    layer0_outputs(567) <= not((inputs(213)) or (inputs(239)));
    layer0_outputs(568) <= (inputs(150)) xor (inputs(177));
    layer0_outputs(569) <= (inputs(242)) and not (inputs(184));
    layer0_outputs(570) <= (inputs(221)) and not (inputs(174));
    layer0_outputs(571) <= not(inputs(160)) or (inputs(78));
    layer0_outputs(572) <= not(inputs(57)) or (inputs(35));
    layer0_outputs(573) <= not((inputs(62)) or (inputs(24)));
    layer0_outputs(574) <= (inputs(82)) or (inputs(74));
    layer0_outputs(575) <= not(inputs(243));
    layer0_outputs(576) <= inputs(30);
    layer0_outputs(577) <= (inputs(236)) and not (inputs(82));
    layer0_outputs(578) <= '0';
    layer0_outputs(579) <= not((inputs(226)) and (inputs(219)));
    layer0_outputs(580) <= (inputs(114)) and not (inputs(233));
    layer0_outputs(581) <= (inputs(105)) and not (inputs(31));
    layer0_outputs(582) <= inputs(246);
    layer0_outputs(583) <= not((inputs(104)) xor (inputs(63)));
    layer0_outputs(584) <= not(inputs(202));
    layer0_outputs(585) <= (inputs(212)) or (inputs(194));
    layer0_outputs(586) <= (inputs(151)) and not (inputs(18));
    layer0_outputs(587) <= not((inputs(75)) or (inputs(85)));
    layer0_outputs(588) <= (inputs(42)) and not (inputs(211));
    layer0_outputs(589) <= not(inputs(133));
    layer0_outputs(590) <= inputs(118);
    layer0_outputs(591) <= '0';
    layer0_outputs(592) <= (inputs(26)) xor (inputs(219));
    layer0_outputs(593) <= (inputs(175)) or (inputs(79));
    layer0_outputs(594) <= (inputs(94)) xor (inputs(47));
    layer0_outputs(595) <= not((inputs(231)) or (inputs(97)));
    layer0_outputs(596) <= (inputs(93)) and not (inputs(122));
    layer0_outputs(597) <= (inputs(25)) and not (inputs(222));
    layer0_outputs(598) <= not((inputs(47)) and (inputs(111)));
    layer0_outputs(599) <= not(inputs(187));
    layer0_outputs(600) <= inputs(185);
    layer0_outputs(601) <= (inputs(233)) or (inputs(177));
    layer0_outputs(602) <= not(inputs(143));
    layer0_outputs(603) <= not((inputs(194)) and (inputs(205)));
    layer0_outputs(604) <= inputs(192);
    layer0_outputs(605) <= (inputs(50)) or (inputs(24));
    layer0_outputs(606) <= '1';
    layer0_outputs(607) <= not(inputs(164)) or (inputs(106));
    layer0_outputs(608) <= not((inputs(44)) xor (inputs(137)));
    layer0_outputs(609) <= not((inputs(226)) or (inputs(119)));
    layer0_outputs(610) <= '1';
    layer0_outputs(611) <= (inputs(151)) xor (inputs(45));
    layer0_outputs(612) <= (inputs(209)) and not (inputs(176));
    layer0_outputs(613) <= not((inputs(224)) xor (inputs(34)));
    layer0_outputs(614) <= (inputs(254)) or (inputs(167));
    layer0_outputs(615) <= not(inputs(148));
    layer0_outputs(616) <= (inputs(51)) and (inputs(130));
    layer0_outputs(617) <= (inputs(168)) or (inputs(88));
    layer0_outputs(618) <= (inputs(125)) or (inputs(124));
    layer0_outputs(619) <= not(inputs(23));
    layer0_outputs(620) <= (inputs(197)) or (inputs(75));
    layer0_outputs(621) <= (inputs(69)) or (inputs(175));
    layer0_outputs(622) <= (inputs(42)) and not (inputs(129));
    layer0_outputs(623) <= (inputs(145)) or (inputs(174));
    layer0_outputs(624) <= not(inputs(169)) or (inputs(78));
    layer0_outputs(625) <= (inputs(195)) and not (inputs(25));
    layer0_outputs(626) <= inputs(171);
    layer0_outputs(627) <= inputs(96);
    layer0_outputs(628) <= not((inputs(239)) xor (inputs(26)));
    layer0_outputs(629) <= (inputs(197)) and not (inputs(10));
    layer0_outputs(630) <= (inputs(195)) or (inputs(42));
    layer0_outputs(631) <= inputs(144);
    layer0_outputs(632) <= (inputs(29)) xor (inputs(68));
    layer0_outputs(633) <= not((inputs(25)) or (inputs(247)));
    layer0_outputs(634) <= inputs(101);
    layer0_outputs(635) <= not(inputs(7)) or (inputs(44));
    layer0_outputs(636) <= inputs(34);
    layer0_outputs(637) <= not(inputs(229)) or (inputs(175));
    layer0_outputs(638) <= not(inputs(228));
    layer0_outputs(639) <= not(inputs(45)) or (inputs(186));
    layer0_outputs(640) <= not(inputs(230)) or (inputs(183));
    layer0_outputs(641) <= inputs(124);
    layer0_outputs(642) <= not(inputs(41)) or (inputs(203));
    layer0_outputs(643) <= '0';
    layer0_outputs(644) <= inputs(133);
    layer0_outputs(645) <= (inputs(152)) and not (inputs(128));
    layer0_outputs(646) <= '0';
    layer0_outputs(647) <= not(inputs(26));
    layer0_outputs(648) <= not(inputs(216));
    layer0_outputs(649) <= not(inputs(95)) or (inputs(84));
    layer0_outputs(650) <= not((inputs(22)) or (inputs(150)));
    layer0_outputs(651) <= (inputs(145)) or (inputs(213));
    layer0_outputs(652) <= (inputs(68)) and not (inputs(208));
    layer0_outputs(653) <= (inputs(103)) or (inputs(234));
    layer0_outputs(654) <= inputs(86);
    layer0_outputs(655) <= not((inputs(124)) or (inputs(241)));
    layer0_outputs(656) <= not((inputs(125)) or (inputs(197)));
    layer0_outputs(657) <= inputs(89);
    layer0_outputs(658) <= '0';
    layer0_outputs(659) <= '0';
    layer0_outputs(660) <= not(inputs(136));
    layer0_outputs(661) <= inputs(198);
    layer0_outputs(662) <= (inputs(143)) and not (inputs(70));
    layer0_outputs(663) <= inputs(194);
    layer0_outputs(664) <= not((inputs(2)) xor (inputs(188)));
    layer0_outputs(665) <= not(inputs(30)) or (inputs(48));
    layer0_outputs(666) <= (inputs(49)) and (inputs(126));
    layer0_outputs(667) <= not(inputs(84));
    layer0_outputs(668) <= '0';
    layer0_outputs(669) <= (inputs(104)) and (inputs(24));
    layer0_outputs(670) <= (inputs(130)) xor (inputs(252));
    layer0_outputs(671) <= (inputs(177)) and not (inputs(45));
    layer0_outputs(672) <= inputs(115);
    layer0_outputs(673) <= not(inputs(59));
    layer0_outputs(674) <= (inputs(206)) or (inputs(61));
    layer0_outputs(675) <= not(inputs(148)) or (inputs(66));
    layer0_outputs(676) <= inputs(233);
    layer0_outputs(677) <= not(inputs(158)) or (inputs(255));
    layer0_outputs(678) <= inputs(127);
    layer0_outputs(679) <= not(inputs(231));
    layer0_outputs(680) <= (inputs(189)) and (inputs(2));
    layer0_outputs(681) <= inputs(248);
    layer0_outputs(682) <= not((inputs(207)) or (inputs(95)));
    layer0_outputs(683) <= not((inputs(78)) or (inputs(37)));
    layer0_outputs(684) <= inputs(123);
    layer0_outputs(685) <= inputs(176);
    layer0_outputs(686) <= '0';
    layer0_outputs(687) <= not((inputs(194)) or (inputs(56)));
    layer0_outputs(688) <= (inputs(6)) and not (inputs(72));
    layer0_outputs(689) <= not(inputs(143));
    layer0_outputs(690) <= (inputs(54)) or (inputs(170));
    layer0_outputs(691) <= not((inputs(110)) xor (inputs(66)));
    layer0_outputs(692) <= not((inputs(160)) xor (inputs(235)));
    layer0_outputs(693) <= not(inputs(16));
    layer0_outputs(694) <= (inputs(179)) and (inputs(29));
    layer0_outputs(695) <= (inputs(122)) and not (inputs(62));
    layer0_outputs(696) <= (inputs(164)) and not (inputs(143));
    layer0_outputs(697) <= not(inputs(245));
    layer0_outputs(698) <= not(inputs(162));
    layer0_outputs(699) <= not((inputs(20)) or (inputs(89)));
    layer0_outputs(700) <= not((inputs(219)) xor (inputs(102)));
    layer0_outputs(701) <= not(inputs(38)) or (inputs(8));
    layer0_outputs(702) <= (inputs(203)) xor (inputs(172));
    layer0_outputs(703) <= not((inputs(72)) xor (inputs(23)));
    layer0_outputs(704) <= (inputs(134)) or (inputs(119));
    layer0_outputs(705) <= not((inputs(42)) or (inputs(108)));
    layer0_outputs(706) <= inputs(93);
    layer0_outputs(707) <= '1';
    layer0_outputs(708) <= inputs(166);
    layer0_outputs(709) <= not(inputs(244));
    layer0_outputs(710) <= (inputs(117)) or (inputs(140));
    layer0_outputs(711) <= '0';
    layer0_outputs(712) <= not((inputs(16)) xor (inputs(67)));
    layer0_outputs(713) <= not((inputs(208)) and (inputs(34)));
    layer0_outputs(714) <= (inputs(38)) and not (inputs(70));
    layer0_outputs(715) <= not(inputs(126));
    layer0_outputs(716) <= not((inputs(255)) or (inputs(14)));
    layer0_outputs(717) <= (inputs(145)) or (inputs(139));
    layer0_outputs(718) <= (inputs(159)) and not (inputs(219));
    layer0_outputs(719) <= not(inputs(45)) or (inputs(187));
    layer0_outputs(720) <= (inputs(99)) and not (inputs(42));
    layer0_outputs(721) <= not(inputs(228)) or (inputs(253));
    layer0_outputs(722) <= not((inputs(232)) or (inputs(75)));
    layer0_outputs(723) <= not((inputs(145)) or (inputs(195)));
    layer0_outputs(724) <= not(inputs(93)) or (inputs(22));
    layer0_outputs(725) <= (inputs(142)) and (inputs(30));
    layer0_outputs(726) <= inputs(196);
    layer0_outputs(727) <= (inputs(122)) and not (inputs(104));
    layer0_outputs(728) <= (inputs(17)) and not (inputs(102));
    layer0_outputs(729) <= '1';
    layer0_outputs(730) <= not(inputs(205)) or (inputs(250));
    layer0_outputs(731) <= '1';
    layer0_outputs(732) <= not(inputs(247)) or (inputs(142));
    layer0_outputs(733) <= not((inputs(159)) xor (inputs(156)));
    layer0_outputs(734) <= (inputs(23)) xor (inputs(171));
    layer0_outputs(735) <= not(inputs(115)) or (inputs(51));
    layer0_outputs(736) <= (inputs(34)) and not (inputs(114));
    layer0_outputs(737) <= (inputs(247)) xor (inputs(8));
    layer0_outputs(738) <= inputs(35);
    layer0_outputs(739) <= inputs(90);
    layer0_outputs(740) <= not(inputs(150));
    layer0_outputs(741) <= not(inputs(18)) or (inputs(229));
    layer0_outputs(742) <= not((inputs(178)) or (inputs(57)));
    layer0_outputs(743) <= '0';
    layer0_outputs(744) <= not(inputs(10)) or (inputs(245));
    layer0_outputs(745) <= (inputs(173)) or (inputs(165));
    layer0_outputs(746) <= not((inputs(144)) and (inputs(176)));
    layer0_outputs(747) <= not((inputs(92)) or (inputs(124)));
    layer0_outputs(748) <= (inputs(255)) and not (inputs(94));
    layer0_outputs(749) <= not(inputs(163)) or (inputs(234));
    layer0_outputs(750) <= not(inputs(119)) or (inputs(235));
    layer0_outputs(751) <= not(inputs(76));
    layer0_outputs(752) <= not((inputs(246)) or (inputs(141)));
    layer0_outputs(753) <= not(inputs(40));
    layer0_outputs(754) <= inputs(119);
    layer0_outputs(755) <= (inputs(28)) and not (inputs(113));
    layer0_outputs(756) <= not(inputs(177));
    layer0_outputs(757) <= (inputs(43)) and (inputs(227));
    layer0_outputs(758) <= (inputs(128)) or (inputs(104));
    layer0_outputs(759) <= not(inputs(36));
    layer0_outputs(760) <= (inputs(244)) xor (inputs(126));
    layer0_outputs(761) <= not((inputs(195)) or (inputs(172)));
    layer0_outputs(762) <= not(inputs(61)) or (inputs(14));
    layer0_outputs(763) <= (inputs(155)) and not (inputs(41));
    layer0_outputs(764) <= not(inputs(103));
    layer0_outputs(765) <= (inputs(178)) xor (inputs(51));
    layer0_outputs(766) <= (inputs(225)) and not (inputs(104));
    layer0_outputs(767) <= not((inputs(251)) xor (inputs(186)));
    layer0_outputs(768) <= (inputs(105)) and not (inputs(134));
    layer0_outputs(769) <= '1';
    layer0_outputs(770) <= (inputs(38)) and not (inputs(160));
    layer0_outputs(771) <= not((inputs(18)) or (inputs(110)));
    layer0_outputs(772) <= not(inputs(236));
    layer0_outputs(773) <= not(inputs(15)) or (inputs(247));
    layer0_outputs(774) <= inputs(59);
    layer0_outputs(775) <= (inputs(119)) or (inputs(178));
    layer0_outputs(776) <= '1';
    layer0_outputs(777) <= not((inputs(51)) xor (inputs(226)));
    layer0_outputs(778) <= not((inputs(143)) and (inputs(105)));
    layer0_outputs(779) <= (inputs(127)) or (inputs(68));
    layer0_outputs(780) <= (inputs(16)) and not (inputs(3));
    layer0_outputs(781) <= (inputs(230)) or (inputs(136));
    layer0_outputs(782) <= (inputs(125)) xor (inputs(182));
    layer0_outputs(783) <= not(inputs(211));
    layer0_outputs(784) <= not((inputs(75)) or (inputs(203)));
    layer0_outputs(785) <= not(inputs(253)) or (inputs(18));
    layer0_outputs(786) <= inputs(31);
    layer0_outputs(787) <= not((inputs(252)) and (inputs(45)));
    layer0_outputs(788) <= (inputs(110)) and not (inputs(67));
    layer0_outputs(789) <= not((inputs(68)) and (inputs(52)));
    layer0_outputs(790) <= not((inputs(186)) and (inputs(151)));
    layer0_outputs(791) <= (inputs(227)) xor (inputs(137));
    layer0_outputs(792) <= not((inputs(129)) or (inputs(125)));
    layer0_outputs(793) <= (inputs(224)) or (inputs(148));
    layer0_outputs(794) <= (inputs(111)) and (inputs(94));
    layer0_outputs(795) <= not(inputs(149)) or (inputs(175));
    layer0_outputs(796) <= not((inputs(75)) xor (inputs(43)));
    layer0_outputs(797) <= (inputs(172)) or (inputs(190));
    layer0_outputs(798) <= (inputs(84)) and not (inputs(112));
    layer0_outputs(799) <= (inputs(13)) and (inputs(154));
    layer0_outputs(800) <= (inputs(20)) or (inputs(220));
    layer0_outputs(801) <= not((inputs(93)) or (inputs(107)));
    layer0_outputs(802) <= inputs(26);
    layer0_outputs(803) <= (inputs(200)) and not (inputs(69));
    layer0_outputs(804) <= (inputs(224)) xor (inputs(132));
    layer0_outputs(805) <= inputs(135);
    layer0_outputs(806) <= not(inputs(168));
    layer0_outputs(807) <= (inputs(56)) and not (inputs(47));
    layer0_outputs(808) <= (inputs(66)) or (inputs(186));
    layer0_outputs(809) <= not((inputs(248)) xor (inputs(69)));
    layer0_outputs(810) <= (inputs(167)) or (inputs(136));
    layer0_outputs(811) <= (inputs(176)) xor (inputs(152));
    layer0_outputs(812) <= not(inputs(221)) or (inputs(146));
    layer0_outputs(813) <= (inputs(78)) and not (inputs(184));
    layer0_outputs(814) <= (inputs(80)) or (inputs(220));
    layer0_outputs(815) <= inputs(218);
    layer0_outputs(816) <= (inputs(164)) xor (inputs(150));
    layer0_outputs(817) <= not((inputs(198)) and (inputs(198)));
    layer0_outputs(818) <= (inputs(42)) and not (inputs(111));
    layer0_outputs(819) <= inputs(24);
    layer0_outputs(820) <= not(inputs(243)) or (inputs(178));
    layer0_outputs(821) <= (inputs(152)) and not (inputs(33));
    layer0_outputs(822) <= not((inputs(94)) and (inputs(203)));
    layer0_outputs(823) <= not((inputs(28)) or (inputs(124)));
    layer0_outputs(824) <= inputs(141);
    layer0_outputs(825) <= not(inputs(125));
    layer0_outputs(826) <= (inputs(113)) or (inputs(101));
    layer0_outputs(827) <= inputs(47);
    layer0_outputs(828) <= '0';
    layer0_outputs(829) <= (inputs(80)) and (inputs(207));
    layer0_outputs(830) <= (inputs(254)) or (inputs(9));
    layer0_outputs(831) <= inputs(243);
    layer0_outputs(832) <= not(inputs(37)) or (inputs(11));
    layer0_outputs(833) <= '1';
    layer0_outputs(834) <= (inputs(248)) and not (inputs(72));
    layer0_outputs(835) <= not(inputs(170));
    layer0_outputs(836) <= (inputs(142)) and not (inputs(177));
    layer0_outputs(837) <= (inputs(89)) or (inputs(34));
    layer0_outputs(838) <= not((inputs(250)) xor (inputs(18)));
    layer0_outputs(839) <= not(inputs(50));
    layer0_outputs(840) <= (inputs(202)) or (inputs(71));
    layer0_outputs(841) <= (inputs(205)) and (inputs(225));
    layer0_outputs(842) <= (inputs(28)) and not (inputs(176));
    layer0_outputs(843) <= (inputs(19)) and not (inputs(212));
    layer0_outputs(844) <= inputs(0);
    layer0_outputs(845) <= (inputs(186)) and not (inputs(14));
    layer0_outputs(846) <= not((inputs(10)) or (inputs(180)));
    layer0_outputs(847) <= not(inputs(20));
    layer0_outputs(848) <= not((inputs(140)) xor (inputs(245)));
    layer0_outputs(849) <= not(inputs(132)) or (inputs(193));
    layer0_outputs(850) <= not(inputs(61));
    layer0_outputs(851) <= (inputs(158)) or (inputs(72));
    layer0_outputs(852) <= (inputs(139)) xor (inputs(30));
    layer0_outputs(853) <= not((inputs(163)) xor (inputs(157)));
    layer0_outputs(854) <= inputs(229);
    layer0_outputs(855) <= (inputs(149)) and not (inputs(27));
    layer0_outputs(856) <= inputs(137);
    layer0_outputs(857) <= inputs(49);
    layer0_outputs(858) <= (inputs(158)) xor (inputs(6));
    layer0_outputs(859) <= (inputs(81)) and not (inputs(72));
    layer0_outputs(860) <= (inputs(128)) and not (inputs(172));
    layer0_outputs(861) <= inputs(118);
    layer0_outputs(862) <= (inputs(145)) and not (inputs(249));
    layer0_outputs(863) <= (inputs(28)) and not (inputs(143));
    layer0_outputs(864) <= not(inputs(22));
    layer0_outputs(865) <= not(inputs(69)) or (inputs(0));
    layer0_outputs(866) <= inputs(206);
    layer0_outputs(867) <= inputs(54);
    layer0_outputs(868) <= not(inputs(58)) or (inputs(229));
    layer0_outputs(869) <= not(inputs(94)) or (inputs(205));
    layer0_outputs(870) <= not(inputs(138)) or (inputs(192));
    layer0_outputs(871) <= not(inputs(99)) or (inputs(252));
    layer0_outputs(872) <= not(inputs(72)) or (inputs(207));
    layer0_outputs(873) <= (inputs(238)) or (inputs(220));
    layer0_outputs(874) <= '0';
    layer0_outputs(875) <= not((inputs(223)) xor (inputs(58)));
    layer0_outputs(876) <= not(inputs(121)) or (inputs(240));
    layer0_outputs(877) <= (inputs(165)) or (inputs(120));
    layer0_outputs(878) <= not(inputs(116)) or (inputs(58));
    layer0_outputs(879) <= not((inputs(108)) or (inputs(121)));
    layer0_outputs(880) <= inputs(207);
    layer0_outputs(881) <= '0';
    layer0_outputs(882) <= (inputs(227)) or (inputs(255));
    layer0_outputs(883) <= (inputs(206)) and (inputs(35));
    layer0_outputs(884) <= (inputs(195)) xor (inputs(62));
    layer0_outputs(885) <= (inputs(80)) and not (inputs(158));
    layer0_outputs(886) <= '0';
    layer0_outputs(887) <= not((inputs(5)) xor (inputs(156)));
    layer0_outputs(888) <= inputs(117);
    layer0_outputs(889) <= (inputs(121)) and not (inputs(196));
    layer0_outputs(890) <= (inputs(210)) xor (inputs(136));
    layer0_outputs(891) <= not(inputs(65));
    layer0_outputs(892) <= not(inputs(44));
    layer0_outputs(893) <= (inputs(56)) and (inputs(91));
    layer0_outputs(894) <= inputs(73);
    layer0_outputs(895) <= (inputs(119)) or (inputs(134));
    layer0_outputs(896) <= '0';
    layer0_outputs(897) <= not((inputs(82)) or (inputs(153)));
    layer0_outputs(898) <= not((inputs(70)) and (inputs(7)));
    layer0_outputs(899) <= inputs(170);
    layer0_outputs(900) <= not(inputs(140));
    layer0_outputs(901) <= inputs(227);
    layer0_outputs(902) <= (inputs(21)) or (inputs(20));
    layer0_outputs(903) <= (inputs(250)) xor (inputs(148));
    layer0_outputs(904) <= not((inputs(209)) and (inputs(10)));
    layer0_outputs(905) <= (inputs(81)) and not (inputs(129));
    layer0_outputs(906) <= not((inputs(118)) or (inputs(149)));
    layer0_outputs(907) <= not((inputs(81)) or (inputs(22)));
    layer0_outputs(908) <= '0';
    layer0_outputs(909) <= (inputs(250)) xor (inputs(87));
    layer0_outputs(910) <= (inputs(33)) and (inputs(169));
    layer0_outputs(911) <= inputs(71);
    layer0_outputs(912) <= inputs(214);
    layer0_outputs(913) <= inputs(22);
    layer0_outputs(914) <= not(inputs(218));
    layer0_outputs(915) <= not(inputs(242)) or (inputs(205));
    layer0_outputs(916) <= not((inputs(161)) or (inputs(227)));
    layer0_outputs(917) <= not((inputs(7)) or (inputs(24)));
    layer0_outputs(918) <= inputs(208);
    layer0_outputs(919) <= (inputs(94)) xor (inputs(5));
    layer0_outputs(920) <= (inputs(193)) xor (inputs(123));
    layer0_outputs(921) <= not(inputs(122));
    layer0_outputs(922) <= not(inputs(225));
    layer0_outputs(923) <= '0';
    layer0_outputs(924) <= '1';
    layer0_outputs(925) <= (inputs(231)) and not (inputs(200));
    layer0_outputs(926) <= '0';
    layer0_outputs(927) <= '1';
    layer0_outputs(928) <= not(inputs(138)) or (inputs(151));
    layer0_outputs(929) <= '0';
    layer0_outputs(930) <= '1';
    layer0_outputs(931) <= '1';
    layer0_outputs(932) <= (inputs(229)) and not (inputs(187));
    layer0_outputs(933) <= '1';
    layer0_outputs(934) <= not((inputs(81)) or (inputs(184)));
    layer0_outputs(935) <= (inputs(185)) and not (inputs(214));
    layer0_outputs(936) <= not((inputs(92)) or (inputs(182)));
    layer0_outputs(937) <= (inputs(215)) and not (inputs(194));
    layer0_outputs(938) <= inputs(74);
    layer0_outputs(939) <= (inputs(87)) and not (inputs(179));
    layer0_outputs(940) <= (inputs(94)) and not (inputs(80));
    layer0_outputs(941) <= not(inputs(185));
    layer0_outputs(942) <= inputs(218);
    layer0_outputs(943) <= not(inputs(230)) or (inputs(26));
    layer0_outputs(944) <= inputs(119);
    layer0_outputs(945) <= not(inputs(174)) or (inputs(79));
    layer0_outputs(946) <= not(inputs(135));
    layer0_outputs(947) <= '1';
    layer0_outputs(948) <= not((inputs(96)) xor (inputs(153)));
    layer0_outputs(949) <= not(inputs(202)) or (inputs(1));
    layer0_outputs(950) <= (inputs(207)) and not (inputs(19));
    layer0_outputs(951) <= '1';
    layer0_outputs(952) <= not((inputs(63)) and (inputs(193)));
    layer0_outputs(953) <= (inputs(239)) xor (inputs(80));
    layer0_outputs(954) <= (inputs(42)) and (inputs(191));
    layer0_outputs(955) <= not((inputs(76)) xor (inputs(103)));
    layer0_outputs(956) <= not((inputs(71)) xor (inputs(236)));
    layer0_outputs(957) <= (inputs(66)) and not (inputs(31));
    layer0_outputs(958) <= (inputs(170)) or (inputs(239));
    layer0_outputs(959) <= (inputs(112)) and (inputs(253));
    layer0_outputs(960) <= not((inputs(91)) and (inputs(79)));
    layer0_outputs(961) <= not(inputs(163));
    layer0_outputs(962) <= not(inputs(24)) or (inputs(78));
    layer0_outputs(963) <= (inputs(140)) and not (inputs(253));
    layer0_outputs(964) <= (inputs(204)) and not (inputs(22));
    layer0_outputs(965) <= '0';
    layer0_outputs(966) <= not((inputs(231)) or (inputs(163)));
    layer0_outputs(967) <= (inputs(170)) and not (inputs(195));
    layer0_outputs(968) <= '0';
    layer0_outputs(969) <= '0';
    layer0_outputs(970) <= not(inputs(70)) or (inputs(62));
    layer0_outputs(971) <= not(inputs(114));
    layer0_outputs(972) <= not(inputs(81));
    layer0_outputs(973) <= (inputs(87)) and not (inputs(213));
    layer0_outputs(974) <= '0';
    layer0_outputs(975) <= inputs(182);
    layer0_outputs(976) <= (inputs(31)) xor (inputs(14));
    layer0_outputs(977) <= not(inputs(156)) or (inputs(52));
    layer0_outputs(978) <= not(inputs(204));
    layer0_outputs(979) <= (inputs(105)) xor (inputs(211));
    layer0_outputs(980) <= (inputs(164)) or (inputs(125));
    layer0_outputs(981) <= not(inputs(193)) or (inputs(12));
    layer0_outputs(982) <= not(inputs(5));
    layer0_outputs(983) <= inputs(194);
    layer0_outputs(984) <= inputs(106);
    layer0_outputs(985) <= not(inputs(72));
    layer0_outputs(986) <= '1';
    layer0_outputs(987) <= inputs(113);
    layer0_outputs(988) <= '0';
    layer0_outputs(989) <= not(inputs(223)) or (inputs(36));
    layer0_outputs(990) <= not(inputs(185)) or (inputs(233));
    layer0_outputs(991) <= '1';
    layer0_outputs(992) <= (inputs(53)) and not (inputs(78));
    layer0_outputs(993) <= not(inputs(167)) or (inputs(84));
    layer0_outputs(994) <= not((inputs(111)) xor (inputs(85)));
    layer0_outputs(995) <= not(inputs(61));
    layer0_outputs(996) <= '0';
    layer0_outputs(997) <= not(inputs(14));
    layer0_outputs(998) <= not(inputs(21)) or (inputs(130));
    layer0_outputs(999) <= (inputs(106)) and not (inputs(196));
    layer0_outputs(1000) <= not(inputs(112)) or (inputs(34));
    layer0_outputs(1001) <= inputs(142);
    layer0_outputs(1002) <= (inputs(171)) xor (inputs(205));
    layer0_outputs(1003) <= (inputs(119)) xor (inputs(150));
    layer0_outputs(1004) <= (inputs(11)) xor (inputs(157));
    layer0_outputs(1005) <= '0';
    layer0_outputs(1006) <= not((inputs(73)) or (inputs(101)));
    layer0_outputs(1007) <= not(inputs(63));
    layer0_outputs(1008) <= '0';
    layer0_outputs(1009) <= '0';
    layer0_outputs(1010) <= '1';
    layer0_outputs(1011) <= not(inputs(12));
    layer0_outputs(1012) <= (inputs(114)) or (inputs(50));
    layer0_outputs(1013) <= '0';
    layer0_outputs(1014) <= (inputs(226)) xor (inputs(119));
    layer0_outputs(1015) <= not((inputs(47)) or (inputs(145)));
    layer0_outputs(1016) <= not((inputs(98)) and (inputs(14)));
    layer0_outputs(1017) <= not((inputs(250)) xor (inputs(197)));
    layer0_outputs(1018) <= not((inputs(45)) and (inputs(250)));
    layer0_outputs(1019) <= (inputs(167)) and (inputs(12));
    layer0_outputs(1020) <= (inputs(131)) and not (inputs(225));
    layer0_outputs(1021) <= not((inputs(201)) xor (inputs(232)));
    layer0_outputs(1022) <= (inputs(156)) or (inputs(205));
    layer0_outputs(1023) <= '1';
    layer0_outputs(1024) <= not((inputs(254)) and (inputs(240)));
    layer0_outputs(1025) <= (inputs(199)) and (inputs(157));
    layer0_outputs(1026) <= not(inputs(55));
    layer0_outputs(1027) <= not((inputs(203)) or (inputs(197)));
    layer0_outputs(1028) <= not(inputs(18));
    layer0_outputs(1029) <= not((inputs(145)) and (inputs(25)));
    layer0_outputs(1030) <= not(inputs(8)) or (inputs(134));
    layer0_outputs(1031) <= inputs(107);
    layer0_outputs(1032) <= not(inputs(19));
    layer0_outputs(1033) <= inputs(172);
    layer0_outputs(1034) <= (inputs(74)) and not (inputs(40));
    layer0_outputs(1035) <= inputs(226);
    layer0_outputs(1036) <= (inputs(18)) and not (inputs(185));
    layer0_outputs(1037) <= not((inputs(17)) or (inputs(150)));
    layer0_outputs(1038) <= '0';
    layer0_outputs(1039) <= (inputs(137)) and not (inputs(248));
    layer0_outputs(1040) <= not(inputs(164));
    layer0_outputs(1041) <= (inputs(146)) and not (inputs(33));
    layer0_outputs(1042) <= not(inputs(86)) or (inputs(242));
    layer0_outputs(1043) <= (inputs(85)) or (inputs(221));
    layer0_outputs(1044) <= '1';
    layer0_outputs(1045) <= not(inputs(70));
    layer0_outputs(1046) <= not(inputs(189)) or (inputs(200));
    layer0_outputs(1047) <= (inputs(240)) xor (inputs(153));
    layer0_outputs(1048) <= (inputs(102)) and not (inputs(34));
    layer0_outputs(1049) <= not(inputs(24)) or (inputs(0));
    layer0_outputs(1050) <= '0';
    layer0_outputs(1051) <= (inputs(58)) and not (inputs(32));
    layer0_outputs(1052) <= not(inputs(205));
    layer0_outputs(1053) <= (inputs(170)) or (inputs(156));
    layer0_outputs(1054) <= (inputs(60)) xor (inputs(15));
    layer0_outputs(1055) <= not(inputs(175));
    layer0_outputs(1056) <= not(inputs(244));
    layer0_outputs(1057) <= (inputs(5)) xor (inputs(220));
    layer0_outputs(1058) <= not(inputs(199)) or (inputs(247));
    layer0_outputs(1059) <= inputs(151);
    layer0_outputs(1060) <= not(inputs(81));
    layer0_outputs(1061) <= not(inputs(76)) or (inputs(78));
    layer0_outputs(1062) <= inputs(123);
    layer0_outputs(1063) <= inputs(234);
    layer0_outputs(1064) <= not((inputs(224)) or (inputs(164)));
    layer0_outputs(1065) <= '0';
    layer0_outputs(1066) <= not(inputs(140)) or (inputs(232));
    layer0_outputs(1067) <= (inputs(191)) and (inputs(114));
    layer0_outputs(1068) <= '0';
    layer0_outputs(1069) <= '0';
    layer0_outputs(1070) <= not(inputs(220)) or (inputs(89));
    layer0_outputs(1071) <= (inputs(178)) and not (inputs(129));
    layer0_outputs(1072) <= not((inputs(31)) xor (inputs(141)));
    layer0_outputs(1073) <= not(inputs(82));
    layer0_outputs(1074) <= inputs(113);
    layer0_outputs(1075) <= not(inputs(214));
    layer0_outputs(1076) <= inputs(64);
    layer0_outputs(1077) <= not((inputs(212)) xor (inputs(112)));
    layer0_outputs(1078) <= (inputs(168)) and not (inputs(120));
    layer0_outputs(1079) <= not((inputs(223)) xor (inputs(193)));
    layer0_outputs(1080) <= inputs(140);
    layer0_outputs(1081) <= not(inputs(168)) or (inputs(134));
    layer0_outputs(1082) <= not((inputs(10)) or (inputs(76)));
    layer0_outputs(1083) <= '1';
    layer0_outputs(1084) <= not((inputs(229)) or (inputs(58)));
    layer0_outputs(1085) <= (inputs(1)) and (inputs(30));
    layer0_outputs(1086) <= (inputs(153)) and not (inputs(198));
    layer0_outputs(1087) <= inputs(52);
    layer0_outputs(1088) <= inputs(189);
    layer0_outputs(1089) <= not((inputs(170)) or (inputs(40)));
    layer0_outputs(1090) <= not(inputs(24)) or (inputs(201));
    layer0_outputs(1091) <= not(inputs(43));
    layer0_outputs(1092) <= (inputs(241)) xor (inputs(204));
    layer0_outputs(1093) <= (inputs(177)) and not (inputs(210));
    layer0_outputs(1094) <= not(inputs(165)) or (inputs(40));
    layer0_outputs(1095) <= (inputs(238)) or (inputs(140));
    layer0_outputs(1096) <= inputs(85);
    layer0_outputs(1097) <= inputs(238);
    layer0_outputs(1098) <= not(inputs(24));
    layer0_outputs(1099) <= inputs(220);
    layer0_outputs(1100) <= inputs(180);
    layer0_outputs(1101) <= not(inputs(107)) or (inputs(232));
    layer0_outputs(1102) <= (inputs(32)) or (inputs(44));
    layer0_outputs(1103) <= not(inputs(123));
    layer0_outputs(1104) <= not(inputs(149));
    layer0_outputs(1105) <= (inputs(53)) and not (inputs(151));
    layer0_outputs(1106) <= '1';
    layer0_outputs(1107) <= (inputs(183)) or (inputs(223));
    layer0_outputs(1108) <= not(inputs(125));
    layer0_outputs(1109) <= inputs(166);
    layer0_outputs(1110) <= not(inputs(162)) or (inputs(4));
    layer0_outputs(1111) <= (inputs(12)) and (inputs(210));
    layer0_outputs(1112) <= not(inputs(47));
    layer0_outputs(1113) <= inputs(5);
    layer0_outputs(1114) <= (inputs(110)) or (inputs(187));
    layer0_outputs(1115) <= not((inputs(136)) and (inputs(39)));
    layer0_outputs(1116) <= not(inputs(215)) or (inputs(51));
    layer0_outputs(1117) <= not(inputs(254));
    layer0_outputs(1118) <= '0';
    layer0_outputs(1119) <= inputs(112);
    layer0_outputs(1120) <= '0';
    layer0_outputs(1121) <= not(inputs(222)) or (inputs(8));
    layer0_outputs(1122) <= (inputs(68)) and (inputs(44));
    layer0_outputs(1123) <= not((inputs(188)) or (inputs(114)));
    layer0_outputs(1124) <= not(inputs(176));
    layer0_outputs(1125) <= not(inputs(83));
    layer0_outputs(1126) <= inputs(43);
    layer0_outputs(1127) <= (inputs(24)) and (inputs(118));
    layer0_outputs(1128) <= (inputs(79)) xor (inputs(145));
    layer0_outputs(1129) <= '1';
    layer0_outputs(1130) <= '1';
    layer0_outputs(1131) <= not(inputs(157)) or (inputs(211));
    layer0_outputs(1132) <= not(inputs(46)) or (inputs(97));
    layer0_outputs(1133) <= (inputs(14)) and (inputs(185));
    layer0_outputs(1134) <= (inputs(224)) and not (inputs(99));
    layer0_outputs(1135) <= (inputs(153)) xor (inputs(254));
    layer0_outputs(1136) <= (inputs(244)) and not (inputs(46));
    layer0_outputs(1137) <= not((inputs(247)) xor (inputs(168)));
    layer0_outputs(1138) <= (inputs(153)) or (inputs(18));
    layer0_outputs(1139) <= '1';
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= inputs(31);
    layer0_outputs(1142) <= not((inputs(121)) or (inputs(83)));
    layer0_outputs(1143) <= not((inputs(135)) or (inputs(210)));
    layer0_outputs(1144) <= not((inputs(9)) xor (inputs(201)));
    layer0_outputs(1145) <= (inputs(0)) and not (inputs(230));
    layer0_outputs(1146) <= (inputs(60)) xor (inputs(100));
    layer0_outputs(1147) <= not(inputs(231)) or (inputs(51));
    layer0_outputs(1148) <= (inputs(149)) and (inputs(15));
    layer0_outputs(1149) <= (inputs(243)) xor (inputs(192));
    layer0_outputs(1150) <= (inputs(200)) and not (inputs(188));
    layer0_outputs(1151) <= inputs(121);
    layer0_outputs(1152) <= inputs(135);
    layer0_outputs(1153) <= inputs(151);
    layer0_outputs(1154) <= not((inputs(117)) or (inputs(203)));
    layer0_outputs(1155) <= not(inputs(139)) or (inputs(107));
    layer0_outputs(1156) <= not(inputs(231));
    layer0_outputs(1157) <= (inputs(63)) xor (inputs(28));
    layer0_outputs(1158) <= not((inputs(61)) and (inputs(80)));
    layer0_outputs(1159) <= (inputs(251)) and (inputs(115));
    layer0_outputs(1160) <= (inputs(151)) and not (inputs(253));
    layer0_outputs(1161) <= (inputs(102)) or (inputs(44));
    layer0_outputs(1162) <= (inputs(223)) and not (inputs(36));
    layer0_outputs(1163) <= not(inputs(125));
    layer0_outputs(1164) <= (inputs(171)) and (inputs(172));
    layer0_outputs(1165) <= (inputs(157)) or (inputs(122));
    layer0_outputs(1166) <= inputs(88);
    layer0_outputs(1167) <= '0';
    layer0_outputs(1168) <= (inputs(182)) and not (inputs(235));
    layer0_outputs(1169) <= (inputs(85)) and not (inputs(73));
    layer0_outputs(1170) <= not(inputs(27));
    layer0_outputs(1171) <= (inputs(104)) and not (inputs(15));
    layer0_outputs(1172) <= (inputs(105)) or (inputs(89));
    layer0_outputs(1173) <= '0';
    layer0_outputs(1174) <= (inputs(6)) or (inputs(166));
    layer0_outputs(1175) <= '1';
    layer0_outputs(1176) <= not(inputs(73)) or (inputs(210));
    layer0_outputs(1177) <= (inputs(217)) and (inputs(65));
    layer0_outputs(1178) <= not(inputs(50));
    layer0_outputs(1179) <= not(inputs(40));
    layer0_outputs(1180) <= (inputs(253)) xor (inputs(150));
    layer0_outputs(1181) <= (inputs(78)) or (inputs(117));
    layer0_outputs(1182) <= not(inputs(78));
    layer0_outputs(1183) <= inputs(99);
    layer0_outputs(1184) <= not(inputs(42)) or (inputs(131));
    layer0_outputs(1185) <= not(inputs(25)) or (inputs(250));
    layer0_outputs(1186) <= (inputs(1)) and (inputs(24));
    layer0_outputs(1187) <= (inputs(216)) and not (inputs(79));
    layer0_outputs(1188) <= inputs(43);
    layer0_outputs(1189) <= (inputs(110)) or (inputs(192));
    layer0_outputs(1190) <= (inputs(237)) xor (inputs(227));
    layer0_outputs(1191) <= (inputs(25)) and not (inputs(159));
    layer0_outputs(1192) <= not((inputs(114)) and (inputs(70)));
    layer0_outputs(1193) <= not(inputs(52));
    layer0_outputs(1194) <= not(inputs(145)) or (inputs(238));
    layer0_outputs(1195) <= '0';
    layer0_outputs(1196) <= not((inputs(71)) xor (inputs(75)));
    layer0_outputs(1197) <= inputs(56);
    layer0_outputs(1198) <= (inputs(204)) or (inputs(203));
    layer0_outputs(1199) <= not((inputs(216)) and (inputs(234)));
    layer0_outputs(1200) <= (inputs(191)) xor (inputs(189));
    layer0_outputs(1201) <= not(inputs(61)) or (inputs(254));
    layer0_outputs(1202) <= not(inputs(112)) or (inputs(192));
    layer0_outputs(1203) <= not(inputs(43));
    layer0_outputs(1204) <= inputs(150);
    layer0_outputs(1205) <= (inputs(90)) and not (inputs(239));
    layer0_outputs(1206) <= not(inputs(225)) or (inputs(200));
    layer0_outputs(1207) <= (inputs(48)) and not (inputs(98));
    layer0_outputs(1208) <= inputs(179);
    layer0_outputs(1209) <= (inputs(201)) or (inputs(148));
    layer0_outputs(1210) <= not(inputs(206));
    layer0_outputs(1211) <= not((inputs(56)) or (inputs(143)));
    layer0_outputs(1212) <= not((inputs(98)) xor (inputs(37)));
    layer0_outputs(1213) <= (inputs(193)) and (inputs(166));
    layer0_outputs(1214) <= (inputs(214)) and not (inputs(26));
    layer0_outputs(1215) <= '1';
    layer0_outputs(1216) <= inputs(227);
    layer0_outputs(1217) <= inputs(239);
    layer0_outputs(1218) <= '1';
    layer0_outputs(1219) <= not((inputs(44)) or (inputs(161)));
    layer0_outputs(1220) <= (inputs(251)) and not (inputs(38));
    layer0_outputs(1221) <= (inputs(193)) and not (inputs(52));
    layer0_outputs(1222) <= (inputs(29)) and not (inputs(144));
    layer0_outputs(1223) <= (inputs(155)) xor (inputs(22));
    layer0_outputs(1224) <= (inputs(104)) and not (inputs(79));
    layer0_outputs(1225) <= inputs(41);
    layer0_outputs(1226) <= not(inputs(84));
    layer0_outputs(1227) <= not(inputs(197));
    layer0_outputs(1228) <= not(inputs(151));
    layer0_outputs(1229) <= not(inputs(143)) or (inputs(119));
    layer0_outputs(1230) <= (inputs(245)) and not (inputs(198));
    layer0_outputs(1231) <= not(inputs(236)) or (inputs(202));
    layer0_outputs(1232) <= inputs(246);
    layer0_outputs(1233) <= (inputs(52)) and not (inputs(24));
    layer0_outputs(1234) <= not((inputs(172)) and (inputs(66)));
    layer0_outputs(1235) <= (inputs(235)) or (inputs(135));
    layer0_outputs(1236) <= not((inputs(176)) xor (inputs(44)));
    layer0_outputs(1237) <= not((inputs(109)) and (inputs(112)));
    layer0_outputs(1238) <= (inputs(173)) and (inputs(239));
    layer0_outputs(1239) <= (inputs(200)) xor (inputs(96));
    layer0_outputs(1240) <= not((inputs(161)) xor (inputs(25)));
    layer0_outputs(1241) <= inputs(218);
    layer0_outputs(1242) <= not((inputs(192)) xor (inputs(142)));
    layer0_outputs(1243) <= not(inputs(143)) or (inputs(3));
    layer0_outputs(1244) <= (inputs(207)) xor (inputs(103));
    layer0_outputs(1245) <= (inputs(108)) and not (inputs(253));
    layer0_outputs(1246) <= not((inputs(193)) and (inputs(5)));
    layer0_outputs(1247) <= (inputs(58)) or (inputs(38));
    layer0_outputs(1248) <= not(inputs(220));
    layer0_outputs(1249) <= not((inputs(237)) or (inputs(90)));
    layer0_outputs(1250) <= (inputs(197)) or (inputs(83));
    layer0_outputs(1251) <= inputs(168);
    layer0_outputs(1252) <= not(inputs(240));
    layer0_outputs(1253) <= not((inputs(182)) or (inputs(164)));
    layer0_outputs(1254) <= (inputs(111)) xor (inputs(215));
    layer0_outputs(1255) <= (inputs(48)) or (inputs(147));
    layer0_outputs(1256) <= (inputs(126)) xor (inputs(93));
    layer0_outputs(1257) <= not(inputs(215));
    layer0_outputs(1258) <= (inputs(90)) or (inputs(126));
    layer0_outputs(1259) <= not((inputs(147)) or (inputs(184)));
    layer0_outputs(1260) <= (inputs(239)) xor (inputs(78));
    layer0_outputs(1261) <= '0';
    layer0_outputs(1262) <= (inputs(73)) or (inputs(130));
    layer0_outputs(1263) <= not((inputs(111)) and (inputs(126)));
    layer0_outputs(1264) <= inputs(137);
    layer0_outputs(1265) <= not(inputs(92));
    layer0_outputs(1266) <= (inputs(170)) and not (inputs(75));
    layer0_outputs(1267) <= (inputs(17)) or (inputs(3));
    layer0_outputs(1268) <= inputs(182);
    layer0_outputs(1269) <= (inputs(88)) and (inputs(83));
    layer0_outputs(1270) <= '0';
    layer0_outputs(1271) <= inputs(136);
    layer0_outputs(1272) <= (inputs(159)) and not (inputs(228));
    layer0_outputs(1273) <= (inputs(216)) or (inputs(94));
    layer0_outputs(1274) <= (inputs(138)) xor (inputs(41));
    layer0_outputs(1275) <= (inputs(27)) and not (inputs(77));
    layer0_outputs(1276) <= '1';
    layer0_outputs(1277) <= (inputs(33)) and not (inputs(38));
    layer0_outputs(1278) <= (inputs(187)) and not (inputs(18));
    layer0_outputs(1279) <= not(inputs(213)) or (inputs(80));
    layer0_outputs(1280) <= inputs(52);
    layer0_outputs(1281) <= (inputs(34)) or (inputs(230));
    layer0_outputs(1282) <= not((inputs(234)) or (inputs(132)));
    layer0_outputs(1283) <= (inputs(166)) xor (inputs(0));
    layer0_outputs(1284) <= '0';
    layer0_outputs(1285) <= (inputs(97)) and (inputs(89));
    layer0_outputs(1286) <= not(inputs(136));
    layer0_outputs(1287) <= inputs(3);
    layer0_outputs(1288) <= inputs(1);
    layer0_outputs(1289) <= (inputs(221)) or (inputs(32));
    layer0_outputs(1290) <= not(inputs(233)) or (inputs(54));
    layer0_outputs(1291) <= (inputs(156)) xor (inputs(2));
    layer0_outputs(1292) <= not(inputs(61));
    layer0_outputs(1293) <= not(inputs(146));
    layer0_outputs(1294) <= (inputs(162)) or (inputs(34));
    layer0_outputs(1295) <= not(inputs(77));
    layer0_outputs(1296) <= inputs(12);
    layer0_outputs(1297) <= '1';
    layer0_outputs(1298) <= not(inputs(209)) or (inputs(41));
    layer0_outputs(1299) <= (inputs(255)) xor (inputs(18));
    layer0_outputs(1300) <= (inputs(11)) or (inputs(208));
    layer0_outputs(1301) <= not((inputs(186)) or (inputs(116)));
    layer0_outputs(1302) <= (inputs(99)) and not (inputs(36));
    layer0_outputs(1303) <= inputs(148);
    layer0_outputs(1304) <= inputs(116);
    layer0_outputs(1305) <= not((inputs(37)) xor (inputs(209)));
    layer0_outputs(1306) <= inputs(156);
    layer0_outputs(1307) <= not((inputs(178)) or (inputs(140)));
    layer0_outputs(1308) <= (inputs(67)) and not (inputs(38));
    layer0_outputs(1309) <= not(inputs(158)) or (inputs(255));
    layer0_outputs(1310) <= not(inputs(36));
    layer0_outputs(1311) <= not(inputs(254)) or (inputs(26));
    layer0_outputs(1312) <= not(inputs(113));
    layer0_outputs(1313) <= (inputs(184)) xor (inputs(243));
    layer0_outputs(1314) <= (inputs(151)) and not (inputs(7));
    layer0_outputs(1315) <= not(inputs(87)) or (inputs(221));
    layer0_outputs(1316) <= (inputs(104)) and not (inputs(92));
    layer0_outputs(1317) <= not(inputs(223)) or (inputs(110));
    layer0_outputs(1318) <= not(inputs(184)) or (inputs(225));
    layer0_outputs(1319) <= (inputs(110)) and not (inputs(107));
    layer0_outputs(1320) <= (inputs(106)) or (inputs(145));
    layer0_outputs(1321) <= (inputs(116)) and not (inputs(117));
    layer0_outputs(1322) <= (inputs(48)) xor (inputs(16));
    layer0_outputs(1323) <= (inputs(60)) xor (inputs(66));
    layer0_outputs(1324) <= (inputs(91)) or (inputs(145));
    layer0_outputs(1325) <= (inputs(94)) and not (inputs(189));
    layer0_outputs(1326) <= not(inputs(159));
    layer0_outputs(1327) <= (inputs(2)) or (inputs(87));
    layer0_outputs(1328) <= not(inputs(4)) or (inputs(81));
    layer0_outputs(1329) <= (inputs(59)) and not (inputs(62));
    layer0_outputs(1330) <= (inputs(199)) xor (inputs(113));
    layer0_outputs(1331) <= not(inputs(190));
    layer0_outputs(1332) <= '0';
    layer0_outputs(1333) <= not(inputs(79)) or (inputs(225));
    layer0_outputs(1334) <= not(inputs(92));
    layer0_outputs(1335) <= (inputs(102)) or (inputs(94));
    layer0_outputs(1336) <= not((inputs(51)) or (inputs(37)));
    layer0_outputs(1337) <= inputs(77);
    layer0_outputs(1338) <= (inputs(211)) xor (inputs(186));
    layer0_outputs(1339) <= '1';
    layer0_outputs(1340) <= '1';
    layer0_outputs(1341) <= '0';
    layer0_outputs(1342) <= not(inputs(120)) or (inputs(44));
    layer0_outputs(1343) <= inputs(149);
    layer0_outputs(1344) <= (inputs(128)) and (inputs(230));
    layer0_outputs(1345) <= (inputs(40)) or (inputs(53));
    layer0_outputs(1346) <= not((inputs(194)) and (inputs(220)));
    layer0_outputs(1347) <= not(inputs(119));
    layer0_outputs(1348) <= inputs(11);
    layer0_outputs(1349) <= not((inputs(24)) or (inputs(25)));
    layer0_outputs(1350) <= not(inputs(220)) or (inputs(177));
    layer0_outputs(1351) <= inputs(70);
    layer0_outputs(1352) <= (inputs(235)) or (inputs(11));
    layer0_outputs(1353) <= not(inputs(49));
    layer0_outputs(1354) <= inputs(192);
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= not(inputs(103)) or (inputs(178));
    layer0_outputs(1357) <= inputs(64);
    layer0_outputs(1358) <= (inputs(34)) and not (inputs(60));
    layer0_outputs(1359) <= not(inputs(108));
    layer0_outputs(1360) <= (inputs(51)) or (inputs(170));
    layer0_outputs(1361) <= (inputs(247)) or (inputs(116));
    layer0_outputs(1362) <= not((inputs(255)) and (inputs(27)));
    layer0_outputs(1363) <= not((inputs(188)) and (inputs(142)));
    layer0_outputs(1364) <= not((inputs(9)) and (inputs(46)));
    layer0_outputs(1365) <= inputs(106);
    layer0_outputs(1366) <= not((inputs(47)) or (inputs(222)));
    layer0_outputs(1367) <= '0';
    layer0_outputs(1368) <= '0';
    layer0_outputs(1369) <= not(inputs(220));
    layer0_outputs(1370) <= inputs(147);
    layer0_outputs(1371) <= '1';
    layer0_outputs(1372) <= (inputs(249)) or (inputs(229));
    layer0_outputs(1373) <= not(inputs(159)) or (inputs(155));
    layer0_outputs(1374) <= not((inputs(233)) and (inputs(110)));
    layer0_outputs(1375) <= '0';
    layer0_outputs(1376) <= not((inputs(160)) or (inputs(66)));
    layer0_outputs(1377) <= (inputs(89)) and (inputs(158));
    layer0_outputs(1378) <= not((inputs(39)) xor (inputs(128)));
    layer0_outputs(1379) <= not((inputs(97)) or (inputs(231)));
    layer0_outputs(1380) <= (inputs(207)) or (inputs(157));
    layer0_outputs(1381) <= not((inputs(147)) or (inputs(109)));
    layer0_outputs(1382) <= not(inputs(132));
    layer0_outputs(1383) <= not((inputs(45)) or (inputs(87)));
    layer0_outputs(1384) <= inputs(119);
    layer0_outputs(1385) <= not(inputs(115));
    layer0_outputs(1386) <= '0';
    layer0_outputs(1387) <= not(inputs(167));
    layer0_outputs(1388) <= (inputs(118)) or (inputs(237));
    layer0_outputs(1389) <= (inputs(122)) or (inputs(15));
    layer0_outputs(1390) <= '0';
    layer0_outputs(1391) <= not(inputs(70)) or (inputs(135));
    layer0_outputs(1392) <= (inputs(15)) and not (inputs(226));
    layer0_outputs(1393) <= not(inputs(105)) or (inputs(99));
    layer0_outputs(1394) <= inputs(42);
    layer0_outputs(1395) <= not(inputs(89));
    layer0_outputs(1396) <= not((inputs(191)) and (inputs(100)));
    layer0_outputs(1397) <= not(inputs(7)) or (inputs(27));
    layer0_outputs(1398) <= (inputs(21)) and (inputs(133));
    layer0_outputs(1399) <= (inputs(116)) and not (inputs(70));
    layer0_outputs(1400) <= (inputs(126)) or (inputs(6));
    layer0_outputs(1401) <= (inputs(173)) and (inputs(193));
    layer0_outputs(1402) <= not((inputs(67)) or (inputs(246)));
    layer0_outputs(1403) <= not(inputs(71)) or (inputs(125));
    layer0_outputs(1404) <= '0';
    layer0_outputs(1405) <= '0';
    layer0_outputs(1406) <= (inputs(140)) and (inputs(22));
    layer0_outputs(1407) <= (inputs(84)) or (inputs(108));
    layer0_outputs(1408) <= not((inputs(132)) or (inputs(138)));
    layer0_outputs(1409) <= '1';
    layer0_outputs(1410) <= not((inputs(161)) or (inputs(138)));
    layer0_outputs(1411) <= (inputs(96)) and not (inputs(255));
    layer0_outputs(1412) <= '1';
    layer0_outputs(1413) <= not(inputs(172));
    layer0_outputs(1414) <= '1';
    layer0_outputs(1415) <= '1';
    layer0_outputs(1416) <= (inputs(123)) and not (inputs(37));
    layer0_outputs(1417) <= (inputs(41)) and not (inputs(254));
    layer0_outputs(1418) <= not(inputs(239));
    layer0_outputs(1419) <= (inputs(65)) and not (inputs(83));
    layer0_outputs(1420) <= (inputs(102)) and not (inputs(250));
    layer0_outputs(1421) <= (inputs(144)) and (inputs(178));
    layer0_outputs(1422) <= not(inputs(132));
    layer0_outputs(1423) <= not((inputs(181)) xor (inputs(159)));
    layer0_outputs(1424) <= (inputs(114)) and not (inputs(83));
    layer0_outputs(1425) <= not((inputs(116)) xor (inputs(114)));
    layer0_outputs(1426) <= inputs(174);
    layer0_outputs(1427) <= (inputs(244)) xor (inputs(159));
    layer0_outputs(1428) <= not(inputs(64));
    layer0_outputs(1429) <= (inputs(66)) and (inputs(59));
    layer0_outputs(1430) <= not(inputs(108)) or (inputs(8));
    layer0_outputs(1431) <= not(inputs(150)) or (inputs(224));
    layer0_outputs(1432) <= not(inputs(236)) or (inputs(83));
    layer0_outputs(1433) <= not(inputs(58)) or (inputs(95));
    layer0_outputs(1434) <= not(inputs(29)) or (inputs(154));
    layer0_outputs(1435) <= not(inputs(112)) or (inputs(0));
    layer0_outputs(1436) <= not(inputs(125)) or (inputs(26));
    layer0_outputs(1437) <= (inputs(214)) xor (inputs(78));
    layer0_outputs(1438) <= not((inputs(106)) and (inputs(188)));
    layer0_outputs(1439) <= '0';
    layer0_outputs(1440) <= (inputs(104)) and not (inputs(232));
    layer0_outputs(1441) <= not((inputs(25)) xor (inputs(152)));
    layer0_outputs(1442) <= not(inputs(91));
    layer0_outputs(1443) <= '0';
    layer0_outputs(1444) <= not(inputs(65));
    layer0_outputs(1445) <= not(inputs(34));
    layer0_outputs(1446) <= not((inputs(188)) and (inputs(4)));
    layer0_outputs(1447) <= not(inputs(178));
    layer0_outputs(1448) <= not(inputs(235));
    layer0_outputs(1449) <= inputs(225);
    layer0_outputs(1450) <= not(inputs(238)) or (inputs(193));
    layer0_outputs(1451) <= (inputs(235)) or (inputs(214));
    layer0_outputs(1452) <= not(inputs(128));
    layer0_outputs(1453) <= inputs(239);
    layer0_outputs(1454) <= (inputs(121)) xor (inputs(232));
    layer0_outputs(1455) <= not((inputs(245)) or (inputs(49)));
    layer0_outputs(1456) <= (inputs(13)) and (inputs(64));
    layer0_outputs(1457) <= '0';
    layer0_outputs(1458) <= not(inputs(36)) or (inputs(90));
    layer0_outputs(1459) <= not(inputs(215));
    layer0_outputs(1460) <= inputs(1);
    layer0_outputs(1461) <= not((inputs(121)) or (inputs(98)));
    layer0_outputs(1462) <= (inputs(63)) and not (inputs(246));
    layer0_outputs(1463) <= not(inputs(130));
    layer0_outputs(1464) <= (inputs(203)) and not (inputs(139));
    layer0_outputs(1465) <= not(inputs(164));
    layer0_outputs(1466) <= inputs(76);
    layer0_outputs(1467) <= not((inputs(173)) xor (inputs(170)));
    layer0_outputs(1468) <= inputs(149);
    layer0_outputs(1469) <= not(inputs(68)) or (inputs(210));
    layer0_outputs(1470) <= not(inputs(165));
    layer0_outputs(1471) <= (inputs(184)) and not (inputs(144));
    layer0_outputs(1472) <= (inputs(29)) xor (inputs(221));
    layer0_outputs(1473) <= not((inputs(39)) and (inputs(55)));
    layer0_outputs(1474) <= not(inputs(70));
    layer0_outputs(1475) <= '1';
    layer0_outputs(1476) <= not(inputs(196)) or (inputs(229));
    layer0_outputs(1477) <= not(inputs(128));
    layer0_outputs(1478) <= '1';
    layer0_outputs(1479) <= not((inputs(49)) xor (inputs(13)));
    layer0_outputs(1480) <= (inputs(102)) and not (inputs(205));
    layer0_outputs(1481) <= not(inputs(154));
    layer0_outputs(1482) <= (inputs(168)) and (inputs(143));
    layer0_outputs(1483) <= (inputs(120)) or (inputs(182));
    layer0_outputs(1484) <= (inputs(206)) xor (inputs(196));
    layer0_outputs(1485) <= inputs(133);
    layer0_outputs(1486) <= (inputs(0)) or (inputs(110));
    layer0_outputs(1487) <= not((inputs(190)) xor (inputs(140)));
    layer0_outputs(1488) <= (inputs(98)) xor (inputs(218));
    layer0_outputs(1489) <= inputs(205);
    layer0_outputs(1490) <= inputs(213);
    layer0_outputs(1491) <= inputs(193);
    layer0_outputs(1492) <= not(inputs(224)) or (inputs(247));
    layer0_outputs(1493) <= (inputs(46)) and not (inputs(9));
    layer0_outputs(1494) <= '0';
    layer0_outputs(1495) <= not((inputs(64)) and (inputs(243)));
    layer0_outputs(1496) <= not((inputs(168)) or (inputs(249)));
    layer0_outputs(1497) <= not(inputs(30)) or (inputs(112));
    layer0_outputs(1498) <= inputs(93);
    layer0_outputs(1499) <= (inputs(164)) and not (inputs(100));
    layer0_outputs(1500) <= inputs(135);
    layer0_outputs(1501) <= not((inputs(48)) or (inputs(46)));
    layer0_outputs(1502) <= inputs(127);
    layer0_outputs(1503) <= not((inputs(212)) or (inputs(33)));
    layer0_outputs(1504) <= not((inputs(191)) xor (inputs(125)));
    layer0_outputs(1505) <= not((inputs(109)) and (inputs(246)));
    layer0_outputs(1506) <= (inputs(204)) and not (inputs(131));
    layer0_outputs(1507) <= not((inputs(203)) and (inputs(175)));
    layer0_outputs(1508) <= not(inputs(204));
    layer0_outputs(1509) <= not(inputs(19));
    layer0_outputs(1510) <= not(inputs(201)) or (inputs(211));
    layer0_outputs(1511) <= (inputs(100)) or (inputs(174));
    layer0_outputs(1512) <= not(inputs(77));
    layer0_outputs(1513) <= not(inputs(188));
    layer0_outputs(1514) <= (inputs(248)) and not (inputs(35));
    layer0_outputs(1515) <= not(inputs(192)) or (inputs(134));
    layer0_outputs(1516) <= not((inputs(166)) or (inputs(176)));
    layer0_outputs(1517) <= inputs(74);
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= not((inputs(66)) xor (inputs(231)));
    layer0_outputs(1520) <= (inputs(105)) and not (inputs(83));
    layer0_outputs(1521) <= not(inputs(17));
    layer0_outputs(1522) <= inputs(230);
    layer0_outputs(1523) <= not(inputs(187)) or (inputs(24));
    layer0_outputs(1524) <= '1';
    layer0_outputs(1525) <= (inputs(119)) and (inputs(155));
    layer0_outputs(1526) <= inputs(171);
    layer0_outputs(1527) <= not(inputs(195)) or (inputs(216));
    layer0_outputs(1528) <= '1';
    layer0_outputs(1529) <= not(inputs(16));
    layer0_outputs(1530) <= (inputs(167)) and not (inputs(17));
    layer0_outputs(1531) <= (inputs(48)) and (inputs(171));
    layer0_outputs(1532) <= (inputs(56)) and not (inputs(30));
    layer0_outputs(1533) <= not(inputs(14)) or (inputs(24));
    layer0_outputs(1534) <= not((inputs(94)) and (inputs(192)));
    layer0_outputs(1535) <= (inputs(216)) and (inputs(73));
    layer0_outputs(1536) <= '1';
    layer0_outputs(1537) <= (inputs(46)) xor (inputs(132));
    layer0_outputs(1538) <= inputs(93);
    layer0_outputs(1539) <= (inputs(144)) and (inputs(210));
    layer0_outputs(1540) <= (inputs(210)) and not (inputs(99));
    layer0_outputs(1541) <= (inputs(33)) or (inputs(104));
    layer0_outputs(1542) <= (inputs(4)) xor (inputs(99));
    layer0_outputs(1543) <= (inputs(111)) or (inputs(181));
    layer0_outputs(1544) <= (inputs(139)) or (inputs(68));
    layer0_outputs(1545) <= (inputs(206)) and (inputs(25));
    layer0_outputs(1546) <= inputs(161);
    layer0_outputs(1547) <= '0';
    layer0_outputs(1548) <= not((inputs(70)) or (inputs(99)));
    layer0_outputs(1549) <= (inputs(29)) and not (inputs(189));
    layer0_outputs(1550) <= not((inputs(164)) xor (inputs(141)));
    layer0_outputs(1551) <= not(inputs(141));
    layer0_outputs(1552) <= (inputs(131)) and not (inputs(194));
    layer0_outputs(1553) <= (inputs(237)) and (inputs(178));
    layer0_outputs(1554) <= (inputs(20)) and not (inputs(218));
    layer0_outputs(1555) <= inputs(18);
    layer0_outputs(1556) <= inputs(183);
    layer0_outputs(1557) <= not(inputs(230)) or (inputs(21));
    layer0_outputs(1558) <= not(inputs(9));
    layer0_outputs(1559) <= not((inputs(120)) xor (inputs(92)));
    layer0_outputs(1560) <= (inputs(197)) or (inputs(14));
    layer0_outputs(1561) <= not((inputs(180)) or (inputs(181)));
    layer0_outputs(1562) <= not(inputs(152));
    layer0_outputs(1563) <= not((inputs(36)) and (inputs(219)));
    layer0_outputs(1564) <= (inputs(246)) and not (inputs(86));
    layer0_outputs(1565) <= not(inputs(223)) or (inputs(161));
    layer0_outputs(1566) <= not(inputs(130));
    layer0_outputs(1567) <= not(inputs(2));
    layer0_outputs(1568) <= (inputs(82)) and (inputs(157));
    layer0_outputs(1569) <= inputs(137);
    layer0_outputs(1570) <= inputs(105);
    layer0_outputs(1571) <= '1';
    layer0_outputs(1572) <= not((inputs(58)) or (inputs(4)));
    layer0_outputs(1573) <= (inputs(127)) xor (inputs(17));
    layer0_outputs(1574) <= not((inputs(202)) xor (inputs(85)));
    layer0_outputs(1575) <= (inputs(209)) xor (inputs(164));
    layer0_outputs(1576) <= not(inputs(112));
    layer0_outputs(1577) <= not(inputs(120));
    layer0_outputs(1578) <= '1';
    layer0_outputs(1579) <= not((inputs(11)) or (inputs(168)));
    layer0_outputs(1580) <= not((inputs(196)) or (inputs(96)));
    layer0_outputs(1581) <= '1';
    layer0_outputs(1582) <= inputs(181);
    layer0_outputs(1583) <= (inputs(225)) or (inputs(161));
    layer0_outputs(1584) <= (inputs(138)) and not (inputs(105));
    layer0_outputs(1585) <= inputs(87);
    layer0_outputs(1586) <= inputs(100);
    layer0_outputs(1587) <= not(inputs(118));
    layer0_outputs(1588) <= not((inputs(126)) or (inputs(180)));
    layer0_outputs(1589) <= (inputs(246)) or (inputs(34));
    layer0_outputs(1590) <= inputs(34);
    layer0_outputs(1591) <= (inputs(186)) or (inputs(177));
    layer0_outputs(1592) <= not(inputs(178));
    layer0_outputs(1593) <= not(inputs(17));
    layer0_outputs(1594) <= not(inputs(74)) or (inputs(57));
    layer0_outputs(1595) <= not(inputs(195)) or (inputs(135));
    layer0_outputs(1596) <= not(inputs(231)) or (inputs(217));
    layer0_outputs(1597) <= '0';
    layer0_outputs(1598) <= not((inputs(29)) or (inputs(166)));
    layer0_outputs(1599) <= not((inputs(255)) xor (inputs(77)));
    layer0_outputs(1600) <= (inputs(43)) or (inputs(85));
    layer0_outputs(1601) <= inputs(83);
    layer0_outputs(1602) <= (inputs(234)) and not (inputs(97));
    layer0_outputs(1603) <= not(inputs(213)) or (inputs(13));
    layer0_outputs(1604) <= not(inputs(5)) or (inputs(255));
    layer0_outputs(1605) <= inputs(217);
    layer0_outputs(1606) <= not(inputs(30)) or (inputs(96));
    layer0_outputs(1607) <= inputs(94);
    layer0_outputs(1608) <= not((inputs(211)) and (inputs(200)));
    layer0_outputs(1609) <= not(inputs(247)) or (inputs(52));
    layer0_outputs(1610) <= '0';
    layer0_outputs(1611) <= not(inputs(59)) or (inputs(168));
    layer0_outputs(1612) <= not((inputs(209)) or (inputs(61)));
    layer0_outputs(1613) <= (inputs(198)) and (inputs(105));
    layer0_outputs(1614) <= not((inputs(33)) or (inputs(160)));
    layer0_outputs(1615) <= not(inputs(23)) or (inputs(202));
    layer0_outputs(1616) <= (inputs(131)) and not (inputs(68));
    layer0_outputs(1617) <= (inputs(195)) and (inputs(3));
    layer0_outputs(1618) <= not((inputs(239)) or (inputs(95)));
    layer0_outputs(1619) <= '1';
    layer0_outputs(1620) <= not(inputs(133)) or (inputs(187));
    layer0_outputs(1621) <= not(inputs(180));
    layer0_outputs(1622) <= (inputs(247)) and not (inputs(221));
    layer0_outputs(1623) <= (inputs(58)) and not (inputs(34));
    layer0_outputs(1624) <= inputs(175);
    layer0_outputs(1625) <= not(inputs(164)) or (inputs(244));
    layer0_outputs(1626) <= inputs(205);
    layer0_outputs(1627) <= (inputs(139)) or (inputs(14));
    layer0_outputs(1628) <= (inputs(1)) xor (inputs(69));
    layer0_outputs(1629) <= (inputs(14)) and not (inputs(76));
    layer0_outputs(1630) <= not((inputs(110)) or (inputs(121)));
    layer0_outputs(1631) <= not(inputs(183)) or (inputs(73));
    layer0_outputs(1632) <= inputs(190);
    layer0_outputs(1633) <= not(inputs(58));
    layer0_outputs(1634) <= (inputs(102)) and not (inputs(221));
    layer0_outputs(1635) <= not((inputs(72)) xor (inputs(195)));
    layer0_outputs(1636) <= (inputs(159)) and (inputs(179));
    layer0_outputs(1637) <= inputs(104);
    layer0_outputs(1638) <= (inputs(254)) xor (inputs(6));
    layer0_outputs(1639) <= (inputs(27)) and (inputs(195));
    layer0_outputs(1640) <= not(inputs(245)) or (inputs(15));
    layer0_outputs(1641) <= (inputs(185)) or (inputs(131));
    layer0_outputs(1642) <= not((inputs(41)) or (inputs(189)));
    layer0_outputs(1643) <= not((inputs(57)) or (inputs(159)));
    layer0_outputs(1644) <= inputs(64);
    layer0_outputs(1645) <= not((inputs(215)) and (inputs(152)));
    layer0_outputs(1646) <= not((inputs(142)) xor (inputs(144)));
    layer0_outputs(1647) <= not(inputs(197)) or (inputs(244));
    layer0_outputs(1648) <= not(inputs(130)) or (inputs(104));
    layer0_outputs(1649) <= (inputs(164)) and (inputs(57));
    layer0_outputs(1650) <= (inputs(253)) xor (inputs(186));
    layer0_outputs(1651) <= (inputs(124)) and not (inputs(177));
    layer0_outputs(1652) <= '1';
    layer0_outputs(1653) <= (inputs(125)) xor (inputs(174));
    layer0_outputs(1654) <= '1';
    layer0_outputs(1655) <= not(inputs(188)) or (inputs(91));
    layer0_outputs(1656) <= (inputs(70)) or (inputs(120));
    layer0_outputs(1657) <= not(inputs(110)) or (inputs(245));
    layer0_outputs(1658) <= (inputs(2)) and not (inputs(127));
    layer0_outputs(1659) <= (inputs(221)) and not (inputs(25));
    layer0_outputs(1660) <= not(inputs(144)) or (inputs(141));
    layer0_outputs(1661) <= (inputs(96)) and (inputs(6));
    layer0_outputs(1662) <= not((inputs(173)) and (inputs(214)));
    layer0_outputs(1663) <= not((inputs(100)) and (inputs(21)));
    layer0_outputs(1664) <= (inputs(204)) or (inputs(212));
    layer0_outputs(1665) <= not((inputs(47)) and (inputs(82)));
    layer0_outputs(1666) <= not((inputs(231)) xor (inputs(230)));
    layer0_outputs(1667) <= (inputs(185)) and not (inputs(66));
    layer0_outputs(1668) <= not((inputs(9)) xor (inputs(33)));
    layer0_outputs(1669) <= not(inputs(153));
    layer0_outputs(1670) <= (inputs(157)) or (inputs(11));
    layer0_outputs(1671) <= not((inputs(205)) xor (inputs(50)));
    layer0_outputs(1672) <= not(inputs(235)) or (inputs(253));
    layer0_outputs(1673) <= (inputs(230)) or (inputs(121));
    layer0_outputs(1674) <= not((inputs(95)) and (inputs(119)));
    layer0_outputs(1675) <= not(inputs(112)) or (inputs(163));
    layer0_outputs(1676) <= (inputs(129)) and not (inputs(49));
    layer0_outputs(1677) <= '0';
    layer0_outputs(1678) <= not((inputs(250)) or (inputs(90)));
    layer0_outputs(1679) <= '0';
    layer0_outputs(1680) <= (inputs(183)) xor (inputs(143));
    layer0_outputs(1681) <= inputs(208);
    layer0_outputs(1682) <= (inputs(209)) and not (inputs(133));
    layer0_outputs(1683) <= not((inputs(39)) xor (inputs(41)));
    layer0_outputs(1684) <= not((inputs(94)) xor (inputs(50)));
    layer0_outputs(1685) <= not((inputs(22)) xor (inputs(234)));
    layer0_outputs(1686) <= not((inputs(105)) xor (inputs(231)));
    layer0_outputs(1687) <= not(inputs(133));
    layer0_outputs(1688) <= not(inputs(200)) or (inputs(233));
    layer0_outputs(1689) <= inputs(96);
    layer0_outputs(1690) <= not((inputs(190)) and (inputs(13)));
    layer0_outputs(1691) <= inputs(22);
    layer0_outputs(1692) <= not((inputs(242)) or (inputs(147)));
    layer0_outputs(1693) <= not((inputs(89)) or (inputs(57)));
    layer0_outputs(1694) <= '0';
    layer0_outputs(1695) <= not(inputs(107)) or (inputs(26));
    layer0_outputs(1696) <= not((inputs(85)) and (inputs(83)));
    layer0_outputs(1697) <= inputs(190);
    layer0_outputs(1698) <= (inputs(109)) xor (inputs(244));
    layer0_outputs(1699) <= inputs(220);
    layer0_outputs(1700) <= not(inputs(49));
    layer0_outputs(1701) <= (inputs(88)) and not (inputs(80));
    layer0_outputs(1702) <= '0';
    layer0_outputs(1703) <= (inputs(99)) and (inputs(15));
    layer0_outputs(1704) <= '0';
    layer0_outputs(1705) <= '0';
    layer0_outputs(1706) <= (inputs(241)) xor (inputs(214));
    layer0_outputs(1707) <= not(inputs(8)) or (inputs(175));
    layer0_outputs(1708) <= inputs(85);
    layer0_outputs(1709) <= not(inputs(70)) or (inputs(123));
    layer0_outputs(1710) <= (inputs(122)) and (inputs(9));
    layer0_outputs(1711) <= '0';
    layer0_outputs(1712) <= '1';
    layer0_outputs(1713) <= '0';
    layer0_outputs(1714) <= not(inputs(194));
    layer0_outputs(1715) <= '0';
    layer0_outputs(1716) <= not(inputs(68)) or (inputs(8));
    layer0_outputs(1717) <= not(inputs(121));
    layer0_outputs(1718) <= not(inputs(188)) or (inputs(233));
    layer0_outputs(1719) <= (inputs(87)) and (inputs(115));
    layer0_outputs(1720) <= (inputs(159)) and not (inputs(191));
    layer0_outputs(1721) <= inputs(147);
    layer0_outputs(1722) <= inputs(231);
    layer0_outputs(1723) <= not(inputs(207));
    layer0_outputs(1724) <= inputs(73);
    layer0_outputs(1725) <= inputs(180);
    layer0_outputs(1726) <= (inputs(67)) and not (inputs(47));
    layer0_outputs(1727) <= (inputs(83)) or (inputs(51));
    layer0_outputs(1728) <= not(inputs(118)) or (inputs(240));
    layer0_outputs(1729) <= (inputs(53)) or (inputs(64));
    layer0_outputs(1730) <= (inputs(146)) or (inputs(105));
    layer0_outputs(1731) <= not(inputs(202));
    layer0_outputs(1732) <= not((inputs(60)) or (inputs(72)));
    layer0_outputs(1733) <= not(inputs(124)) or (inputs(16));
    layer0_outputs(1734) <= (inputs(64)) or (inputs(36));
    layer0_outputs(1735) <= not(inputs(226)) or (inputs(196));
    layer0_outputs(1736) <= not(inputs(117));
    layer0_outputs(1737) <= not(inputs(248));
    layer0_outputs(1738) <= not(inputs(59)) or (inputs(160));
    layer0_outputs(1739) <= inputs(214);
    layer0_outputs(1740) <= inputs(197);
    layer0_outputs(1741) <= inputs(72);
    layer0_outputs(1742) <= not((inputs(117)) and (inputs(66)));
    layer0_outputs(1743) <= not(inputs(183)) or (inputs(203));
    layer0_outputs(1744) <= '1';
    layer0_outputs(1745) <= not(inputs(15)) or (inputs(100));
    layer0_outputs(1746) <= (inputs(76)) or (inputs(134));
    layer0_outputs(1747) <= '1';
    layer0_outputs(1748) <= (inputs(142)) and (inputs(220));
    layer0_outputs(1749) <= not(inputs(219)) or (inputs(229));
    layer0_outputs(1750) <= not((inputs(76)) or (inputs(78)));
    layer0_outputs(1751) <= not(inputs(87)) or (inputs(127));
    layer0_outputs(1752) <= not((inputs(96)) and (inputs(72)));
    layer0_outputs(1753) <= not((inputs(150)) or (inputs(106)));
    layer0_outputs(1754) <= (inputs(247)) or (inputs(73));
    layer0_outputs(1755) <= not((inputs(143)) xor (inputs(212)));
    layer0_outputs(1756) <= '1';
    layer0_outputs(1757) <= not((inputs(61)) or (inputs(101)));
    layer0_outputs(1758) <= (inputs(44)) and not (inputs(202));
    layer0_outputs(1759) <= inputs(124);
    layer0_outputs(1760) <= (inputs(116)) and not (inputs(235));
    layer0_outputs(1761) <= (inputs(40)) or (inputs(194));
    layer0_outputs(1762) <= not((inputs(40)) or (inputs(204)));
    layer0_outputs(1763) <= not(inputs(168)) or (inputs(225));
    layer0_outputs(1764) <= (inputs(84)) xor (inputs(186));
    layer0_outputs(1765) <= not((inputs(53)) xor (inputs(100)));
    layer0_outputs(1766) <= (inputs(205)) and not (inputs(170));
    layer0_outputs(1767) <= not((inputs(169)) or (inputs(229)));
    layer0_outputs(1768) <= not(inputs(22));
    layer0_outputs(1769) <= not((inputs(248)) and (inputs(225)));
    layer0_outputs(1770) <= not(inputs(244)) or (inputs(28));
    layer0_outputs(1771) <= not(inputs(242)) or (inputs(70));
    layer0_outputs(1772) <= (inputs(243)) or (inputs(54));
    layer0_outputs(1773) <= (inputs(88)) and not (inputs(148));
    layer0_outputs(1774) <= inputs(187);
    layer0_outputs(1775) <= inputs(255);
    layer0_outputs(1776) <= not((inputs(233)) and (inputs(94)));
    layer0_outputs(1777) <= (inputs(144)) or (inputs(161));
    layer0_outputs(1778) <= not(inputs(215)) or (inputs(175));
    layer0_outputs(1779) <= inputs(208);
    layer0_outputs(1780) <= inputs(27);
    layer0_outputs(1781) <= not(inputs(57));
    layer0_outputs(1782) <= not(inputs(61)) or (inputs(58));
    layer0_outputs(1783) <= not(inputs(10)) or (inputs(204));
    layer0_outputs(1784) <= not(inputs(180));
    layer0_outputs(1785) <= not((inputs(197)) or (inputs(35)));
    layer0_outputs(1786) <= not(inputs(234));
    layer0_outputs(1787) <= not(inputs(182));
    layer0_outputs(1788) <= not((inputs(105)) or (inputs(159)));
    layer0_outputs(1789) <= not(inputs(208));
    layer0_outputs(1790) <= not((inputs(41)) or (inputs(44)));
    layer0_outputs(1791) <= (inputs(201)) and not (inputs(35));
    layer0_outputs(1792) <= inputs(45);
    layer0_outputs(1793) <= (inputs(226)) or (inputs(242));
    layer0_outputs(1794) <= not((inputs(34)) and (inputs(78)));
    layer0_outputs(1795) <= (inputs(57)) and (inputs(3));
    layer0_outputs(1796) <= not(inputs(177));
    layer0_outputs(1797) <= not(inputs(36)) or (inputs(103));
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= not((inputs(75)) xor (inputs(35)));
    layer0_outputs(1800) <= not((inputs(31)) or (inputs(2)));
    layer0_outputs(1801) <= (inputs(69)) and not (inputs(200));
    layer0_outputs(1802) <= not((inputs(156)) and (inputs(21)));
    layer0_outputs(1803) <= not((inputs(25)) xor (inputs(49)));
    layer0_outputs(1804) <= '0';
    layer0_outputs(1805) <= not((inputs(64)) or (inputs(20)));
    layer0_outputs(1806) <= not(inputs(57)) or (inputs(230));
    layer0_outputs(1807) <= inputs(190);
    layer0_outputs(1808) <= not(inputs(37)) or (inputs(124));
    layer0_outputs(1809) <= (inputs(46)) or (inputs(179));
    layer0_outputs(1810) <= not((inputs(6)) or (inputs(135)));
    layer0_outputs(1811) <= (inputs(26)) or (inputs(182));
    layer0_outputs(1812) <= inputs(27);
    layer0_outputs(1813) <= (inputs(244)) and not (inputs(132));
    layer0_outputs(1814) <= (inputs(86)) and not (inputs(190));
    layer0_outputs(1815) <= not((inputs(221)) or (inputs(89)));
    layer0_outputs(1816) <= '0';
    layer0_outputs(1817) <= (inputs(62)) and not (inputs(11));
    layer0_outputs(1818) <= not((inputs(230)) xor (inputs(71)));
    layer0_outputs(1819) <= not((inputs(243)) and (inputs(163)));
    layer0_outputs(1820) <= not(inputs(218)) or (inputs(213));
    layer0_outputs(1821) <= not(inputs(88)) or (inputs(70));
    layer0_outputs(1822) <= not((inputs(120)) xor (inputs(37)));
    layer0_outputs(1823) <= not((inputs(176)) or (inputs(180)));
    layer0_outputs(1824) <= (inputs(128)) and (inputs(192));
    layer0_outputs(1825) <= (inputs(36)) xor (inputs(56));
    layer0_outputs(1826) <= not((inputs(36)) xor (inputs(82)));
    layer0_outputs(1827) <= '1';
    layer0_outputs(1828) <= inputs(56);
    layer0_outputs(1829) <= not((inputs(93)) or (inputs(21)));
    layer0_outputs(1830) <= not(inputs(116)) or (inputs(253));
    layer0_outputs(1831) <= (inputs(44)) and not (inputs(24));
    layer0_outputs(1832) <= inputs(133);
    layer0_outputs(1833) <= not(inputs(221)) or (inputs(190));
    layer0_outputs(1834) <= (inputs(146)) or (inputs(19));
    layer0_outputs(1835) <= not(inputs(180));
    layer0_outputs(1836) <= not((inputs(22)) and (inputs(38)));
    layer0_outputs(1837) <= inputs(196);
    layer0_outputs(1838) <= inputs(151);
    layer0_outputs(1839) <= (inputs(240)) or (inputs(95));
    layer0_outputs(1840) <= (inputs(195)) and not (inputs(40));
    layer0_outputs(1841) <= (inputs(205)) and not (inputs(204));
    layer0_outputs(1842) <= '0';
    layer0_outputs(1843) <= not(inputs(156)) or (inputs(208));
    layer0_outputs(1844) <= not((inputs(235)) xor (inputs(49)));
    layer0_outputs(1845) <= not(inputs(13));
    layer0_outputs(1846) <= not(inputs(119)) or (inputs(207));
    layer0_outputs(1847) <= not((inputs(52)) xor (inputs(150)));
    layer0_outputs(1848) <= inputs(234);
    layer0_outputs(1849) <= (inputs(50)) and (inputs(127));
    layer0_outputs(1850) <= not((inputs(77)) xor (inputs(254)));
    layer0_outputs(1851) <= (inputs(140)) and not (inputs(171));
    layer0_outputs(1852) <= (inputs(217)) and (inputs(114));
    layer0_outputs(1853) <= (inputs(144)) or (inputs(149));
    layer0_outputs(1854) <= (inputs(75)) or (inputs(61));
    layer0_outputs(1855) <= '1';
    layer0_outputs(1856) <= '0';
    layer0_outputs(1857) <= not(inputs(7));
    layer0_outputs(1858) <= not(inputs(18)) or (inputs(70));
    layer0_outputs(1859) <= '1';
    layer0_outputs(1860) <= (inputs(36)) and not (inputs(62));
    layer0_outputs(1861) <= '1';
    layer0_outputs(1862) <= inputs(253);
    layer0_outputs(1863) <= (inputs(128)) or (inputs(128));
    layer0_outputs(1864) <= not(inputs(87));
    layer0_outputs(1865) <= inputs(212);
    layer0_outputs(1866) <= '1';
    layer0_outputs(1867) <= not((inputs(79)) and (inputs(47)));
    layer0_outputs(1868) <= (inputs(98)) and not (inputs(36));
    layer0_outputs(1869) <= (inputs(80)) and not (inputs(75));
    layer0_outputs(1870) <= inputs(213);
    layer0_outputs(1871) <= not((inputs(62)) and (inputs(186)));
    layer0_outputs(1872) <= (inputs(145)) xor (inputs(112));
    layer0_outputs(1873) <= not(inputs(181)) or (inputs(128));
    layer0_outputs(1874) <= not((inputs(210)) xor (inputs(140)));
    layer0_outputs(1875) <= (inputs(155)) and not (inputs(65));
    layer0_outputs(1876) <= (inputs(202)) and (inputs(40));
    layer0_outputs(1877) <= '1';
    layer0_outputs(1878) <= (inputs(61)) and (inputs(46));
    layer0_outputs(1879) <= (inputs(181)) or (inputs(191));
    layer0_outputs(1880) <= (inputs(0)) xor (inputs(202));
    layer0_outputs(1881) <= inputs(122);
    layer0_outputs(1882) <= '1';
    layer0_outputs(1883) <= '1';
    layer0_outputs(1884) <= not((inputs(134)) or (inputs(129)));
    layer0_outputs(1885) <= not(inputs(25));
    layer0_outputs(1886) <= (inputs(42)) and (inputs(39));
    layer0_outputs(1887) <= not((inputs(69)) and (inputs(59)));
    layer0_outputs(1888) <= (inputs(212)) xor (inputs(253));
    layer0_outputs(1889) <= inputs(255);
    layer0_outputs(1890) <= not((inputs(172)) or (inputs(239)));
    layer0_outputs(1891) <= inputs(240);
    layer0_outputs(1892) <= (inputs(15)) and not (inputs(9));
    layer0_outputs(1893) <= (inputs(146)) and not (inputs(2));
    layer0_outputs(1894) <= (inputs(58)) and not (inputs(250));
    layer0_outputs(1895) <= (inputs(37)) and (inputs(108));
    layer0_outputs(1896) <= (inputs(71)) or (inputs(32));
    layer0_outputs(1897) <= not((inputs(233)) or (inputs(96)));
    layer0_outputs(1898) <= (inputs(209)) xor (inputs(249));
    layer0_outputs(1899) <= inputs(166);
    layer0_outputs(1900) <= not(inputs(52));
    layer0_outputs(1901) <= (inputs(123)) and (inputs(211));
    layer0_outputs(1902) <= not(inputs(218)) or (inputs(29));
    layer0_outputs(1903) <= (inputs(17)) and not (inputs(237));
    layer0_outputs(1904) <= '0';
    layer0_outputs(1905) <= not((inputs(183)) or (inputs(122)));
    layer0_outputs(1906) <= inputs(244);
    layer0_outputs(1907) <= '0';
    layer0_outputs(1908) <= not(inputs(222)) or (inputs(216));
    layer0_outputs(1909) <= inputs(87);
    layer0_outputs(1910) <= not((inputs(108)) or (inputs(135)));
    layer0_outputs(1911) <= (inputs(145)) and not (inputs(110));
    layer0_outputs(1912) <= not(inputs(17));
    layer0_outputs(1913) <= (inputs(53)) and not (inputs(10));
    layer0_outputs(1914) <= not(inputs(230));
    layer0_outputs(1915) <= not((inputs(206)) and (inputs(37)));
    layer0_outputs(1916) <= not(inputs(80)) or (inputs(46));
    layer0_outputs(1917) <= '0';
    layer0_outputs(1918) <= inputs(119);
    layer0_outputs(1919) <= not(inputs(215)) or (inputs(7));
    layer0_outputs(1920) <= (inputs(12)) and not (inputs(217));
    layer0_outputs(1921) <= not(inputs(72));
    layer0_outputs(1922) <= not(inputs(212)) or (inputs(234));
    layer0_outputs(1923) <= (inputs(44)) and not (inputs(46));
    layer0_outputs(1924) <= not(inputs(201)) or (inputs(46));
    layer0_outputs(1925) <= not((inputs(102)) or (inputs(133)));
    layer0_outputs(1926) <= not(inputs(89)) or (inputs(132));
    layer0_outputs(1927) <= (inputs(21)) or (inputs(149));
    layer0_outputs(1928) <= not((inputs(149)) xor (inputs(224)));
    layer0_outputs(1929) <= not((inputs(69)) xor (inputs(161)));
    layer0_outputs(1930) <= (inputs(179)) and not (inputs(47));
    layer0_outputs(1931) <= not(inputs(112)) or (inputs(214));
    layer0_outputs(1932) <= not(inputs(176));
    layer0_outputs(1933) <= inputs(106);
    layer0_outputs(1934) <= (inputs(115)) xor (inputs(226));
    layer0_outputs(1935) <= inputs(5);
    layer0_outputs(1936) <= not(inputs(34));
    layer0_outputs(1937) <= not((inputs(46)) xor (inputs(213)));
    layer0_outputs(1938) <= (inputs(159)) or (inputs(197));
    layer0_outputs(1939) <= inputs(51);
    layer0_outputs(1940) <= (inputs(221)) and (inputs(26));
    layer0_outputs(1941) <= (inputs(132)) and not (inputs(200));
    layer0_outputs(1942) <= '0';
    layer0_outputs(1943) <= not((inputs(93)) or (inputs(72)));
    layer0_outputs(1944) <= (inputs(121)) or (inputs(107));
    layer0_outputs(1945) <= not(inputs(119));
    layer0_outputs(1946) <= not((inputs(189)) and (inputs(65)));
    layer0_outputs(1947) <= inputs(160);
    layer0_outputs(1948) <= '1';
    layer0_outputs(1949) <= (inputs(99)) xor (inputs(74));
    layer0_outputs(1950) <= inputs(140);
    layer0_outputs(1951) <= (inputs(64)) and (inputs(46));
    layer0_outputs(1952) <= '1';
    layer0_outputs(1953) <= not((inputs(73)) xor (inputs(112)));
    layer0_outputs(1954) <= (inputs(59)) or (inputs(173));
    layer0_outputs(1955) <= not((inputs(108)) or (inputs(64)));
    layer0_outputs(1956) <= inputs(190);
    layer0_outputs(1957) <= (inputs(106)) and not (inputs(127));
    layer0_outputs(1958) <= (inputs(6)) or (inputs(151));
    layer0_outputs(1959) <= (inputs(6)) xor (inputs(152));
    layer0_outputs(1960) <= not(inputs(35));
    layer0_outputs(1961) <= '0';
    layer0_outputs(1962) <= not(inputs(240)) or (inputs(99));
    layer0_outputs(1963) <= (inputs(117)) xor (inputs(242));
    layer0_outputs(1964) <= not((inputs(204)) xor (inputs(2)));
    layer0_outputs(1965) <= (inputs(130)) or (inputs(200));
    layer0_outputs(1966) <= (inputs(214)) or (inputs(74));
    layer0_outputs(1967) <= not(inputs(181));
    layer0_outputs(1968) <= inputs(136);
    layer0_outputs(1969) <= (inputs(248)) and not (inputs(45));
    layer0_outputs(1970) <= (inputs(156)) or (inputs(242));
    layer0_outputs(1971) <= (inputs(231)) or (inputs(116));
    layer0_outputs(1972) <= inputs(165);
    layer0_outputs(1973) <= '0';
    layer0_outputs(1974) <= inputs(2);
    layer0_outputs(1975) <= (inputs(31)) and not (inputs(219));
    layer0_outputs(1976) <= not(inputs(245)) or (inputs(181));
    layer0_outputs(1977) <= not((inputs(31)) and (inputs(122)));
    layer0_outputs(1978) <= not((inputs(181)) xor (inputs(60)));
    layer0_outputs(1979) <= inputs(196);
    layer0_outputs(1980) <= not(inputs(117));
    layer0_outputs(1981) <= not((inputs(231)) or (inputs(18)));
    layer0_outputs(1982) <= (inputs(179)) and not (inputs(17));
    layer0_outputs(1983) <= (inputs(155)) or (inputs(179));
    layer0_outputs(1984) <= (inputs(105)) and not (inputs(84));
    layer0_outputs(1985) <= inputs(164);
    layer0_outputs(1986) <= (inputs(28)) or (inputs(163));
    layer0_outputs(1987) <= not(inputs(142));
    layer0_outputs(1988) <= inputs(250);
    layer0_outputs(1989) <= not(inputs(102)) or (inputs(102));
    layer0_outputs(1990) <= (inputs(120)) and not (inputs(1));
    layer0_outputs(1991) <= not(inputs(56)) or (inputs(184));
    layer0_outputs(1992) <= inputs(113);
    layer0_outputs(1993) <= (inputs(230)) or (inputs(76));
    layer0_outputs(1994) <= (inputs(211)) and not (inputs(228));
    layer0_outputs(1995) <= not((inputs(109)) xor (inputs(26)));
    layer0_outputs(1996) <= not(inputs(28));
    layer0_outputs(1997) <= (inputs(243)) or (inputs(137));
    layer0_outputs(1998) <= not(inputs(107));
    layer0_outputs(1999) <= '0';
    layer0_outputs(2000) <= (inputs(109)) or (inputs(124));
    layer0_outputs(2001) <= not(inputs(96)) or (inputs(86));
    layer0_outputs(2002) <= not((inputs(28)) xor (inputs(192)));
    layer0_outputs(2003) <= inputs(32);
    layer0_outputs(2004) <= not(inputs(165));
    layer0_outputs(2005) <= inputs(175);
    layer0_outputs(2006) <= not(inputs(61)) or (inputs(9));
    layer0_outputs(2007) <= not((inputs(156)) or (inputs(208)));
    layer0_outputs(2008) <= '1';
    layer0_outputs(2009) <= not((inputs(131)) xor (inputs(239)));
    layer0_outputs(2010) <= not(inputs(189));
    layer0_outputs(2011) <= inputs(146);
    layer0_outputs(2012) <= not((inputs(125)) and (inputs(3)));
    layer0_outputs(2013) <= (inputs(216)) or (inputs(14));
    layer0_outputs(2014) <= not(inputs(34)) or (inputs(189));
    layer0_outputs(2015) <= (inputs(137)) xor (inputs(193));
    layer0_outputs(2016) <= inputs(132);
    layer0_outputs(2017) <= (inputs(145)) and (inputs(253));
    layer0_outputs(2018) <= not(inputs(36));
    layer0_outputs(2019) <= not((inputs(10)) and (inputs(13)));
    layer0_outputs(2020) <= not((inputs(223)) or (inputs(191)));
    layer0_outputs(2021) <= not(inputs(231)) or (inputs(36));
    layer0_outputs(2022) <= not((inputs(158)) or (inputs(201)));
    layer0_outputs(2023) <= (inputs(91)) or (inputs(132));
    layer0_outputs(2024) <= not((inputs(171)) xor (inputs(91)));
    layer0_outputs(2025) <= (inputs(63)) or (inputs(23));
    layer0_outputs(2026) <= (inputs(64)) and not (inputs(48));
    layer0_outputs(2027) <= '0';
    layer0_outputs(2028) <= not((inputs(129)) xor (inputs(67)));
    layer0_outputs(2029) <= inputs(117);
    layer0_outputs(2030) <= not((inputs(51)) xor (inputs(99)));
    layer0_outputs(2031) <= not((inputs(169)) xor (inputs(113)));
    layer0_outputs(2032) <= '1';
    layer0_outputs(2033) <= (inputs(185)) and (inputs(105));
    layer0_outputs(2034) <= not((inputs(73)) or (inputs(15)));
    layer0_outputs(2035) <= not(inputs(86));
    layer0_outputs(2036) <= not((inputs(38)) or (inputs(3)));
    layer0_outputs(2037) <= inputs(73);
    layer0_outputs(2038) <= inputs(154);
    layer0_outputs(2039) <= (inputs(188)) or (inputs(166));
    layer0_outputs(2040) <= (inputs(17)) and not (inputs(164));
    layer0_outputs(2041) <= not((inputs(75)) xor (inputs(150)));
    layer0_outputs(2042) <= inputs(14);
    layer0_outputs(2043) <= '1';
    layer0_outputs(2044) <= not((inputs(163)) or (inputs(7)));
    layer0_outputs(2045) <= (inputs(246)) and not (inputs(163));
    layer0_outputs(2046) <= not(inputs(236));
    layer0_outputs(2047) <= (inputs(26)) or (inputs(106));
    layer0_outputs(2048) <= not((inputs(78)) or (inputs(143)));
    layer0_outputs(2049) <= (inputs(35)) and not (inputs(206));
    layer0_outputs(2050) <= (inputs(144)) and (inputs(241));
    layer0_outputs(2051) <= (inputs(147)) xor (inputs(149));
    layer0_outputs(2052) <= not(inputs(194)) or (inputs(87));
    layer0_outputs(2053) <= (inputs(255)) xor (inputs(59));
    layer0_outputs(2054) <= '0';
    layer0_outputs(2055) <= inputs(103);
    layer0_outputs(2056) <= not(inputs(203)) or (inputs(42));
    layer0_outputs(2057) <= not((inputs(18)) and (inputs(139)));
    layer0_outputs(2058) <= not((inputs(32)) and (inputs(52)));
    layer0_outputs(2059) <= inputs(44);
    layer0_outputs(2060) <= inputs(103);
    layer0_outputs(2061) <= not(inputs(254)) or (inputs(103));
    layer0_outputs(2062) <= (inputs(200)) xor (inputs(246));
    layer0_outputs(2063) <= inputs(56);
    layer0_outputs(2064) <= not(inputs(238)) or (inputs(123));
    layer0_outputs(2065) <= (inputs(99)) and not (inputs(225));
    layer0_outputs(2066) <= not(inputs(220)) or (inputs(150));
    layer0_outputs(2067) <= '0';
    layer0_outputs(2068) <= inputs(180);
    layer0_outputs(2069) <= inputs(14);
    layer0_outputs(2070) <= inputs(167);
    layer0_outputs(2071) <= not(inputs(87));
    layer0_outputs(2072) <= inputs(179);
    layer0_outputs(2073) <= not((inputs(141)) and (inputs(165)));
    layer0_outputs(2074) <= (inputs(57)) xor (inputs(48));
    layer0_outputs(2075) <= (inputs(90)) and not (inputs(147));
    layer0_outputs(2076) <= (inputs(76)) or (inputs(173));
    layer0_outputs(2077) <= not((inputs(48)) or (inputs(210)));
    layer0_outputs(2078) <= not(inputs(255));
    layer0_outputs(2079) <= inputs(182);
    layer0_outputs(2080) <= inputs(224);
    layer0_outputs(2081) <= inputs(196);
    layer0_outputs(2082) <= (inputs(180)) and not (inputs(79));
    layer0_outputs(2083) <= inputs(163);
    layer0_outputs(2084) <= inputs(16);
    layer0_outputs(2085) <= not((inputs(97)) and (inputs(15)));
    layer0_outputs(2086) <= (inputs(250)) and not (inputs(243));
    layer0_outputs(2087) <= inputs(78);
    layer0_outputs(2088) <= (inputs(170)) or (inputs(186));
    layer0_outputs(2089) <= not((inputs(125)) or (inputs(173)));
    layer0_outputs(2090) <= not(inputs(189)) or (inputs(245));
    layer0_outputs(2091) <= not(inputs(165)) or (inputs(60));
    layer0_outputs(2092) <= inputs(42);
    layer0_outputs(2093) <= not(inputs(101)) or (inputs(50));
    layer0_outputs(2094) <= not(inputs(249));
    layer0_outputs(2095) <= not((inputs(75)) and (inputs(7)));
    layer0_outputs(2096) <= not((inputs(248)) or (inputs(130)));
    layer0_outputs(2097) <= inputs(255);
    layer0_outputs(2098) <= '1';
    layer0_outputs(2099) <= not(inputs(31)) or (inputs(51));
    layer0_outputs(2100) <= not((inputs(39)) and (inputs(142)));
    layer0_outputs(2101) <= (inputs(203)) or (inputs(83));
    layer0_outputs(2102) <= (inputs(164)) and (inputs(208));
    layer0_outputs(2103) <= not(inputs(54));
    layer0_outputs(2104) <= (inputs(33)) xor (inputs(163));
    layer0_outputs(2105) <= not(inputs(32)) or (inputs(246));
    layer0_outputs(2106) <= (inputs(193)) and not (inputs(43));
    layer0_outputs(2107) <= (inputs(86)) or (inputs(28));
    layer0_outputs(2108) <= (inputs(181)) and not (inputs(249));
    layer0_outputs(2109) <= not((inputs(249)) and (inputs(242)));
    layer0_outputs(2110) <= '0';
    layer0_outputs(2111) <= inputs(72);
    layer0_outputs(2112) <= not(inputs(141)) or (inputs(239));
    layer0_outputs(2113) <= (inputs(126)) and not (inputs(216));
    layer0_outputs(2114) <= inputs(29);
    layer0_outputs(2115) <= '1';
    layer0_outputs(2116) <= '1';
    layer0_outputs(2117) <= (inputs(67)) or (inputs(53));
    layer0_outputs(2118) <= not(inputs(33));
    layer0_outputs(2119) <= not((inputs(196)) xor (inputs(39)));
    layer0_outputs(2120) <= (inputs(59)) xor (inputs(146));
    layer0_outputs(2121) <= (inputs(206)) and not (inputs(23));
    layer0_outputs(2122) <= '0';
    layer0_outputs(2123) <= inputs(92);
    layer0_outputs(2124) <= not(inputs(174)) or (inputs(85));
    layer0_outputs(2125) <= not(inputs(224));
    layer0_outputs(2126) <= inputs(151);
    layer0_outputs(2127) <= (inputs(51)) and not (inputs(41));
    layer0_outputs(2128) <= '1';
    layer0_outputs(2129) <= (inputs(242)) or (inputs(83));
    layer0_outputs(2130) <= '0';
    layer0_outputs(2131) <= not(inputs(247));
    layer0_outputs(2132) <= not((inputs(228)) or (inputs(183)));
    layer0_outputs(2133) <= not(inputs(62));
    layer0_outputs(2134) <= inputs(168);
    layer0_outputs(2135) <= not(inputs(24));
    layer0_outputs(2136) <= (inputs(74)) or (inputs(246));
    layer0_outputs(2137) <= (inputs(103)) and not (inputs(72));
    layer0_outputs(2138) <= (inputs(53)) and (inputs(53));
    layer0_outputs(2139) <= not((inputs(16)) or (inputs(42)));
    layer0_outputs(2140) <= (inputs(165)) and not (inputs(31));
    layer0_outputs(2141) <= not((inputs(22)) and (inputs(95)));
    layer0_outputs(2142) <= '1';
    layer0_outputs(2143) <= (inputs(77)) or (inputs(13));
    layer0_outputs(2144) <= not(inputs(112)) or (inputs(144));
    layer0_outputs(2145) <= inputs(139);
    layer0_outputs(2146) <= inputs(163);
    layer0_outputs(2147) <= not((inputs(71)) xor (inputs(214)));
    layer0_outputs(2148) <= (inputs(101)) and not (inputs(179));
    layer0_outputs(2149) <= '0';
    layer0_outputs(2150) <= not(inputs(196));
    layer0_outputs(2151) <= inputs(71);
    layer0_outputs(2152) <= (inputs(215)) and not (inputs(41));
    layer0_outputs(2153) <= (inputs(186)) and not (inputs(86));
    layer0_outputs(2154) <= (inputs(158)) and not (inputs(206));
    layer0_outputs(2155) <= inputs(162);
    layer0_outputs(2156) <= inputs(227);
    layer0_outputs(2157) <= not(inputs(87));
    layer0_outputs(2158) <= not((inputs(188)) xor (inputs(87)));
    layer0_outputs(2159) <= (inputs(68)) and not (inputs(148));
    layer0_outputs(2160) <= (inputs(235)) xor (inputs(51));
    layer0_outputs(2161) <= (inputs(174)) and not (inputs(234));
    layer0_outputs(2162) <= not((inputs(67)) or (inputs(47)));
    layer0_outputs(2163) <= not(inputs(158)) or (inputs(114));
    layer0_outputs(2164) <= inputs(249);
    layer0_outputs(2165) <= (inputs(105)) and not (inputs(99));
    layer0_outputs(2166) <= not(inputs(149));
    layer0_outputs(2167) <= (inputs(59)) and (inputs(39));
    layer0_outputs(2168) <= inputs(111);
    layer0_outputs(2169) <= inputs(219);
    layer0_outputs(2170) <= not(inputs(119)) or (inputs(230));
    layer0_outputs(2171) <= not((inputs(216)) xor (inputs(58)));
    layer0_outputs(2172) <= (inputs(124)) and (inputs(111));
    layer0_outputs(2173) <= not((inputs(248)) and (inputs(168)));
    layer0_outputs(2174) <= (inputs(192)) and (inputs(6));
    layer0_outputs(2175) <= '1';
    layer0_outputs(2176) <= (inputs(94)) and not (inputs(94));
    layer0_outputs(2177) <= (inputs(211)) and not (inputs(132));
    layer0_outputs(2178) <= (inputs(199)) and not (inputs(194));
    layer0_outputs(2179) <= inputs(18);
    layer0_outputs(2180) <= (inputs(208)) and not (inputs(227));
    layer0_outputs(2181) <= not(inputs(80)) or (inputs(50));
    layer0_outputs(2182) <= inputs(229);
    layer0_outputs(2183) <= not((inputs(216)) or (inputs(128)));
    layer0_outputs(2184) <= (inputs(83)) and not (inputs(129));
    layer0_outputs(2185) <= (inputs(138)) and not (inputs(191));
    layer0_outputs(2186) <= inputs(165);
    layer0_outputs(2187) <= (inputs(177)) and not (inputs(64));
    layer0_outputs(2188) <= not(inputs(83));
    layer0_outputs(2189) <= (inputs(106)) or (inputs(49));
    layer0_outputs(2190) <= not(inputs(140)) or (inputs(123));
    layer0_outputs(2191) <= inputs(52);
    layer0_outputs(2192) <= (inputs(171)) or (inputs(22));
    layer0_outputs(2193) <= not(inputs(203));
    layer0_outputs(2194) <= not((inputs(242)) and (inputs(165)));
    layer0_outputs(2195) <= (inputs(134)) or (inputs(59));
    layer0_outputs(2196) <= '0';
    layer0_outputs(2197) <= not(inputs(172));
    layer0_outputs(2198) <= (inputs(14)) xor (inputs(2));
    layer0_outputs(2199) <= not((inputs(56)) or (inputs(194)));
    layer0_outputs(2200) <= not((inputs(176)) and (inputs(121)));
    layer0_outputs(2201) <= inputs(51);
    layer0_outputs(2202) <= (inputs(227)) and not (inputs(156));
    layer0_outputs(2203) <= not(inputs(21)) or (inputs(216));
    layer0_outputs(2204) <= not(inputs(162)) or (inputs(246));
    layer0_outputs(2205) <= not(inputs(9));
    layer0_outputs(2206) <= (inputs(194)) or (inputs(96));
    layer0_outputs(2207) <= '1';
    layer0_outputs(2208) <= not(inputs(214));
    layer0_outputs(2209) <= not(inputs(199)) or (inputs(61));
    layer0_outputs(2210) <= not(inputs(199));
    layer0_outputs(2211) <= '0';
    layer0_outputs(2212) <= (inputs(74)) and not (inputs(36));
    layer0_outputs(2213) <= (inputs(4)) xor (inputs(140));
    layer0_outputs(2214) <= not((inputs(83)) or (inputs(74)));
    layer0_outputs(2215) <= (inputs(222)) and (inputs(248));
    layer0_outputs(2216) <= not((inputs(156)) or (inputs(170)));
    layer0_outputs(2217) <= not(inputs(69));
    layer0_outputs(2218) <= inputs(166);
    layer0_outputs(2219) <= (inputs(52)) and not (inputs(10));
    layer0_outputs(2220) <= (inputs(246)) xor (inputs(194));
    layer0_outputs(2221) <= (inputs(163)) and not (inputs(161));
    layer0_outputs(2222) <= not(inputs(165));
    layer0_outputs(2223) <= not(inputs(138)) or (inputs(47));
    layer0_outputs(2224) <= (inputs(100)) and not (inputs(113));
    layer0_outputs(2225) <= (inputs(209)) or (inputs(27));
    layer0_outputs(2226) <= '0';
    layer0_outputs(2227) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(2228) <= (inputs(216)) xor (inputs(18));
    layer0_outputs(2229) <= not(inputs(92)) or (inputs(210));
    layer0_outputs(2230) <= not((inputs(87)) and (inputs(207)));
    layer0_outputs(2231) <= not(inputs(247)) or (inputs(161));
    layer0_outputs(2232) <= not((inputs(160)) or (inputs(33)));
    layer0_outputs(2233) <= (inputs(27)) and not (inputs(130));
    layer0_outputs(2234) <= inputs(16);
    layer0_outputs(2235) <= (inputs(233)) and not (inputs(206));
    layer0_outputs(2236) <= not(inputs(215));
    layer0_outputs(2237) <= (inputs(244)) and (inputs(219));
    layer0_outputs(2238) <= not(inputs(21));
    layer0_outputs(2239) <= (inputs(182)) and not (inputs(17));
    layer0_outputs(2240) <= (inputs(66)) or (inputs(244));
    layer0_outputs(2241) <= not(inputs(116));
    layer0_outputs(2242) <= not((inputs(122)) or (inputs(98)));
    layer0_outputs(2243) <= not(inputs(241));
    layer0_outputs(2244) <= '1';
    layer0_outputs(2245) <= inputs(186);
    layer0_outputs(2246) <= not(inputs(88));
    layer0_outputs(2247) <= (inputs(239)) and (inputs(177));
    layer0_outputs(2248) <= not(inputs(147));
    layer0_outputs(2249) <= (inputs(66)) and not (inputs(169));
    layer0_outputs(2250) <= inputs(26);
    layer0_outputs(2251) <= '1';
    layer0_outputs(2252) <= (inputs(153)) or (inputs(171));
    layer0_outputs(2253) <= not(inputs(111));
    layer0_outputs(2254) <= '1';
    layer0_outputs(2255) <= (inputs(41)) and not (inputs(85));
    layer0_outputs(2256) <= (inputs(172)) xor (inputs(4));
    layer0_outputs(2257) <= (inputs(153)) and not (inputs(41));
    layer0_outputs(2258) <= (inputs(166)) and not (inputs(213));
    layer0_outputs(2259) <= not(inputs(254)) or (inputs(31));
    layer0_outputs(2260) <= (inputs(64)) or (inputs(112));
    layer0_outputs(2261) <= '0';
    layer0_outputs(2262) <= not(inputs(153));
    layer0_outputs(2263) <= not((inputs(6)) and (inputs(204)));
    layer0_outputs(2264) <= (inputs(222)) or (inputs(86));
    layer0_outputs(2265) <= (inputs(58)) and not (inputs(226));
    layer0_outputs(2266) <= not(inputs(72)) or (inputs(93));
    layer0_outputs(2267) <= not(inputs(82)) or (inputs(115));
    layer0_outputs(2268) <= not(inputs(202));
    layer0_outputs(2269) <= (inputs(160)) and not (inputs(96));
    layer0_outputs(2270) <= '0';
    layer0_outputs(2271) <= not((inputs(224)) or (inputs(180)));
    layer0_outputs(2272) <= not(inputs(3));
    layer0_outputs(2273) <= not(inputs(80)) or (inputs(98));
    layer0_outputs(2274) <= (inputs(49)) and not (inputs(104));
    layer0_outputs(2275) <= (inputs(249)) and not (inputs(32));
    layer0_outputs(2276) <= (inputs(104)) and not (inputs(144));
    layer0_outputs(2277) <= not(inputs(170));
    layer0_outputs(2278) <= not((inputs(159)) or (inputs(99)));
    layer0_outputs(2279) <= not(inputs(96));
    layer0_outputs(2280) <= not((inputs(192)) xor (inputs(104)));
    layer0_outputs(2281) <= not(inputs(136));
    layer0_outputs(2282) <= (inputs(241)) and not (inputs(199));
    layer0_outputs(2283) <= not(inputs(95));
    layer0_outputs(2284) <= (inputs(110)) xor (inputs(78));
    layer0_outputs(2285) <= not((inputs(170)) and (inputs(52)));
    layer0_outputs(2286) <= not(inputs(244));
    layer0_outputs(2287) <= inputs(166);
    layer0_outputs(2288) <= not(inputs(17)) or (inputs(125));
    layer0_outputs(2289) <= not(inputs(58)) or (inputs(142));
    layer0_outputs(2290) <= inputs(241);
    layer0_outputs(2291) <= inputs(153);
    layer0_outputs(2292) <= not(inputs(97));
    layer0_outputs(2293) <= not((inputs(37)) and (inputs(13)));
    layer0_outputs(2294) <= not(inputs(173)) or (inputs(82));
    layer0_outputs(2295) <= (inputs(97)) and (inputs(11));
    layer0_outputs(2296) <= not(inputs(116));
    layer0_outputs(2297) <= not(inputs(240));
    layer0_outputs(2298) <= not(inputs(141)) or (inputs(143));
    layer0_outputs(2299) <= not(inputs(137)) or (inputs(84));
    layer0_outputs(2300) <= inputs(69);
    layer0_outputs(2301) <= not((inputs(156)) or (inputs(195)));
    layer0_outputs(2302) <= (inputs(151)) or (inputs(82));
    layer0_outputs(2303) <= not(inputs(191));
    layer0_outputs(2304) <= not((inputs(71)) or (inputs(255)));
    layer0_outputs(2305) <= not((inputs(14)) or (inputs(99)));
    layer0_outputs(2306) <= not(inputs(58)) or (inputs(193));
    layer0_outputs(2307) <= (inputs(150)) xor (inputs(109));
    layer0_outputs(2308) <= not(inputs(168));
    layer0_outputs(2309) <= not(inputs(80)) or (inputs(244));
    layer0_outputs(2310) <= (inputs(152)) and not (inputs(38));
    layer0_outputs(2311) <= not((inputs(71)) and (inputs(187)));
    layer0_outputs(2312) <= not(inputs(70));
    layer0_outputs(2313) <= not(inputs(16)) or (inputs(65));
    layer0_outputs(2314) <= not((inputs(227)) xor (inputs(129)));
    layer0_outputs(2315) <= not((inputs(160)) and (inputs(195)));
    layer0_outputs(2316) <= not(inputs(57)) or (inputs(99));
    layer0_outputs(2317) <= inputs(86);
    layer0_outputs(2318) <= (inputs(187)) or (inputs(233));
    layer0_outputs(2319) <= (inputs(192)) or (inputs(73));
    layer0_outputs(2320) <= inputs(180);
    layer0_outputs(2321) <= inputs(180);
    layer0_outputs(2322) <= not(inputs(216)) or (inputs(86));
    layer0_outputs(2323) <= (inputs(100)) and not (inputs(155));
    layer0_outputs(2324) <= '0';
    layer0_outputs(2325) <= (inputs(23)) and not (inputs(130));
    layer0_outputs(2326) <= (inputs(16)) or (inputs(121));
    layer0_outputs(2327) <= (inputs(4)) xor (inputs(229));
    layer0_outputs(2328) <= not(inputs(123));
    layer0_outputs(2329) <= '0';
    layer0_outputs(2330) <= (inputs(231)) and not (inputs(110));
    layer0_outputs(2331) <= (inputs(44)) and (inputs(43));
    layer0_outputs(2332) <= (inputs(231)) or (inputs(106));
    layer0_outputs(2333) <= inputs(207);
    layer0_outputs(2334) <= (inputs(133)) and not (inputs(104));
    layer0_outputs(2335) <= not(inputs(215)) or (inputs(157));
    layer0_outputs(2336) <= (inputs(169)) and not (inputs(184));
    layer0_outputs(2337) <= '0';
    layer0_outputs(2338) <= not((inputs(67)) or (inputs(29)));
    layer0_outputs(2339) <= (inputs(171)) and not (inputs(4));
    layer0_outputs(2340) <= (inputs(119)) and not (inputs(23));
    layer0_outputs(2341) <= not(inputs(91));
    layer0_outputs(2342) <= (inputs(243)) xor (inputs(245));
    layer0_outputs(2343) <= inputs(180);
    layer0_outputs(2344) <= inputs(155);
    layer0_outputs(2345) <= (inputs(156)) and not (inputs(177));
    layer0_outputs(2346) <= (inputs(118)) and not (inputs(82));
    layer0_outputs(2347) <= not(inputs(2)) or (inputs(90));
    layer0_outputs(2348) <= not(inputs(80)) or (inputs(40));
    layer0_outputs(2349) <= inputs(139);
    layer0_outputs(2350) <= not((inputs(118)) or (inputs(111)));
    layer0_outputs(2351) <= not((inputs(137)) xor (inputs(36)));
    layer0_outputs(2352) <= (inputs(19)) xor (inputs(4));
    layer0_outputs(2353) <= not((inputs(66)) xor (inputs(247)));
    layer0_outputs(2354) <= not((inputs(19)) and (inputs(172)));
    layer0_outputs(2355) <= not(inputs(188)) or (inputs(253));
    layer0_outputs(2356) <= '1';
    layer0_outputs(2357) <= not(inputs(109));
    layer0_outputs(2358) <= not(inputs(151)) or (inputs(106));
    layer0_outputs(2359) <= not(inputs(122));
    layer0_outputs(2360) <= (inputs(196)) and not (inputs(253));
    layer0_outputs(2361) <= not((inputs(233)) or (inputs(52)));
    layer0_outputs(2362) <= (inputs(97)) xor (inputs(10));
    layer0_outputs(2363) <= not((inputs(76)) xor (inputs(242)));
    layer0_outputs(2364) <= not(inputs(146));
    layer0_outputs(2365) <= inputs(101);
    layer0_outputs(2366) <= not((inputs(66)) or (inputs(82)));
    layer0_outputs(2367) <= not(inputs(55));
    layer0_outputs(2368) <= not(inputs(191));
    layer0_outputs(2369) <= (inputs(54)) and not (inputs(109));
    layer0_outputs(2370) <= not(inputs(90));
    layer0_outputs(2371) <= not((inputs(90)) or (inputs(234)));
    layer0_outputs(2372) <= not((inputs(69)) or (inputs(74)));
    layer0_outputs(2373) <= (inputs(45)) and not (inputs(47));
    layer0_outputs(2374) <= not((inputs(193)) or (inputs(146)));
    layer0_outputs(2375) <= '1';
    layer0_outputs(2376) <= inputs(251);
    layer0_outputs(2377) <= (inputs(204)) or (inputs(52));
    layer0_outputs(2378) <= inputs(233);
    layer0_outputs(2379) <= not(inputs(117)) or (inputs(69));
    layer0_outputs(2380) <= (inputs(119)) and not (inputs(11));
    layer0_outputs(2381) <= not(inputs(152));
    layer0_outputs(2382) <= '1';
    layer0_outputs(2383) <= '0';
    layer0_outputs(2384) <= (inputs(2)) and not (inputs(247));
    layer0_outputs(2385) <= not((inputs(239)) xor (inputs(100)));
    layer0_outputs(2386) <= not((inputs(176)) or (inputs(27)));
    layer0_outputs(2387) <= (inputs(38)) and not (inputs(143));
    layer0_outputs(2388) <= (inputs(162)) or (inputs(57));
    layer0_outputs(2389) <= not(inputs(167)) or (inputs(232));
    layer0_outputs(2390) <= not((inputs(203)) or (inputs(222)));
    layer0_outputs(2391) <= not(inputs(140)) or (inputs(212));
    layer0_outputs(2392) <= not(inputs(187));
    layer0_outputs(2393) <= not(inputs(52)) or (inputs(111));
    layer0_outputs(2394) <= '1';
    layer0_outputs(2395) <= inputs(100);
    layer0_outputs(2396) <= (inputs(201)) and not (inputs(230));
    layer0_outputs(2397) <= inputs(191);
    layer0_outputs(2398) <= not((inputs(79)) xor (inputs(186)));
    layer0_outputs(2399) <= not(inputs(169));
    layer0_outputs(2400) <= not(inputs(77)) or (inputs(169));
    layer0_outputs(2401) <= not((inputs(101)) or (inputs(143)));
    layer0_outputs(2402) <= (inputs(250)) xor (inputs(217));
    layer0_outputs(2403) <= inputs(30);
    layer0_outputs(2404) <= (inputs(170)) xor (inputs(126));
    layer0_outputs(2405) <= inputs(164);
    layer0_outputs(2406) <= (inputs(220)) or (inputs(53));
    layer0_outputs(2407) <= not(inputs(204)) or (inputs(223));
    layer0_outputs(2408) <= '1';
    layer0_outputs(2409) <= (inputs(77)) xor (inputs(108));
    layer0_outputs(2410) <= '1';
    layer0_outputs(2411) <= inputs(162);
    layer0_outputs(2412) <= not(inputs(67)) or (inputs(231));
    layer0_outputs(2413) <= not((inputs(2)) and (inputs(223)));
    layer0_outputs(2414) <= not(inputs(170)) or (inputs(169));
    layer0_outputs(2415) <= inputs(77);
    layer0_outputs(2416) <= (inputs(135)) and not (inputs(45));
    layer0_outputs(2417) <= inputs(244);
    layer0_outputs(2418) <= (inputs(247)) or (inputs(111));
    layer0_outputs(2419) <= not((inputs(227)) and (inputs(0)));
    layer0_outputs(2420) <= '1';
    layer0_outputs(2421) <= not(inputs(123));
    layer0_outputs(2422) <= (inputs(94)) or (inputs(122));
    layer0_outputs(2423) <= inputs(167);
    layer0_outputs(2424) <= not((inputs(202)) and (inputs(54)));
    layer0_outputs(2425) <= (inputs(200)) and (inputs(190));
    layer0_outputs(2426) <= not(inputs(54));
    layer0_outputs(2427) <= '1';
    layer0_outputs(2428) <= not(inputs(250)) or (inputs(154));
    layer0_outputs(2429) <= (inputs(8)) or (inputs(58));
    layer0_outputs(2430) <= (inputs(88)) or (inputs(174));
    layer0_outputs(2431) <= not(inputs(166)) or (inputs(50));
    layer0_outputs(2432) <= inputs(108);
    layer0_outputs(2433) <= '1';
    layer0_outputs(2434) <= (inputs(74)) and not (inputs(239));
    layer0_outputs(2435) <= inputs(73);
    layer0_outputs(2436) <= '1';
    layer0_outputs(2437) <= '0';
    layer0_outputs(2438) <= not((inputs(13)) xor (inputs(235)));
    layer0_outputs(2439) <= '1';
    layer0_outputs(2440) <= not(inputs(171));
    layer0_outputs(2441) <= not(inputs(200)) or (inputs(217));
    layer0_outputs(2442) <= inputs(81);
    layer0_outputs(2443) <= not((inputs(33)) xor (inputs(184)));
    layer0_outputs(2444) <= not(inputs(216));
    layer0_outputs(2445) <= inputs(21);
    layer0_outputs(2446) <= (inputs(61)) xor (inputs(80));
    layer0_outputs(2447) <= (inputs(224)) and (inputs(224));
    layer0_outputs(2448) <= not((inputs(13)) and (inputs(220)));
    layer0_outputs(2449) <= '0';
    layer0_outputs(2450) <= (inputs(15)) xor (inputs(8));
    layer0_outputs(2451) <= inputs(3);
    layer0_outputs(2452) <= (inputs(141)) or (inputs(153));
    layer0_outputs(2453) <= not((inputs(133)) xor (inputs(204)));
    layer0_outputs(2454) <= not(inputs(17)) or (inputs(217));
    layer0_outputs(2455) <= inputs(221);
    layer0_outputs(2456) <= not(inputs(9)) or (inputs(214));
    layer0_outputs(2457) <= (inputs(84)) xor (inputs(170));
    layer0_outputs(2458) <= not((inputs(200)) and (inputs(11)));
    layer0_outputs(2459) <= not(inputs(219)) or (inputs(12));
    layer0_outputs(2460) <= (inputs(248)) or (inputs(106));
    layer0_outputs(2461) <= (inputs(105)) or (inputs(176));
    layer0_outputs(2462) <= not((inputs(210)) or (inputs(106)));
    layer0_outputs(2463) <= '0';
    layer0_outputs(2464) <= not((inputs(141)) xor (inputs(28)));
    layer0_outputs(2465) <= not((inputs(77)) or (inputs(56)));
    layer0_outputs(2466) <= inputs(168);
    layer0_outputs(2467) <= not(inputs(216));
    layer0_outputs(2468) <= inputs(122);
    layer0_outputs(2469) <= not((inputs(173)) or (inputs(159)));
    layer0_outputs(2470) <= not(inputs(155)) or (inputs(20));
    layer0_outputs(2471) <= not(inputs(179));
    layer0_outputs(2472) <= not(inputs(34));
    layer0_outputs(2473) <= not(inputs(77)) or (inputs(188));
    layer0_outputs(2474) <= not((inputs(78)) or (inputs(114)));
    layer0_outputs(2475) <= not((inputs(86)) and (inputs(228)));
    layer0_outputs(2476) <= not((inputs(95)) xor (inputs(96)));
    layer0_outputs(2477) <= not(inputs(138));
    layer0_outputs(2478) <= '1';
    layer0_outputs(2479) <= not(inputs(29));
    layer0_outputs(2480) <= not(inputs(75));
    layer0_outputs(2481) <= (inputs(171)) and not (inputs(97));
    layer0_outputs(2482) <= (inputs(200)) xor (inputs(31));
    layer0_outputs(2483) <= not((inputs(186)) or (inputs(179)));
    layer0_outputs(2484) <= not(inputs(105));
    layer0_outputs(2485) <= '0';
    layer0_outputs(2486) <= (inputs(81)) and not (inputs(111));
    layer0_outputs(2487) <= not((inputs(230)) and (inputs(59)));
    layer0_outputs(2488) <= '1';
    layer0_outputs(2489) <= not(inputs(135));
    layer0_outputs(2490) <= not(inputs(2)) or (inputs(28));
    layer0_outputs(2491) <= not(inputs(158));
    layer0_outputs(2492) <= (inputs(85)) or (inputs(74));
    layer0_outputs(2493) <= not(inputs(217)) or (inputs(114));
    layer0_outputs(2494) <= (inputs(106)) xor (inputs(150));
    layer0_outputs(2495) <= (inputs(154)) and not (inputs(183));
    layer0_outputs(2496) <= (inputs(220)) or (inputs(227));
    layer0_outputs(2497) <= (inputs(223)) xor (inputs(109));
    layer0_outputs(2498) <= not(inputs(81));
    layer0_outputs(2499) <= (inputs(91)) and not (inputs(24));
    layer0_outputs(2500) <= '1';
    layer0_outputs(2501) <= inputs(152);
    layer0_outputs(2502) <= inputs(179);
    layer0_outputs(2503) <= (inputs(76)) and not (inputs(51));
    layer0_outputs(2504) <= not((inputs(164)) xor (inputs(35)));
    layer0_outputs(2505) <= '1';
    layer0_outputs(2506) <= not((inputs(225)) or (inputs(9)));
    layer0_outputs(2507) <= (inputs(155)) and not (inputs(106));
    layer0_outputs(2508) <= (inputs(128)) and (inputs(192));
    layer0_outputs(2509) <= '0';
    layer0_outputs(2510) <= not(inputs(6)) or (inputs(75));
    layer0_outputs(2511) <= '0';
    layer0_outputs(2512) <= '0';
    layer0_outputs(2513) <= '1';
    layer0_outputs(2514) <= (inputs(139)) and not (inputs(190));
    layer0_outputs(2515) <= inputs(188);
    layer0_outputs(2516) <= not((inputs(28)) or (inputs(52)));
    layer0_outputs(2517) <= '1';
    layer0_outputs(2518) <= not((inputs(88)) or (inputs(81)));
    layer0_outputs(2519) <= not(inputs(84));
    layer0_outputs(2520) <= not(inputs(24));
    layer0_outputs(2521) <= inputs(184);
    layer0_outputs(2522) <= (inputs(184)) and (inputs(73));
    layer0_outputs(2523) <= '1';
    layer0_outputs(2524) <= (inputs(247)) or (inputs(24));
    layer0_outputs(2525) <= (inputs(124)) and (inputs(79));
    layer0_outputs(2526) <= (inputs(134)) and not (inputs(160));
    layer0_outputs(2527) <= (inputs(255)) and (inputs(173));
    layer0_outputs(2528) <= not((inputs(210)) xor (inputs(75)));
    layer0_outputs(2529) <= '1';
    layer0_outputs(2530) <= not(inputs(226));
    layer0_outputs(2531) <= not(inputs(209)) or (inputs(23));
    layer0_outputs(2532) <= not(inputs(196));
    layer0_outputs(2533) <= not((inputs(80)) and (inputs(62)));
    layer0_outputs(2534) <= (inputs(66)) and not (inputs(125));
    layer0_outputs(2535) <= inputs(216);
    layer0_outputs(2536) <= not((inputs(97)) and (inputs(36)));
    layer0_outputs(2537) <= '1';
    layer0_outputs(2538) <= not((inputs(200)) or (inputs(181)));
    layer0_outputs(2539) <= '0';
    layer0_outputs(2540) <= (inputs(66)) and not (inputs(53));
    layer0_outputs(2541) <= '1';
    layer0_outputs(2542) <= '1';
    layer0_outputs(2543) <= not(inputs(182)) or (inputs(61));
    layer0_outputs(2544) <= (inputs(159)) and not (inputs(159));
    layer0_outputs(2545) <= not((inputs(192)) or (inputs(244)));
    layer0_outputs(2546) <= (inputs(56)) and not (inputs(99));
    layer0_outputs(2547) <= not(inputs(100));
    layer0_outputs(2548) <= '0';
    layer0_outputs(2549) <= not((inputs(56)) or (inputs(38)));
    layer0_outputs(2550) <= '0';
    layer0_outputs(2551) <= not((inputs(159)) xor (inputs(94)));
    layer0_outputs(2552) <= not((inputs(142)) or (inputs(245)));
    layer0_outputs(2553) <= (inputs(42)) and not (inputs(230));
    layer0_outputs(2554) <= not((inputs(130)) or (inputs(29)));
    layer0_outputs(2555) <= not(inputs(89)) or (inputs(220));
    layer0_outputs(2556) <= not(inputs(225)) or (inputs(171));
    layer0_outputs(2557) <= (inputs(156)) xor (inputs(188));
    layer0_outputs(2558) <= (inputs(167)) and not (inputs(162));
    layer0_outputs(2559) <= (inputs(169)) or (inputs(153));
    layer0_outputs(2560) <= not(inputs(13));
    layer0_outputs(2561) <= (inputs(192)) and not (inputs(132));
    layer0_outputs(2562) <= not(inputs(84)) or (inputs(46));
    layer0_outputs(2563) <= (inputs(51)) and (inputs(37));
    layer0_outputs(2564) <= not(inputs(124)) or (inputs(204));
    layer0_outputs(2565) <= inputs(86);
    layer0_outputs(2566) <= not((inputs(58)) and (inputs(217)));
    layer0_outputs(2567) <= (inputs(238)) or (inputs(75));
    layer0_outputs(2568) <= (inputs(26)) and not (inputs(83));
    layer0_outputs(2569) <= '1';
    layer0_outputs(2570) <= not(inputs(45)) or (inputs(54));
    layer0_outputs(2571) <= (inputs(95)) and not (inputs(4));
    layer0_outputs(2572) <= not(inputs(105)) or (inputs(43));
    layer0_outputs(2573) <= not(inputs(165));
    layer0_outputs(2574) <= (inputs(229)) or (inputs(219));
    layer0_outputs(2575) <= not((inputs(1)) and (inputs(60)));
    layer0_outputs(2576) <= (inputs(138)) and not (inputs(37));
    layer0_outputs(2577) <= not(inputs(224));
    layer0_outputs(2578) <= not(inputs(53));
    layer0_outputs(2579) <= inputs(36);
    layer0_outputs(2580) <= not(inputs(91)) or (inputs(3));
    layer0_outputs(2581) <= inputs(26);
    layer0_outputs(2582) <= inputs(211);
    layer0_outputs(2583) <= not(inputs(55)) or (inputs(94));
    layer0_outputs(2584) <= (inputs(124)) and not (inputs(111));
    layer0_outputs(2585) <= (inputs(218)) xor (inputs(242));
    layer0_outputs(2586) <= not((inputs(245)) or (inputs(158)));
    layer0_outputs(2587) <= (inputs(156)) xor (inputs(62));
    layer0_outputs(2588) <= inputs(134);
    layer0_outputs(2589) <= inputs(8);
    layer0_outputs(2590) <= inputs(155);
    layer0_outputs(2591) <= not((inputs(46)) or (inputs(245)));
    layer0_outputs(2592) <= (inputs(55)) or (inputs(41));
    layer0_outputs(2593) <= not((inputs(88)) or (inputs(253)));
    layer0_outputs(2594) <= inputs(136);
    layer0_outputs(2595) <= not((inputs(223)) and (inputs(223)));
    layer0_outputs(2596) <= (inputs(86)) or (inputs(234));
    layer0_outputs(2597) <= (inputs(246)) and (inputs(29));
    layer0_outputs(2598) <= inputs(60);
    layer0_outputs(2599) <= '0';
    layer0_outputs(2600) <= (inputs(90)) and not (inputs(41));
    layer0_outputs(2601) <= not((inputs(61)) and (inputs(226)));
    layer0_outputs(2602) <= inputs(18);
    layer0_outputs(2603) <= '1';
    layer0_outputs(2604) <= not(inputs(63)) or (inputs(207));
    layer0_outputs(2605) <= (inputs(43)) and (inputs(246));
    layer0_outputs(2606) <= not((inputs(82)) xor (inputs(1)));
    layer0_outputs(2607) <= not((inputs(194)) xor (inputs(145)));
    layer0_outputs(2608) <= (inputs(193)) xor (inputs(237));
    layer0_outputs(2609) <= not(inputs(200)) or (inputs(122));
    layer0_outputs(2610) <= not(inputs(57));
    layer0_outputs(2611) <= not(inputs(53));
    layer0_outputs(2612) <= (inputs(80)) xor (inputs(113));
    layer0_outputs(2613) <= not(inputs(191)) or (inputs(251));
    layer0_outputs(2614) <= inputs(57);
    layer0_outputs(2615) <= not(inputs(186)) or (inputs(248));
    layer0_outputs(2616) <= (inputs(80)) xor (inputs(125));
    layer0_outputs(2617) <= inputs(28);
    layer0_outputs(2618) <= not(inputs(26)) or (inputs(18));
    layer0_outputs(2619) <= '0';
    layer0_outputs(2620) <= (inputs(240)) and not (inputs(47));
    layer0_outputs(2621) <= inputs(93);
    layer0_outputs(2622) <= not(inputs(64));
    layer0_outputs(2623) <= (inputs(161)) xor (inputs(254));
    layer0_outputs(2624) <= inputs(44);
    layer0_outputs(2625) <= (inputs(127)) and not (inputs(79));
    layer0_outputs(2626) <= not(inputs(113));
    layer0_outputs(2627) <= inputs(236);
    layer0_outputs(2628) <= inputs(221);
    layer0_outputs(2629) <= (inputs(141)) or (inputs(116));
    layer0_outputs(2630) <= (inputs(210)) and not (inputs(142));
    layer0_outputs(2631) <= '0';
    layer0_outputs(2632) <= (inputs(189)) and not (inputs(61));
    layer0_outputs(2633) <= (inputs(142)) and not (inputs(150));
    layer0_outputs(2634) <= not((inputs(132)) or (inputs(85)));
    layer0_outputs(2635) <= (inputs(94)) or (inputs(219));
    layer0_outputs(2636) <= (inputs(114)) xor (inputs(90));
    layer0_outputs(2637) <= (inputs(75)) and not (inputs(106));
    layer0_outputs(2638) <= (inputs(12)) or (inputs(88));
    layer0_outputs(2639) <= (inputs(178)) or (inputs(163));
    layer0_outputs(2640) <= (inputs(39)) and not (inputs(209));
    layer0_outputs(2641) <= not(inputs(92));
    layer0_outputs(2642) <= (inputs(170)) or (inputs(77));
    layer0_outputs(2643) <= '1';
    layer0_outputs(2644) <= '0';
    layer0_outputs(2645) <= not(inputs(63));
    layer0_outputs(2646) <= not(inputs(149));
    layer0_outputs(2647) <= (inputs(153)) and not (inputs(198));
    layer0_outputs(2648) <= inputs(90);
    layer0_outputs(2649) <= (inputs(241)) xor (inputs(199));
    layer0_outputs(2650) <= not(inputs(4)) or (inputs(63));
    layer0_outputs(2651) <= (inputs(219)) and (inputs(241));
    layer0_outputs(2652) <= '1';
    layer0_outputs(2653) <= not(inputs(89)) or (inputs(171));
    layer0_outputs(2654) <= (inputs(224)) or (inputs(162));
    layer0_outputs(2655) <= (inputs(32)) xor (inputs(89));
    layer0_outputs(2656) <= inputs(62);
    layer0_outputs(2657) <= not(inputs(207));
    layer0_outputs(2658) <= not(inputs(54));
    layer0_outputs(2659) <= not(inputs(94));
    layer0_outputs(2660) <= inputs(160);
    layer0_outputs(2661) <= not(inputs(63));
    layer0_outputs(2662) <= (inputs(158)) and not (inputs(209));
    layer0_outputs(2663) <= not(inputs(193));
    layer0_outputs(2664) <= inputs(215);
    layer0_outputs(2665) <= (inputs(92)) and not (inputs(150));
    layer0_outputs(2666) <= inputs(12);
    layer0_outputs(2667) <= not(inputs(88));
    layer0_outputs(2668) <= not(inputs(141)) or (inputs(149));
    layer0_outputs(2669) <= '1';
    layer0_outputs(2670) <= '1';
    layer0_outputs(2671) <= (inputs(155)) xor (inputs(242));
    layer0_outputs(2672) <= not((inputs(80)) and (inputs(111)));
    layer0_outputs(2673) <= (inputs(10)) xor (inputs(167));
    layer0_outputs(2674) <= (inputs(162)) and (inputs(17));
    layer0_outputs(2675) <= not(inputs(207));
    layer0_outputs(2676) <= (inputs(70)) and not (inputs(178));
    layer0_outputs(2677) <= (inputs(63)) or (inputs(84));
    layer0_outputs(2678) <= not(inputs(120));
    layer0_outputs(2679) <= (inputs(93)) xor (inputs(221));
    layer0_outputs(2680) <= not((inputs(81)) xor (inputs(156)));
    layer0_outputs(2681) <= '0';
    layer0_outputs(2682) <= (inputs(53)) and not (inputs(209));
    layer0_outputs(2683) <= not((inputs(18)) or (inputs(160)));
    layer0_outputs(2684) <= inputs(223);
    layer0_outputs(2685) <= not(inputs(117)) or (inputs(41));
    layer0_outputs(2686) <= not((inputs(58)) and (inputs(182)));
    layer0_outputs(2687) <= (inputs(171)) or (inputs(181));
    layer0_outputs(2688) <= (inputs(211)) or (inputs(245));
    layer0_outputs(2689) <= not((inputs(4)) or (inputs(224)));
    layer0_outputs(2690) <= (inputs(47)) and (inputs(255));
    layer0_outputs(2691) <= '0';
    layer0_outputs(2692) <= not(inputs(88));
    layer0_outputs(2693) <= (inputs(237)) or (inputs(33));
    layer0_outputs(2694) <= (inputs(2)) xor (inputs(95));
    layer0_outputs(2695) <= not(inputs(196));
    layer0_outputs(2696) <= not(inputs(171)) or (inputs(81));
    layer0_outputs(2697) <= inputs(137);
    layer0_outputs(2698) <= '1';
    layer0_outputs(2699) <= not(inputs(59)) or (inputs(47));
    layer0_outputs(2700) <= (inputs(16)) or (inputs(218));
    layer0_outputs(2701) <= '0';
    layer0_outputs(2702) <= not(inputs(73)) or (inputs(248));
    layer0_outputs(2703) <= not(inputs(47)) or (inputs(196));
    layer0_outputs(2704) <= (inputs(183)) and not (inputs(182));
    layer0_outputs(2705) <= not(inputs(137));
    layer0_outputs(2706) <= not(inputs(207)) or (inputs(80));
    layer0_outputs(2707) <= '0';
    layer0_outputs(2708) <= not(inputs(92));
    layer0_outputs(2709) <= (inputs(184)) and (inputs(14));
    layer0_outputs(2710) <= not(inputs(108)) or (inputs(23));
    layer0_outputs(2711) <= (inputs(66)) or (inputs(141));
    layer0_outputs(2712) <= (inputs(10)) xor (inputs(123));
    layer0_outputs(2713) <= inputs(63);
    layer0_outputs(2714) <= '0';
    layer0_outputs(2715) <= (inputs(114)) and (inputs(61));
    layer0_outputs(2716) <= (inputs(207)) and not (inputs(76));
    layer0_outputs(2717) <= not((inputs(216)) or (inputs(145)));
    layer0_outputs(2718) <= not(inputs(157));
    layer0_outputs(2719) <= '0';
    layer0_outputs(2720) <= (inputs(168)) and not (inputs(226));
    layer0_outputs(2721) <= not(inputs(115)) or (inputs(114));
    layer0_outputs(2722) <= (inputs(53)) and not (inputs(232));
    layer0_outputs(2723) <= not(inputs(159)) or (inputs(45));
    layer0_outputs(2724) <= inputs(173);
    layer0_outputs(2725) <= (inputs(121)) and not (inputs(5));
    layer0_outputs(2726) <= not(inputs(39));
    layer0_outputs(2727) <= not((inputs(153)) or (inputs(144)));
    layer0_outputs(2728) <= not((inputs(186)) xor (inputs(60)));
    layer0_outputs(2729) <= (inputs(239)) or (inputs(234));
    layer0_outputs(2730) <= not(inputs(249));
    layer0_outputs(2731) <= not(inputs(252)) or (inputs(188));
    layer0_outputs(2732) <= (inputs(36)) and not (inputs(226));
    layer0_outputs(2733) <= not(inputs(88)) or (inputs(152));
    layer0_outputs(2734) <= '0';
    layer0_outputs(2735) <= not(inputs(7)) or (inputs(175));
    layer0_outputs(2736) <= (inputs(217)) or (inputs(127));
    layer0_outputs(2737) <= (inputs(65)) xor (inputs(105));
    layer0_outputs(2738) <= not((inputs(146)) xor (inputs(255)));
    layer0_outputs(2739) <= not(inputs(7));
    layer0_outputs(2740) <= not((inputs(128)) or (inputs(157)));
    layer0_outputs(2741) <= (inputs(8)) and not (inputs(20));
    layer0_outputs(2742) <= (inputs(81)) and not (inputs(13));
    layer0_outputs(2743) <= inputs(206);
    layer0_outputs(2744) <= not(inputs(124));
    layer0_outputs(2745) <= not((inputs(21)) xor (inputs(10)));
    layer0_outputs(2746) <= not(inputs(26));
    layer0_outputs(2747) <= (inputs(49)) and (inputs(249));
    layer0_outputs(2748) <= not(inputs(20));
    layer0_outputs(2749) <= (inputs(91)) or (inputs(36));
    layer0_outputs(2750) <= not(inputs(100));
    layer0_outputs(2751) <= (inputs(171)) and not (inputs(123));
    layer0_outputs(2752) <= (inputs(221)) and not (inputs(165));
    layer0_outputs(2753) <= (inputs(121)) and not (inputs(109));
    layer0_outputs(2754) <= not((inputs(169)) and (inputs(237)));
    layer0_outputs(2755) <= inputs(130);
    layer0_outputs(2756) <= (inputs(193)) and (inputs(11));
    layer0_outputs(2757) <= not((inputs(16)) or (inputs(104)));
    layer0_outputs(2758) <= (inputs(70)) and not (inputs(177));
    layer0_outputs(2759) <= '0';
    layer0_outputs(2760) <= '1';
    layer0_outputs(2761) <= '1';
    layer0_outputs(2762) <= (inputs(124)) xor (inputs(240));
    layer0_outputs(2763) <= not((inputs(101)) xor (inputs(201)));
    layer0_outputs(2764) <= inputs(66);
    layer0_outputs(2765) <= not(inputs(74));
    layer0_outputs(2766) <= (inputs(240)) and not (inputs(228));
    layer0_outputs(2767) <= not((inputs(36)) or (inputs(194)));
    layer0_outputs(2768) <= (inputs(157)) and (inputs(237));
    layer0_outputs(2769) <= not(inputs(150));
    layer0_outputs(2770) <= inputs(61);
    layer0_outputs(2771) <= (inputs(242)) or (inputs(50));
    layer0_outputs(2772) <= (inputs(142)) and not (inputs(193));
    layer0_outputs(2773) <= (inputs(66)) and not (inputs(169));
    layer0_outputs(2774) <= inputs(76);
    layer0_outputs(2775) <= (inputs(226)) and (inputs(252));
    layer0_outputs(2776) <= (inputs(65)) xor (inputs(223));
    layer0_outputs(2777) <= (inputs(64)) xor (inputs(197));
    layer0_outputs(2778) <= not(inputs(211));
    layer0_outputs(2779) <= not((inputs(115)) or (inputs(216)));
    layer0_outputs(2780) <= not(inputs(174));
    layer0_outputs(2781) <= (inputs(103)) and not (inputs(37));
    layer0_outputs(2782) <= not((inputs(143)) or (inputs(41)));
    layer0_outputs(2783) <= (inputs(5)) and not (inputs(18));
    layer0_outputs(2784) <= (inputs(157)) and not (inputs(14));
    layer0_outputs(2785) <= inputs(71);
    layer0_outputs(2786) <= inputs(134);
    layer0_outputs(2787) <= not(inputs(32));
    layer0_outputs(2788) <= not((inputs(131)) and (inputs(172)));
    layer0_outputs(2789) <= inputs(141);
    layer0_outputs(2790) <= '1';
    layer0_outputs(2791) <= (inputs(220)) or (inputs(164));
    layer0_outputs(2792) <= (inputs(181)) and not (inputs(96));
    layer0_outputs(2793) <= inputs(24);
    layer0_outputs(2794) <= not(inputs(122)) or (inputs(46));
    layer0_outputs(2795) <= (inputs(42)) and (inputs(233));
    layer0_outputs(2796) <= not((inputs(88)) or (inputs(231)));
    layer0_outputs(2797) <= '0';
    layer0_outputs(2798) <= not(inputs(114)) or (inputs(42));
    layer0_outputs(2799) <= inputs(201);
    layer0_outputs(2800) <= (inputs(184)) xor (inputs(78));
    layer0_outputs(2801) <= not(inputs(21));
    layer0_outputs(2802) <= (inputs(199)) and not (inputs(238));
    layer0_outputs(2803) <= (inputs(33)) xor (inputs(155));
    layer0_outputs(2804) <= '1';
    layer0_outputs(2805) <= not((inputs(191)) xor (inputs(114)));
    layer0_outputs(2806) <= inputs(163);
    layer0_outputs(2807) <= (inputs(154)) or (inputs(172));
    layer0_outputs(2808) <= not(inputs(4));
    layer0_outputs(2809) <= not((inputs(71)) xor (inputs(151)));
    layer0_outputs(2810) <= inputs(104);
    layer0_outputs(2811) <= (inputs(174)) xor (inputs(34));
    layer0_outputs(2812) <= not(inputs(121)) or (inputs(234));
    layer0_outputs(2813) <= not((inputs(166)) or (inputs(40)));
    layer0_outputs(2814) <= '0';
    layer0_outputs(2815) <= (inputs(247)) or (inputs(45));
    layer0_outputs(2816) <= not((inputs(12)) or (inputs(180)));
    layer0_outputs(2817) <= (inputs(177)) and (inputs(219));
    layer0_outputs(2818) <= not(inputs(137));
    layer0_outputs(2819) <= (inputs(41)) and not (inputs(43));
    layer0_outputs(2820) <= (inputs(85)) and (inputs(31));
    layer0_outputs(2821) <= not(inputs(29));
    layer0_outputs(2822) <= (inputs(164)) or (inputs(137));
    layer0_outputs(2823) <= (inputs(102)) or (inputs(246));
    layer0_outputs(2824) <= not(inputs(120));
    layer0_outputs(2825) <= (inputs(86)) xor (inputs(79));
    layer0_outputs(2826) <= not((inputs(187)) or (inputs(194)));
    layer0_outputs(2827) <= inputs(199);
    layer0_outputs(2828) <= (inputs(164)) or (inputs(158));
    layer0_outputs(2829) <= (inputs(247)) and not (inputs(7));
    layer0_outputs(2830) <= (inputs(78)) or (inputs(60));
    layer0_outputs(2831) <= inputs(52);
    layer0_outputs(2832) <= (inputs(233)) and not (inputs(16));
    layer0_outputs(2833) <= (inputs(110)) and not (inputs(250));
    layer0_outputs(2834) <= not(inputs(171));
    layer0_outputs(2835) <= not(inputs(251)) or (inputs(241));
    layer0_outputs(2836) <= not((inputs(19)) and (inputs(113)));
    layer0_outputs(2837) <= not((inputs(127)) xor (inputs(208)));
    layer0_outputs(2838) <= not(inputs(115)) or (inputs(229));
    layer0_outputs(2839) <= (inputs(254)) or (inputs(133));
    layer0_outputs(2840) <= not((inputs(184)) and (inputs(107)));
    layer0_outputs(2841) <= (inputs(112)) xor (inputs(188));
    layer0_outputs(2842) <= '1';
    layer0_outputs(2843) <= (inputs(243)) and (inputs(26));
    layer0_outputs(2844) <= '0';
    layer0_outputs(2845) <= not(inputs(240));
    layer0_outputs(2846) <= (inputs(118)) or (inputs(182));
    layer0_outputs(2847) <= not((inputs(13)) or (inputs(210)));
    layer0_outputs(2848) <= '1';
    layer0_outputs(2849) <= '1';
    layer0_outputs(2850) <= not(inputs(227)) or (inputs(88));
    layer0_outputs(2851) <= inputs(130);
    layer0_outputs(2852) <= (inputs(160)) xor (inputs(149));
    layer0_outputs(2853) <= (inputs(236)) or (inputs(69));
    layer0_outputs(2854) <= inputs(49);
    layer0_outputs(2855) <= (inputs(238)) xor (inputs(223));
    layer0_outputs(2856) <= (inputs(81)) or (inputs(182));
    layer0_outputs(2857) <= (inputs(54)) xor (inputs(206));
    layer0_outputs(2858) <= not((inputs(191)) or (inputs(183)));
    layer0_outputs(2859) <= (inputs(200)) and not (inputs(163));
    layer0_outputs(2860) <= (inputs(104)) xor (inputs(112));
    layer0_outputs(2861) <= (inputs(186)) or (inputs(246));
    layer0_outputs(2862) <= (inputs(141)) and not (inputs(8));
    layer0_outputs(2863) <= '1';
    layer0_outputs(2864) <= not(inputs(94)) or (inputs(227));
    layer0_outputs(2865) <= (inputs(202)) or (inputs(38));
    layer0_outputs(2866) <= not((inputs(74)) xor (inputs(176)));
    layer0_outputs(2867) <= not(inputs(115)) or (inputs(184));
    layer0_outputs(2868) <= not((inputs(233)) xor (inputs(102)));
    layer0_outputs(2869) <= not(inputs(171)) or (inputs(128));
    layer0_outputs(2870) <= '0';
    layer0_outputs(2871) <= inputs(194);
    layer0_outputs(2872) <= (inputs(136)) and not (inputs(209));
    layer0_outputs(2873) <= not(inputs(223)) or (inputs(78));
    layer0_outputs(2874) <= '0';
    layer0_outputs(2875) <= not((inputs(196)) and (inputs(21)));
    layer0_outputs(2876) <= '0';
    layer0_outputs(2877) <= (inputs(127)) xor (inputs(63));
    layer0_outputs(2878) <= (inputs(157)) or (inputs(233));
    layer0_outputs(2879) <= not(inputs(181)) or (inputs(111));
    layer0_outputs(2880) <= not((inputs(225)) xor (inputs(161)));
    layer0_outputs(2881) <= not(inputs(22));
    layer0_outputs(2882) <= not((inputs(170)) or (inputs(59)));
    layer0_outputs(2883) <= '0';
    layer0_outputs(2884) <= '1';
    layer0_outputs(2885) <= (inputs(105)) or (inputs(194));
    layer0_outputs(2886) <= not(inputs(234));
    layer0_outputs(2887) <= (inputs(156)) xor (inputs(254));
    layer0_outputs(2888) <= inputs(124);
    layer0_outputs(2889) <= inputs(174);
    layer0_outputs(2890) <= inputs(204);
    layer0_outputs(2891) <= not(inputs(74)) or (inputs(28));
    layer0_outputs(2892) <= (inputs(118)) xor (inputs(19));
    layer0_outputs(2893) <= not((inputs(105)) and (inputs(50)));
    layer0_outputs(2894) <= (inputs(150)) or (inputs(178));
    layer0_outputs(2895) <= inputs(30);
    layer0_outputs(2896) <= not(inputs(222)) or (inputs(46));
    layer0_outputs(2897) <= not((inputs(91)) or (inputs(65)));
    layer0_outputs(2898) <= inputs(78);
    layer0_outputs(2899) <= (inputs(135)) and not (inputs(158));
    layer0_outputs(2900) <= (inputs(38)) or (inputs(231));
    layer0_outputs(2901) <= (inputs(171)) or (inputs(56));
    layer0_outputs(2902) <= not(inputs(123)) or (inputs(35));
    layer0_outputs(2903) <= (inputs(239)) or (inputs(108));
    layer0_outputs(2904) <= inputs(52);
    layer0_outputs(2905) <= '1';
    layer0_outputs(2906) <= '0';
    layer0_outputs(2907) <= (inputs(118)) or (inputs(145));
    layer0_outputs(2908) <= '1';
    layer0_outputs(2909) <= not(inputs(126));
    layer0_outputs(2910) <= inputs(224);
    layer0_outputs(2911) <= (inputs(230)) and not (inputs(86));
    layer0_outputs(2912) <= not((inputs(170)) xor (inputs(17)));
    layer0_outputs(2913) <= (inputs(57)) and not (inputs(44));
    layer0_outputs(2914) <= not(inputs(179));
    layer0_outputs(2915) <= not(inputs(252));
    layer0_outputs(2916) <= (inputs(167)) or (inputs(174));
    layer0_outputs(2917) <= (inputs(106)) and not (inputs(156));
    layer0_outputs(2918) <= (inputs(23)) or (inputs(155));
    layer0_outputs(2919) <= '0';
    layer0_outputs(2920) <= not(inputs(135)) or (inputs(236));
    layer0_outputs(2921) <= (inputs(15)) and (inputs(108));
    layer0_outputs(2922) <= not((inputs(203)) xor (inputs(4)));
    layer0_outputs(2923) <= not(inputs(156));
    layer0_outputs(2924) <= not(inputs(209));
    layer0_outputs(2925) <= '1';
    layer0_outputs(2926) <= not((inputs(176)) or (inputs(197)));
    layer0_outputs(2927) <= not(inputs(49));
    layer0_outputs(2928) <= '0';
    layer0_outputs(2929) <= (inputs(68)) and not (inputs(1));
    layer0_outputs(2930) <= inputs(165);
    layer0_outputs(2931) <= inputs(206);
    layer0_outputs(2932) <= (inputs(74)) and not (inputs(125));
    layer0_outputs(2933) <= not((inputs(208)) or (inputs(253)));
    layer0_outputs(2934) <= not(inputs(121));
    layer0_outputs(2935) <= (inputs(85)) or (inputs(147));
    layer0_outputs(2936) <= (inputs(229)) and not (inputs(62));
    layer0_outputs(2937) <= inputs(1);
    layer0_outputs(2938) <= '0';
    layer0_outputs(2939) <= not(inputs(206)) or (inputs(94));
    layer0_outputs(2940) <= not(inputs(123)) or (inputs(128));
    layer0_outputs(2941) <= (inputs(126)) or (inputs(73));
    layer0_outputs(2942) <= not((inputs(237)) or (inputs(234)));
    layer0_outputs(2943) <= not((inputs(99)) xor (inputs(242)));
    layer0_outputs(2944) <= not((inputs(235)) or (inputs(234)));
    layer0_outputs(2945) <= inputs(108);
    layer0_outputs(2946) <= '0';
    layer0_outputs(2947) <= not((inputs(128)) and (inputs(181)));
    layer0_outputs(2948) <= not(inputs(92));
    layer0_outputs(2949) <= not((inputs(146)) and (inputs(51)));
    layer0_outputs(2950) <= not(inputs(180)) or (inputs(63));
    layer0_outputs(2951) <= (inputs(88)) or (inputs(82));
    layer0_outputs(2952) <= (inputs(91)) or (inputs(115));
    layer0_outputs(2953) <= not(inputs(192));
    layer0_outputs(2954) <= (inputs(169)) xor (inputs(87));
    layer0_outputs(2955) <= (inputs(171)) and not (inputs(75));
    layer0_outputs(2956) <= (inputs(184)) and not (inputs(229));
    layer0_outputs(2957) <= not(inputs(182)) or (inputs(95));
    layer0_outputs(2958) <= not(inputs(54));
    layer0_outputs(2959) <= (inputs(100)) and not (inputs(62));
    layer0_outputs(2960) <= inputs(102);
    layer0_outputs(2961) <= (inputs(57)) xor (inputs(111));
    layer0_outputs(2962) <= not(inputs(190)) or (inputs(47));
    layer0_outputs(2963) <= not(inputs(240)) or (inputs(29));
    layer0_outputs(2964) <= (inputs(164)) or (inputs(51));
    layer0_outputs(2965) <= not((inputs(253)) xor (inputs(217)));
    layer0_outputs(2966) <= (inputs(145)) and (inputs(145));
    layer0_outputs(2967) <= '1';
    layer0_outputs(2968) <= not((inputs(201)) and (inputs(215)));
    layer0_outputs(2969) <= '1';
    layer0_outputs(2970) <= (inputs(222)) xor (inputs(47));
    layer0_outputs(2971) <= '1';
    layer0_outputs(2972) <= (inputs(68)) and not (inputs(40));
    layer0_outputs(2973) <= inputs(234);
    layer0_outputs(2974) <= not(inputs(103)) or (inputs(227));
    layer0_outputs(2975) <= inputs(168);
    layer0_outputs(2976) <= not(inputs(152)) or (inputs(99));
    layer0_outputs(2977) <= (inputs(18)) and (inputs(143));
    layer0_outputs(2978) <= inputs(51);
    layer0_outputs(2979) <= not(inputs(61)) or (inputs(175));
    layer0_outputs(2980) <= not(inputs(164)) or (inputs(45));
    layer0_outputs(2981) <= not(inputs(124));
    layer0_outputs(2982) <= not((inputs(14)) xor (inputs(48)));
    layer0_outputs(2983) <= (inputs(139)) or (inputs(172));
    layer0_outputs(2984) <= (inputs(82)) or (inputs(106));
    layer0_outputs(2985) <= (inputs(218)) or (inputs(86));
    layer0_outputs(2986) <= '0';
    layer0_outputs(2987) <= not(inputs(32)) or (inputs(250));
    layer0_outputs(2988) <= (inputs(216)) or (inputs(223));
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= inputs(127);
    layer0_outputs(2991) <= (inputs(181)) xor (inputs(82));
    layer0_outputs(2992) <= inputs(193);
    layer0_outputs(2993) <= not((inputs(105)) or (inputs(60)));
    layer0_outputs(2994) <= not((inputs(137)) xor (inputs(143)));
    layer0_outputs(2995) <= (inputs(43)) xor (inputs(206));
    layer0_outputs(2996) <= (inputs(1)) and not (inputs(139));
    layer0_outputs(2997) <= (inputs(212)) or (inputs(28));
    layer0_outputs(2998) <= not((inputs(99)) and (inputs(170)));
    layer0_outputs(2999) <= not(inputs(201));
    layer0_outputs(3000) <= not((inputs(90)) or (inputs(209)));
    layer0_outputs(3001) <= inputs(241);
    layer0_outputs(3002) <= '0';
    layer0_outputs(3003) <= '0';
    layer0_outputs(3004) <= not(inputs(120));
    layer0_outputs(3005) <= '0';
    layer0_outputs(3006) <= not((inputs(154)) or (inputs(160)));
    layer0_outputs(3007) <= (inputs(253)) and (inputs(123));
    layer0_outputs(3008) <= (inputs(184)) and (inputs(129));
    layer0_outputs(3009) <= (inputs(148)) and not (inputs(92));
    layer0_outputs(3010) <= '0';
    layer0_outputs(3011) <= (inputs(152)) and not (inputs(113));
    layer0_outputs(3012) <= (inputs(105)) or (inputs(216));
    layer0_outputs(3013) <= not(inputs(249));
    layer0_outputs(3014) <= not(inputs(133));
    layer0_outputs(3015) <= (inputs(208)) xor (inputs(198));
    layer0_outputs(3016) <= (inputs(217)) or (inputs(229));
    layer0_outputs(3017) <= inputs(192);
    layer0_outputs(3018) <= (inputs(234)) and (inputs(14));
    layer0_outputs(3019) <= not((inputs(67)) xor (inputs(106)));
    layer0_outputs(3020) <= not((inputs(117)) or (inputs(231)));
    layer0_outputs(3021) <= not((inputs(47)) xor (inputs(232)));
    layer0_outputs(3022) <= (inputs(224)) and not (inputs(221));
    layer0_outputs(3023) <= inputs(87);
    layer0_outputs(3024) <= inputs(180);
    layer0_outputs(3025) <= not((inputs(169)) or (inputs(191)));
    layer0_outputs(3026) <= (inputs(122)) or (inputs(227));
    layer0_outputs(3027) <= (inputs(95)) xor (inputs(119));
    layer0_outputs(3028) <= inputs(164);
    layer0_outputs(3029) <= not((inputs(210)) and (inputs(177)));
    layer0_outputs(3030) <= not(inputs(252));
    layer0_outputs(3031) <= (inputs(198)) and (inputs(87));
    layer0_outputs(3032) <= not(inputs(10));
    layer0_outputs(3033) <= not((inputs(90)) or (inputs(63)));
    layer0_outputs(3034) <= (inputs(221)) and not (inputs(204));
    layer0_outputs(3035) <= not(inputs(30));
    layer0_outputs(3036) <= not(inputs(172));
    layer0_outputs(3037) <= not((inputs(154)) xor (inputs(23)));
    layer0_outputs(3038) <= (inputs(82)) and not (inputs(91));
    layer0_outputs(3039) <= not((inputs(94)) or (inputs(185)));
    layer0_outputs(3040) <= (inputs(74)) and not (inputs(39));
    layer0_outputs(3041) <= not((inputs(154)) or (inputs(242)));
    layer0_outputs(3042) <= (inputs(100)) and not (inputs(174));
    layer0_outputs(3043) <= not(inputs(31)) or (inputs(185));
    layer0_outputs(3044) <= '1';
    layer0_outputs(3045) <= (inputs(246)) xor (inputs(59));
    layer0_outputs(3046) <= not(inputs(126));
    layer0_outputs(3047) <= not((inputs(247)) or (inputs(38)));
    layer0_outputs(3048) <= (inputs(223)) or (inputs(186));
    layer0_outputs(3049) <= not((inputs(54)) xor (inputs(163)));
    layer0_outputs(3050) <= not((inputs(85)) and (inputs(73)));
    layer0_outputs(3051) <= not((inputs(210)) xor (inputs(40)));
    layer0_outputs(3052) <= inputs(116);
    layer0_outputs(3053) <= (inputs(13)) and not (inputs(228));
    layer0_outputs(3054) <= not(inputs(148));
    layer0_outputs(3055) <= (inputs(89)) and not (inputs(170));
    layer0_outputs(3056) <= '1';
    layer0_outputs(3057) <= inputs(134);
    layer0_outputs(3058) <= (inputs(3)) and (inputs(22));
    layer0_outputs(3059) <= not(inputs(28));
    layer0_outputs(3060) <= '0';
    layer0_outputs(3061) <= (inputs(137)) and (inputs(84));
    layer0_outputs(3062) <= not((inputs(106)) and (inputs(73)));
    layer0_outputs(3063) <= not(inputs(149));
    layer0_outputs(3064) <= (inputs(212)) and not (inputs(190));
    layer0_outputs(3065) <= not((inputs(218)) and (inputs(93)));
    layer0_outputs(3066) <= inputs(160);
    layer0_outputs(3067) <= (inputs(40)) and not (inputs(179));
    layer0_outputs(3068) <= not(inputs(50));
    layer0_outputs(3069) <= not((inputs(229)) or (inputs(140)));
    layer0_outputs(3070) <= (inputs(209)) xor (inputs(197));
    layer0_outputs(3071) <= not(inputs(66)) or (inputs(26));
    layer0_outputs(3072) <= '1';
    layer0_outputs(3073) <= '1';
    layer0_outputs(3074) <= (inputs(188)) xor (inputs(93));
    layer0_outputs(3075) <= not(inputs(155));
    layer0_outputs(3076) <= (inputs(50)) and not (inputs(100));
    layer0_outputs(3077) <= not((inputs(120)) and (inputs(84)));
    layer0_outputs(3078) <= not((inputs(120)) or (inputs(36)));
    layer0_outputs(3079) <= '0';
    layer0_outputs(3080) <= inputs(249);
    layer0_outputs(3081) <= not(inputs(16));
    layer0_outputs(3082) <= inputs(121);
    layer0_outputs(3083) <= (inputs(186)) and not (inputs(78));
    layer0_outputs(3084) <= (inputs(204)) and not (inputs(113));
    layer0_outputs(3085) <= (inputs(147)) and (inputs(16));
    layer0_outputs(3086) <= '1';
    layer0_outputs(3087) <= not(inputs(41)) or (inputs(210));
    layer0_outputs(3088) <= not((inputs(126)) xor (inputs(158)));
    layer0_outputs(3089) <= not(inputs(204));
    layer0_outputs(3090) <= not(inputs(63)) or (inputs(149));
    layer0_outputs(3091) <= (inputs(196)) and not (inputs(107));
    layer0_outputs(3092) <= '0';
    layer0_outputs(3093) <= inputs(125);
    layer0_outputs(3094) <= not((inputs(221)) xor (inputs(14)));
    layer0_outputs(3095) <= inputs(132);
    layer0_outputs(3096) <= (inputs(46)) and not (inputs(192));
    layer0_outputs(3097) <= not(inputs(150)) or (inputs(157));
    layer0_outputs(3098) <= (inputs(102)) and not (inputs(177));
    layer0_outputs(3099) <= (inputs(131)) xor (inputs(131));
    layer0_outputs(3100) <= not((inputs(55)) or (inputs(182)));
    layer0_outputs(3101) <= not(inputs(97)) or (inputs(227));
    layer0_outputs(3102) <= not((inputs(113)) or (inputs(140)));
    layer0_outputs(3103) <= not((inputs(237)) or (inputs(9)));
    layer0_outputs(3104) <= not((inputs(17)) or (inputs(29)));
    layer0_outputs(3105) <= not((inputs(15)) or (inputs(56)));
    layer0_outputs(3106) <= (inputs(240)) or (inputs(248));
    layer0_outputs(3107) <= (inputs(93)) xor (inputs(223));
    layer0_outputs(3108) <= not(inputs(61)) or (inputs(190));
    layer0_outputs(3109) <= (inputs(237)) xor (inputs(232));
    layer0_outputs(3110) <= (inputs(173)) and (inputs(107));
    layer0_outputs(3111) <= inputs(149);
    layer0_outputs(3112) <= (inputs(119)) xor (inputs(126));
    layer0_outputs(3113) <= inputs(41);
    layer0_outputs(3114) <= not(inputs(91)) or (inputs(45));
    layer0_outputs(3115) <= not(inputs(239)) or (inputs(36));
    layer0_outputs(3116) <= (inputs(1)) xor (inputs(205));
    layer0_outputs(3117) <= not((inputs(239)) or (inputs(198)));
    layer0_outputs(3118) <= (inputs(196)) xor (inputs(112));
    layer0_outputs(3119) <= not(inputs(26)) or (inputs(76));
    layer0_outputs(3120) <= not((inputs(40)) and (inputs(31)));
    layer0_outputs(3121) <= '1';
    layer0_outputs(3122) <= not(inputs(23));
    layer0_outputs(3123) <= (inputs(54)) or (inputs(78));
    layer0_outputs(3124) <= '0';
    layer0_outputs(3125) <= (inputs(121)) and (inputs(16));
    layer0_outputs(3126) <= not(inputs(140));
    layer0_outputs(3127) <= not(inputs(83));
    layer0_outputs(3128) <= (inputs(37)) and not (inputs(241));
    layer0_outputs(3129) <= not((inputs(159)) xor (inputs(19)));
    layer0_outputs(3130) <= (inputs(142)) or (inputs(183));
    layer0_outputs(3131) <= (inputs(44)) xor (inputs(81));
    layer0_outputs(3132) <= '0';
    layer0_outputs(3133) <= not(inputs(112));
    layer0_outputs(3134) <= (inputs(26)) and not (inputs(58));
    layer0_outputs(3135) <= (inputs(232)) and not (inputs(60));
    layer0_outputs(3136) <= not(inputs(104)) or (inputs(53));
    layer0_outputs(3137) <= not(inputs(120));
    layer0_outputs(3138) <= '0';
    layer0_outputs(3139) <= inputs(79);
    layer0_outputs(3140) <= not((inputs(130)) xor (inputs(53)));
    layer0_outputs(3141) <= not(inputs(250));
    layer0_outputs(3142) <= (inputs(122)) or (inputs(202));
    layer0_outputs(3143) <= not((inputs(125)) xor (inputs(202)));
    layer0_outputs(3144) <= not((inputs(188)) and (inputs(249)));
    layer0_outputs(3145) <= (inputs(57)) or (inputs(109));
    layer0_outputs(3146) <= not((inputs(174)) xor (inputs(181)));
    layer0_outputs(3147) <= not(inputs(190)) or (inputs(76));
    layer0_outputs(3148) <= inputs(134);
    layer0_outputs(3149) <= (inputs(148)) and (inputs(121));
    layer0_outputs(3150) <= not(inputs(233)) or (inputs(240));
    layer0_outputs(3151) <= not(inputs(68));
    layer0_outputs(3152) <= (inputs(170)) xor (inputs(241));
    layer0_outputs(3153) <= not((inputs(81)) or (inputs(69)));
    layer0_outputs(3154) <= inputs(37);
    layer0_outputs(3155) <= not((inputs(234)) or (inputs(46)));
    layer0_outputs(3156) <= not(inputs(139)) or (inputs(18));
    layer0_outputs(3157) <= not(inputs(109));
    layer0_outputs(3158) <= not((inputs(191)) or (inputs(182)));
    layer0_outputs(3159) <= not((inputs(241)) xor (inputs(151)));
    layer0_outputs(3160) <= (inputs(10)) or (inputs(240));
    layer0_outputs(3161) <= inputs(38);
    layer0_outputs(3162) <= not(inputs(184)) or (inputs(203));
    layer0_outputs(3163) <= (inputs(110)) and (inputs(44));
    layer0_outputs(3164) <= (inputs(195)) and not (inputs(76));
    layer0_outputs(3165) <= (inputs(33)) and not (inputs(70));
    layer0_outputs(3166) <= '1';
    layer0_outputs(3167) <= '1';
    layer0_outputs(3168) <= (inputs(95)) and not (inputs(63));
    layer0_outputs(3169) <= (inputs(153)) and not (inputs(110));
    layer0_outputs(3170) <= not(inputs(165));
    layer0_outputs(3171) <= (inputs(230)) and not (inputs(123));
    layer0_outputs(3172) <= (inputs(29)) and not (inputs(206));
    layer0_outputs(3173) <= (inputs(35)) and not (inputs(233));
    layer0_outputs(3174) <= not(inputs(132));
    layer0_outputs(3175) <= not((inputs(220)) or (inputs(223)));
    layer0_outputs(3176) <= (inputs(26)) or (inputs(189));
    layer0_outputs(3177) <= inputs(147);
    layer0_outputs(3178) <= not(inputs(172));
    layer0_outputs(3179) <= '1';
    layer0_outputs(3180) <= (inputs(108)) xor (inputs(63));
    layer0_outputs(3181) <= not(inputs(79)) or (inputs(169));
    layer0_outputs(3182) <= inputs(230);
    layer0_outputs(3183) <= not(inputs(59)) or (inputs(192));
    layer0_outputs(3184) <= (inputs(145)) and not (inputs(171));
    layer0_outputs(3185) <= (inputs(194)) or (inputs(70));
    layer0_outputs(3186) <= not(inputs(228));
    layer0_outputs(3187) <= not((inputs(146)) and (inputs(1)));
    layer0_outputs(3188) <= (inputs(248)) or (inputs(138));
    layer0_outputs(3189) <= not(inputs(218)) or (inputs(249));
    layer0_outputs(3190) <= (inputs(51)) and not (inputs(24));
    layer0_outputs(3191) <= not((inputs(142)) or (inputs(109)));
    layer0_outputs(3192) <= inputs(50);
    layer0_outputs(3193) <= '1';
    layer0_outputs(3194) <= (inputs(160)) or (inputs(143));
    layer0_outputs(3195) <= (inputs(191)) and (inputs(120));
    layer0_outputs(3196) <= inputs(145);
    layer0_outputs(3197) <= (inputs(187)) or (inputs(31));
    layer0_outputs(3198) <= not((inputs(230)) xor (inputs(95)));
    layer0_outputs(3199) <= not(inputs(221)) or (inputs(34));
    layer0_outputs(3200) <= inputs(90);
    layer0_outputs(3201) <= not((inputs(135)) xor (inputs(248)));
    layer0_outputs(3202) <= inputs(179);
    layer0_outputs(3203) <= (inputs(8)) xor (inputs(52));
    layer0_outputs(3204) <= not(inputs(176));
    layer0_outputs(3205) <= inputs(15);
    layer0_outputs(3206) <= (inputs(35)) and not (inputs(227));
    layer0_outputs(3207) <= inputs(104);
    layer0_outputs(3208) <= (inputs(115)) or (inputs(40));
    layer0_outputs(3209) <= '1';
    layer0_outputs(3210) <= '0';
    layer0_outputs(3211) <= (inputs(152)) xor (inputs(30));
    layer0_outputs(3212) <= not(inputs(2)) or (inputs(91));
    layer0_outputs(3213) <= not((inputs(217)) and (inputs(56)));
    layer0_outputs(3214) <= (inputs(56)) and not (inputs(55));
    layer0_outputs(3215) <= (inputs(17)) and not (inputs(7));
    layer0_outputs(3216) <= (inputs(54)) and not (inputs(126));
    layer0_outputs(3217) <= not((inputs(113)) and (inputs(34)));
    layer0_outputs(3218) <= (inputs(183)) and not (inputs(67));
    layer0_outputs(3219) <= (inputs(213)) and not (inputs(76));
    layer0_outputs(3220) <= '0';
    layer0_outputs(3221) <= (inputs(252)) or (inputs(96));
    layer0_outputs(3222) <= not(inputs(146)) or (inputs(165));
    layer0_outputs(3223) <= (inputs(86)) and not (inputs(154));
    layer0_outputs(3224) <= inputs(196);
    layer0_outputs(3225) <= not(inputs(74));
    layer0_outputs(3226) <= (inputs(232)) or (inputs(101));
    layer0_outputs(3227) <= (inputs(61)) xor (inputs(51));
    layer0_outputs(3228) <= (inputs(37)) and not (inputs(157));
    layer0_outputs(3229) <= not((inputs(230)) xor (inputs(243)));
    layer0_outputs(3230) <= (inputs(102)) and not (inputs(103));
    layer0_outputs(3231) <= not((inputs(107)) xor (inputs(15)));
    layer0_outputs(3232) <= not((inputs(118)) or (inputs(189)));
    layer0_outputs(3233) <= inputs(12);
    layer0_outputs(3234) <= not((inputs(194)) xor (inputs(144)));
    layer0_outputs(3235) <= (inputs(213)) or (inputs(11));
    layer0_outputs(3236) <= not(inputs(220));
    layer0_outputs(3237) <= (inputs(178)) and not (inputs(200));
    layer0_outputs(3238) <= (inputs(72)) xor (inputs(245));
    layer0_outputs(3239) <= (inputs(197)) xor (inputs(161));
    layer0_outputs(3240) <= '1';
    layer0_outputs(3241) <= not((inputs(143)) or (inputs(97)));
    layer0_outputs(3242) <= inputs(148);
    layer0_outputs(3243) <= not(inputs(13)) or (inputs(36));
    layer0_outputs(3244) <= (inputs(151)) and not (inputs(64));
    layer0_outputs(3245) <= '0';
    layer0_outputs(3246) <= (inputs(179)) and not (inputs(231));
    layer0_outputs(3247) <= '1';
    layer0_outputs(3248) <= not((inputs(241)) xor (inputs(92)));
    layer0_outputs(3249) <= not((inputs(52)) xor (inputs(2)));
    layer0_outputs(3250) <= (inputs(164)) or (inputs(252));
    layer0_outputs(3251) <= not((inputs(1)) and (inputs(240)));
    layer0_outputs(3252) <= (inputs(233)) and (inputs(5));
    layer0_outputs(3253) <= (inputs(215)) or (inputs(251));
    layer0_outputs(3254) <= '1';
    layer0_outputs(3255) <= '0';
    layer0_outputs(3256) <= (inputs(147)) or (inputs(211));
    layer0_outputs(3257) <= not(inputs(216));
    layer0_outputs(3258) <= (inputs(42)) or (inputs(198));
    layer0_outputs(3259) <= '1';
    layer0_outputs(3260) <= not(inputs(165));
    layer0_outputs(3261) <= not(inputs(61));
    layer0_outputs(3262) <= inputs(133);
    layer0_outputs(3263) <= '0';
    layer0_outputs(3264) <= not(inputs(126));
    layer0_outputs(3265) <= '1';
    layer0_outputs(3266) <= not(inputs(120));
    layer0_outputs(3267) <= not(inputs(150));
    layer0_outputs(3268) <= (inputs(10)) xor (inputs(37));
    layer0_outputs(3269) <= not(inputs(143)) or (inputs(69));
    layer0_outputs(3270) <= not(inputs(246));
    layer0_outputs(3271) <= not((inputs(84)) xor (inputs(144)));
    layer0_outputs(3272) <= inputs(64);
    layer0_outputs(3273) <= not(inputs(51));
    layer0_outputs(3274) <= inputs(246);
    layer0_outputs(3275) <= (inputs(173)) xor (inputs(3));
    layer0_outputs(3276) <= inputs(106);
    layer0_outputs(3277) <= not(inputs(11));
    layer0_outputs(3278) <= not((inputs(105)) and (inputs(69)));
    layer0_outputs(3279) <= '1';
    layer0_outputs(3280) <= not(inputs(126)) or (inputs(68));
    layer0_outputs(3281) <= (inputs(23)) xor (inputs(209));
    layer0_outputs(3282) <= '0';
    layer0_outputs(3283) <= (inputs(5)) and not (inputs(129));
    layer0_outputs(3284) <= not((inputs(101)) or (inputs(60)));
    layer0_outputs(3285) <= not(inputs(133));
    layer0_outputs(3286) <= (inputs(81)) and (inputs(232));
    layer0_outputs(3287) <= not(inputs(86)) or (inputs(38));
    layer0_outputs(3288) <= (inputs(73)) and (inputs(87));
    layer0_outputs(3289) <= not((inputs(244)) xor (inputs(124)));
    layer0_outputs(3290) <= inputs(148);
    layer0_outputs(3291) <= not(inputs(149));
    layer0_outputs(3292) <= inputs(88);
    layer0_outputs(3293) <= not((inputs(140)) or (inputs(196)));
    layer0_outputs(3294) <= '0';
    layer0_outputs(3295) <= not((inputs(2)) or (inputs(147)));
    layer0_outputs(3296) <= (inputs(200)) and not (inputs(32));
    layer0_outputs(3297) <= not((inputs(234)) and (inputs(212)));
    layer0_outputs(3298) <= '0';
    layer0_outputs(3299) <= inputs(216);
    layer0_outputs(3300) <= not((inputs(188)) and (inputs(5)));
    layer0_outputs(3301) <= '0';
    layer0_outputs(3302) <= not((inputs(35)) xor (inputs(191)));
    layer0_outputs(3303) <= not((inputs(186)) xor (inputs(65)));
    layer0_outputs(3304) <= (inputs(164)) or (inputs(195));
    layer0_outputs(3305) <= inputs(133);
    layer0_outputs(3306) <= not((inputs(20)) xor (inputs(179)));
    layer0_outputs(3307) <= (inputs(225)) and not (inputs(193));
    layer0_outputs(3308) <= (inputs(28)) or (inputs(132));
    layer0_outputs(3309) <= not((inputs(100)) xor (inputs(136)));
    layer0_outputs(3310) <= not(inputs(122)) or (inputs(202));
    layer0_outputs(3311) <= not(inputs(228));
    layer0_outputs(3312) <= not((inputs(9)) and (inputs(70)));
    layer0_outputs(3313) <= (inputs(220)) and not (inputs(178));
    layer0_outputs(3314) <= '1';
    layer0_outputs(3315) <= inputs(116);
    layer0_outputs(3316) <= inputs(86);
    layer0_outputs(3317) <= inputs(200);
    layer0_outputs(3318) <= (inputs(193)) xor (inputs(18));
    layer0_outputs(3319) <= not(inputs(234));
    layer0_outputs(3320) <= not(inputs(221)) or (inputs(109));
    layer0_outputs(3321) <= (inputs(33)) xor (inputs(71));
    layer0_outputs(3322) <= '0';
    layer0_outputs(3323) <= (inputs(71)) and (inputs(193));
    layer0_outputs(3324) <= not(inputs(37)) or (inputs(228));
    layer0_outputs(3325) <= (inputs(79)) xor (inputs(2));
    layer0_outputs(3326) <= '1';
    layer0_outputs(3327) <= inputs(33);
    layer0_outputs(3328) <= (inputs(33)) and (inputs(193));
    layer0_outputs(3329) <= (inputs(218)) and (inputs(206));
    layer0_outputs(3330) <= (inputs(102)) or (inputs(6));
    layer0_outputs(3331) <= (inputs(160)) and not (inputs(247));
    layer0_outputs(3332) <= (inputs(192)) xor (inputs(126));
    layer0_outputs(3333) <= '0';
    layer0_outputs(3334) <= not((inputs(64)) or (inputs(142)));
    layer0_outputs(3335) <= not((inputs(210)) xor (inputs(204)));
    layer0_outputs(3336) <= inputs(153);
    layer0_outputs(3337) <= (inputs(244)) and not (inputs(82));
    layer0_outputs(3338) <= not(inputs(76));
    layer0_outputs(3339) <= not(inputs(79)) or (inputs(33));
    layer0_outputs(3340) <= inputs(46);
    layer0_outputs(3341) <= (inputs(56)) and not (inputs(150));
    layer0_outputs(3342) <= (inputs(223)) and not (inputs(25));
    layer0_outputs(3343) <= '0';
    layer0_outputs(3344) <= (inputs(161)) or (inputs(156));
    layer0_outputs(3345) <= not(inputs(136));
    layer0_outputs(3346) <= not(inputs(184));
    layer0_outputs(3347) <= not(inputs(45));
    layer0_outputs(3348) <= not((inputs(8)) and (inputs(111)));
    layer0_outputs(3349) <= (inputs(65)) and not (inputs(139));
    layer0_outputs(3350) <= (inputs(192)) or (inputs(137));
    layer0_outputs(3351) <= not(inputs(201)) or (inputs(61));
    layer0_outputs(3352) <= not(inputs(197));
    layer0_outputs(3353) <= not((inputs(9)) or (inputs(179)));
    layer0_outputs(3354) <= (inputs(208)) or (inputs(208));
    layer0_outputs(3355) <= (inputs(119)) and not (inputs(40));
    layer0_outputs(3356) <= '1';
    layer0_outputs(3357) <= (inputs(29)) and not (inputs(51));
    layer0_outputs(3358) <= inputs(224);
    layer0_outputs(3359) <= not(inputs(128));
    layer0_outputs(3360) <= inputs(64);
    layer0_outputs(3361) <= '1';
    layer0_outputs(3362) <= not((inputs(176)) and (inputs(221)));
    layer0_outputs(3363) <= '0';
    layer0_outputs(3364) <= not((inputs(223)) xor (inputs(113)));
    layer0_outputs(3365) <= (inputs(151)) and not (inputs(67));
    layer0_outputs(3366) <= not(inputs(200)) or (inputs(210));
    layer0_outputs(3367) <= '1';
    layer0_outputs(3368) <= not(inputs(76)) or (inputs(48));
    layer0_outputs(3369) <= not((inputs(206)) xor (inputs(139)));
    layer0_outputs(3370) <= '0';
    layer0_outputs(3371) <= inputs(90);
    layer0_outputs(3372) <= not((inputs(187)) and (inputs(74)));
    layer0_outputs(3373) <= inputs(251);
    layer0_outputs(3374) <= not(inputs(69));
    layer0_outputs(3375) <= not(inputs(40)) or (inputs(141));
    layer0_outputs(3376) <= '0';
    layer0_outputs(3377) <= not((inputs(160)) and (inputs(254)));
    layer0_outputs(3378) <= not((inputs(192)) and (inputs(121)));
    layer0_outputs(3379) <= (inputs(238)) and not (inputs(24));
    layer0_outputs(3380) <= (inputs(31)) and not (inputs(104));
    layer0_outputs(3381) <= inputs(150);
    layer0_outputs(3382) <= '1';
    layer0_outputs(3383) <= (inputs(195)) and not (inputs(103));
    layer0_outputs(3384) <= inputs(207);
    layer0_outputs(3385) <= not(inputs(182));
    layer0_outputs(3386) <= not((inputs(10)) xor (inputs(168)));
    layer0_outputs(3387) <= (inputs(179)) and not (inputs(12));
    layer0_outputs(3388) <= inputs(128);
    layer0_outputs(3389) <= not(inputs(237)) or (inputs(172));
    layer0_outputs(3390) <= inputs(203);
    layer0_outputs(3391) <= inputs(95);
    layer0_outputs(3392) <= not(inputs(133)) or (inputs(227));
    layer0_outputs(3393) <= not((inputs(183)) or (inputs(16)));
    layer0_outputs(3394) <= not(inputs(106));
    layer0_outputs(3395) <= (inputs(183)) and not (inputs(52));
    layer0_outputs(3396) <= not((inputs(198)) or (inputs(165)));
    layer0_outputs(3397) <= (inputs(140)) and not (inputs(174));
    layer0_outputs(3398) <= not(inputs(9)) or (inputs(223));
    layer0_outputs(3399) <= (inputs(176)) xor (inputs(44));
    layer0_outputs(3400) <= inputs(11);
    layer0_outputs(3401) <= not((inputs(59)) and (inputs(88)));
    layer0_outputs(3402) <= '1';
    layer0_outputs(3403) <= '1';
    layer0_outputs(3404) <= not((inputs(172)) or (inputs(241)));
    layer0_outputs(3405) <= not(inputs(16)) or (inputs(210));
    layer0_outputs(3406) <= (inputs(219)) and not (inputs(185));
    layer0_outputs(3407) <= (inputs(11)) xor (inputs(187));
    layer0_outputs(3408) <= (inputs(28)) and not (inputs(130));
    layer0_outputs(3409) <= not((inputs(123)) xor (inputs(140)));
    layer0_outputs(3410) <= (inputs(213)) xor (inputs(220));
    layer0_outputs(3411) <= not(inputs(97));
    layer0_outputs(3412) <= '0';
    layer0_outputs(3413) <= not(inputs(46));
    layer0_outputs(3414) <= not(inputs(45)) or (inputs(144));
    layer0_outputs(3415) <= (inputs(65)) and not (inputs(17));
    layer0_outputs(3416) <= inputs(81);
    layer0_outputs(3417) <= (inputs(235)) xor (inputs(19));
    layer0_outputs(3418) <= not((inputs(131)) or (inputs(108)));
    layer0_outputs(3419) <= inputs(59);
    layer0_outputs(3420) <= inputs(109);
    layer0_outputs(3421) <= (inputs(210)) and not (inputs(192));
    layer0_outputs(3422) <= not(inputs(135)) or (inputs(88));
    layer0_outputs(3423) <= not((inputs(113)) xor (inputs(229)));
    layer0_outputs(3424) <= '0';
    layer0_outputs(3425) <= not(inputs(254)) or (inputs(250));
    layer0_outputs(3426) <= not(inputs(130));
    layer0_outputs(3427) <= (inputs(44)) and not (inputs(246));
    layer0_outputs(3428) <= (inputs(58)) and (inputs(239));
    layer0_outputs(3429) <= (inputs(133)) or (inputs(217));
    layer0_outputs(3430) <= not(inputs(16));
    layer0_outputs(3431) <= not((inputs(191)) and (inputs(118)));
    layer0_outputs(3432) <= (inputs(45)) or (inputs(154));
    layer0_outputs(3433) <= not((inputs(156)) or (inputs(254)));
    layer0_outputs(3434) <= (inputs(229)) and not (inputs(235));
    layer0_outputs(3435) <= (inputs(41)) or (inputs(133));
    layer0_outputs(3436) <= not(inputs(47)) or (inputs(85));
    layer0_outputs(3437) <= not((inputs(79)) or (inputs(53)));
    layer0_outputs(3438) <= (inputs(93)) xor (inputs(187));
    layer0_outputs(3439) <= (inputs(144)) or (inputs(139));
    layer0_outputs(3440) <= (inputs(41)) or (inputs(147));
    layer0_outputs(3441) <= inputs(105);
    layer0_outputs(3442) <= (inputs(163)) and not (inputs(64));
    layer0_outputs(3443) <= not(inputs(67)) or (inputs(244));
    layer0_outputs(3444) <= '0';
    layer0_outputs(3445) <= (inputs(198)) or (inputs(195));
    layer0_outputs(3446) <= (inputs(108)) or (inputs(165));
    layer0_outputs(3447) <= (inputs(99)) and not (inputs(207));
    layer0_outputs(3448) <= not((inputs(39)) xor (inputs(22)));
    layer0_outputs(3449) <= inputs(191);
    layer0_outputs(3450) <= not((inputs(142)) or (inputs(148)));
    layer0_outputs(3451) <= not((inputs(249)) or (inputs(140)));
    layer0_outputs(3452) <= not(inputs(55)) or (inputs(228));
    layer0_outputs(3453) <= (inputs(68)) xor (inputs(133));
    layer0_outputs(3454) <= not((inputs(245)) and (inputs(9)));
    layer0_outputs(3455) <= inputs(226);
    layer0_outputs(3456) <= (inputs(243)) and not (inputs(239));
    layer0_outputs(3457) <= inputs(67);
    layer0_outputs(3458) <= (inputs(80)) and not (inputs(123));
    layer0_outputs(3459) <= (inputs(198)) and not (inputs(65));
    layer0_outputs(3460) <= not((inputs(44)) or (inputs(119)));
    layer0_outputs(3461) <= not(inputs(26)) or (inputs(202));
    layer0_outputs(3462) <= (inputs(122)) or (inputs(48));
    layer0_outputs(3463) <= inputs(200);
    layer0_outputs(3464) <= (inputs(144)) and (inputs(69));
    layer0_outputs(3465) <= '1';
    layer0_outputs(3466) <= (inputs(178)) and (inputs(127));
    layer0_outputs(3467) <= not((inputs(157)) xor (inputs(204)));
    layer0_outputs(3468) <= (inputs(108)) and not (inputs(43));
    layer0_outputs(3469) <= inputs(30);
    layer0_outputs(3470) <= not(inputs(128)) or (inputs(74));
    layer0_outputs(3471) <= '1';
    layer0_outputs(3472) <= (inputs(133)) xor (inputs(221));
    layer0_outputs(3473) <= (inputs(28)) and not (inputs(235));
    layer0_outputs(3474) <= '0';
    layer0_outputs(3475) <= (inputs(51)) or (inputs(196));
    layer0_outputs(3476) <= inputs(20);
    layer0_outputs(3477) <= inputs(180);
    layer0_outputs(3478) <= inputs(154);
    layer0_outputs(3479) <= (inputs(5)) and (inputs(145));
    layer0_outputs(3480) <= '0';
    layer0_outputs(3481) <= (inputs(220)) xor (inputs(212));
    layer0_outputs(3482) <= (inputs(13)) and not (inputs(168));
    layer0_outputs(3483) <= (inputs(140)) and not (inputs(170));
    layer0_outputs(3484) <= (inputs(151)) and not (inputs(228));
    layer0_outputs(3485) <= (inputs(251)) or (inputs(234));
    layer0_outputs(3486) <= not(inputs(14));
    layer0_outputs(3487) <= (inputs(6)) and (inputs(93));
    layer0_outputs(3488) <= (inputs(238)) and not (inputs(97));
    layer0_outputs(3489) <= not(inputs(0)) or (inputs(27));
    layer0_outputs(3490) <= not((inputs(1)) or (inputs(162)));
    layer0_outputs(3491) <= not((inputs(196)) or (inputs(174)));
    layer0_outputs(3492) <= (inputs(59)) and not (inputs(48));
    layer0_outputs(3493) <= not(inputs(213));
    layer0_outputs(3494) <= not(inputs(162)) or (inputs(28));
    layer0_outputs(3495) <= not((inputs(76)) and (inputs(76)));
    layer0_outputs(3496) <= not(inputs(136)) or (inputs(144));
    layer0_outputs(3497) <= not(inputs(182)) or (inputs(75));
    layer0_outputs(3498) <= '0';
    layer0_outputs(3499) <= not((inputs(68)) xor (inputs(204)));
    layer0_outputs(3500) <= (inputs(125)) or (inputs(80));
    layer0_outputs(3501) <= inputs(219);
    layer0_outputs(3502) <= inputs(128);
    layer0_outputs(3503) <= '1';
    layer0_outputs(3504) <= inputs(102);
    layer0_outputs(3505) <= not(inputs(35)) or (inputs(227));
    layer0_outputs(3506) <= '0';
    layer0_outputs(3507) <= not((inputs(177)) and (inputs(188)));
    layer0_outputs(3508) <= not(inputs(106));
    layer0_outputs(3509) <= not(inputs(215));
    layer0_outputs(3510) <= not(inputs(196)) or (inputs(161));
    layer0_outputs(3511) <= not(inputs(236)) or (inputs(115));
    layer0_outputs(3512) <= (inputs(48)) or (inputs(38));
    layer0_outputs(3513) <= not((inputs(161)) xor (inputs(198)));
    layer0_outputs(3514) <= not((inputs(109)) or (inputs(213)));
    layer0_outputs(3515) <= inputs(76);
    layer0_outputs(3516) <= inputs(53);
    layer0_outputs(3517) <= inputs(222);
    layer0_outputs(3518) <= (inputs(141)) and not (inputs(91));
    layer0_outputs(3519) <= (inputs(129)) and (inputs(101));
    layer0_outputs(3520) <= (inputs(221)) and not (inputs(33));
    layer0_outputs(3521) <= not(inputs(156));
    layer0_outputs(3522) <= (inputs(206)) or (inputs(163));
    layer0_outputs(3523) <= (inputs(235)) xor (inputs(36));
    layer0_outputs(3524) <= inputs(99);
    layer0_outputs(3525) <= '1';
    layer0_outputs(3526) <= not(inputs(121));
    layer0_outputs(3527) <= (inputs(36)) xor (inputs(215));
    layer0_outputs(3528) <= not(inputs(93)) or (inputs(168));
    layer0_outputs(3529) <= '0';
    layer0_outputs(3530) <= (inputs(161)) or (inputs(37));
    layer0_outputs(3531) <= inputs(57);
    layer0_outputs(3532) <= (inputs(196)) and not (inputs(108));
    layer0_outputs(3533) <= '1';
    layer0_outputs(3534) <= not((inputs(228)) and (inputs(8)));
    layer0_outputs(3535) <= not((inputs(63)) or (inputs(198)));
    layer0_outputs(3536) <= not(inputs(143)) or (inputs(223));
    layer0_outputs(3537) <= (inputs(175)) or (inputs(124));
    layer0_outputs(3538) <= inputs(165);
    layer0_outputs(3539) <= not(inputs(104));
    layer0_outputs(3540) <= not((inputs(30)) or (inputs(107)));
    layer0_outputs(3541) <= not(inputs(9));
    layer0_outputs(3542) <= (inputs(185)) or (inputs(70));
    layer0_outputs(3543) <= inputs(59);
    layer0_outputs(3544) <= not((inputs(175)) or (inputs(3)));
    layer0_outputs(3545) <= not((inputs(73)) xor (inputs(250)));
    layer0_outputs(3546) <= (inputs(202)) or (inputs(20));
    layer0_outputs(3547) <= inputs(235);
    layer0_outputs(3548) <= not(inputs(112));
    layer0_outputs(3549) <= (inputs(112)) and not (inputs(116));
    layer0_outputs(3550) <= (inputs(153)) or (inputs(0));
    layer0_outputs(3551) <= inputs(66);
    layer0_outputs(3552) <= (inputs(252)) or (inputs(19));
    layer0_outputs(3553) <= inputs(180);
    layer0_outputs(3554) <= not((inputs(21)) xor (inputs(206)));
    layer0_outputs(3555) <= (inputs(202)) and not (inputs(21));
    layer0_outputs(3556) <= not(inputs(218));
    layer0_outputs(3557) <= not((inputs(48)) or (inputs(116)));
    layer0_outputs(3558) <= not(inputs(213));
    layer0_outputs(3559) <= not(inputs(12));
    layer0_outputs(3560) <= not((inputs(57)) xor (inputs(158)));
    layer0_outputs(3561) <= (inputs(204)) or (inputs(192));
    layer0_outputs(3562) <= '0';
    layer0_outputs(3563) <= not(inputs(102));
    layer0_outputs(3564) <= not((inputs(180)) xor (inputs(32)));
    layer0_outputs(3565) <= (inputs(242)) or (inputs(175));
    layer0_outputs(3566) <= inputs(186);
    layer0_outputs(3567) <= not(inputs(219)) or (inputs(30));
    layer0_outputs(3568) <= not((inputs(54)) xor (inputs(111)));
    layer0_outputs(3569) <= '1';
    layer0_outputs(3570) <= (inputs(5)) and not (inputs(30));
    layer0_outputs(3571) <= (inputs(237)) and (inputs(20));
    layer0_outputs(3572) <= not((inputs(142)) and (inputs(181)));
    layer0_outputs(3573) <= not((inputs(171)) xor (inputs(188)));
    layer0_outputs(3574) <= not((inputs(15)) xor (inputs(104)));
    layer0_outputs(3575) <= not(inputs(113));
    layer0_outputs(3576) <= (inputs(89)) and not (inputs(164));
    layer0_outputs(3577) <= (inputs(143)) or (inputs(56));
    layer0_outputs(3578) <= not(inputs(235));
    layer0_outputs(3579) <= not((inputs(78)) or (inputs(88)));
    layer0_outputs(3580) <= inputs(152);
    layer0_outputs(3581) <= not(inputs(30));
    layer0_outputs(3582) <= (inputs(200)) xor (inputs(47));
    layer0_outputs(3583) <= not((inputs(234)) or (inputs(98)));
    layer0_outputs(3584) <= not(inputs(6)) or (inputs(95));
    layer0_outputs(3585) <= not(inputs(237)) or (inputs(233));
    layer0_outputs(3586) <= not(inputs(202));
    layer0_outputs(3587) <= not((inputs(211)) or (inputs(69)));
    layer0_outputs(3588) <= (inputs(34)) or (inputs(90));
    layer0_outputs(3589) <= not(inputs(203));
    layer0_outputs(3590) <= not((inputs(178)) or (inputs(72)));
    layer0_outputs(3591) <= not(inputs(201));
    layer0_outputs(3592) <= not(inputs(106)) or (inputs(224));
    layer0_outputs(3593) <= not((inputs(218)) and (inputs(78)));
    layer0_outputs(3594) <= not((inputs(152)) or (inputs(108)));
    layer0_outputs(3595) <= (inputs(185)) and not (inputs(34));
    layer0_outputs(3596) <= (inputs(251)) and not (inputs(141));
    layer0_outputs(3597) <= (inputs(203)) or (inputs(52));
    layer0_outputs(3598) <= (inputs(204)) and not (inputs(112));
    layer0_outputs(3599) <= (inputs(135)) and not (inputs(79));
    layer0_outputs(3600) <= '1';
    layer0_outputs(3601) <= (inputs(137)) and not (inputs(95));
    layer0_outputs(3602) <= (inputs(75)) or (inputs(211));
    layer0_outputs(3603) <= (inputs(59)) and not (inputs(177));
    layer0_outputs(3604) <= not((inputs(68)) xor (inputs(126)));
    layer0_outputs(3605) <= not((inputs(205)) or (inputs(52)));
    layer0_outputs(3606) <= (inputs(190)) or (inputs(4));
    layer0_outputs(3607) <= not((inputs(248)) and (inputs(37)));
    layer0_outputs(3608) <= not(inputs(183));
    layer0_outputs(3609) <= not(inputs(46));
    layer0_outputs(3610) <= (inputs(189)) or (inputs(164));
    layer0_outputs(3611) <= (inputs(36)) and (inputs(129));
    layer0_outputs(3612) <= (inputs(122)) and not (inputs(158));
    layer0_outputs(3613) <= not((inputs(186)) or (inputs(41)));
    layer0_outputs(3614) <= '0';
    layer0_outputs(3615) <= (inputs(135)) or (inputs(52));
    layer0_outputs(3616) <= '1';
    layer0_outputs(3617) <= not((inputs(173)) xor (inputs(63)));
    layer0_outputs(3618) <= not((inputs(166)) xor (inputs(2)));
    layer0_outputs(3619) <= not((inputs(14)) or (inputs(76)));
    layer0_outputs(3620) <= '0';
    layer0_outputs(3621) <= not(inputs(199)) or (inputs(11));
    layer0_outputs(3622) <= inputs(69);
    layer0_outputs(3623) <= not(inputs(133)) or (inputs(5));
    layer0_outputs(3624) <= not(inputs(160)) or (inputs(250));
    layer0_outputs(3625) <= (inputs(71)) or (inputs(233));
    layer0_outputs(3626) <= (inputs(142)) or (inputs(165));
    layer0_outputs(3627) <= not((inputs(10)) xor (inputs(90)));
    layer0_outputs(3628) <= not(inputs(124));
    layer0_outputs(3629) <= not(inputs(52));
    layer0_outputs(3630) <= not((inputs(236)) and (inputs(0)));
    layer0_outputs(3631) <= (inputs(192)) xor (inputs(245));
    layer0_outputs(3632) <= not(inputs(151));
    layer0_outputs(3633) <= inputs(196);
    layer0_outputs(3634) <= inputs(94);
    layer0_outputs(3635) <= inputs(102);
    layer0_outputs(3636) <= (inputs(95)) and (inputs(107));
    layer0_outputs(3637) <= (inputs(18)) and (inputs(160));
    layer0_outputs(3638) <= (inputs(201)) and (inputs(24));
    layer0_outputs(3639) <= not(inputs(227)) or (inputs(96));
    layer0_outputs(3640) <= not((inputs(118)) or (inputs(100)));
    layer0_outputs(3641) <= (inputs(158)) and (inputs(174));
    layer0_outputs(3642) <= inputs(147);
    layer0_outputs(3643) <= inputs(190);
    layer0_outputs(3644) <= (inputs(50)) and (inputs(96));
    layer0_outputs(3645) <= (inputs(2)) xor (inputs(188));
    layer0_outputs(3646) <= (inputs(201)) or (inputs(161));
    layer0_outputs(3647) <= not(inputs(33));
    layer0_outputs(3648) <= (inputs(23)) and (inputs(225));
    layer0_outputs(3649) <= not((inputs(103)) or (inputs(86)));
    layer0_outputs(3650) <= not(inputs(73));
    layer0_outputs(3651) <= not((inputs(95)) xor (inputs(232)));
    layer0_outputs(3652) <= inputs(108);
    layer0_outputs(3653) <= (inputs(202)) and not (inputs(19));
    layer0_outputs(3654) <= not(inputs(46));
    layer0_outputs(3655) <= not((inputs(36)) xor (inputs(120)));
    layer0_outputs(3656) <= '0';
    layer0_outputs(3657) <= '1';
    layer0_outputs(3658) <= not(inputs(197)) or (inputs(127));
    layer0_outputs(3659) <= (inputs(127)) and not (inputs(125));
    layer0_outputs(3660) <= not(inputs(138));
    layer0_outputs(3661) <= '1';
    layer0_outputs(3662) <= not(inputs(100));
    layer0_outputs(3663) <= inputs(76);
    layer0_outputs(3664) <= (inputs(42)) or (inputs(25));
    layer0_outputs(3665) <= (inputs(30)) xor (inputs(109));
    layer0_outputs(3666) <= inputs(177);
    layer0_outputs(3667) <= (inputs(229)) and (inputs(2));
    layer0_outputs(3668) <= (inputs(79)) or (inputs(55));
    layer0_outputs(3669) <= '0';
    layer0_outputs(3670) <= not(inputs(152));
    layer0_outputs(3671) <= '0';
    layer0_outputs(3672) <= not((inputs(81)) xor (inputs(51)));
    layer0_outputs(3673) <= not((inputs(82)) and (inputs(130)));
    layer0_outputs(3674) <= not((inputs(234)) xor (inputs(195)));
    layer0_outputs(3675) <= not(inputs(111)) or (inputs(53));
    layer0_outputs(3676) <= not(inputs(60));
    layer0_outputs(3677) <= not((inputs(145)) and (inputs(25)));
    layer0_outputs(3678) <= not(inputs(79)) or (inputs(59));
    layer0_outputs(3679) <= not(inputs(148)) or (inputs(221));
    layer0_outputs(3680) <= not((inputs(251)) and (inputs(119)));
    layer0_outputs(3681) <= not((inputs(166)) xor (inputs(0)));
    layer0_outputs(3682) <= not(inputs(48));
    layer0_outputs(3683) <= not((inputs(7)) or (inputs(223)));
    layer0_outputs(3684) <= '1';
    layer0_outputs(3685) <= (inputs(115)) and not (inputs(161));
    layer0_outputs(3686) <= not(inputs(29));
    layer0_outputs(3687) <= inputs(152);
    layer0_outputs(3688) <= not(inputs(10)) or (inputs(213));
    layer0_outputs(3689) <= (inputs(90)) or (inputs(171));
    layer0_outputs(3690) <= not(inputs(202));
    layer0_outputs(3691) <= (inputs(175)) xor (inputs(152));
    layer0_outputs(3692) <= (inputs(22)) and not (inputs(227));
    layer0_outputs(3693) <= inputs(197);
    layer0_outputs(3694) <= inputs(21);
    layer0_outputs(3695) <= not(inputs(93));
    layer0_outputs(3696) <= (inputs(253)) and not (inputs(55));
    layer0_outputs(3697) <= not(inputs(213));
    layer0_outputs(3698) <= not((inputs(141)) xor (inputs(28)));
    layer0_outputs(3699) <= not(inputs(164));
    layer0_outputs(3700) <= not(inputs(143)) or (inputs(6));
    layer0_outputs(3701) <= (inputs(136)) and not (inputs(172));
    layer0_outputs(3702) <= (inputs(165)) xor (inputs(1));
    layer0_outputs(3703) <= not(inputs(65));
    layer0_outputs(3704) <= not((inputs(163)) or (inputs(214)));
    layer0_outputs(3705) <= not((inputs(13)) or (inputs(62)));
    layer0_outputs(3706) <= '0';
    layer0_outputs(3707) <= not(inputs(128));
    layer0_outputs(3708) <= (inputs(185)) or (inputs(37));
    layer0_outputs(3709) <= not(inputs(120)) or (inputs(81));
    layer0_outputs(3710) <= not(inputs(241)) or (inputs(52));
    layer0_outputs(3711) <= inputs(53);
    layer0_outputs(3712) <= '0';
    layer0_outputs(3713) <= not(inputs(178)) or (inputs(175));
    layer0_outputs(3714) <= (inputs(75)) and not (inputs(222));
    layer0_outputs(3715) <= (inputs(178)) or (inputs(179));
    layer0_outputs(3716) <= not((inputs(62)) or (inputs(180)));
    layer0_outputs(3717) <= (inputs(12)) and not (inputs(211));
    layer0_outputs(3718) <= (inputs(162)) and not (inputs(232));
    layer0_outputs(3719) <= '0';
    layer0_outputs(3720) <= (inputs(108)) and (inputs(179));
    layer0_outputs(3721) <= (inputs(160)) or (inputs(18));
    layer0_outputs(3722) <= inputs(235);
    layer0_outputs(3723) <= '0';
    layer0_outputs(3724) <= (inputs(186)) and not (inputs(221));
    layer0_outputs(3725) <= inputs(224);
    layer0_outputs(3726) <= not(inputs(93));
    layer0_outputs(3727) <= not((inputs(236)) and (inputs(74)));
    layer0_outputs(3728) <= (inputs(46)) or (inputs(55));
    layer0_outputs(3729) <= not(inputs(116)) or (inputs(37));
    layer0_outputs(3730) <= inputs(199);
    layer0_outputs(3731) <= '0';
    layer0_outputs(3732) <= (inputs(215)) and not (inputs(142));
    layer0_outputs(3733) <= (inputs(183)) and not (inputs(184));
    layer0_outputs(3734) <= '0';
    layer0_outputs(3735) <= not((inputs(28)) xor (inputs(247)));
    layer0_outputs(3736) <= not((inputs(142)) or (inputs(100)));
    layer0_outputs(3737) <= '1';
    layer0_outputs(3738) <= (inputs(126)) and (inputs(91));
    layer0_outputs(3739) <= (inputs(160)) and not (inputs(255));
    layer0_outputs(3740) <= (inputs(10)) or (inputs(215));
    layer0_outputs(3741) <= (inputs(186)) or (inputs(4));
    layer0_outputs(3742) <= '1';
    layer0_outputs(3743) <= not((inputs(108)) or (inputs(239)));
    layer0_outputs(3744) <= not((inputs(6)) or (inputs(251)));
    layer0_outputs(3745) <= not((inputs(105)) or (inputs(98)));
    layer0_outputs(3746) <= not(inputs(2)) or (inputs(238));
    layer0_outputs(3747) <= not((inputs(170)) or (inputs(10)));
    layer0_outputs(3748) <= (inputs(150)) or (inputs(37));
    layer0_outputs(3749) <= not(inputs(170));
    layer0_outputs(3750) <= '0';
    layer0_outputs(3751) <= inputs(178);
    layer0_outputs(3752) <= (inputs(235)) or (inputs(248));
    layer0_outputs(3753) <= not((inputs(132)) xor (inputs(28)));
    layer0_outputs(3754) <= not(inputs(162)) or (inputs(150));
    layer0_outputs(3755) <= inputs(100);
    layer0_outputs(3756) <= not((inputs(235)) or (inputs(191)));
    layer0_outputs(3757) <= not((inputs(38)) or (inputs(181)));
    layer0_outputs(3758) <= not((inputs(203)) or (inputs(91)));
    layer0_outputs(3759) <= inputs(5);
    layer0_outputs(3760) <= not(inputs(48));
    layer0_outputs(3761) <= not((inputs(40)) xor (inputs(86)));
    layer0_outputs(3762) <= not((inputs(144)) xor (inputs(197)));
    layer0_outputs(3763) <= not(inputs(35)) or (inputs(207));
    layer0_outputs(3764) <= not(inputs(48)) or (inputs(243));
    layer0_outputs(3765) <= inputs(115);
    layer0_outputs(3766) <= not((inputs(100)) xor (inputs(232)));
    layer0_outputs(3767) <= not(inputs(168)) or (inputs(158));
    layer0_outputs(3768) <= not(inputs(203)) or (inputs(187));
    layer0_outputs(3769) <= not(inputs(247)) or (inputs(120));
    layer0_outputs(3770) <= (inputs(140)) or (inputs(41));
    layer0_outputs(3771) <= inputs(253);
    layer0_outputs(3772) <= not((inputs(83)) and (inputs(57)));
    layer0_outputs(3773) <= '1';
    layer0_outputs(3774) <= not(inputs(120)) or (inputs(162));
    layer0_outputs(3775) <= (inputs(168)) xor (inputs(159));
    layer0_outputs(3776) <= not(inputs(202));
    layer0_outputs(3777) <= not(inputs(156)) or (inputs(2));
    layer0_outputs(3778) <= inputs(138);
    layer0_outputs(3779) <= (inputs(48)) and not (inputs(206));
    layer0_outputs(3780) <= '0';
    layer0_outputs(3781) <= inputs(132);
    layer0_outputs(3782) <= not(inputs(171)) or (inputs(130));
    layer0_outputs(3783) <= (inputs(80)) or (inputs(250));
    layer0_outputs(3784) <= (inputs(26)) or (inputs(248));
    layer0_outputs(3785) <= not((inputs(120)) and (inputs(58)));
    layer0_outputs(3786) <= (inputs(105)) xor (inputs(46));
    layer0_outputs(3787) <= (inputs(133)) and not (inputs(92));
    layer0_outputs(3788) <= not((inputs(169)) or (inputs(67)));
    layer0_outputs(3789) <= not(inputs(46));
    layer0_outputs(3790) <= inputs(78);
    layer0_outputs(3791) <= (inputs(170)) and not (inputs(228));
    layer0_outputs(3792) <= inputs(195);
    layer0_outputs(3793) <= (inputs(109)) or (inputs(116));
    layer0_outputs(3794) <= (inputs(204)) and not (inputs(99));
    layer0_outputs(3795) <= inputs(250);
    layer0_outputs(3796) <= '1';
    layer0_outputs(3797) <= not((inputs(4)) and (inputs(180)));
    layer0_outputs(3798) <= inputs(101);
    layer0_outputs(3799) <= inputs(87);
    layer0_outputs(3800) <= (inputs(126)) or (inputs(125));
    layer0_outputs(3801) <= (inputs(163)) and not (inputs(6));
    layer0_outputs(3802) <= inputs(131);
    layer0_outputs(3803) <= not((inputs(15)) or (inputs(215)));
    layer0_outputs(3804) <= not((inputs(55)) or (inputs(240)));
    layer0_outputs(3805) <= inputs(153);
    layer0_outputs(3806) <= (inputs(119)) and (inputs(71));
    layer0_outputs(3807) <= (inputs(157)) and not (inputs(63));
    layer0_outputs(3808) <= (inputs(240)) and not (inputs(144));
    layer0_outputs(3809) <= not(inputs(129)) or (inputs(141));
    layer0_outputs(3810) <= '1';
    layer0_outputs(3811) <= inputs(164);
    layer0_outputs(3812) <= '1';
    layer0_outputs(3813) <= '1';
    layer0_outputs(3814) <= not(inputs(100));
    layer0_outputs(3815) <= (inputs(101)) or (inputs(8));
    layer0_outputs(3816) <= (inputs(11)) and not (inputs(58));
    layer0_outputs(3817) <= not((inputs(22)) and (inputs(131)));
    layer0_outputs(3818) <= not(inputs(188)) or (inputs(198));
    layer0_outputs(3819) <= (inputs(71)) or (inputs(181));
    layer0_outputs(3820) <= (inputs(58)) and not (inputs(250));
    layer0_outputs(3821) <= (inputs(206)) and not (inputs(206));
    layer0_outputs(3822) <= not((inputs(227)) xor (inputs(182)));
    layer0_outputs(3823) <= not(inputs(121));
    layer0_outputs(3824) <= not(inputs(209));
    layer0_outputs(3825) <= not(inputs(187)) or (inputs(77));
    layer0_outputs(3826) <= (inputs(203)) and (inputs(162));
    layer0_outputs(3827) <= (inputs(183)) and not (inputs(32));
    layer0_outputs(3828) <= inputs(30);
    layer0_outputs(3829) <= '1';
    layer0_outputs(3830) <= (inputs(36)) or (inputs(195));
    layer0_outputs(3831) <= inputs(11);
    layer0_outputs(3832) <= not((inputs(101)) or (inputs(219)));
    layer0_outputs(3833) <= (inputs(43)) xor (inputs(159));
    layer0_outputs(3834) <= not(inputs(32)) or (inputs(220));
    layer0_outputs(3835) <= not(inputs(43)) or (inputs(39));
    layer0_outputs(3836) <= inputs(117);
    layer0_outputs(3837) <= (inputs(164)) or (inputs(110));
    layer0_outputs(3838) <= inputs(31);
    layer0_outputs(3839) <= '0';
    layer0_outputs(3840) <= not(inputs(91)) or (inputs(23));
    layer0_outputs(3841) <= not(inputs(1)) or (inputs(216));
    layer0_outputs(3842) <= (inputs(237)) xor (inputs(125));
    layer0_outputs(3843) <= not(inputs(132));
    layer0_outputs(3844) <= (inputs(118)) and not (inputs(2));
    layer0_outputs(3845) <= not(inputs(45));
    layer0_outputs(3846) <= (inputs(149)) and (inputs(186));
    layer0_outputs(3847) <= (inputs(88)) and not (inputs(9));
    layer0_outputs(3848) <= not(inputs(105));
    layer0_outputs(3849) <= (inputs(33)) and not (inputs(8));
    layer0_outputs(3850) <= (inputs(2)) and (inputs(253));
    layer0_outputs(3851) <= (inputs(53)) or (inputs(8));
    layer0_outputs(3852) <= not(inputs(24)) or (inputs(101));
    layer0_outputs(3853) <= not((inputs(244)) and (inputs(74)));
    layer0_outputs(3854) <= (inputs(51)) and not (inputs(193));
    layer0_outputs(3855) <= (inputs(36)) or (inputs(22));
    layer0_outputs(3856) <= not(inputs(24));
    layer0_outputs(3857) <= not((inputs(218)) xor (inputs(186)));
    layer0_outputs(3858) <= inputs(159);
    layer0_outputs(3859) <= (inputs(124)) and not (inputs(48));
    layer0_outputs(3860) <= (inputs(137)) and not (inputs(3));
    layer0_outputs(3861) <= (inputs(215)) and not (inputs(242));
    layer0_outputs(3862) <= not(inputs(238)) or (inputs(10));
    layer0_outputs(3863) <= '1';
    layer0_outputs(3864) <= (inputs(158)) and not (inputs(28));
    layer0_outputs(3865) <= not(inputs(126));
    layer0_outputs(3866) <= inputs(30);
    layer0_outputs(3867) <= (inputs(157)) or (inputs(129));
    layer0_outputs(3868) <= not(inputs(12)) or (inputs(77));
    layer0_outputs(3869) <= (inputs(76)) xor (inputs(5));
    layer0_outputs(3870) <= '0';
    layer0_outputs(3871) <= (inputs(92)) and (inputs(18));
    layer0_outputs(3872) <= not(inputs(78)) or (inputs(228));
    layer0_outputs(3873) <= (inputs(118)) or (inputs(200));
    layer0_outputs(3874) <= inputs(85);
    layer0_outputs(3875) <= '1';
    layer0_outputs(3876) <= not((inputs(144)) or (inputs(121)));
    layer0_outputs(3877) <= not((inputs(144)) or (inputs(110)));
    layer0_outputs(3878) <= (inputs(30)) xor (inputs(55));
    layer0_outputs(3879) <= (inputs(114)) or (inputs(101));
    layer0_outputs(3880) <= not(inputs(56)) or (inputs(29));
    layer0_outputs(3881) <= not(inputs(102)) or (inputs(238));
    layer0_outputs(3882) <= (inputs(117)) and not (inputs(153));
    layer0_outputs(3883) <= (inputs(249)) or (inputs(22));
    layer0_outputs(3884) <= '0';
    layer0_outputs(3885) <= (inputs(198)) or (inputs(204));
    layer0_outputs(3886) <= not((inputs(118)) xor (inputs(147)));
    layer0_outputs(3887) <= '0';
    layer0_outputs(3888) <= (inputs(186)) or (inputs(129));
    layer0_outputs(3889) <= not(inputs(40)) or (inputs(0));
    layer0_outputs(3890) <= (inputs(180)) and not (inputs(212));
    layer0_outputs(3891) <= (inputs(10)) or (inputs(113));
    layer0_outputs(3892) <= not(inputs(185));
    layer0_outputs(3893) <= not(inputs(158));
    layer0_outputs(3894) <= not((inputs(212)) or (inputs(153)));
    layer0_outputs(3895) <= inputs(85);
    layer0_outputs(3896) <= not(inputs(90)) or (inputs(157));
    layer0_outputs(3897) <= not((inputs(221)) xor (inputs(194)));
    layer0_outputs(3898) <= inputs(71);
    layer0_outputs(3899) <= inputs(15);
    layer0_outputs(3900) <= (inputs(243)) and (inputs(29));
    layer0_outputs(3901) <= not(inputs(175)) or (inputs(128));
    layer0_outputs(3902) <= not((inputs(37)) or (inputs(227)));
    layer0_outputs(3903) <= not((inputs(204)) or (inputs(249)));
    layer0_outputs(3904) <= (inputs(142)) and not (inputs(137));
    layer0_outputs(3905) <= not(inputs(42)) or (inputs(104));
    layer0_outputs(3906) <= '1';
    layer0_outputs(3907) <= (inputs(11)) xor (inputs(20));
    layer0_outputs(3908) <= not(inputs(213)) or (inputs(24));
    layer0_outputs(3909) <= not((inputs(115)) and (inputs(131)));
    layer0_outputs(3910) <= not(inputs(104)) or (inputs(22));
    layer0_outputs(3911) <= not((inputs(58)) xor (inputs(3)));
    layer0_outputs(3912) <= not((inputs(152)) or (inputs(30)));
    layer0_outputs(3913) <= (inputs(226)) and not (inputs(205));
    layer0_outputs(3914) <= not((inputs(26)) xor (inputs(92)));
    layer0_outputs(3915) <= (inputs(161)) and not (inputs(213));
    layer0_outputs(3916) <= not(inputs(218)) or (inputs(212));
    layer0_outputs(3917) <= (inputs(231)) and (inputs(157));
    layer0_outputs(3918) <= not(inputs(137)) or (inputs(217));
    layer0_outputs(3919) <= not(inputs(92)) or (inputs(68));
    layer0_outputs(3920) <= '0';
    layer0_outputs(3921) <= (inputs(58)) and not (inputs(44));
    layer0_outputs(3922) <= (inputs(130)) and not (inputs(48));
    layer0_outputs(3923) <= not((inputs(108)) or (inputs(75)));
    layer0_outputs(3924) <= '1';
    layer0_outputs(3925) <= not((inputs(174)) and (inputs(29)));
    layer0_outputs(3926) <= inputs(147);
    layer0_outputs(3927) <= '1';
    layer0_outputs(3928) <= (inputs(197)) or (inputs(158));
    layer0_outputs(3929) <= inputs(42);
    layer0_outputs(3930) <= '1';
    layer0_outputs(3931) <= not(inputs(77));
    layer0_outputs(3932) <= '1';
    layer0_outputs(3933) <= inputs(180);
    layer0_outputs(3934) <= not(inputs(134));
    layer0_outputs(3935) <= '0';
    layer0_outputs(3936) <= not((inputs(233)) and (inputs(37)));
    layer0_outputs(3937) <= not((inputs(239)) xor (inputs(153)));
    layer0_outputs(3938) <= not(inputs(100)) or (inputs(94));
    layer0_outputs(3939) <= inputs(68);
    layer0_outputs(3940) <= not(inputs(29));
    layer0_outputs(3941) <= (inputs(239)) and (inputs(25));
    layer0_outputs(3942) <= (inputs(40)) and (inputs(96));
    layer0_outputs(3943) <= (inputs(23)) or (inputs(109));
    layer0_outputs(3944) <= (inputs(159)) and (inputs(27));
    layer0_outputs(3945) <= (inputs(9)) and not (inputs(34));
    layer0_outputs(3946) <= not(inputs(32)) or (inputs(11));
    layer0_outputs(3947) <= not(inputs(225));
    layer0_outputs(3948) <= inputs(169);
    layer0_outputs(3949) <= not(inputs(246));
    layer0_outputs(3950) <= not((inputs(104)) or (inputs(75)));
    layer0_outputs(3951) <= (inputs(213)) xor (inputs(72));
    layer0_outputs(3952) <= not(inputs(128));
    layer0_outputs(3953) <= not((inputs(205)) and (inputs(158)));
    layer0_outputs(3954) <= not((inputs(248)) or (inputs(185)));
    layer0_outputs(3955) <= (inputs(139)) and not (inputs(228));
    layer0_outputs(3956) <= (inputs(203)) and not (inputs(180));
    layer0_outputs(3957) <= (inputs(172)) or (inputs(210));
    layer0_outputs(3958) <= not(inputs(11));
    layer0_outputs(3959) <= inputs(134);
    layer0_outputs(3960) <= not(inputs(55)) or (inputs(255));
    layer0_outputs(3961) <= '0';
    layer0_outputs(3962) <= (inputs(68)) and not (inputs(198));
    layer0_outputs(3963) <= not((inputs(49)) or (inputs(54)));
    layer0_outputs(3964) <= (inputs(49)) xor (inputs(135));
    layer0_outputs(3965) <= not(inputs(131));
    layer0_outputs(3966) <= not((inputs(121)) or (inputs(114)));
    layer0_outputs(3967) <= inputs(78);
    layer0_outputs(3968) <= '0';
    layer0_outputs(3969) <= (inputs(62)) and not (inputs(211));
    layer0_outputs(3970) <= '1';
    layer0_outputs(3971) <= not(inputs(93));
    layer0_outputs(3972) <= (inputs(148)) xor (inputs(116));
    layer0_outputs(3973) <= (inputs(216)) and not (inputs(35));
    layer0_outputs(3974) <= (inputs(133)) xor (inputs(95));
    layer0_outputs(3975) <= (inputs(3)) and not (inputs(192));
    layer0_outputs(3976) <= (inputs(240)) and not (inputs(80));
    layer0_outputs(3977) <= (inputs(35)) and not (inputs(124));
    layer0_outputs(3978) <= (inputs(106)) and not (inputs(157));
    layer0_outputs(3979) <= not((inputs(146)) xor (inputs(184)));
    layer0_outputs(3980) <= (inputs(228)) and not (inputs(251));
    layer0_outputs(3981) <= (inputs(134)) and not (inputs(184));
    layer0_outputs(3982) <= inputs(128);
    layer0_outputs(3983) <= not(inputs(77));
    layer0_outputs(3984) <= (inputs(73)) and (inputs(64));
    layer0_outputs(3985) <= not(inputs(191)) or (inputs(51));
    layer0_outputs(3986) <= inputs(40);
    layer0_outputs(3987) <= '1';
    layer0_outputs(3988) <= (inputs(190)) or (inputs(132));
    layer0_outputs(3989) <= (inputs(53)) and not (inputs(45));
    layer0_outputs(3990) <= '1';
    layer0_outputs(3991) <= not((inputs(14)) xor (inputs(107)));
    layer0_outputs(3992) <= (inputs(104)) and (inputs(151));
    layer0_outputs(3993) <= not(inputs(236));
    layer0_outputs(3994) <= inputs(113);
    layer0_outputs(3995) <= (inputs(37)) and not (inputs(181));
    layer0_outputs(3996) <= (inputs(107)) and not (inputs(177));
    layer0_outputs(3997) <= (inputs(184)) or (inputs(174));
    layer0_outputs(3998) <= not((inputs(142)) and (inputs(8)));
    layer0_outputs(3999) <= not(inputs(41)) or (inputs(160));
    layer0_outputs(4000) <= not(inputs(205));
    layer0_outputs(4001) <= not(inputs(89)) or (inputs(185));
    layer0_outputs(4002) <= (inputs(110)) or (inputs(120));
    layer0_outputs(4003) <= inputs(248);
    layer0_outputs(4004) <= not(inputs(224));
    layer0_outputs(4005) <= inputs(115);
    layer0_outputs(4006) <= not((inputs(114)) or (inputs(162)));
    layer0_outputs(4007) <= not(inputs(229)) or (inputs(1));
    layer0_outputs(4008) <= (inputs(87)) or (inputs(252));
    layer0_outputs(4009) <= (inputs(214)) and not (inputs(50));
    layer0_outputs(4010) <= (inputs(11)) xor (inputs(156));
    layer0_outputs(4011) <= (inputs(231)) or (inputs(55));
    layer0_outputs(4012) <= (inputs(77)) or (inputs(238));
    layer0_outputs(4013) <= not((inputs(216)) or (inputs(130)));
    layer0_outputs(4014) <= not((inputs(227)) or (inputs(89)));
    layer0_outputs(4015) <= '0';
    layer0_outputs(4016) <= '1';
    layer0_outputs(4017) <= (inputs(112)) or (inputs(151));
    layer0_outputs(4018) <= '0';
    layer0_outputs(4019) <= (inputs(91)) and (inputs(134));
    layer0_outputs(4020) <= not(inputs(155)) or (inputs(235));
    layer0_outputs(4021) <= (inputs(202)) or (inputs(4));
    layer0_outputs(4022) <= '0';
    layer0_outputs(4023) <= not((inputs(179)) or (inputs(32)));
    layer0_outputs(4024) <= not(inputs(252)) or (inputs(144));
    layer0_outputs(4025) <= (inputs(224)) and not (inputs(235));
    layer0_outputs(4026) <= (inputs(47)) xor (inputs(136));
    layer0_outputs(4027) <= not((inputs(14)) or (inputs(139)));
    layer0_outputs(4028) <= not((inputs(67)) xor (inputs(92)));
    layer0_outputs(4029) <= inputs(215);
    layer0_outputs(4030) <= not(inputs(170)) or (inputs(84));
    layer0_outputs(4031) <= (inputs(33)) and not (inputs(47));
    layer0_outputs(4032) <= '1';
    layer0_outputs(4033) <= inputs(101);
    layer0_outputs(4034) <= not((inputs(116)) xor (inputs(149)));
    layer0_outputs(4035) <= not((inputs(161)) or (inputs(251)));
    layer0_outputs(4036) <= (inputs(214)) or (inputs(111));
    layer0_outputs(4037) <= not(inputs(175));
    layer0_outputs(4038) <= not((inputs(38)) or (inputs(203)));
    layer0_outputs(4039) <= (inputs(236)) or (inputs(153));
    layer0_outputs(4040) <= not((inputs(58)) or (inputs(184)));
    layer0_outputs(4041) <= not((inputs(0)) or (inputs(37)));
    layer0_outputs(4042) <= not(inputs(147));
    layer0_outputs(4043) <= not((inputs(1)) or (inputs(208)));
    layer0_outputs(4044) <= not(inputs(75)) or (inputs(184));
    layer0_outputs(4045) <= not(inputs(178));
    layer0_outputs(4046) <= (inputs(94)) or (inputs(9));
    layer0_outputs(4047) <= not(inputs(184));
    layer0_outputs(4048) <= (inputs(56)) and (inputs(26));
    layer0_outputs(4049) <= not((inputs(81)) xor (inputs(25)));
    layer0_outputs(4050) <= (inputs(190)) and not (inputs(123));
    layer0_outputs(4051) <= not(inputs(227));
    layer0_outputs(4052) <= not((inputs(122)) or (inputs(19)));
    layer0_outputs(4053) <= not(inputs(109)) or (inputs(149));
    layer0_outputs(4054) <= inputs(146);
    layer0_outputs(4055) <= not(inputs(41));
    layer0_outputs(4056) <= not((inputs(248)) xor (inputs(167)));
    layer0_outputs(4057) <= not((inputs(109)) xor (inputs(174)));
    layer0_outputs(4058) <= not((inputs(21)) and (inputs(79)));
    layer0_outputs(4059) <= '0';
    layer0_outputs(4060) <= not((inputs(75)) xor (inputs(244)));
    layer0_outputs(4061) <= '0';
    layer0_outputs(4062) <= (inputs(80)) or (inputs(170));
    layer0_outputs(4063) <= not(inputs(58)) or (inputs(237));
    layer0_outputs(4064) <= '0';
    layer0_outputs(4065) <= (inputs(76)) and not (inputs(129));
    layer0_outputs(4066) <= inputs(26);
    layer0_outputs(4067) <= (inputs(15)) and (inputs(49));
    layer0_outputs(4068) <= not(inputs(254));
    layer0_outputs(4069) <= not(inputs(254)) or (inputs(130));
    layer0_outputs(4070) <= not(inputs(82));
    layer0_outputs(4071) <= not(inputs(138)) or (inputs(196));
    layer0_outputs(4072) <= (inputs(80)) and not (inputs(209));
    layer0_outputs(4073) <= (inputs(237)) and not (inputs(43));
    layer0_outputs(4074) <= (inputs(189)) or (inputs(132));
    layer0_outputs(4075) <= (inputs(148)) xor (inputs(202));
    layer0_outputs(4076) <= '0';
    layer0_outputs(4077) <= (inputs(62)) and not (inputs(202));
    layer0_outputs(4078) <= inputs(114);
    layer0_outputs(4079) <= not(inputs(46)) or (inputs(142));
    layer0_outputs(4080) <= not(inputs(105)) or (inputs(237));
    layer0_outputs(4081) <= inputs(42);
    layer0_outputs(4082) <= not(inputs(66)) or (inputs(117));
    layer0_outputs(4083) <= inputs(60);
    layer0_outputs(4084) <= '1';
    layer0_outputs(4085) <= inputs(169);
    layer0_outputs(4086) <= not(inputs(183));
    layer0_outputs(4087) <= inputs(196);
    layer0_outputs(4088) <= not((inputs(178)) and (inputs(240)));
    layer0_outputs(4089) <= (inputs(161)) and (inputs(191));
    layer0_outputs(4090) <= (inputs(153)) and not (inputs(213));
    layer0_outputs(4091) <= not((inputs(209)) and (inputs(79)));
    layer0_outputs(4092) <= (inputs(204)) xor (inputs(222));
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= not(inputs(174)) or (inputs(126));
    layer0_outputs(4095) <= not(inputs(102));
    layer0_outputs(4096) <= '0';
    layer0_outputs(4097) <= '1';
    layer0_outputs(4098) <= inputs(134);
    layer0_outputs(4099) <= not(inputs(204));
    layer0_outputs(4100) <= '1';
    layer0_outputs(4101) <= (inputs(221)) and (inputs(124));
    layer0_outputs(4102) <= (inputs(24)) xor (inputs(16));
    layer0_outputs(4103) <= (inputs(134)) or (inputs(77));
    layer0_outputs(4104) <= not((inputs(25)) and (inputs(224)));
    layer0_outputs(4105) <= inputs(121);
    layer0_outputs(4106) <= inputs(73);
    layer0_outputs(4107) <= (inputs(21)) or (inputs(155));
    layer0_outputs(4108) <= inputs(81);
    layer0_outputs(4109) <= not((inputs(197)) or (inputs(219)));
    layer0_outputs(4110) <= (inputs(166)) and not (inputs(133));
    layer0_outputs(4111) <= not(inputs(85));
    layer0_outputs(4112) <= (inputs(190)) and (inputs(189));
    layer0_outputs(4113) <= not(inputs(65)) or (inputs(90));
    layer0_outputs(4114) <= not((inputs(233)) or (inputs(126)));
    layer0_outputs(4115) <= (inputs(192)) and not (inputs(16));
    layer0_outputs(4116) <= not(inputs(54));
    layer0_outputs(4117) <= not(inputs(214)) or (inputs(251));
    layer0_outputs(4118) <= not((inputs(255)) and (inputs(49)));
    layer0_outputs(4119) <= not((inputs(166)) and (inputs(150)));
    layer0_outputs(4120) <= (inputs(198)) and not (inputs(10));
    layer0_outputs(4121) <= inputs(77);
    layer0_outputs(4122) <= inputs(247);
    layer0_outputs(4123) <= '1';
    layer0_outputs(4124) <= (inputs(131)) and not (inputs(207));
    layer0_outputs(4125) <= not(inputs(29)) or (inputs(30));
    layer0_outputs(4126) <= not(inputs(149)) or (inputs(96));
    layer0_outputs(4127) <= not(inputs(63));
    layer0_outputs(4128) <= not((inputs(62)) or (inputs(189)));
    layer0_outputs(4129) <= inputs(132);
    layer0_outputs(4130) <= not(inputs(241)) or (inputs(152));
    layer0_outputs(4131) <= inputs(134);
    layer0_outputs(4132) <= not((inputs(148)) and (inputs(30)));
    layer0_outputs(4133) <= (inputs(175)) and (inputs(111));
    layer0_outputs(4134) <= (inputs(75)) xor (inputs(189));
    layer0_outputs(4135) <= not(inputs(197));
    layer0_outputs(4136) <= inputs(193);
    layer0_outputs(4137) <= inputs(45);
    layer0_outputs(4138) <= not(inputs(52));
    layer0_outputs(4139) <= (inputs(11)) and not (inputs(75));
    layer0_outputs(4140) <= (inputs(211)) and not (inputs(251));
    layer0_outputs(4141) <= not((inputs(179)) or (inputs(107)));
    layer0_outputs(4142) <= not((inputs(42)) and (inputs(19)));
    layer0_outputs(4143) <= not(inputs(46)) or (inputs(79));
    layer0_outputs(4144) <= inputs(78);
    layer0_outputs(4145) <= inputs(221);
    layer0_outputs(4146) <= not(inputs(113));
    layer0_outputs(4147) <= (inputs(173)) or (inputs(43));
    layer0_outputs(4148) <= inputs(82);
    layer0_outputs(4149) <= not(inputs(43)) or (inputs(49));
    layer0_outputs(4150) <= (inputs(0)) or (inputs(133));
    layer0_outputs(4151) <= not((inputs(16)) xor (inputs(235)));
    layer0_outputs(4152) <= not(inputs(20));
    layer0_outputs(4153) <= not(inputs(20)) or (inputs(217));
    layer0_outputs(4154) <= '0';
    layer0_outputs(4155) <= not((inputs(221)) or (inputs(215)));
    layer0_outputs(4156) <= not((inputs(43)) and (inputs(72)));
    layer0_outputs(4157) <= (inputs(202)) and not (inputs(81));
    layer0_outputs(4158) <= not(inputs(203)) or (inputs(89));
    layer0_outputs(4159) <= (inputs(141)) and not (inputs(25));
    layer0_outputs(4160) <= inputs(41);
    layer0_outputs(4161) <= not(inputs(206));
    layer0_outputs(4162) <= inputs(137);
    layer0_outputs(4163) <= (inputs(80)) or (inputs(182));
    layer0_outputs(4164) <= not(inputs(234));
    layer0_outputs(4165) <= (inputs(9)) and not (inputs(248));
    layer0_outputs(4166) <= not((inputs(175)) and (inputs(130)));
    layer0_outputs(4167) <= not(inputs(53)) or (inputs(24));
    layer0_outputs(4168) <= inputs(70);
    layer0_outputs(4169) <= not(inputs(135));
    layer0_outputs(4170) <= (inputs(34)) and not (inputs(137));
    layer0_outputs(4171) <= (inputs(109)) or (inputs(53));
    layer0_outputs(4172) <= '0';
    layer0_outputs(4173) <= (inputs(20)) or (inputs(225));
    layer0_outputs(4174) <= not((inputs(80)) xor (inputs(255)));
    layer0_outputs(4175) <= inputs(43);
    layer0_outputs(4176) <= not((inputs(54)) or (inputs(36)));
    layer0_outputs(4177) <= (inputs(156)) and not (inputs(63));
    layer0_outputs(4178) <= (inputs(235)) and (inputs(57));
    layer0_outputs(4179) <= (inputs(141)) and not (inputs(30));
    layer0_outputs(4180) <= not((inputs(206)) xor (inputs(64)));
    layer0_outputs(4181) <= (inputs(0)) and not (inputs(77));
    layer0_outputs(4182) <= not((inputs(97)) or (inputs(40)));
    layer0_outputs(4183) <= not(inputs(152));
    layer0_outputs(4184) <= not(inputs(30)) or (inputs(213));
    layer0_outputs(4185) <= not(inputs(56));
    layer0_outputs(4186) <= (inputs(215)) and not (inputs(174));
    layer0_outputs(4187) <= not(inputs(105)) or (inputs(139));
    layer0_outputs(4188) <= inputs(185);
    layer0_outputs(4189) <= not((inputs(102)) or (inputs(15)));
    layer0_outputs(4190) <= inputs(76);
    layer0_outputs(4191) <= not((inputs(15)) xor (inputs(113)));
    layer0_outputs(4192) <= (inputs(47)) and (inputs(223));
    layer0_outputs(4193) <= not((inputs(151)) xor (inputs(127)));
    layer0_outputs(4194) <= not(inputs(217));
    layer0_outputs(4195) <= (inputs(107)) and (inputs(27));
    layer0_outputs(4196) <= (inputs(95)) and not (inputs(165));
    layer0_outputs(4197) <= inputs(80);
    layer0_outputs(4198) <= not(inputs(148));
    layer0_outputs(4199) <= not(inputs(58));
    layer0_outputs(4200) <= not((inputs(115)) xor (inputs(111)));
    layer0_outputs(4201) <= (inputs(156)) or (inputs(156));
    layer0_outputs(4202) <= inputs(180);
    layer0_outputs(4203) <= (inputs(98)) or (inputs(104));
    layer0_outputs(4204) <= not((inputs(56)) xor (inputs(71)));
    layer0_outputs(4205) <= (inputs(210)) and not (inputs(15));
    layer0_outputs(4206) <= not(inputs(9)) or (inputs(187));
    layer0_outputs(4207) <= not((inputs(19)) or (inputs(171)));
    layer0_outputs(4208) <= inputs(76);
    layer0_outputs(4209) <= not((inputs(212)) or (inputs(36)));
    layer0_outputs(4210) <= not(inputs(27));
    layer0_outputs(4211) <= (inputs(207)) and not (inputs(57));
    layer0_outputs(4212) <= not(inputs(77));
    layer0_outputs(4213) <= inputs(19);
    layer0_outputs(4214) <= inputs(208);
    layer0_outputs(4215) <= (inputs(92)) or (inputs(249));
    layer0_outputs(4216) <= not(inputs(89));
    layer0_outputs(4217) <= '0';
    layer0_outputs(4218) <= not(inputs(121)) or (inputs(5));
    layer0_outputs(4219) <= (inputs(18)) or (inputs(131));
    layer0_outputs(4220) <= (inputs(182)) or (inputs(66));
    layer0_outputs(4221) <= inputs(185);
    layer0_outputs(4222) <= not((inputs(27)) xor (inputs(38)));
    layer0_outputs(4223) <= (inputs(53)) xor (inputs(46));
    layer0_outputs(4224) <= not((inputs(107)) or (inputs(41)));
    layer0_outputs(4225) <= '0';
    layer0_outputs(4226) <= not((inputs(241)) or (inputs(179)));
    layer0_outputs(4227) <= (inputs(146)) and not (inputs(62));
    layer0_outputs(4228) <= not((inputs(104)) or (inputs(94)));
    layer0_outputs(4229) <= not((inputs(0)) xor (inputs(61)));
    layer0_outputs(4230) <= inputs(171);
    layer0_outputs(4231) <= not(inputs(227)) or (inputs(158));
    layer0_outputs(4232) <= not((inputs(80)) or (inputs(58)));
    layer0_outputs(4233) <= (inputs(189)) and not (inputs(235));
    layer0_outputs(4234) <= not(inputs(116));
    layer0_outputs(4235) <= inputs(161);
    layer0_outputs(4236) <= (inputs(124)) and not (inputs(3));
    layer0_outputs(4237) <= (inputs(198)) and not (inputs(226));
    layer0_outputs(4238) <= not((inputs(66)) or (inputs(255)));
    layer0_outputs(4239) <= inputs(215);
    layer0_outputs(4240) <= not(inputs(39)) or (inputs(61));
    layer0_outputs(4241) <= (inputs(114)) or (inputs(91));
    layer0_outputs(4242) <= '0';
    layer0_outputs(4243) <= '1';
    layer0_outputs(4244) <= (inputs(102)) and (inputs(126));
    layer0_outputs(4245) <= not(inputs(192)) or (inputs(69));
    layer0_outputs(4246) <= not((inputs(27)) and (inputs(160)));
    layer0_outputs(4247) <= (inputs(41)) and not (inputs(206));
    layer0_outputs(4248) <= not((inputs(163)) or (inputs(73)));
    layer0_outputs(4249) <= inputs(52);
    layer0_outputs(4250) <= inputs(191);
    layer0_outputs(4251) <= '1';
    layer0_outputs(4252) <= (inputs(122)) and not (inputs(56));
    layer0_outputs(4253) <= not(inputs(43)) or (inputs(71));
    layer0_outputs(4254) <= (inputs(34)) or (inputs(191));
    layer0_outputs(4255) <= not(inputs(90)) or (inputs(220));
    layer0_outputs(4256) <= not(inputs(181)) or (inputs(125));
    layer0_outputs(4257) <= inputs(79);
    layer0_outputs(4258) <= inputs(242);
    layer0_outputs(4259) <= '0';
    layer0_outputs(4260) <= inputs(87);
    layer0_outputs(4261) <= inputs(227);
    layer0_outputs(4262) <= inputs(206);
    layer0_outputs(4263) <= '1';
    layer0_outputs(4264) <= not(inputs(190));
    layer0_outputs(4265) <= (inputs(98)) and not (inputs(63));
    layer0_outputs(4266) <= (inputs(177)) xor (inputs(8));
    layer0_outputs(4267) <= (inputs(211)) and not (inputs(193));
    layer0_outputs(4268) <= not(inputs(9));
    layer0_outputs(4269) <= (inputs(219)) xor (inputs(30));
    layer0_outputs(4270) <= not((inputs(195)) and (inputs(244)));
    layer0_outputs(4271) <= (inputs(191)) or (inputs(37));
    layer0_outputs(4272) <= (inputs(118)) and not (inputs(2));
    layer0_outputs(4273) <= (inputs(6)) or (inputs(83));
    layer0_outputs(4274) <= not(inputs(242));
    layer0_outputs(4275) <= not(inputs(213)) or (inputs(67));
    layer0_outputs(4276) <= not((inputs(192)) xor (inputs(44)));
    layer0_outputs(4277) <= not(inputs(117));
    layer0_outputs(4278) <= '1';
    layer0_outputs(4279) <= (inputs(58)) xor (inputs(89));
    layer0_outputs(4280) <= (inputs(12)) xor (inputs(236));
    layer0_outputs(4281) <= not(inputs(185));
    layer0_outputs(4282) <= '0';
    layer0_outputs(4283) <= not((inputs(108)) xor (inputs(82)));
    layer0_outputs(4284) <= not((inputs(230)) or (inputs(6)));
    layer0_outputs(4285) <= not(inputs(240));
    layer0_outputs(4286) <= (inputs(39)) xor (inputs(9));
    layer0_outputs(4287) <= not(inputs(191)) or (inputs(236));
    layer0_outputs(4288) <= (inputs(105)) or (inputs(65));
    layer0_outputs(4289) <= not(inputs(67));
    layer0_outputs(4290) <= (inputs(56)) and not (inputs(61));
    layer0_outputs(4291) <= not((inputs(198)) and (inputs(95)));
    layer0_outputs(4292) <= inputs(172);
    layer0_outputs(4293) <= inputs(97);
    layer0_outputs(4294) <= not((inputs(12)) xor (inputs(96)));
    layer0_outputs(4295) <= inputs(158);
    layer0_outputs(4296) <= not((inputs(25)) and (inputs(194)));
    layer0_outputs(4297) <= not((inputs(121)) or (inputs(61)));
    layer0_outputs(4298) <= not((inputs(57)) or (inputs(221)));
    layer0_outputs(4299) <= '1';
    layer0_outputs(4300) <= (inputs(242)) and not (inputs(212));
    layer0_outputs(4301) <= inputs(155);
    layer0_outputs(4302) <= (inputs(157)) or (inputs(79));
    layer0_outputs(4303) <= (inputs(34)) or (inputs(221));
    layer0_outputs(4304) <= inputs(166);
    layer0_outputs(4305) <= (inputs(253)) and not (inputs(236));
    layer0_outputs(4306) <= not((inputs(64)) or (inputs(198)));
    layer0_outputs(4307) <= (inputs(160)) and not (inputs(218));
    layer0_outputs(4308) <= not((inputs(183)) and (inputs(18)));
    layer0_outputs(4309) <= not((inputs(202)) or (inputs(121)));
    layer0_outputs(4310) <= (inputs(155)) and (inputs(127));
    layer0_outputs(4311) <= (inputs(28)) and not (inputs(8));
    layer0_outputs(4312) <= not((inputs(15)) and (inputs(67)));
    layer0_outputs(4313) <= not((inputs(96)) xor (inputs(76)));
    layer0_outputs(4314) <= '0';
    layer0_outputs(4315) <= (inputs(119)) and not (inputs(44));
    layer0_outputs(4316) <= '0';
    layer0_outputs(4317) <= not((inputs(89)) and (inputs(94)));
    layer0_outputs(4318) <= not((inputs(149)) xor (inputs(63)));
    layer0_outputs(4319) <= (inputs(114)) or (inputs(171));
    layer0_outputs(4320) <= not(inputs(116));
    layer0_outputs(4321) <= inputs(82);
    layer0_outputs(4322) <= (inputs(138)) xor (inputs(178));
    layer0_outputs(4323) <= not(inputs(107));
    layer0_outputs(4324) <= not((inputs(203)) or (inputs(167)));
    layer0_outputs(4325) <= (inputs(99)) and (inputs(19));
    layer0_outputs(4326) <= '0';
    layer0_outputs(4327) <= not((inputs(22)) or (inputs(70)));
    layer0_outputs(4328) <= (inputs(164)) and not (inputs(76));
    layer0_outputs(4329) <= (inputs(119)) and (inputs(195));
    layer0_outputs(4330) <= (inputs(21)) xor (inputs(255));
    layer0_outputs(4331) <= inputs(16);
    layer0_outputs(4332) <= not(inputs(68)) or (inputs(146));
    layer0_outputs(4333) <= (inputs(80)) or (inputs(48));
    layer0_outputs(4334) <= (inputs(89)) and (inputs(190));
    layer0_outputs(4335) <= not(inputs(155)) or (inputs(60));
    layer0_outputs(4336) <= not(inputs(147)) or (inputs(14));
    layer0_outputs(4337) <= not(inputs(120));
    layer0_outputs(4338) <= inputs(73);
    layer0_outputs(4339) <= not(inputs(55));
    layer0_outputs(4340) <= (inputs(102)) and not (inputs(65));
    layer0_outputs(4341) <= (inputs(148)) xor (inputs(174));
    layer0_outputs(4342) <= (inputs(199)) and not (inputs(25));
    layer0_outputs(4343) <= (inputs(155)) and (inputs(130));
    layer0_outputs(4344) <= not((inputs(212)) or (inputs(97)));
    layer0_outputs(4345) <= (inputs(25)) and not (inputs(180));
    layer0_outputs(4346) <= inputs(220);
    layer0_outputs(4347) <= inputs(108);
    layer0_outputs(4348) <= (inputs(80)) and not (inputs(82));
    layer0_outputs(4349) <= not((inputs(3)) xor (inputs(131)));
    layer0_outputs(4350) <= not(inputs(138));
    layer0_outputs(4351) <= not((inputs(13)) xor (inputs(118)));
    layer0_outputs(4352) <= (inputs(56)) and not (inputs(230));
    layer0_outputs(4353) <= inputs(5);
    layer0_outputs(4354) <= not((inputs(102)) or (inputs(143)));
    layer0_outputs(4355) <= inputs(91);
    layer0_outputs(4356) <= not((inputs(149)) or (inputs(60)));
    layer0_outputs(4357) <= not((inputs(94)) or (inputs(11)));
    layer0_outputs(4358) <= not((inputs(38)) or (inputs(234)));
    layer0_outputs(4359) <= not((inputs(12)) and (inputs(209)));
    layer0_outputs(4360) <= (inputs(38)) or (inputs(164));
    layer0_outputs(4361) <= '0';
    layer0_outputs(4362) <= (inputs(174)) and not (inputs(28));
    layer0_outputs(4363) <= (inputs(137)) or (inputs(33));
    layer0_outputs(4364) <= not(inputs(140));
    layer0_outputs(4365) <= not((inputs(221)) xor (inputs(236)));
    layer0_outputs(4366) <= (inputs(48)) xor (inputs(51));
    layer0_outputs(4367) <= '1';
    layer0_outputs(4368) <= (inputs(210)) or (inputs(72));
    layer0_outputs(4369) <= not((inputs(174)) and (inputs(24)));
    layer0_outputs(4370) <= (inputs(69)) xor (inputs(0));
    layer0_outputs(4371) <= '0';
    layer0_outputs(4372) <= not(inputs(151));
    layer0_outputs(4373) <= (inputs(189)) and not (inputs(218));
    layer0_outputs(4374) <= (inputs(181)) and (inputs(54));
    layer0_outputs(4375) <= '0';
    layer0_outputs(4376) <= '0';
    layer0_outputs(4377) <= not(inputs(156));
    layer0_outputs(4378) <= (inputs(78)) and not (inputs(227));
    layer0_outputs(4379) <= (inputs(234)) xor (inputs(226));
    layer0_outputs(4380) <= not(inputs(70));
    layer0_outputs(4381) <= not((inputs(12)) xor (inputs(71)));
    layer0_outputs(4382) <= inputs(192);
    layer0_outputs(4383) <= not(inputs(252)) or (inputs(11));
    layer0_outputs(4384) <= not((inputs(39)) or (inputs(252)));
    layer0_outputs(4385) <= not(inputs(220));
    layer0_outputs(4386) <= not(inputs(110)) or (inputs(220));
    layer0_outputs(4387) <= not((inputs(79)) xor (inputs(6)));
    layer0_outputs(4388) <= (inputs(1)) xor (inputs(117));
    layer0_outputs(4389) <= '0';
    layer0_outputs(4390) <= not(inputs(5));
    layer0_outputs(4391) <= (inputs(195)) and (inputs(7));
    layer0_outputs(4392) <= not(inputs(126)) or (inputs(250));
    layer0_outputs(4393) <= (inputs(108)) and (inputs(25));
    layer0_outputs(4394) <= not(inputs(147)) or (inputs(23));
    layer0_outputs(4395) <= inputs(56);
    layer0_outputs(4396) <= (inputs(105)) or (inputs(54));
    layer0_outputs(4397) <= not(inputs(238));
    layer0_outputs(4398) <= '0';
    layer0_outputs(4399) <= not((inputs(156)) xor (inputs(232)));
    layer0_outputs(4400) <= inputs(99);
    layer0_outputs(4401) <= not(inputs(247)) or (inputs(0));
    layer0_outputs(4402) <= not(inputs(57)) or (inputs(136));
    layer0_outputs(4403) <= inputs(142);
    layer0_outputs(4404) <= '0';
    layer0_outputs(4405) <= (inputs(217)) and not (inputs(79));
    layer0_outputs(4406) <= not(inputs(85));
    layer0_outputs(4407) <= (inputs(198)) and not (inputs(236));
    layer0_outputs(4408) <= (inputs(103)) and not (inputs(240));
    layer0_outputs(4409) <= '1';
    layer0_outputs(4410) <= not((inputs(29)) and (inputs(193)));
    layer0_outputs(4411) <= '1';
    layer0_outputs(4412) <= inputs(147);
    layer0_outputs(4413) <= not(inputs(58)) or (inputs(10));
    layer0_outputs(4414) <= inputs(238);
    layer0_outputs(4415) <= (inputs(244)) and not (inputs(172));
    layer0_outputs(4416) <= (inputs(79)) xor (inputs(55));
    layer0_outputs(4417) <= not(inputs(65)) or (inputs(8));
    layer0_outputs(4418) <= (inputs(228)) and not (inputs(32));
    layer0_outputs(4419) <= inputs(6);
    layer0_outputs(4420) <= not((inputs(82)) xor (inputs(214)));
    layer0_outputs(4421) <= (inputs(102)) and not (inputs(243));
    layer0_outputs(4422) <= not(inputs(173));
    layer0_outputs(4423) <= not(inputs(128)) or (inputs(97));
    layer0_outputs(4424) <= not((inputs(89)) or (inputs(171)));
    layer0_outputs(4425) <= (inputs(64)) and not (inputs(0));
    layer0_outputs(4426) <= not((inputs(149)) and (inputs(176)));
    layer0_outputs(4427) <= (inputs(64)) and not (inputs(148));
    layer0_outputs(4428) <= '0';
    layer0_outputs(4429) <= (inputs(84)) xor (inputs(164));
    layer0_outputs(4430) <= (inputs(10)) xor (inputs(122));
    layer0_outputs(4431) <= (inputs(149)) and not (inputs(50));
    layer0_outputs(4432) <= not((inputs(49)) and (inputs(110)));
    layer0_outputs(4433) <= not(inputs(119));
    layer0_outputs(4434) <= not(inputs(180)) or (inputs(52));
    layer0_outputs(4435) <= '1';
    layer0_outputs(4436) <= not(inputs(8));
    layer0_outputs(4437) <= not(inputs(189));
    layer0_outputs(4438) <= (inputs(87)) xor (inputs(251));
    layer0_outputs(4439) <= not(inputs(67)) or (inputs(17));
    layer0_outputs(4440) <= '1';
    layer0_outputs(4441) <= not((inputs(219)) or (inputs(83)));
    layer0_outputs(4442) <= inputs(19);
    layer0_outputs(4443) <= not((inputs(107)) or (inputs(122)));
    layer0_outputs(4444) <= '0';
    layer0_outputs(4445) <= (inputs(21)) and not (inputs(177));
    layer0_outputs(4446) <= not(inputs(212)) or (inputs(80));
    layer0_outputs(4447) <= not((inputs(142)) xor (inputs(183)));
    layer0_outputs(4448) <= inputs(199);
    layer0_outputs(4449) <= inputs(122);
    layer0_outputs(4450) <= not(inputs(228)) or (inputs(45));
    layer0_outputs(4451) <= not(inputs(132));
    layer0_outputs(4452) <= (inputs(181)) and not (inputs(50));
    layer0_outputs(4453) <= not((inputs(230)) or (inputs(45)));
    layer0_outputs(4454) <= '1';
    layer0_outputs(4455) <= not((inputs(205)) or (inputs(131)));
    layer0_outputs(4456) <= '1';
    layer0_outputs(4457) <= '1';
    layer0_outputs(4458) <= inputs(195);
    layer0_outputs(4459) <= '1';
    layer0_outputs(4460) <= not((inputs(146)) xor (inputs(194)));
    layer0_outputs(4461) <= (inputs(100)) or (inputs(91));
    layer0_outputs(4462) <= not(inputs(131));
    layer0_outputs(4463) <= '0';
    layer0_outputs(4464) <= (inputs(202)) and not (inputs(214));
    layer0_outputs(4465) <= inputs(216);
    layer0_outputs(4466) <= (inputs(115)) and not (inputs(32));
    layer0_outputs(4467) <= not((inputs(0)) and (inputs(124)));
    layer0_outputs(4468) <= not(inputs(23));
    layer0_outputs(4469) <= (inputs(254)) and not (inputs(68));
    layer0_outputs(4470) <= not((inputs(222)) or (inputs(187)));
    layer0_outputs(4471) <= not((inputs(74)) or (inputs(197)));
    layer0_outputs(4472) <= (inputs(131)) or (inputs(148));
    layer0_outputs(4473) <= not(inputs(41)) or (inputs(83));
    layer0_outputs(4474) <= (inputs(24)) xor (inputs(88));
    layer0_outputs(4475) <= (inputs(51)) and (inputs(161));
    layer0_outputs(4476) <= not((inputs(3)) or (inputs(201)));
    layer0_outputs(4477) <= not(inputs(96)) or (inputs(179));
    layer0_outputs(4478) <= not(inputs(31)) or (inputs(17));
    layer0_outputs(4479) <= (inputs(179)) or (inputs(174));
    layer0_outputs(4480) <= not(inputs(210));
    layer0_outputs(4481) <= not((inputs(118)) and (inputs(177)));
    layer0_outputs(4482) <= '1';
    layer0_outputs(4483) <= '1';
    layer0_outputs(4484) <= not(inputs(216)) or (inputs(114));
    layer0_outputs(4485) <= not((inputs(52)) and (inputs(228)));
    layer0_outputs(4486) <= (inputs(225)) and not (inputs(227));
    layer0_outputs(4487) <= inputs(244);
    layer0_outputs(4488) <= not((inputs(218)) xor (inputs(252)));
    layer0_outputs(4489) <= not(inputs(254)) or (inputs(56));
    layer0_outputs(4490) <= (inputs(104)) or (inputs(233));
    layer0_outputs(4491) <= not(inputs(229));
    layer0_outputs(4492) <= not((inputs(29)) xor (inputs(117)));
    layer0_outputs(4493) <= (inputs(163)) xor (inputs(57));
    layer0_outputs(4494) <= inputs(43);
    layer0_outputs(4495) <= not((inputs(191)) xor (inputs(178)));
    layer0_outputs(4496) <= not(inputs(134)) or (inputs(155));
    layer0_outputs(4497) <= not(inputs(87));
    layer0_outputs(4498) <= not((inputs(7)) xor (inputs(177)));
    layer0_outputs(4499) <= not(inputs(11)) or (inputs(202));
    layer0_outputs(4500) <= not(inputs(92));
    layer0_outputs(4501) <= not(inputs(117));
    layer0_outputs(4502) <= not(inputs(28)) or (inputs(23));
    layer0_outputs(4503) <= not(inputs(45));
    layer0_outputs(4504) <= not(inputs(138));
    layer0_outputs(4505) <= not(inputs(31)) or (inputs(9));
    layer0_outputs(4506) <= (inputs(116)) or (inputs(20));
    layer0_outputs(4507) <= '1';
    layer0_outputs(4508) <= not((inputs(209)) or (inputs(165)));
    layer0_outputs(4509) <= not(inputs(18));
    layer0_outputs(4510) <= not(inputs(216)) or (inputs(249));
    layer0_outputs(4511) <= not((inputs(75)) and (inputs(99)));
    layer0_outputs(4512) <= '0';
    layer0_outputs(4513) <= '0';
    layer0_outputs(4514) <= '0';
    layer0_outputs(4515) <= (inputs(135)) and not (inputs(139));
    layer0_outputs(4516) <= not(inputs(92));
    layer0_outputs(4517) <= not((inputs(197)) xor (inputs(126)));
    layer0_outputs(4518) <= inputs(183);
    layer0_outputs(4519) <= (inputs(106)) or (inputs(36));
    layer0_outputs(4520) <= not((inputs(45)) and (inputs(214)));
    layer0_outputs(4521) <= (inputs(224)) and (inputs(56));
    layer0_outputs(4522) <= (inputs(244)) or (inputs(128));
    layer0_outputs(4523) <= '1';
    layer0_outputs(4524) <= not(inputs(154));
    layer0_outputs(4525) <= not((inputs(148)) xor (inputs(179)));
    layer0_outputs(4526) <= (inputs(99)) and (inputs(225));
    layer0_outputs(4527) <= not(inputs(123));
    layer0_outputs(4528) <= not((inputs(212)) or (inputs(66)));
    layer0_outputs(4529) <= not((inputs(130)) and (inputs(94)));
    layer0_outputs(4530) <= not(inputs(194)) or (inputs(125));
    layer0_outputs(4531) <= not(inputs(253));
    layer0_outputs(4532) <= (inputs(245)) and not (inputs(188));
    layer0_outputs(4533) <= (inputs(207)) and not (inputs(164));
    layer0_outputs(4534) <= (inputs(100)) and (inputs(206));
    layer0_outputs(4535) <= '0';
    layer0_outputs(4536) <= not(inputs(56));
    layer0_outputs(4537) <= not((inputs(78)) and (inputs(189)));
    layer0_outputs(4538) <= inputs(167);
    layer0_outputs(4539) <= (inputs(2)) and not (inputs(39));
    layer0_outputs(4540) <= inputs(14);
    layer0_outputs(4541) <= not(inputs(66));
    layer0_outputs(4542) <= not(inputs(186));
    layer0_outputs(4543) <= (inputs(7)) xor (inputs(198));
    layer0_outputs(4544) <= not(inputs(241));
    layer0_outputs(4545) <= inputs(233);
    layer0_outputs(4546) <= '1';
    layer0_outputs(4547) <= not(inputs(8));
    layer0_outputs(4548) <= not((inputs(244)) or (inputs(205)));
    layer0_outputs(4549) <= (inputs(142)) xor (inputs(48));
    layer0_outputs(4550) <= (inputs(105)) or (inputs(172));
    layer0_outputs(4551) <= not(inputs(162)) or (inputs(86));
    layer0_outputs(4552) <= (inputs(25)) xor (inputs(5));
    layer0_outputs(4553) <= '1';
    layer0_outputs(4554) <= (inputs(2)) and not (inputs(54));
    layer0_outputs(4555) <= not(inputs(72));
    layer0_outputs(4556) <= (inputs(134)) and not (inputs(67));
    layer0_outputs(4557) <= inputs(178);
    layer0_outputs(4558) <= not(inputs(142)) or (inputs(201));
    layer0_outputs(4559) <= '1';
    layer0_outputs(4560) <= (inputs(157)) xor (inputs(129));
    layer0_outputs(4561) <= not((inputs(121)) xor (inputs(65)));
    layer0_outputs(4562) <= not(inputs(80)) or (inputs(0));
    layer0_outputs(4563) <= inputs(76);
    layer0_outputs(4564) <= '0';
    layer0_outputs(4565) <= '0';
    layer0_outputs(4566) <= not((inputs(246)) or (inputs(36)));
    layer0_outputs(4567) <= (inputs(141)) or (inputs(108));
    layer0_outputs(4568) <= (inputs(126)) and not (inputs(231));
    layer0_outputs(4569) <= not(inputs(73));
    layer0_outputs(4570) <= '1';
    layer0_outputs(4571) <= not((inputs(157)) or (inputs(35)));
    layer0_outputs(4572) <= not((inputs(43)) and (inputs(194)));
    layer0_outputs(4573) <= not((inputs(24)) xor (inputs(136)));
    layer0_outputs(4574) <= (inputs(21)) or (inputs(162));
    layer0_outputs(4575) <= not((inputs(29)) or (inputs(65)));
    layer0_outputs(4576) <= (inputs(38)) or (inputs(155));
    layer0_outputs(4577) <= not(inputs(72)) or (inputs(52));
    layer0_outputs(4578) <= not(inputs(231));
    layer0_outputs(4579) <= (inputs(88)) and not (inputs(36));
    layer0_outputs(4580) <= (inputs(116)) and not (inputs(159));
    layer0_outputs(4581) <= (inputs(83)) or (inputs(140));
    layer0_outputs(4582) <= not(inputs(98)) or (inputs(162));
    layer0_outputs(4583) <= (inputs(37)) or (inputs(129));
    layer0_outputs(4584) <= '0';
    layer0_outputs(4585) <= inputs(236);
    layer0_outputs(4586) <= not((inputs(50)) and (inputs(4)));
    layer0_outputs(4587) <= (inputs(156)) xor (inputs(227));
    layer0_outputs(4588) <= (inputs(25)) or (inputs(182));
    layer0_outputs(4589) <= (inputs(92)) and (inputs(7));
    layer0_outputs(4590) <= (inputs(156)) and not (inputs(18));
    layer0_outputs(4591) <= inputs(154);
    layer0_outputs(4592) <= (inputs(114)) and not (inputs(159));
    layer0_outputs(4593) <= inputs(166);
    layer0_outputs(4594) <= (inputs(252)) and (inputs(132));
    layer0_outputs(4595) <= not((inputs(134)) and (inputs(199)));
    layer0_outputs(4596) <= (inputs(108)) or (inputs(200));
    layer0_outputs(4597) <= (inputs(99)) or (inputs(209));
    layer0_outputs(4598) <= not(inputs(150)) or (inputs(66));
    layer0_outputs(4599) <= not((inputs(32)) or (inputs(221)));
    layer0_outputs(4600) <= (inputs(75)) and not (inputs(196));
    layer0_outputs(4601) <= not(inputs(101)) or (inputs(13));
    layer0_outputs(4602) <= inputs(251);
    layer0_outputs(4603) <= inputs(225);
    layer0_outputs(4604) <= not((inputs(149)) or (inputs(171)));
    layer0_outputs(4605) <= inputs(195);
    layer0_outputs(4606) <= inputs(198);
    layer0_outputs(4607) <= not(inputs(57));
    layer0_outputs(4608) <= (inputs(104)) or (inputs(211));
    layer0_outputs(4609) <= not((inputs(59)) or (inputs(75)));
    layer0_outputs(4610) <= '1';
    layer0_outputs(4611) <= not((inputs(45)) and (inputs(206)));
    layer0_outputs(4612) <= inputs(37);
    layer0_outputs(4613) <= (inputs(11)) or (inputs(214));
    layer0_outputs(4614) <= (inputs(35)) xor (inputs(198));
    layer0_outputs(4615) <= (inputs(70)) and not (inputs(103));
    layer0_outputs(4616) <= (inputs(141)) or (inputs(188));
    layer0_outputs(4617) <= inputs(226);
    layer0_outputs(4618) <= '0';
    layer0_outputs(4619) <= (inputs(12)) and not (inputs(28));
    layer0_outputs(4620) <= not(inputs(217));
    layer0_outputs(4621) <= (inputs(88)) xor (inputs(180));
    layer0_outputs(4622) <= not(inputs(252)) or (inputs(9));
    layer0_outputs(4623) <= (inputs(46)) and not (inputs(145));
    layer0_outputs(4624) <= not((inputs(231)) and (inputs(220)));
    layer0_outputs(4625) <= (inputs(158)) xor (inputs(192));
    layer0_outputs(4626) <= not((inputs(253)) or (inputs(3)));
    layer0_outputs(4627) <= (inputs(3)) xor (inputs(143));
    layer0_outputs(4628) <= not(inputs(18));
    layer0_outputs(4629) <= (inputs(213)) or (inputs(145));
    layer0_outputs(4630) <= inputs(40);
    layer0_outputs(4631) <= not((inputs(112)) and (inputs(210)));
    layer0_outputs(4632) <= not((inputs(142)) xor (inputs(58)));
    layer0_outputs(4633) <= (inputs(155)) or (inputs(251));
    layer0_outputs(4634) <= (inputs(222)) or (inputs(97));
    layer0_outputs(4635) <= (inputs(250)) and (inputs(244));
    layer0_outputs(4636) <= (inputs(48)) and not (inputs(29));
    layer0_outputs(4637) <= not(inputs(178));
    layer0_outputs(4638) <= '0';
    layer0_outputs(4639) <= inputs(136);
    layer0_outputs(4640) <= (inputs(99)) or (inputs(116));
    layer0_outputs(4641) <= inputs(218);
    layer0_outputs(4642) <= inputs(19);
    layer0_outputs(4643) <= not(inputs(248));
    layer0_outputs(4644) <= (inputs(196)) xor (inputs(176));
    layer0_outputs(4645) <= not(inputs(166)) or (inputs(81));
    layer0_outputs(4646) <= (inputs(94)) and not (inputs(160));
    layer0_outputs(4647) <= (inputs(246)) xor (inputs(98));
    layer0_outputs(4648) <= not(inputs(108));
    layer0_outputs(4649) <= (inputs(136)) and not (inputs(36));
    layer0_outputs(4650) <= not((inputs(234)) or (inputs(13)));
    layer0_outputs(4651) <= inputs(233);
    layer0_outputs(4652) <= inputs(150);
    layer0_outputs(4653) <= (inputs(158)) and (inputs(33));
    layer0_outputs(4654) <= not((inputs(201)) and (inputs(49)));
    layer0_outputs(4655) <= not((inputs(79)) xor (inputs(110)));
    layer0_outputs(4656) <= (inputs(132)) and not (inputs(211));
    layer0_outputs(4657) <= not((inputs(197)) xor (inputs(189)));
    layer0_outputs(4658) <= not(inputs(1)) or (inputs(155));
    layer0_outputs(4659) <= not(inputs(44));
    layer0_outputs(4660) <= not(inputs(11)) or (inputs(205));
    layer0_outputs(4661) <= not(inputs(240)) or (inputs(78));
    layer0_outputs(4662) <= (inputs(39)) and not (inputs(28));
    layer0_outputs(4663) <= '0';
    layer0_outputs(4664) <= (inputs(105)) and (inputs(196));
    layer0_outputs(4665) <= not((inputs(129)) and (inputs(109)));
    layer0_outputs(4666) <= (inputs(29)) xor (inputs(4));
    layer0_outputs(4667) <= not((inputs(43)) xor (inputs(60)));
    layer0_outputs(4668) <= not(inputs(238)) or (inputs(187));
    layer0_outputs(4669) <= not(inputs(92));
    layer0_outputs(4670) <= not(inputs(56)) or (inputs(119));
    layer0_outputs(4671) <= (inputs(52)) and not (inputs(247));
    layer0_outputs(4672) <= (inputs(59)) and not (inputs(248));
    layer0_outputs(4673) <= (inputs(214)) and not (inputs(64));
    layer0_outputs(4674) <= not(inputs(130)) or (inputs(153));
    layer0_outputs(4675) <= '1';
    layer0_outputs(4676) <= not((inputs(238)) and (inputs(142)));
    layer0_outputs(4677) <= '0';
    layer0_outputs(4678) <= inputs(250);
    layer0_outputs(4679) <= (inputs(7)) and (inputs(40));
    layer0_outputs(4680) <= not((inputs(165)) or (inputs(84)));
    layer0_outputs(4681) <= '0';
    layer0_outputs(4682) <= inputs(6);
    layer0_outputs(4683) <= (inputs(166)) and not (inputs(49));
    layer0_outputs(4684) <= '1';
    layer0_outputs(4685) <= inputs(93);
    layer0_outputs(4686) <= (inputs(96)) and not (inputs(217));
    layer0_outputs(4687) <= not((inputs(232)) or (inputs(249)));
    layer0_outputs(4688) <= (inputs(24)) or (inputs(182));
    layer0_outputs(4689) <= (inputs(158)) and not (inputs(47));
    layer0_outputs(4690) <= not((inputs(57)) or (inputs(33)));
    layer0_outputs(4691) <= not((inputs(228)) and (inputs(208)));
    layer0_outputs(4692) <= inputs(121);
    layer0_outputs(4693) <= (inputs(155)) and not (inputs(228));
    layer0_outputs(4694) <= (inputs(87)) xor (inputs(49));
    layer0_outputs(4695) <= not(inputs(65));
    layer0_outputs(4696) <= (inputs(243)) or (inputs(247));
    layer0_outputs(4697) <= (inputs(38)) or (inputs(29));
    layer0_outputs(4698) <= not(inputs(94)) or (inputs(176));
    layer0_outputs(4699) <= not(inputs(217));
    layer0_outputs(4700) <= inputs(180);
    layer0_outputs(4701) <= (inputs(29)) and not (inputs(36));
    layer0_outputs(4702) <= not(inputs(157));
    layer0_outputs(4703) <= '1';
    layer0_outputs(4704) <= inputs(215);
    layer0_outputs(4705) <= inputs(212);
    layer0_outputs(4706) <= not((inputs(230)) and (inputs(44)));
    layer0_outputs(4707) <= inputs(124);
    layer0_outputs(4708) <= inputs(133);
    layer0_outputs(4709) <= (inputs(113)) and (inputs(123));
    layer0_outputs(4710) <= (inputs(94)) or (inputs(207));
    layer0_outputs(4711) <= not(inputs(150)) or (inputs(60));
    layer0_outputs(4712) <= inputs(141);
    layer0_outputs(4713) <= not(inputs(19));
    layer0_outputs(4714) <= not(inputs(145)) or (inputs(146));
    layer0_outputs(4715) <= (inputs(31)) and not (inputs(44));
    layer0_outputs(4716) <= not((inputs(163)) and (inputs(67)));
    layer0_outputs(4717) <= not(inputs(136)) or (inputs(115));
    layer0_outputs(4718) <= not(inputs(0)) or (inputs(249));
    layer0_outputs(4719) <= not(inputs(104)) or (inputs(93));
    layer0_outputs(4720) <= not(inputs(55)) or (inputs(81));
    layer0_outputs(4721) <= '1';
    layer0_outputs(4722) <= inputs(86);
    layer0_outputs(4723) <= not(inputs(127)) or (inputs(115));
    layer0_outputs(4724) <= not(inputs(167));
    layer0_outputs(4725) <= '1';
    layer0_outputs(4726) <= not((inputs(155)) or (inputs(124)));
    layer0_outputs(4727) <= not((inputs(97)) or (inputs(206)));
    layer0_outputs(4728) <= (inputs(145)) and not (inputs(252));
    layer0_outputs(4729) <= not((inputs(144)) xor (inputs(215)));
    layer0_outputs(4730) <= '1';
    layer0_outputs(4731) <= not(inputs(169));
    layer0_outputs(4732) <= (inputs(236)) xor (inputs(120));
    layer0_outputs(4733) <= (inputs(105)) xor (inputs(16));
    layer0_outputs(4734) <= (inputs(119)) and not (inputs(51));
    layer0_outputs(4735) <= (inputs(202)) and not (inputs(110));
    layer0_outputs(4736) <= (inputs(184)) xor (inputs(129));
    layer0_outputs(4737) <= inputs(165);
    layer0_outputs(4738) <= not(inputs(84)) or (inputs(73));
    layer0_outputs(4739) <= not((inputs(22)) and (inputs(227)));
    layer0_outputs(4740) <= (inputs(141)) and not (inputs(133));
    layer0_outputs(4741) <= not(inputs(92)) or (inputs(252));
    layer0_outputs(4742) <= (inputs(15)) and (inputs(109));
    layer0_outputs(4743) <= inputs(198);
    layer0_outputs(4744) <= inputs(46);
    layer0_outputs(4745) <= (inputs(144)) and not (inputs(83));
    layer0_outputs(4746) <= (inputs(10)) and not (inputs(236));
    layer0_outputs(4747) <= '1';
    layer0_outputs(4748) <= (inputs(251)) and not (inputs(192));
    layer0_outputs(4749) <= not((inputs(119)) or (inputs(77)));
    layer0_outputs(4750) <= '1';
    layer0_outputs(4751) <= not((inputs(222)) xor (inputs(137)));
    layer0_outputs(4752) <= (inputs(72)) and not (inputs(194));
    layer0_outputs(4753) <= not(inputs(25));
    layer0_outputs(4754) <= (inputs(42)) or (inputs(190));
    layer0_outputs(4755) <= (inputs(111)) or (inputs(110));
    layer0_outputs(4756) <= (inputs(72)) and not (inputs(120));
    layer0_outputs(4757) <= not(inputs(166));
    layer0_outputs(4758) <= (inputs(243)) and not (inputs(101));
    layer0_outputs(4759) <= not(inputs(200));
    layer0_outputs(4760) <= not(inputs(181));
    layer0_outputs(4761) <= not((inputs(194)) or (inputs(164)));
    layer0_outputs(4762) <= not(inputs(141)) or (inputs(82));
    layer0_outputs(4763) <= not((inputs(38)) and (inputs(44)));
    layer0_outputs(4764) <= (inputs(162)) or (inputs(55));
    layer0_outputs(4765) <= inputs(107);
    layer0_outputs(4766) <= not(inputs(182)) or (inputs(161));
    layer0_outputs(4767) <= not((inputs(236)) xor (inputs(107)));
    layer0_outputs(4768) <= not(inputs(227)) or (inputs(130));
    layer0_outputs(4769) <= (inputs(207)) and not (inputs(243));
    layer0_outputs(4770) <= (inputs(133)) and not (inputs(242));
    layer0_outputs(4771) <= not(inputs(176));
    layer0_outputs(4772) <= inputs(47);
    layer0_outputs(4773) <= not((inputs(29)) and (inputs(208)));
    layer0_outputs(4774) <= not((inputs(252)) or (inputs(129)));
    layer0_outputs(4775) <= (inputs(59)) and not (inputs(81));
    layer0_outputs(4776) <= inputs(212);
    layer0_outputs(4777) <= inputs(39);
    layer0_outputs(4778) <= (inputs(28)) xor (inputs(149));
    layer0_outputs(4779) <= '1';
    layer0_outputs(4780) <= not(inputs(116));
    layer0_outputs(4781) <= not((inputs(18)) or (inputs(40)));
    layer0_outputs(4782) <= not((inputs(102)) xor (inputs(253)));
    layer0_outputs(4783) <= not((inputs(95)) xor (inputs(144)));
    layer0_outputs(4784) <= (inputs(67)) and (inputs(209));
    layer0_outputs(4785) <= (inputs(177)) and (inputs(50));
    layer0_outputs(4786) <= not(inputs(248));
    layer0_outputs(4787) <= not((inputs(243)) and (inputs(124)));
    layer0_outputs(4788) <= not((inputs(244)) or (inputs(196)));
    layer0_outputs(4789) <= (inputs(167)) or (inputs(17));
    layer0_outputs(4790) <= not((inputs(219)) or (inputs(137)));
    layer0_outputs(4791) <= not(inputs(218)) or (inputs(201));
    layer0_outputs(4792) <= '0';
    layer0_outputs(4793) <= (inputs(85)) or (inputs(228));
    layer0_outputs(4794) <= not((inputs(157)) or (inputs(228)));
    layer0_outputs(4795) <= not(inputs(27)) or (inputs(20));
    layer0_outputs(4796) <= not(inputs(242));
    layer0_outputs(4797) <= (inputs(5)) and not (inputs(83));
    layer0_outputs(4798) <= (inputs(104)) and not (inputs(230));
    layer0_outputs(4799) <= inputs(29);
    layer0_outputs(4800) <= inputs(152);
    layer0_outputs(4801) <= not((inputs(46)) or (inputs(115)));
    layer0_outputs(4802) <= not((inputs(161)) xor (inputs(71)));
    layer0_outputs(4803) <= not(inputs(111));
    layer0_outputs(4804) <= not(inputs(167));
    layer0_outputs(4805) <= not((inputs(165)) or (inputs(57)));
    layer0_outputs(4806) <= (inputs(216)) and not (inputs(221));
    layer0_outputs(4807) <= not((inputs(180)) or (inputs(62)));
    layer0_outputs(4808) <= not(inputs(139)) or (inputs(193));
    layer0_outputs(4809) <= not((inputs(175)) or (inputs(31)));
    layer0_outputs(4810) <= '0';
    layer0_outputs(4811) <= not(inputs(173)) or (inputs(207));
    layer0_outputs(4812) <= not((inputs(229)) or (inputs(106)));
    layer0_outputs(4813) <= not(inputs(70)) or (inputs(237));
    layer0_outputs(4814) <= (inputs(247)) and not (inputs(176));
    layer0_outputs(4815) <= (inputs(16)) and (inputs(50));
    layer0_outputs(4816) <= inputs(201);
    layer0_outputs(4817) <= (inputs(120)) and not (inputs(238));
    layer0_outputs(4818) <= not(inputs(61));
    layer0_outputs(4819) <= inputs(173);
    layer0_outputs(4820) <= not((inputs(134)) xor (inputs(63)));
    layer0_outputs(4821) <= (inputs(64)) and not (inputs(79));
    layer0_outputs(4822) <= inputs(178);
    layer0_outputs(4823) <= not((inputs(149)) xor (inputs(166)));
    layer0_outputs(4824) <= (inputs(115)) or (inputs(112));
    layer0_outputs(4825) <= not((inputs(4)) or (inputs(60)));
    layer0_outputs(4826) <= not((inputs(172)) or (inputs(190)));
    layer0_outputs(4827) <= not((inputs(149)) or (inputs(133)));
    layer0_outputs(4828) <= '0';
    layer0_outputs(4829) <= (inputs(216)) or (inputs(165));
    layer0_outputs(4830) <= (inputs(84)) or (inputs(93));
    layer0_outputs(4831) <= not(inputs(62)) or (inputs(98));
    layer0_outputs(4832) <= '0';
    layer0_outputs(4833) <= not(inputs(37)) or (inputs(65));
    layer0_outputs(4834) <= (inputs(29)) and not (inputs(115));
    layer0_outputs(4835) <= (inputs(167)) xor (inputs(87));
    layer0_outputs(4836) <= '0';
    layer0_outputs(4837) <= not((inputs(68)) and (inputs(70)));
    layer0_outputs(4838) <= inputs(108);
    layer0_outputs(4839) <= not((inputs(126)) xor (inputs(181)));
    layer0_outputs(4840) <= not(inputs(127));
    layer0_outputs(4841) <= inputs(167);
    layer0_outputs(4842) <= inputs(3);
    layer0_outputs(4843) <= not((inputs(28)) xor (inputs(189)));
    layer0_outputs(4844) <= not((inputs(63)) or (inputs(158)));
    layer0_outputs(4845) <= (inputs(247)) and (inputs(34));
    layer0_outputs(4846) <= inputs(145);
    layer0_outputs(4847) <= '0';
    layer0_outputs(4848) <= inputs(13);
    layer0_outputs(4849) <= not((inputs(31)) or (inputs(34)));
    layer0_outputs(4850) <= '1';
    layer0_outputs(4851) <= inputs(188);
    layer0_outputs(4852) <= not((inputs(98)) and (inputs(219)));
    layer0_outputs(4853) <= (inputs(38)) or (inputs(236));
    layer0_outputs(4854) <= (inputs(139)) and (inputs(49));
    layer0_outputs(4855) <= (inputs(95)) xor (inputs(124));
    layer0_outputs(4856) <= not(inputs(182));
    layer0_outputs(4857) <= (inputs(125)) xor (inputs(48));
    layer0_outputs(4858) <= inputs(217);
    layer0_outputs(4859) <= not((inputs(199)) or (inputs(19)));
    layer0_outputs(4860) <= (inputs(110)) and not (inputs(103));
    layer0_outputs(4861) <= (inputs(126)) xor (inputs(166));
    layer0_outputs(4862) <= not((inputs(129)) or (inputs(97)));
    layer0_outputs(4863) <= not((inputs(115)) or (inputs(43)));
    layer0_outputs(4864) <= '1';
    layer0_outputs(4865) <= not(inputs(183)) or (inputs(110));
    layer0_outputs(4866) <= '0';
    layer0_outputs(4867) <= inputs(116);
    layer0_outputs(4868) <= (inputs(109)) and not (inputs(223));
    layer0_outputs(4869) <= '0';
    layer0_outputs(4870) <= (inputs(138)) and (inputs(168));
    layer0_outputs(4871) <= not(inputs(214)) or (inputs(199));
    layer0_outputs(4872) <= inputs(131);
    layer0_outputs(4873) <= not(inputs(12)) or (inputs(135));
    layer0_outputs(4874) <= not(inputs(196));
    layer0_outputs(4875) <= not(inputs(165));
    layer0_outputs(4876) <= not((inputs(139)) xor (inputs(179)));
    layer0_outputs(4877) <= (inputs(21)) and (inputs(177));
    layer0_outputs(4878) <= not((inputs(3)) or (inputs(74)));
    layer0_outputs(4879) <= (inputs(23)) and not (inputs(64));
    layer0_outputs(4880) <= inputs(201);
    layer0_outputs(4881) <= (inputs(91)) or (inputs(93));
    layer0_outputs(4882) <= (inputs(178)) xor (inputs(209));
    layer0_outputs(4883) <= (inputs(65)) and not (inputs(121));
    layer0_outputs(4884) <= inputs(149);
    layer0_outputs(4885) <= not((inputs(251)) xor (inputs(83)));
    layer0_outputs(4886) <= inputs(192);
    layer0_outputs(4887) <= (inputs(255)) and (inputs(254));
    layer0_outputs(4888) <= not(inputs(236));
    layer0_outputs(4889) <= '1';
    layer0_outputs(4890) <= (inputs(204)) and not (inputs(238));
    layer0_outputs(4891) <= (inputs(209)) and not (inputs(242));
    layer0_outputs(4892) <= not((inputs(5)) or (inputs(55)));
    layer0_outputs(4893) <= '0';
    layer0_outputs(4894) <= not(inputs(19));
    layer0_outputs(4895) <= '1';
    layer0_outputs(4896) <= not((inputs(70)) or (inputs(61)));
    layer0_outputs(4897) <= (inputs(122)) and not (inputs(170));
    layer0_outputs(4898) <= not(inputs(215)) or (inputs(209));
    layer0_outputs(4899) <= not(inputs(190)) or (inputs(157));
    layer0_outputs(4900) <= (inputs(245)) or (inputs(186));
    layer0_outputs(4901) <= not(inputs(152));
    layer0_outputs(4902) <= not(inputs(113));
    layer0_outputs(4903) <= (inputs(70)) and not (inputs(174));
    layer0_outputs(4904) <= not((inputs(143)) xor (inputs(151)));
    layer0_outputs(4905) <= not(inputs(53));
    layer0_outputs(4906) <= not(inputs(182));
    layer0_outputs(4907) <= (inputs(192)) and not (inputs(21));
    layer0_outputs(4908) <= not(inputs(160)) or (inputs(89));
    layer0_outputs(4909) <= not(inputs(240));
    layer0_outputs(4910) <= inputs(113);
    layer0_outputs(4911) <= inputs(151);
    layer0_outputs(4912) <= not((inputs(156)) and (inputs(127)));
    layer0_outputs(4913) <= (inputs(221)) and not (inputs(88));
    layer0_outputs(4914) <= not(inputs(137)) or (inputs(163));
    layer0_outputs(4915) <= not((inputs(212)) and (inputs(34)));
    layer0_outputs(4916) <= (inputs(166)) and not (inputs(228));
    layer0_outputs(4917) <= inputs(192);
    layer0_outputs(4918) <= not(inputs(5));
    layer0_outputs(4919) <= '1';
    layer0_outputs(4920) <= not(inputs(222)) or (inputs(103));
    layer0_outputs(4921) <= not(inputs(212)) or (inputs(52));
    layer0_outputs(4922) <= not((inputs(177)) or (inputs(139)));
    layer0_outputs(4923) <= (inputs(23)) or (inputs(95));
    layer0_outputs(4924) <= not((inputs(228)) or (inputs(146)));
    layer0_outputs(4925) <= (inputs(172)) and (inputs(17));
    layer0_outputs(4926) <= not(inputs(47)) or (inputs(214));
    layer0_outputs(4927) <= not(inputs(120));
    layer0_outputs(4928) <= not(inputs(224));
    layer0_outputs(4929) <= not((inputs(148)) xor (inputs(222)));
    layer0_outputs(4930) <= not((inputs(11)) and (inputs(219)));
    layer0_outputs(4931) <= not(inputs(201));
    layer0_outputs(4932) <= not((inputs(126)) and (inputs(73)));
    layer0_outputs(4933) <= not(inputs(65)) or (inputs(232));
    layer0_outputs(4934) <= not(inputs(142));
    layer0_outputs(4935) <= not(inputs(89));
    layer0_outputs(4936) <= (inputs(161)) xor (inputs(7));
    layer0_outputs(4937) <= inputs(188);
    layer0_outputs(4938) <= not((inputs(10)) and (inputs(83)));
    layer0_outputs(4939) <= not(inputs(76));
    layer0_outputs(4940) <= not((inputs(178)) or (inputs(181)));
    layer0_outputs(4941) <= (inputs(178)) and not (inputs(218));
    layer0_outputs(4942) <= not(inputs(170));
    layer0_outputs(4943) <= not(inputs(35));
    layer0_outputs(4944) <= (inputs(170)) or (inputs(68));
    layer0_outputs(4945) <= inputs(217);
    layer0_outputs(4946) <= (inputs(110)) xor (inputs(80));
    layer0_outputs(4947) <= not(inputs(177));
    layer0_outputs(4948) <= (inputs(45)) and not (inputs(161));
    layer0_outputs(4949) <= not((inputs(189)) or (inputs(217)));
    layer0_outputs(4950) <= (inputs(73)) or (inputs(128));
    layer0_outputs(4951) <= not(inputs(7));
    layer0_outputs(4952) <= not((inputs(146)) and (inputs(163)));
    layer0_outputs(4953) <= (inputs(71)) or (inputs(87));
    layer0_outputs(4954) <= not((inputs(48)) xor (inputs(127)));
    layer0_outputs(4955) <= (inputs(155)) or (inputs(107));
    layer0_outputs(4956) <= not(inputs(65));
    layer0_outputs(4957) <= not((inputs(117)) xor (inputs(132)));
    layer0_outputs(4958) <= not(inputs(57)) or (inputs(88));
    layer0_outputs(4959) <= (inputs(234)) and (inputs(46));
    layer0_outputs(4960) <= (inputs(190)) and (inputs(50));
    layer0_outputs(4961) <= not(inputs(164));
    layer0_outputs(4962) <= (inputs(189)) xor (inputs(88));
    layer0_outputs(4963) <= (inputs(4)) and (inputs(198));
    layer0_outputs(4964) <= not((inputs(178)) xor (inputs(54)));
    layer0_outputs(4965) <= not((inputs(0)) xor (inputs(151)));
    layer0_outputs(4966) <= (inputs(168)) and not (inputs(221));
    layer0_outputs(4967) <= (inputs(237)) and not (inputs(17));
    layer0_outputs(4968) <= not(inputs(146));
    layer0_outputs(4969) <= not(inputs(208)) or (inputs(141));
    layer0_outputs(4970) <= (inputs(202)) and not (inputs(141));
    layer0_outputs(4971) <= not(inputs(86));
    layer0_outputs(4972) <= not((inputs(217)) or (inputs(201)));
    layer0_outputs(4973) <= not((inputs(184)) or (inputs(38)));
    layer0_outputs(4974) <= not((inputs(64)) or (inputs(70)));
    layer0_outputs(4975) <= (inputs(93)) and (inputs(27));
    layer0_outputs(4976) <= (inputs(65)) and not (inputs(52));
    layer0_outputs(4977) <= inputs(61);
    layer0_outputs(4978) <= (inputs(65)) and not (inputs(226));
    layer0_outputs(4979) <= (inputs(82)) and not (inputs(9));
    layer0_outputs(4980) <= not(inputs(146));
    layer0_outputs(4981) <= (inputs(139)) xor (inputs(112));
    layer0_outputs(4982) <= not((inputs(242)) xor (inputs(193)));
    layer0_outputs(4983) <= inputs(63);
    layer0_outputs(4984) <= (inputs(211)) xor (inputs(200));
    layer0_outputs(4985) <= inputs(59);
    layer0_outputs(4986) <= (inputs(143)) and not (inputs(191));
    layer0_outputs(4987) <= inputs(100);
    layer0_outputs(4988) <= (inputs(212)) or (inputs(72));
    layer0_outputs(4989) <= not((inputs(196)) xor (inputs(228)));
    layer0_outputs(4990) <= (inputs(162)) and (inputs(114));
    layer0_outputs(4991) <= (inputs(90)) or (inputs(19));
    layer0_outputs(4992) <= (inputs(93)) and not (inputs(227));
    layer0_outputs(4993) <= (inputs(9)) xor (inputs(217));
    layer0_outputs(4994) <= (inputs(208)) or (inputs(84));
    layer0_outputs(4995) <= not(inputs(149)) or (inputs(236));
    layer0_outputs(4996) <= not(inputs(55)) or (inputs(27));
    layer0_outputs(4997) <= (inputs(108)) and (inputs(59));
    layer0_outputs(4998) <= '0';
    layer0_outputs(4999) <= inputs(170);
    layer0_outputs(5000) <= not((inputs(251)) xor (inputs(161)));
    layer0_outputs(5001) <= '0';
    layer0_outputs(5002) <= (inputs(94)) and not (inputs(25));
    layer0_outputs(5003) <= not(inputs(71));
    layer0_outputs(5004) <= not((inputs(106)) or (inputs(251)));
    layer0_outputs(5005) <= '1';
    layer0_outputs(5006) <= not(inputs(206)) or (inputs(125));
    layer0_outputs(5007) <= not(inputs(182));
    layer0_outputs(5008) <= not(inputs(88)) or (inputs(91));
    layer0_outputs(5009) <= inputs(152);
    layer0_outputs(5010) <= not((inputs(133)) or (inputs(117)));
    layer0_outputs(5011) <= (inputs(176)) and (inputs(222));
    layer0_outputs(5012) <= (inputs(122)) or (inputs(145));
    layer0_outputs(5013) <= (inputs(223)) xor (inputs(45));
    layer0_outputs(5014) <= '1';
    layer0_outputs(5015) <= not((inputs(249)) or (inputs(252)));
    layer0_outputs(5016) <= not(inputs(6)) or (inputs(28));
    layer0_outputs(5017) <= not((inputs(151)) or (inputs(164)));
    layer0_outputs(5018) <= (inputs(55)) xor (inputs(146));
    layer0_outputs(5019) <= not(inputs(55));
    layer0_outputs(5020) <= (inputs(156)) or (inputs(57));
    layer0_outputs(5021) <= inputs(12);
    layer0_outputs(5022) <= (inputs(180)) and not (inputs(97));
    layer0_outputs(5023) <= not(inputs(27)) or (inputs(224));
    layer0_outputs(5024) <= not(inputs(164)) or (inputs(234));
    layer0_outputs(5025) <= inputs(43);
    layer0_outputs(5026) <= not(inputs(215)) or (inputs(177));
    layer0_outputs(5027) <= not(inputs(90)) or (inputs(43));
    layer0_outputs(5028) <= not(inputs(167)) or (inputs(82));
    layer0_outputs(5029) <= inputs(145);
    layer0_outputs(5030) <= not((inputs(50)) or (inputs(205)));
    layer0_outputs(5031) <= (inputs(202)) and (inputs(84));
    layer0_outputs(5032) <= (inputs(121)) and not (inputs(158));
    layer0_outputs(5033) <= (inputs(96)) and not (inputs(168));
    layer0_outputs(5034) <= not(inputs(212)) or (inputs(233));
    layer0_outputs(5035) <= (inputs(255)) and not (inputs(31));
    layer0_outputs(5036) <= (inputs(158)) and not (inputs(234));
    layer0_outputs(5037) <= not(inputs(167));
    layer0_outputs(5038) <= not((inputs(167)) or (inputs(242)));
    layer0_outputs(5039) <= inputs(20);
    layer0_outputs(5040) <= (inputs(162)) xor (inputs(188));
    layer0_outputs(5041) <= not(inputs(76));
    layer0_outputs(5042) <= (inputs(31)) and not (inputs(248));
    layer0_outputs(5043) <= (inputs(252)) and not (inputs(157));
    layer0_outputs(5044) <= inputs(27);
    layer0_outputs(5045) <= not(inputs(85));
    layer0_outputs(5046) <= inputs(179);
    layer0_outputs(5047) <= '0';
    layer0_outputs(5048) <= not(inputs(100)) or (inputs(4));
    layer0_outputs(5049) <= (inputs(162)) or (inputs(189));
    layer0_outputs(5050) <= '1';
    layer0_outputs(5051) <= not(inputs(169));
    layer0_outputs(5052) <= not(inputs(167)) or (inputs(243));
    layer0_outputs(5053) <= (inputs(101)) and not (inputs(200));
    layer0_outputs(5054) <= not((inputs(6)) or (inputs(223)));
    layer0_outputs(5055) <= '1';
    layer0_outputs(5056) <= '0';
    layer0_outputs(5057) <= not((inputs(100)) or (inputs(103)));
    layer0_outputs(5058) <= not(inputs(211)) or (inputs(113));
    layer0_outputs(5059) <= not(inputs(164));
    layer0_outputs(5060) <= inputs(82);
    layer0_outputs(5061) <= not(inputs(212));
    layer0_outputs(5062) <= not(inputs(166));
    layer0_outputs(5063) <= not(inputs(102)) or (inputs(78));
    layer0_outputs(5064) <= not((inputs(109)) or (inputs(142)));
    layer0_outputs(5065) <= (inputs(210)) and not (inputs(195));
    layer0_outputs(5066) <= (inputs(30)) or (inputs(240));
    layer0_outputs(5067) <= not((inputs(12)) or (inputs(178)));
    layer0_outputs(5068) <= (inputs(67)) and (inputs(133));
    layer0_outputs(5069) <= inputs(105);
    layer0_outputs(5070) <= not(inputs(56)) or (inputs(208));
    layer0_outputs(5071) <= (inputs(174)) xor (inputs(236));
    layer0_outputs(5072) <= not((inputs(150)) or (inputs(134)));
    layer0_outputs(5073) <= not(inputs(168)) or (inputs(181));
    layer0_outputs(5074) <= not(inputs(176)) or (inputs(75));
    layer0_outputs(5075) <= inputs(58);
    layer0_outputs(5076) <= not(inputs(137)) or (inputs(44));
    layer0_outputs(5077) <= not(inputs(26)) or (inputs(31));
    layer0_outputs(5078) <= (inputs(121)) and not (inputs(148));
    layer0_outputs(5079) <= '1';
    layer0_outputs(5080) <= not((inputs(111)) xor (inputs(212)));
    layer0_outputs(5081) <= not((inputs(170)) and (inputs(12)));
    layer0_outputs(5082) <= '1';
    layer0_outputs(5083) <= not(inputs(68));
    layer0_outputs(5084) <= not(inputs(166)) or (inputs(146));
    layer0_outputs(5085) <= not(inputs(190));
    layer0_outputs(5086) <= inputs(140);
    layer0_outputs(5087) <= (inputs(133)) xor (inputs(233));
    layer0_outputs(5088) <= (inputs(98)) and not (inputs(188));
    layer0_outputs(5089) <= not(inputs(72));
    layer0_outputs(5090) <= not(inputs(34));
    layer0_outputs(5091) <= not((inputs(164)) or (inputs(205)));
    layer0_outputs(5092) <= '1';
    layer0_outputs(5093) <= (inputs(179)) xor (inputs(149));
    layer0_outputs(5094) <= (inputs(31)) or (inputs(221));
    layer0_outputs(5095) <= (inputs(223)) xor (inputs(154));
    layer0_outputs(5096) <= not((inputs(163)) or (inputs(94)));
    layer0_outputs(5097) <= not(inputs(192));
    layer0_outputs(5098) <= (inputs(65)) and not (inputs(160));
    layer0_outputs(5099) <= (inputs(55)) and not (inputs(243));
    layer0_outputs(5100) <= (inputs(151)) and not (inputs(140));
    layer0_outputs(5101) <= (inputs(68)) and (inputs(126));
    layer0_outputs(5102) <= (inputs(56)) and not (inputs(147));
    layer0_outputs(5103) <= (inputs(55)) and (inputs(165));
    layer0_outputs(5104) <= inputs(56);
    layer0_outputs(5105) <= (inputs(69)) xor (inputs(69));
    layer0_outputs(5106) <= (inputs(86)) or (inputs(238));
    layer0_outputs(5107) <= (inputs(196)) or (inputs(228));
    layer0_outputs(5108) <= not(inputs(169));
    layer0_outputs(5109) <= not((inputs(208)) and (inputs(101)));
    layer0_outputs(5110) <= not(inputs(195)) or (inputs(67));
    layer0_outputs(5111) <= not(inputs(162));
    layer0_outputs(5112) <= (inputs(251)) and not (inputs(5));
    layer0_outputs(5113) <= '0';
    layer0_outputs(5114) <= not(inputs(65));
    layer0_outputs(5115) <= not((inputs(85)) xor (inputs(34)));
    layer0_outputs(5116) <= not(inputs(228));
    layer0_outputs(5117) <= not(inputs(71));
    layer0_outputs(5118) <= inputs(124);
    layer0_outputs(5119) <= not((inputs(200)) xor (inputs(175)));
    layer0_outputs(5120) <= not(inputs(151)) or (inputs(144));
    layer0_outputs(5121) <= inputs(147);
    layer0_outputs(5122) <= not(inputs(175));
    layer0_outputs(5123) <= (inputs(215)) and not (inputs(95));
    layer0_outputs(5124) <= inputs(27);
    layer0_outputs(5125) <= not(inputs(80));
    layer0_outputs(5126) <= (inputs(185)) and not (inputs(128));
    layer0_outputs(5127) <= inputs(150);
    layer0_outputs(5128) <= inputs(85);
    layer0_outputs(5129) <= (inputs(208)) xor (inputs(157));
    layer0_outputs(5130) <= not(inputs(199));
    layer0_outputs(5131) <= inputs(186);
    layer0_outputs(5132) <= inputs(179);
    layer0_outputs(5133) <= inputs(183);
    layer0_outputs(5134) <= (inputs(192)) or (inputs(65));
    layer0_outputs(5135) <= not(inputs(208)) or (inputs(208));
    layer0_outputs(5136) <= not((inputs(113)) xor (inputs(114)));
    layer0_outputs(5137) <= inputs(11);
    layer0_outputs(5138) <= not((inputs(27)) and (inputs(224)));
    layer0_outputs(5139) <= not(inputs(209)) or (inputs(189));
    layer0_outputs(5140) <= '1';
    layer0_outputs(5141) <= not(inputs(106)) or (inputs(26));
    layer0_outputs(5142) <= not((inputs(4)) xor (inputs(248)));
    layer0_outputs(5143) <= not((inputs(240)) xor (inputs(51)));
    layer0_outputs(5144) <= (inputs(220)) or (inputs(193));
    layer0_outputs(5145) <= not((inputs(183)) and (inputs(154)));
    layer0_outputs(5146) <= inputs(127);
    layer0_outputs(5147) <= not(inputs(147));
    layer0_outputs(5148) <= (inputs(24)) xor (inputs(79));
    layer0_outputs(5149) <= (inputs(24)) or (inputs(35));
    layer0_outputs(5150) <= (inputs(226)) xor (inputs(67));
    layer0_outputs(5151) <= '1';
    layer0_outputs(5152) <= inputs(136);
    layer0_outputs(5153) <= inputs(175);
    layer0_outputs(5154) <= (inputs(13)) or (inputs(190));
    layer0_outputs(5155) <= not(inputs(91));
    layer0_outputs(5156) <= (inputs(213)) or (inputs(163));
    layer0_outputs(5157) <= inputs(232);
    layer0_outputs(5158) <= not(inputs(120));
    layer0_outputs(5159) <= not(inputs(36));
    layer0_outputs(5160) <= (inputs(219)) or (inputs(40));
    layer0_outputs(5161) <= (inputs(42)) and not (inputs(68));
    layer0_outputs(5162) <= (inputs(101)) and not (inputs(220));
    layer0_outputs(5163) <= not((inputs(201)) xor (inputs(1)));
    layer0_outputs(5164) <= inputs(229);
    layer0_outputs(5165) <= not(inputs(66)) or (inputs(4));
    layer0_outputs(5166) <= (inputs(143)) xor (inputs(119));
    layer0_outputs(5167) <= (inputs(8)) and not (inputs(90));
    layer0_outputs(5168) <= (inputs(90)) and not (inputs(141));
    layer0_outputs(5169) <= not((inputs(5)) and (inputs(223)));
    layer0_outputs(5170) <= not((inputs(70)) xor (inputs(77)));
    layer0_outputs(5171) <= (inputs(42)) or (inputs(251));
    layer0_outputs(5172) <= not((inputs(108)) or (inputs(182)));
    layer0_outputs(5173) <= (inputs(109)) or (inputs(192));
    layer0_outputs(5174) <= not(inputs(152));
    layer0_outputs(5175) <= not(inputs(94)) or (inputs(250));
    layer0_outputs(5176) <= not(inputs(41)) or (inputs(250));
    layer0_outputs(5177) <= inputs(172);
    layer0_outputs(5178) <= not((inputs(255)) xor (inputs(151)));
    layer0_outputs(5179) <= not((inputs(82)) or (inputs(161)));
    layer0_outputs(5180) <= not(inputs(255));
    layer0_outputs(5181) <= inputs(16);
    layer0_outputs(5182) <= not((inputs(242)) or (inputs(171)));
    layer0_outputs(5183) <= inputs(198);
    layer0_outputs(5184) <= (inputs(180)) or (inputs(42));
    layer0_outputs(5185) <= (inputs(132)) and not (inputs(174));
    layer0_outputs(5186) <= inputs(205);
    layer0_outputs(5187) <= (inputs(69)) and not (inputs(49));
    layer0_outputs(5188) <= not((inputs(114)) xor (inputs(167)));
    layer0_outputs(5189) <= not((inputs(43)) or (inputs(135)));
    layer0_outputs(5190) <= (inputs(19)) xor (inputs(32));
    layer0_outputs(5191) <= not(inputs(175)) or (inputs(69));
    layer0_outputs(5192) <= not(inputs(253)) or (inputs(226));
    layer0_outputs(5193) <= inputs(90);
    layer0_outputs(5194) <= not(inputs(132));
    layer0_outputs(5195) <= '1';
    layer0_outputs(5196) <= not((inputs(187)) xor (inputs(154)));
    layer0_outputs(5197) <= not((inputs(2)) xor (inputs(178)));
    layer0_outputs(5198) <= not((inputs(54)) or (inputs(207)));
    layer0_outputs(5199) <= not((inputs(170)) xor (inputs(217)));
    layer0_outputs(5200) <= (inputs(109)) and not (inputs(244));
    layer0_outputs(5201) <= not((inputs(125)) and (inputs(92)));
    layer0_outputs(5202) <= not((inputs(217)) or (inputs(92)));
    layer0_outputs(5203) <= inputs(102);
    layer0_outputs(5204) <= inputs(197);
    layer0_outputs(5205) <= not((inputs(13)) xor (inputs(42)));
    layer0_outputs(5206) <= not(inputs(69)) or (inputs(59));
    layer0_outputs(5207) <= not((inputs(48)) or (inputs(147)));
    layer0_outputs(5208) <= (inputs(152)) and not (inputs(210));
    layer0_outputs(5209) <= (inputs(174)) or (inputs(229));
    layer0_outputs(5210) <= '0';
    layer0_outputs(5211) <= not(inputs(106)) or (inputs(97));
    layer0_outputs(5212) <= (inputs(183)) and not (inputs(236));
    layer0_outputs(5213) <= (inputs(94)) and not (inputs(144));
    layer0_outputs(5214) <= (inputs(154)) and (inputs(217));
    layer0_outputs(5215) <= not(inputs(168)) or (inputs(194));
    layer0_outputs(5216) <= inputs(167);
    layer0_outputs(5217) <= (inputs(167)) or (inputs(128));
    layer0_outputs(5218) <= not((inputs(113)) or (inputs(217)));
    layer0_outputs(5219) <= inputs(89);
    layer0_outputs(5220) <= inputs(120);
    layer0_outputs(5221) <= inputs(33);
    layer0_outputs(5222) <= not(inputs(69));
    layer0_outputs(5223) <= not((inputs(132)) or (inputs(181)));
    layer0_outputs(5224) <= (inputs(161)) xor (inputs(188));
    layer0_outputs(5225) <= inputs(239);
    layer0_outputs(5226) <= inputs(153);
    layer0_outputs(5227) <= not((inputs(86)) or (inputs(160)));
    layer0_outputs(5228) <= '0';
    layer0_outputs(5229) <= inputs(173);
    layer0_outputs(5230) <= inputs(40);
    layer0_outputs(5231) <= not((inputs(137)) or (inputs(227)));
    layer0_outputs(5232) <= not(inputs(33));
    layer0_outputs(5233) <= (inputs(11)) and (inputs(29));
    layer0_outputs(5234) <= not((inputs(190)) and (inputs(162)));
    layer0_outputs(5235) <= (inputs(184)) and (inputs(142));
    layer0_outputs(5236) <= not(inputs(33)) or (inputs(2));
    layer0_outputs(5237) <= '1';
    layer0_outputs(5238) <= (inputs(76)) xor (inputs(238));
    layer0_outputs(5239) <= (inputs(22)) xor (inputs(175));
    layer0_outputs(5240) <= inputs(53);
    layer0_outputs(5241) <= '1';
    layer0_outputs(5242) <= inputs(25);
    layer0_outputs(5243) <= (inputs(131)) xor (inputs(118));
    layer0_outputs(5244) <= inputs(51);
    layer0_outputs(5245) <= (inputs(210)) and (inputs(75));
    layer0_outputs(5246) <= not(inputs(6)) or (inputs(155));
    layer0_outputs(5247) <= not((inputs(12)) or (inputs(96)));
    layer0_outputs(5248) <= inputs(48);
    layer0_outputs(5249) <= '0';
    layer0_outputs(5250) <= '0';
    layer0_outputs(5251) <= (inputs(3)) xor (inputs(17));
    layer0_outputs(5252) <= '1';
    layer0_outputs(5253) <= (inputs(16)) and not (inputs(45));
    layer0_outputs(5254) <= inputs(87);
    layer0_outputs(5255) <= not(inputs(134)) or (inputs(33));
    layer0_outputs(5256) <= not((inputs(216)) xor (inputs(226)));
    layer0_outputs(5257) <= '0';
    layer0_outputs(5258) <= not(inputs(196)) or (inputs(135));
    layer0_outputs(5259) <= not(inputs(206)) or (inputs(43));
    layer0_outputs(5260) <= not(inputs(177));
    layer0_outputs(5261) <= (inputs(132)) xor (inputs(82));
    layer0_outputs(5262) <= inputs(240);
    layer0_outputs(5263) <= inputs(81);
    layer0_outputs(5264) <= not(inputs(45)) or (inputs(33));
    layer0_outputs(5265) <= not(inputs(67)) or (inputs(237));
    layer0_outputs(5266) <= not((inputs(220)) or (inputs(83)));
    layer0_outputs(5267) <= '1';
    layer0_outputs(5268) <= (inputs(196)) and not (inputs(165));
    layer0_outputs(5269) <= (inputs(82)) xor (inputs(96));
    layer0_outputs(5270) <= not(inputs(110));
    layer0_outputs(5271) <= not(inputs(98));
    layer0_outputs(5272) <= not(inputs(254)) or (inputs(14));
    layer0_outputs(5273) <= (inputs(46)) or (inputs(120));
    layer0_outputs(5274) <= not((inputs(165)) or (inputs(195)));
    layer0_outputs(5275) <= not((inputs(45)) xor (inputs(40)));
    layer0_outputs(5276) <= (inputs(22)) and not (inputs(191));
    layer0_outputs(5277) <= not(inputs(52)) or (inputs(219));
    layer0_outputs(5278) <= not(inputs(53));
    layer0_outputs(5279) <= not(inputs(232)) or (inputs(83));
    layer0_outputs(5280) <= (inputs(236)) and not (inputs(5));
    layer0_outputs(5281) <= not(inputs(29));
    layer0_outputs(5282) <= (inputs(119)) and not (inputs(0));
    layer0_outputs(5283) <= (inputs(136)) or (inputs(10));
    layer0_outputs(5284) <= (inputs(246)) or (inputs(60));
    layer0_outputs(5285) <= not(inputs(147)) or (inputs(96));
    layer0_outputs(5286) <= (inputs(71)) and not (inputs(1));
    layer0_outputs(5287) <= (inputs(139)) xor (inputs(129));
    layer0_outputs(5288) <= inputs(1);
    layer0_outputs(5289) <= '1';
    layer0_outputs(5290) <= not(inputs(60));
    layer0_outputs(5291) <= inputs(7);
    layer0_outputs(5292) <= (inputs(136)) and not (inputs(252));
    layer0_outputs(5293) <= not((inputs(238)) or (inputs(100)));
    layer0_outputs(5294) <= not((inputs(108)) or (inputs(140)));
    layer0_outputs(5295) <= (inputs(180)) and not (inputs(138));
    layer0_outputs(5296) <= not((inputs(153)) or (inputs(42)));
    layer0_outputs(5297) <= (inputs(194)) xor (inputs(20));
    layer0_outputs(5298) <= inputs(56);
    layer0_outputs(5299) <= (inputs(182)) or (inputs(47));
    layer0_outputs(5300) <= not(inputs(7));
    layer0_outputs(5301) <= inputs(115);
    layer0_outputs(5302) <= not(inputs(85));
    layer0_outputs(5303) <= (inputs(134)) and not (inputs(83));
    layer0_outputs(5304) <= not(inputs(93)) or (inputs(198));
    layer0_outputs(5305) <= not((inputs(24)) or (inputs(39)));
    layer0_outputs(5306) <= (inputs(189)) or (inputs(196));
    layer0_outputs(5307) <= inputs(139);
    layer0_outputs(5308) <= not(inputs(126)) or (inputs(73));
    layer0_outputs(5309) <= (inputs(26)) xor (inputs(192));
    layer0_outputs(5310) <= '0';
    layer0_outputs(5311) <= '1';
    layer0_outputs(5312) <= (inputs(144)) and not (inputs(255));
    layer0_outputs(5313) <= not((inputs(188)) and (inputs(143)));
    layer0_outputs(5314) <= not((inputs(107)) or (inputs(138)));
    layer0_outputs(5315) <= '0';
    layer0_outputs(5316) <= (inputs(21)) or (inputs(54));
    layer0_outputs(5317) <= (inputs(79)) and not (inputs(232));
    layer0_outputs(5318) <= not((inputs(210)) and (inputs(44)));
    layer0_outputs(5319) <= not(inputs(234));
    layer0_outputs(5320) <= not(inputs(160));
    layer0_outputs(5321) <= inputs(125);
    layer0_outputs(5322) <= not((inputs(78)) xor (inputs(61)));
    layer0_outputs(5323) <= (inputs(214)) and not (inputs(8));
    layer0_outputs(5324) <= '1';
    layer0_outputs(5325) <= not(inputs(92));
    layer0_outputs(5326) <= inputs(208);
    layer0_outputs(5327) <= '1';
    layer0_outputs(5328) <= inputs(151);
    layer0_outputs(5329) <= inputs(27);
    layer0_outputs(5330) <= (inputs(183)) and not (inputs(171));
    layer0_outputs(5331) <= not(inputs(75));
    layer0_outputs(5332) <= (inputs(7)) or (inputs(77));
    layer0_outputs(5333) <= '0';
    layer0_outputs(5334) <= (inputs(180)) and not (inputs(235));
    layer0_outputs(5335) <= '0';
    layer0_outputs(5336) <= not(inputs(87)) or (inputs(146));
    layer0_outputs(5337) <= not(inputs(90));
    layer0_outputs(5338) <= (inputs(184)) and not (inputs(53));
    layer0_outputs(5339) <= (inputs(211)) and not (inputs(98));
    layer0_outputs(5340) <= (inputs(63)) or (inputs(225));
    layer0_outputs(5341) <= inputs(120);
    layer0_outputs(5342) <= (inputs(57)) and not (inputs(135));
    layer0_outputs(5343) <= (inputs(85)) and not (inputs(60));
    layer0_outputs(5344) <= inputs(198);
    layer0_outputs(5345) <= not(inputs(182)) or (inputs(206));
    layer0_outputs(5346) <= not(inputs(119)) or (inputs(240));
    layer0_outputs(5347) <= inputs(74);
    layer0_outputs(5348) <= (inputs(169)) or (inputs(31));
    layer0_outputs(5349) <= (inputs(241)) and (inputs(194));
    layer0_outputs(5350) <= not(inputs(205));
    layer0_outputs(5351) <= inputs(249);
    layer0_outputs(5352) <= not((inputs(211)) xor (inputs(238)));
    layer0_outputs(5353) <= not((inputs(203)) or (inputs(146)));
    layer0_outputs(5354) <= (inputs(107)) and (inputs(1));
    layer0_outputs(5355) <= not((inputs(77)) and (inputs(242)));
    layer0_outputs(5356) <= not((inputs(62)) xor (inputs(147)));
    layer0_outputs(5357) <= inputs(71);
    layer0_outputs(5358) <= (inputs(40)) or (inputs(120));
    layer0_outputs(5359) <= inputs(136);
    layer0_outputs(5360) <= not(inputs(152)) or (inputs(133));
    layer0_outputs(5361) <= not(inputs(92)) or (inputs(254));
    layer0_outputs(5362) <= (inputs(7)) or (inputs(211));
    layer0_outputs(5363) <= not(inputs(213));
    layer0_outputs(5364) <= (inputs(16)) and not (inputs(96));
    layer0_outputs(5365) <= '0';
    layer0_outputs(5366) <= not(inputs(207)) or (inputs(95));
    layer0_outputs(5367) <= not((inputs(206)) xor (inputs(148)));
    layer0_outputs(5368) <= not((inputs(169)) xor (inputs(67)));
    layer0_outputs(5369) <= not(inputs(117)) or (inputs(136));
    layer0_outputs(5370) <= inputs(17);
    layer0_outputs(5371) <= (inputs(120)) and not (inputs(92));
    layer0_outputs(5372) <= not((inputs(197)) xor (inputs(182)));
    layer0_outputs(5373) <= inputs(121);
    layer0_outputs(5374) <= (inputs(66)) or (inputs(57));
    layer0_outputs(5375) <= (inputs(32)) or (inputs(216));
    layer0_outputs(5376) <= not((inputs(250)) and (inputs(242)));
    layer0_outputs(5377) <= not(inputs(3)) or (inputs(127));
    layer0_outputs(5378) <= not((inputs(129)) or (inputs(194)));
    layer0_outputs(5379) <= inputs(138);
    layer0_outputs(5380) <= not(inputs(82)) or (inputs(223));
    layer0_outputs(5381) <= (inputs(174)) or (inputs(197));
    layer0_outputs(5382) <= '1';
    layer0_outputs(5383) <= not((inputs(92)) or (inputs(74)));
    layer0_outputs(5384) <= not((inputs(21)) and (inputs(204)));
    layer0_outputs(5385) <= '0';
    layer0_outputs(5386) <= inputs(245);
    layer0_outputs(5387) <= inputs(216);
    layer0_outputs(5388) <= (inputs(145)) or (inputs(200));
    layer0_outputs(5389) <= (inputs(60)) xor (inputs(46));
    layer0_outputs(5390) <= not(inputs(215));
    layer0_outputs(5391) <= not((inputs(240)) and (inputs(25)));
    layer0_outputs(5392) <= inputs(41);
    layer0_outputs(5393) <= (inputs(5)) and (inputs(203));
    layer0_outputs(5394) <= not((inputs(41)) xor (inputs(23)));
    layer0_outputs(5395) <= (inputs(144)) and not (inputs(234));
    layer0_outputs(5396) <= inputs(86);
    layer0_outputs(5397) <= not(inputs(165));
    layer0_outputs(5398) <= not((inputs(255)) or (inputs(53)));
    layer0_outputs(5399) <= not((inputs(237)) xor (inputs(213)));
    layer0_outputs(5400) <= not((inputs(188)) or (inputs(22)));
    layer0_outputs(5401) <= (inputs(120)) and not (inputs(85));
    layer0_outputs(5402) <= not((inputs(3)) or (inputs(213)));
    layer0_outputs(5403) <= not((inputs(93)) or (inputs(131)));
    layer0_outputs(5404) <= not((inputs(48)) and (inputs(102)));
    layer0_outputs(5405) <= (inputs(241)) or (inputs(24));
    layer0_outputs(5406) <= not((inputs(177)) xor (inputs(173)));
    layer0_outputs(5407) <= not(inputs(113)) or (inputs(126));
    layer0_outputs(5408) <= '1';
    layer0_outputs(5409) <= inputs(216);
    layer0_outputs(5410) <= inputs(40);
    layer0_outputs(5411) <= not((inputs(219)) and (inputs(112)));
    layer0_outputs(5412) <= '1';
    layer0_outputs(5413) <= inputs(205);
    layer0_outputs(5414) <= '1';
    layer0_outputs(5415) <= (inputs(85)) and not (inputs(140));
    layer0_outputs(5416) <= inputs(181);
    layer0_outputs(5417) <= (inputs(234)) xor (inputs(40));
    layer0_outputs(5418) <= (inputs(198)) and not (inputs(25));
    layer0_outputs(5419) <= (inputs(109)) or (inputs(216));
    layer0_outputs(5420) <= (inputs(142)) or (inputs(167));
    layer0_outputs(5421) <= '0';
    layer0_outputs(5422) <= (inputs(205)) and not (inputs(157));
    layer0_outputs(5423) <= not(inputs(209));
    layer0_outputs(5424) <= inputs(55);
    layer0_outputs(5425) <= inputs(167);
    layer0_outputs(5426) <= (inputs(178)) and not (inputs(89));
    layer0_outputs(5427) <= not(inputs(216)) or (inputs(148));
    layer0_outputs(5428) <= not(inputs(60)) or (inputs(248));
    layer0_outputs(5429) <= not(inputs(89)) or (inputs(118));
    layer0_outputs(5430) <= not(inputs(167));
    layer0_outputs(5431) <= not(inputs(143)) or (inputs(191));
    layer0_outputs(5432) <= not((inputs(36)) xor (inputs(34)));
    layer0_outputs(5433) <= (inputs(120)) xor (inputs(190));
    layer0_outputs(5434) <= (inputs(135)) or (inputs(225));
    layer0_outputs(5435) <= (inputs(202)) and not (inputs(127));
    layer0_outputs(5436) <= not(inputs(157)) or (inputs(107));
    layer0_outputs(5437) <= '0';
    layer0_outputs(5438) <= (inputs(70)) xor (inputs(123));
    layer0_outputs(5439) <= not((inputs(223)) and (inputs(159)));
    layer0_outputs(5440) <= (inputs(183)) xor (inputs(177));
    layer0_outputs(5441) <= inputs(203);
    layer0_outputs(5442) <= not(inputs(121));
    layer0_outputs(5443) <= not(inputs(122));
    layer0_outputs(5444) <= not(inputs(197));
    layer0_outputs(5445) <= (inputs(76)) and not (inputs(17));
    layer0_outputs(5446) <= not(inputs(89)) or (inputs(0));
    layer0_outputs(5447) <= not(inputs(230)) or (inputs(191));
    layer0_outputs(5448) <= not((inputs(242)) or (inputs(189)));
    layer0_outputs(5449) <= not(inputs(110));
    layer0_outputs(5450) <= not((inputs(115)) or (inputs(132)));
    layer0_outputs(5451) <= not(inputs(86));
    layer0_outputs(5452) <= '1';
    layer0_outputs(5453) <= '0';
    layer0_outputs(5454) <= '0';
    layer0_outputs(5455) <= not((inputs(65)) xor (inputs(211)));
    layer0_outputs(5456) <= '1';
    layer0_outputs(5457) <= not(inputs(82)) or (inputs(246));
    layer0_outputs(5458) <= not(inputs(141));
    layer0_outputs(5459) <= not(inputs(84)) or (inputs(158));
    layer0_outputs(5460) <= not((inputs(171)) xor (inputs(148)));
    layer0_outputs(5461) <= '0';
    layer0_outputs(5462) <= (inputs(27)) and not (inputs(97));
    layer0_outputs(5463) <= inputs(105);
    layer0_outputs(5464) <= (inputs(180)) and not (inputs(78));
    layer0_outputs(5465) <= '1';
    layer0_outputs(5466) <= (inputs(54)) or (inputs(151));
    layer0_outputs(5467) <= (inputs(221)) and not (inputs(246));
    layer0_outputs(5468) <= not(inputs(55)) or (inputs(141));
    layer0_outputs(5469) <= (inputs(37)) and not (inputs(38));
    layer0_outputs(5470) <= (inputs(242)) and not (inputs(83));
    layer0_outputs(5471) <= (inputs(82)) xor (inputs(115));
    layer0_outputs(5472) <= (inputs(49)) and (inputs(18));
    layer0_outputs(5473) <= '1';
    layer0_outputs(5474) <= (inputs(159)) xor (inputs(147));
    layer0_outputs(5475) <= not((inputs(80)) xor (inputs(134)));
    layer0_outputs(5476) <= (inputs(138)) and not (inputs(138));
    layer0_outputs(5477) <= (inputs(89)) or (inputs(168));
    layer0_outputs(5478) <= '0';
    layer0_outputs(5479) <= not(inputs(0));
    layer0_outputs(5480) <= not((inputs(172)) or (inputs(177)));
    layer0_outputs(5481) <= not(inputs(197));
    layer0_outputs(5482) <= (inputs(202)) and not (inputs(86));
    layer0_outputs(5483) <= not(inputs(232)) or (inputs(177));
    layer0_outputs(5484) <= not(inputs(132));
    layer0_outputs(5485) <= (inputs(239)) and (inputs(8));
    layer0_outputs(5486) <= not((inputs(76)) or (inputs(148)));
    layer0_outputs(5487) <= (inputs(185)) and not (inputs(51));
    layer0_outputs(5488) <= '0';
    layer0_outputs(5489) <= not((inputs(21)) xor (inputs(6)));
    layer0_outputs(5490) <= '0';
    layer0_outputs(5491) <= not(inputs(26));
    layer0_outputs(5492) <= inputs(51);
    layer0_outputs(5493) <= not((inputs(200)) xor (inputs(4)));
    layer0_outputs(5494) <= (inputs(182)) and not (inputs(55));
    layer0_outputs(5495) <= not((inputs(208)) or (inputs(65)));
    layer0_outputs(5496) <= not(inputs(62));
    layer0_outputs(5497) <= (inputs(251)) xor (inputs(149));
    layer0_outputs(5498) <= not(inputs(207)) or (inputs(80));
    layer0_outputs(5499) <= (inputs(39)) or (inputs(4));
    layer0_outputs(5500) <= not(inputs(207));
    layer0_outputs(5501) <= not((inputs(153)) or (inputs(110)));
    layer0_outputs(5502) <= '0';
    layer0_outputs(5503) <= not(inputs(148));
    layer0_outputs(5504) <= not(inputs(164)) or (inputs(212));
    layer0_outputs(5505) <= inputs(158);
    layer0_outputs(5506) <= inputs(186);
    layer0_outputs(5507) <= not((inputs(249)) or (inputs(7)));
    layer0_outputs(5508) <= (inputs(79)) or (inputs(249));
    layer0_outputs(5509) <= not(inputs(166));
    layer0_outputs(5510) <= (inputs(69)) and not (inputs(238));
    layer0_outputs(5511) <= inputs(145);
    layer0_outputs(5512) <= not(inputs(149)) or (inputs(254));
    layer0_outputs(5513) <= (inputs(188)) and (inputs(34));
    layer0_outputs(5514) <= (inputs(163)) or (inputs(222));
    layer0_outputs(5515) <= not(inputs(45));
    layer0_outputs(5516) <= not((inputs(20)) xor (inputs(97)));
    layer0_outputs(5517) <= not(inputs(16));
    layer0_outputs(5518) <= (inputs(73)) and not (inputs(78));
    layer0_outputs(5519) <= '1';
    layer0_outputs(5520) <= inputs(59);
    layer0_outputs(5521) <= not((inputs(185)) or (inputs(193)));
    layer0_outputs(5522) <= (inputs(55)) or (inputs(154));
    layer0_outputs(5523) <= (inputs(131)) or (inputs(207));
    layer0_outputs(5524) <= (inputs(91)) or (inputs(214));
    layer0_outputs(5525) <= (inputs(63)) and not (inputs(231));
    layer0_outputs(5526) <= (inputs(146)) and not (inputs(79));
    layer0_outputs(5527) <= inputs(75);
    layer0_outputs(5528) <= not((inputs(177)) or (inputs(214)));
    layer0_outputs(5529) <= (inputs(162)) and not (inputs(158));
    layer0_outputs(5530) <= (inputs(167)) or (inputs(20));
    layer0_outputs(5531) <= inputs(245);
    layer0_outputs(5532) <= not((inputs(82)) xor (inputs(200)));
    layer0_outputs(5533) <= '1';
    layer0_outputs(5534) <= inputs(181);
    layer0_outputs(5535) <= inputs(208);
    layer0_outputs(5536) <= (inputs(176)) and (inputs(5));
    layer0_outputs(5537) <= '1';
    layer0_outputs(5538) <= not((inputs(115)) and (inputs(85)));
    layer0_outputs(5539) <= not((inputs(233)) xor (inputs(167)));
    layer0_outputs(5540) <= inputs(8);
    layer0_outputs(5541) <= not((inputs(173)) xor (inputs(159)));
    layer0_outputs(5542) <= '0';
    layer0_outputs(5543) <= not((inputs(19)) and (inputs(47)));
    layer0_outputs(5544) <= (inputs(99)) and not (inputs(193));
    layer0_outputs(5545) <= not(inputs(180));
    layer0_outputs(5546) <= '1';
    layer0_outputs(5547) <= (inputs(235)) or (inputs(210));
    layer0_outputs(5548) <= '0';
    layer0_outputs(5549) <= '0';
    layer0_outputs(5550) <= inputs(229);
    layer0_outputs(5551) <= '0';
    layer0_outputs(5552) <= not(inputs(121)) or (inputs(200));
    layer0_outputs(5553) <= inputs(217);
    layer0_outputs(5554) <= (inputs(48)) and not (inputs(134));
    layer0_outputs(5555) <= inputs(2);
    layer0_outputs(5556) <= not((inputs(218)) xor (inputs(86)));
    layer0_outputs(5557) <= inputs(232);
    layer0_outputs(5558) <= (inputs(184)) and not (inputs(197));
    layer0_outputs(5559) <= not(inputs(4)) or (inputs(139));
    layer0_outputs(5560) <= not(inputs(226));
    layer0_outputs(5561) <= inputs(232);
    layer0_outputs(5562) <= not((inputs(199)) xor (inputs(215)));
    layer0_outputs(5563) <= '0';
    layer0_outputs(5564) <= (inputs(154)) and (inputs(4));
    layer0_outputs(5565) <= (inputs(229)) xor (inputs(244));
    layer0_outputs(5566) <= (inputs(223)) and (inputs(10));
    layer0_outputs(5567) <= '1';
    layer0_outputs(5568) <= not(inputs(167));
    layer0_outputs(5569) <= '0';
    layer0_outputs(5570) <= '1';
    layer0_outputs(5571) <= not((inputs(84)) or (inputs(247)));
    layer0_outputs(5572) <= not(inputs(86));
    layer0_outputs(5573) <= not(inputs(48)) or (inputs(64));
    layer0_outputs(5574) <= not(inputs(222)) or (inputs(99));
    layer0_outputs(5575) <= (inputs(54)) or (inputs(140));
    layer0_outputs(5576) <= (inputs(151)) and not (inputs(233));
    layer0_outputs(5577) <= (inputs(20)) xor (inputs(117));
    layer0_outputs(5578) <= not((inputs(88)) xor (inputs(155)));
    layer0_outputs(5579) <= (inputs(235)) and not (inputs(118));
    layer0_outputs(5580) <= '0';
    layer0_outputs(5581) <= not(inputs(126)) or (inputs(127));
    layer0_outputs(5582) <= not((inputs(123)) and (inputs(223)));
    layer0_outputs(5583) <= not((inputs(215)) or (inputs(233)));
    layer0_outputs(5584) <= not((inputs(147)) or (inputs(91)));
    layer0_outputs(5585) <= inputs(31);
    layer0_outputs(5586) <= (inputs(241)) xor (inputs(152));
    layer0_outputs(5587) <= (inputs(38)) and not (inputs(158));
    layer0_outputs(5588) <= '0';
    layer0_outputs(5589) <= (inputs(74)) xor (inputs(211));
    layer0_outputs(5590) <= (inputs(192)) or (inputs(172));
    layer0_outputs(5591) <= inputs(171);
    layer0_outputs(5592) <= (inputs(242)) and not (inputs(14));
    layer0_outputs(5593) <= inputs(166);
    layer0_outputs(5594) <= not((inputs(30)) and (inputs(222)));
    layer0_outputs(5595) <= not(inputs(139));
    layer0_outputs(5596) <= (inputs(202)) xor (inputs(185));
    layer0_outputs(5597) <= not(inputs(126)) or (inputs(242));
    layer0_outputs(5598) <= (inputs(252)) or (inputs(73));
    layer0_outputs(5599) <= (inputs(17)) xor (inputs(63));
    layer0_outputs(5600) <= not(inputs(26)) or (inputs(175));
    layer0_outputs(5601) <= not(inputs(126));
    layer0_outputs(5602) <= (inputs(66)) and not (inputs(180));
    layer0_outputs(5603) <= not((inputs(26)) or (inputs(155)));
    layer0_outputs(5604) <= (inputs(9)) and not (inputs(46));
    layer0_outputs(5605) <= not(inputs(185)) or (inputs(212));
    layer0_outputs(5606) <= not(inputs(252)) or (inputs(41));
    layer0_outputs(5607) <= not(inputs(211)) or (inputs(49));
    layer0_outputs(5608) <= not(inputs(115)) or (inputs(215));
    layer0_outputs(5609) <= (inputs(209)) or (inputs(147));
    layer0_outputs(5610) <= not((inputs(103)) or (inputs(27)));
    layer0_outputs(5611) <= (inputs(24)) and not (inputs(254));
    layer0_outputs(5612) <= not(inputs(209));
    layer0_outputs(5613) <= (inputs(71)) and not (inputs(148));
    layer0_outputs(5614) <= (inputs(158)) and not (inputs(253));
    layer0_outputs(5615) <= inputs(16);
    layer0_outputs(5616) <= (inputs(167)) and not (inputs(236));
    layer0_outputs(5617) <= (inputs(252)) and (inputs(241));
    layer0_outputs(5618) <= (inputs(135)) and not (inputs(45));
    layer0_outputs(5619) <= '1';
    layer0_outputs(5620) <= not(inputs(34));
    layer0_outputs(5621) <= (inputs(214)) or (inputs(251));
    layer0_outputs(5622) <= inputs(51);
    layer0_outputs(5623) <= (inputs(148)) and not (inputs(128));
    layer0_outputs(5624) <= not((inputs(118)) or (inputs(54)));
    layer0_outputs(5625) <= (inputs(216)) and (inputs(243));
    layer0_outputs(5626) <= '1';
    layer0_outputs(5627) <= (inputs(32)) xor (inputs(119));
    layer0_outputs(5628) <= inputs(55);
    layer0_outputs(5629) <= (inputs(139)) xor (inputs(47));
    layer0_outputs(5630) <= (inputs(7)) or (inputs(107));
    layer0_outputs(5631) <= not((inputs(146)) xor (inputs(158)));
    layer0_outputs(5632) <= inputs(123);
    layer0_outputs(5633) <= not(inputs(65)) or (inputs(65));
    layer0_outputs(5634) <= inputs(204);
    layer0_outputs(5635) <= '1';
    layer0_outputs(5636) <= not(inputs(1)) or (inputs(216));
    layer0_outputs(5637) <= inputs(207);
    layer0_outputs(5638) <= (inputs(155)) and not (inputs(114));
    layer0_outputs(5639) <= not(inputs(188)) or (inputs(148));
    layer0_outputs(5640) <= inputs(77);
    layer0_outputs(5641) <= not((inputs(187)) or (inputs(44)));
    layer0_outputs(5642) <= not((inputs(204)) xor (inputs(58)));
    layer0_outputs(5643) <= not(inputs(155)) or (inputs(139));
    layer0_outputs(5644) <= not(inputs(90));
    layer0_outputs(5645) <= inputs(151);
    layer0_outputs(5646) <= not((inputs(72)) xor (inputs(252)));
    layer0_outputs(5647) <= '0';
    layer0_outputs(5648) <= (inputs(156)) and (inputs(201));
    layer0_outputs(5649) <= (inputs(202)) or (inputs(60));
    layer0_outputs(5650) <= not(inputs(213));
    layer0_outputs(5651) <= '0';
    layer0_outputs(5652) <= not((inputs(53)) xor (inputs(173)));
    layer0_outputs(5653) <= (inputs(232)) xor (inputs(27));
    layer0_outputs(5654) <= not(inputs(127));
    layer0_outputs(5655) <= not(inputs(182)) or (inputs(75));
    layer0_outputs(5656) <= '0';
    layer0_outputs(5657) <= (inputs(168)) and not (inputs(94));
    layer0_outputs(5658) <= '1';
    layer0_outputs(5659) <= not(inputs(197));
    layer0_outputs(5660) <= not((inputs(144)) xor (inputs(114)));
    layer0_outputs(5661) <= not((inputs(210)) xor (inputs(64)));
    layer0_outputs(5662) <= (inputs(28)) and not (inputs(123));
    layer0_outputs(5663) <= not(inputs(116));
    layer0_outputs(5664) <= '1';
    layer0_outputs(5665) <= '1';
    layer0_outputs(5666) <= inputs(220);
    layer0_outputs(5667) <= '0';
    layer0_outputs(5668) <= not((inputs(194)) or (inputs(180)));
    layer0_outputs(5669) <= '0';
    layer0_outputs(5670) <= not((inputs(137)) xor (inputs(139)));
    layer0_outputs(5671) <= '1';
    layer0_outputs(5672) <= (inputs(55)) or (inputs(42));
    layer0_outputs(5673) <= not((inputs(20)) or (inputs(140)));
    layer0_outputs(5674) <= (inputs(75)) xor (inputs(238));
    layer0_outputs(5675) <= not(inputs(5)) or (inputs(60));
    layer0_outputs(5676) <= (inputs(40)) and not (inputs(63));
    layer0_outputs(5677) <= not((inputs(170)) or (inputs(244)));
    layer0_outputs(5678) <= (inputs(250)) and not (inputs(215));
    layer0_outputs(5679) <= '1';
    layer0_outputs(5680) <= inputs(82);
    layer0_outputs(5681) <= not((inputs(254)) xor (inputs(40)));
    layer0_outputs(5682) <= inputs(210);
    layer0_outputs(5683) <= (inputs(117)) or (inputs(55));
    layer0_outputs(5684) <= (inputs(107)) or (inputs(132));
    layer0_outputs(5685) <= (inputs(236)) and not (inputs(202));
    layer0_outputs(5686) <= not(inputs(13));
    layer0_outputs(5687) <= not(inputs(66));
    layer0_outputs(5688) <= (inputs(101)) xor (inputs(14));
    layer0_outputs(5689) <= not(inputs(124));
    layer0_outputs(5690) <= not((inputs(48)) or (inputs(7)));
    layer0_outputs(5691) <= '1';
    layer0_outputs(5692) <= (inputs(50)) xor (inputs(92));
    layer0_outputs(5693) <= not(inputs(125));
    layer0_outputs(5694) <= '1';
    layer0_outputs(5695) <= inputs(39);
    layer0_outputs(5696) <= (inputs(124)) xor (inputs(30));
    layer0_outputs(5697) <= not(inputs(103));
    layer0_outputs(5698) <= not((inputs(221)) and (inputs(29)));
    layer0_outputs(5699) <= inputs(254);
    layer0_outputs(5700) <= not(inputs(44));
    layer0_outputs(5701) <= (inputs(53)) or (inputs(67));
    layer0_outputs(5702) <= '1';
    layer0_outputs(5703) <= '1';
    layer0_outputs(5704) <= not(inputs(79)) or (inputs(88));
    layer0_outputs(5705) <= not((inputs(108)) or (inputs(20)));
    layer0_outputs(5706) <= (inputs(9)) or (inputs(243));
    layer0_outputs(5707) <= inputs(31);
    layer0_outputs(5708) <= inputs(150);
    layer0_outputs(5709) <= (inputs(201)) and (inputs(86));
    layer0_outputs(5710) <= not((inputs(125)) and (inputs(233)));
    layer0_outputs(5711) <= inputs(140);
    layer0_outputs(5712) <= (inputs(206)) and not (inputs(114));
    layer0_outputs(5713) <= '0';
    layer0_outputs(5714) <= not(inputs(24)) or (inputs(33));
    layer0_outputs(5715) <= not((inputs(0)) or (inputs(75)));
    layer0_outputs(5716) <= (inputs(23)) and not (inputs(80));
    layer0_outputs(5717) <= not(inputs(52));
    layer0_outputs(5718) <= not(inputs(21));
    layer0_outputs(5719) <= (inputs(212)) and (inputs(241));
    layer0_outputs(5720) <= not(inputs(209));
    layer0_outputs(5721) <= '0';
    layer0_outputs(5722) <= (inputs(47)) and not (inputs(213));
    layer0_outputs(5723) <= (inputs(204)) or (inputs(167));
    layer0_outputs(5724) <= '1';
    layer0_outputs(5725) <= (inputs(95)) and not (inputs(86));
    layer0_outputs(5726) <= (inputs(232)) or (inputs(17));
    layer0_outputs(5727) <= not(inputs(6));
    layer0_outputs(5728) <= inputs(79);
    layer0_outputs(5729) <= (inputs(122)) and not (inputs(97));
    layer0_outputs(5730) <= '1';
    layer0_outputs(5731) <= not((inputs(123)) or (inputs(167)));
    layer0_outputs(5732) <= not(inputs(163));
    layer0_outputs(5733) <= (inputs(42)) and not (inputs(74));
    layer0_outputs(5734) <= (inputs(235)) xor (inputs(237));
    layer0_outputs(5735) <= not(inputs(178)) or (inputs(191));
    layer0_outputs(5736) <= not((inputs(75)) and (inputs(244)));
    layer0_outputs(5737) <= inputs(28);
    layer0_outputs(5738) <= not((inputs(217)) xor (inputs(211)));
    layer0_outputs(5739) <= not((inputs(164)) or (inputs(243)));
    layer0_outputs(5740) <= not(inputs(120)) or (inputs(131));
    layer0_outputs(5741) <= inputs(97);
    layer0_outputs(5742) <= (inputs(9)) or (inputs(93));
    layer0_outputs(5743) <= (inputs(36)) and not (inputs(163));
    layer0_outputs(5744) <= not((inputs(51)) xor (inputs(23)));
    layer0_outputs(5745) <= not(inputs(70));
    layer0_outputs(5746) <= (inputs(19)) and not (inputs(92));
    layer0_outputs(5747) <= '0';
    layer0_outputs(5748) <= not(inputs(88));
    layer0_outputs(5749) <= not((inputs(165)) xor (inputs(63)));
    layer0_outputs(5750) <= not(inputs(47));
    layer0_outputs(5751) <= (inputs(169)) or (inputs(134));
    layer0_outputs(5752) <= (inputs(195)) or (inputs(68));
    layer0_outputs(5753) <= inputs(190);
    layer0_outputs(5754) <= not((inputs(228)) xor (inputs(34)));
    layer0_outputs(5755) <= not((inputs(191)) xor (inputs(252)));
    layer0_outputs(5756) <= not(inputs(207));
    layer0_outputs(5757) <= (inputs(69)) and (inputs(1));
    layer0_outputs(5758) <= not(inputs(142)) or (inputs(222));
    layer0_outputs(5759) <= not((inputs(110)) or (inputs(190)));
    layer0_outputs(5760) <= (inputs(227)) or (inputs(113));
    layer0_outputs(5761) <= not(inputs(146)) or (inputs(119));
    layer0_outputs(5762) <= (inputs(170)) and not (inputs(183));
    layer0_outputs(5763) <= not(inputs(239));
    layer0_outputs(5764) <= not(inputs(133));
    layer0_outputs(5765) <= not(inputs(97)) or (inputs(22));
    layer0_outputs(5766) <= inputs(229);
    layer0_outputs(5767) <= (inputs(70)) or (inputs(89));
    layer0_outputs(5768) <= (inputs(106)) and (inputs(191));
    layer0_outputs(5769) <= (inputs(8)) and (inputs(45));
    layer0_outputs(5770) <= not(inputs(122));
    layer0_outputs(5771) <= (inputs(104)) and not (inputs(27));
    layer0_outputs(5772) <= '1';
    layer0_outputs(5773) <= (inputs(222)) and not (inputs(206));
    layer0_outputs(5774) <= inputs(4);
    layer0_outputs(5775) <= not(inputs(143)) or (inputs(73));
    layer0_outputs(5776) <= (inputs(124)) and not (inputs(189));
    layer0_outputs(5777) <= (inputs(252)) and not (inputs(212));
    layer0_outputs(5778) <= not(inputs(85)) or (inputs(129));
    layer0_outputs(5779) <= not(inputs(60));
    layer0_outputs(5780) <= not(inputs(137)) or (inputs(157));
    layer0_outputs(5781) <= not(inputs(204)) or (inputs(232));
    layer0_outputs(5782) <= not(inputs(51)) or (inputs(84));
    layer0_outputs(5783) <= not((inputs(249)) or (inputs(168)));
    layer0_outputs(5784) <= not(inputs(104));
    layer0_outputs(5785) <= (inputs(15)) and not (inputs(127));
    layer0_outputs(5786) <= (inputs(156)) and not (inputs(61));
    layer0_outputs(5787) <= not((inputs(176)) or (inputs(198)));
    layer0_outputs(5788) <= not(inputs(127));
    layer0_outputs(5789) <= not(inputs(106));
    layer0_outputs(5790) <= inputs(200);
    layer0_outputs(5791) <= '0';
    layer0_outputs(5792) <= (inputs(210)) or (inputs(181));
    layer0_outputs(5793) <= not(inputs(81));
    layer0_outputs(5794) <= not((inputs(181)) or (inputs(35)));
    layer0_outputs(5795) <= not(inputs(97));
    layer0_outputs(5796) <= inputs(44);
    layer0_outputs(5797) <= not((inputs(67)) and (inputs(87)));
    layer0_outputs(5798) <= not(inputs(6)) or (inputs(244));
    layer0_outputs(5799) <= not((inputs(43)) xor (inputs(21)));
    layer0_outputs(5800) <= (inputs(78)) and (inputs(51));
    layer0_outputs(5801) <= not((inputs(95)) or (inputs(14)));
    layer0_outputs(5802) <= not(inputs(229)) or (inputs(81));
    layer0_outputs(5803) <= (inputs(91)) xor (inputs(105));
    layer0_outputs(5804) <= (inputs(232)) and not (inputs(101));
    layer0_outputs(5805) <= not(inputs(161)) or (inputs(34));
    layer0_outputs(5806) <= not(inputs(24)) or (inputs(212));
    layer0_outputs(5807) <= not((inputs(148)) and (inputs(67)));
    layer0_outputs(5808) <= (inputs(41)) and not (inputs(85));
    layer0_outputs(5809) <= '1';
    layer0_outputs(5810) <= not(inputs(73));
    layer0_outputs(5811) <= not((inputs(23)) or (inputs(196)));
    layer0_outputs(5812) <= (inputs(144)) xor (inputs(186));
    layer0_outputs(5813) <= not(inputs(50)) or (inputs(22));
    layer0_outputs(5814) <= (inputs(221)) and not (inputs(103));
    layer0_outputs(5815) <= not(inputs(217)) or (inputs(92));
    layer0_outputs(5816) <= not(inputs(42)) or (inputs(143));
    layer0_outputs(5817) <= not(inputs(68));
    layer0_outputs(5818) <= (inputs(224)) or (inputs(53));
    layer0_outputs(5819) <= (inputs(242)) xor (inputs(4));
    layer0_outputs(5820) <= '1';
    layer0_outputs(5821) <= not((inputs(103)) and (inputs(79)));
    layer0_outputs(5822) <= inputs(60);
    layer0_outputs(5823) <= (inputs(129)) and not (inputs(14));
    layer0_outputs(5824) <= inputs(32);
    layer0_outputs(5825) <= (inputs(58)) or (inputs(97));
    layer0_outputs(5826) <= (inputs(17)) and not (inputs(38));
    layer0_outputs(5827) <= (inputs(107)) xor (inputs(230));
    layer0_outputs(5828) <= not(inputs(34)) or (inputs(99));
    layer0_outputs(5829) <= not((inputs(57)) or (inputs(94)));
    layer0_outputs(5830) <= (inputs(124)) or (inputs(16));
    layer0_outputs(5831) <= inputs(80);
    layer0_outputs(5832) <= (inputs(228)) and not (inputs(154));
    layer0_outputs(5833) <= not(inputs(249));
    layer0_outputs(5834) <= '0';
    layer0_outputs(5835) <= (inputs(226)) xor (inputs(104));
    layer0_outputs(5836) <= inputs(136);
    layer0_outputs(5837) <= not((inputs(32)) xor (inputs(134)));
    layer0_outputs(5838) <= inputs(86);
    layer0_outputs(5839) <= (inputs(141)) and not (inputs(130));
    layer0_outputs(5840) <= not(inputs(46));
    layer0_outputs(5841) <= not((inputs(189)) or (inputs(237)));
    layer0_outputs(5842) <= (inputs(19)) xor (inputs(22));
    layer0_outputs(5843) <= not((inputs(3)) xor (inputs(44)));
    layer0_outputs(5844) <= '0';
    layer0_outputs(5845) <= not((inputs(141)) or (inputs(157)));
    layer0_outputs(5846) <= (inputs(245)) xor (inputs(43));
    layer0_outputs(5847) <= (inputs(97)) and (inputs(32));
    layer0_outputs(5848) <= (inputs(118)) xor (inputs(142));
    layer0_outputs(5849) <= not((inputs(6)) xor (inputs(248)));
    layer0_outputs(5850) <= inputs(27);
    layer0_outputs(5851) <= not((inputs(152)) xor (inputs(20)));
    layer0_outputs(5852) <= not((inputs(19)) xor (inputs(93)));
    layer0_outputs(5853) <= (inputs(233)) and (inputs(39));
    layer0_outputs(5854) <= not((inputs(28)) or (inputs(217)));
    layer0_outputs(5855) <= (inputs(210)) and (inputs(145));
    layer0_outputs(5856) <= (inputs(227)) or (inputs(147));
    layer0_outputs(5857) <= (inputs(91)) or (inputs(228));
    layer0_outputs(5858) <= not((inputs(136)) or (inputs(135)));
    layer0_outputs(5859) <= (inputs(242)) and not (inputs(95));
    layer0_outputs(5860) <= inputs(136);
    layer0_outputs(5861) <= (inputs(201)) and not (inputs(16));
    layer0_outputs(5862) <= not(inputs(117));
    layer0_outputs(5863) <= '0';
    layer0_outputs(5864) <= (inputs(71)) and not (inputs(155));
    layer0_outputs(5865) <= (inputs(124)) and not (inputs(55));
    layer0_outputs(5866) <= not(inputs(37));
    layer0_outputs(5867) <= not((inputs(204)) or (inputs(200)));
    layer0_outputs(5868) <= (inputs(191)) xor (inputs(93));
    layer0_outputs(5869) <= (inputs(48)) and not (inputs(7));
    layer0_outputs(5870) <= not(inputs(172)) or (inputs(61));
    layer0_outputs(5871) <= not((inputs(174)) and (inputs(45)));
    layer0_outputs(5872) <= inputs(17);
    layer0_outputs(5873) <= not(inputs(166));
    layer0_outputs(5874) <= not(inputs(22));
    layer0_outputs(5875) <= not(inputs(137)) or (inputs(68));
    layer0_outputs(5876) <= (inputs(163)) and not (inputs(26));
    layer0_outputs(5877) <= not(inputs(119));
    layer0_outputs(5878) <= (inputs(45)) and not (inputs(252));
    layer0_outputs(5879) <= (inputs(140)) and not (inputs(73));
    layer0_outputs(5880) <= '0';
    layer0_outputs(5881) <= (inputs(155)) and not (inputs(75));
    layer0_outputs(5882) <= not(inputs(4)) or (inputs(248));
    layer0_outputs(5883) <= inputs(184);
    layer0_outputs(5884) <= (inputs(219)) and not (inputs(240));
    layer0_outputs(5885) <= (inputs(47)) xor (inputs(155));
    layer0_outputs(5886) <= not(inputs(68));
    layer0_outputs(5887) <= '1';
    layer0_outputs(5888) <= not(inputs(254)) or (inputs(209));
    layer0_outputs(5889) <= not((inputs(254)) xor (inputs(221)));
    layer0_outputs(5890) <= inputs(16);
    layer0_outputs(5891) <= not((inputs(17)) xor (inputs(8)));
    layer0_outputs(5892) <= (inputs(139)) or (inputs(133));
    layer0_outputs(5893) <= '0';
    layer0_outputs(5894) <= not(inputs(126)) or (inputs(236));
    layer0_outputs(5895) <= (inputs(180)) xor (inputs(11));
    layer0_outputs(5896) <= '1';
    layer0_outputs(5897) <= inputs(152);
    layer0_outputs(5898) <= not((inputs(82)) and (inputs(165)));
    layer0_outputs(5899) <= inputs(115);
    layer0_outputs(5900) <= not((inputs(53)) or (inputs(128)));
    layer0_outputs(5901) <= (inputs(168)) and (inputs(46));
    layer0_outputs(5902) <= inputs(218);
    layer0_outputs(5903) <= not(inputs(39));
    layer0_outputs(5904) <= inputs(162);
    layer0_outputs(5905) <= not(inputs(165));
    layer0_outputs(5906) <= inputs(155);
    layer0_outputs(5907) <= not((inputs(131)) or (inputs(153)));
    layer0_outputs(5908) <= not(inputs(58));
    layer0_outputs(5909) <= (inputs(146)) or (inputs(17));
    layer0_outputs(5910) <= not(inputs(91)) or (inputs(187));
    layer0_outputs(5911) <= not((inputs(108)) and (inputs(63)));
    layer0_outputs(5912) <= inputs(231);
    layer0_outputs(5913) <= not(inputs(40)) or (inputs(250));
    layer0_outputs(5914) <= (inputs(60)) and (inputs(224));
    layer0_outputs(5915) <= (inputs(229)) and not (inputs(46));
    layer0_outputs(5916) <= not(inputs(226)) or (inputs(253));
    layer0_outputs(5917) <= inputs(98);
    layer0_outputs(5918) <= (inputs(149)) xor (inputs(144));
    layer0_outputs(5919) <= inputs(16);
    layer0_outputs(5920) <= not(inputs(54)) or (inputs(193));
    layer0_outputs(5921) <= (inputs(15)) and (inputs(62));
    layer0_outputs(5922) <= not(inputs(169));
    layer0_outputs(5923) <= (inputs(96)) or (inputs(164));
    layer0_outputs(5924) <= (inputs(252)) xor (inputs(8));
    layer0_outputs(5925) <= not(inputs(88));
    layer0_outputs(5926) <= not(inputs(65));
    layer0_outputs(5927) <= inputs(133);
    layer0_outputs(5928) <= (inputs(126)) or (inputs(70));
    layer0_outputs(5929) <= (inputs(215)) or (inputs(9));
    layer0_outputs(5930) <= (inputs(96)) and not (inputs(39));
    layer0_outputs(5931) <= '1';
    layer0_outputs(5932) <= (inputs(229)) xor (inputs(237));
    layer0_outputs(5933) <= (inputs(173)) and not (inputs(105));
    layer0_outputs(5934) <= not((inputs(161)) and (inputs(130)));
    layer0_outputs(5935) <= not(inputs(59));
    layer0_outputs(5936) <= (inputs(9)) and not (inputs(44));
    layer0_outputs(5937) <= inputs(211);
    layer0_outputs(5938) <= '0';
    layer0_outputs(5939) <= inputs(57);
    layer0_outputs(5940) <= inputs(176);
    layer0_outputs(5941) <= '1';
    layer0_outputs(5942) <= not((inputs(141)) xor (inputs(213)));
    layer0_outputs(5943) <= not(inputs(204));
    layer0_outputs(5944) <= not((inputs(156)) or (inputs(3)));
    layer0_outputs(5945) <= not(inputs(117)) or (inputs(209));
    layer0_outputs(5946) <= inputs(86);
    layer0_outputs(5947) <= (inputs(107)) xor (inputs(228));
    layer0_outputs(5948) <= not((inputs(12)) xor (inputs(174)));
    layer0_outputs(5949) <= (inputs(56)) and not (inputs(130));
    layer0_outputs(5950) <= (inputs(129)) and not (inputs(141));
    layer0_outputs(5951) <= (inputs(71)) and not (inputs(28));
    layer0_outputs(5952) <= '0';
    layer0_outputs(5953) <= (inputs(134)) and not (inputs(25));
    layer0_outputs(5954) <= (inputs(191)) and not (inputs(158));
    layer0_outputs(5955) <= '1';
    layer0_outputs(5956) <= '0';
    layer0_outputs(5957) <= (inputs(64)) or (inputs(99));
    layer0_outputs(5958) <= not(inputs(68));
    layer0_outputs(5959) <= (inputs(108)) and (inputs(36));
    layer0_outputs(5960) <= inputs(60);
    layer0_outputs(5961) <= not(inputs(17));
    layer0_outputs(5962) <= not((inputs(30)) and (inputs(228)));
    layer0_outputs(5963) <= not((inputs(134)) or (inputs(27)));
    layer0_outputs(5964) <= inputs(132);
    layer0_outputs(5965) <= inputs(167);
    layer0_outputs(5966) <= inputs(45);
    layer0_outputs(5967) <= not((inputs(8)) and (inputs(232)));
    layer0_outputs(5968) <= (inputs(159)) or (inputs(158));
    layer0_outputs(5969) <= not((inputs(165)) xor (inputs(88)));
    layer0_outputs(5970) <= not((inputs(183)) xor (inputs(193)));
    layer0_outputs(5971) <= '0';
    layer0_outputs(5972) <= not((inputs(94)) and (inputs(35)));
    layer0_outputs(5973) <= not(inputs(108)) or (inputs(24));
    layer0_outputs(5974) <= not(inputs(26));
    layer0_outputs(5975) <= (inputs(240)) and not (inputs(112));
    layer0_outputs(5976) <= '0';
    layer0_outputs(5977) <= not((inputs(120)) or (inputs(250)));
    layer0_outputs(5978) <= not((inputs(0)) or (inputs(195)));
    layer0_outputs(5979) <= inputs(128);
    layer0_outputs(5980) <= inputs(222);
    layer0_outputs(5981) <= (inputs(138)) xor (inputs(7));
    layer0_outputs(5982) <= not(inputs(59));
    layer0_outputs(5983) <= inputs(150);
    layer0_outputs(5984) <= (inputs(115)) and not (inputs(133));
    layer0_outputs(5985) <= not(inputs(191));
    layer0_outputs(5986) <= inputs(250);
    layer0_outputs(5987) <= (inputs(165)) and not (inputs(80));
    layer0_outputs(5988) <= (inputs(152)) xor (inputs(116));
    layer0_outputs(5989) <= '0';
    layer0_outputs(5990) <= not(inputs(115));
    layer0_outputs(5991) <= inputs(249);
    layer0_outputs(5992) <= not((inputs(205)) or (inputs(188)));
    layer0_outputs(5993) <= not((inputs(42)) xor (inputs(30)));
    layer0_outputs(5994) <= not(inputs(83));
    layer0_outputs(5995) <= (inputs(155)) or (inputs(62));
    layer0_outputs(5996) <= not((inputs(233)) or (inputs(134)));
    layer0_outputs(5997) <= (inputs(169)) and not (inputs(148));
    layer0_outputs(5998) <= not(inputs(128));
    layer0_outputs(5999) <= (inputs(8)) and not (inputs(126));
    layer0_outputs(6000) <= not((inputs(222)) and (inputs(17)));
    layer0_outputs(6001) <= not(inputs(204)) or (inputs(252));
    layer0_outputs(6002) <= (inputs(112)) and (inputs(101));
    layer0_outputs(6003) <= (inputs(135)) and not (inputs(51));
    layer0_outputs(6004) <= inputs(64);
    layer0_outputs(6005) <= not((inputs(111)) xor (inputs(94)));
    layer0_outputs(6006) <= (inputs(230)) and not (inputs(186));
    layer0_outputs(6007) <= not((inputs(127)) and (inputs(68)));
    layer0_outputs(6008) <= (inputs(19)) or (inputs(238));
    layer0_outputs(6009) <= inputs(172);
    layer0_outputs(6010) <= (inputs(76)) and not (inputs(49));
    layer0_outputs(6011) <= not((inputs(30)) or (inputs(114)));
    layer0_outputs(6012) <= '0';
    layer0_outputs(6013) <= not((inputs(239)) xor (inputs(162)));
    layer0_outputs(6014) <= not((inputs(27)) xor (inputs(191)));
    layer0_outputs(6015) <= inputs(176);
    layer0_outputs(6016) <= inputs(17);
    layer0_outputs(6017) <= (inputs(96)) and (inputs(217));
    layer0_outputs(6018) <= inputs(146);
    layer0_outputs(6019) <= not((inputs(215)) and (inputs(121)));
    layer0_outputs(6020) <= (inputs(100)) and not (inputs(2));
    layer0_outputs(6021) <= '1';
    layer0_outputs(6022) <= (inputs(8)) and not (inputs(46));
    layer0_outputs(6023) <= '1';
    layer0_outputs(6024) <= (inputs(54)) and not (inputs(199));
    layer0_outputs(6025) <= not(inputs(19)) or (inputs(78));
    layer0_outputs(6026) <= (inputs(233)) xor (inputs(214));
    layer0_outputs(6027) <= (inputs(180)) and not (inputs(27));
    layer0_outputs(6028) <= not(inputs(95));
    layer0_outputs(6029) <= not((inputs(51)) and (inputs(175)));
    layer0_outputs(6030) <= not((inputs(9)) or (inputs(7)));
    layer0_outputs(6031) <= (inputs(220)) and not (inputs(94));
    layer0_outputs(6032) <= not((inputs(163)) or (inputs(139)));
    layer0_outputs(6033) <= not(inputs(247)) or (inputs(103));
    layer0_outputs(6034) <= '0';
    layer0_outputs(6035) <= (inputs(192)) or (inputs(3));
    layer0_outputs(6036) <= not((inputs(98)) or (inputs(90)));
    layer0_outputs(6037) <= (inputs(174)) xor (inputs(151));
    layer0_outputs(6038) <= not(inputs(232));
    layer0_outputs(6039) <= not(inputs(68));
    layer0_outputs(6040) <= (inputs(80)) and not (inputs(111));
    layer0_outputs(6041) <= not((inputs(135)) or (inputs(93)));
    layer0_outputs(6042) <= not(inputs(150)) or (inputs(90));
    layer0_outputs(6043) <= inputs(51);
    layer0_outputs(6044) <= inputs(236);
    layer0_outputs(6045) <= not((inputs(174)) and (inputs(242)));
    layer0_outputs(6046) <= not(inputs(139)) or (inputs(89));
    layer0_outputs(6047) <= (inputs(193)) and not (inputs(72));
    layer0_outputs(6048) <= inputs(40);
    layer0_outputs(6049) <= not((inputs(63)) and (inputs(239)));
    layer0_outputs(6050) <= not(inputs(50)) or (inputs(32));
    layer0_outputs(6051) <= (inputs(158)) or (inputs(183));
    layer0_outputs(6052) <= (inputs(115)) and not (inputs(2));
    layer0_outputs(6053) <= (inputs(119)) and not (inputs(80));
    layer0_outputs(6054) <= not(inputs(89));
    layer0_outputs(6055) <= (inputs(67)) or (inputs(77));
    layer0_outputs(6056) <= (inputs(63)) xor (inputs(216));
    layer0_outputs(6057) <= not(inputs(15));
    layer0_outputs(6058) <= not((inputs(0)) xor (inputs(144)));
    layer0_outputs(6059) <= '0';
    layer0_outputs(6060) <= not((inputs(84)) xor (inputs(201)));
    layer0_outputs(6061) <= (inputs(21)) xor (inputs(170));
    layer0_outputs(6062) <= inputs(185);
    layer0_outputs(6063) <= not(inputs(85)) or (inputs(181));
    layer0_outputs(6064) <= (inputs(70)) or (inputs(76));
    layer0_outputs(6065) <= not((inputs(92)) or (inputs(57)));
    layer0_outputs(6066) <= not(inputs(214)) or (inputs(159));
    layer0_outputs(6067) <= (inputs(170)) and not (inputs(149));
    layer0_outputs(6068) <= (inputs(69)) xor (inputs(8));
    layer0_outputs(6069) <= not(inputs(133)) or (inputs(112));
    layer0_outputs(6070) <= not(inputs(250)) or (inputs(91));
    layer0_outputs(6071) <= (inputs(151)) xor (inputs(120));
    layer0_outputs(6072) <= not(inputs(166)) or (inputs(236));
    layer0_outputs(6073) <= not((inputs(26)) or (inputs(105)));
    layer0_outputs(6074) <= not(inputs(172));
    layer0_outputs(6075) <= '1';
    layer0_outputs(6076) <= not((inputs(171)) xor (inputs(51)));
    layer0_outputs(6077) <= '0';
    layer0_outputs(6078) <= (inputs(101)) or (inputs(78));
    layer0_outputs(6079) <= inputs(173);
    layer0_outputs(6080) <= not(inputs(43));
    layer0_outputs(6081) <= (inputs(172)) or (inputs(207));
    layer0_outputs(6082) <= not(inputs(102));
    layer0_outputs(6083) <= (inputs(214)) or (inputs(55));
    layer0_outputs(6084) <= (inputs(220)) or (inputs(202));
    layer0_outputs(6085) <= not((inputs(237)) or (inputs(156)));
    layer0_outputs(6086) <= inputs(70);
    layer0_outputs(6087) <= inputs(172);
    layer0_outputs(6088) <= (inputs(23)) and (inputs(43));
    layer0_outputs(6089) <= (inputs(240)) and not (inputs(29));
    layer0_outputs(6090) <= (inputs(153)) and not (inputs(199));
    layer0_outputs(6091) <= inputs(134);
    layer0_outputs(6092) <= (inputs(134)) and not (inputs(217));
    layer0_outputs(6093) <= not(inputs(30));
    layer0_outputs(6094) <= not(inputs(54));
    layer0_outputs(6095) <= inputs(122);
    layer0_outputs(6096) <= (inputs(41)) xor (inputs(28));
    layer0_outputs(6097) <= not((inputs(18)) or (inputs(179)));
    layer0_outputs(6098) <= not(inputs(125)) or (inputs(222));
    layer0_outputs(6099) <= (inputs(92)) and (inputs(194));
    layer0_outputs(6100) <= inputs(82);
    layer0_outputs(6101) <= not((inputs(238)) and (inputs(98)));
    layer0_outputs(6102) <= (inputs(52)) or (inputs(253));
    layer0_outputs(6103) <= not((inputs(78)) or (inputs(3)));
    layer0_outputs(6104) <= inputs(86);
    layer0_outputs(6105) <= not((inputs(76)) and (inputs(12)));
    layer0_outputs(6106) <= not((inputs(38)) xor (inputs(66)));
    layer0_outputs(6107) <= not(inputs(217)) or (inputs(15));
    layer0_outputs(6108) <= (inputs(254)) and (inputs(121));
    layer0_outputs(6109) <= (inputs(178)) xor (inputs(202));
    layer0_outputs(6110) <= (inputs(31)) and (inputs(222));
    layer0_outputs(6111) <= not(inputs(137)) or (inputs(23));
    layer0_outputs(6112) <= not((inputs(147)) and (inputs(131)));
    layer0_outputs(6113) <= not((inputs(151)) or (inputs(226)));
    layer0_outputs(6114) <= (inputs(105)) and (inputs(72));
    layer0_outputs(6115) <= not((inputs(197)) or (inputs(52)));
    layer0_outputs(6116) <= (inputs(112)) and not (inputs(219));
    layer0_outputs(6117) <= (inputs(165)) or (inputs(191));
    layer0_outputs(6118) <= (inputs(55)) and not (inputs(115));
    layer0_outputs(6119) <= not(inputs(223)) or (inputs(13));
    layer0_outputs(6120) <= not(inputs(242)) or (inputs(82));
    layer0_outputs(6121) <= inputs(119);
    layer0_outputs(6122) <= not((inputs(207)) xor (inputs(168)));
    layer0_outputs(6123) <= (inputs(48)) or (inputs(187));
    layer0_outputs(6124) <= inputs(85);
    layer0_outputs(6125) <= inputs(230);
    layer0_outputs(6126) <= '1';
    layer0_outputs(6127) <= not((inputs(109)) xor (inputs(240)));
    layer0_outputs(6128) <= not((inputs(182)) xor (inputs(193)));
    layer0_outputs(6129) <= '1';
    layer0_outputs(6130) <= (inputs(153)) or (inputs(194));
    layer0_outputs(6131) <= inputs(79);
    layer0_outputs(6132) <= inputs(64);
    layer0_outputs(6133) <= inputs(113);
    layer0_outputs(6134) <= not(inputs(116)) or (inputs(33));
    layer0_outputs(6135) <= not(inputs(128));
    layer0_outputs(6136) <= not(inputs(90)) or (inputs(141));
    layer0_outputs(6137) <= not(inputs(149));
    layer0_outputs(6138) <= (inputs(205)) and not (inputs(221));
    layer0_outputs(6139) <= '0';
    layer0_outputs(6140) <= (inputs(70)) or (inputs(148));
    layer0_outputs(6141) <= not(inputs(36)) or (inputs(246));
    layer0_outputs(6142) <= not((inputs(63)) xor (inputs(181)));
    layer0_outputs(6143) <= inputs(33);
    layer0_outputs(6144) <= inputs(29);
    layer0_outputs(6145) <= inputs(224);
    layer0_outputs(6146) <= inputs(206);
    layer0_outputs(6147) <= (inputs(248)) and not (inputs(155));
    layer0_outputs(6148) <= (inputs(251)) xor (inputs(25));
    layer0_outputs(6149) <= (inputs(15)) and (inputs(41));
    layer0_outputs(6150) <= not(inputs(143));
    layer0_outputs(6151) <= '1';
    layer0_outputs(6152) <= (inputs(134)) xor (inputs(254));
    layer0_outputs(6153) <= not(inputs(138));
    layer0_outputs(6154) <= not((inputs(152)) and (inputs(246)));
    layer0_outputs(6155) <= not((inputs(168)) xor (inputs(222)));
    layer0_outputs(6156) <= not((inputs(228)) xor (inputs(213)));
    layer0_outputs(6157) <= not((inputs(160)) xor (inputs(111)));
    layer0_outputs(6158) <= inputs(245);
    layer0_outputs(6159) <= not((inputs(20)) or (inputs(94)));
    layer0_outputs(6160) <= not(inputs(47)) or (inputs(193));
    layer0_outputs(6161) <= inputs(117);
    layer0_outputs(6162) <= not((inputs(18)) xor (inputs(107)));
    layer0_outputs(6163) <= not(inputs(96));
    layer0_outputs(6164) <= not(inputs(60));
    layer0_outputs(6165) <= (inputs(8)) or (inputs(41));
    layer0_outputs(6166) <= '0';
    layer0_outputs(6167) <= (inputs(195)) xor (inputs(165));
    layer0_outputs(6168) <= (inputs(155)) and not (inputs(63));
    layer0_outputs(6169) <= not((inputs(66)) xor (inputs(162)));
    layer0_outputs(6170) <= not((inputs(53)) and (inputs(129)));
    layer0_outputs(6171) <= '0';
    layer0_outputs(6172) <= (inputs(8)) and (inputs(140));
    layer0_outputs(6173) <= inputs(229);
    layer0_outputs(6174) <= inputs(60);
    layer0_outputs(6175) <= (inputs(166)) or (inputs(149));
    layer0_outputs(6176) <= not(inputs(118));
    layer0_outputs(6177) <= not((inputs(189)) or (inputs(111)));
    layer0_outputs(6178) <= '1';
    layer0_outputs(6179) <= not(inputs(77)) or (inputs(75));
    layer0_outputs(6180) <= (inputs(141)) xor (inputs(250));
    layer0_outputs(6181) <= (inputs(121)) and not (inputs(44));
    layer0_outputs(6182) <= not(inputs(220)) or (inputs(11));
    layer0_outputs(6183) <= not(inputs(55)) or (inputs(235));
    layer0_outputs(6184) <= '1';
    layer0_outputs(6185) <= '1';
    layer0_outputs(6186) <= (inputs(59)) and not (inputs(23));
    layer0_outputs(6187) <= (inputs(75)) and not (inputs(160));
    layer0_outputs(6188) <= not((inputs(90)) and (inputs(182)));
    layer0_outputs(6189) <= not(inputs(43));
    layer0_outputs(6190) <= (inputs(205)) or (inputs(136));
    layer0_outputs(6191) <= inputs(245);
    layer0_outputs(6192) <= not((inputs(28)) xor (inputs(62)));
    layer0_outputs(6193) <= not((inputs(210)) or (inputs(74)));
    layer0_outputs(6194) <= not((inputs(41)) or (inputs(207)));
    layer0_outputs(6195) <= not(inputs(149)) or (inputs(79));
    layer0_outputs(6196) <= (inputs(63)) and not (inputs(73));
    layer0_outputs(6197) <= (inputs(26)) or (inputs(234));
    layer0_outputs(6198) <= '0';
    layer0_outputs(6199) <= not(inputs(178));
    layer0_outputs(6200) <= not(inputs(50));
    layer0_outputs(6201) <= (inputs(116)) xor (inputs(225));
    layer0_outputs(6202) <= (inputs(190)) xor (inputs(53));
    layer0_outputs(6203) <= not((inputs(111)) xor (inputs(56)));
    layer0_outputs(6204) <= not((inputs(48)) and (inputs(1)));
    layer0_outputs(6205) <= (inputs(134)) xor (inputs(239));
    layer0_outputs(6206) <= (inputs(201)) and not (inputs(67));
    layer0_outputs(6207) <= not(inputs(225));
    layer0_outputs(6208) <= not(inputs(137));
    layer0_outputs(6209) <= (inputs(251)) xor (inputs(46));
    layer0_outputs(6210) <= not(inputs(90));
    layer0_outputs(6211) <= not(inputs(2));
    layer0_outputs(6212) <= not((inputs(95)) xor (inputs(25)));
    layer0_outputs(6213) <= (inputs(235)) and not (inputs(36));
    layer0_outputs(6214) <= not((inputs(15)) xor (inputs(130)));
    layer0_outputs(6215) <= '0';
    layer0_outputs(6216) <= not(inputs(4));
    layer0_outputs(6217) <= not(inputs(210));
    layer0_outputs(6218) <= '0';
    layer0_outputs(6219) <= inputs(172);
    layer0_outputs(6220) <= not(inputs(163));
    layer0_outputs(6221) <= not(inputs(82)) or (inputs(240));
    layer0_outputs(6222) <= (inputs(167)) and (inputs(83));
    layer0_outputs(6223) <= (inputs(176)) xor (inputs(19));
    layer0_outputs(6224) <= not(inputs(174));
    layer0_outputs(6225) <= (inputs(248)) and (inputs(56));
    layer0_outputs(6226) <= (inputs(215)) and not (inputs(236));
    layer0_outputs(6227) <= not((inputs(197)) or (inputs(77)));
    layer0_outputs(6228) <= (inputs(87)) and not (inputs(126));
    layer0_outputs(6229) <= not((inputs(221)) or (inputs(80)));
    layer0_outputs(6230) <= inputs(181);
    layer0_outputs(6231) <= '0';
    layer0_outputs(6232) <= (inputs(35)) or (inputs(254));
    layer0_outputs(6233) <= (inputs(246)) and (inputs(147));
    layer0_outputs(6234) <= (inputs(90)) or (inputs(66));
    layer0_outputs(6235) <= not((inputs(125)) xor (inputs(108)));
    layer0_outputs(6236) <= (inputs(200)) xor (inputs(44));
    layer0_outputs(6237) <= not(inputs(238)) or (inputs(24));
    layer0_outputs(6238) <= '1';
    layer0_outputs(6239) <= not(inputs(177)) or (inputs(147));
    layer0_outputs(6240) <= not((inputs(201)) xor (inputs(125)));
    layer0_outputs(6241) <= not((inputs(35)) xor (inputs(136)));
    layer0_outputs(6242) <= (inputs(124)) or (inputs(51));
    layer0_outputs(6243) <= '1';
    layer0_outputs(6244) <= (inputs(242)) or (inputs(97));
    layer0_outputs(6245) <= not((inputs(12)) xor (inputs(137)));
    layer0_outputs(6246) <= not((inputs(123)) and (inputs(99)));
    layer0_outputs(6247) <= not((inputs(177)) and (inputs(1)));
    layer0_outputs(6248) <= '0';
    layer0_outputs(6249) <= inputs(215);
    layer0_outputs(6250) <= inputs(172);
    layer0_outputs(6251) <= (inputs(156)) or (inputs(155));
    layer0_outputs(6252) <= '1';
    layer0_outputs(6253) <= (inputs(1)) and not (inputs(252));
    layer0_outputs(6254) <= (inputs(88)) xor (inputs(12));
    layer0_outputs(6255) <= not((inputs(145)) xor (inputs(59)));
    layer0_outputs(6256) <= (inputs(109)) and not (inputs(254));
    layer0_outputs(6257) <= (inputs(241)) and (inputs(166));
    layer0_outputs(6258) <= (inputs(119)) xor (inputs(20));
    layer0_outputs(6259) <= (inputs(47)) or (inputs(50));
    layer0_outputs(6260) <= inputs(174);
    layer0_outputs(6261) <= (inputs(90)) and (inputs(163));
    layer0_outputs(6262) <= not((inputs(160)) and (inputs(63)));
    layer0_outputs(6263) <= not(inputs(150)) or (inputs(81));
    layer0_outputs(6264) <= inputs(237);
    layer0_outputs(6265) <= not(inputs(50)) or (inputs(223));
    layer0_outputs(6266) <= not((inputs(30)) or (inputs(94)));
    layer0_outputs(6267) <= (inputs(111)) and not (inputs(15));
    layer0_outputs(6268) <= (inputs(18)) xor (inputs(122));
    layer0_outputs(6269) <= not(inputs(186));
    layer0_outputs(6270) <= not(inputs(131));
    layer0_outputs(6271) <= '0';
    layer0_outputs(6272) <= not((inputs(68)) xor (inputs(130)));
    layer0_outputs(6273) <= not(inputs(149));
    layer0_outputs(6274) <= (inputs(31)) and (inputs(214));
    layer0_outputs(6275) <= not(inputs(38)) or (inputs(50));
    layer0_outputs(6276) <= inputs(185);
    layer0_outputs(6277) <= not((inputs(127)) xor (inputs(217)));
    layer0_outputs(6278) <= not(inputs(203));
    layer0_outputs(6279) <= (inputs(138)) xor (inputs(50));
    layer0_outputs(6280) <= (inputs(236)) and (inputs(16));
    layer0_outputs(6281) <= (inputs(249)) and (inputs(157));
    layer0_outputs(6282) <= not(inputs(119)) or (inputs(232));
    layer0_outputs(6283) <= inputs(190);
    layer0_outputs(6284) <= (inputs(102)) and not (inputs(226));
    layer0_outputs(6285) <= (inputs(17)) or (inputs(220));
    layer0_outputs(6286) <= not(inputs(247)) or (inputs(78));
    layer0_outputs(6287) <= (inputs(62)) and not (inputs(4));
    layer0_outputs(6288) <= (inputs(220)) and not (inputs(129));
    layer0_outputs(6289) <= not(inputs(16)) or (inputs(8));
    layer0_outputs(6290) <= (inputs(175)) or (inputs(253));
    layer0_outputs(6291) <= not(inputs(60));
    layer0_outputs(6292) <= (inputs(253)) and (inputs(163));
    layer0_outputs(6293) <= '0';
    layer0_outputs(6294) <= (inputs(26)) and not (inputs(73));
    layer0_outputs(6295) <= (inputs(71)) and not (inputs(107));
    layer0_outputs(6296) <= not(inputs(135));
    layer0_outputs(6297) <= not(inputs(173));
    layer0_outputs(6298) <= inputs(36);
    layer0_outputs(6299) <= (inputs(224)) or (inputs(57));
    layer0_outputs(6300) <= not(inputs(50));
    layer0_outputs(6301) <= not(inputs(23));
    layer0_outputs(6302) <= (inputs(54)) and not (inputs(209));
    layer0_outputs(6303) <= (inputs(58)) or (inputs(120));
    layer0_outputs(6304) <= not((inputs(226)) or (inputs(68)));
    layer0_outputs(6305) <= (inputs(119)) and not (inputs(174));
    layer0_outputs(6306) <= '0';
    layer0_outputs(6307) <= not((inputs(107)) xor (inputs(81)));
    layer0_outputs(6308) <= not(inputs(62));
    layer0_outputs(6309) <= '0';
    layer0_outputs(6310) <= (inputs(251)) xor (inputs(248));
    layer0_outputs(6311) <= not((inputs(62)) and (inputs(91)));
    layer0_outputs(6312) <= (inputs(199)) and not (inputs(102));
    layer0_outputs(6313) <= not((inputs(89)) or (inputs(241)));
    layer0_outputs(6314) <= not((inputs(179)) xor (inputs(65)));
    layer0_outputs(6315) <= not(inputs(245));
    layer0_outputs(6316) <= not(inputs(143));
    layer0_outputs(6317) <= not((inputs(161)) or (inputs(37)));
    layer0_outputs(6318) <= (inputs(209)) and (inputs(238));
    layer0_outputs(6319) <= (inputs(182)) xor (inputs(247));
    layer0_outputs(6320) <= not((inputs(55)) or (inputs(12)));
    layer0_outputs(6321) <= not((inputs(125)) xor (inputs(193)));
    layer0_outputs(6322) <= (inputs(198)) and (inputs(131));
    layer0_outputs(6323) <= (inputs(50)) and not (inputs(237));
    layer0_outputs(6324) <= '0';
    layer0_outputs(6325) <= not(inputs(29));
    layer0_outputs(6326) <= (inputs(104)) or (inputs(166));
    layer0_outputs(6327) <= (inputs(133)) or (inputs(22));
    layer0_outputs(6328) <= (inputs(253)) xor (inputs(208));
    layer0_outputs(6329) <= (inputs(47)) and not (inputs(39));
    layer0_outputs(6330) <= '0';
    layer0_outputs(6331) <= (inputs(250)) and not (inputs(230));
    layer0_outputs(6332) <= inputs(58);
    layer0_outputs(6333) <= (inputs(71)) and not (inputs(210));
    layer0_outputs(6334) <= (inputs(56)) and not (inputs(133));
    layer0_outputs(6335) <= (inputs(93)) and not (inputs(147));
    layer0_outputs(6336) <= (inputs(215)) or (inputs(227));
    layer0_outputs(6337) <= (inputs(96)) and (inputs(100));
    layer0_outputs(6338) <= (inputs(108)) or (inputs(88));
    layer0_outputs(6339) <= not(inputs(126)) or (inputs(184));
    layer0_outputs(6340) <= (inputs(214)) xor (inputs(120));
    layer0_outputs(6341) <= not(inputs(198));
    layer0_outputs(6342) <= not(inputs(132));
    layer0_outputs(6343) <= (inputs(35)) and not (inputs(81));
    layer0_outputs(6344) <= '0';
    layer0_outputs(6345) <= '1';
    layer0_outputs(6346) <= '1';
    layer0_outputs(6347) <= not(inputs(89));
    layer0_outputs(6348) <= (inputs(11)) and (inputs(139));
    layer0_outputs(6349) <= (inputs(49)) and (inputs(132));
    layer0_outputs(6350) <= (inputs(74)) or (inputs(160));
    layer0_outputs(6351) <= not((inputs(156)) or (inputs(190)));
    layer0_outputs(6352) <= not(inputs(29));
    layer0_outputs(6353) <= (inputs(114)) and not (inputs(219));
    layer0_outputs(6354) <= '0';
    layer0_outputs(6355) <= (inputs(93)) or (inputs(77));
    layer0_outputs(6356) <= not((inputs(153)) or (inputs(131)));
    layer0_outputs(6357) <= not((inputs(163)) xor (inputs(15)));
    layer0_outputs(6358) <= not(inputs(167));
    layer0_outputs(6359) <= not(inputs(79));
    layer0_outputs(6360) <= not(inputs(153)) or (inputs(201));
    layer0_outputs(6361) <= '1';
    layer0_outputs(6362) <= (inputs(210)) and not (inputs(113));
    layer0_outputs(6363) <= (inputs(73)) and not (inputs(22));
    layer0_outputs(6364) <= inputs(237);
    layer0_outputs(6365) <= not(inputs(40));
    layer0_outputs(6366) <= (inputs(110)) and (inputs(0));
    layer0_outputs(6367) <= inputs(40);
    layer0_outputs(6368) <= (inputs(125)) or (inputs(151));
    layer0_outputs(6369) <= '0';
    layer0_outputs(6370) <= not(inputs(98));
    layer0_outputs(6371) <= not(inputs(35)) or (inputs(39));
    layer0_outputs(6372) <= not((inputs(109)) or (inputs(205)));
    layer0_outputs(6373) <= (inputs(236)) and not (inputs(108));
    layer0_outputs(6374) <= not(inputs(247)) or (inputs(21));
    layer0_outputs(6375) <= '0';
    layer0_outputs(6376) <= not(inputs(60)) or (inputs(247));
    layer0_outputs(6377) <= inputs(149);
    layer0_outputs(6378) <= (inputs(97)) or (inputs(148));
    layer0_outputs(6379) <= '1';
    layer0_outputs(6380) <= '1';
    layer0_outputs(6381) <= not((inputs(189)) and (inputs(150)));
    layer0_outputs(6382) <= (inputs(210)) or (inputs(98));
    layer0_outputs(6383) <= (inputs(212)) and not (inputs(114));
    layer0_outputs(6384) <= (inputs(248)) or (inputs(153));
    layer0_outputs(6385) <= (inputs(241)) or (inputs(137));
    layer0_outputs(6386) <= not(inputs(82)) or (inputs(35));
    layer0_outputs(6387) <= not(inputs(102)) or (inputs(253));
    layer0_outputs(6388) <= inputs(5);
    layer0_outputs(6389) <= (inputs(22)) xor (inputs(41));
    layer0_outputs(6390) <= (inputs(97)) xor (inputs(241));
    layer0_outputs(6391) <= inputs(102);
    layer0_outputs(6392) <= (inputs(83)) or (inputs(97));
    layer0_outputs(6393) <= inputs(124);
    layer0_outputs(6394) <= '0';
    layer0_outputs(6395) <= (inputs(200)) xor (inputs(33));
    layer0_outputs(6396) <= not(inputs(139));
    layer0_outputs(6397) <= not(inputs(138)) or (inputs(144));
    layer0_outputs(6398) <= not(inputs(47));
    layer0_outputs(6399) <= not((inputs(230)) xor (inputs(191)));
    layer0_outputs(6400) <= not(inputs(141));
    layer0_outputs(6401) <= inputs(210);
    layer0_outputs(6402) <= '1';
    layer0_outputs(6403) <= inputs(167);
    layer0_outputs(6404) <= (inputs(221)) and not (inputs(19));
    layer0_outputs(6405) <= not((inputs(28)) xor (inputs(11)));
    layer0_outputs(6406) <= not((inputs(22)) or (inputs(191)));
    layer0_outputs(6407) <= not((inputs(86)) or (inputs(231)));
    layer0_outputs(6408) <= (inputs(90)) or (inputs(14));
    layer0_outputs(6409) <= '0';
    layer0_outputs(6410) <= not((inputs(77)) or (inputs(15)));
    layer0_outputs(6411) <= not((inputs(52)) or (inputs(141)));
    layer0_outputs(6412) <= not((inputs(131)) or (inputs(1)));
    layer0_outputs(6413) <= (inputs(166)) and not (inputs(131));
    layer0_outputs(6414) <= (inputs(153)) and not (inputs(162));
    layer0_outputs(6415) <= not((inputs(247)) or (inputs(123)));
    layer0_outputs(6416) <= (inputs(44)) and (inputs(74));
    layer0_outputs(6417) <= (inputs(55)) and not (inputs(64));
    layer0_outputs(6418) <= '1';
    layer0_outputs(6419) <= not((inputs(130)) and (inputs(188)));
    layer0_outputs(6420) <= (inputs(246)) and not (inputs(82));
    layer0_outputs(6421) <= not(inputs(249));
    layer0_outputs(6422) <= not(inputs(22));
    layer0_outputs(6423) <= not((inputs(215)) or (inputs(115)));
    layer0_outputs(6424) <= not((inputs(141)) or (inputs(23)));
    layer0_outputs(6425) <= (inputs(111)) and not (inputs(218));
    layer0_outputs(6426) <= not(inputs(175)) or (inputs(203));
    layer0_outputs(6427) <= not(inputs(168));
    layer0_outputs(6428) <= (inputs(147)) or (inputs(201));
    layer0_outputs(6429) <= not((inputs(141)) xor (inputs(187)));
    layer0_outputs(6430) <= not((inputs(91)) and (inputs(120)));
    layer0_outputs(6431) <= not(inputs(199));
    layer0_outputs(6432) <= inputs(167);
    layer0_outputs(6433) <= '1';
    layer0_outputs(6434) <= not(inputs(173));
    layer0_outputs(6435) <= (inputs(242)) and (inputs(39));
    layer0_outputs(6436) <= (inputs(26)) and not (inputs(8));
    layer0_outputs(6437) <= (inputs(155)) and not (inputs(2));
    layer0_outputs(6438) <= not(inputs(213));
    layer0_outputs(6439) <= not(inputs(127)) or (inputs(0));
    layer0_outputs(6440) <= not(inputs(138));
    layer0_outputs(6441) <= not((inputs(5)) xor (inputs(157)));
    layer0_outputs(6442) <= inputs(87);
    layer0_outputs(6443) <= not(inputs(94));
    layer0_outputs(6444) <= (inputs(150)) or (inputs(233));
    layer0_outputs(6445) <= (inputs(18)) xor (inputs(176));
    layer0_outputs(6446) <= (inputs(182)) and not (inputs(49));
    layer0_outputs(6447) <= (inputs(231)) or (inputs(13));
    layer0_outputs(6448) <= not(inputs(7));
    layer0_outputs(6449) <= (inputs(70)) and not (inputs(87));
    layer0_outputs(6450) <= (inputs(191)) and not (inputs(34));
    layer0_outputs(6451) <= not((inputs(113)) or (inputs(244)));
    layer0_outputs(6452) <= not(inputs(225));
    layer0_outputs(6453) <= not(inputs(105));
    layer0_outputs(6454) <= (inputs(226)) and (inputs(10));
    layer0_outputs(6455) <= (inputs(80)) or (inputs(139));
    layer0_outputs(6456) <= (inputs(187)) or (inputs(171));
    layer0_outputs(6457) <= not(inputs(33));
    layer0_outputs(6458) <= (inputs(118)) and not (inputs(50));
    layer0_outputs(6459) <= not(inputs(71)) or (inputs(118));
    layer0_outputs(6460) <= '1';
    layer0_outputs(6461) <= not(inputs(100));
    layer0_outputs(6462) <= not((inputs(70)) and (inputs(97)));
    layer0_outputs(6463) <= not(inputs(75)) or (inputs(160));
    layer0_outputs(6464) <= not(inputs(136));
    layer0_outputs(6465) <= not(inputs(113)) or (inputs(42));
    layer0_outputs(6466) <= inputs(223);
    layer0_outputs(6467) <= (inputs(106)) and not (inputs(19));
    layer0_outputs(6468) <= not(inputs(154)) or (inputs(213));
    layer0_outputs(6469) <= (inputs(214)) or (inputs(50));
    layer0_outputs(6470) <= inputs(74);
    layer0_outputs(6471) <= not(inputs(147));
    layer0_outputs(6472) <= not(inputs(195)) or (inputs(0));
    layer0_outputs(6473) <= (inputs(180)) or (inputs(165));
    layer0_outputs(6474) <= not((inputs(115)) or (inputs(110)));
    layer0_outputs(6475) <= (inputs(237)) and (inputs(176));
    layer0_outputs(6476) <= (inputs(230)) and not (inputs(21));
    layer0_outputs(6477) <= (inputs(173)) and (inputs(49));
    layer0_outputs(6478) <= (inputs(202)) xor (inputs(47));
    layer0_outputs(6479) <= not((inputs(224)) xor (inputs(53)));
    layer0_outputs(6480) <= not((inputs(193)) and (inputs(30)));
    layer0_outputs(6481) <= not(inputs(149)) or (inputs(35));
    layer0_outputs(6482) <= not(inputs(106)) or (inputs(87));
    layer0_outputs(6483) <= not(inputs(218)) or (inputs(51));
    layer0_outputs(6484) <= '1';
    layer0_outputs(6485) <= (inputs(15)) or (inputs(56));
    layer0_outputs(6486) <= not((inputs(17)) or (inputs(136)));
    layer0_outputs(6487) <= not(inputs(94));
    layer0_outputs(6488) <= (inputs(106)) and not (inputs(10));
    layer0_outputs(6489) <= not(inputs(85)) or (inputs(151));
    layer0_outputs(6490) <= '0';
    layer0_outputs(6491) <= (inputs(97)) and not (inputs(108));
    layer0_outputs(6492) <= inputs(131);
    layer0_outputs(6493) <= not((inputs(53)) xor (inputs(41)));
    layer0_outputs(6494) <= (inputs(174)) and not (inputs(63));
    layer0_outputs(6495) <= not(inputs(232)) or (inputs(207));
    layer0_outputs(6496) <= not(inputs(85));
    layer0_outputs(6497) <= not((inputs(220)) xor (inputs(173)));
    layer0_outputs(6498) <= not(inputs(83)) or (inputs(14));
    layer0_outputs(6499) <= not(inputs(165));
    layer0_outputs(6500) <= (inputs(153)) and not (inputs(144));
    layer0_outputs(6501) <= not(inputs(213));
    layer0_outputs(6502) <= not((inputs(158)) xor (inputs(4)));
    layer0_outputs(6503) <= (inputs(181)) or (inputs(4));
    layer0_outputs(6504) <= not((inputs(57)) or (inputs(174)));
    layer0_outputs(6505) <= not((inputs(252)) and (inputs(227)));
    layer0_outputs(6506) <= not(inputs(235));
    layer0_outputs(6507) <= inputs(183);
    layer0_outputs(6508) <= not(inputs(83));
    layer0_outputs(6509) <= not((inputs(35)) xor (inputs(230)));
    layer0_outputs(6510) <= (inputs(77)) and not (inputs(169));
    layer0_outputs(6511) <= inputs(239);
    layer0_outputs(6512) <= (inputs(127)) and not (inputs(240));
    layer0_outputs(6513) <= not(inputs(182));
    layer0_outputs(6514) <= (inputs(181)) and not (inputs(236));
    layer0_outputs(6515) <= (inputs(129)) or (inputs(224));
    layer0_outputs(6516) <= '0';
    layer0_outputs(6517) <= not(inputs(237)) or (inputs(159));
    layer0_outputs(6518) <= '1';
    layer0_outputs(6519) <= not((inputs(78)) xor (inputs(7)));
    layer0_outputs(6520) <= not(inputs(217));
    layer0_outputs(6521) <= (inputs(155)) or (inputs(71));
    layer0_outputs(6522) <= '0';
    layer0_outputs(6523) <= not((inputs(75)) and (inputs(228)));
    layer0_outputs(6524) <= not((inputs(232)) and (inputs(200)));
    layer0_outputs(6525) <= not((inputs(210)) and (inputs(129)));
    layer0_outputs(6526) <= not((inputs(78)) xor (inputs(55)));
    layer0_outputs(6527) <= (inputs(9)) or (inputs(151));
    layer0_outputs(6528) <= inputs(75);
    layer0_outputs(6529) <= (inputs(146)) and not (inputs(125));
    layer0_outputs(6530) <= not((inputs(212)) or (inputs(53)));
    layer0_outputs(6531) <= inputs(236);
    layer0_outputs(6532) <= (inputs(183)) or (inputs(3));
    layer0_outputs(6533) <= inputs(166);
    layer0_outputs(6534) <= inputs(109);
    layer0_outputs(6535) <= not(inputs(151)) or (inputs(105));
    layer0_outputs(6536) <= not((inputs(241)) xor (inputs(204)));
    layer0_outputs(6537) <= (inputs(107)) or (inputs(214));
    layer0_outputs(6538) <= not(inputs(74)) or (inputs(208));
    layer0_outputs(6539) <= not(inputs(213)) or (inputs(241));
    layer0_outputs(6540) <= not(inputs(229)) or (inputs(113));
    layer0_outputs(6541) <= (inputs(211)) or (inputs(47));
    layer0_outputs(6542) <= not((inputs(145)) xor (inputs(249)));
    layer0_outputs(6543) <= '1';
    layer0_outputs(6544) <= not((inputs(188)) or (inputs(171)));
    layer0_outputs(6545) <= (inputs(67)) and (inputs(225));
    layer0_outputs(6546) <= not((inputs(37)) or (inputs(166)));
    layer0_outputs(6547) <= not((inputs(95)) xor (inputs(127)));
    layer0_outputs(6548) <= not(inputs(148));
    layer0_outputs(6549) <= (inputs(142)) xor (inputs(213));
    layer0_outputs(6550) <= (inputs(224)) or (inputs(92));
    layer0_outputs(6551) <= not(inputs(148)) or (inputs(205));
    layer0_outputs(6552) <= (inputs(111)) xor (inputs(33));
    layer0_outputs(6553) <= not(inputs(171)) or (inputs(198));
    layer0_outputs(6554) <= inputs(9);
    layer0_outputs(6555) <= inputs(125);
    layer0_outputs(6556) <= '0';
    layer0_outputs(6557) <= not((inputs(235)) or (inputs(82)));
    layer0_outputs(6558) <= not(inputs(176));
    layer0_outputs(6559) <= not(inputs(142)) or (inputs(252));
    layer0_outputs(6560) <= inputs(180);
    layer0_outputs(6561) <= not((inputs(141)) or (inputs(185)));
    layer0_outputs(6562) <= not(inputs(210)) or (inputs(215));
    layer0_outputs(6563) <= not(inputs(79));
    layer0_outputs(6564) <= not((inputs(106)) and (inputs(210)));
    layer0_outputs(6565) <= not(inputs(209)) or (inputs(255));
    layer0_outputs(6566) <= not((inputs(163)) or (inputs(187)));
    layer0_outputs(6567) <= not((inputs(65)) xor (inputs(227)));
    layer0_outputs(6568) <= not(inputs(168));
    layer0_outputs(6569) <= (inputs(155)) or (inputs(54));
    layer0_outputs(6570) <= (inputs(133)) and not (inputs(193));
    layer0_outputs(6571) <= (inputs(59)) or (inputs(202));
    layer0_outputs(6572) <= not(inputs(142)) or (inputs(18));
    layer0_outputs(6573) <= not((inputs(187)) or (inputs(240)));
    layer0_outputs(6574) <= (inputs(153)) and not (inputs(211));
    layer0_outputs(6575) <= not((inputs(66)) or (inputs(204)));
    layer0_outputs(6576) <= (inputs(0)) and not (inputs(145));
    layer0_outputs(6577) <= inputs(151);
    layer0_outputs(6578) <= not(inputs(193));
    layer0_outputs(6579) <= (inputs(217)) or (inputs(162));
    layer0_outputs(6580) <= (inputs(230)) and not (inputs(36));
    layer0_outputs(6581) <= (inputs(122)) and not (inputs(44));
    layer0_outputs(6582) <= (inputs(216)) or (inputs(173));
    layer0_outputs(6583) <= not((inputs(197)) and (inputs(226)));
    layer0_outputs(6584) <= (inputs(67)) xor (inputs(127));
    layer0_outputs(6585) <= inputs(96);
    layer0_outputs(6586) <= not((inputs(51)) or (inputs(53)));
    layer0_outputs(6587) <= (inputs(122)) or (inputs(202));
    layer0_outputs(6588) <= not(inputs(230));
    layer0_outputs(6589) <= (inputs(76)) and (inputs(191));
    layer0_outputs(6590) <= (inputs(39)) or (inputs(148));
    layer0_outputs(6591) <= not((inputs(82)) or (inputs(76)));
    layer0_outputs(6592) <= inputs(165);
    layer0_outputs(6593) <= not((inputs(153)) xor (inputs(64)));
    layer0_outputs(6594) <= not(inputs(235));
    layer0_outputs(6595) <= (inputs(20)) and (inputs(209));
    layer0_outputs(6596) <= not(inputs(122));
    layer0_outputs(6597) <= (inputs(50)) and (inputs(39));
    layer0_outputs(6598) <= (inputs(111)) or (inputs(107));
    layer0_outputs(6599) <= not((inputs(195)) xor (inputs(211)));
    layer0_outputs(6600) <= (inputs(20)) or (inputs(141));
    layer0_outputs(6601) <= (inputs(164)) and not (inputs(57));
    layer0_outputs(6602) <= (inputs(56)) or (inputs(124));
    layer0_outputs(6603) <= inputs(135);
    layer0_outputs(6604) <= not((inputs(30)) or (inputs(31)));
    layer0_outputs(6605) <= inputs(139);
    layer0_outputs(6606) <= (inputs(108)) and not (inputs(80));
    layer0_outputs(6607) <= '1';
    layer0_outputs(6608) <= not(inputs(170)) or (inputs(214));
    layer0_outputs(6609) <= inputs(200);
    layer0_outputs(6610) <= not((inputs(229)) xor (inputs(14)));
    layer0_outputs(6611) <= inputs(177);
    layer0_outputs(6612) <= not(inputs(238)) or (inputs(30));
    layer0_outputs(6613) <= '1';
    layer0_outputs(6614) <= '0';
    layer0_outputs(6615) <= not((inputs(223)) or (inputs(1)));
    layer0_outputs(6616) <= not((inputs(139)) or (inputs(212)));
    layer0_outputs(6617) <= inputs(155);
    layer0_outputs(6618) <= not((inputs(17)) and (inputs(232)));
    layer0_outputs(6619) <= not((inputs(170)) or (inputs(61)));
    layer0_outputs(6620) <= not((inputs(23)) and (inputs(60)));
    layer0_outputs(6621) <= inputs(145);
    layer0_outputs(6622) <= (inputs(38)) xor (inputs(205));
    layer0_outputs(6623) <= not(inputs(102)) or (inputs(120));
    layer0_outputs(6624) <= '0';
    layer0_outputs(6625) <= not(inputs(137));
    layer0_outputs(6626) <= not(inputs(183)) or (inputs(77));
    layer0_outputs(6627) <= not(inputs(13));
    layer0_outputs(6628) <= (inputs(243)) and not (inputs(240));
    layer0_outputs(6629) <= not((inputs(61)) and (inputs(158)));
    layer0_outputs(6630) <= (inputs(147)) and not (inputs(208));
    layer0_outputs(6631) <= (inputs(167)) and (inputs(67));
    layer0_outputs(6632) <= (inputs(100)) or (inputs(115));
    layer0_outputs(6633) <= not(inputs(252)) or (inputs(113));
    layer0_outputs(6634) <= not(inputs(24)) or (inputs(11));
    layer0_outputs(6635) <= (inputs(115)) xor (inputs(206));
    layer0_outputs(6636) <= (inputs(14)) xor (inputs(201));
    layer0_outputs(6637) <= not(inputs(229));
    layer0_outputs(6638) <= not(inputs(108));
    layer0_outputs(6639) <= not((inputs(37)) and (inputs(169)));
    layer0_outputs(6640) <= not(inputs(67));
    layer0_outputs(6641) <= (inputs(189)) and not (inputs(98));
    layer0_outputs(6642) <= not(inputs(247));
    layer0_outputs(6643) <= not((inputs(225)) or (inputs(174)));
    layer0_outputs(6644) <= (inputs(196)) and not (inputs(145));
    layer0_outputs(6645) <= '1';
    layer0_outputs(6646) <= not(inputs(84)) or (inputs(128));
    layer0_outputs(6647) <= inputs(168);
    layer0_outputs(6648) <= not((inputs(39)) xor (inputs(219)));
    layer0_outputs(6649) <= (inputs(110)) xor (inputs(103));
    layer0_outputs(6650) <= (inputs(141)) xor (inputs(50));
    layer0_outputs(6651) <= not((inputs(105)) or (inputs(244)));
    layer0_outputs(6652) <= '1';
    layer0_outputs(6653) <= (inputs(208)) and (inputs(187));
    layer0_outputs(6654) <= (inputs(157)) xor (inputs(117));
    layer0_outputs(6655) <= (inputs(52)) and not (inputs(63));
    layer0_outputs(6656) <= not((inputs(93)) or (inputs(216)));
    layer0_outputs(6657) <= inputs(172);
    layer0_outputs(6658) <= inputs(138);
    layer0_outputs(6659) <= '1';
    layer0_outputs(6660) <= not(inputs(5));
    layer0_outputs(6661) <= not((inputs(39)) or (inputs(27)));
    layer0_outputs(6662) <= (inputs(182)) and (inputs(144));
    layer0_outputs(6663) <= not((inputs(83)) or (inputs(153)));
    layer0_outputs(6664) <= not(inputs(123)) or (inputs(224));
    layer0_outputs(6665) <= (inputs(164)) and not (inputs(155));
    layer0_outputs(6666) <= (inputs(27)) and not (inputs(88));
    layer0_outputs(6667) <= inputs(80);
    layer0_outputs(6668) <= not(inputs(121)) or (inputs(7));
    layer0_outputs(6669) <= (inputs(225)) and not (inputs(15));
    layer0_outputs(6670) <= not((inputs(4)) xor (inputs(84)));
    layer0_outputs(6671) <= (inputs(24)) and not (inputs(81));
    layer0_outputs(6672) <= (inputs(28)) and not (inputs(119));
    layer0_outputs(6673) <= (inputs(238)) or (inputs(19));
    layer0_outputs(6674) <= (inputs(111)) or (inputs(23));
    layer0_outputs(6675) <= inputs(117);
    layer0_outputs(6676) <= inputs(250);
    layer0_outputs(6677) <= not(inputs(74)) or (inputs(217));
    layer0_outputs(6678) <= '1';
    layer0_outputs(6679) <= '0';
    layer0_outputs(6680) <= (inputs(35)) and not (inputs(101));
    layer0_outputs(6681) <= (inputs(181)) xor (inputs(237));
    layer0_outputs(6682) <= (inputs(212)) and not (inputs(130));
    layer0_outputs(6683) <= inputs(85);
    layer0_outputs(6684) <= (inputs(5)) and not (inputs(135));
    layer0_outputs(6685) <= (inputs(208)) and not (inputs(60));
    layer0_outputs(6686) <= not((inputs(106)) or (inputs(226)));
    layer0_outputs(6687) <= not((inputs(189)) or (inputs(246)));
    layer0_outputs(6688) <= (inputs(66)) and not (inputs(43));
    layer0_outputs(6689) <= not((inputs(66)) or (inputs(204)));
    layer0_outputs(6690) <= inputs(122);
    layer0_outputs(6691) <= not(inputs(151)) or (inputs(154));
    layer0_outputs(6692) <= (inputs(56)) and not (inputs(175));
    layer0_outputs(6693) <= not(inputs(179));
    layer0_outputs(6694) <= (inputs(133)) or (inputs(71));
    layer0_outputs(6695) <= (inputs(245)) or (inputs(208));
    layer0_outputs(6696) <= inputs(217);
    layer0_outputs(6697) <= (inputs(215)) xor (inputs(28));
    layer0_outputs(6698) <= not((inputs(254)) or (inputs(137)));
    layer0_outputs(6699) <= (inputs(141)) and not (inputs(248));
    layer0_outputs(6700) <= not(inputs(143)) or (inputs(62));
    layer0_outputs(6701) <= not((inputs(242)) or (inputs(134)));
    layer0_outputs(6702) <= (inputs(126)) and (inputs(81));
    layer0_outputs(6703) <= not((inputs(21)) xor (inputs(240)));
    layer0_outputs(6704) <= not(inputs(244));
    layer0_outputs(6705) <= not(inputs(94)) or (inputs(152));
    layer0_outputs(6706) <= not(inputs(125));
    layer0_outputs(6707) <= '0';
    layer0_outputs(6708) <= (inputs(176)) or (inputs(158));
    layer0_outputs(6709) <= not(inputs(242)) or (inputs(3));
    layer0_outputs(6710) <= (inputs(189)) or (inputs(196));
    layer0_outputs(6711) <= '1';
    layer0_outputs(6712) <= '1';
    layer0_outputs(6713) <= inputs(170);
    layer0_outputs(6714) <= not(inputs(163));
    layer0_outputs(6715) <= (inputs(32)) and not (inputs(146));
    layer0_outputs(6716) <= inputs(23);
    layer0_outputs(6717) <= not((inputs(0)) xor (inputs(93)));
    layer0_outputs(6718) <= '0';
    layer0_outputs(6719) <= (inputs(191)) and not (inputs(14));
    layer0_outputs(6720) <= '0';
    layer0_outputs(6721) <= '1';
    layer0_outputs(6722) <= (inputs(38)) and not (inputs(115));
    layer0_outputs(6723) <= inputs(165);
    layer0_outputs(6724) <= '1';
    layer0_outputs(6725) <= (inputs(146)) and (inputs(216));
    layer0_outputs(6726) <= not(inputs(69)) or (inputs(94));
    layer0_outputs(6727) <= '1';
    layer0_outputs(6728) <= inputs(140);
    layer0_outputs(6729) <= (inputs(92)) and not (inputs(147));
    layer0_outputs(6730) <= not(inputs(188));
    layer0_outputs(6731) <= not(inputs(67));
    layer0_outputs(6732) <= inputs(251);
    layer0_outputs(6733) <= not(inputs(155)) or (inputs(62));
    layer0_outputs(6734) <= '0';
    layer0_outputs(6735) <= not(inputs(138)) or (inputs(146));
    layer0_outputs(6736) <= not(inputs(215));
    layer0_outputs(6737) <= not((inputs(235)) and (inputs(47)));
    layer0_outputs(6738) <= not(inputs(186));
    layer0_outputs(6739) <= (inputs(247)) xor (inputs(61));
    layer0_outputs(6740) <= (inputs(178)) xor (inputs(95));
    layer0_outputs(6741) <= (inputs(12)) and (inputs(30));
    layer0_outputs(6742) <= not((inputs(7)) and (inputs(143)));
    layer0_outputs(6743) <= '0';
    layer0_outputs(6744) <= not((inputs(147)) xor (inputs(62)));
    layer0_outputs(6745) <= not(inputs(221));
    layer0_outputs(6746) <= '0';
    layer0_outputs(6747) <= not((inputs(189)) or (inputs(21)));
    layer0_outputs(6748) <= inputs(102);
    layer0_outputs(6749) <= not((inputs(65)) and (inputs(61)));
    layer0_outputs(6750) <= not((inputs(213)) xor (inputs(111)));
    layer0_outputs(6751) <= not(inputs(109));
    layer0_outputs(6752) <= not(inputs(145));
    layer0_outputs(6753) <= (inputs(218)) or (inputs(29));
    layer0_outputs(6754) <= inputs(153);
    layer0_outputs(6755) <= not((inputs(250)) xor (inputs(183)));
    layer0_outputs(6756) <= inputs(89);
    layer0_outputs(6757) <= inputs(88);
    layer0_outputs(6758) <= not(inputs(114));
    layer0_outputs(6759) <= not((inputs(84)) and (inputs(253)));
    layer0_outputs(6760) <= (inputs(48)) or (inputs(36));
    layer0_outputs(6761) <= (inputs(219)) xor (inputs(39));
    layer0_outputs(6762) <= not((inputs(181)) xor (inputs(22)));
    layer0_outputs(6763) <= not((inputs(176)) xor (inputs(135)));
    layer0_outputs(6764) <= (inputs(13)) or (inputs(50));
    layer0_outputs(6765) <= (inputs(74)) or (inputs(162));
    layer0_outputs(6766) <= (inputs(33)) and not (inputs(245));
    layer0_outputs(6767) <= inputs(67);
    layer0_outputs(6768) <= '1';
    layer0_outputs(6769) <= not((inputs(183)) xor (inputs(161)));
    layer0_outputs(6770) <= not(inputs(145));
    layer0_outputs(6771) <= not((inputs(180)) or (inputs(249)));
    layer0_outputs(6772) <= not((inputs(219)) or (inputs(118)));
    layer0_outputs(6773) <= inputs(222);
    layer0_outputs(6774) <= inputs(104);
    layer0_outputs(6775) <= not((inputs(129)) and (inputs(98)));
    layer0_outputs(6776) <= inputs(204);
    layer0_outputs(6777) <= not((inputs(24)) xor (inputs(176)));
    layer0_outputs(6778) <= (inputs(25)) and (inputs(49));
    layer0_outputs(6779) <= not((inputs(250)) xor (inputs(229)));
    layer0_outputs(6780) <= not(inputs(190)) or (inputs(87));
    layer0_outputs(6781) <= (inputs(235)) or (inputs(229));
    layer0_outputs(6782) <= (inputs(164)) and not (inputs(225));
    layer0_outputs(6783) <= not(inputs(230));
    layer0_outputs(6784) <= not(inputs(252));
    layer0_outputs(6785) <= (inputs(169)) and (inputs(0));
    layer0_outputs(6786) <= not((inputs(85)) xor (inputs(238)));
    layer0_outputs(6787) <= '0';
    layer0_outputs(6788) <= (inputs(122)) xor (inputs(19));
    layer0_outputs(6789) <= not(inputs(101)) or (inputs(132));
    layer0_outputs(6790) <= (inputs(129)) or (inputs(183));
    layer0_outputs(6791) <= inputs(174);
    layer0_outputs(6792) <= not(inputs(138)) or (inputs(195));
    layer0_outputs(6793) <= (inputs(48)) and not (inputs(183));
    layer0_outputs(6794) <= not((inputs(248)) xor (inputs(74)));
    layer0_outputs(6795) <= not(inputs(103));
    layer0_outputs(6796) <= (inputs(154)) xor (inputs(3));
    layer0_outputs(6797) <= (inputs(45)) or (inputs(194));
    layer0_outputs(6798) <= '1';
    layer0_outputs(6799) <= (inputs(82)) xor (inputs(180));
    layer0_outputs(6800) <= '1';
    layer0_outputs(6801) <= (inputs(3)) and not (inputs(140));
    layer0_outputs(6802) <= not((inputs(220)) and (inputs(89)));
    layer0_outputs(6803) <= (inputs(102)) and not (inputs(174));
    layer0_outputs(6804) <= not(inputs(127));
    layer0_outputs(6805) <= (inputs(57)) and (inputs(148));
    layer0_outputs(6806) <= '0';
    layer0_outputs(6807) <= not((inputs(218)) and (inputs(11)));
    layer0_outputs(6808) <= not(inputs(88));
    layer0_outputs(6809) <= (inputs(26)) or (inputs(148));
    layer0_outputs(6810) <= (inputs(149)) or (inputs(57));
    layer0_outputs(6811) <= (inputs(167)) xor (inputs(207));
    layer0_outputs(6812) <= not(inputs(186)) or (inputs(130));
    layer0_outputs(6813) <= (inputs(191)) or (inputs(68));
    layer0_outputs(6814) <= not((inputs(241)) or (inputs(171)));
    layer0_outputs(6815) <= inputs(44);
    layer0_outputs(6816) <= (inputs(111)) or (inputs(146));
    layer0_outputs(6817) <= (inputs(254)) or (inputs(234));
    layer0_outputs(6818) <= not((inputs(208)) and (inputs(254)));
    layer0_outputs(6819) <= not(inputs(130));
    layer0_outputs(6820) <= not((inputs(179)) and (inputs(125)));
    layer0_outputs(6821) <= not(inputs(97));
    layer0_outputs(6822) <= not((inputs(246)) and (inputs(187)));
    layer0_outputs(6823) <= (inputs(20)) and not (inputs(119));
    layer0_outputs(6824) <= (inputs(242)) and not (inputs(127));
    layer0_outputs(6825) <= (inputs(164)) and not (inputs(145));
    layer0_outputs(6826) <= (inputs(236)) xor (inputs(229));
    layer0_outputs(6827) <= not(inputs(181));
    layer0_outputs(6828) <= (inputs(111)) and (inputs(41));
    layer0_outputs(6829) <= inputs(145);
    layer0_outputs(6830) <= not(inputs(239)) or (inputs(4));
    layer0_outputs(6831) <= not((inputs(185)) or (inputs(35)));
    layer0_outputs(6832) <= not(inputs(151)) or (inputs(146));
    layer0_outputs(6833) <= inputs(118);
    layer0_outputs(6834) <= '1';
    layer0_outputs(6835) <= not((inputs(241)) or (inputs(139)));
    layer0_outputs(6836) <= not((inputs(254)) xor (inputs(137)));
    layer0_outputs(6837) <= not(inputs(7)) or (inputs(169));
    layer0_outputs(6838) <= not(inputs(150)) or (inputs(240));
    layer0_outputs(6839) <= not((inputs(39)) or (inputs(212)));
    layer0_outputs(6840) <= (inputs(11)) xor (inputs(21));
    layer0_outputs(6841) <= not(inputs(118)) or (inputs(190));
    layer0_outputs(6842) <= not((inputs(226)) and (inputs(175)));
    layer0_outputs(6843) <= not((inputs(98)) xor (inputs(167)));
    layer0_outputs(6844) <= inputs(166);
    layer0_outputs(6845) <= '0';
    layer0_outputs(6846) <= inputs(205);
    layer0_outputs(6847) <= inputs(30);
    layer0_outputs(6848) <= (inputs(187)) or (inputs(62));
    layer0_outputs(6849) <= not((inputs(155)) or (inputs(69)));
    layer0_outputs(6850) <= (inputs(0)) or (inputs(39));
    layer0_outputs(6851) <= not((inputs(170)) or (inputs(219)));
    layer0_outputs(6852) <= inputs(149);
    layer0_outputs(6853) <= inputs(90);
    layer0_outputs(6854) <= not(inputs(163));
    layer0_outputs(6855) <= not((inputs(27)) and (inputs(2)));
    layer0_outputs(6856) <= (inputs(138)) and (inputs(218));
    layer0_outputs(6857) <= not(inputs(134)) or (inputs(245));
    layer0_outputs(6858) <= not((inputs(13)) xor (inputs(76)));
    layer0_outputs(6859) <= '0';
    layer0_outputs(6860) <= not((inputs(224)) xor (inputs(52)));
    layer0_outputs(6861) <= inputs(86);
    layer0_outputs(6862) <= (inputs(26)) or (inputs(176));
    layer0_outputs(6863) <= not((inputs(253)) or (inputs(104)));
    layer0_outputs(6864) <= (inputs(246)) or (inputs(115));
    layer0_outputs(6865) <= not(inputs(192));
    layer0_outputs(6866) <= not((inputs(149)) xor (inputs(132)));
    layer0_outputs(6867) <= inputs(121);
    layer0_outputs(6868) <= not(inputs(167)) or (inputs(232));
    layer0_outputs(6869) <= inputs(29);
    layer0_outputs(6870) <= not(inputs(148)) or (inputs(69));
    layer0_outputs(6871) <= not(inputs(90)) or (inputs(87));
    layer0_outputs(6872) <= not(inputs(101));
    layer0_outputs(6873) <= inputs(250);
    layer0_outputs(6874) <= (inputs(40)) and not (inputs(104));
    layer0_outputs(6875) <= not(inputs(105));
    layer0_outputs(6876) <= not(inputs(218));
    layer0_outputs(6877) <= not(inputs(120));
    layer0_outputs(6878) <= (inputs(75)) and not (inputs(43));
    layer0_outputs(6879) <= (inputs(249)) and not (inputs(10));
    layer0_outputs(6880) <= not(inputs(87)) or (inputs(34));
    layer0_outputs(6881) <= not((inputs(187)) or (inputs(58)));
    layer0_outputs(6882) <= inputs(127);
    layer0_outputs(6883) <= '1';
    layer0_outputs(6884) <= not((inputs(222)) xor (inputs(59)));
    layer0_outputs(6885) <= '0';
    layer0_outputs(6886) <= (inputs(89)) or (inputs(157));
    layer0_outputs(6887) <= (inputs(12)) xor (inputs(138));
    layer0_outputs(6888) <= not((inputs(241)) and (inputs(168)));
    layer0_outputs(6889) <= inputs(35);
    layer0_outputs(6890) <= not(inputs(23));
    layer0_outputs(6891) <= inputs(1);
    layer0_outputs(6892) <= (inputs(252)) and not (inputs(156));
    layer0_outputs(6893) <= '1';
    layer0_outputs(6894) <= not(inputs(27));
    layer0_outputs(6895) <= inputs(14);
    layer0_outputs(6896) <= not(inputs(249)) or (inputs(129));
    layer0_outputs(6897) <= '0';
    layer0_outputs(6898) <= inputs(77);
    layer0_outputs(6899) <= not(inputs(232));
    layer0_outputs(6900) <= inputs(123);
    layer0_outputs(6901) <= (inputs(152)) and not (inputs(110));
    layer0_outputs(6902) <= not(inputs(86)) or (inputs(228));
    layer0_outputs(6903) <= not(inputs(255));
    layer0_outputs(6904) <= not((inputs(93)) and (inputs(173)));
    layer0_outputs(6905) <= not((inputs(239)) xor (inputs(108)));
    layer0_outputs(6906) <= not(inputs(110));
    layer0_outputs(6907) <= not(inputs(93)) or (inputs(71));
    layer0_outputs(6908) <= (inputs(70)) or (inputs(254));
    layer0_outputs(6909) <= (inputs(235)) xor (inputs(222));
    layer0_outputs(6910) <= not((inputs(242)) xor (inputs(42)));
    layer0_outputs(6911) <= (inputs(77)) xor (inputs(230));
    layer0_outputs(6912) <= '1';
    layer0_outputs(6913) <= inputs(207);
    layer0_outputs(6914) <= (inputs(129)) or (inputs(176));
    layer0_outputs(6915) <= (inputs(189)) or (inputs(178));
    layer0_outputs(6916) <= not(inputs(204)) or (inputs(106));
    layer0_outputs(6917) <= not(inputs(143)) or (inputs(170));
    layer0_outputs(6918) <= '0';
    layer0_outputs(6919) <= not((inputs(238)) or (inputs(166)));
    layer0_outputs(6920) <= (inputs(8)) and not (inputs(12));
    layer0_outputs(6921) <= '1';
    layer0_outputs(6922) <= not(inputs(22));
    layer0_outputs(6923) <= (inputs(181)) and not (inputs(102));
    layer0_outputs(6924) <= (inputs(162)) and not (inputs(176));
    layer0_outputs(6925) <= (inputs(112)) and not (inputs(201));
    layer0_outputs(6926) <= not((inputs(7)) or (inputs(96)));
    layer0_outputs(6927) <= not((inputs(94)) or (inputs(149)));
    layer0_outputs(6928) <= (inputs(61)) xor (inputs(80));
    layer0_outputs(6929) <= (inputs(244)) and (inputs(227));
    layer0_outputs(6930) <= (inputs(88)) and not (inputs(156));
    layer0_outputs(6931) <= not(inputs(237));
    layer0_outputs(6932) <= not((inputs(76)) or (inputs(74)));
    layer0_outputs(6933) <= (inputs(37)) or (inputs(9));
    layer0_outputs(6934) <= (inputs(237)) or (inputs(107));
    layer0_outputs(6935) <= not(inputs(163)) or (inputs(112));
    layer0_outputs(6936) <= inputs(50);
    layer0_outputs(6937) <= not(inputs(70));
    layer0_outputs(6938) <= not((inputs(251)) and (inputs(188)));
    layer0_outputs(6939) <= not((inputs(69)) or (inputs(28)));
    layer0_outputs(6940) <= not(inputs(248)) or (inputs(44));
    layer0_outputs(6941) <= not(inputs(76));
    layer0_outputs(6942) <= not(inputs(64)) or (inputs(110));
    layer0_outputs(6943) <= (inputs(202)) and not (inputs(82));
    layer0_outputs(6944) <= (inputs(50)) and (inputs(249));
    layer0_outputs(6945) <= (inputs(184)) and not (inputs(117));
    layer0_outputs(6946) <= not(inputs(87));
    layer0_outputs(6947) <= (inputs(81)) xor (inputs(124));
    layer0_outputs(6948) <= not(inputs(153));
    layer0_outputs(6949) <= inputs(158);
    layer0_outputs(6950) <= inputs(157);
    layer0_outputs(6951) <= not((inputs(12)) or (inputs(250)));
    layer0_outputs(6952) <= (inputs(179)) or (inputs(104));
    layer0_outputs(6953) <= inputs(136);
    layer0_outputs(6954) <= (inputs(87)) or (inputs(116));
    layer0_outputs(6955) <= inputs(91);
    layer0_outputs(6956) <= not(inputs(7)) or (inputs(87));
    layer0_outputs(6957) <= (inputs(246)) and (inputs(51));
    layer0_outputs(6958) <= not(inputs(194));
    layer0_outputs(6959) <= not((inputs(201)) and (inputs(167)));
    layer0_outputs(6960) <= (inputs(230)) and not (inputs(34));
    layer0_outputs(6961) <= not((inputs(103)) or (inputs(236)));
    layer0_outputs(6962) <= not(inputs(88)) or (inputs(4));
    layer0_outputs(6963) <= (inputs(56)) or (inputs(156));
    layer0_outputs(6964) <= not((inputs(246)) xor (inputs(207)));
    layer0_outputs(6965) <= (inputs(6)) and not (inputs(79));
    layer0_outputs(6966) <= '0';
    layer0_outputs(6967) <= (inputs(153)) and not (inputs(123));
    layer0_outputs(6968) <= not((inputs(133)) xor (inputs(84)));
    layer0_outputs(6969) <= (inputs(12)) and not (inputs(242));
    layer0_outputs(6970) <= '0';
    layer0_outputs(6971) <= '0';
    layer0_outputs(6972) <= not((inputs(120)) or (inputs(239)));
    layer0_outputs(6973) <= '0';
    layer0_outputs(6974) <= (inputs(216)) and not (inputs(63));
    layer0_outputs(6975) <= not((inputs(187)) or (inputs(202)));
    layer0_outputs(6976) <= not((inputs(169)) xor (inputs(161)));
    layer0_outputs(6977) <= not((inputs(127)) or (inputs(112)));
    layer0_outputs(6978) <= inputs(139);
    layer0_outputs(6979) <= (inputs(16)) and (inputs(224));
    layer0_outputs(6980) <= not((inputs(146)) or (inputs(210)));
    layer0_outputs(6981) <= not((inputs(33)) and (inputs(193)));
    layer0_outputs(6982) <= '1';
    layer0_outputs(6983) <= (inputs(96)) or (inputs(117));
    layer0_outputs(6984) <= inputs(30);
    layer0_outputs(6985) <= inputs(63);
    layer0_outputs(6986) <= (inputs(203)) xor (inputs(79));
    layer0_outputs(6987) <= not(inputs(233));
    layer0_outputs(6988) <= not(inputs(210)) or (inputs(224));
    layer0_outputs(6989) <= inputs(139);
    layer0_outputs(6990) <= not(inputs(177)) or (inputs(53));
    layer0_outputs(6991) <= (inputs(2)) xor (inputs(248));
    layer0_outputs(6992) <= not((inputs(55)) or (inputs(48)));
    layer0_outputs(6993) <= inputs(199);
    layer0_outputs(6994) <= not((inputs(53)) and (inputs(14)));
    layer0_outputs(6995) <= (inputs(135)) and not (inputs(22));
    layer0_outputs(6996) <= not((inputs(202)) or (inputs(42)));
    layer0_outputs(6997) <= '0';
    layer0_outputs(6998) <= not((inputs(96)) and (inputs(237)));
    layer0_outputs(6999) <= not(inputs(78));
    layer0_outputs(7000) <= not(inputs(119));
    layer0_outputs(7001) <= (inputs(189)) or (inputs(176));
    layer0_outputs(7002) <= not((inputs(139)) and (inputs(64)));
    layer0_outputs(7003) <= not(inputs(167)) or (inputs(214));
    layer0_outputs(7004) <= (inputs(55)) or (inputs(57));
    layer0_outputs(7005) <= (inputs(70)) and not (inputs(6));
    layer0_outputs(7006) <= not(inputs(105));
    layer0_outputs(7007) <= (inputs(60)) and not (inputs(167));
    layer0_outputs(7008) <= not(inputs(116)) or (inputs(209));
    layer0_outputs(7009) <= (inputs(30)) or (inputs(134));
    layer0_outputs(7010) <= (inputs(204)) or (inputs(72));
    layer0_outputs(7011) <= (inputs(22)) and not (inputs(106));
    layer0_outputs(7012) <= not(inputs(218)) or (inputs(45));
    layer0_outputs(7013) <= not(inputs(166));
    layer0_outputs(7014) <= (inputs(232)) or (inputs(179));
    layer0_outputs(7015) <= (inputs(108)) xor (inputs(225));
    layer0_outputs(7016) <= inputs(141);
    layer0_outputs(7017) <= not(inputs(146)) or (inputs(81));
    layer0_outputs(7018) <= not(inputs(225));
    layer0_outputs(7019) <= (inputs(53)) or (inputs(168));
    layer0_outputs(7020) <= inputs(255);
    layer0_outputs(7021) <= (inputs(211)) and not (inputs(204));
    layer0_outputs(7022) <= not(inputs(235));
    layer0_outputs(7023) <= not(inputs(61)) or (inputs(26));
    layer0_outputs(7024) <= not((inputs(192)) and (inputs(202)));
    layer0_outputs(7025) <= (inputs(174)) and not (inputs(14));
    layer0_outputs(7026) <= (inputs(45)) xor (inputs(218));
    layer0_outputs(7027) <= inputs(144);
    layer0_outputs(7028) <= (inputs(140)) and not (inputs(226));
    layer0_outputs(7029) <= (inputs(79)) xor (inputs(50));
    layer0_outputs(7030) <= not((inputs(146)) and (inputs(247)));
    layer0_outputs(7031) <= (inputs(107)) and not (inputs(185));
    layer0_outputs(7032) <= not(inputs(39)) or (inputs(139));
    layer0_outputs(7033) <= not(inputs(127));
    layer0_outputs(7034) <= not((inputs(47)) or (inputs(219)));
    layer0_outputs(7035) <= (inputs(35)) or (inputs(202));
    layer0_outputs(7036) <= inputs(154);
    layer0_outputs(7037) <= (inputs(162)) xor (inputs(111));
    layer0_outputs(7038) <= not((inputs(164)) and (inputs(136)));
    layer0_outputs(7039) <= not((inputs(26)) and (inputs(236)));
    layer0_outputs(7040) <= inputs(160);
    layer0_outputs(7041) <= '1';
    layer0_outputs(7042) <= not(inputs(243));
    layer0_outputs(7043) <= not(inputs(185));
    layer0_outputs(7044) <= inputs(216);
    layer0_outputs(7045) <= not((inputs(117)) xor (inputs(2)));
    layer0_outputs(7046) <= inputs(214);
    layer0_outputs(7047) <= not((inputs(39)) xor (inputs(19)));
    layer0_outputs(7048) <= (inputs(145)) and not (inputs(84));
    layer0_outputs(7049) <= not((inputs(1)) and (inputs(207)));
    layer0_outputs(7050) <= (inputs(74)) xor (inputs(160));
    layer0_outputs(7051) <= (inputs(93)) and not (inputs(27));
    layer0_outputs(7052) <= not(inputs(189));
    layer0_outputs(7053) <= not((inputs(119)) and (inputs(197)));
    layer0_outputs(7054) <= inputs(107);
    layer0_outputs(7055) <= not(inputs(81));
    layer0_outputs(7056) <= (inputs(93)) or (inputs(35));
    layer0_outputs(7057) <= not((inputs(53)) xor (inputs(213)));
    layer0_outputs(7058) <= inputs(185);
    layer0_outputs(7059) <= '0';
    layer0_outputs(7060) <= (inputs(209)) and not (inputs(219));
    layer0_outputs(7061) <= inputs(119);
    layer0_outputs(7062) <= not(inputs(8)) or (inputs(161));
    layer0_outputs(7063) <= (inputs(20)) and not (inputs(51));
    layer0_outputs(7064) <= inputs(181);
    layer0_outputs(7065) <= not((inputs(53)) and (inputs(87)));
    layer0_outputs(7066) <= inputs(194);
    layer0_outputs(7067) <= not((inputs(10)) or (inputs(90)));
    layer0_outputs(7068) <= not((inputs(63)) or (inputs(247)));
    layer0_outputs(7069) <= '1';
    layer0_outputs(7070) <= not(inputs(102));
    layer0_outputs(7071) <= not((inputs(160)) and (inputs(31)));
    layer0_outputs(7072) <= (inputs(35)) and not (inputs(206));
    layer0_outputs(7073) <= '0';
    layer0_outputs(7074) <= not(inputs(104)) or (inputs(45));
    layer0_outputs(7075) <= inputs(197);
    layer0_outputs(7076) <= not(inputs(22)) or (inputs(8));
    layer0_outputs(7077) <= '0';
    layer0_outputs(7078) <= (inputs(69)) xor (inputs(27));
    layer0_outputs(7079) <= inputs(180);
    layer0_outputs(7080) <= not(inputs(224)) or (inputs(178));
    layer0_outputs(7081) <= not(inputs(215));
    layer0_outputs(7082) <= (inputs(221)) and (inputs(159));
    layer0_outputs(7083) <= not(inputs(11));
    layer0_outputs(7084) <= (inputs(222)) or (inputs(98));
    layer0_outputs(7085) <= (inputs(189)) xor (inputs(11));
    layer0_outputs(7086) <= not((inputs(76)) or (inputs(179)));
    layer0_outputs(7087) <= not(inputs(70)) or (inputs(251));
    layer0_outputs(7088) <= '0';
    layer0_outputs(7089) <= not((inputs(228)) or (inputs(96)));
    layer0_outputs(7090) <= not(inputs(72)) or (inputs(52));
    layer0_outputs(7091) <= (inputs(243)) and not (inputs(183));
    layer0_outputs(7092) <= not((inputs(249)) or (inputs(97)));
    layer0_outputs(7093) <= not((inputs(157)) and (inputs(42)));
    layer0_outputs(7094) <= inputs(102);
    layer0_outputs(7095) <= not((inputs(40)) xor (inputs(101)));
    layer0_outputs(7096) <= '0';
    layer0_outputs(7097) <= (inputs(227)) and not (inputs(4));
    layer0_outputs(7098) <= (inputs(33)) and (inputs(115));
    layer0_outputs(7099) <= not((inputs(32)) or (inputs(197)));
    layer0_outputs(7100) <= not((inputs(237)) or (inputs(160)));
    layer0_outputs(7101) <= not(inputs(166)) or (inputs(234));
    layer0_outputs(7102) <= (inputs(197)) and not (inputs(67));
    layer0_outputs(7103) <= (inputs(237)) and not (inputs(232));
    layer0_outputs(7104) <= (inputs(225)) and not (inputs(56));
    layer0_outputs(7105) <= (inputs(177)) and not (inputs(199));
    layer0_outputs(7106) <= '1';
    layer0_outputs(7107) <= not((inputs(73)) and (inputs(34)));
    layer0_outputs(7108) <= not((inputs(142)) or (inputs(233)));
    layer0_outputs(7109) <= (inputs(9)) xor (inputs(55));
    layer0_outputs(7110) <= inputs(84);
    layer0_outputs(7111) <= not(inputs(57));
    layer0_outputs(7112) <= (inputs(247)) and not (inputs(191));
    layer0_outputs(7113) <= not((inputs(189)) or (inputs(31)));
    layer0_outputs(7114) <= not((inputs(208)) xor (inputs(20)));
    layer0_outputs(7115) <= not(inputs(216)) or (inputs(0));
    layer0_outputs(7116) <= '0';
    layer0_outputs(7117) <= not(inputs(106));
    layer0_outputs(7118) <= not(inputs(82)) or (inputs(243));
    layer0_outputs(7119) <= (inputs(50)) and not (inputs(218));
    layer0_outputs(7120) <= (inputs(231)) or (inputs(173));
    layer0_outputs(7121) <= not((inputs(85)) or (inputs(123)));
    layer0_outputs(7122) <= inputs(234);
    layer0_outputs(7123) <= (inputs(63)) or (inputs(168));
    layer0_outputs(7124) <= not(inputs(225)) or (inputs(151));
    layer0_outputs(7125) <= not((inputs(93)) or (inputs(157)));
    layer0_outputs(7126) <= (inputs(123)) and not (inputs(186));
    layer0_outputs(7127) <= (inputs(47)) and not (inputs(177));
    layer0_outputs(7128) <= (inputs(242)) or (inputs(207));
    layer0_outputs(7129) <= (inputs(12)) or (inputs(138));
    layer0_outputs(7130) <= (inputs(82)) and (inputs(156));
    layer0_outputs(7131) <= not(inputs(172));
    layer0_outputs(7132) <= inputs(6);
    layer0_outputs(7133) <= not((inputs(124)) and (inputs(106)));
    layer0_outputs(7134) <= not(inputs(53)) or (inputs(48));
    layer0_outputs(7135) <= (inputs(158)) xor (inputs(127));
    layer0_outputs(7136) <= not(inputs(16)) or (inputs(78));
    layer0_outputs(7137) <= (inputs(144)) or (inputs(18));
    layer0_outputs(7138) <= inputs(87);
    layer0_outputs(7139) <= (inputs(184)) and not (inputs(205));
    layer0_outputs(7140) <= (inputs(76)) or (inputs(216));
    layer0_outputs(7141) <= inputs(152);
    layer0_outputs(7142) <= (inputs(247)) or (inputs(157));
    layer0_outputs(7143) <= (inputs(129)) and not (inputs(210));
    layer0_outputs(7144) <= not(inputs(34));
    layer0_outputs(7145) <= '1';
    layer0_outputs(7146) <= not((inputs(60)) and (inputs(205)));
    layer0_outputs(7147) <= not((inputs(88)) xor (inputs(208)));
    layer0_outputs(7148) <= not(inputs(187));
    layer0_outputs(7149) <= (inputs(159)) xor (inputs(9));
    layer0_outputs(7150) <= (inputs(151)) and not (inputs(251));
    layer0_outputs(7151) <= not((inputs(210)) xor (inputs(40)));
    layer0_outputs(7152) <= not(inputs(188));
    layer0_outputs(7153) <= (inputs(86)) and not (inputs(106));
    layer0_outputs(7154) <= inputs(93);
    layer0_outputs(7155) <= inputs(73);
    layer0_outputs(7156) <= inputs(136);
    layer0_outputs(7157) <= not(inputs(200));
    layer0_outputs(7158) <= '1';
    layer0_outputs(7159) <= not((inputs(212)) xor (inputs(163)));
    layer0_outputs(7160) <= not((inputs(69)) xor (inputs(86)));
    layer0_outputs(7161) <= not(inputs(199)) or (inputs(188));
    layer0_outputs(7162) <= not(inputs(154));
    layer0_outputs(7163) <= inputs(25);
    layer0_outputs(7164) <= (inputs(185)) and not (inputs(236));
    layer0_outputs(7165) <= (inputs(126)) xor (inputs(16));
    layer0_outputs(7166) <= not(inputs(170));
    layer0_outputs(7167) <= not(inputs(104)) or (inputs(172));
    layer0_outputs(7168) <= not(inputs(204)) or (inputs(238));
    layer0_outputs(7169) <= not((inputs(54)) or (inputs(234)));
    layer0_outputs(7170) <= (inputs(234)) xor (inputs(79));
    layer0_outputs(7171) <= not(inputs(241)) or (inputs(16));
    layer0_outputs(7172) <= (inputs(115)) and (inputs(78));
    layer0_outputs(7173) <= not((inputs(32)) or (inputs(78)));
    layer0_outputs(7174) <= not(inputs(136)) or (inputs(186));
    layer0_outputs(7175) <= inputs(137);
    layer0_outputs(7176) <= '0';
    layer0_outputs(7177) <= not(inputs(5));
    layer0_outputs(7178) <= (inputs(24)) and not (inputs(140));
    layer0_outputs(7179) <= not(inputs(138)) or (inputs(25));
    layer0_outputs(7180) <= (inputs(254)) and not (inputs(250));
    layer0_outputs(7181) <= not(inputs(108)) or (inputs(72));
    layer0_outputs(7182) <= not((inputs(214)) xor (inputs(24)));
    layer0_outputs(7183) <= (inputs(168)) xor (inputs(245));
    layer0_outputs(7184) <= inputs(187);
    layer0_outputs(7185) <= (inputs(254)) xor (inputs(55));
    layer0_outputs(7186) <= '0';
    layer0_outputs(7187) <= inputs(59);
    layer0_outputs(7188) <= not(inputs(32)) or (inputs(115));
    layer0_outputs(7189) <= (inputs(161)) xor (inputs(99));
    layer0_outputs(7190) <= (inputs(199)) xor (inputs(128));
    layer0_outputs(7191) <= inputs(241);
    layer0_outputs(7192) <= not(inputs(95)) or (inputs(19));
    layer0_outputs(7193) <= (inputs(193)) xor (inputs(32));
    layer0_outputs(7194) <= (inputs(5)) and (inputs(149));
    layer0_outputs(7195) <= (inputs(215)) and not (inputs(164));
    layer0_outputs(7196) <= not((inputs(101)) and (inputs(101)));
    layer0_outputs(7197) <= inputs(6);
    layer0_outputs(7198) <= not((inputs(132)) or (inputs(109)));
    layer0_outputs(7199) <= (inputs(186)) and not (inputs(162));
    layer0_outputs(7200) <= not(inputs(154));
    layer0_outputs(7201) <= not((inputs(187)) or (inputs(216)));
    layer0_outputs(7202) <= '1';
    layer0_outputs(7203) <= inputs(63);
    layer0_outputs(7204) <= not(inputs(148)) or (inputs(241));
    layer0_outputs(7205) <= '1';
    layer0_outputs(7206) <= not(inputs(152)) or (inputs(68));
    layer0_outputs(7207) <= inputs(246);
    layer0_outputs(7208) <= (inputs(105)) or (inputs(98));
    layer0_outputs(7209) <= (inputs(153)) and not (inputs(50));
    layer0_outputs(7210) <= not(inputs(46));
    layer0_outputs(7211) <= inputs(62);
    layer0_outputs(7212) <= (inputs(4)) xor (inputs(178));
    layer0_outputs(7213) <= (inputs(136)) and not (inputs(125));
    layer0_outputs(7214) <= not(inputs(52));
    layer0_outputs(7215) <= not((inputs(251)) and (inputs(126)));
    layer0_outputs(7216) <= not((inputs(164)) or (inputs(226)));
    layer0_outputs(7217) <= (inputs(16)) or (inputs(103));
    layer0_outputs(7218) <= not(inputs(110)) or (inputs(211));
    layer0_outputs(7219) <= not(inputs(212));
    layer0_outputs(7220) <= not((inputs(9)) or (inputs(186)));
    layer0_outputs(7221) <= (inputs(104)) and (inputs(40));
    layer0_outputs(7222) <= (inputs(2)) and not (inputs(209));
    layer0_outputs(7223) <= not((inputs(125)) and (inputs(85)));
    layer0_outputs(7224) <= not((inputs(15)) and (inputs(75)));
    layer0_outputs(7225) <= '1';
    layer0_outputs(7226) <= not(inputs(176));
    layer0_outputs(7227) <= (inputs(54)) and not (inputs(100));
    layer0_outputs(7228) <= (inputs(240)) or (inputs(103));
    layer0_outputs(7229) <= not(inputs(109)) or (inputs(123));
    layer0_outputs(7230) <= (inputs(130)) and not (inputs(251));
    layer0_outputs(7231) <= (inputs(162)) and (inputs(100));
    layer0_outputs(7232) <= not(inputs(136)) or (inputs(76));
    layer0_outputs(7233) <= not((inputs(90)) and (inputs(180)));
    layer0_outputs(7234) <= inputs(217);
    layer0_outputs(7235) <= not(inputs(91)) or (inputs(27));
    layer0_outputs(7236) <= not(inputs(100)) or (inputs(131));
    layer0_outputs(7237) <= (inputs(150)) and not (inputs(219));
    layer0_outputs(7238) <= '0';
    layer0_outputs(7239) <= (inputs(42)) and (inputs(2));
    layer0_outputs(7240) <= (inputs(254)) and (inputs(8));
    layer0_outputs(7241) <= '1';
    layer0_outputs(7242) <= not(inputs(207)) or (inputs(1));
    layer0_outputs(7243) <= (inputs(73)) and not (inputs(147));
    layer0_outputs(7244) <= '1';
    layer0_outputs(7245) <= inputs(188);
    layer0_outputs(7246) <= not((inputs(134)) xor (inputs(46)));
    layer0_outputs(7247) <= not(inputs(180)) or (inputs(4));
    layer0_outputs(7248) <= (inputs(212)) or (inputs(67));
    layer0_outputs(7249) <= inputs(167);
    layer0_outputs(7250) <= (inputs(26)) and (inputs(144));
    layer0_outputs(7251) <= not(inputs(242));
    layer0_outputs(7252) <= not((inputs(168)) or (inputs(190)));
    layer0_outputs(7253) <= not((inputs(31)) and (inputs(23)));
    layer0_outputs(7254) <= not(inputs(47));
    layer0_outputs(7255) <= not((inputs(73)) or (inputs(31)));
    layer0_outputs(7256) <= '1';
    layer0_outputs(7257) <= inputs(60);
    layer0_outputs(7258) <= (inputs(3)) xor (inputs(150));
    layer0_outputs(7259) <= not((inputs(84)) and (inputs(51)));
    layer0_outputs(7260) <= (inputs(123)) xor (inputs(89));
    layer0_outputs(7261) <= not(inputs(111)) or (inputs(157));
    layer0_outputs(7262) <= inputs(163);
    layer0_outputs(7263) <= (inputs(77)) and (inputs(82));
    layer0_outputs(7264) <= not(inputs(116));
    layer0_outputs(7265) <= (inputs(182)) or (inputs(189));
    layer0_outputs(7266) <= (inputs(219)) xor (inputs(59));
    layer0_outputs(7267) <= (inputs(248)) and (inputs(64));
    layer0_outputs(7268) <= inputs(72);
    layer0_outputs(7269) <= not(inputs(56));
    layer0_outputs(7270) <= '0';
    layer0_outputs(7271) <= not(inputs(34)) or (inputs(137));
    layer0_outputs(7272) <= not(inputs(132)) or (inputs(176));
    layer0_outputs(7273) <= '0';
    layer0_outputs(7274) <= not(inputs(149));
    layer0_outputs(7275) <= inputs(149);
    layer0_outputs(7276) <= not((inputs(13)) xor (inputs(171)));
    layer0_outputs(7277) <= (inputs(11)) or (inputs(147));
    layer0_outputs(7278) <= inputs(190);
    layer0_outputs(7279) <= not(inputs(38));
    layer0_outputs(7280) <= (inputs(162)) xor (inputs(91));
    layer0_outputs(7281) <= not(inputs(10)) or (inputs(52));
    layer0_outputs(7282) <= (inputs(179)) or (inputs(137));
    layer0_outputs(7283) <= inputs(126);
    layer0_outputs(7284) <= not((inputs(71)) xor (inputs(136)));
    layer0_outputs(7285) <= (inputs(106)) and not (inputs(97));
    layer0_outputs(7286) <= inputs(129);
    layer0_outputs(7287) <= (inputs(251)) xor (inputs(24));
    layer0_outputs(7288) <= not((inputs(177)) xor (inputs(155)));
    layer0_outputs(7289) <= inputs(121);
    layer0_outputs(7290) <= not((inputs(241)) or (inputs(95)));
    layer0_outputs(7291) <= '0';
    layer0_outputs(7292) <= not(inputs(24)) or (inputs(240));
    layer0_outputs(7293) <= (inputs(122)) and not (inputs(244));
    layer0_outputs(7294) <= not(inputs(154));
    layer0_outputs(7295) <= inputs(2);
    layer0_outputs(7296) <= '1';
    layer0_outputs(7297) <= '0';
    layer0_outputs(7298) <= not(inputs(39));
    layer0_outputs(7299) <= not((inputs(33)) or (inputs(70)));
    layer0_outputs(7300) <= (inputs(172)) or (inputs(212));
    layer0_outputs(7301) <= inputs(182);
    layer0_outputs(7302) <= not(inputs(166));
    layer0_outputs(7303) <= not((inputs(67)) or (inputs(156)));
    layer0_outputs(7304) <= not(inputs(238)) or (inputs(212));
    layer0_outputs(7305) <= not((inputs(0)) xor (inputs(17)));
    layer0_outputs(7306) <= (inputs(241)) and not (inputs(211));
    layer0_outputs(7307) <= '1';
    layer0_outputs(7308) <= (inputs(205)) and (inputs(32));
    layer0_outputs(7309) <= not(inputs(137)) or (inputs(62));
    layer0_outputs(7310) <= not(inputs(56));
    layer0_outputs(7311) <= not(inputs(70));
    layer0_outputs(7312) <= (inputs(142)) and not (inputs(143));
    layer0_outputs(7313) <= '0';
    layer0_outputs(7314) <= '1';
    layer0_outputs(7315) <= (inputs(69)) or (inputs(173));
    layer0_outputs(7316) <= not(inputs(194)) or (inputs(118));
    layer0_outputs(7317) <= not((inputs(204)) xor (inputs(208)));
    layer0_outputs(7318) <= inputs(192);
    layer0_outputs(7319) <= (inputs(234)) and (inputs(252));
    layer0_outputs(7320) <= (inputs(191)) or (inputs(113));
    layer0_outputs(7321) <= not((inputs(224)) or (inputs(78)));
    layer0_outputs(7322) <= not((inputs(9)) or (inputs(200)));
    layer0_outputs(7323) <= not(inputs(49));
    layer0_outputs(7324) <= not(inputs(160)) or (inputs(47));
    layer0_outputs(7325) <= not((inputs(136)) xor (inputs(222)));
    layer0_outputs(7326) <= (inputs(214)) xor (inputs(239));
    layer0_outputs(7327) <= (inputs(12)) and not (inputs(196));
    layer0_outputs(7328) <= (inputs(104)) or (inputs(85));
    layer0_outputs(7329) <= not(inputs(184));
    layer0_outputs(7330) <= not(inputs(78));
    layer0_outputs(7331) <= (inputs(35)) xor (inputs(245));
    layer0_outputs(7332) <= not((inputs(81)) or (inputs(198)));
    layer0_outputs(7333) <= '0';
    layer0_outputs(7334) <= not(inputs(70));
    layer0_outputs(7335) <= (inputs(131)) and not (inputs(130));
    layer0_outputs(7336) <= inputs(90);
    layer0_outputs(7337) <= (inputs(138)) and not (inputs(233));
    layer0_outputs(7338) <= not((inputs(61)) xor (inputs(220)));
    layer0_outputs(7339) <= (inputs(254)) or (inputs(23));
    layer0_outputs(7340) <= (inputs(40)) and not (inputs(243));
    layer0_outputs(7341) <= not((inputs(206)) or (inputs(202)));
    layer0_outputs(7342) <= not(inputs(178));
    layer0_outputs(7343) <= not(inputs(5)) or (inputs(102));
    layer0_outputs(7344) <= (inputs(102)) or (inputs(179));
    layer0_outputs(7345) <= not(inputs(91));
    layer0_outputs(7346) <= (inputs(83)) or (inputs(68));
    layer0_outputs(7347) <= '0';
    layer0_outputs(7348) <= not((inputs(66)) xor (inputs(207)));
    layer0_outputs(7349) <= not((inputs(152)) or (inputs(59)));
    layer0_outputs(7350) <= not((inputs(59)) and (inputs(0)));
    layer0_outputs(7351) <= not(inputs(39)) or (inputs(115));
    layer0_outputs(7352) <= not((inputs(128)) xor (inputs(242)));
    layer0_outputs(7353) <= not(inputs(210)) or (inputs(248));
    layer0_outputs(7354) <= inputs(20);
    layer0_outputs(7355) <= not(inputs(175));
    layer0_outputs(7356) <= not((inputs(129)) and (inputs(24)));
    layer0_outputs(7357) <= not((inputs(18)) and (inputs(88)));
    layer0_outputs(7358) <= not(inputs(153));
    layer0_outputs(7359) <= inputs(115);
    layer0_outputs(7360) <= (inputs(214)) or (inputs(205));
    layer0_outputs(7361) <= '1';
    layer0_outputs(7362) <= '1';
    layer0_outputs(7363) <= not((inputs(204)) or (inputs(178)));
    layer0_outputs(7364) <= '1';
    layer0_outputs(7365) <= not((inputs(194)) and (inputs(97)));
    layer0_outputs(7366) <= not(inputs(173)) or (inputs(200));
    layer0_outputs(7367) <= not(inputs(57));
    layer0_outputs(7368) <= (inputs(208)) xor (inputs(233));
    layer0_outputs(7369) <= not(inputs(54));
    layer0_outputs(7370) <= '0';
    layer0_outputs(7371) <= not((inputs(241)) and (inputs(197)));
    layer0_outputs(7372) <= (inputs(187)) xor (inputs(203));
    layer0_outputs(7373) <= not((inputs(231)) or (inputs(172)));
    layer0_outputs(7374) <= not((inputs(88)) and (inputs(69)));
    layer0_outputs(7375) <= (inputs(224)) and (inputs(126));
    layer0_outputs(7376) <= not(inputs(91)) or (inputs(107));
    layer0_outputs(7377) <= '1';
    layer0_outputs(7378) <= not(inputs(139));
    layer0_outputs(7379) <= inputs(198);
    layer0_outputs(7380) <= (inputs(38)) or (inputs(10));
    layer0_outputs(7381) <= (inputs(185)) and (inputs(3));
    layer0_outputs(7382) <= inputs(211);
    layer0_outputs(7383) <= not((inputs(36)) or (inputs(222)));
    layer0_outputs(7384) <= not((inputs(0)) or (inputs(154)));
    layer0_outputs(7385) <= not((inputs(156)) and (inputs(101)));
    layer0_outputs(7386) <= '1';
    layer0_outputs(7387) <= not((inputs(180)) xor (inputs(234)));
    layer0_outputs(7388) <= (inputs(41)) or (inputs(57));
    layer0_outputs(7389) <= not(inputs(240));
    layer0_outputs(7390) <= inputs(44);
    layer0_outputs(7391) <= (inputs(230)) or (inputs(181));
    layer0_outputs(7392) <= (inputs(149)) and not (inputs(222));
    layer0_outputs(7393) <= (inputs(225)) and not (inputs(64));
    layer0_outputs(7394) <= inputs(117);
    layer0_outputs(7395) <= not((inputs(48)) and (inputs(29)));
    layer0_outputs(7396) <= not(inputs(181));
    layer0_outputs(7397) <= not((inputs(125)) and (inputs(91)));
    layer0_outputs(7398) <= (inputs(4)) xor (inputs(210));
    layer0_outputs(7399) <= (inputs(169)) and not (inputs(97));
    layer0_outputs(7400) <= inputs(167);
    layer0_outputs(7401) <= '0';
    layer0_outputs(7402) <= not((inputs(82)) xor (inputs(129)));
    layer0_outputs(7403) <= inputs(196);
    layer0_outputs(7404) <= '0';
    layer0_outputs(7405) <= not((inputs(143)) or (inputs(231)));
    layer0_outputs(7406) <= (inputs(12)) or (inputs(84));
    layer0_outputs(7407) <= not(inputs(223));
    layer0_outputs(7408) <= inputs(99);
    layer0_outputs(7409) <= '0';
    layer0_outputs(7410) <= '1';
    layer0_outputs(7411) <= not(inputs(138));
    layer0_outputs(7412) <= not((inputs(38)) xor (inputs(20)));
    layer0_outputs(7413) <= '0';
    layer0_outputs(7414) <= not((inputs(213)) and (inputs(145)));
    layer0_outputs(7415) <= (inputs(140)) and not (inputs(195));
    layer0_outputs(7416) <= (inputs(111)) xor (inputs(153));
    layer0_outputs(7417) <= inputs(67);
    layer0_outputs(7418) <= (inputs(162)) or (inputs(72));
    layer0_outputs(7419) <= inputs(237);
    layer0_outputs(7420) <= inputs(165);
    layer0_outputs(7421) <= (inputs(69)) xor (inputs(47));
    layer0_outputs(7422) <= '0';
    layer0_outputs(7423) <= (inputs(41)) and not (inputs(61));
    layer0_outputs(7424) <= '1';
    layer0_outputs(7425) <= not(inputs(218)) or (inputs(162));
    layer0_outputs(7426) <= not(inputs(128)) or (inputs(166));
    layer0_outputs(7427) <= (inputs(49)) and (inputs(211));
    layer0_outputs(7428) <= '1';
    layer0_outputs(7429) <= not(inputs(178)) or (inputs(49));
    layer0_outputs(7430) <= inputs(95);
    layer0_outputs(7431) <= not((inputs(236)) or (inputs(231)));
    layer0_outputs(7432) <= '0';
    layer0_outputs(7433) <= not(inputs(3));
    layer0_outputs(7434) <= '1';
    layer0_outputs(7435) <= not((inputs(31)) or (inputs(192)));
    layer0_outputs(7436) <= inputs(245);
    layer0_outputs(7437) <= not(inputs(250)) or (inputs(75));
    layer0_outputs(7438) <= inputs(155);
    layer0_outputs(7439) <= (inputs(95)) or (inputs(213));
    layer0_outputs(7440) <= (inputs(189)) and not (inputs(3));
    layer0_outputs(7441) <= not(inputs(94)) or (inputs(6));
    layer0_outputs(7442) <= not((inputs(188)) or (inputs(214)));
    layer0_outputs(7443) <= inputs(189);
    layer0_outputs(7444) <= (inputs(7)) or (inputs(56));
    layer0_outputs(7445) <= (inputs(204)) and not (inputs(161));
    layer0_outputs(7446) <= not((inputs(97)) and (inputs(70)));
    layer0_outputs(7447) <= not(inputs(209));
    layer0_outputs(7448) <= (inputs(253)) xor (inputs(180));
    layer0_outputs(7449) <= not(inputs(181));
    layer0_outputs(7450) <= (inputs(53)) or (inputs(184));
    layer0_outputs(7451) <= not((inputs(57)) or (inputs(171)));
    layer0_outputs(7452) <= not(inputs(48)) or (inputs(177));
    layer0_outputs(7453) <= (inputs(244)) xor (inputs(236));
    layer0_outputs(7454) <= (inputs(209)) and (inputs(173));
    layer0_outputs(7455) <= (inputs(28)) or (inputs(122));
    layer0_outputs(7456) <= not(inputs(164));
    layer0_outputs(7457) <= (inputs(120)) and not (inputs(249));
    layer0_outputs(7458) <= (inputs(117)) and not (inputs(41));
    layer0_outputs(7459) <= (inputs(32)) xor (inputs(58));
    layer0_outputs(7460) <= not((inputs(56)) or (inputs(240)));
    layer0_outputs(7461) <= not(inputs(117)) or (inputs(89));
    layer0_outputs(7462) <= not((inputs(44)) or (inputs(113)));
    layer0_outputs(7463) <= not(inputs(206)) or (inputs(206));
    layer0_outputs(7464) <= (inputs(51)) and (inputs(143));
    layer0_outputs(7465) <= (inputs(13)) and not (inputs(95));
    layer0_outputs(7466) <= not(inputs(139));
    layer0_outputs(7467) <= (inputs(235)) and (inputs(123));
    layer0_outputs(7468) <= (inputs(89)) and (inputs(215));
    layer0_outputs(7469) <= '1';
    layer0_outputs(7470) <= (inputs(192)) and not (inputs(194));
    layer0_outputs(7471) <= not((inputs(101)) or (inputs(154)));
    layer0_outputs(7472) <= '1';
    layer0_outputs(7473) <= '1';
    layer0_outputs(7474) <= not((inputs(83)) and (inputs(12)));
    layer0_outputs(7475) <= not(inputs(13)) or (inputs(60));
    layer0_outputs(7476) <= (inputs(102)) or (inputs(102));
    layer0_outputs(7477) <= not(inputs(207));
    layer0_outputs(7478) <= inputs(69);
    layer0_outputs(7479) <= (inputs(79)) and not (inputs(156));
    layer0_outputs(7480) <= (inputs(46)) or (inputs(54));
    layer0_outputs(7481) <= (inputs(116)) and not (inputs(96));
    layer0_outputs(7482) <= not(inputs(201)) or (inputs(5));
    layer0_outputs(7483) <= not(inputs(148));
    layer0_outputs(7484) <= (inputs(214)) and (inputs(97));
    layer0_outputs(7485) <= inputs(188);
    layer0_outputs(7486) <= (inputs(238)) or (inputs(20));
    layer0_outputs(7487) <= not(inputs(204));
    layer0_outputs(7488) <= not(inputs(222)) or (inputs(91));
    layer0_outputs(7489) <= not(inputs(249)) or (inputs(73));
    layer0_outputs(7490) <= (inputs(138)) and not (inputs(5));
    layer0_outputs(7491) <= not(inputs(86));
    layer0_outputs(7492) <= not(inputs(151));
    layer0_outputs(7493) <= not((inputs(140)) xor (inputs(191)));
    layer0_outputs(7494) <= not(inputs(127));
    layer0_outputs(7495) <= not(inputs(71));
    layer0_outputs(7496) <= (inputs(22)) and not (inputs(50));
    layer0_outputs(7497) <= inputs(178);
    layer0_outputs(7498) <= (inputs(99)) or (inputs(50));
    layer0_outputs(7499) <= not(inputs(21));
    layer0_outputs(7500) <= (inputs(7)) and (inputs(188));
    layer0_outputs(7501) <= (inputs(110)) xor (inputs(121));
    layer0_outputs(7502) <= not(inputs(109)) or (inputs(190));
    layer0_outputs(7503) <= not((inputs(251)) xor (inputs(247)));
    layer0_outputs(7504) <= (inputs(201)) xor (inputs(238));
    layer0_outputs(7505) <= not((inputs(247)) xor (inputs(151)));
    layer0_outputs(7506) <= (inputs(43)) or (inputs(78));
    layer0_outputs(7507) <= not(inputs(31));
    layer0_outputs(7508) <= inputs(68);
    layer0_outputs(7509) <= not((inputs(159)) xor (inputs(239)));
    layer0_outputs(7510) <= (inputs(241)) and (inputs(61));
    layer0_outputs(7511) <= not(inputs(98)) or (inputs(222));
    layer0_outputs(7512) <= (inputs(203)) or (inputs(31));
    layer0_outputs(7513) <= (inputs(81)) xor (inputs(213));
    layer0_outputs(7514) <= (inputs(155)) or (inputs(191));
    layer0_outputs(7515) <= inputs(209);
    layer0_outputs(7516) <= '1';
    layer0_outputs(7517) <= not(inputs(244)) or (inputs(125));
    layer0_outputs(7518) <= not((inputs(204)) xor (inputs(32)));
    layer0_outputs(7519) <= (inputs(140)) and (inputs(116));
    layer0_outputs(7520) <= not(inputs(67));
    layer0_outputs(7521) <= not((inputs(249)) and (inputs(38)));
    layer0_outputs(7522) <= not(inputs(167)) or (inputs(237));
    layer0_outputs(7523) <= (inputs(135)) xor (inputs(72));
    layer0_outputs(7524) <= (inputs(136)) and not (inputs(227));
    layer0_outputs(7525) <= inputs(224);
    layer0_outputs(7526) <= inputs(3);
    layer0_outputs(7527) <= not(inputs(1)) or (inputs(178));
    layer0_outputs(7528) <= (inputs(195)) and (inputs(234));
    layer0_outputs(7529) <= not((inputs(241)) or (inputs(136)));
    layer0_outputs(7530) <= '1';
    layer0_outputs(7531) <= (inputs(109)) or (inputs(165));
    layer0_outputs(7532) <= '0';
    layer0_outputs(7533) <= (inputs(77)) and not (inputs(224));
    layer0_outputs(7534) <= not(inputs(39));
    layer0_outputs(7535) <= (inputs(151)) and not (inputs(132));
    layer0_outputs(7536) <= not((inputs(28)) or (inputs(93)));
    layer0_outputs(7537) <= (inputs(226)) or (inputs(212));
    layer0_outputs(7538) <= not(inputs(110));
    layer0_outputs(7539) <= '1';
    layer0_outputs(7540) <= (inputs(173)) or (inputs(91));
    layer0_outputs(7541) <= not((inputs(103)) or (inputs(83)));
    layer0_outputs(7542) <= (inputs(118)) or (inputs(38));
    layer0_outputs(7543) <= (inputs(189)) and (inputs(19));
    layer0_outputs(7544) <= (inputs(89)) and (inputs(71));
    layer0_outputs(7545) <= (inputs(241)) and (inputs(146));
    layer0_outputs(7546) <= (inputs(149)) or (inputs(140));
    layer0_outputs(7547) <= not(inputs(156)) or (inputs(97));
    layer0_outputs(7548) <= not((inputs(215)) or (inputs(191)));
    layer0_outputs(7549) <= not(inputs(118)) or (inputs(173));
    layer0_outputs(7550) <= not((inputs(184)) or (inputs(252)));
    layer0_outputs(7551) <= inputs(231);
    layer0_outputs(7552) <= inputs(62);
    layer0_outputs(7553) <= '0';
    layer0_outputs(7554) <= inputs(111);
    layer0_outputs(7555) <= (inputs(163)) and not (inputs(21));
    layer0_outputs(7556) <= not(inputs(55)) or (inputs(46));
    layer0_outputs(7557) <= not((inputs(206)) xor (inputs(124)));
    layer0_outputs(7558) <= '0';
    layer0_outputs(7559) <= not(inputs(133)) or (inputs(159));
    layer0_outputs(7560) <= (inputs(179)) and not (inputs(219));
    layer0_outputs(7561) <= not(inputs(58));
    layer0_outputs(7562) <= (inputs(215)) and not (inputs(202));
    layer0_outputs(7563) <= '1';
    layer0_outputs(7564) <= not((inputs(25)) and (inputs(50)));
    layer0_outputs(7565) <= '1';
    layer0_outputs(7566) <= (inputs(50)) and not (inputs(113));
    layer0_outputs(7567) <= (inputs(81)) and not (inputs(46));
    layer0_outputs(7568) <= not(inputs(131));
    layer0_outputs(7569) <= (inputs(126)) xor (inputs(214));
    layer0_outputs(7570) <= (inputs(38)) and not (inputs(135));
    layer0_outputs(7571) <= not(inputs(77));
    layer0_outputs(7572) <= not((inputs(116)) or (inputs(17)));
    layer0_outputs(7573) <= inputs(20);
    layer0_outputs(7574) <= not(inputs(121)) or (inputs(200));
    layer0_outputs(7575) <= inputs(234);
    layer0_outputs(7576) <= inputs(7);
    layer0_outputs(7577) <= inputs(136);
    layer0_outputs(7578) <= (inputs(195)) or (inputs(130));
    layer0_outputs(7579) <= not(inputs(208));
    layer0_outputs(7580) <= not(inputs(89));
    layer0_outputs(7581) <= not(inputs(25)) or (inputs(84));
    layer0_outputs(7582) <= not((inputs(30)) and (inputs(249)));
    layer0_outputs(7583) <= not((inputs(62)) or (inputs(142)));
    layer0_outputs(7584) <= inputs(152);
    layer0_outputs(7585) <= (inputs(178)) or (inputs(53));
    layer0_outputs(7586) <= (inputs(166)) xor (inputs(62));
    layer0_outputs(7587) <= (inputs(136)) and not (inputs(243));
    layer0_outputs(7588) <= (inputs(216)) and not (inputs(238));
    layer0_outputs(7589) <= '0';
    layer0_outputs(7590) <= (inputs(243)) and not (inputs(49));
    layer0_outputs(7591) <= not((inputs(196)) or (inputs(124)));
    layer0_outputs(7592) <= (inputs(98)) or (inputs(1));
    layer0_outputs(7593) <= not(inputs(57));
    layer0_outputs(7594) <= (inputs(201)) and (inputs(242));
    layer0_outputs(7595) <= not((inputs(227)) and (inputs(97)));
    layer0_outputs(7596) <= inputs(207);
    layer0_outputs(7597) <= (inputs(116)) and not (inputs(112));
    layer0_outputs(7598) <= not(inputs(190));
    layer0_outputs(7599) <= inputs(98);
    layer0_outputs(7600) <= not((inputs(242)) or (inputs(245)));
    layer0_outputs(7601) <= (inputs(190)) and (inputs(235));
    layer0_outputs(7602) <= '0';
    layer0_outputs(7603) <= not((inputs(255)) xor (inputs(230)));
    layer0_outputs(7604) <= inputs(251);
    layer0_outputs(7605) <= (inputs(151)) and not (inputs(19));
    layer0_outputs(7606) <= (inputs(42)) and not (inputs(59));
    layer0_outputs(7607) <= inputs(118);
    layer0_outputs(7608) <= '1';
    layer0_outputs(7609) <= (inputs(244)) xor (inputs(158));
    layer0_outputs(7610) <= not(inputs(103)) or (inputs(69));
    layer0_outputs(7611) <= not((inputs(6)) and (inputs(64)));
    layer0_outputs(7612) <= not((inputs(75)) or (inputs(147)));
    layer0_outputs(7613) <= not(inputs(87)) or (inputs(184));
    layer0_outputs(7614) <= (inputs(151)) or (inputs(130));
    layer0_outputs(7615) <= (inputs(167)) or (inputs(46));
    layer0_outputs(7616) <= not(inputs(174));
    layer0_outputs(7617) <= not(inputs(223));
    layer0_outputs(7618) <= inputs(94);
    layer0_outputs(7619) <= inputs(10);
    layer0_outputs(7620) <= '0';
    layer0_outputs(7621) <= inputs(40);
    layer0_outputs(7622) <= inputs(35);
    layer0_outputs(7623) <= not((inputs(129)) or (inputs(124)));
    layer0_outputs(7624) <= (inputs(233)) and not (inputs(48));
    layer0_outputs(7625) <= '0';
    layer0_outputs(7626) <= (inputs(38)) and not (inputs(191));
    layer0_outputs(7627) <= (inputs(154)) xor (inputs(99));
    layer0_outputs(7628) <= not((inputs(105)) or (inputs(233)));
    layer0_outputs(7629) <= (inputs(231)) and not (inputs(243));
    layer0_outputs(7630) <= (inputs(207)) xor (inputs(18));
    layer0_outputs(7631) <= not(inputs(24)) or (inputs(156));
    layer0_outputs(7632) <= (inputs(108)) and not (inputs(150));
    layer0_outputs(7633) <= not(inputs(239));
    layer0_outputs(7634) <= inputs(58);
    layer0_outputs(7635) <= not(inputs(102)) or (inputs(14));
    layer0_outputs(7636) <= not(inputs(57)) or (inputs(33));
    layer0_outputs(7637) <= not(inputs(78));
    layer0_outputs(7638) <= not(inputs(214));
    layer0_outputs(7639) <= inputs(118);
    layer0_outputs(7640) <= not(inputs(159)) or (inputs(203));
    layer0_outputs(7641) <= '1';
    layer0_outputs(7642) <= (inputs(255)) or (inputs(140));
    layer0_outputs(7643) <= (inputs(236)) and not (inputs(249));
    layer0_outputs(7644) <= not((inputs(13)) or (inputs(150)));
    layer0_outputs(7645) <= (inputs(153)) xor (inputs(19));
    layer0_outputs(7646) <= '1';
    layer0_outputs(7647) <= not(inputs(138)) or (inputs(18));
    layer0_outputs(7648) <= not((inputs(222)) xor (inputs(91)));
    layer0_outputs(7649) <= not((inputs(193)) xor (inputs(31)));
    layer0_outputs(7650) <= not(inputs(69));
    layer0_outputs(7651) <= (inputs(40)) and not (inputs(16));
    layer0_outputs(7652) <= not((inputs(32)) and (inputs(233)));
    layer0_outputs(7653) <= not(inputs(182));
    layer0_outputs(7654) <= not(inputs(97));
    layer0_outputs(7655) <= '1';
    layer0_outputs(7656) <= (inputs(44)) xor (inputs(54));
    layer0_outputs(7657) <= '1';
    layer0_outputs(7658) <= (inputs(112)) and not (inputs(85));
    layer0_outputs(7659) <= inputs(74);
    layer0_outputs(7660) <= (inputs(201)) xor (inputs(190));
    layer0_outputs(7661) <= not((inputs(231)) and (inputs(18)));
    layer0_outputs(7662) <= not(inputs(181));
    layer0_outputs(7663) <= '0';
    layer0_outputs(7664) <= '0';
    layer0_outputs(7665) <= (inputs(179)) or (inputs(187));
    layer0_outputs(7666) <= (inputs(44)) or (inputs(77));
    layer0_outputs(7667) <= not((inputs(180)) or (inputs(20)));
    layer0_outputs(7668) <= '0';
    layer0_outputs(7669) <= not((inputs(208)) and (inputs(186)));
    layer0_outputs(7670) <= not((inputs(190)) or (inputs(215)));
    layer0_outputs(7671) <= inputs(85);
    layer0_outputs(7672) <= (inputs(171)) and (inputs(88));
    layer0_outputs(7673) <= not((inputs(107)) or (inputs(220)));
    layer0_outputs(7674) <= (inputs(103)) xor (inputs(200));
    layer0_outputs(7675) <= not((inputs(106)) or (inputs(250)));
    layer0_outputs(7676) <= inputs(0);
    layer0_outputs(7677) <= not(inputs(163));
    layer0_outputs(7678) <= (inputs(47)) and (inputs(80));
    layer0_outputs(7679) <= not(inputs(128)) or (inputs(200));
    layer0_outputs(7680) <= not(inputs(9));
    layer0_outputs(7681) <= '1';
    layer0_outputs(7682) <= not((inputs(134)) xor (inputs(204)));
    layer0_outputs(7683) <= (inputs(211)) and (inputs(205));
    layer0_outputs(7684) <= inputs(43);
    layer0_outputs(7685) <= not(inputs(54));
    layer0_outputs(7686) <= (inputs(163)) xor (inputs(95));
    layer0_outputs(7687) <= not((inputs(79)) or (inputs(139)));
    layer0_outputs(7688) <= inputs(164);
    layer0_outputs(7689) <= (inputs(252)) and not (inputs(162));
    layer0_outputs(7690) <= not((inputs(57)) xor (inputs(67)));
    layer0_outputs(7691) <= (inputs(15)) xor (inputs(8));
    layer0_outputs(7692) <= (inputs(11)) and not (inputs(182));
    layer0_outputs(7693) <= not((inputs(113)) and (inputs(52)));
    layer0_outputs(7694) <= (inputs(207)) and not (inputs(52));
    layer0_outputs(7695) <= (inputs(223)) xor (inputs(85));
    layer0_outputs(7696) <= (inputs(123)) or (inputs(42));
    layer0_outputs(7697) <= inputs(247);
    layer0_outputs(7698) <= not((inputs(15)) xor (inputs(231)));
    layer0_outputs(7699) <= not((inputs(103)) xor (inputs(115)));
    layer0_outputs(7700) <= inputs(140);
    layer0_outputs(7701) <= not(inputs(179)) or (inputs(1));
    layer0_outputs(7702) <= inputs(119);
    layer0_outputs(7703) <= not((inputs(173)) xor (inputs(88)));
    layer0_outputs(7704) <= inputs(157);
    layer0_outputs(7705) <= (inputs(208)) and not (inputs(154));
    layer0_outputs(7706) <= inputs(124);
    layer0_outputs(7707) <= not(inputs(37)) or (inputs(100));
    layer0_outputs(7708) <= not(inputs(100)) or (inputs(150));
    layer0_outputs(7709) <= not(inputs(233));
    layer0_outputs(7710) <= (inputs(225)) or (inputs(115));
    layer0_outputs(7711) <= not((inputs(226)) and (inputs(51)));
    layer0_outputs(7712) <= not(inputs(243));
    layer0_outputs(7713) <= not((inputs(11)) xor (inputs(190)));
    layer0_outputs(7714) <= (inputs(28)) xor (inputs(244));
    layer0_outputs(7715) <= (inputs(139)) or (inputs(9));
    layer0_outputs(7716) <= not((inputs(175)) and (inputs(124)));
    layer0_outputs(7717) <= '0';
    layer0_outputs(7718) <= not(inputs(192)) or (inputs(42));
    layer0_outputs(7719) <= not((inputs(16)) or (inputs(58)));
    layer0_outputs(7720) <= not((inputs(11)) or (inputs(166)));
    layer0_outputs(7721) <= not((inputs(66)) xor (inputs(158)));
    layer0_outputs(7722) <= not((inputs(36)) or (inputs(98)));
    layer0_outputs(7723) <= (inputs(101)) or (inputs(255));
    layer0_outputs(7724) <= '1';
    layer0_outputs(7725) <= inputs(198);
    layer0_outputs(7726) <= not((inputs(240)) xor (inputs(217)));
    layer0_outputs(7727) <= (inputs(173)) xor (inputs(32));
    layer0_outputs(7728) <= inputs(193);
    layer0_outputs(7729) <= not((inputs(91)) and (inputs(49)));
    layer0_outputs(7730) <= inputs(55);
    layer0_outputs(7731) <= (inputs(27)) and not (inputs(53));
    layer0_outputs(7732) <= '1';
    layer0_outputs(7733) <= not((inputs(69)) xor (inputs(31)));
    layer0_outputs(7734) <= (inputs(153)) and not (inputs(228));
    layer0_outputs(7735) <= not(inputs(170));
    layer0_outputs(7736) <= (inputs(110)) or (inputs(53));
    layer0_outputs(7737) <= inputs(43);
    layer0_outputs(7738) <= not(inputs(194));
    layer0_outputs(7739) <= not(inputs(55));
    layer0_outputs(7740) <= not((inputs(58)) and (inputs(177)));
    layer0_outputs(7741) <= inputs(145);
    layer0_outputs(7742) <= (inputs(187)) and (inputs(174));
    layer0_outputs(7743) <= (inputs(183)) or (inputs(36));
    layer0_outputs(7744) <= not((inputs(3)) and (inputs(122)));
    layer0_outputs(7745) <= not((inputs(132)) or (inputs(99)));
    layer0_outputs(7746) <= inputs(6);
    layer0_outputs(7747) <= not(inputs(109)) or (inputs(222));
    layer0_outputs(7748) <= (inputs(183)) or (inputs(22));
    layer0_outputs(7749) <= (inputs(148)) and (inputs(225));
    layer0_outputs(7750) <= (inputs(95)) and not (inputs(41));
    layer0_outputs(7751) <= not((inputs(138)) xor (inputs(190)));
    layer0_outputs(7752) <= not(inputs(233)) or (inputs(43));
    layer0_outputs(7753) <= (inputs(226)) and not (inputs(203));
    layer0_outputs(7754) <= inputs(157);
    layer0_outputs(7755) <= not((inputs(156)) xor (inputs(148)));
    layer0_outputs(7756) <= (inputs(13)) and not (inputs(143));
    layer0_outputs(7757) <= (inputs(180)) and not (inputs(15));
    layer0_outputs(7758) <= '0';
    layer0_outputs(7759) <= (inputs(87)) and not (inputs(189));
    layer0_outputs(7760) <= '1';
    layer0_outputs(7761) <= not((inputs(132)) or (inputs(134)));
    layer0_outputs(7762) <= (inputs(118)) and not (inputs(147));
    layer0_outputs(7763) <= inputs(56);
    layer0_outputs(7764) <= not((inputs(239)) xor (inputs(20)));
    layer0_outputs(7765) <= '1';
    layer0_outputs(7766) <= not((inputs(46)) or (inputs(76)));
    layer0_outputs(7767) <= (inputs(102)) or (inputs(149));
    layer0_outputs(7768) <= not(inputs(233)) or (inputs(134));
    layer0_outputs(7769) <= '1';
    layer0_outputs(7770) <= not(inputs(187)) or (inputs(78));
    layer0_outputs(7771) <= (inputs(6)) or (inputs(36));
    layer0_outputs(7772) <= (inputs(31)) and not (inputs(39));
    layer0_outputs(7773) <= (inputs(4)) and (inputs(35));
    layer0_outputs(7774) <= '1';
    layer0_outputs(7775) <= not((inputs(86)) xor (inputs(80)));
    layer0_outputs(7776) <= (inputs(28)) xor (inputs(202));
    layer0_outputs(7777) <= '1';
    layer0_outputs(7778) <= (inputs(249)) and (inputs(122));
    layer0_outputs(7779) <= inputs(223);
    layer0_outputs(7780) <= not(inputs(103));
    layer0_outputs(7781) <= not((inputs(199)) xor (inputs(211)));
    layer0_outputs(7782) <= not((inputs(103)) or (inputs(24)));
    layer0_outputs(7783) <= not(inputs(136)) or (inputs(10));
    layer0_outputs(7784) <= not((inputs(25)) xor (inputs(160)));
    layer0_outputs(7785) <= not(inputs(124));
    layer0_outputs(7786) <= (inputs(195)) xor (inputs(127));
    layer0_outputs(7787) <= not((inputs(17)) xor (inputs(0)));
    layer0_outputs(7788) <= not((inputs(3)) xor (inputs(156)));
    layer0_outputs(7789) <= (inputs(1)) or (inputs(163));
    layer0_outputs(7790) <= (inputs(84)) and (inputs(234));
    layer0_outputs(7791) <= not((inputs(232)) and (inputs(95)));
    layer0_outputs(7792) <= not((inputs(10)) or (inputs(36)));
    layer0_outputs(7793) <= inputs(38);
    layer0_outputs(7794) <= not((inputs(36)) xor (inputs(181)));
    layer0_outputs(7795) <= '0';
    layer0_outputs(7796) <= not((inputs(206)) or (inputs(163)));
    layer0_outputs(7797) <= not(inputs(197)) or (inputs(134));
    layer0_outputs(7798) <= '0';
    layer0_outputs(7799) <= not(inputs(140)) or (inputs(249));
    layer0_outputs(7800) <= not(inputs(86));
    layer0_outputs(7801) <= not(inputs(121)) or (inputs(40));
    layer0_outputs(7802) <= inputs(55);
    layer0_outputs(7803) <= (inputs(131)) and not (inputs(84));
    layer0_outputs(7804) <= (inputs(73)) or (inputs(41));
    layer0_outputs(7805) <= not(inputs(66));
    layer0_outputs(7806) <= not((inputs(12)) and (inputs(36)));
    layer0_outputs(7807) <= (inputs(85)) and not (inputs(57));
    layer0_outputs(7808) <= inputs(72);
    layer0_outputs(7809) <= inputs(189);
    layer0_outputs(7810) <= (inputs(155)) or (inputs(173));
    layer0_outputs(7811) <= '0';
    layer0_outputs(7812) <= not(inputs(84)) or (inputs(221));
    layer0_outputs(7813) <= '1';
    layer0_outputs(7814) <= (inputs(229)) or (inputs(57));
    layer0_outputs(7815) <= (inputs(107)) or (inputs(171));
    layer0_outputs(7816) <= inputs(227);
    layer0_outputs(7817) <= not((inputs(120)) xor (inputs(14)));
    layer0_outputs(7818) <= '1';
    layer0_outputs(7819) <= not(inputs(118));
    layer0_outputs(7820) <= not(inputs(17));
    layer0_outputs(7821) <= '1';
    layer0_outputs(7822) <= inputs(66);
    layer0_outputs(7823) <= not((inputs(107)) xor (inputs(113)));
    layer0_outputs(7824) <= not((inputs(221)) and (inputs(225)));
    layer0_outputs(7825) <= (inputs(224)) and not (inputs(234));
    layer0_outputs(7826) <= not(inputs(85)) or (inputs(172));
    layer0_outputs(7827) <= (inputs(187)) and not (inputs(213));
    layer0_outputs(7828) <= not((inputs(80)) and (inputs(29)));
    layer0_outputs(7829) <= (inputs(245)) and (inputs(241));
    layer0_outputs(7830) <= not(inputs(104));
    layer0_outputs(7831) <= not((inputs(39)) or (inputs(72)));
    layer0_outputs(7832) <= '1';
    layer0_outputs(7833) <= (inputs(150)) or (inputs(107));
    layer0_outputs(7834) <= not(inputs(240));
    layer0_outputs(7835) <= inputs(10);
    layer0_outputs(7836) <= '0';
    layer0_outputs(7837) <= not(inputs(47)) or (inputs(3));
    layer0_outputs(7838) <= not((inputs(192)) or (inputs(241)));
    layer0_outputs(7839) <= not(inputs(69));
    layer0_outputs(7840) <= inputs(188);
    layer0_outputs(7841) <= inputs(155);
    layer0_outputs(7842) <= inputs(70);
    layer0_outputs(7843) <= not(inputs(158));
    layer0_outputs(7844) <= not((inputs(156)) xor (inputs(218)));
    layer0_outputs(7845) <= '1';
    layer0_outputs(7846) <= not(inputs(38));
    layer0_outputs(7847) <= (inputs(221)) and not (inputs(26));
    layer0_outputs(7848) <= '1';
    layer0_outputs(7849) <= not(inputs(108));
    layer0_outputs(7850) <= (inputs(33)) xor (inputs(86));
    layer0_outputs(7851) <= not(inputs(105)) or (inputs(0));
    layer0_outputs(7852) <= not(inputs(244)) or (inputs(92));
    layer0_outputs(7853) <= (inputs(27)) or (inputs(137));
    layer0_outputs(7854) <= not((inputs(90)) and (inputs(168)));
    layer0_outputs(7855) <= (inputs(136)) xor (inputs(23));
    layer0_outputs(7856) <= '1';
    layer0_outputs(7857) <= inputs(90);
    layer0_outputs(7858) <= (inputs(101)) and not (inputs(138));
    layer0_outputs(7859) <= not((inputs(181)) or (inputs(19)));
    layer0_outputs(7860) <= (inputs(13)) or (inputs(131));
    layer0_outputs(7861) <= (inputs(239)) or (inputs(98));
    layer0_outputs(7862) <= (inputs(130)) xor (inputs(205));
    layer0_outputs(7863) <= not(inputs(184)) or (inputs(244));
    layer0_outputs(7864) <= not((inputs(98)) and (inputs(82)));
    layer0_outputs(7865) <= (inputs(230)) or (inputs(244));
    layer0_outputs(7866) <= not((inputs(115)) and (inputs(193)));
    layer0_outputs(7867) <= not((inputs(201)) xor (inputs(196)));
    layer0_outputs(7868) <= not((inputs(159)) xor (inputs(231)));
    layer0_outputs(7869) <= not((inputs(175)) xor (inputs(48)));
    layer0_outputs(7870) <= not(inputs(47));
    layer0_outputs(7871) <= not(inputs(65)) or (inputs(99));
    layer0_outputs(7872) <= not(inputs(118));
    layer0_outputs(7873) <= not((inputs(149)) xor (inputs(111)));
    layer0_outputs(7874) <= (inputs(165)) and not (inputs(69));
    layer0_outputs(7875) <= not((inputs(229)) xor (inputs(22)));
    layer0_outputs(7876) <= inputs(142);
    layer0_outputs(7877) <= '1';
    layer0_outputs(7878) <= (inputs(134)) and (inputs(159));
    layer0_outputs(7879) <= not(inputs(105));
    layer0_outputs(7880) <= (inputs(218)) and not (inputs(14));
    layer0_outputs(7881) <= (inputs(183)) and not (inputs(91));
    layer0_outputs(7882) <= not((inputs(6)) xor (inputs(31)));
    layer0_outputs(7883) <= inputs(135);
    layer0_outputs(7884) <= not(inputs(100)) or (inputs(82));
    layer0_outputs(7885) <= not((inputs(112)) or (inputs(179)));
    layer0_outputs(7886) <= not((inputs(83)) and (inputs(160)));
    layer0_outputs(7887) <= not((inputs(52)) or (inputs(102)));
    layer0_outputs(7888) <= (inputs(14)) and not (inputs(150));
    layer0_outputs(7889) <= not((inputs(91)) xor (inputs(7)));
    layer0_outputs(7890) <= not((inputs(169)) xor (inputs(81)));
    layer0_outputs(7891) <= (inputs(193)) and (inputs(246));
    layer0_outputs(7892) <= inputs(27);
    layer0_outputs(7893) <= not((inputs(121)) and (inputs(56)));
    layer0_outputs(7894) <= inputs(175);
    layer0_outputs(7895) <= not(inputs(32)) or (inputs(56));
    layer0_outputs(7896) <= not(inputs(163));
    layer0_outputs(7897) <= '1';
    layer0_outputs(7898) <= not(inputs(119));
    layer0_outputs(7899) <= '0';
    layer0_outputs(7900) <= inputs(119);
    layer0_outputs(7901) <= not(inputs(148));
    layer0_outputs(7902) <= inputs(160);
    layer0_outputs(7903) <= not((inputs(71)) and (inputs(209)));
    layer0_outputs(7904) <= not(inputs(123));
    layer0_outputs(7905) <= (inputs(178)) xor (inputs(211));
    layer0_outputs(7906) <= (inputs(75)) and (inputs(57));
    layer0_outputs(7907) <= not((inputs(135)) or (inputs(119)));
    layer0_outputs(7908) <= inputs(101);
    layer0_outputs(7909) <= not((inputs(143)) xor (inputs(12)));
    layer0_outputs(7910) <= (inputs(243)) and not (inputs(222));
    layer0_outputs(7911) <= (inputs(255)) and not (inputs(40));
    layer0_outputs(7912) <= not((inputs(242)) and (inputs(68)));
    layer0_outputs(7913) <= inputs(168);
    layer0_outputs(7914) <= not((inputs(153)) or (inputs(27)));
    layer0_outputs(7915) <= (inputs(174)) or (inputs(179));
    layer0_outputs(7916) <= inputs(82);
    layer0_outputs(7917) <= inputs(130);
    layer0_outputs(7918) <= (inputs(254)) or (inputs(240));
    layer0_outputs(7919) <= not((inputs(208)) xor (inputs(201)));
    layer0_outputs(7920) <= not(inputs(138)) or (inputs(157));
    layer0_outputs(7921) <= not(inputs(131)) or (inputs(26));
    layer0_outputs(7922) <= '0';
    layer0_outputs(7923) <= (inputs(163)) and not (inputs(107));
    layer0_outputs(7924) <= (inputs(176)) xor (inputs(109));
    layer0_outputs(7925) <= not((inputs(218)) xor (inputs(231)));
    layer0_outputs(7926) <= (inputs(187)) and not (inputs(204));
    layer0_outputs(7927) <= not(inputs(210)) or (inputs(43));
    layer0_outputs(7928) <= '1';
    layer0_outputs(7929) <= not(inputs(138));
    layer0_outputs(7930) <= inputs(154);
    layer0_outputs(7931) <= (inputs(153)) and not (inputs(202));
    layer0_outputs(7932) <= not(inputs(121)) or (inputs(206));
    layer0_outputs(7933) <= '0';
    layer0_outputs(7934) <= not(inputs(89)) or (inputs(192));
    layer0_outputs(7935) <= inputs(92);
    layer0_outputs(7936) <= inputs(19);
    layer0_outputs(7937) <= (inputs(155)) xor (inputs(68));
    layer0_outputs(7938) <= not(inputs(252)) or (inputs(83));
    layer0_outputs(7939) <= not((inputs(59)) and (inputs(162)));
    layer0_outputs(7940) <= (inputs(54)) or (inputs(34));
    layer0_outputs(7941) <= (inputs(250)) xor (inputs(156));
    layer0_outputs(7942) <= not((inputs(186)) or (inputs(187)));
    layer0_outputs(7943) <= not((inputs(72)) or (inputs(103)));
    layer0_outputs(7944) <= not(inputs(148));
    layer0_outputs(7945) <= (inputs(218)) or (inputs(135));
    layer0_outputs(7946) <= (inputs(152)) and not (inputs(199));
    layer0_outputs(7947) <= not(inputs(179));
    layer0_outputs(7948) <= (inputs(126)) and (inputs(175));
    layer0_outputs(7949) <= (inputs(3)) and not (inputs(229));
    layer0_outputs(7950) <= not(inputs(255)) or (inputs(138));
    layer0_outputs(7951) <= not(inputs(169)) or (inputs(223));
    layer0_outputs(7952) <= not((inputs(171)) or (inputs(22)));
    layer0_outputs(7953) <= not((inputs(26)) or (inputs(138)));
    layer0_outputs(7954) <= not(inputs(166));
    layer0_outputs(7955) <= (inputs(180)) or (inputs(129));
    layer0_outputs(7956) <= (inputs(174)) and not (inputs(66));
    layer0_outputs(7957) <= not(inputs(199)) or (inputs(99));
    layer0_outputs(7958) <= '1';
    layer0_outputs(7959) <= (inputs(75)) and not (inputs(246));
    layer0_outputs(7960) <= '1';
    layer0_outputs(7961) <= '1';
    layer0_outputs(7962) <= not(inputs(240));
    layer0_outputs(7963) <= not(inputs(99)) or (inputs(43));
    layer0_outputs(7964) <= not(inputs(112)) or (inputs(240));
    layer0_outputs(7965) <= (inputs(147)) and not (inputs(177));
    layer0_outputs(7966) <= '0';
    layer0_outputs(7967) <= not(inputs(7));
    layer0_outputs(7968) <= not((inputs(76)) or (inputs(215)));
    layer0_outputs(7969) <= inputs(162);
    layer0_outputs(7970) <= (inputs(113)) or (inputs(12));
    layer0_outputs(7971) <= (inputs(186)) and not (inputs(154));
    layer0_outputs(7972) <= inputs(92);
    layer0_outputs(7973) <= not(inputs(42));
    layer0_outputs(7974) <= '0';
    layer0_outputs(7975) <= not(inputs(197));
    layer0_outputs(7976) <= not(inputs(242)) or (inputs(96));
    layer0_outputs(7977) <= not((inputs(216)) and (inputs(114)));
    layer0_outputs(7978) <= not(inputs(75));
    layer0_outputs(7979) <= not(inputs(86));
    layer0_outputs(7980) <= (inputs(180)) or (inputs(78));
    layer0_outputs(7981) <= not(inputs(146)) or (inputs(4));
    layer0_outputs(7982) <= (inputs(41)) or (inputs(166));
    layer0_outputs(7983) <= not(inputs(165));
    layer0_outputs(7984) <= not((inputs(228)) xor (inputs(55)));
    layer0_outputs(7985) <= not(inputs(173));
    layer0_outputs(7986) <= (inputs(239)) and not (inputs(242));
    layer0_outputs(7987) <= not((inputs(2)) or (inputs(66)));
    layer0_outputs(7988) <= not(inputs(153)) or (inputs(175));
    layer0_outputs(7989) <= not((inputs(152)) xor (inputs(21)));
    layer0_outputs(7990) <= inputs(255);
    layer0_outputs(7991) <= '1';
    layer0_outputs(7992) <= '0';
    layer0_outputs(7993) <= inputs(31);
    layer0_outputs(7994) <= (inputs(144)) xor (inputs(142));
    layer0_outputs(7995) <= not(inputs(108)) or (inputs(22));
    layer0_outputs(7996) <= not((inputs(41)) and (inputs(210)));
    layer0_outputs(7997) <= (inputs(13)) xor (inputs(97));
    layer0_outputs(7998) <= (inputs(168)) and not (inputs(93));
    layer0_outputs(7999) <= inputs(242);
    layer0_outputs(8000) <= not(inputs(192)) or (inputs(153));
    layer0_outputs(8001) <= not(inputs(6)) or (inputs(237));
    layer0_outputs(8002) <= not((inputs(115)) xor (inputs(200)));
    layer0_outputs(8003) <= '1';
    layer0_outputs(8004) <= (inputs(80)) or (inputs(10));
    layer0_outputs(8005) <= '1';
    layer0_outputs(8006) <= (inputs(98)) or (inputs(143));
    layer0_outputs(8007) <= '0';
    layer0_outputs(8008) <= not(inputs(143)) or (inputs(199));
    layer0_outputs(8009) <= '1';
    layer0_outputs(8010) <= not((inputs(232)) xor (inputs(112)));
    layer0_outputs(8011) <= '1';
    layer0_outputs(8012) <= (inputs(32)) or (inputs(109));
    layer0_outputs(8013) <= not(inputs(169));
    layer0_outputs(8014) <= not((inputs(210)) and (inputs(140)));
    layer0_outputs(8015) <= (inputs(75)) and (inputs(78));
    layer0_outputs(8016) <= (inputs(92)) and not (inputs(236));
    layer0_outputs(8017) <= not((inputs(196)) xor (inputs(80)));
    layer0_outputs(8018) <= inputs(37);
    layer0_outputs(8019) <= not(inputs(177));
    layer0_outputs(8020) <= inputs(142);
    layer0_outputs(8021) <= '1';
    layer0_outputs(8022) <= (inputs(223)) and not (inputs(160));
    layer0_outputs(8023) <= '0';
    layer0_outputs(8024) <= not((inputs(13)) or (inputs(135)));
    layer0_outputs(8025) <= not((inputs(216)) and (inputs(168)));
    layer0_outputs(8026) <= (inputs(95)) and (inputs(81));
    layer0_outputs(8027) <= (inputs(252)) or (inputs(151));
    layer0_outputs(8028) <= not(inputs(158));
    layer0_outputs(8029) <= (inputs(21)) and not (inputs(98));
    layer0_outputs(8030) <= (inputs(60)) or (inputs(198));
    layer0_outputs(8031) <= not((inputs(5)) xor (inputs(160)));
    layer0_outputs(8032) <= (inputs(129)) or (inputs(171));
    layer0_outputs(8033) <= (inputs(68)) xor (inputs(82));
    layer0_outputs(8034) <= not(inputs(159)) or (inputs(253));
    layer0_outputs(8035) <= '1';
    layer0_outputs(8036) <= inputs(150);
    layer0_outputs(8037) <= inputs(33);
    layer0_outputs(8038) <= '1';
    layer0_outputs(8039) <= not(inputs(85));
    layer0_outputs(8040) <= '1';
    layer0_outputs(8041) <= not(inputs(217)) or (inputs(133));
    layer0_outputs(8042) <= (inputs(48)) xor (inputs(176));
    layer0_outputs(8043) <= (inputs(87)) and not (inputs(81));
    layer0_outputs(8044) <= not((inputs(19)) or (inputs(199)));
    layer0_outputs(8045) <= inputs(76);
    layer0_outputs(8046) <= not((inputs(2)) xor (inputs(187)));
    layer0_outputs(8047) <= not(inputs(37));
    layer0_outputs(8048) <= not(inputs(76)) or (inputs(40));
    layer0_outputs(8049) <= '0';
    layer0_outputs(8050) <= (inputs(66)) and not (inputs(96));
    layer0_outputs(8051) <= (inputs(251)) and not (inputs(247));
    layer0_outputs(8052) <= (inputs(86)) or (inputs(94));
    layer0_outputs(8053) <= not((inputs(110)) xor (inputs(172)));
    layer0_outputs(8054) <= not((inputs(141)) and (inputs(13)));
    layer0_outputs(8055) <= not(inputs(215)) or (inputs(244));
    layer0_outputs(8056) <= '1';
    layer0_outputs(8057) <= not(inputs(106)) or (inputs(25));
    layer0_outputs(8058) <= '0';
    layer0_outputs(8059) <= (inputs(243)) and (inputs(50));
    layer0_outputs(8060) <= not((inputs(214)) and (inputs(214)));
    layer0_outputs(8061) <= not((inputs(232)) xor (inputs(49)));
    layer0_outputs(8062) <= not((inputs(174)) xor (inputs(237)));
    layer0_outputs(8063) <= (inputs(34)) and not (inputs(61));
    layer0_outputs(8064) <= not(inputs(88));
    layer0_outputs(8065) <= not(inputs(83));
    layer0_outputs(8066) <= inputs(118);
    layer0_outputs(8067) <= (inputs(8)) or (inputs(157));
    layer0_outputs(8068) <= inputs(138);
    layer0_outputs(8069) <= (inputs(22)) and not (inputs(98));
    layer0_outputs(8070) <= not(inputs(22)) or (inputs(169));
    layer0_outputs(8071) <= not(inputs(109));
    layer0_outputs(8072) <= not(inputs(168)) or (inputs(147));
    layer0_outputs(8073) <= not((inputs(7)) and (inputs(182)));
    layer0_outputs(8074) <= not((inputs(151)) or (inputs(24)));
    layer0_outputs(8075) <= not((inputs(159)) xor (inputs(242)));
    layer0_outputs(8076) <= '0';
    layer0_outputs(8077) <= (inputs(151)) and (inputs(17));
    layer0_outputs(8078) <= inputs(197);
    layer0_outputs(8079) <= not(inputs(121)) or (inputs(92));
    layer0_outputs(8080) <= not(inputs(164));
    layer0_outputs(8081) <= not((inputs(120)) or (inputs(209)));
    layer0_outputs(8082) <= not((inputs(97)) or (inputs(220)));
    layer0_outputs(8083) <= inputs(102);
    layer0_outputs(8084) <= (inputs(93)) or (inputs(118));
    layer0_outputs(8085) <= not(inputs(236));
    layer0_outputs(8086) <= not(inputs(82)) or (inputs(82));
    layer0_outputs(8087) <= not((inputs(83)) or (inputs(137)));
    layer0_outputs(8088) <= not((inputs(12)) xor (inputs(105)));
    layer0_outputs(8089) <= not((inputs(69)) xor (inputs(184)));
    layer0_outputs(8090) <= (inputs(109)) and not (inputs(22));
    layer0_outputs(8091) <= not((inputs(93)) or (inputs(146)));
    layer0_outputs(8092) <= not((inputs(230)) or (inputs(154)));
    layer0_outputs(8093) <= not((inputs(105)) or (inputs(90)));
    layer0_outputs(8094) <= '0';
    layer0_outputs(8095) <= not(inputs(96)) or (inputs(209));
    layer0_outputs(8096) <= not(inputs(84));
    layer0_outputs(8097) <= (inputs(199)) or (inputs(177));
    layer0_outputs(8098) <= not(inputs(138)) or (inputs(144));
    layer0_outputs(8099) <= not(inputs(212));
    layer0_outputs(8100) <= (inputs(56)) or (inputs(133));
    layer0_outputs(8101) <= not(inputs(106));
    layer0_outputs(8102) <= not((inputs(233)) and (inputs(129)));
    layer0_outputs(8103) <= not(inputs(24)) or (inputs(142));
    layer0_outputs(8104) <= not(inputs(127)) or (inputs(3));
    layer0_outputs(8105) <= not((inputs(55)) or (inputs(238)));
    layer0_outputs(8106) <= not(inputs(109));
    layer0_outputs(8107) <= '1';
    layer0_outputs(8108) <= not((inputs(204)) xor (inputs(213)));
    layer0_outputs(8109) <= (inputs(23)) xor (inputs(181));
    layer0_outputs(8110) <= inputs(70);
    layer0_outputs(8111) <= (inputs(255)) and not (inputs(207));
    layer0_outputs(8112) <= inputs(41);
    layer0_outputs(8113) <= (inputs(74)) and (inputs(72));
    layer0_outputs(8114) <= not((inputs(174)) or (inputs(223)));
    layer0_outputs(8115) <= (inputs(238)) and not (inputs(127));
    layer0_outputs(8116) <= not(inputs(194));
    layer0_outputs(8117) <= not(inputs(90));
    layer0_outputs(8118) <= (inputs(231)) or (inputs(103));
    layer0_outputs(8119) <= not(inputs(225));
    layer0_outputs(8120) <= '1';
    layer0_outputs(8121) <= not((inputs(146)) xor (inputs(38)));
    layer0_outputs(8122) <= (inputs(147)) and (inputs(118));
    layer0_outputs(8123) <= not(inputs(94)) or (inputs(177));
    layer0_outputs(8124) <= '1';
    layer0_outputs(8125) <= (inputs(215)) and not (inputs(101));
    layer0_outputs(8126) <= '1';
    layer0_outputs(8127) <= inputs(155);
    layer0_outputs(8128) <= not(inputs(117));
    layer0_outputs(8129) <= not((inputs(243)) xor (inputs(54)));
    layer0_outputs(8130) <= (inputs(37)) and (inputs(254));
    layer0_outputs(8131) <= (inputs(122)) and not (inputs(94));
    layer0_outputs(8132) <= not(inputs(91));
    layer0_outputs(8133) <= not((inputs(39)) or (inputs(31)));
    layer0_outputs(8134) <= '0';
    layer0_outputs(8135) <= not(inputs(207)) or (inputs(221));
    layer0_outputs(8136) <= not((inputs(35)) or (inputs(110)));
    layer0_outputs(8137) <= inputs(14);
    layer0_outputs(8138) <= (inputs(229)) and (inputs(135));
    layer0_outputs(8139) <= (inputs(215)) and not (inputs(167));
    layer0_outputs(8140) <= (inputs(196)) or (inputs(52));
    layer0_outputs(8141) <= not((inputs(214)) xor (inputs(95)));
    layer0_outputs(8142) <= '0';
    layer0_outputs(8143) <= (inputs(167)) and not (inputs(64));
    layer0_outputs(8144) <= (inputs(165)) or (inputs(213));
    layer0_outputs(8145) <= inputs(59);
    layer0_outputs(8146) <= not((inputs(48)) xor (inputs(250)));
    layer0_outputs(8147) <= not((inputs(245)) xor (inputs(4)));
    layer0_outputs(8148) <= inputs(171);
    layer0_outputs(8149) <= not(inputs(66)) or (inputs(156));
    layer0_outputs(8150) <= not(inputs(131));
    layer0_outputs(8151) <= not((inputs(160)) xor (inputs(185)));
    layer0_outputs(8152) <= '0';
    layer0_outputs(8153) <= not((inputs(9)) or (inputs(53)));
    layer0_outputs(8154) <= (inputs(207)) and (inputs(107));
    layer0_outputs(8155) <= inputs(60);
    layer0_outputs(8156) <= inputs(108);
    layer0_outputs(8157) <= inputs(15);
    layer0_outputs(8158) <= not((inputs(155)) and (inputs(200)));
    layer0_outputs(8159) <= inputs(154);
    layer0_outputs(8160) <= (inputs(199)) and (inputs(224));
    layer0_outputs(8161) <= not(inputs(49)) or (inputs(69));
    layer0_outputs(8162) <= '0';
    layer0_outputs(8163) <= (inputs(240)) and not (inputs(191));
    layer0_outputs(8164) <= not(inputs(53)) or (inputs(251));
    layer0_outputs(8165) <= (inputs(56)) and not (inputs(50));
    layer0_outputs(8166) <= not((inputs(86)) xor (inputs(229)));
    layer0_outputs(8167) <= not((inputs(2)) and (inputs(71)));
    layer0_outputs(8168) <= '1';
    layer0_outputs(8169) <= (inputs(255)) or (inputs(142));
    layer0_outputs(8170) <= not((inputs(25)) xor (inputs(90)));
    layer0_outputs(8171) <= not(inputs(110));
    layer0_outputs(8172) <= (inputs(212)) xor (inputs(110));
    layer0_outputs(8173) <= inputs(18);
    layer0_outputs(8174) <= (inputs(47)) or (inputs(38));
    layer0_outputs(8175) <= (inputs(22)) or (inputs(78));
    layer0_outputs(8176) <= not(inputs(205));
    layer0_outputs(8177) <= inputs(111);
    layer0_outputs(8178) <= inputs(139);
    layer0_outputs(8179) <= inputs(240);
    layer0_outputs(8180) <= (inputs(31)) or (inputs(236));
    layer0_outputs(8181) <= (inputs(224)) and not (inputs(126));
    layer0_outputs(8182) <= not((inputs(207)) and (inputs(61)));
    layer0_outputs(8183) <= inputs(168);
    layer0_outputs(8184) <= inputs(250);
    layer0_outputs(8185) <= (inputs(179)) and not (inputs(89));
    layer0_outputs(8186) <= not(inputs(16)) or (inputs(170));
    layer0_outputs(8187) <= (inputs(110)) and (inputs(107));
    layer0_outputs(8188) <= (inputs(200)) and not (inputs(177));
    layer0_outputs(8189) <= not(inputs(4)) or (inputs(134));
    layer0_outputs(8190) <= not(inputs(188)) or (inputs(253));
    layer0_outputs(8191) <= '1';
    layer0_outputs(8192) <= not((inputs(78)) xor (inputs(19)));
    layer0_outputs(8193) <= not((inputs(54)) or (inputs(74)));
    layer0_outputs(8194) <= inputs(104);
    layer0_outputs(8195) <= not((inputs(73)) and (inputs(142)));
    layer0_outputs(8196) <= inputs(67);
    layer0_outputs(8197) <= '0';
    layer0_outputs(8198) <= not(inputs(159));
    layer0_outputs(8199) <= (inputs(145)) xor (inputs(29));
    layer0_outputs(8200) <= not(inputs(159)) or (inputs(217));
    layer0_outputs(8201) <= not(inputs(188)) or (inputs(35));
    layer0_outputs(8202) <= '1';
    layer0_outputs(8203) <= (inputs(71)) xor (inputs(77));
    layer0_outputs(8204) <= (inputs(101)) or (inputs(97));
    layer0_outputs(8205) <= inputs(169);
    layer0_outputs(8206) <= (inputs(217)) and not (inputs(3));
    layer0_outputs(8207) <= (inputs(172)) or (inputs(194));
    layer0_outputs(8208) <= inputs(89);
    layer0_outputs(8209) <= inputs(46);
    layer0_outputs(8210) <= not((inputs(29)) xor (inputs(199)));
    layer0_outputs(8211) <= not(inputs(192));
    layer0_outputs(8212) <= not(inputs(113)) or (inputs(176));
    layer0_outputs(8213) <= (inputs(190)) and not (inputs(210));
    layer0_outputs(8214) <= not((inputs(169)) xor (inputs(64)));
    layer0_outputs(8215) <= not(inputs(222)) or (inputs(128));
    layer0_outputs(8216) <= not(inputs(162));
    layer0_outputs(8217) <= '1';
    layer0_outputs(8218) <= inputs(108);
    layer0_outputs(8219) <= not(inputs(206)) or (inputs(125));
    layer0_outputs(8220) <= '1';
    layer0_outputs(8221) <= (inputs(119)) and not (inputs(205));
    layer0_outputs(8222) <= not(inputs(48)) or (inputs(46));
    layer0_outputs(8223) <= (inputs(63)) xor (inputs(219));
    layer0_outputs(8224) <= not(inputs(24)) or (inputs(176));
    layer0_outputs(8225) <= not(inputs(71));
    layer0_outputs(8226) <= inputs(19);
    layer0_outputs(8227) <= (inputs(48)) or (inputs(252));
    layer0_outputs(8228) <= inputs(240);
    layer0_outputs(8229) <= (inputs(64)) and (inputs(161));
    layer0_outputs(8230) <= inputs(160);
    layer0_outputs(8231) <= not(inputs(111)) or (inputs(178));
    layer0_outputs(8232) <= (inputs(226)) xor (inputs(180));
    layer0_outputs(8233) <= (inputs(205)) xor (inputs(59));
    layer0_outputs(8234) <= inputs(100);
    layer0_outputs(8235) <= (inputs(133)) or (inputs(62));
    layer0_outputs(8236) <= not(inputs(58)) or (inputs(34));
    layer0_outputs(8237) <= (inputs(134)) and (inputs(126));
    layer0_outputs(8238) <= inputs(140);
    layer0_outputs(8239) <= (inputs(158)) xor (inputs(252));
    layer0_outputs(8240) <= not(inputs(247)) or (inputs(99));
    layer0_outputs(8241) <= not((inputs(154)) or (inputs(117)));
    layer0_outputs(8242) <= not(inputs(156));
    layer0_outputs(8243) <= not(inputs(107));
    layer0_outputs(8244) <= not((inputs(208)) and (inputs(97)));
    layer0_outputs(8245) <= '0';
    layer0_outputs(8246) <= inputs(188);
    layer0_outputs(8247) <= not((inputs(116)) xor (inputs(3)));
    layer0_outputs(8248) <= '1';
    layer0_outputs(8249) <= inputs(106);
    layer0_outputs(8250) <= not((inputs(225)) xor (inputs(202)));
    layer0_outputs(8251) <= not(inputs(148)) or (inputs(110));
    layer0_outputs(8252) <= (inputs(166)) and not (inputs(66));
    layer0_outputs(8253) <= (inputs(165)) xor (inputs(225));
    layer0_outputs(8254) <= not(inputs(27)) or (inputs(234));
    layer0_outputs(8255) <= (inputs(194)) xor (inputs(175));
    layer0_outputs(8256) <= not(inputs(37));
    layer0_outputs(8257) <= not(inputs(204));
    layer0_outputs(8258) <= (inputs(55)) or (inputs(52));
    layer0_outputs(8259) <= '1';
    layer0_outputs(8260) <= (inputs(199)) xor (inputs(5));
    layer0_outputs(8261) <= not(inputs(188)) or (inputs(109));
    layer0_outputs(8262) <= (inputs(219)) or (inputs(145));
    layer0_outputs(8263) <= not(inputs(218));
    layer0_outputs(8264) <= '0';
    layer0_outputs(8265) <= not(inputs(37)) or (inputs(13));
    layer0_outputs(8266) <= (inputs(88)) or (inputs(79));
    layer0_outputs(8267) <= (inputs(114)) or (inputs(91));
    layer0_outputs(8268) <= (inputs(42)) and not (inputs(143));
    layer0_outputs(8269) <= not(inputs(197)) or (inputs(207));
    layer0_outputs(8270) <= not(inputs(88));
    layer0_outputs(8271) <= not((inputs(96)) or (inputs(219)));
    layer0_outputs(8272) <= (inputs(116)) or (inputs(45));
    layer0_outputs(8273) <= not((inputs(132)) or (inputs(131)));
    layer0_outputs(8274) <= '1';
    layer0_outputs(8275) <= not(inputs(63));
    layer0_outputs(8276) <= (inputs(93)) and (inputs(67));
    layer0_outputs(8277) <= '1';
    layer0_outputs(8278) <= not(inputs(82));
    layer0_outputs(8279) <= not((inputs(142)) or (inputs(159)));
    layer0_outputs(8280) <= not(inputs(225)) or (inputs(11));
    layer0_outputs(8281) <= inputs(53);
    layer0_outputs(8282) <= (inputs(182)) and not (inputs(80));
    layer0_outputs(8283) <= '1';
    layer0_outputs(8284) <= not(inputs(165));
    layer0_outputs(8285) <= not(inputs(55));
    layer0_outputs(8286) <= (inputs(241)) xor (inputs(233));
    layer0_outputs(8287) <= not((inputs(245)) and (inputs(245)));
    layer0_outputs(8288) <= '1';
    layer0_outputs(8289) <= not(inputs(134)) or (inputs(35));
    layer0_outputs(8290) <= not(inputs(77));
    layer0_outputs(8291) <= (inputs(131)) or (inputs(45));
    layer0_outputs(8292) <= not((inputs(168)) xor (inputs(170)));
    layer0_outputs(8293) <= not(inputs(72)) or (inputs(193));
    layer0_outputs(8294) <= not(inputs(104)) or (inputs(223));
    layer0_outputs(8295) <= not(inputs(147)) or (inputs(48));
    layer0_outputs(8296) <= not((inputs(252)) and (inputs(113)));
    layer0_outputs(8297) <= (inputs(28)) and (inputs(206));
    layer0_outputs(8298) <= (inputs(123)) or (inputs(124));
    layer0_outputs(8299) <= (inputs(108)) and (inputs(244));
    layer0_outputs(8300) <= (inputs(143)) xor (inputs(200));
    layer0_outputs(8301) <= not((inputs(219)) xor (inputs(70)));
    layer0_outputs(8302) <= (inputs(38)) and not (inputs(249));
    layer0_outputs(8303) <= not(inputs(194));
    layer0_outputs(8304) <= not((inputs(158)) or (inputs(224)));
    layer0_outputs(8305) <= not((inputs(137)) xor (inputs(53)));
    layer0_outputs(8306) <= '1';
    layer0_outputs(8307) <= not(inputs(208));
    layer0_outputs(8308) <= inputs(136);
    layer0_outputs(8309) <= (inputs(227)) or (inputs(254));
    layer0_outputs(8310) <= '1';
    layer0_outputs(8311) <= (inputs(222)) and not (inputs(21));
    layer0_outputs(8312) <= not(inputs(28)) or (inputs(63));
    layer0_outputs(8313) <= inputs(211);
    layer0_outputs(8314) <= (inputs(70)) or (inputs(203));
    layer0_outputs(8315) <= not((inputs(54)) or (inputs(211)));
    layer0_outputs(8316) <= not(inputs(249)) or (inputs(72));
    layer0_outputs(8317) <= (inputs(230)) or (inputs(162));
    layer0_outputs(8318) <= not((inputs(21)) or (inputs(200)));
    layer0_outputs(8319) <= (inputs(120)) and not (inputs(165));
    layer0_outputs(8320) <= not(inputs(41)) or (inputs(213));
    layer0_outputs(8321) <= not((inputs(49)) and (inputs(254)));
    layer0_outputs(8322) <= '1';
    layer0_outputs(8323) <= not((inputs(16)) or (inputs(75)));
    layer0_outputs(8324) <= not((inputs(138)) xor (inputs(98)));
    layer0_outputs(8325) <= not(inputs(200));
    layer0_outputs(8326) <= not(inputs(145)) or (inputs(206));
    layer0_outputs(8327) <= '1';
    layer0_outputs(8328) <= not((inputs(181)) xor (inputs(218)));
    layer0_outputs(8329) <= '0';
    layer0_outputs(8330) <= inputs(6);
    layer0_outputs(8331) <= not((inputs(25)) xor (inputs(112)));
    layer0_outputs(8332) <= not((inputs(141)) and (inputs(35)));
    layer0_outputs(8333) <= not(inputs(160));
    layer0_outputs(8334) <= (inputs(167)) and not (inputs(155));
    layer0_outputs(8335) <= not(inputs(222)) or (inputs(43));
    layer0_outputs(8336) <= (inputs(33)) xor (inputs(125));
    layer0_outputs(8337) <= (inputs(25)) and not (inputs(222));
    layer0_outputs(8338) <= inputs(121);
    layer0_outputs(8339) <= (inputs(250)) or (inputs(52));
    layer0_outputs(8340) <= not(inputs(39)) or (inputs(248));
    layer0_outputs(8341) <= (inputs(56)) and not (inputs(242));
    layer0_outputs(8342) <= not(inputs(116));
    layer0_outputs(8343) <= not(inputs(23));
    layer0_outputs(8344) <= not((inputs(124)) or (inputs(123)));
    layer0_outputs(8345) <= not(inputs(150));
    layer0_outputs(8346) <= not(inputs(237)) or (inputs(90));
    layer0_outputs(8347) <= inputs(107);
    layer0_outputs(8348) <= not((inputs(14)) xor (inputs(136)));
    layer0_outputs(8349) <= not(inputs(51));
    layer0_outputs(8350) <= inputs(182);
    layer0_outputs(8351) <= not(inputs(247)) or (inputs(44));
    layer0_outputs(8352) <= not(inputs(254));
    layer0_outputs(8353) <= (inputs(82)) or (inputs(245));
    layer0_outputs(8354) <= not((inputs(136)) xor (inputs(143)));
    layer0_outputs(8355) <= not(inputs(116));
    layer0_outputs(8356) <= not(inputs(89));
    layer0_outputs(8357) <= '0';
    layer0_outputs(8358) <= not((inputs(97)) xor (inputs(131)));
    layer0_outputs(8359) <= '0';
    layer0_outputs(8360) <= inputs(55);
    layer0_outputs(8361) <= not(inputs(132)) or (inputs(174));
    layer0_outputs(8362) <= inputs(104);
    layer0_outputs(8363) <= not(inputs(242)) or (inputs(168));
    layer0_outputs(8364) <= not(inputs(111)) or (inputs(47));
    layer0_outputs(8365) <= (inputs(150)) and not (inputs(25));
    layer0_outputs(8366) <= (inputs(49)) or (inputs(233));
    layer0_outputs(8367) <= not((inputs(163)) or (inputs(206)));
    layer0_outputs(8368) <= inputs(200);
    layer0_outputs(8369) <= '1';
    layer0_outputs(8370) <= '1';
    layer0_outputs(8371) <= not(inputs(73));
    layer0_outputs(8372) <= inputs(27);
    layer0_outputs(8373) <= not((inputs(22)) xor (inputs(61)));
    layer0_outputs(8374) <= '0';
    layer0_outputs(8375) <= not(inputs(105));
    layer0_outputs(8376) <= not((inputs(154)) or (inputs(233)));
    layer0_outputs(8377) <= (inputs(65)) and (inputs(205));
    layer0_outputs(8378) <= not(inputs(83));
    layer0_outputs(8379) <= not(inputs(227)) or (inputs(18));
    layer0_outputs(8380) <= (inputs(30)) and not (inputs(33));
    layer0_outputs(8381) <= not(inputs(130)) or (inputs(64));
    layer0_outputs(8382) <= not(inputs(177)) or (inputs(249));
    layer0_outputs(8383) <= inputs(130);
    layer0_outputs(8384) <= (inputs(106)) xor (inputs(190));
    layer0_outputs(8385) <= not((inputs(143)) and (inputs(219)));
    layer0_outputs(8386) <= (inputs(86)) and not (inputs(150));
    layer0_outputs(8387) <= inputs(27);
    layer0_outputs(8388) <= not(inputs(89));
    layer0_outputs(8389) <= (inputs(229)) or (inputs(139));
    layer0_outputs(8390) <= (inputs(216)) and (inputs(34));
    layer0_outputs(8391) <= (inputs(92)) and (inputs(158));
    layer0_outputs(8392) <= inputs(28);
    layer0_outputs(8393) <= not(inputs(89));
    layer0_outputs(8394) <= (inputs(54)) or (inputs(185));
    layer0_outputs(8395) <= '1';
    layer0_outputs(8396) <= '1';
    layer0_outputs(8397) <= '1';
    layer0_outputs(8398) <= not((inputs(45)) and (inputs(40)));
    layer0_outputs(8399) <= not((inputs(241)) and (inputs(176)));
    layer0_outputs(8400) <= not((inputs(46)) and (inputs(20)));
    layer0_outputs(8401) <= not(inputs(3)) or (inputs(207));
    layer0_outputs(8402) <= inputs(213);
    layer0_outputs(8403) <= (inputs(106)) xor (inputs(124));
    layer0_outputs(8404) <= '0';
    layer0_outputs(8405) <= not(inputs(117)) or (inputs(244));
    layer0_outputs(8406) <= (inputs(196)) or (inputs(211));
    layer0_outputs(8407) <= (inputs(238)) and (inputs(70));
    layer0_outputs(8408) <= not((inputs(137)) or (inputs(65)));
    layer0_outputs(8409) <= inputs(0);
    layer0_outputs(8410) <= inputs(226);
    layer0_outputs(8411) <= not(inputs(218)) or (inputs(30));
    layer0_outputs(8412) <= inputs(62);
    layer0_outputs(8413) <= inputs(78);
    layer0_outputs(8414) <= (inputs(73)) or (inputs(172));
    layer0_outputs(8415) <= inputs(15);
    layer0_outputs(8416) <= (inputs(43)) and (inputs(9));
    layer0_outputs(8417) <= not(inputs(135)) or (inputs(223));
    layer0_outputs(8418) <= not(inputs(134)) or (inputs(107));
    layer0_outputs(8419) <= (inputs(207)) and not (inputs(44));
    layer0_outputs(8420) <= (inputs(21)) and not (inputs(46));
    layer0_outputs(8421) <= (inputs(140)) and not (inputs(188));
    layer0_outputs(8422) <= not((inputs(249)) or (inputs(201)));
    layer0_outputs(8423) <= not((inputs(102)) or (inputs(27)));
    layer0_outputs(8424) <= inputs(143);
    layer0_outputs(8425) <= inputs(136);
    layer0_outputs(8426) <= (inputs(179)) or (inputs(239));
    layer0_outputs(8427) <= not(inputs(1));
    layer0_outputs(8428) <= not(inputs(67)) or (inputs(98));
    layer0_outputs(8429) <= '1';
    layer0_outputs(8430) <= '1';
    layer0_outputs(8431) <= not(inputs(116)) or (inputs(39));
    layer0_outputs(8432) <= (inputs(67)) xor (inputs(46));
    layer0_outputs(8433) <= (inputs(99)) xor (inputs(132));
    layer0_outputs(8434) <= not((inputs(111)) xor (inputs(73)));
    layer0_outputs(8435) <= '0';
    layer0_outputs(8436) <= (inputs(122)) and not (inputs(158));
    layer0_outputs(8437) <= not(inputs(180));
    layer0_outputs(8438) <= not(inputs(104)) or (inputs(150));
    layer0_outputs(8439) <= not(inputs(175));
    layer0_outputs(8440) <= '1';
    layer0_outputs(8441) <= not(inputs(250)) or (inputs(3));
    layer0_outputs(8442) <= not(inputs(195)) or (inputs(133));
    layer0_outputs(8443) <= (inputs(212)) xor (inputs(197));
    layer0_outputs(8444) <= not((inputs(137)) or (inputs(5)));
    layer0_outputs(8445) <= '0';
    layer0_outputs(8446) <= not((inputs(1)) or (inputs(231)));
    layer0_outputs(8447) <= '0';
    layer0_outputs(8448) <= not(inputs(49)) or (inputs(68));
    layer0_outputs(8449) <= inputs(208);
    layer0_outputs(8450) <= (inputs(177)) and not (inputs(29));
    layer0_outputs(8451) <= (inputs(168)) and not (inputs(190));
    layer0_outputs(8452) <= '0';
    layer0_outputs(8453) <= not((inputs(38)) xor (inputs(93)));
    layer0_outputs(8454) <= inputs(220);
    layer0_outputs(8455) <= '0';
    layer0_outputs(8456) <= not(inputs(196));
    layer0_outputs(8457) <= not((inputs(117)) or (inputs(125)));
    layer0_outputs(8458) <= not((inputs(40)) or (inputs(0)));
    layer0_outputs(8459) <= (inputs(90)) and (inputs(139));
    layer0_outputs(8460) <= not((inputs(9)) or (inputs(55)));
    layer0_outputs(8461) <= not((inputs(159)) or (inputs(153)));
    layer0_outputs(8462) <= not(inputs(137));
    layer0_outputs(8463) <= (inputs(114)) or (inputs(56));
    layer0_outputs(8464) <= inputs(25);
    layer0_outputs(8465) <= (inputs(103)) and not (inputs(208));
    layer0_outputs(8466) <= '0';
    layer0_outputs(8467) <= not((inputs(135)) or (inputs(195)));
    layer0_outputs(8468) <= inputs(79);
    layer0_outputs(8469) <= '0';
    layer0_outputs(8470) <= (inputs(157)) and (inputs(91));
    layer0_outputs(8471) <= '1';
    layer0_outputs(8472) <= not(inputs(26)) or (inputs(255));
    layer0_outputs(8473) <= '0';
    layer0_outputs(8474) <= not((inputs(29)) or (inputs(92)));
    layer0_outputs(8475) <= (inputs(83)) or (inputs(20));
    layer0_outputs(8476) <= '0';
    layer0_outputs(8477) <= (inputs(232)) and not (inputs(215));
    layer0_outputs(8478) <= (inputs(219)) or (inputs(130));
    layer0_outputs(8479) <= inputs(118);
    layer0_outputs(8480) <= (inputs(252)) or (inputs(228));
    layer0_outputs(8481) <= not((inputs(174)) or (inputs(167)));
    layer0_outputs(8482) <= not((inputs(238)) xor (inputs(101)));
    layer0_outputs(8483) <= inputs(252);
    layer0_outputs(8484) <= not(inputs(126));
    layer0_outputs(8485) <= (inputs(193)) and (inputs(223));
    layer0_outputs(8486) <= (inputs(223)) or (inputs(224));
    layer0_outputs(8487) <= not((inputs(20)) or (inputs(236)));
    layer0_outputs(8488) <= not(inputs(218));
    layer0_outputs(8489) <= (inputs(193)) or (inputs(125));
    layer0_outputs(8490) <= (inputs(118)) or (inputs(166));
    layer0_outputs(8491) <= '0';
    layer0_outputs(8492) <= not(inputs(100));
    layer0_outputs(8493) <= not((inputs(183)) or (inputs(243)));
    layer0_outputs(8494) <= (inputs(132)) and not (inputs(230));
    layer0_outputs(8495) <= (inputs(77)) or (inputs(172));
    layer0_outputs(8496) <= not((inputs(93)) and (inputs(217)));
    layer0_outputs(8497) <= '1';
    layer0_outputs(8498) <= not(inputs(132)) or (inputs(98));
    layer0_outputs(8499) <= not((inputs(176)) xor (inputs(107)));
    layer0_outputs(8500) <= (inputs(49)) or (inputs(68));
    layer0_outputs(8501) <= (inputs(235)) xor (inputs(142));
    layer0_outputs(8502) <= not(inputs(187)) or (inputs(11));
    layer0_outputs(8503) <= (inputs(70)) and (inputs(2));
    layer0_outputs(8504) <= (inputs(195)) or (inputs(35));
    layer0_outputs(8505) <= inputs(90);
    layer0_outputs(8506) <= inputs(102);
    layer0_outputs(8507) <= '1';
    layer0_outputs(8508) <= (inputs(0)) and not (inputs(31));
    layer0_outputs(8509) <= inputs(84);
    layer0_outputs(8510) <= inputs(47);
    layer0_outputs(8511) <= '0';
    layer0_outputs(8512) <= (inputs(136)) xor (inputs(158));
    layer0_outputs(8513) <= not(inputs(57));
    layer0_outputs(8514) <= inputs(144);
    layer0_outputs(8515) <= (inputs(119)) or (inputs(25));
    layer0_outputs(8516) <= not((inputs(6)) xor (inputs(17)));
    layer0_outputs(8517) <= (inputs(255)) and not (inputs(68));
    layer0_outputs(8518) <= '0';
    layer0_outputs(8519) <= not((inputs(139)) or (inputs(127)));
    layer0_outputs(8520) <= not(inputs(242));
    layer0_outputs(8521) <= (inputs(45)) or (inputs(67));
    layer0_outputs(8522) <= not((inputs(9)) or (inputs(208)));
    layer0_outputs(8523) <= inputs(247);
    layer0_outputs(8524) <= (inputs(131)) xor (inputs(166));
    layer0_outputs(8525) <= not((inputs(220)) or (inputs(164)));
    layer0_outputs(8526) <= (inputs(84)) or (inputs(252));
    layer0_outputs(8527) <= inputs(208);
    layer0_outputs(8528) <= not((inputs(132)) or (inputs(117)));
    layer0_outputs(8529) <= not((inputs(12)) and (inputs(20)));
    layer0_outputs(8530) <= inputs(122);
    layer0_outputs(8531) <= (inputs(194)) xor (inputs(165));
    layer0_outputs(8532) <= not(inputs(221));
    layer0_outputs(8533) <= not((inputs(249)) and (inputs(224)));
    layer0_outputs(8534) <= not(inputs(88)) or (inputs(11));
    layer0_outputs(8535) <= not((inputs(149)) xor (inputs(105)));
    layer0_outputs(8536) <= '0';
    layer0_outputs(8537) <= inputs(190);
    layer0_outputs(8538) <= (inputs(115)) and not (inputs(50));
    layer0_outputs(8539) <= not(inputs(10));
    layer0_outputs(8540) <= inputs(189);
    layer0_outputs(8541) <= '1';
    layer0_outputs(8542) <= (inputs(6)) and not (inputs(74));
    layer0_outputs(8543) <= inputs(231);
    layer0_outputs(8544) <= '1';
    layer0_outputs(8545) <= not(inputs(148)) or (inputs(15));
    layer0_outputs(8546) <= inputs(189);
    layer0_outputs(8547) <= inputs(17);
    layer0_outputs(8548) <= (inputs(158)) or (inputs(221));
    layer0_outputs(8549) <= (inputs(6)) and not (inputs(107));
    layer0_outputs(8550) <= (inputs(1)) and not (inputs(161));
    layer0_outputs(8551) <= '1';
    layer0_outputs(8552) <= not(inputs(200));
    layer0_outputs(8553) <= not((inputs(244)) and (inputs(125)));
    layer0_outputs(8554) <= not(inputs(166)) or (inputs(110));
    layer0_outputs(8555) <= not((inputs(226)) and (inputs(237)));
    layer0_outputs(8556) <= not(inputs(173)) or (inputs(66));
    layer0_outputs(8557) <= not(inputs(35)) or (inputs(204));
    layer0_outputs(8558) <= (inputs(26)) and (inputs(204));
    layer0_outputs(8559) <= not(inputs(180)) or (inputs(10));
    layer0_outputs(8560) <= not(inputs(121));
    layer0_outputs(8561) <= (inputs(108)) and (inputs(72));
    layer0_outputs(8562) <= (inputs(43)) or (inputs(206));
    layer0_outputs(8563) <= (inputs(214)) and (inputs(55));
    layer0_outputs(8564) <= not(inputs(79)) or (inputs(213));
    layer0_outputs(8565) <= not(inputs(104)) or (inputs(206));
    layer0_outputs(8566) <= (inputs(222)) or (inputs(255));
    layer0_outputs(8567) <= not(inputs(245));
    layer0_outputs(8568) <= not((inputs(161)) xor (inputs(118)));
    layer0_outputs(8569) <= not((inputs(243)) or (inputs(67)));
    layer0_outputs(8570) <= not((inputs(115)) or (inputs(185)));
    layer0_outputs(8571) <= not(inputs(33));
    layer0_outputs(8572) <= (inputs(121)) and not (inputs(39));
    layer0_outputs(8573) <= (inputs(184)) and not (inputs(152));
    layer0_outputs(8574) <= (inputs(139)) and not (inputs(221));
    layer0_outputs(8575) <= not(inputs(157)) or (inputs(177));
    layer0_outputs(8576) <= not(inputs(150)) or (inputs(20));
    layer0_outputs(8577) <= not((inputs(7)) and (inputs(172)));
    layer0_outputs(8578) <= inputs(90);
    layer0_outputs(8579) <= not(inputs(255));
    layer0_outputs(8580) <= not((inputs(250)) or (inputs(181)));
    layer0_outputs(8581) <= (inputs(145)) or (inputs(185));
    layer0_outputs(8582) <= not((inputs(101)) or (inputs(95)));
    layer0_outputs(8583) <= not(inputs(52));
    layer0_outputs(8584) <= not((inputs(226)) and (inputs(212)));
    layer0_outputs(8585) <= not(inputs(179));
    layer0_outputs(8586) <= inputs(138);
    layer0_outputs(8587) <= not(inputs(154));
    layer0_outputs(8588) <= (inputs(84)) or (inputs(93));
    layer0_outputs(8589) <= inputs(208);
    layer0_outputs(8590) <= (inputs(99)) and (inputs(254));
    layer0_outputs(8591) <= inputs(63);
    layer0_outputs(8592) <= (inputs(228)) or (inputs(81));
    layer0_outputs(8593) <= (inputs(146)) and not (inputs(134));
    layer0_outputs(8594) <= not((inputs(84)) xor (inputs(171)));
    layer0_outputs(8595) <= not((inputs(214)) xor (inputs(22)));
    layer0_outputs(8596) <= not(inputs(224));
    layer0_outputs(8597) <= not(inputs(146));
    layer0_outputs(8598) <= inputs(210);
    layer0_outputs(8599) <= not(inputs(56));
    layer0_outputs(8600) <= (inputs(239)) and not (inputs(211));
    layer0_outputs(8601) <= not(inputs(56));
    layer0_outputs(8602) <= not(inputs(127));
    layer0_outputs(8603) <= not((inputs(168)) xor (inputs(144)));
    layer0_outputs(8604) <= not(inputs(151));
    layer0_outputs(8605) <= not(inputs(41));
    layer0_outputs(8606) <= inputs(51);
    layer0_outputs(8607) <= not((inputs(39)) xor (inputs(37)));
    layer0_outputs(8608) <= inputs(150);
    layer0_outputs(8609) <= not(inputs(175)) or (inputs(220));
    layer0_outputs(8610) <= not((inputs(131)) and (inputs(64)));
    layer0_outputs(8611) <= not((inputs(250)) or (inputs(185)));
    layer0_outputs(8612) <= (inputs(114)) and not (inputs(248));
    layer0_outputs(8613) <= not(inputs(152)) or (inputs(162));
    layer0_outputs(8614) <= not((inputs(234)) xor (inputs(51)));
    layer0_outputs(8615) <= not(inputs(133)) or (inputs(162));
    layer0_outputs(8616) <= (inputs(85)) and not (inputs(195));
    layer0_outputs(8617) <= not((inputs(67)) and (inputs(223)));
    layer0_outputs(8618) <= not((inputs(135)) or (inputs(138)));
    layer0_outputs(8619) <= '1';
    layer0_outputs(8620) <= not(inputs(154)) or (inputs(25));
    layer0_outputs(8621) <= (inputs(113)) and (inputs(251));
    layer0_outputs(8622) <= (inputs(196)) or (inputs(195));
    layer0_outputs(8623) <= not(inputs(245)) or (inputs(248));
    layer0_outputs(8624) <= not((inputs(183)) or (inputs(24)));
    layer0_outputs(8625) <= '0';
    layer0_outputs(8626) <= inputs(228);
    layer0_outputs(8627) <= (inputs(166)) and not (inputs(237));
    layer0_outputs(8628) <= (inputs(233)) or (inputs(32));
    layer0_outputs(8629) <= not((inputs(165)) and (inputs(208)));
    layer0_outputs(8630) <= inputs(21);
    layer0_outputs(8631) <= not(inputs(152));
    layer0_outputs(8632) <= not((inputs(47)) xor (inputs(173)));
    layer0_outputs(8633) <= (inputs(236)) or (inputs(106));
    layer0_outputs(8634) <= not(inputs(58)) or (inputs(160));
    layer0_outputs(8635) <= not(inputs(34)) or (inputs(127));
    layer0_outputs(8636) <= (inputs(124)) and not (inputs(105));
    layer0_outputs(8637) <= inputs(77);
    layer0_outputs(8638) <= not(inputs(232));
    layer0_outputs(8639) <= (inputs(196)) and not (inputs(29));
    layer0_outputs(8640) <= (inputs(129)) xor (inputs(202));
    layer0_outputs(8641) <= not(inputs(101)) or (inputs(42));
    layer0_outputs(8642) <= inputs(171);
    layer0_outputs(8643) <= not(inputs(132));
    layer0_outputs(8644) <= not(inputs(10));
    layer0_outputs(8645) <= (inputs(52)) and not (inputs(17));
    layer0_outputs(8646) <= not((inputs(206)) or (inputs(12)));
    layer0_outputs(8647) <= (inputs(99)) xor (inputs(253));
    layer0_outputs(8648) <= inputs(35);
    layer0_outputs(8649) <= '0';
    layer0_outputs(8650) <= (inputs(53)) and not (inputs(110));
    layer0_outputs(8651) <= (inputs(140)) or (inputs(93));
    layer0_outputs(8652) <= not(inputs(123));
    layer0_outputs(8653) <= (inputs(49)) and not (inputs(14));
    layer0_outputs(8654) <= inputs(11);
    layer0_outputs(8655) <= inputs(93);
    layer0_outputs(8656) <= not((inputs(239)) or (inputs(37)));
    layer0_outputs(8657) <= not(inputs(167)) or (inputs(38));
    layer0_outputs(8658) <= not(inputs(223)) or (inputs(84));
    layer0_outputs(8659) <= (inputs(147)) and not (inputs(211));
    layer0_outputs(8660) <= not(inputs(148));
    layer0_outputs(8661) <= not((inputs(69)) and (inputs(61)));
    layer0_outputs(8662) <= not(inputs(50)) or (inputs(65));
    layer0_outputs(8663) <= not((inputs(248)) and (inputs(192)));
    layer0_outputs(8664) <= (inputs(155)) and not (inputs(166));
    layer0_outputs(8665) <= inputs(87);
    layer0_outputs(8666) <= (inputs(117)) and not (inputs(133));
    layer0_outputs(8667) <= (inputs(193)) and (inputs(34));
    layer0_outputs(8668) <= inputs(155);
    layer0_outputs(8669) <= not((inputs(225)) xor (inputs(43)));
    layer0_outputs(8670) <= not((inputs(77)) or (inputs(65)));
    layer0_outputs(8671) <= not((inputs(177)) xor (inputs(161)));
    layer0_outputs(8672) <= not(inputs(108));
    layer0_outputs(8673) <= not(inputs(147)) or (inputs(5));
    layer0_outputs(8674) <= not(inputs(131)) or (inputs(62));
    layer0_outputs(8675) <= not((inputs(136)) or (inputs(231)));
    layer0_outputs(8676) <= not((inputs(35)) or (inputs(42)));
    layer0_outputs(8677) <= (inputs(73)) and not (inputs(27));
    layer0_outputs(8678) <= inputs(248);
    layer0_outputs(8679) <= not(inputs(164)) or (inputs(95));
    layer0_outputs(8680) <= inputs(186);
    layer0_outputs(8681) <= '0';
    layer0_outputs(8682) <= not(inputs(245)) or (inputs(209));
    layer0_outputs(8683) <= not(inputs(226)) or (inputs(238));
    layer0_outputs(8684) <= (inputs(47)) or (inputs(2));
    layer0_outputs(8685) <= not((inputs(212)) xor (inputs(114)));
    layer0_outputs(8686) <= not((inputs(192)) and (inputs(146)));
    layer0_outputs(8687) <= not(inputs(5)) or (inputs(149));
    layer0_outputs(8688) <= '1';
    layer0_outputs(8689) <= (inputs(234)) and not (inputs(156));
    layer0_outputs(8690) <= '0';
    layer0_outputs(8691) <= not(inputs(182));
    layer0_outputs(8692) <= inputs(249);
    layer0_outputs(8693) <= (inputs(166)) and not (inputs(189));
    layer0_outputs(8694) <= not((inputs(80)) and (inputs(127)));
    layer0_outputs(8695) <= not(inputs(198));
    layer0_outputs(8696) <= '1';
    layer0_outputs(8697) <= '1';
    layer0_outputs(8698) <= not((inputs(232)) or (inputs(166)));
    layer0_outputs(8699) <= not((inputs(24)) and (inputs(217)));
    layer0_outputs(8700) <= inputs(9);
    layer0_outputs(8701) <= not((inputs(92)) and (inputs(96)));
    layer0_outputs(8702) <= (inputs(25)) xor (inputs(146));
    layer0_outputs(8703) <= (inputs(246)) and (inputs(6));
    layer0_outputs(8704) <= not((inputs(170)) xor (inputs(249)));
    layer0_outputs(8705) <= inputs(183);
    layer0_outputs(8706) <= inputs(128);
    layer0_outputs(8707) <= not((inputs(28)) xor (inputs(153)));
    layer0_outputs(8708) <= inputs(26);
    layer0_outputs(8709) <= not((inputs(244)) xor (inputs(243)));
    layer0_outputs(8710) <= not(inputs(9)) or (inputs(247));
    layer0_outputs(8711) <= (inputs(191)) and not (inputs(114));
    layer0_outputs(8712) <= not((inputs(176)) and (inputs(2)));
    layer0_outputs(8713) <= not(inputs(5));
    layer0_outputs(8714) <= (inputs(58)) or (inputs(111));
    layer0_outputs(8715) <= not(inputs(44)) or (inputs(75));
    layer0_outputs(8716) <= not(inputs(57)) or (inputs(61));
    layer0_outputs(8717) <= not((inputs(232)) and (inputs(175)));
    layer0_outputs(8718) <= '1';
    layer0_outputs(8719) <= (inputs(235)) xor (inputs(223));
    layer0_outputs(8720) <= (inputs(158)) or (inputs(167));
    layer0_outputs(8721) <= not((inputs(199)) xor (inputs(96)));
    layer0_outputs(8722) <= not((inputs(182)) xor (inputs(209)));
    layer0_outputs(8723) <= '1';
    layer0_outputs(8724) <= not((inputs(201)) xor (inputs(36)));
    layer0_outputs(8725) <= (inputs(200)) and not (inputs(48));
    layer0_outputs(8726) <= (inputs(112)) and not (inputs(40));
    layer0_outputs(8727) <= not((inputs(194)) or (inputs(130)));
    layer0_outputs(8728) <= not(inputs(110)) or (inputs(96));
    layer0_outputs(8729) <= '0';
    layer0_outputs(8730) <= (inputs(119)) xor (inputs(21));
    layer0_outputs(8731) <= not(inputs(104));
    layer0_outputs(8732) <= not((inputs(69)) or (inputs(23)));
    layer0_outputs(8733) <= inputs(117);
    layer0_outputs(8734) <= not(inputs(153)) or (inputs(197));
    layer0_outputs(8735) <= not(inputs(95)) or (inputs(48));
    layer0_outputs(8736) <= (inputs(226)) or (inputs(20));
    layer0_outputs(8737) <= not(inputs(59));
    layer0_outputs(8738) <= inputs(18);
    layer0_outputs(8739) <= not((inputs(117)) and (inputs(3)));
    layer0_outputs(8740) <= '0';
    layer0_outputs(8741) <= '0';
    layer0_outputs(8742) <= inputs(187);
    layer0_outputs(8743) <= (inputs(253)) or (inputs(125));
    layer0_outputs(8744) <= not(inputs(97)) or (inputs(233));
    layer0_outputs(8745) <= '0';
    layer0_outputs(8746) <= (inputs(34)) and (inputs(221));
    layer0_outputs(8747) <= not(inputs(135)) or (inputs(102));
    layer0_outputs(8748) <= not((inputs(6)) or (inputs(165)));
    layer0_outputs(8749) <= not((inputs(188)) or (inputs(151)));
    layer0_outputs(8750) <= inputs(199);
    layer0_outputs(8751) <= not(inputs(126));
    layer0_outputs(8752) <= not((inputs(111)) or (inputs(252)));
    layer0_outputs(8753) <= not(inputs(114)) or (inputs(60));
    layer0_outputs(8754) <= not((inputs(117)) and (inputs(58)));
    layer0_outputs(8755) <= (inputs(142)) xor (inputs(162));
    layer0_outputs(8756) <= not((inputs(224)) and (inputs(105)));
    layer0_outputs(8757) <= not(inputs(52)) or (inputs(15));
    layer0_outputs(8758) <= not(inputs(12));
    layer0_outputs(8759) <= not(inputs(91));
    layer0_outputs(8760) <= not(inputs(106));
    layer0_outputs(8761) <= (inputs(218)) and not (inputs(82));
    layer0_outputs(8762) <= not(inputs(125)) or (inputs(226));
    layer0_outputs(8763) <= (inputs(189)) and (inputs(66));
    layer0_outputs(8764) <= not(inputs(134)) or (inputs(22));
    layer0_outputs(8765) <= not((inputs(240)) or (inputs(172)));
    layer0_outputs(8766) <= (inputs(51)) and (inputs(37));
    layer0_outputs(8767) <= inputs(77);
    layer0_outputs(8768) <= not((inputs(199)) or (inputs(181)));
    layer0_outputs(8769) <= (inputs(91)) xor (inputs(112));
    layer0_outputs(8770) <= inputs(35);
    layer0_outputs(8771) <= not((inputs(225)) or (inputs(114)));
    layer0_outputs(8772) <= not((inputs(133)) or (inputs(93)));
    layer0_outputs(8773) <= not((inputs(66)) and (inputs(231)));
    layer0_outputs(8774) <= not((inputs(172)) or (inputs(220)));
    layer0_outputs(8775) <= not(inputs(148)) or (inputs(227));
    layer0_outputs(8776) <= inputs(253);
    layer0_outputs(8777) <= not((inputs(74)) and (inputs(188)));
    layer0_outputs(8778) <= inputs(153);
    layer0_outputs(8779) <= (inputs(34)) xor (inputs(44));
    layer0_outputs(8780) <= not(inputs(166));
    layer0_outputs(8781) <= (inputs(214)) and not (inputs(66));
    layer0_outputs(8782) <= not((inputs(27)) or (inputs(119)));
    layer0_outputs(8783) <= '1';
    layer0_outputs(8784) <= not((inputs(179)) or (inputs(155)));
    layer0_outputs(8785) <= not((inputs(58)) and (inputs(210)));
    layer0_outputs(8786) <= '0';
    layer0_outputs(8787) <= '0';
    layer0_outputs(8788) <= not(inputs(60));
    layer0_outputs(8789) <= inputs(95);
    layer0_outputs(8790) <= (inputs(239)) and (inputs(221));
    layer0_outputs(8791) <= (inputs(168)) and not (inputs(97));
    layer0_outputs(8792) <= not(inputs(7));
    layer0_outputs(8793) <= not(inputs(145)) or (inputs(25));
    layer0_outputs(8794) <= not(inputs(135));
    layer0_outputs(8795) <= not(inputs(162)) or (inputs(62));
    layer0_outputs(8796) <= '1';
    layer0_outputs(8797) <= (inputs(167)) xor (inputs(29));
    layer0_outputs(8798) <= inputs(209);
    layer0_outputs(8799) <= not(inputs(124)) or (inputs(110));
    layer0_outputs(8800) <= not((inputs(93)) or (inputs(116)));
    layer0_outputs(8801) <= not((inputs(146)) xor (inputs(159)));
    layer0_outputs(8802) <= not((inputs(125)) or (inputs(180)));
    layer0_outputs(8803) <= inputs(89);
    layer0_outputs(8804) <= (inputs(208)) or (inputs(59));
    layer0_outputs(8805) <= not((inputs(145)) xor (inputs(153)));
    layer0_outputs(8806) <= '0';
    layer0_outputs(8807) <= not((inputs(43)) xor (inputs(88)));
    layer0_outputs(8808) <= '0';
    layer0_outputs(8809) <= '1';
    layer0_outputs(8810) <= inputs(112);
    layer0_outputs(8811) <= not((inputs(29)) xor (inputs(243)));
    layer0_outputs(8812) <= not(inputs(125));
    layer0_outputs(8813) <= not((inputs(85)) or (inputs(174)));
    layer0_outputs(8814) <= not(inputs(29));
    layer0_outputs(8815) <= not(inputs(89));
    layer0_outputs(8816) <= (inputs(132)) or (inputs(211));
    layer0_outputs(8817) <= not(inputs(91)) or (inputs(46));
    layer0_outputs(8818) <= not((inputs(187)) xor (inputs(110)));
    layer0_outputs(8819) <= inputs(187);
    layer0_outputs(8820) <= inputs(163);
    layer0_outputs(8821) <= not((inputs(183)) and (inputs(146)));
    layer0_outputs(8822) <= not(inputs(130)) or (inputs(27));
    layer0_outputs(8823) <= (inputs(135)) and not (inputs(107));
    layer0_outputs(8824) <= inputs(3);
    layer0_outputs(8825) <= not(inputs(184)) or (inputs(186));
    layer0_outputs(8826) <= (inputs(112)) and not (inputs(193));
    layer0_outputs(8827) <= (inputs(141)) or (inputs(28));
    layer0_outputs(8828) <= inputs(129);
    layer0_outputs(8829) <= not((inputs(99)) xor (inputs(25)));
    layer0_outputs(8830) <= not(inputs(123));
    layer0_outputs(8831) <= (inputs(53)) and not (inputs(112));
    layer0_outputs(8832) <= not((inputs(183)) and (inputs(7)));
    layer0_outputs(8833) <= not((inputs(93)) or (inputs(213)));
    layer0_outputs(8834) <= not((inputs(75)) or (inputs(50)));
    layer0_outputs(8835) <= '0';
    layer0_outputs(8836) <= (inputs(180)) and not (inputs(97));
    layer0_outputs(8837) <= inputs(237);
    layer0_outputs(8838) <= (inputs(166)) and not (inputs(100));
    layer0_outputs(8839) <= not((inputs(47)) xor (inputs(172)));
    layer0_outputs(8840) <= not((inputs(82)) and (inputs(218)));
    layer0_outputs(8841) <= not((inputs(66)) and (inputs(0)));
    layer0_outputs(8842) <= not((inputs(101)) or (inputs(188)));
    layer0_outputs(8843) <= not(inputs(40));
    layer0_outputs(8844) <= not((inputs(160)) or (inputs(135)));
    layer0_outputs(8845) <= not((inputs(41)) or (inputs(96)));
    layer0_outputs(8846) <= inputs(9);
    layer0_outputs(8847) <= (inputs(136)) xor (inputs(45));
    layer0_outputs(8848) <= (inputs(220)) and not (inputs(197));
    layer0_outputs(8849) <= not((inputs(209)) and (inputs(18)));
    layer0_outputs(8850) <= '1';
    layer0_outputs(8851) <= (inputs(248)) or (inputs(86));
    layer0_outputs(8852) <= not(inputs(188));
    layer0_outputs(8853) <= (inputs(152)) and not (inputs(6));
    layer0_outputs(8854) <= (inputs(238)) or (inputs(225));
    layer0_outputs(8855) <= inputs(85);
    layer0_outputs(8856) <= inputs(137);
    layer0_outputs(8857) <= not((inputs(141)) or (inputs(12)));
    layer0_outputs(8858) <= not(inputs(91)) or (inputs(137));
    layer0_outputs(8859) <= not((inputs(3)) and (inputs(227)));
    layer0_outputs(8860) <= '1';
    layer0_outputs(8861) <= not((inputs(189)) or (inputs(172)));
    layer0_outputs(8862) <= inputs(159);
    layer0_outputs(8863) <= not(inputs(216)) or (inputs(42));
    layer0_outputs(8864) <= not(inputs(70)) or (inputs(215));
    layer0_outputs(8865) <= (inputs(194)) and (inputs(184));
    layer0_outputs(8866) <= '1';
    layer0_outputs(8867) <= (inputs(169)) xor (inputs(51));
    layer0_outputs(8868) <= (inputs(193)) and not (inputs(237));
    layer0_outputs(8869) <= not((inputs(107)) xor (inputs(177)));
    layer0_outputs(8870) <= (inputs(247)) and not (inputs(225));
    layer0_outputs(8871) <= (inputs(107)) and not (inputs(212));
    layer0_outputs(8872) <= '0';
    layer0_outputs(8873) <= (inputs(150)) and not (inputs(50));
    layer0_outputs(8874) <= inputs(14);
    layer0_outputs(8875) <= (inputs(166)) and (inputs(196));
    layer0_outputs(8876) <= (inputs(123)) and not (inputs(54));
    layer0_outputs(8877) <= not(inputs(164));
    layer0_outputs(8878) <= not(inputs(254));
    layer0_outputs(8879) <= not((inputs(170)) xor (inputs(82)));
    layer0_outputs(8880) <= not((inputs(225)) xor (inputs(72)));
    layer0_outputs(8881) <= not((inputs(69)) or (inputs(173)));
    layer0_outputs(8882) <= not(inputs(248)) or (inputs(27));
    layer0_outputs(8883) <= not(inputs(202));
    layer0_outputs(8884) <= (inputs(220)) and not (inputs(135));
    layer0_outputs(8885) <= inputs(151);
    layer0_outputs(8886) <= not(inputs(244));
    layer0_outputs(8887) <= not(inputs(92));
    layer0_outputs(8888) <= not((inputs(31)) or (inputs(183)));
    layer0_outputs(8889) <= (inputs(222)) or (inputs(53));
    layer0_outputs(8890) <= (inputs(168)) or (inputs(176));
    layer0_outputs(8891) <= '0';
    layer0_outputs(8892) <= (inputs(205)) and (inputs(111));
    layer0_outputs(8893) <= not((inputs(234)) or (inputs(13)));
    layer0_outputs(8894) <= not(inputs(13)) or (inputs(58));
    layer0_outputs(8895) <= (inputs(82)) and (inputs(9));
    layer0_outputs(8896) <= not(inputs(110)) or (inputs(173));
    layer0_outputs(8897) <= inputs(122);
    layer0_outputs(8898) <= not((inputs(16)) or (inputs(113)));
    layer0_outputs(8899) <= (inputs(12)) and not (inputs(163));
    layer0_outputs(8900) <= (inputs(195)) or (inputs(156));
    layer0_outputs(8901) <= not((inputs(155)) or (inputs(41)));
    layer0_outputs(8902) <= not(inputs(102)) or (inputs(232));
    layer0_outputs(8903) <= not((inputs(142)) or (inputs(97)));
    layer0_outputs(8904) <= (inputs(122)) or (inputs(147));
    layer0_outputs(8905) <= inputs(180);
    layer0_outputs(8906) <= (inputs(152)) xor (inputs(246));
    layer0_outputs(8907) <= not(inputs(172)) or (inputs(175));
    layer0_outputs(8908) <= (inputs(158)) and not (inputs(99));
    layer0_outputs(8909) <= not(inputs(195));
    layer0_outputs(8910) <= inputs(143);
    layer0_outputs(8911) <= not(inputs(243));
    layer0_outputs(8912) <= '0';
    layer0_outputs(8913) <= not(inputs(32));
    layer0_outputs(8914) <= not(inputs(250));
    layer0_outputs(8915) <= inputs(205);
    layer0_outputs(8916) <= (inputs(172)) and not (inputs(92));
    layer0_outputs(8917) <= not((inputs(58)) or (inputs(69)));
    layer0_outputs(8918) <= inputs(8);
    layer0_outputs(8919) <= (inputs(106)) or (inputs(10));
    layer0_outputs(8920) <= not(inputs(238)) or (inputs(187));
    layer0_outputs(8921) <= inputs(18);
    layer0_outputs(8922) <= (inputs(232)) and not (inputs(27));
    layer0_outputs(8923) <= (inputs(74)) or (inputs(8));
    layer0_outputs(8924) <= (inputs(203)) and (inputs(43));
    layer0_outputs(8925) <= not(inputs(76));
    layer0_outputs(8926) <= not((inputs(141)) or (inputs(90)));
    layer0_outputs(8927) <= not(inputs(24));
    layer0_outputs(8928) <= (inputs(103)) and not (inputs(79));
    layer0_outputs(8929) <= (inputs(207)) and (inputs(81));
    layer0_outputs(8930) <= '0';
    layer0_outputs(8931) <= not(inputs(70));
    layer0_outputs(8932) <= (inputs(128)) and not (inputs(234));
    layer0_outputs(8933) <= inputs(34);
    layer0_outputs(8934) <= not((inputs(115)) xor (inputs(238)));
    layer0_outputs(8935) <= not(inputs(180));
    layer0_outputs(8936) <= '1';
    layer0_outputs(8937) <= (inputs(198)) or (inputs(84));
    layer0_outputs(8938) <= not(inputs(90));
    layer0_outputs(8939) <= not(inputs(72));
    layer0_outputs(8940) <= not(inputs(171));
    layer0_outputs(8941) <= not(inputs(38)) or (inputs(93));
    layer0_outputs(8942) <= inputs(20);
    layer0_outputs(8943) <= (inputs(104)) and not (inputs(158));
    layer0_outputs(8944) <= not(inputs(33));
    layer0_outputs(8945) <= not(inputs(77)) or (inputs(40));
    layer0_outputs(8946) <= not(inputs(121));
    layer0_outputs(8947) <= not(inputs(22));
    layer0_outputs(8948) <= (inputs(185)) or (inputs(121));
    layer0_outputs(8949) <= (inputs(206)) or (inputs(77));
    layer0_outputs(8950) <= (inputs(20)) and not (inputs(131));
    layer0_outputs(8951) <= not((inputs(63)) xor (inputs(12)));
    layer0_outputs(8952) <= not(inputs(78)) or (inputs(26));
    layer0_outputs(8953) <= (inputs(198)) and (inputs(198));
    layer0_outputs(8954) <= not(inputs(100));
    layer0_outputs(8955) <= (inputs(244)) and (inputs(220));
    layer0_outputs(8956) <= not(inputs(104)) or (inputs(50));
    layer0_outputs(8957) <= (inputs(116)) and not (inputs(210));
    layer0_outputs(8958) <= inputs(228);
    layer0_outputs(8959) <= inputs(245);
    layer0_outputs(8960) <= inputs(228);
    layer0_outputs(8961) <= not(inputs(161)) or (inputs(200));
    layer0_outputs(8962) <= not((inputs(0)) xor (inputs(138)));
    layer0_outputs(8963) <= not((inputs(231)) or (inputs(8)));
    layer0_outputs(8964) <= (inputs(229)) and not (inputs(243));
    layer0_outputs(8965) <= (inputs(104)) and (inputs(1));
    layer0_outputs(8966) <= (inputs(229)) and (inputs(83));
    layer0_outputs(8967) <= not((inputs(216)) or (inputs(232)));
    layer0_outputs(8968) <= '1';
    layer0_outputs(8969) <= (inputs(186)) xor (inputs(200));
    layer0_outputs(8970) <= inputs(138);
    layer0_outputs(8971) <= '1';
    layer0_outputs(8972) <= not((inputs(1)) or (inputs(123)));
    layer0_outputs(8973) <= '0';
    layer0_outputs(8974) <= not((inputs(137)) and (inputs(14)));
    layer0_outputs(8975) <= (inputs(233)) and not (inputs(46));
    layer0_outputs(8976) <= (inputs(145)) and not (inputs(53));
    layer0_outputs(8977) <= not(inputs(191)) or (inputs(213));
    layer0_outputs(8978) <= not(inputs(49)) or (inputs(130));
    layer0_outputs(8979) <= not((inputs(142)) and (inputs(35)));
    layer0_outputs(8980) <= inputs(53);
    layer0_outputs(8981) <= '1';
    layer0_outputs(8982) <= not(inputs(132)) or (inputs(118));
    layer0_outputs(8983) <= (inputs(240)) and (inputs(210));
    layer0_outputs(8984) <= not((inputs(225)) or (inputs(199)));
    layer0_outputs(8985) <= inputs(228);
    layer0_outputs(8986) <= not(inputs(125)) or (inputs(57));
    layer0_outputs(8987) <= inputs(148);
    layer0_outputs(8988) <= not(inputs(13));
    layer0_outputs(8989) <= (inputs(198)) and not (inputs(5));
    layer0_outputs(8990) <= not((inputs(48)) or (inputs(127)));
    layer0_outputs(8991) <= (inputs(102)) or (inputs(124));
    layer0_outputs(8992) <= not((inputs(88)) or (inputs(104)));
    layer0_outputs(8993) <= not(inputs(247)) or (inputs(13));
    layer0_outputs(8994) <= inputs(144);
    layer0_outputs(8995) <= (inputs(100)) and not (inputs(17));
    layer0_outputs(8996) <= (inputs(19)) xor (inputs(172));
    layer0_outputs(8997) <= inputs(164);
    layer0_outputs(8998) <= (inputs(219)) and (inputs(153));
    layer0_outputs(8999) <= (inputs(194)) and not (inputs(31));
    layer0_outputs(9000) <= '0';
    layer0_outputs(9001) <= not(inputs(112)) or (inputs(179));
    layer0_outputs(9002) <= inputs(52);
    layer0_outputs(9003) <= (inputs(127)) or (inputs(157));
    layer0_outputs(9004) <= not((inputs(46)) or (inputs(78)));
    layer0_outputs(9005) <= '1';
    layer0_outputs(9006) <= not(inputs(191));
    layer0_outputs(9007) <= not((inputs(171)) or (inputs(19)));
    layer0_outputs(9008) <= not(inputs(104)) or (inputs(204));
    layer0_outputs(9009) <= '0';
    layer0_outputs(9010) <= (inputs(86)) or (inputs(133));
    layer0_outputs(9011) <= (inputs(122)) xor (inputs(113));
    layer0_outputs(9012) <= '1';
    layer0_outputs(9013) <= inputs(123);
    layer0_outputs(9014) <= (inputs(202)) and not (inputs(87));
    layer0_outputs(9015) <= not((inputs(138)) xor (inputs(21)));
    layer0_outputs(9016) <= (inputs(77)) and not (inputs(241));
    layer0_outputs(9017) <= not((inputs(255)) and (inputs(203)));
    layer0_outputs(9018) <= not((inputs(39)) or (inputs(220)));
    layer0_outputs(9019) <= '1';
    layer0_outputs(9020) <= (inputs(246)) and (inputs(22));
    layer0_outputs(9021) <= (inputs(38)) and not (inputs(131));
    layer0_outputs(9022) <= (inputs(197)) and not (inputs(199));
    layer0_outputs(9023) <= inputs(141);
    layer0_outputs(9024) <= inputs(249);
    layer0_outputs(9025) <= '1';
    layer0_outputs(9026) <= not(inputs(87));
    layer0_outputs(9027) <= not((inputs(241)) or (inputs(80)));
    layer0_outputs(9028) <= '0';
    layer0_outputs(9029) <= (inputs(63)) or (inputs(78));
    layer0_outputs(9030) <= '0';
    layer0_outputs(9031) <= not(inputs(170)) or (inputs(144));
    layer0_outputs(9032) <= (inputs(9)) and (inputs(5));
    layer0_outputs(9033) <= (inputs(202)) or (inputs(226));
    layer0_outputs(9034) <= not(inputs(86));
    layer0_outputs(9035) <= (inputs(73)) and (inputs(30));
    layer0_outputs(9036) <= not(inputs(181)) or (inputs(23));
    layer0_outputs(9037) <= not((inputs(86)) xor (inputs(19)));
    layer0_outputs(9038) <= not(inputs(84));
    layer0_outputs(9039) <= inputs(162);
    layer0_outputs(9040) <= inputs(189);
    layer0_outputs(9041) <= (inputs(158)) and not (inputs(45));
    layer0_outputs(9042) <= not((inputs(0)) or (inputs(161)));
    layer0_outputs(9043) <= not((inputs(43)) or (inputs(25)));
    layer0_outputs(9044) <= not(inputs(203));
    layer0_outputs(9045) <= inputs(106);
    layer0_outputs(9046) <= not((inputs(253)) or (inputs(212)));
    layer0_outputs(9047) <= not(inputs(169)) or (inputs(89));
    layer0_outputs(9048) <= not(inputs(202));
    layer0_outputs(9049) <= inputs(156);
    layer0_outputs(9050) <= not((inputs(7)) and (inputs(234)));
    layer0_outputs(9051) <= not(inputs(37));
    layer0_outputs(9052) <= (inputs(198)) and not (inputs(130));
    layer0_outputs(9053) <= not(inputs(192)) or (inputs(155));
    layer0_outputs(9054) <= (inputs(150)) xor (inputs(131));
    layer0_outputs(9055) <= not(inputs(20)) or (inputs(84));
    layer0_outputs(9056) <= inputs(36);
    layer0_outputs(9057) <= not((inputs(54)) or (inputs(183)));
    layer0_outputs(9058) <= not((inputs(24)) xor (inputs(208)));
    layer0_outputs(9059) <= (inputs(65)) and (inputs(43));
    layer0_outputs(9060) <= (inputs(237)) xor (inputs(86));
    layer0_outputs(9061) <= not(inputs(175));
    layer0_outputs(9062) <= not(inputs(27)) or (inputs(32));
    layer0_outputs(9063) <= not(inputs(126));
    layer0_outputs(9064) <= inputs(108);
    layer0_outputs(9065) <= not((inputs(161)) xor (inputs(94)));
    layer0_outputs(9066) <= '1';
    layer0_outputs(9067) <= (inputs(140)) or (inputs(159));
    layer0_outputs(9068) <= (inputs(54)) and not (inputs(10));
    layer0_outputs(9069) <= not(inputs(77));
    layer0_outputs(9070) <= (inputs(152)) or (inputs(205));
    layer0_outputs(9071) <= (inputs(210)) and not (inputs(157));
    layer0_outputs(9072) <= not(inputs(53)) or (inputs(94));
    layer0_outputs(9073) <= not(inputs(111));
    layer0_outputs(9074) <= (inputs(172)) and (inputs(239));
    layer0_outputs(9075) <= not(inputs(103)) or (inputs(201));
    layer0_outputs(9076) <= not((inputs(193)) xor (inputs(14)));
    layer0_outputs(9077) <= (inputs(45)) and not (inputs(16));
    layer0_outputs(9078) <= '0';
    layer0_outputs(9079) <= '0';
    layer0_outputs(9080) <= (inputs(6)) xor (inputs(247));
    layer0_outputs(9081) <= not(inputs(65)) or (inputs(46));
    layer0_outputs(9082) <= not(inputs(58)) or (inputs(238));
    layer0_outputs(9083) <= not((inputs(253)) or (inputs(220)));
    layer0_outputs(9084) <= '0';
    layer0_outputs(9085) <= inputs(23);
    layer0_outputs(9086) <= '1';
    layer0_outputs(9087) <= not((inputs(14)) or (inputs(30)));
    layer0_outputs(9088) <= not(inputs(230));
    layer0_outputs(9089) <= not(inputs(77)) or (inputs(11));
    layer0_outputs(9090) <= not((inputs(235)) xor (inputs(150)));
    layer0_outputs(9091) <= not((inputs(178)) xor (inputs(74)));
    layer0_outputs(9092) <= '1';
    layer0_outputs(9093) <= inputs(48);
    layer0_outputs(9094) <= not((inputs(132)) xor (inputs(150)));
    layer0_outputs(9095) <= (inputs(58)) xor (inputs(248));
    layer0_outputs(9096) <= not(inputs(213));
    layer0_outputs(9097) <= inputs(13);
    layer0_outputs(9098) <= inputs(83);
    layer0_outputs(9099) <= '0';
    layer0_outputs(9100) <= not(inputs(195)) or (inputs(96));
    layer0_outputs(9101) <= not(inputs(110)) or (inputs(6));
    layer0_outputs(9102) <= (inputs(169)) or (inputs(3));
    layer0_outputs(9103) <= (inputs(110)) and not (inputs(78));
    layer0_outputs(9104) <= inputs(58);
    layer0_outputs(9105) <= (inputs(66)) or (inputs(68));
    layer0_outputs(9106) <= inputs(226);
    layer0_outputs(9107) <= not((inputs(166)) xor (inputs(160)));
    layer0_outputs(9108) <= '0';
    layer0_outputs(9109) <= (inputs(159)) or (inputs(128));
    layer0_outputs(9110) <= (inputs(235)) and not (inputs(24));
    layer0_outputs(9111) <= '1';
    layer0_outputs(9112) <= not(inputs(98));
    layer0_outputs(9113) <= (inputs(14)) xor (inputs(164));
    layer0_outputs(9114) <= (inputs(240)) and not (inputs(65));
    layer0_outputs(9115) <= inputs(161);
    layer0_outputs(9116) <= not(inputs(45));
    layer0_outputs(9117) <= (inputs(27)) or (inputs(118));
    layer0_outputs(9118) <= (inputs(153)) and not (inputs(40));
    layer0_outputs(9119) <= not((inputs(204)) or (inputs(238)));
    layer0_outputs(9120) <= '0';
    layer0_outputs(9121) <= not((inputs(236)) or (inputs(1)));
    layer0_outputs(9122) <= inputs(101);
    layer0_outputs(9123) <= '0';
    layer0_outputs(9124) <= not(inputs(135)) or (inputs(130));
    layer0_outputs(9125) <= (inputs(178)) xor (inputs(218));
    layer0_outputs(9126) <= not(inputs(231)) or (inputs(2));
    layer0_outputs(9127) <= inputs(158);
    layer0_outputs(9128) <= not((inputs(116)) and (inputs(214)));
    layer0_outputs(9129) <= '0';
    layer0_outputs(9130) <= not((inputs(19)) xor (inputs(246)));
    layer0_outputs(9131) <= not(inputs(5)) or (inputs(248));
    layer0_outputs(9132) <= inputs(179);
    layer0_outputs(9133) <= (inputs(192)) and not (inputs(58));
    layer0_outputs(9134) <= (inputs(174)) or (inputs(17));
    layer0_outputs(9135) <= not((inputs(95)) xor (inputs(61)));
    layer0_outputs(9136) <= inputs(140);
    layer0_outputs(9137) <= not(inputs(211)) or (inputs(183));
    layer0_outputs(9138) <= (inputs(217)) and (inputs(79));
    layer0_outputs(9139) <= (inputs(65)) xor (inputs(111));
    layer0_outputs(9140) <= (inputs(16)) and (inputs(161));
    layer0_outputs(9141) <= not(inputs(206));
    layer0_outputs(9142) <= (inputs(35)) and not (inputs(206));
    layer0_outputs(9143) <= (inputs(151)) xor (inputs(202));
    layer0_outputs(9144) <= not(inputs(245));
    layer0_outputs(9145) <= inputs(181);
    layer0_outputs(9146) <= not((inputs(14)) xor (inputs(189)));
    layer0_outputs(9147) <= (inputs(118)) or (inputs(138));
    layer0_outputs(9148) <= not((inputs(196)) or (inputs(63)));
    layer0_outputs(9149) <= not(inputs(33)) or (inputs(3));
    layer0_outputs(9150) <= not(inputs(88)) or (inputs(220));
    layer0_outputs(9151) <= (inputs(23)) or (inputs(141));
    layer0_outputs(9152) <= not((inputs(86)) or (inputs(60)));
    layer0_outputs(9153) <= (inputs(166)) and not (inputs(1));
    layer0_outputs(9154) <= (inputs(181)) and not (inputs(144));
    layer0_outputs(9155) <= (inputs(250)) and not (inputs(44));
    layer0_outputs(9156) <= not(inputs(205)) or (inputs(207));
    layer0_outputs(9157) <= inputs(153);
    layer0_outputs(9158) <= not(inputs(135)) or (inputs(41));
    layer0_outputs(9159) <= (inputs(173)) or (inputs(244));
    layer0_outputs(9160) <= (inputs(29)) xor (inputs(137));
    layer0_outputs(9161) <= not((inputs(13)) or (inputs(239)));
    layer0_outputs(9162) <= not(inputs(226));
    layer0_outputs(9163) <= inputs(150);
    layer0_outputs(9164) <= not((inputs(30)) and (inputs(138)));
    layer0_outputs(9165) <= '1';
    layer0_outputs(9166) <= inputs(251);
    layer0_outputs(9167) <= (inputs(226)) or (inputs(117));
    layer0_outputs(9168) <= not(inputs(153)) or (inputs(19));
    layer0_outputs(9169) <= (inputs(242)) xor (inputs(185));
    layer0_outputs(9170) <= (inputs(52)) or (inputs(210));
    layer0_outputs(9171) <= not((inputs(223)) or (inputs(155)));
    layer0_outputs(9172) <= (inputs(187)) xor (inputs(109));
    layer0_outputs(9173) <= not(inputs(3));
    layer0_outputs(9174) <= not((inputs(251)) and (inputs(104)));
    layer0_outputs(9175) <= inputs(9);
    layer0_outputs(9176) <= inputs(211);
    layer0_outputs(9177) <= not((inputs(145)) xor (inputs(210)));
    layer0_outputs(9178) <= not((inputs(209)) and (inputs(246)));
    layer0_outputs(9179) <= (inputs(180)) and not (inputs(176));
    layer0_outputs(9180) <= (inputs(74)) and not (inputs(144));
    layer0_outputs(9181) <= (inputs(120)) or (inputs(26));
    layer0_outputs(9182) <= (inputs(13)) or (inputs(102));
    layer0_outputs(9183) <= not(inputs(131)) or (inputs(94));
    layer0_outputs(9184) <= (inputs(212)) xor (inputs(102));
    layer0_outputs(9185) <= not((inputs(14)) xor (inputs(129)));
    layer0_outputs(9186) <= (inputs(101)) and not (inputs(4));
    layer0_outputs(9187) <= not(inputs(204));
    layer0_outputs(9188) <= not((inputs(151)) or (inputs(111)));
    layer0_outputs(9189) <= (inputs(182)) and (inputs(246));
    layer0_outputs(9190) <= not((inputs(225)) and (inputs(191)));
    layer0_outputs(9191) <= not(inputs(107)) or (inputs(58));
    layer0_outputs(9192) <= not((inputs(250)) and (inputs(85)));
    layer0_outputs(9193) <= not((inputs(88)) or (inputs(93)));
    layer0_outputs(9194) <= inputs(45);
    layer0_outputs(9195) <= (inputs(103)) and not (inputs(130));
    layer0_outputs(9196) <= not((inputs(7)) or (inputs(151)));
    layer0_outputs(9197) <= (inputs(0)) and not (inputs(122));
    layer0_outputs(9198) <= inputs(78);
    layer0_outputs(9199) <= not(inputs(196));
    layer0_outputs(9200) <= not((inputs(253)) xor (inputs(248)));
    layer0_outputs(9201) <= (inputs(237)) and not (inputs(68));
    layer0_outputs(9202) <= not(inputs(5));
    layer0_outputs(9203) <= '0';
    layer0_outputs(9204) <= not((inputs(45)) or (inputs(209)));
    layer0_outputs(9205) <= not(inputs(150));
    layer0_outputs(9206) <= inputs(126);
    layer0_outputs(9207) <= '0';
    layer0_outputs(9208) <= not(inputs(89)) or (inputs(9));
    layer0_outputs(9209) <= not(inputs(97)) or (inputs(231));
    layer0_outputs(9210) <= inputs(150);
    layer0_outputs(9211) <= not(inputs(136)) or (inputs(78));
    layer0_outputs(9212) <= inputs(235);
    layer0_outputs(9213) <= not(inputs(172));
    layer0_outputs(9214) <= (inputs(122)) and (inputs(81));
    layer0_outputs(9215) <= not(inputs(112)) or (inputs(54));
    layer0_outputs(9216) <= '0';
    layer0_outputs(9217) <= not((inputs(123)) or (inputs(73)));
    layer0_outputs(9218) <= (inputs(190)) xor (inputs(147));
    layer0_outputs(9219) <= (inputs(17)) or (inputs(195));
    layer0_outputs(9220) <= inputs(132);
    layer0_outputs(9221) <= (inputs(147)) and not (inputs(52));
    layer0_outputs(9222) <= not((inputs(153)) xor (inputs(155)));
    layer0_outputs(9223) <= inputs(122);
    layer0_outputs(9224) <= not(inputs(136)) or (inputs(133));
    layer0_outputs(9225) <= not((inputs(127)) xor (inputs(149)));
    layer0_outputs(9226) <= not(inputs(120)) or (inputs(51));
    layer0_outputs(9227) <= '0';
    layer0_outputs(9228) <= '0';
    layer0_outputs(9229) <= not((inputs(117)) or (inputs(33)));
    layer0_outputs(9230) <= inputs(222);
    layer0_outputs(9231) <= not((inputs(98)) xor (inputs(33)));
    layer0_outputs(9232) <= not(inputs(119));
    layer0_outputs(9233) <= '1';
    layer0_outputs(9234) <= inputs(81);
    layer0_outputs(9235) <= (inputs(170)) xor (inputs(99));
    layer0_outputs(9236) <= not((inputs(159)) xor (inputs(4)));
    layer0_outputs(9237) <= not(inputs(227));
    layer0_outputs(9238) <= not((inputs(253)) xor (inputs(204)));
    layer0_outputs(9239) <= not(inputs(11)) or (inputs(86));
    layer0_outputs(9240) <= not(inputs(41)) or (inputs(40));
    layer0_outputs(9241) <= inputs(35);
    layer0_outputs(9242) <= (inputs(21)) or (inputs(216));
    layer0_outputs(9243) <= inputs(126);
    layer0_outputs(9244) <= (inputs(75)) or (inputs(98));
    layer0_outputs(9245) <= not((inputs(222)) or (inputs(79)));
    layer0_outputs(9246) <= (inputs(115)) or (inputs(78));
    layer0_outputs(9247) <= (inputs(45)) and not (inputs(136));
    layer0_outputs(9248) <= not((inputs(93)) and (inputs(131)));
    layer0_outputs(9249) <= not(inputs(195));
    layer0_outputs(9250) <= (inputs(160)) or (inputs(88));
    layer0_outputs(9251) <= not(inputs(91));
    layer0_outputs(9252) <= not((inputs(27)) or (inputs(165)));
    layer0_outputs(9253) <= not(inputs(109)) or (inputs(195));
    layer0_outputs(9254) <= not(inputs(224)) or (inputs(120));
    layer0_outputs(9255) <= (inputs(113)) and not (inputs(120));
    layer0_outputs(9256) <= (inputs(145)) xor (inputs(182));
    layer0_outputs(9257) <= not((inputs(148)) or (inputs(6)));
    layer0_outputs(9258) <= not(inputs(34)) or (inputs(174));
    layer0_outputs(9259) <= not(inputs(84)) or (inputs(6));
    layer0_outputs(9260) <= '0';
    layer0_outputs(9261) <= (inputs(61)) and not (inputs(183));
    layer0_outputs(9262) <= not((inputs(33)) or (inputs(7)));
    layer0_outputs(9263) <= (inputs(13)) xor (inputs(187));
    layer0_outputs(9264) <= not(inputs(141));
    layer0_outputs(9265) <= not(inputs(92)) or (inputs(154));
    layer0_outputs(9266) <= not(inputs(183)) or (inputs(230));
    layer0_outputs(9267) <= not(inputs(168)) or (inputs(57));
    layer0_outputs(9268) <= not((inputs(75)) or (inputs(196)));
    layer0_outputs(9269) <= '1';
    layer0_outputs(9270) <= (inputs(39)) or (inputs(142));
    layer0_outputs(9271) <= inputs(227);
    layer0_outputs(9272) <= inputs(112);
    layer0_outputs(9273) <= not((inputs(229)) or (inputs(201)));
    layer0_outputs(9274) <= (inputs(123)) xor (inputs(253));
    layer0_outputs(9275) <= not(inputs(100));
    layer0_outputs(9276) <= not(inputs(113)) or (inputs(1));
    layer0_outputs(9277) <= inputs(166);
    layer0_outputs(9278) <= not((inputs(95)) or (inputs(127)));
    layer0_outputs(9279) <= not((inputs(155)) xor (inputs(95)));
    layer0_outputs(9280) <= '0';
    layer0_outputs(9281) <= (inputs(113)) xor (inputs(28));
    layer0_outputs(9282) <= (inputs(110)) and not (inputs(30));
    layer0_outputs(9283) <= (inputs(39)) xor (inputs(198));
    layer0_outputs(9284) <= '0';
    layer0_outputs(9285) <= not(inputs(117)) or (inputs(199));
    layer0_outputs(9286) <= (inputs(22)) or (inputs(157));
    layer0_outputs(9287) <= not(inputs(123)) or (inputs(194));
    layer0_outputs(9288) <= not(inputs(242));
    layer0_outputs(9289) <= (inputs(152)) or (inputs(203));
    layer0_outputs(9290) <= '0';
    layer0_outputs(9291) <= inputs(193);
    layer0_outputs(9292) <= '0';
    layer0_outputs(9293) <= not(inputs(43)) or (inputs(113));
    layer0_outputs(9294) <= inputs(38);
    layer0_outputs(9295) <= (inputs(50)) and not (inputs(205));
    layer0_outputs(9296) <= not(inputs(91)) or (inputs(222));
    layer0_outputs(9297) <= not((inputs(146)) or (inputs(15)));
    layer0_outputs(9298) <= not(inputs(111)) or (inputs(65));
    layer0_outputs(9299) <= (inputs(174)) and (inputs(51));
    layer0_outputs(9300) <= (inputs(216)) or (inputs(15));
    layer0_outputs(9301) <= not((inputs(48)) xor (inputs(125)));
    layer0_outputs(9302) <= inputs(151);
    layer0_outputs(9303) <= (inputs(17)) and not (inputs(226));
    layer0_outputs(9304) <= not(inputs(151));
    layer0_outputs(9305) <= not((inputs(4)) xor (inputs(152)));
    layer0_outputs(9306) <= not(inputs(74)) or (inputs(122));
    layer0_outputs(9307) <= not((inputs(72)) and (inputs(128)));
    layer0_outputs(9308) <= not((inputs(148)) xor (inputs(223)));
    layer0_outputs(9309) <= not((inputs(231)) xor (inputs(229)));
    layer0_outputs(9310) <= inputs(223);
    layer0_outputs(9311) <= inputs(2);
    layer0_outputs(9312) <= not((inputs(61)) and (inputs(247)));
    layer0_outputs(9313) <= (inputs(55)) and not (inputs(82));
    layer0_outputs(9314) <= not((inputs(158)) xor (inputs(34)));
    layer0_outputs(9315) <= inputs(187);
    layer0_outputs(9316) <= inputs(249);
    layer0_outputs(9317) <= not((inputs(31)) xor (inputs(166)));
    layer0_outputs(9318) <= (inputs(112)) and (inputs(208));
    layer0_outputs(9319) <= '0';
    layer0_outputs(9320) <= not(inputs(213));
    layer0_outputs(9321) <= not(inputs(137));
    layer0_outputs(9322) <= (inputs(2)) or (inputs(187));
    layer0_outputs(9323) <= inputs(247);
    layer0_outputs(9324) <= (inputs(227)) and not (inputs(126));
    layer0_outputs(9325) <= not(inputs(251)) or (inputs(192));
    layer0_outputs(9326) <= not((inputs(229)) or (inputs(64)));
    layer0_outputs(9327) <= (inputs(24)) and not (inputs(2));
    layer0_outputs(9328) <= not((inputs(93)) xor (inputs(107)));
    layer0_outputs(9329) <= '0';
    layer0_outputs(9330) <= (inputs(68)) and not (inputs(234));
    layer0_outputs(9331) <= not(inputs(162)) or (inputs(140));
    layer0_outputs(9332) <= not((inputs(184)) xor (inputs(80)));
    layer0_outputs(9333) <= not((inputs(158)) xor (inputs(141)));
    layer0_outputs(9334) <= not(inputs(148)) or (inputs(110));
    layer0_outputs(9335) <= inputs(151);
    layer0_outputs(9336) <= not((inputs(166)) or (inputs(29)));
    layer0_outputs(9337) <= (inputs(254)) and (inputs(46));
    layer0_outputs(9338) <= not((inputs(30)) and (inputs(174)));
    layer0_outputs(9339) <= inputs(103);
    layer0_outputs(9340) <= not(inputs(74)) or (inputs(45));
    layer0_outputs(9341) <= (inputs(63)) xor (inputs(165));
    layer0_outputs(9342) <= (inputs(86)) and not (inputs(226));
    layer0_outputs(9343) <= not(inputs(239));
    layer0_outputs(9344) <= '0';
    layer0_outputs(9345) <= (inputs(93)) and (inputs(199));
    layer0_outputs(9346) <= not(inputs(238));
    layer0_outputs(9347) <= not((inputs(66)) or (inputs(125)));
    layer0_outputs(9348) <= inputs(228);
    layer0_outputs(9349) <= (inputs(192)) and not (inputs(0));
    layer0_outputs(9350) <= inputs(250);
    layer0_outputs(9351) <= inputs(149);
    layer0_outputs(9352) <= inputs(199);
    layer0_outputs(9353) <= not(inputs(111)) or (inputs(118));
    layer0_outputs(9354) <= inputs(56);
    layer0_outputs(9355) <= not(inputs(220));
    layer0_outputs(9356) <= not(inputs(64)) or (inputs(114));
    layer0_outputs(9357) <= (inputs(242)) xor (inputs(12));
    layer0_outputs(9358) <= not(inputs(32)) or (inputs(208));
    layer0_outputs(9359) <= '0';
    layer0_outputs(9360) <= (inputs(123)) and not (inputs(95));
    layer0_outputs(9361) <= inputs(140);
    layer0_outputs(9362) <= not(inputs(12)) or (inputs(14));
    layer0_outputs(9363) <= not(inputs(57));
    layer0_outputs(9364) <= (inputs(194)) xor (inputs(22));
    layer0_outputs(9365) <= (inputs(164)) or (inputs(60));
    layer0_outputs(9366) <= (inputs(120)) xor (inputs(209));
    layer0_outputs(9367) <= (inputs(221)) or (inputs(67));
    layer0_outputs(9368) <= not(inputs(122)) or (inputs(190));
    layer0_outputs(9369) <= not((inputs(152)) or (inputs(96)));
    layer0_outputs(9370) <= not(inputs(253)) or (inputs(18));
    layer0_outputs(9371) <= (inputs(72)) and (inputs(177));
    layer0_outputs(9372) <= (inputs(0)) and (inputs(141));
    layer0_outputs(9373) <= not(inputs(157)) or (inputs(146));
    layer0_outputs(9374) <= (inputs(38)) xor (inputs(11));
    layer0_outputs(9375) <= (inputs(234)) xor (inputs(104));
    layer0_outputs(9376) <= (inputs(229)) and not (inputs(128));
    layer0_outputs(9377) <= not(inputs(98)) or (inputs(85));
    layer0_outputs(9378) <= not(inputs(70)) or (inputs(169));
    layer0_outputs(9379) <= not((inputs(235)) xor (inputs(222)));
    layer0_outputs(9380) <= '1';
    layer0_outputs(9381) <= (inputs(119)) and not (inputs(174));
    layer0_outputs(9382) <= not((inputs(121)) or (inputs(170)));
    layer0_outputs(9383) <= (inputs(36)) or (inputs(181));
    layer0_outputs(9384) <= not(inputs(167)) or (inputs(125));
    layer0_outputs(9385) <= not((inputs(13)) or (inputs(122)));
    layer0_outputs(9386) <= not(inputs(56)) or (inputs(228));
    layer0_outputs(9387) <= (inputs(228)) and not (inputs(159));
    layer0_outputs(9388) <= not(inputs(207)) or (inputs(181));
    layer0_outputs(9389) <= inputs(178);
    layer0_outputs(9390) <= '1';
    layer0_outputs(9391) <= not((inputs(162)) xor (inputs(126)));
    layer0_outputs(9392) <= not(inputs(89));
    layer0_outputs(9393) <= not((inputs(193)) or (inputs(161)));
    layer0_outputs(9394) <= '1';
    layer0_outputs(9395) <= (inputs(163)) and not (inputs(129));
    layer0_outputs(9396) <= not(inputs(106));
    layer0_outputs(9397) <= not((inputs(49)) xor (inputs(169)));
    layer0_outputs(9398) <= not(inputs(7));
    layer0_outputs(9399) <= (inputs(92)) or (inputs(34));
    layer0_outputs(9400) <= (inputs(24)) xor (inputs(177));
    layer0_outputs(9401) <= (inputs(56)) xor (inputs(47));
    layer0_outputs(9402) <= not(inputs(107)) or (inputs(79));
    layer0_outputs(9403) <= not(inputs(199));
    layer0_outputs(9404) <= inputs(247);
    layer0_outputs(9405) <= '0';
    layer0_outputs(9406) <= (inputs(234)) and not (inputs(14));
    layer0_outputs(9407) <= (inputs(167)) xor (inputs(111));
    layer0_outputs(9408) <= '1';
    layer0_outputs(9409) <= not(inputs(100));
    layer0_outputs(9410) <= '0';
    layer0_outputs(9411) <= (inputs(19)) or (inputs(178));
    layer0_outputs(9412) <= not((inputs(232)) or (inputs(87)));
    layer0_outputs(9413) <= not(inputs(218));
    layer0_outputs(9414) <= not(inputs(74)) or (inputs(216));
    layer0_outputs(9415) <= (inputs(116)) xor (inputs(10));
    layer0_outputs(9416) <= (inputs(89)) and not (inputs(123));
    layer0_outputs(9417) <= inputs(86);
    layer0_outputs(9418) <= not((inputs(101)) or (inputs(236)));
    layer0_outputs(9419) <= (inputs(165)) and not (inputs(177));
    layer0_outputs(9420) <= not((inputs(165)) or (inputs(25)));
    layer0_outputs(9421) <= (inputs(120)) and (inputs(241));
    layer0_outputs(9422) <= (inputs(101)) xor (inputs(141));
    layer0_outputs(9423) <= not((inputs(26)) and (inputs(242)));
    layer0_outputs(9424) <= '1';
    layer0_outputs(9425) <= inputs(132);
    layer0_outputs(9426) <= (inputs(96)) and not (inputs(199));
    layer0_outputs(9427) <= not((inputs(62)) or (inputs(123)));
    layer0_outputs(9428) <= not(inputs(95)) or (inputs(216));
    layer0_outputs(9429) <= not(inputs(61));
    layer0_outputs(9430) <= inputs(216);
    layer0_outputs(9431) <= (inputs(54)) and not (inputs(66));
    layer0_outputs(9432) <= not((inputs(226)) or (inputs(5)));
    layer0_outputs(9433) <= '0';
    layer0_outputs(9434) <= inputs(128);
    layer0_outputs(9435) <= inputs(204);
    layer0_outputs(9436) <= not(inputs(142));
    layer0_outputs(9437) <= not((inputs(36)) or (inputs(164)));
    layer0_outputs(9438) <= not((inputs(26)) xor (inputs(133)));
    layer0_outputs(9439) <= not((inputs(182)) xor (inputs(224)));
    layer0_outputs(9440) <= not((inputs(96)) or (inputs(4)));
    layer0_outputs(9441) <= not(inputs(201)) or (inputs(76));
    layer0_outputs(9442) <= not((inputs(254)) xor (inputs(191)));
    layer0_outputs(9443) <= (inputs(31)) or (inputs(37));
    layer0_outputs(9444) <= (inputs(37)) or (inputs(243));
    layer0_outputs(9445) <= '0';
    layer0_outputs(9446) <= (inputs(37)) and not (inputs(27));
    layer0_outputs(9447) <= not(inputs(13));
    layer0_outputs(9448) <= not((inputs(55)) and (inputs(129)));
    layer0_outputs(9449) <= (inputs(194)) and (inputs(19));
    layer0_outputs(9450) <= not((inputs(92)) xor (inputs(89)));
    layer0_outputs(9451) <= (inputs(211)) and not (inputs(158));
    layer0_outputs(9452) <= inputs(6);
    layer0_outputs(9453) <= (inputs(197)) or (inputs(203));
    layer0_outputs(9454) <= not((inputs(165)) or (inputs(184)));
    layer0_outputs(9455) <= not(inputs(170)) or (inputs(210));
    layer0_outputs(9456) <= not((inputs(15)) xor (inputs(166)));
    layer0_outputs(9457) <= (inputs(2)) or (inputs(96));
    layer0_outputs(9458) <= (inputs(23)) xor (inputs(42));
    layer0_outputs(9459) <= inputs(250);
    layer0_outputs(9460) <= not((inputs(82)) or (inputs(193)));
    layer0_outputs(9461) <= (inputs(182)) xor (inputs(243));
    layer0_outputs(9462) <= inputs(67);
    layer0_outputs(9463) <= not(inputs(186)) or (inputs(121));
    layer0_outputs(9464) <= inputs(196);
    layer0_outputs(9465) <= not(inputs(154));
    layer0_outputs(9466) <= not(inputs(85));
    layer0_outputs(9467) <= (inputs(250)) or (inputs(100));
    layer0_outputs(9468) <= not(inputs(176));
    layer0_outputs(9469) <= '0';
    layer0_outputs(9470) <= (inputs(255)) xor (inputs(62));
    layer0_outputs(9471) <= not((inputs(230)) and (inputs(18)));
    layer0_outputs(9472) <= not((inputs(55)) and (inputs(44)));
    layer0_outputs(9473) <= not(inputs(136));
    layer0_outputs(9474) <= not(inputs(76));
    layer0_outputs(9475) <= not(inputs(106)) or (inputs(226));
    layer0_outputs(9476) <= (inputs(66)) and not (inputs(125));
    layer0_outputs(9477) <= not(inputs(101));
    layer0_outputs(9478) <= not(inputs(120));
    layer0_outputs(9479) <= '0';
    layer0_outputs(9480) <= not((inputs(21)) xor (inputs(2)));
    layer0_outputs(9481) <= not(inputs(130)) or (inputs(254));
    layer0_outputs(9482) <= not(inputs(182));
    layer0_outputs(9483) <= not((inputs(7)) and (inputs(255)));
    layer0_outputs(9484) <= not((inputs(232)) or (inputs(101)));
    layer0_outputs(9485) <= not((inputs(196)) or (inputs(186)));
    layer0_outputs(9486) <= (inputs(55)) and not (inputs(252));
    layer0_outputs(9487) <= not((inputs(87)) xor (inputs(169)));
    layer0_outputs(9488) <= (inputs(169)) and not (inputs(197));
    layer0_outputs(9489) <= not(inputs(114)) or (inputs(197));
    layer0_outputs(9490) <= (inputs(48)) xor (inputs(74));
    layer0_outputs(9491) <= (inputs(183)) and not (inputs(164));
    layer0_outputs(9492) <= '0';
    layer0_outputs(9493) <= '0';
    layer0_outputs(9494) <= (inputs(149)) xor (inputs(109));
    layer0_outputs(9495) <= '0';
    layer0_outputs(9496) <= (inputs(171)) and (inputs(189));
    layer0_outputs(9497) <= not((inputs(148)) xor (inputs(9)));
    layer0_outputs(9498) <= not((inputs(190)) or (inputs(72)));
    layer0_outputs(9499) <= not((inputs(235)) xor (inputs(147)));
    layer0_outputs(9500) <= not(inputs(58));
    layer0_outputs(9501) <= (inputs(157)) and not (inputs(90));
    layer0_outputs(9502) <= not((inputs(91)) xor (inputs(4)));
    layer0_outputs(9503) <= inputs(244);
    layer0_outputs(9504) <= inputs(189);
    layer0_outputs(9505) <= (inputs(55)) and not (inputs(95));
    layer0_outputs(9506) <= not(inputs(55)) or (inputs(91));
    layer0_outputs(9507) <= '1';
    layer0_outputs(9508) <= inputs(169);
    layer0_outputs(9509) <= '1';
    layer0_outputs(9510) <= not((inputs(235)) or (inputs(169)));
    layer0_outputs(9511) <= not((inputs(164)) xor (inputs(79)));
    layer0_outputs(9512) <= not((inputs(6)) xor (inputs(25)));
    layer0_outputs(9513) <= (inputs(218)) xor (inputs(234));
    layer0_outputs(9514) <= not((inputs(35)) and (inputs(48)));
    layer0_outputs(9515) <= '1';
    layer0_outputs(9516) <= inputs(25);
    layer0_outputs(9517) <= not(inputs(3));
    layer0_outputs(9518) <= '0';
    layer0_outputs(9519) <= (inputs(116)) or (inputs(48));
    layer0_outputs(9520) <= not(inputs(253)) or (inputs(13));
    layer0_outputs(9521) <= not(inputs(149)) or (inputs(228));
    layer0_outputs(9522) <= not(inputs(99)) or (inputs(14));
    layer0_outputs(9523) <= inputs(68);
    layer0_outputs(9524) <= (inputs(10)) and (inputs(12));
    layer0_outputs(9525) <= (inputs(8)) and (inputs(201));
    layer0_outputs(9526) <= not(inputs(168)) or (inputs(80));
    layer0_outputs(9527) <= not((inputs(116)) or (inputs(29)));
    layer0_outputs(9528) <= (inputs(141)) and not (inputs(35));
    layer0_outputs(9529) <= not((inputs(121)) or (inputs(158)));
    layer0_outputs(9530) <= not(inputs(225)) or (inputs(235));
    layer0_outputs(9531) <= (inputs(145)) xor (inputs(159));
    layer0_outputs(9532) <= (inputs(227)) or (inputs(90));
    layer0_outputs(9533) <= not((inputs(225)) xor (inputs(213)));
    layer0_outputs(9534) <= inputs(251);
    layer0_outputs(9535) <= '1';
    layer0_outputs(9536) <= (inputs(115)) and not (inputs(214));
    layer0_outputs(9537) <= inputs(25);
    layer0_outputs(9538) <= (inputs(252)) or (inputs(18));
    layer0_outputs(9539) <= not(inputs(253));
    layer0_outputs(9540) <= (inputs(5)) or (inputs(211));
    layer0_outputs(9541) <= not((inputs(169)) and (inputs(9)));
    layer0_outputs(9542) <= inputs(196);
    layer0_outputs(9543) <= inputs(214);
    layer0_outputs(9544) <= (inputs(152)) or (inputs(137));
    layer0_outputs(9545) <= (inputs(21)) xor (inputs(1));
    layer0_outputs(9546) <= not(inputs(228));
    layer0_outputs(9547) <= inputs(215);
    layer0_outputs(9548) <= (inputs(209)) and not (inputs(229));
    layer0_outputs(9549) <= inputs(11);
    layer0_outputs(9550) <= not(inputs(155)) or (inputs(75));
    layer0_outputs(9551) <= '1';
    layer0_outputs(9552) <= (inputs(156)) and not (inputs(208));
    layer0_outputs(9553) <= '1';
    layer0_outputs(9554) <= not(inputs(79));
    layer0_outputs(9555) <= (inputs(11)) and not (inputs(248));
    layer0_outputs(9556) <= not(inputs(224));
    layer0_outputs(9557) <= not(inputs(158)) or (inputs(93));
    layer0_outputs(9558) <= inputs(179);
    layer0_outputs(9559) <= (inputs(49)) and not (inputs(85));
    layer0_outputs(9560) <= '1';
    layer0_outputs(9561) <= not((inputs(133)) and (inputs(172)));
    layer0_outputs(9562) <= inputs(213);
    layer0_outputs(9563) <= not((inputs(88)) xor (inputs(191)));
    layer0_outputs(9564) <= not(inputs(190));
    layer0_outputs(9565) <= not(inputs(94));
    layer0_outputs(9566) <= not((inputs(236)) xor (inputs(143)));
    layer0_outputs(9567) <= '1';
    layer0_outputs(9568) <= (inputs(234)) and not (inputs(232));
    layer0_outputs(9569) <= not(inputs(230)) or (inputs(66));
    layer0_outputs(9570) <= not((inputs(215)) or (inputs(130)));
    layer0_outputs(9571) <= not(inputs(54)) or (inputs(132));
    layer0_outputs(9572) <= not(inputs(212));
    layer0_outputs(9573) <= not((inputs(157)) and (inputs(251)));
    layer0_outputs(9574) <= not(inputs(101));
    layer0_outputs(9575) <= (inputs(159)) and not (inputs(228));
    layer0_outputs(9576) <= (inputs(11)) and not (inputs(179));
    layer0_outputs(9577) <= not((inputs(113)) or (inputs(104)));
    layer0_outputs(9578) <= not(inputs(116));
    layer0_outputs(9579) <= not((inputs(197)) or (inputs(58)));
    layer0_outputs(9580) <= (inputs(173)) and not (inputs(80));
    layer0_outputs(9581) <= not((inputs(214)) or (inputs(0)));
    layer0_outputs(9582) <= not(inputs(42));
    layer0_outputs(9583) <= not((inputs(81)) xor (inputs(239)));
    layer0_outputs(9584) <= (inputs(37)) xor (inputs(29));
    layer0_outputs(9585) <= not(inputs(206));
    layer0_outputs(9586) <= not((inputs(55)) or (inputs(16)));
    layer0_outputs(9587) <= inputs(138);
    layer0_outputs(9588) <= not(inputs(73));
    layer0_outputs(9589) <= (inputs(183)) xor (inputs(244));
    layer0_outputs(9590) <= (inputs(113)) and (inputs(193));
    layer0_outputs(9591) <= '1';
    layer0_outputs(9592) <= (inputs(141)) and not (inputs(124));
    layer0_outputs(9593) <= (inputs(17)) and not (inputs(100));
    layer0_outputs(9594) <= not((inputs(110)) or (inputs(115)));
    layer0_outputs(9595) <= (inputs(187)) and not (inputs(150));
    layer0_outputs(9596) <= (inputs(239)) and not (inputs(235));
    layer0_outputs(9597) <= inputs(252);
    layer0_outputs(9598) <= not(inputs(243)) or (inputs(243));
    layer0_outputs(9599) <= not((inputs(253)) xor (inputs(234)));
    layer0_outputs(9600) <= (inputs(106)) and not (inputs(2));
    layer0_outputs(9601) <= '0';
    layer0_outputs(9602) <= (inputs(181)) xor (inputs(143));
    layer0_outputs(9603) <= (inputs(154)) and not (inputs(0));
    layer0_outputs(9604) <= (inputs(178)) xor (inputs(240));
    layer0_outputs(9605) <= not(inputs(163)) or (inputs(202));
    layer0_outputs(9606) <= (inputs(214)) or (inputs(232));
    layer0_outputs(9607) <= inputs(211);
    layer0_outputs(9608) <= (inputs(17)) and (inputs(218));
    layer0_outputs(9609) <= not(inputs(229)) or (inputs(200));
    layer0_outputs(9610) <= (inputs(86)) and (inputs(151));
    layer0_outputs(9611) <= (inputs(15)) and (inputs(248));
    layer0_outputs(9612) <= (inputs(162)) and not (inputs(44));
    layer0_outputs(9613) <= (inputs(254)) xor (inputs(140));
    layer0_outputs(9614) <= (inputs(48)) and (inputs(251));
    layer0_outputs(9615) <= '1';
    layer0_outputs(9616) <= '0';
    layer0_outputs(9617) <= not((inputs(92)) xor (inputs(240)));
    layer0_outputs(9618) <= not((inputs(173)) or (inputs(189)));
    layer0_outputs(9619) <= not(inputs(35));
    layer0_outputs(9620) <= not(inputs(170));
    layer0_outputs(9621) <= (inputs(187)) or (inputs(251));
    layer0_outputs(9622) <= (inputs(45)) or (inputs(234));
    layer0_outputs(9623) <= not(inputs(36));
    layer0_outputs(9624) <= (inputs(25)) or (inputs(137));
    layer0_outputs(9625) <= not(inputs(8)) or (inputs(222));
    layer0_outputs(9626) <= not((inputs(41)) and (inputs(197)));
    layer0_outputs(9627) <= '1';
    layer0_outputs(9628) <= (inputs(216)) or (inputs(244));
    layer0_outputs(9629) <= (inputs(136)) xor (inputs(22));
    layer0_outputs(9630) <= (inputs(26)) or (inputs(59));
    layer0_outputs(9631) <= not(inputs(127));
    layer0_outputs(9632) <= (inputs(231)) or (inputs(74));
    layer0_outputs(9633) <= (inputs(45)) or (inputs(53));
    layer0_outputs(9634) <= not(inputs(196));
    layer0_outputs(9635) <= not(inputs(185)) or (inputs(77));
    layer0_outputs(9636) <= (inputs(68)) xor (inputs(153));
    layer0_outputs(9637) <= (inputs(18)) and not (inputs(54));
    layer0_outputs(9638) <= not(inputs(97));
    layer0_outputs(9639) <= (inputs(67)) or (inputs(59));
    layer0_outputs(9640) <= not((inputs(95)) or (inputs(22)));
    layer0_outputs(9641) <= not((inputs(37)) or (inputs(137)));
    layer0_outputs(9642) <= inputs(107);
    layer0_outputs(9643) <= not(inputs(239)) or (inputs(195));
    layer0_outputs(9644) <= not(inputs(125));
    layer0_outputs(9645) <= inputs(149);
    layer0_outputs(9646) <= inputs(62);
    layer0_outputs(9647) <= not(inputs(118));
    layer0_outputs(9648) <= not(inputs(174)) or (inputs(111));
    layer0_outputs(9649) <= inputs(42);
    layer0_outputs(9650) <= not(inputs(73));
    layer0_outputs(9651) <= not((inputs(200)) and (inputs(161)));
    layer0_outputs(9652) <= not(inputs(162));
    layer0_outputs(9653) <= (inputs(118)) and not (inputs(0));
    layer0_outputs(9654) <= '0';
    layer0_outputs(9655) <= not(inputs(231)) or (inputs(35));
    layer0_outputs(9656) <= (inputs(165)) xor (inputs(176));
    layer0_outputs(9657) <= (inputs(141)) and not (inputs(113));
    layer0_outputs(9658) <= not((inputs(15)) xor (inputs(42)));
    layer0_outputs(9659) <= (inputs(14)) or (inputs(96));
    layer0_outputs(9660) <= not(inputs(106)) or (inputs(171));
    layer0_outputs(9661) <= not(inputs(3)) or (inputs(138));
    layer0_outputs(9662) <= inputs(148);
    layer0_outputs(9663) <= inputs(26);
    layer0_outputs(9664) <= not(inputs(98)) or (inputs(95));
    layer0_outputs(9665) <= not(inputs(175)) or (inputs(24));
    layer0_outputs(9666) <= not(inputs(77));
    layer0_outputs(9667) <= '1';
    layer0_outputs(9668) <= (inputs(216)) xor (inputs(232));
    layer0_outputs(9669) <= not(inputs(91));
    layer0_outputs(9670) <= (inputs(114)) and not (inputs(93));
    layer0_outputs(9671) <= not(inputs(175));
    layer0_outputs(9672) <= '0';
    layer0_outputs(9673) <= (inputs(160)) xor (inputs(155));
    layer0_outputs(9674) <= not(inputs(77)) or (inputs(32));
    layer0_outputs(9675) <= (inputs(71)) and not (inputs(224));
    layer0_outputs(9676) <= not(inputs(187)) or (inputs(119));
    layer0_outputs(9677) <= not((inputs(137)) and (inputs(42)));
    layer0_outputs(9678) <= inputs(94);
    layer0_outputs(9679) <= '0';
    layer0_outputs(9680) <= not(inputs(184)) or (inputs(190));
    layer0_outputs(9681) <= (inputs(177)) and not (inputs(11));
    layer0_outputs(9682) <= not(inputs(185));
    layer0_outputs(9683) <= not((inputs(107)) or (inputs(84)));
    layer0_outputs(9684) <= not((inputs(162)) or (inputs(186)));
    layer0_outputs(9685) <= not(inputs(246));
    layer0_outputs(9686) <= (inputs(210)) and not (inputs(248));
    layer0_outputs(9687) <= inputs(222);
    layer0_outputs(9688) <= not((inputs(178)) or (inputs(162)));
    layer0_outputs(9689) <= not((inputs(10)) or (inputs(116)));
    layer0_outputs(9690) <= not(inputs(76));
    layer0_outputs(9691) <= (inputs(242)) and (inputs(217));
    layer0_outputs(9692) <= (inputs(10)) xor (inputs(20));
    layer0_outputs(9693) <= (inputs(117)) xor (inputs(119));
    layer0_outputs(9694) <= not(inputs(143)) or (inputs(25));
    layer0_outputs(9695) <= (inputs(227)) or (inputs(223));
    layer0_outputs(9696) <= (inputs(76)) and (inputs(49));
    layer0_outputs(9697) <= not(inputs(154)) or (inputs(30));
    layer0_outputs(9698) <= (inputs(20)) and not (inputs(157));
    layer0_outputs(9699) <= not((inputs(8)) and (inputs(92)));
    layer0_outputs(9700) <= not(inputs(113));
    layer0_outputs(9701) <= not(inputs(63)) or (inputs(48));
    layer0_outputs(9702) <= not(inputs(54));
    layer0_outputs(9703) <= not((inputs(81)) xor (inputs(124)));
    layer0_outputs(9704) <= not(inputs(137));
    layer0_outputs(9705) <= (inputs(110)) and (inputs(246));
    layer0_outputs(9706) <= (inputs(16)) or (inputs(148));
    layer0_outputs(9707) <= inputs(77);
    layer0_outputs(9708) <= inputs(77);
    layer0_outputs(9709) <= (inputs(32)) or (inputs(227));
    layer0_outputs(9710) <= not((inputs(128)) and (inputs(171)));
    layer0_outputs(9711) <= (inputs(167)) and not (inputs(121));
    layer0_outputs(9712) <= not(inputs(189));
    layer0_outputs(9713) <= (inputs(105)) and not (inputs(88));
    layer0_outputs(9714) <= not((inputs(25)) or (inputs(95)));
    layer0_outputs(9715) <= inputs(79);
    layer0_outputs(9716) <= not(inputs(225)) or (inputs(251));
    layer0_outputs(9717) <= inputs(71);
    layer0_outputs(9718) <= (inputs(98)) xor (inputs(249));
    layer0_outputs(9719) <= '0';
    layer0_outputs(9720) <= not(inputs(171));
    layer0_outputs(9721) <= not(inputs(198));
    layer0_outputs(9722) <= not(inputs(138));
    layer0_outputs(9723) <= inputs(91);
    layer0_outputs(9724) <= (inputs(235)) and not (inputs(178));
    layer0_outputs(9725) <= not(inputs(203));
    layer0_outputs(9726) <= not(inputs(20)) or (inputs(108));
    layer0_outputs(9727) <= not((inputs(221)) xor (inputs(114)));
    layer0_outputs(9728) <= not(inputs(61));
    layer0_outputs(9729) <= (inputs(129)) and (inputs(75));
    layer0_outputs(9730) <= (inputs(191)) xor (inputs(207));
    layer0_outputs(9731) <= not(inputs(218));
    layer0_outputs(9732) <= inputs(172);
    layer0_outputs(9733) <= (inputs(165)) or (inputs(117));
    layer0_outputs(9734) <= not((inputs(128)) or (inputs(97)));
    layer0_outputs(9735) <= not(inputs(61)) or (inputs(229));
    layer0_outputs(9736) <= not(inputs(218));
    layer0_outputs(9737) <= not((inputs(220)) or (inputs(136)));
    layer0_outputs(9738) <= (inputs(116)) xor (inputs(219));
    layer0_outputs(9739) <= not((inputs(235)) and (inputs(129)));
    layer0_outputs(9740) <= not((inputs(30)) and (inputs(176)));
    layer0_outputs(9741) <= (inputs(136)) and (inputs(173));
    layer0_outputs(9742) <= not((inputs(137)) or (inputs(250)));
    layer0_outputs(9743) <= (inputs(246)) and not (inputs(108));
    layer0_outputs(9744) <= inputs(245);
    layer0_outputs(9745) <= not(inputs(84));
    layer0_outputs(9746) <= not(inputs(39));
    layer0_outputs(9747) <= (inputs(50)) and not (inputs(112));
    layer0_outputs(9748) <= not((inputs(153)) or (inputs(61)));
    layer0_outputs(9749) <= (inputs(25)) and not (inputs(96));
    layer0_outputs(9750) <= (inputs(147)) or (inputs(209));
    layer0_outputs(9751) <= not(inputs(136));
    layer0_outputs(9752) <= '1';
    layer0_outputs(9753) <= not(inputs(138)) or (inputs(237));
    layer0_outputs(9754) <= '0';
    layer0_outputs(9755) <= '1';
    layer0_outputs(9756) <= (inputs(135)) xor (inputs(50));
    layer0_outputs(9757) <= (inputs(210)) and (inputs(12));
    layer0_outputs(9758) <= inputs(126);
    layer0_outputs(9759) <= not((inputs(59)) and (inputs(167)));
    layer0_outputs(9760) <= (inputs(140)) xor (inputs(4));
    layer0_outputs(9761) <= inputs(65);
    layer0_outputs(9762) <= not((inputs(170)) and (inputs(21)));
    layer0_outputs(9763) <= (inputs(231)) and not (inputs(208));
    layer0_outputs(9764) <= '1';
    layer0_outputs(9765) <= not(inputs(6)) or (inputs(169));
    layer0_outputs(9766) <= inputs(77);
    layer0_outputs(9767) <= (inputs(216)) and (inputs(17));
    layer0_outputs(9768) <= not(inputs(182)) or (inputs(174));
    layer0_outputs(9769) <= not(inputs(224)) or (inputs(205));
    layer0_outputs(9770) <= not((inputs(93)) or (inputs(230)));
    layer0_outputs(9771) <= not((inputs(123)) or (inputs(64)));
    layer0_outputs(9772) <= not((inputs(69)) xor (inputs(196)));
    layer0_outputs(9773) <= not(inputs(157)) or (inputs(95));
    layer0_outputs(9774) <= not((inputs(144)) or (inputs(196)));
    layer0_outputs(9775) <= not((inputs(132)) and (inputs(213)));
    layer0_outputs(9776) <= '0';
    layer0_outputs(9777) <= inputs(121);
    layer0_outputs(9778) <= (inputs(13)) xor (inputs(109));
    layer0_outputs(9779) <= inputs(33);
    layer0_outputs(9780) <= (inputs(222)) and not (inputs(243));
    layer0_outputs(9781) <= not(inputs(220));
    layer0_outputs(9782) <= (inputs(20)) or (inputs(42));
    layer0_outputs(9783) <= inputs(108);
    layer0_outputs(9784) <= (inputs(147)) or (inputs(38));
    layer0_outputs(9785) <= (inputs(89)) or (inputs(30));
    layer0_outputs(9786) <= not(inputs(255));
    layer0_outputs(9787) <= not(inputs(116)) or (inputs(20));
    layer0_outputs(9788) <= not((inputs(228)) and (inputs(203)));
    layer0_outputs(9789) <= not(inputs(216));
    layer0_outputs(9790) <= (inputs(228)) and not (inputs(218));
    layer0_outputs(9791) <= not(inputs(25)) or (inputs(128));
    layer0_outputs(9792) <= not((inputs(46)) xor (inputs(98)));
    layer0_outputs(9793) <= inputs(184);
    layer0_outputs(9794) <= not((inputs(186)) xor (inputs(12)));
    layer0_outputs(9795) <= '1';
    layer0_outputs(9796) <= not(inputs(99)) or (inputs(62));
    layer0_outputs(9797) <= not((inputs(93)) xor (inputs(192)));
    layer0_outputs(9798) <= not((inputs(126)) xor (inputs(8)));
    layer0_outputs(9799) <= '1';
    layer0_outputs(9800) <= not(inputs(36)) or (inputs(85));
    layer0_outputs(9801) <= not((inputs(109)) or (inputs(132)));
    layer0_outputs(9802) <= not(inputs(89));
    layer0_outputs(9803) <= (inputs(183)) xor (inputs(255));
    layer0_outputs(9804) <= inputs(206);
    layer0_outputs(9805) <= (inputs(131)) or (inputs(118));
    layer0_outputs(9806) <= not((inputs(5)) or (inputs(16)));
    layer0_outputs(9807) <= inputs(140);
    layer0_outputs(9808) <= '1';
    layer0_outputs(9809) <= not(inputs(183)) or (inputs(12));
    layer0_outputs(9810) <= not(inputs(12));
    layer0_outputs(9811) <= (inputs(24)) xor (inputs(136));
    layer0_outputs(9812) <= (inputs(39)) or (inputs(57));
    layer0_outputs(9813) <= inputs(108);
    layer0_outputs(9814) <= not(inputs(125));
    layer0_outputs(9815) <= not(inputs(57)) or (inputs(227));
    layer0_outputs(9816) <= inputs(250);
    layer0_outputs(9817) <= not((inputs(174)) xor (inputs(232)));
    layer0_outputs(9818) <= inputs(195);
    layer0_outputs(9819) <= (inputs(79)) xor (inputs(58));
    layer0_outputs(9820) <= not((inputs(128)) xor (inputs(45)));
    layer0_outputs(9821) <= not(inputs(178)) or (inputs(184));
    layer0_outputs(9822) <= not((inputs(85)) or (inputs(239)));
    layer0_outputs(9823) <= (inputs(182)) and not (inputs(160));
    layer0_outputs(9824) <= not((inputs(119)) xor (inputs(241)));
    layer0_outputs(9825) <= '0';
    layer0_outputs(9826) <= (inputs(95)) and not (inputs(98));
    layer0_outputs(9827) <= not((inputs(95)) xor (inputs(215)));
    layer0_outputs(9828) <= not(inputs(127));
    layer0_outputs(9829) <= not((inputs(152)) xor (inputs(189)));
    layer0_outputs(9830) <= not(inputs(34)) or (inputs(26));
    layer0_outputs(9831) <= not((inputs(107)) xor (inputs(30)));
    layer0_outputs(9832) <= not((inputs(18)) and (inputs(185)));
    layer0_outputs(9833) <= not(inputs(175)) or (inputs(202));
    layer0_outputs(9834) <= (inputs(215)) xor (inputs(45));
    layer0_outputs(9835) <= not((inputs(101)) and (inputs(23)));
    layer0_outputs(9836) <= (inputs(124)) xor (inputs(93));
    layer0_outputs(9837) <= not(inputs(101));
    layer0_outputs(9838) <= inputs(160);
    layer0_outputs(9839) <= not((inputs(1)) and (inputs(64)));
    layer0_outputs(9840) <= (inputs(109)) or (inputs(211));
    layer0_outputs(9841) <= not((inputs(37)) xor (inputs(3)));
    layer0_outputs(9842) <= inputs(152);
    layer0_outputs(9843) <= not(inputs(154)) or (inputs(174));
    layer0_outputs(9844) <= not(inputs(152));
    layer0_outputs(9845) <= inputs(113);
    layer0_outputs(9846) <= '1';
    layer0_outputs(9847) <= not((inputs(159)) and (inputs(72)));
    layer0_outputs(9848) <= not((inputs(169)) xor (inputs(175)));
    layer0_outputs(9849) <= not(inputs(196)) or (inputs(30));
    layer0_outputs(9850) <= not(inputs(186)) or (inputs(45));
    layer0_outputs(9851) <= not((inputs(94)) xor (inputs(229)));
    layer0_outputs(9852) <= inputs(236);
    layer0_outputs(9853) <= inputs(185);
    layer0_outputs(9854) <= inputs(89);
    layer0_outputs(9855) <= not((inputs(5)) xor (inputs(196)));
    layer0_outputs(9856) <= not((inputs(54)) or (inputs(214)));
    layer0_outputs(9857) <= (inputs(190)) and not (inputs(165));
    layer0_outputs(9858) <= not((inputs(61)) or (inputs(104)));
    layer0_outputs(9859) <= (inputs(119)) and not (inputs(224));
    layer0_outputs(9860) <= not(inputs(71));
    layer0_outputs(9861) <= (inputs(165)) or (inputs(65));
    layer0_outputs(9862) <= not(inputs(129));
    layer0_outputs(9863) <= inputs(133);
    layer0_outputs(9864) <= not(inputs(116));
    layer0_outputs(9865) <= (inputs(17)) and not (inputs(245));
    layer0_outputs(9866) <= not(inputs(104)) or (inputs(76));
    layer0_outputs(9867) <= not((inputs(34)) xor (inputs(101)));
    layer0_outputs(9868) <= not(inputs(210)) or (inputs(65));
    layer0_outputs(9869) <= not(inputs(175));
    layer0_outputs(9870) <= not(inputs(161));
    layer0_outputs(9871) <= inputs(150);
    layer0_outputs(9872) <= not(inputs(232)) or (inputs(24));
    layer0_outputs(9873) <= inputs(220);
    layer0_outputs(9874) <= not(inputs(195));
    layer0_outputs(9875) <= not((inputs(221)) and (inputs(149)));
    layer0_outputs(9876) <= (inputs(58)) and (inputs(175));
    layer0_outputs(9877) <= inputs(3);
    layer0_outputs(9878) <= (inputs(124)) and not (inputs(137));
    layer0_outputs(9879) <= inputs(193);
    layer0_outputs(9880) <= (inputs(91)) xor (inputs(168));
    layer0_outputs(9881) <= (inputs(149)) or (inputs(7));
    layer0_outputs(9882) <= inputs(59);
    layer0_outputs(9883) <= (inputs(56)) and not (inputs(89));
    layer0_outputs(9884) <= inputs(168);
    layer0_outputs(9885) <= not(inputs(247)) or (inputs(190));
    layer0_outputs(9886) <= (inputs(132)) xor (inputs(3));
    layer0_outputs(9887) <= not(inputs(2));
    layer0_outputs(9888) <= inputs(145);
    layer0_outputs(9889) <= (inputs(249)) xor (inputs(184));
    layer0_outputs(9890) <= (inputs(134)) or (inputs(143));
    layer0_outputs(9891) <= inputs(189);
    layer0_outputs(9892) <= inputs(167);
    layer0_outputs(9893) <= not(inputs(137));
    layer0_outputs(9894) <= (inputs(244)) xor (inputs(246));
    layer0_outputs(9895) <= (inputs(198)) and not (inputs(189));
    layer0_outputs(9896) <= not(inputs(126));
    layer0_outputs(9897) <= not(inputs(145));
    layer0_outputs(9898) <= '0';
    layer0_outputs(9899) <= (inputs(247)) xor (inputs(38));
    layer0_outputs(9900) <= not(inputs(204));
    layer0_outputs(9901) <= (inputs(175)) and not (inputs(218));
    layer0_outputs(9902) <= inputs(111);
    layer0_outputs(9903) <= not(inputs(27));
    layer0_outputs(9904) <= not((inputs(67)) and (inputs(82)));
    layer0_outputs(9905) <= (inputs(169)) xor (inputs(10));
    layer0_outputs(9906) <= '0';
    layer0_outputs(9907) <= not(inputs(125)) or (inputs(6));
    layer0_outputs(9908) <= (inputs(130)) or (inputs(72));
    layer0_outputs(9909) <= not(inputs(176)) or (inputs(254));
    layer0_outputs(9910) <= '1';
    layer0_outputs(9911) <= not(inputs(140));
    layer0_outputs(9912) <= (inputs(24)) and (inputs(4));
    layer0_outputs(9913) <= inputs(179);
    layer0_outputs(9914) <= not(inputs(26));
    layer0_outputs(9915) <= (inputs(35)) or (inputs(164));
    layer0_outputs(9916) <= not((inputs(9)) xor (inputs(83)));
    layer0_outputs(9917) <= inputs(235);
    layer0_outputs(9918) <= not((inputs(23)) or (inputs(68)));
    layer0_outputs(9919) <= not((inputs(63)) or (inputs(154)));
    layer0_outputs(9920) <= inputs(129);
    layer0_outputs(9921) <= not(inputs(148));
    layer0_outputs(9922) <= not(inputs(232));
    layer0_outputs(9923) <= (inputs(0)) and not (inputs(236));
    layer0_outputs(9924) <= '0';
    layer0_outputs(9925) <= not(inputs(153)) or (inputs(23));
    layer0_outputs(9926) <= not((inputs(14)) or (inputs(19)));
    layer0_outputs(9927) <= not((inputs(80)) xor (inputs(38)));
    layer0_outputs(9928) <= not(inputs(84));
    layer0_outputs(9929) <= '0';
    layer0_outputs(9930) <= (inputs(54)) xor (inputs(1));
    layer0_outputs(9931) <= not((inputs(236)) xor (inputs(231)));
    layer0_outputs(9932) <= not((inputs(158)) xor (inputs(109)));
    layer0_outputs(9933) <= not(inputs(233));
    layer0_outputs(9934) <= (inputs(120)) xor (inputs(237));
    layer0_outputs(9935) <= inputs(64);
    layer0_outputs(9936) <= (inputs(215)) xor (inputs(253));
    layer0_outputs(9937) <= not(inputs(116));
    layer0_outputs(9938) <= not((inputs(7)) xor (inputs(115)));
    layer0_outputs(9939) <= not(inputs(23));
    layer0_outputs(9940) <= '0';
    layer0_outputs(9941) <= (inputs(156)) or (inputs(154));
    layer0_outputs(9942) <= (inputs(5)) and not (inputs(145));
    layer0_outputs(9943) <= (inputs(164)) or (inputs(202));
    layer0_outputs(9944) <= not(inputs(39)) or (inputs(178));
    layer0_outputs(9945) <= not((inputs(232)) or (inputs(83)));
    layer0_outputs(9946) <= not(inputs(94)) or (inputs(79));
    layer0_outputs(9947) <= not(inputs(17)) or (inputs(238));
    layer0_outputs(9948) <= (inputs(244)) xor (inputs(179));
    layer0_outputs(9949) <= not(inputs(141));
    layer0_outputs(9950) <= not(inputs(209)) or (inputs(64));
    layer0_outputs(9951) <= not((inputs(61)) and (inputs(228)));
    layer0_outputs(9952) <= (inputs(144)) and not (inputs(192));
    layer0_outputs(9953) <= inputs(48);
    layer0_outputs(9954) <= (inputs(172)) and (inputs(96));
    layer0_outputs(9955) <= not((inputs(204)) or (inputs(70)));
    layer0_outputs(9956) <= not(inputs(216));
    layer0_outputs(9957) <= not(inputs(235)) or (inputs(173));
    layer0_outputs(9958) <= (inputs(231)) xor (inputs(1));
    layer0_outputs(9959) <= inputs(29);
    layer0_outputs(9960) <= not(inputs(207)) or (inputs(74));
    layer0_outputs(9961) <= not(inputs(30));
    layer0_outputs(9962) <= not(inputs(145)) or (inputs(87));
    layer0_outputs(9963) <= (inputs(153)) xor (inputs(69));
    layer0_outputs(9964) <= not((inputs(179)) or (inputs(86)));
    layer0_outputs(9965) <= '1';
    layer0_outputs(9966) <= not(inputs(225));
    layer0_outputs(9967) <= not(inputs(179)) or (inputs(103));
    layer0_outputs(9968) <= '0';
    layer0_outputs(9969) <= not(inputs(181));
    layer0_outputs(9970) <= (inputs(241)) xor (inputs(239));
    layer0_outputs(9971) <= not(inputs(151)) or (inputs(147));
    layer0_outputs(9972) <= inputs(65);
    layer0_outputs(9973) <= not(inputs(134));
    layer0_outputs(9974) <= (inputs(191)) xor (inputs(118));
    layer0_outputs(9975) <= not(inputs(134));
    layer0_outputs(9976) <= (inputs(236)) or (inputs(60));
    layer0_outputs(9977) <= (inputs(166)) and not (inputs(105));
    layer0_outputs(9978) <= '0';
    layer0_outputs(9979) <= (inputs(166)) and not (inputs(210));
    layer0_outputs(9980) <= not(inputs(73));
    layer0_outputs(9981) <= '1';
    layer0_outputs(9982) <= not((inputs(94)) or (inputs(241)));
    layer0_outputs(9983) <= not((inputs(197)) xor (inputs(12)));
    layer0_outputs(9984) <= (inputs(133)) and not (inputs(227));
    layer0_outputs(9985) <= (inputs(54)) or (inputs(192));
    layer0_outputs(9986) <= not(inputs(55)) or (inputs(232));
    layer0_outputs(9987) <= not(inputs(225)) or (inputs(222));
    layer0_outputs(9988) <= not(inputs(182)) or (inputs(178));
    layer0_outputs(9989) <= not((inputs(135)) or (inputs(79)));
    layer0_outputs(9990) <= not(inputs(237));
    layer0_outputs(9991) <= (inputs(63)) or (inputs(175));
    layer0_outputs(9992) <= inputs(80);
    layer0_outputs(9993) <= (inputs(60)) or (inputs(75));
    layer0_outputs(9994) <= inputs(72);
    layer0_outputs(9995) <= '0';
    layer0_outputs(9996) <= (inputs(254)) xor (inputs(85));
    layer0_outputs(9997) <= not(inputs(95)) or (inputs(157));
    layer0_outputs(9998) <= not(inputs(95));
    layer0_outputs(9999) <= (inputs(17)) xor (inputs(187));
    layer0_outputs(10000) <= (inputs(161)) and (inputs(76));
    layer0_outputs(10001) <= (inputs(5)) and not (inputs(185));
    layer0_outputs(10002) <= not(inputs(41)) or (inputs(11));
    layer0_outputs(10003) <= not((inputs(206)) xor (inputs(18)));
    layer0_outputs(10004) <= (inputs(230)) and (inputs(38));
    layer0_outputs(10005) <= not((inputs(69)) or (inputs(139)));
    layer0_outputs(10006) <= (inputs(205)) and not (inputs(44));
    layer0_outputs(10007) <= (inputs(208)) and not (inputs(162));
    layer0_outputs(10008) <= not((inputs(167)) or (inputs(242)));
    layer0_outputs(10009) <= (inputs(20)) or (inputs(207));
    layer0_outputs(10010) <= '0';
    layer0_outputs(10011) <= (inputs(176)) xor (inputs(0));
    layer0_outputs(10012) <= not(inputs(61));
    layer0_outputs(10013) <= (inputs(251)) or (inputs(91));
    layer0_outputs(10014) <= not((inputs(82)) or (inputs(213)));
    layer0_outputs(10015) <= (inputs(116)) xor (inputs(27));
    layer0_outputs(10016) <= '0';
    layer0_outputs(10017) <= not((inputs(254)) and (inputs(54)));
    layer0_outputs(10018) <= not(inputs(135)) or (inputs(182));
    layer0_outputs(10019) <= (inputs(10)) or (inputs(11));
    layer0_outputs(10020) <= not(inputs(194));
    layer0_outputs(10021) <= not((inputs(19)) xor (inputs(132)));
    layer0_outputs(10022) <= not(inputs(222));
    layer0_outputs(10023) <= inputs(12);
    layer0_outputs(10024) <= (inputs(194)) and (inputs(123));
    layer0_outputs(10025) <= (inputs(219)) and not (inputs(225));
    layer0_outputs(10026) <= not(inputs(168)) or (inputs(59));
    layer0_outputs(10027) <= (inputs(64)) or (inputs(214));
    layer0_outputs(10028) <= not((inputs(58)) or (inputs(62)));
    layer0_outputs(10029) <= inputs(83);
    layer0_outputs(10030) <= (inputs(150)) or (inputs(144));
    layer0_outputs(10031) <= not((inputs(32)) or (inputs(33)));
    layer0_outputs(10032) <= (inputs(106)) xor (inputs(108));
    layer0_outputs(10033) <= (inputs(196)) or (inputs(9));
    layer0_outputs(10034) <= not(inputs(230));
    layer0_outputs(10035) <= not((inputs(226)) or (inputs(44)));
    layer0_outputs(10036) <= not((inputs(34)) xor (inputs(31)));
    layer0_outputs(10037) <= inputs(174);
    layer0_outputs(10038) <= not((inputs(133)) and (inputs(156)));
    layer0_outputs(10039) <= (inputs(120)) and not (inputs(203));
    layer0_outputs(10040) <= (inputs(15)) xor (inputs(59));
    layer0_outputs(10041) <= (inputs(195)) and (inputs(160));
    layer0_outputs(10042) <= not(inputs(37)) or (inputs(114));
    layer0_outputs(10043) <= not(inputs(211));
    layer0_outputs(10044) <= not((inputs(33)) and (inputs(67)));
    layer0_outputs(10045) <= not(inputs(199)) or (inputs(111));
    layer0_outputs(10046) <= not(inputs(208)) or (inputs(88));
    layer0_outputs(10047) <= not(inputs(19));
    layer0_outputs(10048) <= inputs(36);
    layer0_outputs(10049) <= (inputs(235)) or (inputs(154));
    layer0_outputs(10050) <= not(inputs(72)) or (inputs(35));
    layer0_outputs(10051) <= '0';
    layer0_outputs(10052) <= not(inputs(211));
    layer0_outputs(10053) <= not((inputs(106)) xor (inputs(78)));
    layer0_outputs(10054) <= (inputs(57)) and not (inputs(184));
    layer0_outputs(10055) <= inputs(146);
    layer0_outputs(10056) <= not((inputs(142)) and (inputs(28)));
    layer0_outputs(10057) <= not(inputs(99)) or (inputs(141));
    layer0_outputs(10058) <= (inputs(198)) and not (inputs(158));
    layer0_outputs(10059) <= not((inputs(47)) or (inputs(50)));
    layer0_outputs(10060) <= (inputs(162)) xor (inputs(96));
    layer0_outputs(10061) <= (inputs(86)) or (inputs(109));
    layer0_outputs(10062) <= (inputs(188)) and not (inputs(97));
    layer0_outputs(10063) <= inputs(106);
    layer0_outputs(10064) <= (inputs(147)) or (inputs(92));
    layer0_outputs(10065) <= inputs(190);
    layer0_outputs(10066) <= not((inputs(168)) or (inputs(99)));
    layer0_outputs(10067) <= not(inputs(68));
    layer0_outputs(10068) <= inputs(132);
    layer0_outputs(10069) <= inputs(158);
    layer0_outputs(10070) <= '0';
    layer0_outputs(10071) <= (inputs(143)) or (inputs(227));
    layer0_outputs(10072) <= not(inputs(117));
    layer0_outputs(10073) <= (inputs(206)) or (inputs(58));
    layer0_outputs(10074) <= not(inputs(177));
    layer0_outputs(10075) <= (inputs(66)) xor (inputs(194));
    layer0_outputs(10076) <= not(inputs(98)) or (inputs(100));
    layer0_outputs(10077) <= (inputs(151)) and not (inputs(68));
    layer0_outputs(10078) <= (inputs(88)) and (inputs(100));
    layer0_outputs(10079) <= not((inputs(5)) and (inputs(213)));
    layer0_outputs(10080) <= not((inputs(133)) xor (inputs(34)));
    layer0_outputs(10081) <= (inputs(96)) and not (inputs(103));
    layer0_outputs(10082) <= inputs(155);
    layer0_outputs(10083) <= not(inputs(198));
    layer0_outputs(10084) <= not((inputs(24)) xor (inputs(145)));
    layer0_outputs(10085) <= (inputs(109)) xor (inputs(231));
    layer0_outputs(10086) <= '0';
    layer0_outputs(10087) <= inputs(243);
    layer0_outputs(10088) <= (inputs(3)) xor (inputs(236));
    layer0_outputs(10089) <= (inputs(32)) and not (inputs(219));
    layer0_outputs(10090) <= not((inputs(190)) or (inputs(83)));
    layer0_outputs(10091) <= inputs(118);
    layer0_outputs(10092) <= (inputs(170)) and not (inputs(3));
    layer0_outputs(10093) <= '1';
    layer0_outputs(10094) <= (inputs(122)) and not (inputs(72));
    layer0_outputs(10095) <= (inputs(65)) and not (inputs(3));
    layer0_outputs(10096) <= (inputs(179)) and not (inputs(72));
    layer0_outputs(10097) <= not((inputs(46)) or (inputs(134)));
    layer0_outputs(10098) <= (inputs(99)) and not (inputs(110));
    layer0_outputs(10099) <= inputs(201);
    layer0_outputs(10100) <= inputs(242);
    layer0_outputs(10101) <= inputs(130);
    layer0_outputs(10102) <= not((inputs(247)) or (inputs(13)));
    layer0_outputs(10103) <= not(inputs(76));
    layer0_outputs(10104) <= not(inputs(52));
    layer0_outputs(10105) <= (inputs(189)) or (inputs(117));
    layer0_outputs(10106) <= '1';
    layer0_outputs(10107) <= not((inputs(33)) and (inputs(169)));
    layer0_outputs(10108) <= inputs(132);
    layer0_outputs(10109) <= (inputs(20)) and (inputs(166));
    layer0_outputs(10110) <= (inputs(123)) and not (inputs(252));
    layer0_outputs(10111) <= not(inputs(99));
    layer0_outputs(10112) <= (inputs(135)) or (inputs(143));
    layer0_outputs(10113) <= not(inputs(194));
    layer0_outputs(10114) <= not((inputs(208)) or (inputs(89)));
    layer0_outputs(10115) <= not((inputs(209)) xor (inputs(88)));
    layer0_outputs(10116) <= not(inputs(233));
    layer0_outputs(10117) <= not((inputs(255)) or (inputs(203)));
    layer0_outputs(10118) <= (inputs(73)) and (inputs(60));
    layer0_outputs(10119) <= not(inputs(72)) or (inputs(203));
    layer0_outputs(10120) <= not((inputs(183)) or (inputs(197)));
    layer0_outputs(10121) <= not(inputs(224)) or (inputs(213));
    layer0_outputs(10122) <= not(inputs(81));
    layer0_outputs(10123) <= inputs(229);
    layer0_outputs(10124) <= (inputs(116)) and not (inputs(220));
    layer0_outputs(10125) <= not(inputs(2)) or (inputs(21));
    layer0_outputs(10126) <= (inputs(158)) and not (inputs(213));
    layer0_outputs(10127) <= inputs(180);
    layer0_outputs(10128) <= (inputs(249)) or (inputs(74));
    layer0_outputs(10129) <= (inputs(66)) xor (inputs(39));
    layer0_outputs(10130) <= not(inputs(65)) or (inputs(150));
    layer0_outputs(10131) <= not(inputs(172)) or (inputs(205));
    layer0_outputs(10132) <= (inputs(229)) or (inputs(176));
    layer0_outputs(10133) <= inputs(137);
    layer0_outputs(10134) <= inputs(197);
    layer0_outputs(10135) <= not(inputs(115)) or (inputs(103));
    layer0_outputs(10136) <= '1';
    layer0_outputs(10137) <= not((inputs(85)) and (inputs(24)));
    layer0_outputs(10138) <= inputs(236);
    layer0_outputs(10139) <= not(inputs(77));
    layer0_outputs(10140) <= (inputs(224)) and not (inputs(114));
    layer0_outputs(10141) <= not((inputs(182)) or (inputs(40)));
    layer0_outputs(10142) <= (inputs(188)) and (inputs(213));
    layer0_outputs(10143) <= (inputs(149)) and not (inputs(229));
    layer0_outputs(10144) <= not(inputs(98));
    layer0_outputs(10145) <= not(inputs(114)) or (inputs(136));
    layer0_outputs(10146) <= inputs(118);
    layer0_outputs(10147) <= not((inputs(165)) xor (inputs(18)));
    layer0_outputs(10148) <= inputs(169);
    layer0_outputs(10149) <= not(inputs(129));
    layer0_outputs(10150) <= not((inputs(144)) or (inputs(173)));
    layer0_outputs(10151) <= not(inputs(247));
    layer0_outputs(10152) <= inputs(147);
    layer0_outputs(10153) <= not(inputs(215)) or (inputs(203));
    layer0_outputs(10154) <= not(inputs(193));
    layer0_outputs(10155) <= not(inputs(193)) or (inputs(198));
    layer0_outputs(10156) <= (inputs(146)) and not (inputs(195));
    layer0_outputs(10157) <= not(inputs(59));
    layer0_outputs(10158) <= not(inputs(162));
    layer0_outputs(10159) <= not((inputs(156)) and (inputs(183)));
    layer0_outputs(10160) <= (inputs(156)) and not (inputs(236));
    layer0_outputs(10161) <= not((inputs(18)) xor (inputs(169)));
    layer0_outputs(10162) <= (inputs(89)) or (inputs(161));
    layer0_outputs(10163) <= not((inputs(190)) and (inputs(158)));
    layer0_outputs(10164) <= not(inputs(150));
    layer0_outputs(10165) <= inputs(160);
    layer0_outputs(10166) <= (inputs(92)) and not (inputs(146));
    layer0_outputs(10167) <= not(inputs(88)) or (inputs(109));
    layer0_outputs(10168) <= not(inputs(87)) or (inputs(156));
    layer0_outputs(10169) <= (inputs(228)) or (inputs(50));
    layer0_outputs(10170) <= '0';
    layer0_outputs(10171) <= (inputs(18)) and (inputs(161));
    layer0_outputs(10172) <= inputs(73);
    layer0_outputs(10173) <= not(inputs(88));
    layer0_outputs(10174) <= not((inputs(62)) xor (inputs(23)));
    layer0_outputs(10175) <= not(inputs(196));
    layer0_outputs(10176) <= '0';
    layer0_outputs(10177) <= not(inputs(90));
    layer0_outputs(10178) <= not(inputs(67));
    layer0_outputs(10179) <= not((inputs(181)) or (inputs(1)));
    layer0_outputs(10180) <= (inputs(29)) and not (inputs(246));
    layer0_outputs(10181) <= (inputs(181)) or (inputs(125));
    layer0_outputs(10182) <= (inputs(150)) or (inputs(140));
    layer0_outputs(10183) <= (inputs(207)) and (inputs(126));
    layer0_outputs(10184) <= not((inputs(30)) or (inputs(221)));
    layer0_outputs(10185) <= not((inputs(133)) or (inputs(165)));
    layer0_outputs(10186) <= (inputs(65)) xor (inputs(84));
    layer0_outputs(10187) <= inputs(149);
    layer0_outputs(10188) <= not(inputs(194)) or (inputs(204));
    layer0_outputs(10189) <= not(inputs(41));
    layer0_outputs(10190) <= (inputs(85)) or (inputs(20));
    layer0_outputs(10191) <= not(inputs(60)) or (inputs(238));
    layer0_outputs(10192) <= not((inputs(237)) xor (inputs(35)));
    layer0_outputs(10193) <= not(inputs(134));
    layer0_outputs(10194) <= '1';
    layer0_outputs(10195) <= not(inputs(231));
    layer0_outputs(10196) <= not((inputs(71)) or (inputs(95)));
    layer0_outputs(10197) <= inputs(107);
    layer0_outputs(10198) <= not((inputs(124)) and (inputs(33)));
    layer0_outputs(10199) <= not(inputs(27)) or (inputs(2));
    layer0_outputs(10200) <= (inputs(68)) and not (inputs(190));
    layer0_outputs(10201) <= (inputs(243)) and not (inputs(21));
    layer0_outputs(10202) <= inputs(175);
    layer0_outputs(10203) <= not((inputs(201)) or (inputs(93)));
    layer0_outputs(10204) <= not(inputs(186)) or (inputs(220));
    layer0_outputs(10205) <= not(inputs(153)) or (inputs(198));
    layer0_outputs(10206) <= (inputs(226)) and not (inputs(206));
    layer0_outputs(10207) <= inputs(130);
    layer0_outputs(10208) <= (inputs(40)) and (inputs(46));
    layer0_outputs(10209) <= not(inputs(204)) or (inputs(31));
    layer0_outputs(10210) <= not(inputs(198)) or (inputs(127));
    layer0_outputs(10211) <= not(inputs(28));
    layer0_outputs(10212) <= not((inputs(13)) and (inputs(104)));
    layer0_outputs(10213) <= inputs(237);
    layer0_outputs(10214) <= not(inputs(168));
    layer0_outputs(10215) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(10216) <= '1';
    layer0_outputs(10217) <= (inputs(125)) or (inputs(100));
    layer0_outputs(10218) <= (inputs(16)) xor (inputs(207));
    layer0_outputs(10219) <= not((inputs(30)) xor (inputs(157)));
    layer0_outputs(10220) <= (inputs(236)) and not (inputs(59));
    layer0_outputs(10221) <= not((inputs(29)) xor (inputs(222)));
    layer0_outputs(10222) <= not((inputs(165)) or (inputs(117)));
    layer0_outputs(10223) <= not((inputs(253)) and (inputs(71)));
    layer0_outputs(10224) <= inputs(152);
    layer0_outputs(10225) <= not((inputs(123)) and (inputs(119)));
    layer0_outputs(10226) <= inputs(74);
    layer0_outputs(10227) <= not(inputs(200));
    layer0_outputs(10228) <= (inputs(83)) xor (inputs(42));
    layer0_outputs(10229) <= not((inputs(28)) xor (inputs(213)));
    layer0_outputs(10230) <= inputs(59);
    layer0_outputs(10231) <= not(inputs(249)) or (inputs(206));
    layer0_outputs(10232) <= '1';
    layer0_outputs(10233) <= '1';
    layer0_outputs(10234) <= (inputs(174)) and not (inputs(238));
    layer0_outputs(10235) <= not(inputs(77)) or (inputs(212));
    layer0_outputs(10236) <= (inputs(51)) or (inputs(16));
    layer0_outputs(10237) <= not((inputs(180)) or (inputs(201)));
    layer0_outputs(10238) <= not(inputs(135)) or (inputs(67));
    layer0_outputs(10239) <= (inputs(60)) and not (inputs(108));
    layer1_outputs(0) <= not((layer0_outputs(10085)) or (layer0_outputs(4163)));
    layer1_outputs(1) <= not(layer0_outputs(263));
    layer1_outputs(2) <= layer0_outputs(3956);
    layer1_outputs(3) <= not(layer0_outputs(4563));
    layer1_outputs(4) <= layer0_outputs(632);
    layer1_outputs(5) <= (layer0_outputs(3570)) and (layer0_outputs(6804));
    layer1_outputs(6) <= (layer0_outputs(8299)) and (layer0_outputs(6828));
    layer1_outputs(7) <= layer0_outputs(7655);
    layer1_outputs(8) <= layer0_outputs(1006);
    layer1_outputs(9) <= (layer0_outputs(196)) and not (layer0_outputs(145));
    layer1_outputs(10) <= not((layer0_outputs(5935)) xor (layer0_outputs(5193)));
    layer1_outputs(11) <= (layer0_outputs(5923)) and not (layer0_outputs(1465));
    layer1_outputs(12) <= not((layer0_outputs(95)) or (layer0_outputs(9624)));
    layer1_outputs(13) <= (layer0_outputs(7320)) and not (layer0_outputs(1102));
    layer1_outputs(14) <= layer0_outputs(3686);
    layer1_outputs(15) <= not(layer0_outputs(6382));
    layer1_outputs(16) <= (layer0_outputs(4633)) and not (layer0_outputs(10200));
    layer1_outputs(17) <= not((layer0_outputs(1938)) or (layer0_outputs(9513)));
    layer1_outputs(18) <= '0';
    layer1_outputs(19) <= not((layer0_outputs(2913)) and (layer0_outputs(9137)));
    layer1_outputs(20) <= not(layer0_outputs(9905)) or (layer0_outputs(9772));
    layer1_outputs(21) <= '0';
    layer1_outputs(22) <= (layer0_outputs(6480)) or (layer0_outputs(8866));
    layer1_outputs(23) <= (layer0_outputs(2835)) and not (layer0_outputs(3934));
    layer1_outputs(24) <= not(layer0_outputs(5388)) or (layer0_outputs(4436));
    layer1_outputs(25) <= layer0_outputs(6161);
    layer1_outputs(26) <= not((layer0_outputs(5811)) or (layer0_outputs(6885)));
    layer1_outputs(27) <= not((layer0_outputs(345)) or (layer0_outputs(3449)));
    layer1_outputs(28) <= '0';
    layer1_outputs(29) <= (layer0_outputs(5460)) or (layer0_outputs(6009));
    layer1_outputs(30) <= (layer0_outputs(288)) and (layer0_outputs(10141));
    layer1_outputs(31) <= layer0_outputs(7860);
    layer1_outputs(32) <= not(layer0_outputs(5900));
    layer1_outputs(33) <= not(layer0_outputs(2822)) or (layer0_outputs(9009));
    layer1_outputs(34) <= '0';
    layer1_outputs(35) <= layer0_outputs(1006);
    layer1_outputs(36) <= not((layer0_outputs(7848)) or (layer0_outputs(1639)));
    layer1_outputs(37) <= not(layer0_outputs(7210)) or (layer0_outputs(8446));
    layer1_outputs(38) <= (layer0_outputs(6130)) or (layer0_outputs(5686));
    layer1_outputs(39) <= not((layer0_outputs(6256)) xor (layer0_outputs(8286)));
    layer1_outputs(40) <= not(layer0_outputs(8611));
    layer1_outputs(41) <= (layer0_outputs(2708)) and (layer0_outputs(3903));
    layer1_outputs(42) <= (layer0_outputs(2535)) and not (layer0_outputs(8699));
    layer1_outputs(43) <= (layer0_outputs(4752)) or (layer0_outputs(7689));
    layer1_outputs(44) <= (layer0_outputs(6356)) or (layer0_outputs(895));
    layer1_outputs(45) <= layer0_outputs(8393);
    layer1_outputs(46) <= not(layer0_outputs(3702));
    layer1_outputs(47) <= not(layer0_outputs(368));
    layer1_outputs(48) <= (layer0_outputs(2217)) and (layer0_outputs(1548));
    layer1_outputs(49) <= layer0_outputs(6529);
    layer1_outputs(50) <= not(layer0_outputs(7889));
    layer1_outputs(51) <= '0';
    layer1_outputs(52) <= '0';
    layer1_outputs(53) <= (layer0_outputs(3778)) and not (layer0_outputs(702));
    layer1_outputs(54) <= not(layer0_outputs(2308));
    layer1_outputs(55) <= not(layer0_outputs(9722));
    layer1_outputs(56) <= not(layer0_outputs(6557));
    layer1_outputs(57) <= (layer0_outputs(3005)) and (layer0_outputs(1915));
    layer1_outputs(58) <= (layer0_outputs(8573)) and (layer0_outputs(4627));
    layer1_outputs(59) <= layer0_outputs(4290);
    layer1_outputs(60) <= (layer0_outputs(7109)) or (layer0_outputs(9458));
    layer1_outputs(61) <= not(layer0_outputs(4354));
    layer1_outputs(62) <= '1';
    layer1_outputs(63) <= layer0_outputs(49);
    layer1_outputs(64) <= not((layer0_outputs(5547)) xor (layer0_outputs(1777)));
    layer1_outputs(65) <= layer0_outputs(6274);
    layer1_outputs(66) <= not((layer0_outputs(9520)) or (layer0_outputs(7950)));
    layer1_outputs(67) <= not((layer0_outputs(9191)) or (layer0_outputs(8076)));
    layer1_outputs(68) <= (layer0_outputs(475)) or (layer0_outputs(7397));
    layer1_outputs(69) <= not(layer0_outputs(382));
    layer1_outputs(70) <= (layer0_outputs(779)) or (layer0_outputs(4639));
    layer1_outputs(71) <= '1';
    layer1_outputs(72) <= (layer0_outputs(9318)) and not (layer0_outputs(722));
    layer1_outputs(73) <= not((layer0_outputs(6264)) and (layer0_outputs(6971)));
    layer1_outputs(74) <= not((layer0_outputs(7418)) xor (layer0_outputs(1131)));
    layer1_outputs(75) <= layer0_outputs(141);
    layer1_outputs(76) <= layer0_outputs(9665);
    layer1_outputs(77) <= (layer0_outputs(3279)) or (layer0_outputs(6984));
    layer1_outputs(78) <= (layer0_outputs(4481)) and (layer0_outputs(247));
    layer1_outputs(79) <= not((layer0_outputs(927)) and (layer0_outputs(10029)));
    layer1_outputs(80) <= (layer0_outputs(7008)) and not (layer0_outputs(1982));
    layer1_outputs(81) <= not(layer0_outputs(4109)) or (layer0_outputs(1575));
    layer1_outputs(82) <= not(layer0_outputs(7623));
    layer1_outputs(83) <= '1';
    layer1_outputs(84) <= layer0_outputs(1003);
    layer1_outputs(85) <= not((layer0_outputs(6276)) xor (layer0_outputs(6595)));
    layer1_outputs(86) <= not(layer0_outputs(6997)) or (layer0_outputs(1615));
    layer1_outputs(87) <= layer0_outputs(6805);
    layer1_outputs(88) <= not(layer0_outputs(5019));
    layer1_outputs(89) <= not(layer0_outputs(2580)) or (layer0_outputs(768));
    layer1_outputs(90) <= (layer0_outputs(7250)) and not (layer0_outputs(492));
    layer1_outputs(91) <= (layer0_outputs(3907)) and (layer0_outputs(4267));
    layer1_outputs(92) <= not(layer0_outputs(8885));
    layer1_outputs(93) <= not((layer0_outputs(7129)) or (layer0_outputs(1222)));
    layer1_outputs(94) <= not(layer0_outputs(6698));
    layer1_outputs(95) <= not((layer0_outputs(8179)) or (layer0_outputs(476)));
    layer1_outputs(96) <= not(layer0_outputs(9895)) or (layer0_outputs(3116));
    layer1_outputs(97) <= (layer0_outputs(3476)) xor (layer0_outputs(285));
    layer1_outputs(98) <= '0';
    layer1_outputs(99) <= not(layer0_outputs(5177));
    layer1_outputs(100) <= '1';
    layer1_outputs(101) <= not(layer0_outputs(830));
    layer1_outputs(102) <= not(layer0_outputs(2673));
    layer1_outputs(103) <= not(layer0_outputs(9190)) or (layer0_outputs(1039));
    layer1_outputs(104) <= not(layer0_outputs(3136));
    layer1_outputs(105) <= layer0_outputs(8563);
    layer1_outputs(106) <= layer0_outputs(5899);
    layer1_outputs(107) <= not(layer0_outputs(250)) or (layer0_outputs(4819));
    layer1_outputs(108) <= '1';
    layer1_outputs(109) <= (layer0_outputs(4146)) xor (layer0_outputs(8946));
    layer1_outputs(110) <= layer0_outputs(806);
    layer1_outputs(111) <= not(layer0_outputs(8219));
    layer1_outputs(112) <= not((layer0_outputs(6448)) and (layer0_outputs(9282)));
    layer1_outputs(113) <= not((layer0_outputs(2769)) and (layer0_outputs(5102)));
    layer1_outputs(114) <= layer0_outputs(9319);
    layer1_outputs(115) <= '1';
    layer1_outputs(116) <= not(layer0_outputs(7521)) or (layer0_outputs(7606));
    layer1_outputs(117) <= layer0_outputs(7367);
    layer1_outputs(118) <= layer0_outputs(4855);
    layer1_outputs(119) <= (layer0_outputs(6425)) and (layer0_outputs(8491));
    layer1_outputs(120) <= layer0_outputs(5464);
    layer1_outputs(121) <= layer0_outputs(7423);
    layer1_outputs(122) <= layer0_outputs(450);
    layer1_outputs(123) <= '0';
    layer1_outputs(124) <= (layer0_outputs(9183)) and not (layer0_outputs(3913));
    layer1_outputs(125) <= not((layer0_outputs(8587)) or (layer0_outputs(8576)));
    layer1_outputs(126) <= layer0_outputs(8543);
    layer1_outputs(127) <= not(layer0_outputs(6945));
    layer1_outputs(128) <= (layer0_outputs(9071)) or (layer0_outputs(9543));
    layer1_outputs(129) <= (layer0_outputs(2338)) and not (layer0_outputs(1031));
    layer1_outputs(130) <= not(layer0_outputs(6507));
    layer1_outputs(131) <= layer0_outputs(9160);
    layer1_outputs(132) <= not((layer0_outputs(4844)) and (layer0_outputs(7850)));
    layer1_outputs(133) <= layer0_outputs(3062);
    layer1_outputs(134) <= not(layer0_outputs(1334));
    layer1_outputs(135) <= (layer0_outputs(8164)) and not (layer0_outputs(5272));
    layer1_outputs(136) <= '0';
    layer1_outputs(137) <= not(layer0_outputs(5645));
    layer1_outputs(138) <= layer0_outputs(3114);
    layer1_outputs(139) <= '1';
    layer1_outputs(140) <= '0';
    layer1_outputs(141) <= not(layer0_outputs(5223));
    layer1_outputs(142) <= (layer0_outputs(6182)) and (layer0_outputs(9381));
    layer1_outputs(143) <= (layer0_outputs(2494)) or (layer0_outputs(5333));
    layer1_outputs(144) <= (layer0_outputs(5105)) and not (layer0_outputs(7091));
    layer1_outputs(145) <= (layer0_outputs(27)) and (layer0_outputs(3958));
    layer1_outputs(146) <= not(layer0_outputs(5718)) or (layer0_outputs(2287));
    layer1_outputs(147) <= '1';
    layer1_outputs(148) <= not(layer0_outputs(8099));
    layer1_outputs(149) <= not((layer0_outputs(3186)) xor (layer0_outputs(6069)));
    layer1_outputs(150) <= (layer0_outputs(9576)) and not (layer0_outputs(9711));
    layer1_outputs(151) <= not(layer0_outputs(9699)) or (layer0_outputs(8436));
    layer1_outputs(152) <= not(layer0_outputs(2792));
    layer1_outputs(153) <= not(layer0_outputs(9766)) or (layer0_outputs(9236));
    layer1_outputs(154) <= not(layer0_outputs(1620));
    layer1_outputs(155) <= (layer0_outputs(9392)) and not (layer0_outputs(7702));
    layer1_outputs(156) <= not(layer0_outputs(4220)) or (layer0_outputs(1036));
    layer1_outputs(157) <= (layer0_outputs(1460)) and not (layer0_outputs(814));
    layer1_outputs(158) <= layer0_outputs(6858);
    layer1_outputs(159) <= (layer0_outputs(6106)) and not (layer0_outputs(5316));
    layer1_outputs(160) <= (layer0_outputs(6256)) and not (layer0_outputs(8910));
    layer1_outputs(161) <= (layer0_outputs(8331)) and not (layer0_outputs(1114));
    layer1_outputs(162) <= (layer0_outputs(10213)) and not (layer0_outputs(8322));
    layer1_outputs(163) <= '1';
    layer1_outputs(164) <= '0';
    layer1_outputs(165) <= layer0_outputs(1233);
    layer1_outputs(166) <= not((layer0_outputs(80)) and (layer0_outputs(19)));
    layer1_outputs(167) <= not((layer0_outputs(5255)) and (layer0_outputs(8619)));
    layer1_outputs(168) <= not(layer0_outputs(4606)) or (layer0_outputs(7930));
    layer1_outputs(169) <= not(layer0_outputs(193));
    layer1_outputs(170) <= not((layer0_outputs(224)) xor (layer0_outputs(4440)));
    layer1_outputs(171) <= (layer0_outputs(669)) or (layer0_outputs(857));
    layer1_outputs(172) <= not(layer0_outputs(6162));
    layer1_outputs(173) <= layer0_outputs(4131);
    layer1_outputs(174) <= layer0_outputs(8087);
    layer1_outputs(175) <= layer0_outputs(10010);
    layer1_outputs(176) <= '0';
    layer1_outputs(177) <= '1';
    layer1_outputs(178) <= not(layer0_outputs(9476));
    layer1_outputs(179) <= layer0_outputs(8694);
    layer1_outputs(180) <= not(layer0_outputs(2393));
    layer1_outputs(181) <= (layer0_outputs(2480)) and not (layer0_outputs(3230));
    layer1_outputs(182) <= not(layer0_outputs(2706)) or (layer0_outputs(3633));
    layer1_outputs(183) <= not(layer0_outputs(10061)) or (layer0_outputs(8301));
    layer1_outputs(184) <= not(layer0_outputs(6226)) or (layer0_outputs(6191));
    layer1_outputs(185) <= not(layer0_outputs(7817));
    layer1_outputs(186) <= not(layer0_outputs(2664));
    layer1_outputs(187) <= not(layer0_outputs(5357));
    layer1_outputs(188) <= (layer0_outputs(8703)) and (layer0_outputs(9503));
    layer1_outputs(189) <= layer0_outputs(6736);
    layer1_outputs(190) <= (layer0_outputs(8355)) xor (layer0_outputs(9947));
    layer1_outputs(191) <= not((layer0_outputs(6464)) xor (layer0_outputs(5643)));
    layer1_outputs(192) <= (layer0_outputs(2185)) or (layer0_outputs(9202));
    layer1_outputs(193) <= '0';
    layer1_outputs(194) <= layer0_outputs(3148);
    layer1_outputs(195) <= not(layer0_outputs(8655));
    layer1_outputs(196) <= not(layer0_outputs(6297)) or (layer0_outputs(6657));
    layer1_outputs(197) <= not(layer0_outputs(7746));
    layer1_outputs(198) <= layer0_outputs(614);
    layer1_outputs(199) <= not((layer0_outputs(1557)) and (layer0_outputs(8291)));
    layer1_outputs(200) <= layer0_outputs(2150);
    layer1_outputs(201) <= not((layer0_outputs(10077)) or (layer0_outputs(6600)));
    layer1_outputs(202) <= (layer0_outputs(4859)) and not (layer0_outputs(5124));
    layer1_outputs(203) <= layer0_outputs(3626);
    layer1_outputs(204) <= (layer0_outputs(5110)) and not (layer0_outputs(8444));
    layer1_outputs(205) <= not((layer0_outputs(421)) and (layer0_outputs(9294)));
    layer1_outputs(206) <= not(layer0_outputs(4533));
    layer1_outputs(207) <= not(layer0_outputs(3780));
    layer1_outputs(208) <= not((layer0_outputs(4705)) or (layer0_outputs(2647)));
    layer1_outputs(209) <= (layer0_outputs(7973)) xor (layer0_outputs(7771));
    layer1_outputs(210) <= layer0_outputs(5595);
    layer1_outputs(211) <= not((layer0_outputs(9966)) xor (layer0_outputs(9937)));
    layer1_outputs(212) <= (layer0_outputs(4122)) or (layer0_outputs(1929));
    layer1_outputs(213) <= layer0_outputs(4009);
    layer1_outputs(214) <= not(layer0_outputs(3294));
    layer1_outputs(215) <= layer0_outputs(8852);
    layer1_outputs(216) <= (layer0_outputs(7928)) or (layer0_outputs(4409));
    layer1_outputs(217) <= not((layer0_outputs(2539)) and (layer0_outputs(7834)));
    layer1_outputs(218) <= not(layer0_outputs(685)) or (layer0_outputs(2212));
    layer1_outputs(219) <= not((layer0_outputs(7783)) or (layer0_outputs(4625)));
    layer1_outputs(220) <= not((layer0_outputs(3184)) xor (layer0_outputs(4743)));
    layer1_outputs(221) <= '1';
    layer1_outputs(222) <= layer0_outputs(185);
    layer1_outputs(223) <= not(layer0_outputs(8406)) or (layer0_outputs(8452));
    layer1_outputs(224) <= layer0_outputs(4995);
    layer1_outputs(225) <= layer0_outputs(8206);
    layer1_outputs(226) <= (layer0_outputs(9681)) and not (layer0_outputs(9309));
    layer1_outputs(227) <= (layer0_outputs(5239)) or (layer0_outputs(1157));
    layer1_outputs(228) <= (layer0_outputs(7878)) and not (layer0_outputs(2874));
    layer1_outputs(229) <= layer0_outputs(2004);
    layer1_outputs(230) <= '1';
    layer1_outputs(231) <= not((layer0_outputs(5796)) and (layer0_outputs(4491)));
    layer1_outputs(232) <= layer0_outputs(717);
    layer1_outputs(233) <= '1';
    layer1_outputs(234) <= (layer0_outputs(5937)) and not (layer0_outputs(5035));
    layer1_outputs(235) <= not(layer0_outputs(8095));
    layer1_outputs(236) <= layer0_outputs(4789);
    layer1_outputs(237) <= (layer0_outputs(4130)) or (layer0_outputs(6410));
    layer1_outputs(238) <= (layer0_outputs(3721)) and not (layer0_outputs(5150));
    layer1_outputs(239) <= (layer0_outputs(3391)) xor (layer0_outputs(3985));
    layer1_outputs(240) <= not(layer0_outputs(9658)) or (layer0_outputs(9606));
    layer1_outputs(241) <= not(layer0_outputs(4412));
    layer1_outputs(242) <= not((layer0_outputs(425)) and (layer0_outputs(1277)));
    layer1_outputs(243) <= (layer0_outputs(8233)) xor (layer0_outputs(9713));
    layer1_outputs(244) <= '0';
    layer1_outputs(245) <= layer0_outputs(1306);
    layer1_outputs(246) <= (layer0_outputs(2952)) xor (layer0_outputs(6814));
    layer1_outputs(247) <= not(layer0_outputs(4982)) or (layer0_outputs(8751));
    layer1_outputs(248) <= not(layer0_outputs(2178));
    layer1_outputs(249) <= layer0_outputs(6280);
    layer1_outputs(250) <= (layer0_outputs(4316)) and (layer0_outputs(9041));
    layer1_outputs(251) <= '1';
    layer1_outputs(252) <= not((layer0_outputs(6467)) or (layer0_outputs(1145)));
    layer1_outputs(253) <= not(layer0_outputs(2259)) or (layer0_outputs(8084));
    layer1_outputs(254) <= layer0_outputs(8047);
    layer1_outputs(255) <= (layer0_outputs(3558)) and not (layer0_outputs(5124));
    layer1_outputs(256) <= (layer0_outputs(5516)) xor (layer0_outputs(3391));
    layer1_outputs(257) <= not(layer0_outputs(5527));
    layer1_outputs(258) <= not(layer0_outputs(8442));
    layer1_outputs(259) <= layer0_outputs(2585);
    layer1_outputs(260) <= layer0_outputs(795);
    layer1_outputs(261) <= not(layer0_outputs(7541)) or (layer0_outputs(5944));
    layer1_outputs(262) <= '1';
    layer1_outputs(263) <= layer0_outputs(6527);
    layer1_outputs(264) <= (layer0_outputs(3608)) and not (layer0_outputs(3512));
    layer1_outputs(265) <= not(layer0_outputs(3067));
    layer1_outputs(266) <= not(layer0_outputs(3934));
    layer1_outputs(267) <= (layer0_outputs(7152)) and (layer0_outputs(8475));
    layer1_outputs(268) <= not(layer0_outputs(4403));
    layer1_outputs(269) <= layer0_outputs(1587);
    layer1_outputs(270) <= not(layer0_outputs(5192));
    layer1_outputs(271) <= '0';
    layer1_outputs(272) <= (layer0_outputs(8207)) and not (layer0_outputs(2700));
    layer1_outputs(273) <= not((layer0_outputs(9833)) xor (layer0_outputs(8715)));
    layer1_outputs(274) <= layer0_outputs(5921);
    layer1_outputs(275) <= layer0_outputs(5598);
    layer1_outputs(276) <= not(layer0_outputs(8666));
    layer1_outputs(277) <= (layer0_outputs(3155)) xor (layer0_outputs(9008));
    layer1_outputs(278) <= not(layer0_outputs(3846));
    layer1_outputs(279) <= not((layer0_outputs(6819)) and (layer0_outputs(2705)));
    layer1_outputs(280) <= not((layer0_outputs(9350)) and (layer0_outputs(2990)));
    layer1_outputs(281) <= not(layer0_outputs(8349));
    layer1_outputs(282) <= (layer0_outputs(989)) xor (layer0_outputs(8015));
    layer1_outputs(283) <= layer0_outputs(9320);
    layer1_outputs(284) <= not((layer0_outputs(3318)) or (layer0_outputs(245)));
    layer1_outputs(285) <= (layer0_outputs(2583)) and (layer0_outputs(3498));
    layer1_outputs(286) <= not((layer0_outputs(4192)) or (layer0_outputs(3346)));
    layer1_outputs(287) <= layer0_outputs(10097);
    layer1_outputs(288) <= layer0_outputs(8281);
    layer1_outputs(289) <= '1';
    layer1_outputs(290) <= (layer0_outputs(6014)) and not (layer0_outputs(9984));
    layer1_outputs(291) <= (layer0_outputs(1068)) and not (layer0_outputs(2868));
    layer1_outputs(292) <= '0';
    layer1_outputs(293) <= (layer0_outputs(2975)) and not (layer0_outputs(4616));
    layer1_outputs(294) <= not(layer0_outputs(7596)) or (layer0_outputs(5486));
    layer1_outputs(295) <= layer0_outputs(7997);
    layer1_outputs(296) <= (layer0_outputs(4776)) or (layer0_outputs(2904));
    layer1_outputs(297) <= (layer0_outputs(4852)) and (layer0_outputs(572));
    layer1_outputs(298) <= (layer0_outputs(8229)) and not (layer0_outputs(1142));
    layer1_outputs(299) <= not(layer0_outputs(5087));
    layer1_outputs(300) <= '1';
    layer1_outputs(301) <= not(layer0_outputs(135)) or (layer0_outputs(2334));
    layer1_outputs(302) <= not(layer0_outputs(3491)) or (layer0_outputs(5276));
    layer1_outputs(303) <= (layer0_outputs(6309)) or (layer0_outputs(6540));
    layer1_outputs(304) <= not(layer0_outputs(8790));
    layer1_outputs(305) <= layer0_outputs(4002);
    layer1_outputs(306) <= not(layer0_outputs(1350));
    layer1_outputs(307) <= (layer0_outputs(2716)) and (layer0_outputs(1595));
    layer1_outputs(308) <= (layer0_outputs(6534)) or (layer0_outputs(7872));
    layer1_outputs(309) <= (layer0_outputs(2575)) and (layer0_outputs(3794));
    layer1_outputs(310) <= '1';
    layer1_outputs(311) <= (layer0_outputs(4266)) or (layer0_outputs(8111));
    layer1_outputs(312) <= layer0_outputs(10194);
    layer1_outputs(313) <= not(layer0_outputs(1053)) or (layer0_outputs(2449));
    layer1_outputs(314) <= (layer0_outputs(9777)) and not (layer0_outputs(4360));
    layer1_outputs(315) <= (layer0_outputs(6841)) or (layer0_outputs(9807));
    layer1_outputs(316) <= (layer0_outputs(7192)) and not (layer0_outputs(4974));
    layer1_outputs(317) <= layer0_outputs(9915);
    layer1_outputs(318) <= (layer0_outputs(8725)) xor (layer0_outputs(4065));
    layer1_outputs(319) <= '1';
    layer1_outputs(320) <= layer0_outputs(6992);
    layer1_outputs(321) <= not(layer0_outputs(7457));
    layer1_outputs(322) <= not((layer0_outputs(5353)) and (layer0_outputs(6954)));
    layer1_outputs(323) <= (layer0_outputs(7134)) xor (layer0_outputs(5001));
    layer1_outputs(324) <= (layer0_outputs(5173)) and not (layer0_outputs(10177));
    layer1_outputs(325) <= not((layer0_outputs(7074)) and (layer0_outputs(8842)));
    layer1_outputs(326) <= not((layer0_outputs(7345)) or (layer0_outputs(5680)));
    layer1_outputs(327) <= (layer0_outputs(3986)) or (layer0_outputs(6820));
    layer1_outputs(328) <= (layer0_outputs(1868)) and not (layer0_outputs(6823));
    layer1_outputs(329) <= not(layer0_outputs(2945)) or (layer0_outputs(4182));
    layer1_outputs(330) <= not((layer0_outputs(7895)) and (layer0_outputs(9827)));
    layer1_outputs(331) <= (layer0_outputs(8494)) and not (layer0_outputs(341));
    layer1_outputs(332) <= not(layer0_outputs(1967));
    layer1_outputs(333) <= not(layer0_outputs(837)) or (layer0_outputs(4303));
    layer1_outputs(334) <= layer0_outputs(6908);
    layer1_outputs(335) <= not(layer0_outputs(10234));
    layer1_outputs(336) <= (layer0_outputs(2744)) and not (layer0_outputs(5903));
    layer1_outputs(337) <= '1';
    layer1_outputs(338) <= layer0_outputs(827);
    layer1_outputs(339) <= not(layer0_outputs(9072));
    layer1_outputs(340) <= not(layer0_outputs(4078));
    layer1_outputs(341) <= (layer0_outputs(1616)) and not (layer0_outputs(6932));
    layer1_outputs(342) <= layer0_outputs(5631);
    layer1_outputs(343) <= not(layer0_outputs(3915)) or (layer0_outputs(3103));
    layer1_outputs(344) <= layer0_outputs(5052);
    layer1_outputs(345) <= layer0_outputs(3855);
    layer1_outputs(346) <= layer0_outputs(2912);
    layer1_outputs(347) <= not(layer0_outputs(16)) or (layer0_outputs(6944));
    layer1_outputs(348) <= (layer0_outputs(7480)) and not (layer0_outputs(826));
    layer1_outputs(349) <= not((layer0_outputs(3970)) or (layer0_outputs(2838)));
    layer1_outputs(350) <= '0';
    layer1_outputs(351) <= not(layer0_outputs(6069));
    layer1_outputs(352) <= layer0_outputs(10093);
    layer1_outputs(353) <= (layer0_outputs(9032)) xor (layer0_outputs(8303));
    layer1_outputs(354) <= '0';
    layer1_outputs(355) <= not((layer0_outputs(1693)) or (layer0_outputs(4372)));
    layer1_outputs(356) <= not(layer0_outputs(4305));
    layer1_outputs(357) <= (layer0_outputs(9629)) and not (layer0_outputs(4087));
    layer1_outputs(358) <= (layer0_outputs(1893)) or (layer0_outputs(10032));
    layer1_outputs(359) <= not((layer0_outputs(8942)) xor (layer0_outputs(7628)));
    layer1_outputs(360) <= not(layer0_outputs(4080));
    layer1_outputs(361) <= not(layer0_outputs(9365)) or (layer0_outputs(9404));
    layer1_outputs(362) <= not(layer0_outputs(7219));
    layer1_outputs(363) <= (layer0_outputs(6870)) xor (layer0_outputs(6939));
    layer1_outputs(364) <= not(layer0_outputs(2972));
    layer1_outputs(365) <= not((layer0_outputs(2643)) and (layer0_outputs(3959)));
    layer1_outputs(366) <= not((layer0_outputs(4387)) or (layer0_outputs(1553)));
    layer1_outputs(367) <= not((layer0_outputs(6681)) and (layer0_outputs(9214)));
    layer1_outputs(368) <= layer0_outputs(2960);
    layer1_outputs(369) <= not((layer0_outputs(8473)) and (layer0_outputs(6198)));
    layer1_outputs(370) <= layer0_outputs(9546);
    layer1_outputs(371) <= (layer0_outputs(2995)) and not (layer0_outputs(7262));
    layer1_outputs(372) <= not(layer0_outputs(2040)) or (layer0_outputs(2458));
    layer1_outputs(373) <= layer0_outputs(5413);
    layer1_outputs(374) <= '0';
    layer1_outputs(375) <= not((layer0_outputs(6620)) or (layer0_outputs(1311)));
    layer1_outputs(376) <= not(layer0_outputs(8776)) or (layer0_outputs(899));
    layer1_outputs(377) <= layer0_outputs(7346);
    layer1_outputs(378) <= (layer0_outputs(7052)) and not (layer0_outputs(8795));
    layer1_outputs(379) <= not((layer0_outputs(7788)) and (layer0_outputs(9721)));
    layer1_outputs(380) <= not(layer0_outputs(1315)) or (layer0_outputs(1053));
    layer1_outputs(381) <= not(layer0_outputs(6538));
    layer1_outputs(382) <= not((layer0_outputs(1419)) or (layer0_outputs(7233)));
    layer1_outputs(383) <= not(layer0_outputs(104)) or (layer0_outputs(2898));
    layer1_outputs(384) <= layer0_outputs(9065);
    layer1_outputs(385) <= not(layer0_outputs(2548)) or (layer0_outputs(9998));
    layer1_outputs(386) <= not((layer0_outputs(6546)) and (layer0_outputs(5730)));
    layer1_outputs(387) <= layer0_outputs(6071);
    layer1_outputs(388) <= not(layer0_outputs(2309));
    layer1_outputs(389) <= (layer0_outputs(709)) and (layer0_outputs(5991));
    layer1_outputs(390) <= not(layer0_outputs(7396));
    layer1_outputs(391) <= not(layer0_outputs(4606));
    layer1_outputs(392) <= (layer0_outputs(10131)) and not (layer0_outputs(7686));
    layer1_outputs(393) <= not((layer0_outputs(6259)) or (layer0_outputs(5255)));
    layer1_outputs(394) <= not((layer0_outputs(2574)) and (layer0_outputs(2614)));
    layer1_outputs(395) <= (layer0_outputs(3703)) and not (layer0_outputs(5209));
    layer1_outputs(396) <= layer0_outputs(4434);
    layer1_outputs(397) <= layer0_outputs(5762);
    layer1_outputs(398) <= not(layer0_outputs(10027));
    layer1_outputs(399) <= not(layer0_outputs(1240));
    layer1_outputs(400) <= not((layer0_outputs(6847)) and (layer0_outputs(9593)));
    layer1_outputs(401) <= layer0_outputs(5368);
    layer1_outputs(402) <= not(layer0_outputs(5546)) or (layer0_outputs(7121));
    layer1_outputs(403) <= (layer0_outputs(3006)) xor (layer0_outputs(3657));
    layer1_outputs(404) <= '0';
    layer1_outputs(405) <= (layer0_outputs(2042)) and (layer0_outputs(605));
    layer1_outputs(406) <= '0';
    layer1_outputs(407) <= (layer0_outputs(3164)) xor (layer0_outputs(9686));
    layer1_outputs(408) <= not(layer0_outputs(8090)) or (layer0_outputs(7621));
    layer1_outputs(409) <= '1';
    layer1_outputs(410) <= not(layer0_outputs(6975));
    layer1_outputs(411) <= not(layer0_outputs(2700)) or (layer0_outputs(9586));
    layer1_outputs(412) <= (layer0_outputs(5715)) and not (layer0_outputs(8225));
    layer1_outputs(413) <= (layer0_outputs(7995)) and (layer0_outputs(8959));
    layer1_outputs(414) <= (layer0_outputs(3124)) and not (layer0_outputs(9177));
    layer1_outputs(415) <= '0';
    layer1_outputs(416) <= (layer0_outputs(9727)) and not (layer0_outputs(5350));
    layer1_outputs(417) <= not(layer0_outputs(1508));
    layer1_outputs(418) <= not((layer0_outputs(4383)) or (layer0_outputs(8168)));
    layer1_outputs(419) <= not(layer0_outputs(9552));
    layer1_outputs(420) <= layer0_outputs(2976);
    layer1_outputs(421) <= not(layer0_outputs(10185));
    layer1_outputs(422) <= not((layer0_outputs(2508)) or (layer0_outputs(7433)));
    layer1_outputs(423) <= not((layer0_outputs(3641)) and (layer0_outputs(877)));
    layer1_outputs(424) <= not((layer0_outputs(6537)) or (layer0_outputs(8196)));
    layer1_outputs(425) <= not(layer0_outputs(3807)) or (layer0_outputs(8726));
    layer1_outputs(426) <= not(layer0_outputs(8297));
    layer1_outputs(427) <= not(layer0_outputs(6512)) or (layer0_outputs(4118));
    layer1_outputs(428) <= not(layer0_outputs(1828));
    layer1_outputs(429) <= (layer0_outputs(3128)) or (layer0_outputs(3729));
    layer1_outputs(430) <= (layer0_outputs(8300)) and (layer0_outputs(7897));
    layer1_outputs(431) <= not(layer0_outputs(5577)) or (layer0_outputs(7503));
    layer1_outputs(432) <= not(layer0_outputs(6104));
    layer1_outputs(433) <= not(layer0_outputs(5072));
    layer1_outputs(434) <= not(layer0_outputs(5659));
    layer1_outputs(435) <= not(layer0_outputs(6277));
    layer1_outputs(436) <= layer0_outputs(3693);
    layer1_outputs(437) <= '0';
    layer1_outputs(438) <= '1';
    layer1_outputs(439) <= not(layer0_outputs(9436)) or (layer0_outputs(365));
    layer1_outputs(440) <= (layer0_outputs(8691)) or (layer0_outputs(9231));
    layer1_outputs(441) <= layer0_outputs(8927);
    layer1_outputs(442) <= '0';
    layer1_outputs(443) <= '0';
    layer1_outputs(444) <= (layer0_outputs(7481)) and (layer0_outputs(8287));
    layer1_outputs(445) <= not(layer0_outputs(1315)) or (layer0_outputs(9028));
    layer1_outputs(446) <= not(layer0_outputs(6334));
    layer1_outputs(447) <= '0';
    layer1_outputs(448) <= not(layer0_outputs(9614));
    layer1_outputs(449) <= not(layer0_outputs(4327)) or (layer0_outputs(4700));
    layer1_outputs(450) <= (layer0_outputs(2151)) and not (layer0_outputs(5543));
    layer1_outputs(451) <= '1';
    layer1_outputs(452) <= not((layer0_outputs(5971)) and (layer0_outputs(4994)));
    layer1_outputs(453) <= (layer0_outputs(7114)) and not (layer0_outputs(2287));
    layer1_outputs(454) <= not(layer0_outputs(8440)) or (layer0_outputs(9886));
    layer1_outputs(455) <= layer0_outputs(1197);
    layer1_outputs(456) <= layer0_outputs(7299);
    layer1_outputs(457) <= not(layer0_outputs(645));
    layer1_outputs(458) <= '1';
    layer1_outputs(459) <= (layer0_outputs(1149)) or (layer0_outputs(4341));
    layer1_outputs(460) <= (layer0_outputs(8417)) and not (layer0_outputs(1063));
    layer1_outputs(461) <= (layer0_outputs(4366)) and not (layer0_outputs(4553));
    layer1_outputs(462) <= not(layer0_outputs(7858)) or (layer0_outputs(10021));
    layer1_outputs(463) <= (layer0_outputs(8006)) and not (layer0_outputs(1533));
    layer1_outputs(464) <= not(layer0_outputs(9617));
    layer1_outputs(465) <= not((layer0_outputs(4990)) and (layer0_outputs(3280)));
    layer1_outputs(466) <= not(layer0_outputs(6023)) or (layer0_outputs(6451));
    layer1_outputs(467) <= '1';
    layer1_outputs(468) <= not((layer0_outputs(3672)) and (layer0_outputs(2028)));
    layer1_outputs(469) <= not(layer0_outputs(2055));
    layer1_outputs(470) <= not(layer0_outputs(6631));
    layer1_outputs(471) <= layer0_outputs(2955);
    layer1_outputs(472) <= (layer0_outputs(8550)) and not (layer0_outputs(5626));
    layer1_outputs(473) <= not((layer0_outputs(7153)) or (layer0_outputs(5895)));
    layer1_outputs(474) <= '0';
    layer1_outputs(475) <= not(layer0_outputs(1722));
    layer1_outputs(476) <= not(layer0_outputs(1015)) or (layer0_outputs(7562));
    layer1_outputs(477) <= layer0_outputs(5649);
    layer1_outputs(478) <= not((layer0_outputs(6854)) xor (layer0_outputs(9087)));
    layer1_outputs(479) <= not((layer0_outputs(3067)) and (layer0_outputs(751)));
    layer1_outputs(480) <= not(layer0_outputs(7156)) or (layer0_outputs(6915));
    layer1_outputs(481) <= not(layer0_outputs(2473));
    layer1_outputs(482) <= (layer0_outputs(8390)) and not (layer0_outputs(781));
    layer1_outputs(483) <= not(layer0_outputs(1499)) or (layer0_outputs(7076));
    layer1_outputs(484) <= not(layer0_outputs(4200));
    layer1_outputs(485) <= (layer0_outputs(9674)) or (layer0_outputs(7025));
    layer1_outputs(486) <= not((layer0_outputs(2443)) or (layer0_outputs(10075)));
    layer1_outputs(487) <= not(layer0_outputs(8373)) or (layer0_outputs(8429));
    layer1_outputs(488) <= layer0_outputs(7117);
    layer1_outputs(489) <= (layer0_outputs(10092)) and (layer0_outputs(2591));
    layer1_outputs(490) <= not((layer0_outputs(9903)) xor (layer0_outputs(4879)));
    layer1_outputs(491) <= (layer0_outputs(9167)) or (layer0_outputs(1277));
    layer1_outputs(492) <= not(layer0_outputs(309)) or (layer0_outputs(240));
    layer1_outputs(493) <= '1';
    layer1_outputs(494) <= not((layer0_outputs(2106)) and (layer0_outputs(7527)));
    layer1_outputs(495) <= layer0_outputs(9341);
    layer1_outputs(496) <= (layer0_outputs(186)) and not (layer0_outputs(9144));
    layer1_outputs(497) <= (layer0_outputs(2146)) or (layer0_outputs(10178));
    layer1_outputs(498) <= '0';
    layer1_outputs(499) <= not(layer0_outputs(1756));
    layer1_outputs(500) <= not(layer0_outputs(3762)) or (layer0_outputs(3689));
    layer1_outputs(501) <= (layer0_outputs(5552)) and (layer0_outputs(4008));
    layer1_outputs(502) <= layer0_outputs(4245);
    layer1_outputs(503) <= (layer0_outputs(7172)) and not (layer0_outputs(7610));
    layer1_outputs(504) <= layer0_outputs(6652);
    layer1_outputs(505) <= not(layer0_outputs(4003));
    layer1_outputs(506) <= (layer0_outputs(664)) and (layer0_outputs(1425));
    layer1_outputs(507) <= not((layer0_outputs(8760)) and (layer0_outputs(2303)));
    layer1_outputs(508) <= (layer0_outputs(5903)) and not (layer0_outputs(9845));
    layer1_outputs(509) <= '1';
    layer1_outputs(510) <= layer0_outputs(652);
    layer1_outputs(511) <= not(layer0_outputs(8447));
    layer1_outputs(512) <= (layer0_outputs(7776)) xor (layer0_outputs(4726));
    layer1_outputs(513) <= layer0_outputs(1308);
    layer1_outputs(514) <= not(layer0_outputs(2444)) or (layer0_outputs(9848));
    layer1_outputs(515) <= (layer0_outputs(7805)) and not (layer0_outputs(7855));
    layer1_outputs(516) <= (layer0_outputs(6520)) and (layer0_outputs(3439));
    layer1_outputs(517) <= (layer0_outputs(9207)) and not (layer0_outputs(2758));
    layer1_outputs(518) <= (layer0_outputs(9964)) or (layer0_outputs(7277));
    layer1_outputs(519) <= (layer0_outputs(8892)) and not (layer0_outputs(7462));
    layer1_outputs(520) <= not(layer0_outputs(7844));
    layer1_outputs(521) <= '0';
    layer1_outputs(522) <= not(layer0_outputs(1910));
    layer1_outputs(523) <= not(layer0_outputs(1136));
    layer1_outputs(524) <= (layer0_outputs(2131)) and not (layer0_outputs(4296));
    layer1_outputs(525) <= not((layer0_outputs(10138)) xor (layer0_outputs(6300)));
    layer1_outputs(526) <= (layer0_outputs(9823)) and not (layer0_outputs(7040));
    layer1_outputs(527) <= not(layer0_outputs(4377)) or (layer0_outputs(9014));
    layer1_outputs(528) <= not(layer0_outputs(8177)) or (layer0_outputs(6352));
    layer1_outputs(529) <= not(layer0_outputs(1408));
    layer1_outputs(530) <= not(layer0_outputs(990)) or (layer0_outputs(5297));
    layer1_outputs(531) <= not(layer0_outputs(7175)) or (layer0_outputs(8391));
    layer1_outputs(532) <= (layer0_outputs(6196)) and not (layer0_outputs(5074));
    layer1_outputs(533) <= not(layer0_outputs(8093));
    layer1_outputs(534) <= not((layer0_outputs(115)) or (layer0_outputs(7268)));
    layer1_outputs(535) <= not(layer0_outputs(7589)) or (layer0_outputs(6594));
    layer1_outputs(536) <= layer0_outputs(3441);
    layer1_outputs(537) <= (layer0_outputs(733)) and not (layer0_outputs(9094));
    layer1_outputs(538) <= (layer0_outputs(5096)) or (layer0_outputs(2263));
    layer1_outputs(539) <= (layer0_outputs(207)) and not (layer0_outputs(7622));
    layer1_outputs(540) <= (layer0_outputs(4219)) and not (layer0_outputs(3106));
    layer1_outputs(541) <= (layer0_outputs(8824)) and not (layer0_outputs(5699));
    layer1_outputs(542) <= layer0_outputs(3802);
    layer1_outputs(543) <= '1';
    layer1_outputs(544) <= not(layer0_outputs(161));
    layer1_outputs(545) <= not((layer0_outputs(6034)) xor (layer0_outputs(8698)));
    layer1_outputs(546) <= not((layer0_outputs(214)) and (layer0_outputs(176)));
    layer1_outputs(547) <= layer0_outputs(8422);
    layer1_outputs(548) <= '1';
    layer1_outputs(549) <= not(layer0_outputs(3910));
    layer1_outputs(550) <= layer0_outputs(5524);
    layer1_outputs(551) <= not(layer0_outputs(7428)) or (layer0_outputs(5654));
    layer1_outputs(552) <= not((layer0_outputs(7324)) or (layer0_outputs(8973)));
    layer1_outputs(553) <= not(layer0_outputs(3559)) or (layer0_outputs(108));
    layer1_outputs(554) <= not(layer0_outputs(1982));
    layer1_outputs(555) <= layer0_outputs(9491);
    layer1_outputs(556) <= layer0_outputs(7147);
    layer1_outputs(557) <= not(layer0_outputs(568));
    layer1_outputs(558) <= (layer0_outputs(5491)) and not (layer0_outputs(1924));
    layer1_outputs(559) <= not(layer0_outputs(7190)) or (layer0_outputs(5677));
    layer1_outputs(560) <= not(layer0_outputs(268)) or (layer0_outputs(8914));
    layer1_outputs(561) <= layer0_outputs(4828);
    layer1_outputs(562) <= not(layer0_outputs(5507)) or (layer0_outputs(6697));
    layer1_outputs(563) <= (layer0_outputs(1418)) and (layer0_outputs(2447));
    layer1_outputs(564) <= not((layer0_outputs(5485)) or (layer0_outputs(5739)));
    layer1_outputs(565) <= not(layer0_outputs(10140)) or (layer0_outputs(1736));
    layer1_outputs(566) <= not(layer0_outputs(298)) or (layer0_outputs(247));
    layer1_outputs(567) <= layer0_outputs(8615);
    layer1_outputs(568) <= layer0_outputs(7228);
    layer1_outputs(569) <= (layer0_outputs(5879)) and (layer0_outputs(6309));
    layer1_outputs(570) <= not(layer0_outputs(8606)) or (layer0_outputs(2184));
    layer1_outputs(571) <= not(layer0_outputs(9653));
    layer1_outputs(572) <= not((layer0_outputs(10150)) and (layer0_outputs(9094)));
    layer1_outputs(573) <= not(layer0_outputs(1160));
    layer1_outputs(574) <= (layer0_outputs(5164)) and not (layer0_outputs(3528));
    layer1_outputs(575) <= '0';
    layer1_outputs(576) <= (layer0_outputs(1930)) and not (layer0_outputs(3405));
    layer1_outputs(577) <= layer0_outputs(6755);
    layer1_outputs(578) <= not(layer0_outputs(6661)) or (layer0_outputs(3546));
    layer1_outputs(579) <= not(layer0_outputs(821));
    layer1_outputs(580) <= (layer0_outputs(5515)) and not (layer0_outputs(3893));
    layer1_outputs(581) <= not(layer0_outputs(4430));
    layer1_outputs(582) <= layer0_outputs(4761);
    layer1_outputs(583) <= not(layer0_outputs(5912)) or (layer0_outputs(8629));
    layer1_outputs(584) <= (layer0_outputs(533)) and not (layer0_outputs(5818));
    layer1_outputs(585) <= not(layer0_outputs(8810));
    layer1_outputs(586) <= not((layer0_outputs(719)) xor (layer0_outputs(3441)));
    layer1_outputs(587) <= layer0_outputs(3439);
    layer1_outputs(588) <= (layer0_outputs(3181)) and not (layer0_outputs(4033));
    layer1_outputs(589) <= not(layer0_outputs(4105));
    layer1_outputs(590) <= not((layer0_outputs(9634)) or (layer0_outputs(3328)));
    layer1_outputs(591) <= not(layer0_outputs(6881)) or (layer0_outputs(1078));
    layer1_outputs(592) <= not((layer0_outputs(9964)) or (layer0_outputs(8788)));
    layer1_outputs(593) <= not((layer0_outputs(5825)) and (layer0_outputs(5063)));
    layer1_outputs(594) <= '1';
    layer1_outputs(595) <= not(layer0_outputs(866)) or (layer0_outputs(8090));
    layer1_outputs(596) <= not(layer0_outputs(4826)) or (layer0_outputs(7725));
    layer1_outputs(597) <= layer0_outputs(8211);
    layer1_outputs(598) <= (layer0_outputs(5659)) and (layer0_outputs(8041));
    layer1_outputs(599) <= '0';
    layer1_outputs(600) <= layer0_outputs(7139);
    layer1_outputs(601) <= not((layer0_outputs(4740)) and (layer0_outputs(582)));
    layer1_outputs(602) <= (layer0_outputs(8756)) and (layer0_outputs(1530));
    layer1_outputs(603) <= not(layer0_outputs(1913));
    layer1_outputs(604) <= (layer0_outputs(9685)) or (layer0_outputs(9280));
    layer1_outputs(605) <= '1';
    layer1_outputs(606) <= layer0_outputs(4878);
    layer1_outputs(607) <= (layer0_outputs(1723)) or (layer0_outputs(2254));
    layer1_outputs(608) <= layer0_outputs(289);
    layer1_outputs(609) <= '0';
    layer1_outputs(610) <= (layer0_outputs(643)) or (layer0_outputs(1519));
    layer1_outputs(611) <= layer0_outputs(4073);
    layer1_outputs(612) <= not(layer0_outputs(2680)) or (layer0_outputs(5955));
    layer1_outputs(613) <= not((layer0_outputs(1569)) or (layer0_outputs(8398)));
    layer1_outputs(614) <= (layer0_outputs(139)) and not (layer0_outputs(8271));
    layer1_outputs(615) <= (layer0_outputs(1797)) or (layer0_outputs(3760));
    layer1_outputs(616) <= (layer0_outputs(4397)) and not (layer0_outputs(7136));
    layer1_outputs(617) <= '1';
    layer1_outputs(618) <= not(layer0_outputs(1095)) or (layer0_outputs(4084));
    layer1_outputs(619) <= not(layer0_outputs(1323));
    layer1_outputs(620) <= not(layer0_outputs(1365)) or (layer0_outputs(9930));
    layer1_outputs(621) <= (layer0_outputs(9757)) and not (layer0_outputs(5727));
    layer1_outputs(622) <= not(layer0_outputs(9673));
    layer1_outputs(623) <= not(layer0_outputs(4950)) or (layer0_outputs(9229));
    layer1_outputs(624) <= layer0_outputs(5141);
    layer1_outputs(625) <= not(layer0_outputs(9384));
    layer1_outputs(626) <= not(layer0_outputs(5858)) or (layer0_outputs(1241));
    layer1_outputs(627) <= not((layer0_outputs(2370)) and (layer0_outputs(5155)));
    layer1_outputs(628) <= (layer0_outputs(5911)) and not (layer0_outputs(5826));
    layer1_outputs(629) <= (layer0_outputs(3661)) or (layer0_outputs(10137));
    layer1_outputs(630) <= (layer0_outputs(6448)) or (layer0_outputs(8795));
    layer1_outputs(631) <= '0';
    layer1_outputs(632) <= (layer0_outputs(7510)) and not (layer0_outputs(7354));
    layer1_outputs(633) <= not((layer0_outputs(4722)) xor (layer0_outputs(6584)));
    layer1_outputs(634) <= layer0_outputs(9663);
    layer1_outputs(635) <= not(layer0_outputs(9051));
    layer1_outputs(636) <= not(layer0_outputs(853));
    layer1_outputs(637) <= not(layer0_outputs(2739)) or (layer0_outputs(9870));
    layer1_outputs(638) <= '1';
    layer1_outputs(639) <= not(layer0_outputs(1558)) or (layer0_outputs(5745));
    layer1_outputs(640) <= not((layer0_outputs(2174)) and (layer0_outputs(7042)));
    layer1_outputs(641) <= not((layer0_outputs(8019)) xor (layer0_outputs(6230)));
    layer1_outputs(642) <= '0';
    layer1_outputs(643) <= layer0_outputs(5754);
    layer1_outputs(644) <= (layer0_outputs(158)) or (layer0_outputs(2640));
    layer1_outputs(645) <= not((layer0_outputs(10118)) xor (layer0_outputs(3537)));
    layer1_outputs(646) <= '0';
    layer1_outputs(647) <= (layer0_outputs(9482)) xor (layer0_outputs(4465));
    layer1_outputs(648) <= not((layer0_outputs(5458)) and (layer0_outputs(2394)));
    layer1_outputs(649) <= not(layer0_outputs(7849));
    layer1_outputs(650) <= layer0_outputs(749);
    layer1_outputs(651) <= (layer0_outputs(5175)) or (layer0_outputs(5398));
    layer1_outputs(652) <= (layer0_outputs(7)) or (layer0_outputs(4771));
    layer1_outputs(653) <= not(layer0_outputs(1874)) or (layer0_outputs(6148));
    layer1_outputs(654) <= (layer0_outputs(6654)) and not (layer0_outputs(4289));
    layer1_outputs(655) <= layer0_outputs(4258);
    layer1_outputs(656) <= not(layer0_outputs(3471));
    layer1_outputs(657) <= not(layer0_outputs(650));
    layer1_outputs(658) <= layer0_outputs(3687);
    layer1_outputs(659) <= not((layer0_outputs(4273)) xor (layer0_outputs(7056)));
    layer1_outputs(660) <= not((layer0_outputs(7577)) or (layer0_outputs(9572)));
    layer1_outputs(661) <= not(layer0_outputs(8348)) or (layer0_outputs(70));
    layer1_outputs(662) <= layer0_outputs(2000);
    layer1_outputs(663) <= not((layer0_outputs(2252)) xor (layer0_outputs(8911)));
    layer1_outputs(664) <= (layer0_outputs(416)) and (layer0_outputs(6577));
    layer1_outputs(665) <= layer0_outputs(7140);
    layer1_outputs(666) <= layer0_outputs(3601);
    layer1_outputs(667) <= not(layer0_outputs(192));
    layer1_outputs(668) <= layer0_outputs(1245);
    layer1_outputs(669) <= not(layer0_outputs(8132));
    layer1_outputs(670) <= not(layer0_outputs(2639));
    layer1_outputs(671) <= (layer0_outputs(7071)) xor (layer0_outputs(1295));
    layer1_outputs(672) <= (layer0_outputs(9860)) and (layer0_outputs(5182));
    layer1_outputs(673) <= not((layer0_outputs(3511)) and (layer0_outputs(7359)));
    layer1_outputs(674) <= (layer0_outputs(4972)) and not (layer0_outputs(6569));
    layer1_outputs(675) <= (layer0_outputs(6791)) and not (layer0_outputs(10071));
    layer1_outputs(676) <= (layer0_outputs(4274)) or (layer0_outputs(6517));
    layer1_outputs(677) <= (layer0_outputs(4542)) and not (layer0_outputs(8426));
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= layer0_outputs(2426);
    layer1_outputs(680) <= not(layer0_outputs(4362));
    layer1_outputs(681) <= not(layer0_outputs(6871));
    layer1_outputs(682) <= '1';
    layer1_outputs(683) <= not((layer0_outputs(9347)) and (layer0_outputs(5833)));
    layer1_outputs(684) <= (layer0_outputs(1287)) and not (layer0_outputs(7452));
    layer1_outputs(685) <= '0';
    layer1_outputs(686) <= (layer0_outputs(9751)) xor (layer0_outputs(6848));
    layer1_outputs(687) <= '0';
    layer1_outputs(688) <= (layer0_outputs(6878)) and not (layer0_outputs(1532));
    layer1_outputs(689) <= (layer0_outputs(1685)) and not (layer0_outputs(8453));
    layer1_outputs(690) <= layer0_outputs(7561);
    layer1_outputs(691) <= not((layer0_outputs(869)) xor (layer0_outputs(5507)));
    layer1_outputs(692) <= not((layer0_outputs(890)) or (layer0_outputs(9002)));
    layer1_outputs(693) <= layer0_outputs(5603);
    layer1_outputs(694) <= layer0_outputs(4474);
    layer1_outputs(695) <= (layer0_outputs(8379)) or (layer0_outputs(671));
    layer1_outputs(696) <= not((layer0_outputs(500)) xor (layer0_outputs(5752)));
    layer1_outputs(697) <= (layer0_outputs(1631)) and not (layer0_outputs(1225));
    layer1_outputs(698) <= not(layer0_outputs(9615));
    layer1_outputs(699) <= (layer0_outputs(6779)) and not (layer0_outputs(1900));
    layer1_outputs(700) <= (layer0_outputs(6002)) and not (layer0_outputs(9447));
    layer1_outputs(701) <= not(layer0_outputs(8778));
    layer1_outputs(702) <= not((layer0_outputs(3196)) or (layer0_outputs(9522)));
    layer1_outputs(703) <= (layer0_outputs(8762)) and (layer0_outputs(5826));
    layer1_outputs(704) <= not((layer0_outputs(9157)) xor (layer0_outputs(1560)));
    layer1_outputs(705) <= not((layer0_outputs(4962)) xor (layer0_outputs(1288)));
    layer1_outputs(706) <= '1';
    layer1_outputs(707) <= layer0_outputs(7757);
    layer1_outputs(708) <= not(layer0_outputs(3594));
    layer1_outputs(709) <= not(layer0_outputs(48));
    layer1_outputs(710) <= not(layer0_outputs(3717)) or (layer0_outputs(3317));
    layer1_outputs(711) <= layer0_outputs(6067);
    layer1_outputs(712) <= not((layer0_outputs(7200)) or (layer0_outputs(2504)));
    layer1_outputs(713) <= (layer0_outputs(6093)) and not (layer0_outputs(9275));
    layer1_outputs(714) <= not((layer0_outputs(9765)) or (layer0_outputs(7304)));
    layer1_outputs(715) <= '1';
    layer1_outputs(716) <= layer0_outputs(5591);
    layer1_outputs(717) <= not(layer0_outputs(5527)) or (layer0_outputs(3378));
    layer1_outputs(718) <= '1';
    layer1_outputs(719) <= not((layer0_outputs(862)) and (layer0_outputs(663)));
    layer1_outputs(720) <= layer0_outputs(867);
    layer1_outputs(721) <= not(layer0_outputs(261));
    layer1_outputs(722) <= (layer0_outputs(7730)) and not (layer0_outputs(9378));
    layer1_outputs(723) <= not((layer0_outputs(4672)) xor (layer0_outputs(9095)));
    layer1_outputs(724) <= not(layer0_outputs(7401)) or (layer0_outputs(9762));
    layer1_outputs(725) <= not(layer0_outputs(1351));
    layer1_outputs(726) <= (layer0_outputs(1685)) xor (layer0_outputs(6996));
    layer1_outputs(727) <= '1';
    layer1_outputs(728) <= not(layer0_outputs(8381));
    layer1_outputs(729) <= not(layer0_outputs(1807)) or (layer0_outputs(9703));
    layer1_outputs(730) <= (layer0_outputs(7793)) and not (layer0_outputs(6551));
    layer1_outputs(731) <= layer0_outputs(5562);
    layer1_outputs(732) <= not((layer0_outputs(9946)) and (layer0_outputs(367)));
    layer1_outputs(733) <= (layer0_outputs(2167)) or (layer0_outputs(1669));
    layer1_outputs(734) <= layer0_outputs(2812);
    layer1_outputs(735) <= not(layer0_outputs(4027));
    layer1_outputs(736) <= '0';
    layer1_outputs(737) <= (layer0_outputs(3004)) and (layer0_outputs(6192));
    layer1_outputs(738) <= (layer0_outputs(2172)) and (layer0_outputs(7678));
    layer1_outputs(739) <= not(layer0_outputs(8145));
    layer1_outputs(740) <= not((layer0_outputs(2332)) or (layer0_outputs(3148)));
    layer1_outputs(741) <= not(layer0_outputs(6910));
    layer1_outputs(742) <= (layer0_outputs(6184)) or (layer0_outputs(4999));
    layer1_outputs(743) <= not(layer0_outputs(8622));
    layer1_outputs(744) <= layer0_outputs(1748);
    layer1_outputs(745) <= (layer0_outputs(5517)) and not (layer0_outputs(1403));
    layer1_outputs(746) <= (layer0_outputs(2241)) and not (layer0_outputs(3654));
    layer1_outputs(747) <= not(layer0_outputs(7859));
    layer1_outputs(748) <= '0';
    layer1_outputs(749) <= not((layer0_outputs(3373)) and (layer0_outputs(5882)));
    layer1_outputs(750) <= not(layer0_outputs(2743));
    layer1_outputs(751) <= not(layer0_outputs(2411));
    layer1_outputs(752) <= layer0_outputs(8704);
    layer1_outputs(753) <= not(layer0_outputs(3921));
    layer1_outputs(754) <= layer0_outputs(8515);
    layer1_outputs(755) <= not(layer0_outputs(2291));
    layer1_outputs(756) <= (layer0_outputs(1674)) xor (layer0_outputs(6408));
    layer1_outputs(757) <= not(layer0_outputs(9569)) or (layer0_outputs(9695));
    layer1_outputs(758) <= (layer0_outputs(8199)) or (layer0_outputs(2616));
    layer1_outputs(759) <= not(layer0_outputs(8664));
    layer1_outputs(760) <= (layer0_outputs(5708)) xor (layer0_outputs(1900));
    layer1_outputs(761) <= layer0_outputs(9793);
    layer1_outputs(762) <= not(layer0_outputs(4089)) or (layer0_outputs(1618));
    layer1_outputs(763) <= not((layer0_outputs(4643)) and (layer0_outputs(6288)));
    layer1_outputs(764) <= layer0_outputs(9748);
    layer1_outputs(765) <= (layer0_outputs(9216)) or (layer0_outputs(6368));
    layer1_outputs(766) <= '1';
    layer1_outputs(767) <= layer0_outputs(696);
    layer1_outputs(768) <= '0';
    layer1_outputs(769) <= (layer0_outputs(1387)) and not (layer0_outputs(3811));
    layer1_outputs(770) <= layer0_outputs(6750);
    layer1_outputs(771) <= (layer0_outputs(6478)) and (layer0_outputs(468));
    layer1_outputs(772) <= '1';
    layer1_outputs(773) <= not((layer0_outputs(17)) and (layer0_outputs(8695)));
    layer1_outputs(774) <= not(layer0_outputs(6166)) or (layer0_outputs(6660));
    layer1_outputs(775) <= layer0_outputs(5558);
    layer1_outputs(776) <= '1';
    layer1_outputs(777) <= not(layer0_outputs(2197)) or (layer0_outputs(177));
    layer1_outputs(778) <= not(layer0_outputs(945));
    layer1_outputs(779) <= '1';
    layer1_outputs(780) <= (layer0_outputs(3224)) xor (layer0_outputs(281));
    layer1_outputs(781) <= not(layer0_outputs(1057)) or (layer0_outputs(9652));
    layer1_outputs(782) <= not(layer0_outputs(8079)) or (layer0_outputs(7293));
    layer1_outputs(783) <= not(layer0_outputs(3566));
    layer1_outputs(784) <= (layer0_outputs(9718)) and (layer0_outputs(9611));
    layer1_outputs(785) <= not(layer0_outputs(1208)) or (layer0_outputs(575));
    layer1_outputs(786) <= (layer0_outputs(1813)) and not (layer0_outputs(4815));
    layer1_outputs(787) <= (layer0_outputs(3746)) and not (layer0_outputs(3268));
    layer1_outputs(788) <= (layer0_outputs(422)) or (layer0_outputs(1180));
    layer1_outputs(789) <= '1';
    layer1_outputs(790) <= layer0_outputs(5714);
    layer1_outputs(791) <= not((layer0_outputs(9487)) or (layer0_outputs(8489)));
    layer1_outputs(792) <= layer0_outputs(5892);
    layer1_outputs(793) <= not(layer0_outputs(2418));
    layer1_outputs(794) <= (layer0_outputs(519)) and not (layer0_outputs(651));
    layer1_outputs(795) <= not(layer0_outputs(4462));
    layer1_outputs(796) <= not((layer0_outputs(9403)) xor (layer0_outputs(1241)));
    layer1_outputs(797) <= not((layer0_outputs(3619)) and (layer0_outputs(2466)));
    layer1_outputs(798) <= not((layer0_outputs(3544)) and (layer0_outputs(491)));
    layer1_outputs(799) <= '1';
    layer1_outputs(800) <= not((layer0_outputs(8135)) and (layer0_outputs(9724)));
    layer1_outputs(801) <= (layer0_outputs(2091)) and (layer0_outputs(6232));
    layer1_outputs(802) <= (layer0_outputs(8685)) or (layer0_outputs(8293));
    layer1_outputs(803) <= '1';
    layer1_outputs(804) <= layer0_outputs(8524);
    layer1_outputs(805) <= not(layer0_outputs(7164));
    layer1_outputs(806) <= layer0_outputs(6240);
    layer1_outputs(807) <= not((layer0_outputs(2336)) and (layer0_outputs(6773)));
    layer1_outputs(808) <= not(layer0_outputs(611)) or (layer0_outputs(9769));
    layer1_outputs(809) <= (layer0_outputs(1164)) and not (layer0_outputs(2648));
    layer1_outputs(810) <= not(layer0_outputs(2803));
    layer1_outputs(811) <= not((layer0_outputs(9780)) xor (layer0_outputs(2536)));
    layer1_outputs(812) <= not(layer0_outputs(1669));
    layer1_outputs(813) <= not(layer0_outputs(9833)) or (layer0_outputs(429));
    layer1_outputs(814) <= layer0_outputs(3603);
    layer1_outputs(815) <= layer0_outputs(4812);
    layer1_outputs(816) <= (layer0_outputs(8556)) and not (layer0_outputs(4709));
    layer1_outputs(817) <= (layer0_outputs(857)) or (layer0_outputs(863));
    layer1_outputs(818) <= layer0_outputs(2351);
    layer1_outputs(819) <= not(layer0_outputs(5073));
    layer1_outputs(820) <= not(layer0_outputs(8482)) or (layer0_outputs(8133));
    layer1_outputs(821) <= (layer0_outputs(889)) or (layer0_outputs(10201));
    layer1_outputs(822) <= not(layer0_outputs(3748));
    layer1_outputs(823) <= (layer0_outputs(5385)) and not (layer0_outputs(5000));
    layer1_outputs(824) <= not(layer0_outputs(3267));
    layer1_outputs(825) <= not(layer0_outputs(4357));
    layer1_outputs(826) <= not(layer0_outputs(3881));
    layer1_outputs(827) <= not(layer0_outputs(5860)) or (layer0_outputs(1789));
    layer1_outputs(828) <= layer0_outputs(7839);
    layer1_outputs(829) <= (layer0_outputs(4282)) or (layer0_outputs(7502));
    layer1_outputs(830) <= '1';
    layer1_outputs(831) <= not(layer0_outputs(9328));
    layer1_outputs(832) <= not(layer0_outputs(6970));
    layer1_outputs(833) <= not(layer0_outputs(5292));
    layer1_outputs(834) <= not((layer0_outputs(10117)) and (layer0_outputs(1822)));
    layer1_outputs(835) <= not(layer0_outputs(5424));
    layer1_outputs(836) <= (layer0_outputs(3596)) xor (layer0_outputs(5589));
    layer1_outputs(837) <= not(layer0_outputs(8805));
    layer1_outputs(838) <= not(layer0_outputs(5362));
    layer1_outputs(839) <= not(layer0_outputs(5132));
    layer1_outputs(840) <= not(layer0_outputs(2301));
    layer1_outputs(841) <= not((layer0_outputs(2727)) or (layer0_outputs(1870)));
    layer1_outputs(842) <= not((layer0_outputs(3359)) or (layer0_outputs(3290)));
    layer1_outputs(843) <= (layer0_outputs(3286)) and not (layer0_outputs(3334));
    layer1_outputs(844) <= (layer0_outputs(9480)) and (layer0_outputs(9452));
    layer1_outputs(845) <= not((layer0_outputs(7471)) and (layer0_outputs(1850)));
    layer1_outputs(846) <= (layer0_outputs(9317)) and (layer0_outputs(5364));
    layer1_outputs(847) <= not(layer0_outputs(1561));
    layer1_outputs(848) <= layer0_outputs(5790);
    layer1_outputs(849) <= not(layer0_outputs(6095));
    layer1_outputs(850) <= layer0_outputs(3992);
    layer1_outputs(851) <= not((layer0_outputs(9235)) and (layer0_outputs(9585)));
    layer1_outputs(852) <= not((layer0_outputs(7211)) and (layer0_outputs(209)));
    layer1_outputs(853) <= (layer0_outputs(4766)) xor (layer0_outputs(6764));
    layer1_outputs(854) <= not(layer0_outputs(8433));
    layer1_outputs(855) <= not(layer0_outputs(2578)) or (layer0_outputs(633));
    layer1_outputs(856) <= not((layer0_outputs(9140)) or (layer0_outputs(4644)));
    layer1_outputs(857) <= (layer0_outputs(6342)) and not (layer0_outputs(8554));
    layer1_outputs(858) <= not(layer0_outputs(4769)) or (layer0_outputs(10107));
    layer1_outputs(859) <= '1';
    layer1_outputs(860) <= not(layer0_outputs(8294)) or (layer0_outputs(5112));
    layer1_outputs(861) <= not(layer0_outputs(8423));
    layer1_outputs(862) <= not(layer0_outputs(6666)) or (layer0_outputs(5282));
    layer1_outputs(863) <= (layer0_outputs(6563)) and (layer0_outputs(1043));
    layer1_outputs(864) <= (layer0_outputs(3758)) and not (layer0_outputs(5915));
    layer1_outputs(865) <= layer0_outputs(5018);
    layer1_outputs(866) <= layer0_outputs(2770);
    layer1_outputs(867) <= not(layer0_outputs(2607)) or (layer0_outputs(4734));
    layer1_outputs(868) <= not(layer0_outputs(371));
    layer1_outputs(869) <= layer0_outputs(1199);
    layer1_outputs(870) <= (layer0_outputs(6970)) and not (layer0_outputs(9732));
    layer1_outputs(871) <= not(layer0_outputs(6810));
    layer1_outputs(872) <= not(layer0_outputs(7556)) or (layer0_outputs(988));
    layer1_outputs(873) <= not(layer0_outputs(1839));
    layer1_outputs(874) <= (layer0_outputs(2891)) or (layer0_outputs(6168));
    layer1_outputs(875) <= not(layer0_outputs(1945)) or (layer0_outputs(861));
    layer1_outputs(876) <= (layer0_outputs(6158)) xor (layer0_outputs(1630));
    layer1_outputs(877) <= (layer0_outputs(3256)) and (layer0_outputs(1125));
    layer1_outputs(878) <= (layer0_outputs(9302)) and not (layer0_outputs(7544));
    layer1_outputs(879) <= (layer0_outputs(8443)) and not (layer0_outputs(8574));
    layer1_outputs(880) <= (layer0_outputs(5106)) or (layer0_outputs(4985));
    layer1_outputs(881) <= not(layer0_outputs(7650)) or (layer0_outputs(2604));
    layer1_outputs(882) <= layer0_outputs(8103);
    layer1_outputs(883) <= '0';
    layer1_outputs(884) <= not(layer0_outputs(7581));
    layer1_outputs(885) <= not(layer0_outputs(9716));
    layer1_outputs(886) <= not(layer0_outputs(2877));
    layer1_outputs(887) <= not(layer0_outputs(6737)) or (layer0_outputs(9999));
    layer1_outputs(888) <= (layer0_outputs(2486)) or (layer0_outputs(5407));
    layer1_outputs(889) <= layer0_outputs(9044);
    layer1_outputs(890) <= (layer0_outputs(6769)) or (layer0_outputs(8766));
    layer1_outputs(891) <= layer0_outputs(8388);
    layer1_outputs(892) <= not(layer0_outputs(4304));
    layer1_outputs(893) <= layer0_outputs(8057);
    layer1_outputs(894) <= not((layer0_outputs(4408)) or (layer0_outputs(9706)));
    layer1_outputs(895) <= not((layer0_outputs(1287)) and (layer0_outputs(426)));
    layer1_outputs(896) <= (layer0_outputs(3024)) or (layer0_outputs(9466));
    layer1_outputs(897) <= '1';
    layer1_outputs(898) <= not((layer0_outputs(7564)) or (layer0_outputs(4831)));
    layer1_outputs(899) <= '0';
    layer1_outputs(900) <= '0';
    layer1_outputs(901) <= not(layer0_outputs(6030));
    layer1_outputs(902) <= not((layer0_outputs(3890)) and (layer0_outputs(4910)));
    layer1_outputs(903) <= layer0_outputs(885);
    layer1_outputs(904) <= layer0_outputs(3442);
    layer1_outputs(905) <= layer0_outputs(7640);
    layer1_outputs(906) <= layer0_outputs(5851);
    layer1_outputs(907) <= '0';
    layer1_outputs(908) <= layer0_outputs(4458);
    layer1_outputs(909) <= (layer0_outputs(4418)) or (layer0_outputs(8338));
    layer1_outputs(910) <= not(layer0_outputs(2712)) or (layer0_outputs(7999));
    layer1_outputs(911) <= (layer0_outputs(2988)) and not (layer0_outputs(2330));
    layer1_outputs(912) <= '0';
    layer1_outputs(913) <= not(layer0_outputs(268));
    layer1_outputs(914) <= not(layer0_outputs(3988));
    layer1_outputs(915) <= not(layer0_outputs(7266));
    layer1_outputs(916) <= not(layer0_outputs(1528)) or (layer0_outputs(9073));
    layer1_outputs(917) <= (layer0_outputs(2118)) and (layer0_outputs(763));
    layer1_outputs(918) <= layer0_outputs(9196);
    layer1_outputs(919) <= (layer0_outputs(8721)) and not (layer0_outputs(10123));
    layer1_outputs(920) <= layer0_outputs(8757);
    layer1_outputs(921) <= layer0_outputs(4438);
    layer1_outputs(922) <= not(layer0_outputs(1972));
    layer1_outputs(923) <= layer0_outputs(2436);
    layer1_outputs(924) <= layer0_outputs(5828);
    layer1_outputs(925) <= (layer0_outputs(2629)) or (layer0_outputs(65));
    layer1_outputs(926) <= not((layer0_outputs(680)) xor (layer0_outputs(3515)));
    layer1_outputs(927) <= not(layer0_outputs(1062)) or (layer0_outputs(7605));
    layer1_outputs(928) <= not(layer0_outputs(447));
    layer1_outputs(929) <= not(layer0_outputs(3803)) or (layer0_outputs(10161));
    layer1_outputs(930) <= not(layer0_outputs(8418)) or (layer0_outputs(8584));
    layer1_outputs(931) <= not(layer0_outputs(2647));
    layer1_outputs(932) <= not(layer0_outputs(4935)) or (layer0_outputs(451));
    layer1_outputs(933) <= layer0_outputs(6699);
    layer1_outputs(934) <= layer0_outputs(3028);
    layer1_outputs(935) <= not((layer0_outputs(10055)) xor (layer0_outputs(4212)));
    layer1_outputs(936) <= not(layer0_outputs(8872)) or (layer0_outputs(8192));
    layer1_outputs(937) <= not(layer0_outputs(2084)) or (layer0_outputs(8610));
    layer1_outputs(938) <= (layer0_outputs(8020)) and not (layer0_outputs(2300));
    layer1_outputs(939) <= not((layer0_outputs(3130)) or (layer0_outputs(3726)));
    layer1_outputs(940) <= not(layer0_outputs(753)) or (layer0_outputs(2764));
    layer1_outputs(941) <= layer0_outputs(8747);
    layer1_outputs(942) <= '0';
    layer1_outputs(943) <= not(layer0_outputs(992));
    layer1_outputs(944) <= '1';
    layer1_outputs(945) <= (layer0_outputs(6027)) and not (layer0_outputs(4050));
    layer1_outputs(946) <= not(layer0_outputs(566));
    layer1_outputs(947) <= layer0_outputs(10015);
    layer1_outputs(948) <= not(layer0_outputs(4469));
    layer1_outputs(949) <= layer0_outputs(2945);
    layer1_outputs(950) <= not(layer0_outputs(7757));
    layer1_outputs(951) <= not(layer0_outputs(3246));
    layer1_outputs(952) <= not(layer0_outputs(7110));
    layer1_outputs(953) <= (layer0_outputs(1090)) xor (layer0_outputs(7991));
    layer1_outputs(954) <= not(layer0_outputs(6568)) or (layer0_outputs(5646));
    layer1_outputs(955) <= not(layer0_outputs(3618)) or (layer0_outputs(6244));
    layer1_outputs(956) <= (layer0_outputs(4339)) or (layer0_outputs(8879));
    layer1_outputs(957) <= '0';
    layer1_outputs(958) <= not(layer0_outputs(2559)) or (layer0_outputs(5674));
    layer1_outputs(959) <= (layer0_outputs(8994)) xor (layer0_outputs(8828));
    layer1_outputs(960) <= not(layer0_outputs(9124));
    layer1_outputs(961) <= layer0_outputs(5597);
    layer1_outputs(962) <= not((layer0_outputs(1977)) or (layer0_outputs(5208)));
    layer1_outputs(963) <= (layer0_outputs(4349)) and not (layer0_outputs(4997));
    layer1_outputs(964) <= '0';
    layer1_outputs(965) <= layer0_outputs(6577);
    layer1_outputs(966) <= not(layer0_outputs(2912));
    layer1_outputs(967) <= (layer0_outputs(7819)) and not (layer0_outputs(2957));
    layer1_outputs(968) <= (layer0_outputs(3365)) and not (layer0_outputs(3008));
    layer1_outputs(969) <= (layer0_outputs(10108)) and not (layer0_outputs(1201));
    layer1_outputs(970) <= layer0_outputs(1635);
    layer1_outputs(971) <= layer0_outputs(8045);
    layer1_outputs(972) <= layer0_outputs(9881);
    layer1_outputs(973) <= not(layer0_outputs(4227));
    layer1_outputs(974) <= (layer0_outputs(3365)) and not (layer0_outputs(9272));
    layer1_outputs(975) <= not((layer0_outputs(4810)) or (layer0_outputs(7653)));
    layer1_outputs(976) <= (layer0_outputs(2)) xor (layer0_outputs(9159));
    layer1_outputs(977) <= (layer0_outputs(1586)) or (layer0_outputs(3798));
    layer1_outputs(978) <= layer0_outputs(3401);
    layer1_outputs(979) <= not(layer0_outputs(1782));
    layer1_outputs(980) <= not(layer0_outputs(4770));
    layer1_outputs(981) <= not((layer0_outputs(3943)) xor (layer0_outputs(9953)));
    layer1_outputs(982) <= (layer0_outputs(10172)) or (layer0_outputs(7179));
    layer1_outputs(983) <= layer0_outputs(7242);
    layer1_outputs(984) <= '1';
    layer1_outputs(985) <= not(layer0_outputs(4763)) or (layer0_outputs(7117));
    layer1_outputs(986) <= not(layer0_outputs(4030));
    layer1_outputs(987) <= not(layer0_outputs(1437));
    layer1_outputs(988) <= not((layer0_outputs(7290)) and (layer0_outputs(6258)));
    layer1_outputs(989) <= (layer0_outputs(7795)) and not (layer0_outputs(6938));
    layer1_outputs(990) <= (layer0_outputs(8464)) and not (layer0_outputs(1165));
    layer1_outputs(991) <= not(layer0_outputs(4930)) or (layer0_outputs(8927));
    layer1_outputs(992) <= (layer0_outputs(3504)) or (layer0_outputs(4239));
    layer1_outputs(993) <= not((layer0_outputs(2638)) xor (layer0_outputs(8862)));
    layer1_outputs(994) <= layer0_outputs(960);
    layer1_outputs(995) <= not((layer0_outputs(4553)) and (layer0_outputs(5637)));
    layer1_outputs(996) <= '0';
    layer1_outputs(997) <= not(layer0_outputs(6261)) or (layer0_outputs(6491));
    layer1_outputs(998) <= not(layer0_outputs(8817));
    layer1_outputs(999) <= not((layer0_outputs(7234)) or (layer0_outputs(3604)));
    layer1_outputs(1000) <= not((layer0_outputs(2919)) or (layer0_outputs(6651)));
    layer1_outputs(1001) <= layer0_outputs(2680);
    layer1_outputs(1002) <= not(layer0_outputs(4107)) or (layer0_outputs(1152));
    layer1_outputs(1003) <= (layer0_outputs(7162)) and (layer0_outputs(10235));
    layer1_outputs(1004) <= layer0_outputs(6397);
    layer1_outputs(1005) <= not(layer0_outputs(6190));
    layer1_outputs(1006) <= '0';
    layer1_outputs(1007) <= not((layer0_outputs(1342)) xor (layer0_outputs(5111)));
    layer1_outputs(1008) <= (layer0_outputs(539)) or (layer0_outputs(9519));
    layer1_outputs(1009) <= not(layer0_outputs(8888)) or (layer0_outputs(8489));
    layer1_outputs(1010) <= not(layer0_outputs(2293));
    layer1_outputs(1011) <= (layer0_outputs(7187)) and not (layer0_outputs(4435));
    layer1_outputs(1012) <= not(layer0_outputs(1734));
    layer1_outputs(1013) <= not(layer0_outputs(8801)) or (layer0_outputs(7290));
    layer1_outputs(1014) <= (layer0_outputs(5661)) and not (layer0_outputs(6924));
    layer1_outputs(1015) <= (layer0_outputs(3609)) or (layer0_outputs(4925));
    layer1_outputs(1016) <= (layer0_outputs(7978)) and (layer0_outputs(7201));
    layer1_outputs(1017) <= not((layer0_outputs(3827)) and (layer0_outputs(2399)));
    layer1_outputs(1018) <= layer0_outputs(1980);
    layer1_outputs(1019) <= not(layer0_outputs(3689));
    layer1_outputs(1020) <= not(layer0_outputs(7536)) or (layer0_outputs(676));
    layer1_outputs(1021) <= not((layer0_outputs(2649)) or (layer0_outputs(10046)));
    layer1_outputs(1022) <= not((layer0_outputs(7926)) or (layer0_outputs(6153)));
    layer1_outputs(1023) <= '1';
    layer1_outputs(1024) <= layer0_outputs(8172);
    layer1_outputs(1025) <= layer0_outputs(206);
    layer1_outputs(1026) <= (layer0_outputs(3383)) or (layer0_outputs(8624));
    layer1_outputs(1027) <= not((layer0_outputs(5104)) or (layer0_outputs(7154)));
    layer1_outputs(1028) <= not((layer0_outputs(8126)) or (layer0_outputs(9786)));
    layer1_outputs(1029) <= layer0_outputs(6359);
    layer1_outputs(1030) <= (layer0_outputs(7839)) and not (layer0_outputs(5287));
    layer1_outputs(1031) <= (layer0_outputs(585)) and (layer0_outputs(2026));
    layer1_outputs(1032) <= '0';
    layer1_outputs(1033) <= not(layer0_outputs(5359)) or (layer0_outputs(5632));
    layer1_outputs(1034) <= layer0_outputs(5771);
    layer1_outputs(1035) <= (layer0_outputs(7099)) or (layer0_outputs(5878));
    layer1_outputs(1036) <= not(layer0_outputs(10156));
    layer1_outputs(1037) <= (layer0_outputs(6049)) or (layer0_outputs(6252));
    layer1_outputs(1038) <= not(layer0_outputs(1787)) or (layer0_outputs(9286));
    layer1_outputs(1039) <= layer0_outputs(8318);
    layer1_outputs(1040) <= layer0_outputs(5673);
    layer1_outputs(1041) <= not(layer0_outputs(6128)) or (layer0_outputs(6565));
    layer1_outputs(1042) <= not((layer0_outputs(9119)) and (layer0_outputs(7565)));
    layer1_outputs(1043) <= (layer0_outputs(660)) and not (layer0_outputs(3715));
    layer1_outputs(1044) <= '1';
    layer1_outputs(1045) <= not(layer0_outputs(1610)) or (layer0_outputs(1533));
    layer1_outputs(1046) <= not((layer0_outputs(7694)) and (layer0_outputs(8789)));
    layer1_outputs(1047) <= layer0_outputs(3450);
    layer1_outputs(1048) <= layer0_outputs(1727);
    layer1_outputs(1049) <= '0';
    layer1_outputs(1050) <= not((layer0_outputs(9521)) and (layer0_outputs(4265)));
    layer1_outputs(1051) <= (layer0_outputs(3494)) and (layer0_outputs(618));
    layer1_outputs(1052) <= '0';
    layer1_outputs(1053) <= not(layer0_outputs(1993)) or (layer0_outputs(1030));
    layer1_outputs(1054) <= not((layer0_outputs(9395)) and (layer0_outputs(6668)));
    layer1_outputs(1055) <= not(layer0_outputs(2193));
    layer1_outputs(1056) <= (layer0_outputs(9269)) or (layer0_outputs(427));
    layer1_outputs(1057) <= layer0_outputs(9029);
    layer1_outputs(1058) <= (layer0_outputs(9589)) and (layer0_outputs(3942));
    layer1_outputs(1059) <= (layer0_outputs(5338)) and not (layer0_outputs(3203));
    layer1_outputs(1060) <= (layer0_outputs(1110)) xor (layer0_outputs(3930));
    layer1_outputs(1061) <= not((layer0_outputs(2816)) xor (layer0_outputs(9159)));
    layer1_outputs(1062) <= not(layer0_outputs(851));
    layer1_outputs(1063) <= layer0_outputs(318);
    layer1_outputs(1064) <= layer0_outputs(6786);
    layer1_outputs(1065) <= not(layer0_outputs(5303));
    layer1_outputs(1066) <= not(layer0_outputs(2101));
    layer1_outputs(1067) <= (layer0_outputs(4836)) and not (layer0_outputs(10111));
    layer1_outputs(1068) <= (layer0_outputs(3158)) xor (layer0_outputs(9987));
    layer1_outputs(1069) <= (layer0_outputs(3038)) and (layer0_outputs(8015));
    layer1_outputs(1070) <= (layer0_outputs(7014)) xor (layer0_outputs(6494));
    layer1_outputs(1071) <= not(layer0_outputs(8069));
    layer1_outputs(1072) <= not((layer0_outputs(9478)) and (layer0_outputs(8063)));
    layer1_outputs(1073) <= layer0_outputs(8298);
    layer1_outputs(1074) <= (layer0_outputs(8535)) and (layer0_outputs(4389));
    layer1_outputs(1075) <= '0';
    layer1_outputs(1076) <= not((layer0_outputs(5207)) and (layer0_outputs(6593)));
    layer1_outputs(1077) <= '1';
    layer1_outputs(1078) <= (layer0_outputs(3640)) or (layer0_outputs(5049));
    layer1_outputs(1079) <= (layer0_outputs(3872)) and (layer0_outputs(3447));
    layer1_outputs(1080) <= (layer0_outputs(8338)) and (layer0_outputs(10035));
    layer1_outputs(1081) <= not(layer0_outputs(9145));
    layer1_outputs(1082) <= layer0_outputs(4787);
    layer1_outputs(1083) <= '1';
    layer1_outputs(1084) <= not((layer0_outputs(9018)) xor (layer0_outputs(5319)));
    layer1_outputs(1085) <= (layer0_outputs(9705)) and not (layer0_outputs(6766));
    layer1_outputs(1086) <= '1';
    layer1_outputs(1087) <= (layer0_outputs(10225)) and (layer0_outputs(2562));
    layer1_outputs(1088) <= (layer0_outputs(9078)) and not (layer0_outputs(4762));
    layer1_outputs(1089) <= layer0_outputs(3787);
    layer1_outputs(1090) <= (layer0_outputs(7489)) and not (layer0_outputs(5747));
    layer1_outputs(1091) <= layer0_outputs(2003);
    layer1_outputs(1092) <= (layer0_outputs(9842)) and (layer0_outputs(6003));
    layer1_outputs(1093) <= layer0_outputs(2470);
    layer1_outputs(1094) <= (layer0_outputs(2809)) or (layer0_outputs(6767));
    layer1_outputs(1095) <= not(layer0_outputs(8618));
    layer1_outputs(1096) <= (layer0_outputs(898)) and (layer0_outputs(8548));
    layer1_outputs(1097) <= (layer0_outputs(7648)) and (layer0_outputs(2233));
    layer1_outputs(1098) <= (layer0_outputs(4871)) and not (layer0_outputs(8418));
    layer1_outputs(1099) <= not(layer0_outputs(1211)) or (layer0_outputs(290));
    layer1_outputs(1100) <= (layer0_outputs(3709)) xor (layer0_outputs(3544));
    layer1_outputs(1101) <= (layer0_outputs(4074)) xor (layer0_outputs(910));
    layer1_outputs(1102) <= layer0_outputs(8052);
    layer1_outputs(1103) <= (layer0_outputs(8901)) and not (layer0_outputs(2525));
    layer1_outputs(1104) <= (layer0_outputs(7107)) and not (layer0_outputs(7660));
    layer1_outputs(1105) <= (layer0_outputs(474)) and not (layer0_outputs(6635));
    layer1_outputs(1106) <= not(layer0_outputs(1846));
    layer1_outputs(1107) <= layer0_outputs(1228);
    layer1_outputs(1108) <= (layer0_outputs(6560)) and not (layer0_outputs(6370));
    layer1_outputs(1109) <= (layer0_outputs(8754)) and not (layer0_outputs(2345));
    layer1_outputs(1110) <= not((layer0_outputs(6462)) and (layer0_outputs(6111)));
    layer1_outputs(1111) <= (layer0_outputs(317)) and not (layer0_outputs(6535));
    layer1_outputs(1112) <= layer0_outputs(545);
    layer1_outputs(1113) <= layer0_outputs(7952);
    layer1_outputs(1114) <= not((layer0_outputs(3059)) or (layer0_outputs(6741)));
    layer1_outputs(1115) <= not(layer0_outputs(1995));
    layer1_outputs(1116) <= (layer0_outputs(8649)) and (layer0_outputs(9203));
    layer1_outputs(1117) <= '0';
    layer1_outputs(1118) <= layer0_outputs(8487);
    layer1_outputs(1119) <= '1';
    layer1_outputs(1120) <= not(layer0_outputs(1750));
    layer1_outputs(1121) <= layer0_outputs(5837);
    layer1_outputs(1122) <= layer0_outputs(1024);
    layer1_outputs(1123) <= not((layer0_outputs(7709)) or (layer0_outputs(9213)));
    layer1_outputs(1124) <= layer0_outputs(9289);
    layer1_outputs(1125) <= (layer0_outputs(7077)) and not (layer0_outputs(5202));
    layer1_outputs(1126) <= not((layer0_outputs(8059)) xor (layer0_outputs(9548)));
    layer1_outputs(1127) <= '0';
    layer1_outputs(1128) <= (layer0_outputs(248)) or (layer0_outputs(369));
    layer1_outputs(1129) <= (layer0_outputs(348)) or (layer0_outputs(8444));
    layer1_outputs(1130) <= layer0_outputs(4929);
    layer1_outputs(1131) <= not((layer0_outputs(2974)) and (layer0_outputs(5880)));
    layer1_outputs(1132) <= not((layer0_outputs(568)) or (layer0_outputs(8648)));
    layer1_outputs(1133) <= '1';
    layer1_outputs(1134) <= not(layer0_outputs(6764)) or (layer0_outputs(7415));
    layer1_outputs(1135) <= layer0_outputs(923);
    layer1_outputs(1136) <= (layer0_outputs(6375)) and not (layer0_outputs(4057));
    layer1_outputs(1137) <= not((layer0_outputs(6521)) xor (layer0_outputs(1739)));
    layer1_outputs(1138) <= not(layer0_outputs(6923));
    layer1_outputs(1139) <= (layer0_outputs(2831)) or (layer0_outputs(2092));
    layer1_outputs(1140) <= (layer0_outputs(2977)) and (layer0_outputs(5179));
    layer1_outputs(1141) <= (layer0_outputs(3738)) and (layer0_outputs(7226));
    layer1_outputs(1142) <= not((layer0_outputs(8167)) and (layer0_outputs(397)));
    layer1_outputs(1143) <= '0';
    layer1_outputs(1144) <= not(layer0_outputs(1704)) or (layer0_outputs(950));
    layer1_outputs(1145) <= (layer0_outputs(8885)) or (layer0_outputs(3561));
    layer1_outputs(1146) <= '0';
    layer1_outputs(1147) <= not(layer0_outputs(7986));
    layer1_outputs(1148) <= '1';
    layer1_outputs(1149) <= not(layer0_outputs(2450)) or (layer0_outputs(4311));
    layer1_outputs(1150) <= not(layer0_outputs(9355)) or (layer0_outputs(2697));
    layer1_outputs(1151) <= not(layer0_outputs(4854));
    layer1_outputs(1152) <= not(layer0_outputs(3442));
    layer1_outputs(1153) <= not(layer0_outputs(9502)) or (layer0_outputs(4713));
    layer1_outputs(1154) <= '1';
    layer1_outputs(1155) <= '1';
    layer1_outputs(1156) <= not((layer0_outputs(5099)) or (layer0_outputs(10071)));
    layer1_outputs(1157) <= not(layer0_outputs(7981)) or (layer0_outputs(3646));
    layer1_outputs(1158) <= layer0_outputs(382);
    layer1_outputs(1159) <= not((layer0_outputs(6476)) and (layer0_outputs(3527)));
    layer1_outputs(1160) <= (layer0_outputs(8006)) or (layer0_outputs(3294));
    layer1_outputs(1161) <= (layer0_outputs(5671)) or (layer0_outputs(1984));
    layer1_outputs(1162) <= not((layer0_outputs(5115)) xor (layer0_outputs(9313)));
    layer1_outputs(1163) <= not(layer0_outputs(9847)) or (layer0_outputs(5328));
    layer1_outputs(1164) <= '1';
    layer1_outputs(1165) <= not((layer0_outputs(5489)) or (layer0_outputs(7724)));
    layer1_outputs(1166) <= not(layer0_outputs(9177)) or (layer0_outputs(1825));
    layer1_outputs(1167) <= (layer0_outputs(9749)) or (layer0_outputs(8512));
    layer1_outputs(1168) <= layer0_outputs(2141);
    layer1_outputs(1169) <= not((layer0_outputs(6571)) and (layer0_outputs(9273)));
    layer1_outputs(1170) <= (layer0_outputs(7611)) and not (layer0_outputs(4896));
    layer1_outputs(1171) <= (layer0_outputs(8502)) and not (layer0_outputs(6125));
    layer1_outputs(1172) <= '0';
    layer1_outputs(1173) <= (layer0_outputs(3859)) and (layer0_outputs(3813));
    layer1_outputs(1174) <= (layer0_outputs(3370)) and not (layer0_outputs(1346));
    layer1_outputs(1175) <= layer0_outputs(5883);
    layer1_outputs(1176) <= '0';
    layer1_outputs(1177) <= not(layer0_outputs(8349));
    layer1_outputs(1178) <= (layer0_outputs(339)) or (layer0_outputs(6605));
    layer1_outputs(1179) <= not(layer0_outputs(8613));
    layer1_outputs(1180) <= not((layer0_outputs(8639)) and (layer0_outputs(7868)));
    layer1_outputs(1181) <= not(layer0_outputs(4253));
    layer1_outputs(1182) <= not((layer0_outputs(5385)) and (layer0_outputs(1514)));
    layer1_outputs(1183) <= not((layer0_outputs(709)) and (layer0_outputs(9296)));
    layer1_outputs(1184) <= not(layer0_outputs(6127));
    layer1_outputs(1185) <= (layer0_outputs(760)) xor (layer0_outputs(165));
    layer1_outputs(1186) <= '0';
    layer1_outputs(1187) <= not(layer0_outputs(566)) or (layer0_outputs(3343));
    layer1_outputs(1188) <= not(layer0_outputs(7161));
    layer1_outputs(1189) <= not(layer0_outputs(3888));
    layer1_outputs(1190) <= (layer0_outputs(1374)) and not (layer0_outputs(1655));
    layer1_outputs(1191) <= (layer0_outputs(6349)) xor (layer0_outputs(9496));
    layer1_outputs(1192) <= layer0_outputs(3240);
    layer1_outputs(1193) <= not(layer0_outputs(3502)) or (layer0_outputs(2383));
    layer1_outputs(1194) <= (layer0_outputs(2493)) or (layer0_outputs(7985));
    layer1_outputs(1195) <= layer0_outputs(4279);
    layer1_outputs(1196) <= not(layer0_outputs(7063));
    layer1_outputs(1197) <= layer0_outputs(10097);
    layer1_outputs(1198) <= not(layer0_outputs(10190));
    layer1_outputs(1199) <= not((layer0_outputs(9579)) and (layer0_outputs(2322)));
    layer1_outputs(1200) <= not(layer0_outputs(2404)) or (layer0_outputs(8714));
    layer1_outputs(1201) <= not((layer0_outputs(8019)) xor (layer0_outputs(608)));
    layer1_outputs(1202) <= (layer0_outputs(1826)) or (layer0_outputs(955));
    layer1_outputs(1203) <= (layer0_outputs(5501)) and (layer0_outputs(130));
    layer1_outputs(1204) <= layer0_outputs(825);
    layer1_outputs(1205) <= not((layer0_outputs(10093)) or (layer0_outputs(4392)));
    layer1_outputs(1206) <= layer0_outputs(4973);
    layer1_outputs(1207) <= not(layer0_outputs(6995)) or (layer0_outputs(5531));
    layer1_outputs(1208) <= not(layer0_outputs(7588));
    layer1_outputs(1209) <= not((layer0_outputs(7337)) xor (layer0_outputs(2910)));
    layer1_outputs(1210) <= layer0_outputs(4319);
    layer1_outputs(1211) <= (layer0_outputs(5778)) or (layer0_outputs(6588));
    layer1_outputs(1212) <= not((layer0_outputs(8980)) and (layer0_outputs(5215)));
    layer1_outputs(1213) <= not(layer0_outputs(4215));
    layer1_outputs(1214) <= (layer0_outputs(690)) or (layer0_outputs(209));
    layer1_outputs(1215) <= not(layer0_outputs(7340)) or (layer0_outputs(1012));
    layer1_outputs(1216) <= (layer0_outputs(4170)) or (layer0_outputs(5433));
    layer1_outputs(1217) <= not(layer0_outputs(9158)) or (layer0_outputs(9669));
    layer1_outputs(1218) <= not(layer0_outputs(9322));
    layer1_outputs(1219) <= layer0_outputs(7162);
    layer1_outputs(1220) <= not((layer0_outputs(7398)) xor (layer0_outputs(4394)));
    layer1_outputs(1221) <= (layer0_outputs(9647)) and not (layer0_outputs(3425));
    layer1_outputs(1222) <= (layer0_outputs(5110)) xor (layer0_outputs(8829));
    layer1_outputs(1223) <= not(layer0_outputs(2499));
    layer1_outputs(1224) <= '1';
    layer1_outputs(1225) <= (layer0_outputs(7358)) and not (layer0_outputs(10098));
    layer1_outputs(1226) <= not((layer0_outputs(3303)) or (layer0_outputs(8811)));
    layer1_outputs(1227) <= (layer0_outputs(8295)) xor (layer0_outputs(418));
    layer1_outputs(1228) <= not((layer0_outputs(4010)) xor (layer0_outputs(6884)));
    layer1_outputs(1229) <= not((layer0_outputs(9577)) and (layer0_outputs(8860)));
    layer1_outputs(1230) <= not(layer0_outputs(3542)) or (layer0_outputs(8976));
    layer1_outputs(1231) <= (layer0_outputs(5726)) and (layer0_outputs(9619));
    layer1_outputs(1232) <= layer0_outputs(8258);
    layer1_outputs(1233) <= layer0_outputs(4579);
    layer1_outputs(1234) <= not((layer0_outputs(8710)) or (layer0_outputs(2123)));
    layer1_outputs(1235) <= layer0_outputs(6983);
    layer1_outputs(1236) <= (layer0_outputs(9096)) and not (layer0_outputs(5772));
    layer1_outputs(1237) <= '1';
    layer1_outputs(1238) <= not(layer0_outputs(1198));
    layer1_outputs(1239) <= not(layer0_outputs(9880)) or (layer0_outputs(8997));
    layer1_outputs(1240) <= not((layer0_outputs(2833)) and (layer0_outputs(7586)));
    layer1_outputs(1241) <= layer0_outputs(1684);
    layer1_outputs(1242) <= (layer0_outputs(7518)) xor (layer0_outputs(9027));
    layer1_outputs(1243) <= not(layer0_outputs(4927));
    layer1_outputs(1244) <= layer0_outputs(4347);
    layer1_outputs(1245) <= not((layer0_outputs(8818)) or (layer0_outputs(8898)));
    layer1_outputs(1246) <= '1';
    layer1_outputs(1247) <= layer0_outputs(6724);
    layer1_outputs(1248) <= layer0_outputs(4337);
    layer1_outputs(1249) <= not(layer0_outputs(7677));
    layer1_outputs(1250) <= (layer0_outputs(2770)) or (layer0_outputs(1066));
    layer1_outputs(1251) <= (layer0_outputs(1496)) and not (layer0_outputs(1956));
    layer1_outputs(1252) <= not(layer0_outputs(9218));
    layer1_outputs(1253) <= layer0_outputs(749);
    layer1_outputs(1254) <= not(layer0_outputs(5639)) or (layer0_outputs(1853));
    layer1_outputs(1255) <= (layer0_outputs(1949)) and (layer0_outputs(7001));
    layer1_outputs(1256) <= layer0_outputs(219);
    layer1_outputs(1257) <= not(layer0_outputs(4229)) or (layer0_outputs(8064));
    layer1_outputs(1258) <= layer0_outputs(9291);
    layer1_outputs(1259) <= not(layer0_outputs(9115)) or (layer0_outputs(4496));
    layer1_outputs(1260) <= not(layer0_outputs(3640));
    layer1_outputs(1261) <= not(layer0_outputs(6045));
    layer1_outputs(1262) <= not(layer0_outputs(5247)) or (layer0_outputs(4676));
    layer1_outputs(1263) <= not(layer0_outputs(8492)) or (layer0_outputs(7195));
    layer1_outputs(1264) <= not((layer0_outputs(1677)) and (layer0_outputs(4195)));
    layer1_outputs(1265) <= layer0_outputs(9288);
    layer1_outputs(1266) <= not((layer0_outputs(459)) xor (layer0_outputs(4052)));
    layer1_outputs(1267) <= not(layer0_outputs(6943));
    layer1_outputs(1268) <= not(layer0_outputs(1628)) or (layer0_outputs(3022));
    layer1_outputs(1269) <= (layer0_outputs(4239)) and not (layer0_outputs(6708));
    layer1_outputs(1270) <= not((layer0_outputs(2183)) or (layer0_outputs(5959)));
    layer1_outputs(1271) <= layer0_outputs(9470);
    layer1_outputs(1272) <= layer0_outputs(8148);
    layer1_outputs(1273) <= not(layer0_outputs(5649));
    layer1_outputs(1274) <= not(layer0_outputs(2721)) or (layer0_outputs(9977));
    layer1_outputs(1275) <= (layer0_outputs(8415)) and (layer0_outputs(4801));
    layer1_outputs(1276) <= not((layer0_outputs(1228)) and (layer0_outputs(1702)));
    layer1_outputs(1277) <= (layer0_outputs(3911)) and not (layer0_outputs(1535));
    layer1_outputs(1278) <= '0';
    layer1_outputs(1279) <= not(layer0_outputs(3310));
    layer1_outputs(1280) <= not(layer0_outputs(9748)) or (layer0_outputs(7372));
    layer1_outputs(1281) <= not((layer0_outputs(8497)) and (layer0_outputs(10175)));
    layer1_outputs(1282) <= (layer0_outputs(7703)) and not (layer0_outputs(4773));
    layer1_outputs(1283) <= not(layer0_outputs(2565));
    layer1_outputs(1284) <= '0';
    layer1_outputs(1285) <= not(layer0_outputs(5371));
    layer1_outputs(1286) <= not((layer0_outputs(1417)) and (layer0_outputs(3644)));
    layer1_outputs(1287) <= not(layer0_outputs(4113)) or (layer0_outputs(230));
    layer1_outputs(1288) <= not(layer0_outputs(5586));
    layer1_outputs(1289) <= layer0_outputs(6341);
    layer1_outputs(1290) <= not((layer0_outputs(4660)) and (layer0_outputs(8868)));
    layer1_outputs(1291) <= not(layer0_outputs(1832));
    layer1_outputs(1292) <= (layer0_outputs(7579)) and not (layer0_outputs(4212));
    layer1_outputs(1293) <= '0';
    layer1_outputs(1294) <= (layer0_outputs(3105)) and not (layer0_outputs(9210));
    layer1_outputs(1295) <= layer0_outputs(8210);
    layer1_outputs(1296) <= (layer0_outputs(6526)) or (layer0_outputs(5301));
    layer1_outputs(1297) <= not(layer0_outputs(4346)) or (layer0_outputs(8012));
    layer1_outputs(1298) <= not(layer0_outputs(9863));
    layer1_outputs(1299) <= (layer0_outputs(7381)) and (layer0_outputs(6503));
    layer1_outputs(1300) <= layer0_outputs(5416);
    layer1_outputs(1301) <= (layer0_outputs(4135)) xor (layer0_outputs(1638));
    layer1_outputs(1302) <= not((layer0_outputs(5542)) xor (layer0_outputs(867)));
    layer1_outputs(1303) <= layer0_outputs(1503);
    layer1_outputs(1304) <= (layer0_outputs(6811)) and not (layer0_outputs(7130));
    layer1_outputs(1305) <= layer0_outputs(6701);
    layer1_outputs(1306) <= not(layer0_outputs(6562)) or (layer0_outputs(1741));
    layer1_outputs(1307) <= (layer0_outputs(3575)) xor (layer0_outputs(3473));
    layer1_outputs(1308) <= (layer0_outputs(9262)) and (layer0_outputs(7174));
    layer1_outputs(1309) <= not(layer0_outputs(9282));
    layer1_outputs(1310) <= (layer0_outputs(3564)) and not (layer0_outputs(7626));
    layer1_outputs(1311) <= not((layer0_outputs(7412)) or (layer0_outputs(6292)));
    layer1_outputs(1312) <= layer0_outputs(1347);
    layer1_outputs(1313) <= not((layer0_outputs(4826)) and (layer0_outputs(7627)));
    layer1_outputs(1314) <= layer0_outputs(5188);
    layer1_outputs(1315) <= not((layer0_outputs(3672)) and (layer0_outputs(4086)));
    layer1_outputs(1316) <= not(layer0_outputs(5490)) or (layer0_outputs(1263));
    layer1_outputs(1317) <= (layer0_outputs(5216)) and not (layer0_outputs(6139));
    layer1_outputs(1318) <= not((layer0_outputs(4314)) xor (layer0_outputs(7147)));
    layer1_outputs(1319) <= not((layer0_outputs(3403)) and (layer0_outputs(2560)));
    layer1_outputs(1320) <= (layer0_outputs(3113)) xor (layer0_outputs(1403));
    layer1_outputs(1321) <= (layer0_outputs(2256)) or (layer0_outputs(4218));
    layer1_outputs(1322) <= not(layer0_outputs(290));
    layer1_outputs(1323) <= not(layer0_outputs(4601));
    layer1_outputs(1324) <= not(layer0_outputs(7577));
    layer1_outputs(1325) <= layer0_outputs(4060);
    layer1_outputs(1326) <= not(layer0_outputs(4380));
    layer1_outputs(1327) <= not(layer0_outputs(1781)) or (layer0_outputs(6146));
    layer1_outputs(1328) <= (layer0_outputs(2896)) and not (layer0_outputs(10047));
    layer1_outputs(1329) <= (layer0_outputs(3388)) or (layer0_outputs(9152));
    layer1_outputs(1330) <= layer0_outputs(8151);
    layer1_outputs(1331) <= (layer0_outputs(7086)) and not (layer0_outputs(2456));
    layer1_outputs(1332) <= not(layer0_outputs(2741)) or (layer0_outputs(9572));
    layer1_outputs(1333) <= not((layer0_outputs(8114)) and (layer0_outputs(2676)));
    layer1_outputs(1334) <= (layer0_outputs(3662)) and not (layer0_outputs(3455));
    layer1_outputs(1335) <= (layer0_outputs(4599)) and (layer0_outputs(4823));
    layer1_outputs(1336) <= not(layer0_outputs(2487)) or (layer0_outputs(5275));
    layer1_outputs(1337) <= layer0_outputs(9790);
    layer1_outputs(1338) <= layer0_outputs(6825);
    layer1_outputs(1339) <= not(layer0_outputs(3491));
    layer1_outputs(1340) <= not((layer0_outputs(4685)) xor (layer0_outputs(7163)));
    layer1_outputs(1341) <= layer0_outputs(7026);
    layer1_outputs(1342) <= not(layer0_outputs(5780)) or (layer0_outputs(6213));
    layer1_outputs(1343) <= not((layer0_outputs(5451)) and (layer0_outputs(7718)));
    layer1_outputs(1344) <= not(layer0_outputs(7079));
    layer1_outputs(1345) <= (layer0_outputs(3673)) and not (layer0_outputs(8784));
    layer1_outputs(1346) <= (layer0_outputs(7560)) xor (layer0_outputs(7876));
    layer1_outputs(1347) <= not(layer0_outputs(7997));
    layer1_outputs(1348) <= '0';
    layer1_outputs(1349) <= (layer0_outputs(8936)) and (layer0_outputs(2264));
    layer1_outputs(1350) <= (layer0_outputs(6664)) and not (layer0_outputs(6765));
    layer1_outputs(1351) <= layer0_outputs(1937);
    layer1_outputs(1352) <= not((layer0_outputs(138)) or (layer0_outputs(5621)));
    layer1_outputs(1353) <= not(layer0_outputs(5663));
    layer1_outputs(1354) <= layer0_outputs(7092);
    layer1_outputs(1355) <= not((layer0_outputs(2180)) xor (layer0_outputs(1552)));
    layer1_outputs(1356) <= '1';
    layer1_outputs(1357) <= (layer0_outputs(2958)) and not (layer0_outputs(5658));
    layer1_outputs(1358) <= (layer0_outputs(5767)) and not (layer0_outputs(1732));
    layer1_outputs(1359) <= not(layer0_outputs(8632));
    layer1_outputs(1360) <= not(layer0_outputs(464)) or (layer0_outputs(9008));
    layer1_outputs(1361) <= not((layer0_outputs(99)) and (layer0_outputs(4897)));
    layer1_outputs(1362) <= layer0_outputs(615);
    layer1_outputs(1363) <= (layer0_outputs(6177)) and not (layer0_outputs(1335));
    layer1_outputs(1364) <= layer0_outputs(1156);
    layer1_outputs(1365) <= (layer0_outputs(584)) and not (layer0_outputs(9180));
    layer1_outputs(1366) <= not(layer0_outputs(1409));
    layer1_outputs(1367) <= '0';
    layer1_outputs(1368) <= (layer0_outputs(3229)) and (layer0_outputs(4228));
    layer1_outputs(1369) <= not(layer0_outputs(2468));
    layer1_outputs(1370) <= not(layer0_outputs(6255));
    layer1_outputs(1371) <= not(layer0_outputs(8143)) or (layer0_outputs(6767));
    layer1_outputs(1372) <= not((layer0_outputs(10015)) or (layer0_outputs(9011)));
    layer1_outputs(1373) <= not(layer0_outputs(5480)) or (layer0_outputs(6393));
    layer1_outputs(1374) <= not(layer0_outputs(3336));
    layer1_outputs(1375) <= not(layer0_outputs(321));
    layer1_outputs(1376) <= not(layer0_outputs(110));
    layer1_outputs(1377) <= not((layer0_outputs(3215)) or (layer0_outputs(7632)));
    layer1_outputs(1378) <= not(layer0_outputs(358)) or (layer0_outputs(1743));
    layer1_outputs(1379) <= not((layer0_outputs(275)) or (layer0_outputs(6752)));
    layer1_outputs(1380) <= not(layer0_outputs(4793));
    layer1_outputs(1381) <= layer0_outputs(8526);
    layer1_outputs(1382) <= not(layer0_outputs(1422));
    layer1_outputs(1383) <= (layer0_outputs(3425)) xor (layer0_outputs(7580));
    layer1_outputs(1384) <= (layer0_outputs(6468)) and not (layer0_outputs(4004));
    layer1_outputs(1385) <= not((layer0_outputs(4213)) xor (layer0_outputs(7010)));
    layer1_outputs(1386) <= layer0_outputs(6680);
    layer1_outputs(1387) <= layer0_outputs(6591);
    layer1_outputs(1388) <= (layer0_outputs(3560)) or (layer0_outputs(992));
    layer1_outputs(1389) <= '1';
    layer1_outputs(1390) <= layer0_outputs(682);
    layer1_outputs(1391) <= layer0_outputs(618);
    layer1_outputs(1392) <= (layer0_outputs(8065)) xor (layer0_outputs(6052));
    layer1_outputs(1393) <= (layer0_outputs(8236)) and not (layer0_outputs(1865));
    layer1_outputs(1394) <= (layer0_outputs(1820)) xor (layer0_outputs(6726));
    layer1_outputs(1395) <= (layer0_outputs(5079)) xor (layer0_outputs(1836));
    layer1_outputs(1396) <= '1';
    layer1_outputs(1397) <= (layer0_outputs(5056)) and not (layer0_outputs(4174));
    layer1_outputs(1398) <= layer0_outputs(8925);
    layer1_outputs(1399) <= '0';
    layer1_outputs(1400) <= (layer0_outputs(1920)) xor (layer0_outputs(4873));
    layer1_outputs(1401) <= '1';
    layer1_outputs(1402) <= (layer0_outputs(7435)) or (layer0_outputs(3249));
    layer1_outputs(1403) <= not(layer0_outputs(3234)) or (layer0_outputs(8592));
    layer1_outputs(1404) <= not(layer0_outputs(5438)) or (layer0_outputs(3333));
    layer1_outputs(1405) <= not(layer0_outputs(5946));
    layer1_outputs(1406) <= (layer0_outputs(9139)) or (layer0_outputs(2672));
    layer1_outputs(1407) <= not((layer0_outputs(3922)) and (layer0_outputs(2128)));
    layer1_outputs(1408) <= not((layer0_outputs(7360)) or (layer0_outputs(3595)));
    layer1_outputs(1409) <= layer0_outputs(8842);
    layer1_outputs(1410) <= layer0_outputs(4865);
    layer1_outputs(1411) <= layer0_outputs(647);
    layer1_outputs(1412) <= (layer0_outputs(6073)) and not (layer0_outputs(7018));
    layer1_outputs(1413) <= not(layer0_outputs(3917)) or (layer0_outputs(6419));
    layer1_outputs(1414) <= layer0_outputs(7941);
    layer1_outputs(1415) <= (layer0_outputs(6799)) xor (layer0_outputs(10102));
    layer1_outputs(1416) <= not((layer0_outputs(1633)) or (layer0_outputs(3180)));
    layer1_outputs(1417) <= not((layer0_outputs(6933)) or (layer0_outputs(7358)));
    layer1_outputs(1418) <= (layer0_outputs(9372)) xor (layer0_outputs(9172));
    layer1_outputs(1419) <= not(layer0_outputs(8447)) or (layer0_outputs(5067));
    layer1_outputs(1420) <= '1';
    layer1_outputs(1421) <= not((layer0_outputs(7561)) and (layer0_outputs(5597)));
    layer1_outputs(1422) <= (layer0_outputs(6424)) and not (layer0_outputs(6669));
    layer1_outputs(1423) <= not(layer0_outputs(3053)) or (layer0_outputs(6599));
    layer1_outputs(1424) <= not(layer0_outputs(3133));
    layer1_outputs(1425) <= not(layer0_outputs(5744)) or (layer0_outputs(7582));
    layer1_outputs(1426) <= (layer0_outputs(711)) and not (layer0_outputs(6981));
    layer1_outputs(1427) <= not(layer0_outputs(6085));
    layer1_outputs(1428) <= not((layer0_outputs(1999)) xor (layer0_outputs(3686)));
    layer1_outputs(1429) <= layer0_outputs(4358);
    layer1_outputs(1430) <= not(layer0_outputs(2320));
    layer1_outputs(1431) <= not(layer0_outputs(4556));
    layer1_outputs(1432) <= (layer0_outputs(5567)) and (layer0_outputs(1918));
    layer1_outputs(1433) <= not(layer0_outputs(3484));
    layer1_outputs(1434) <= (layer0_outputs(4589)) and (layer0_outputs(9117));
    layer1_outputs(1435) <= '1';
    layer1_outputs(1436) <= not(layer0_outputs(5286));
    layer1_outputs(1437) <= not((layer0_outputs(3641)) xor (layer0_outputs(8485)));
    layer1_outputs(1438) <= '0';
    layer1_outputs(1439) <= not(layer0_outputs(2164));
    layer1_outputs(1440) <= not((layer0_outputs(2491)) or (layer0_outputs(7552)));
    layer1_outputs(1441) <= (layer0_outputs(700)) and not (layer0_outputs(4092));
    layer1_outputs(1442) <= (layer0_outputs(6491)) and (layer0_outputs(7575));
    layer1_outputs(1443) <= (layer0_outputs(9181)) or (layer0_outputs(5723));
    layer1_outputs(1444) <= (layer0_outputs(2036)) and not (layer0_outputs(9267));
    layer1_outputs(1445) <= '0';
    layer1_outputs(1446) <= (layer0_outputs(5705)) and not (layer0_outputs(2391));
    layer1_outputs(1447) <= (layer0_outputs(6429)) and (layer0_outputs(7214));
    layer1_outputs(1448) <= (layer0_outputs(5077)) xor (layer0_outputs(5637));
    layer1_outputs(1449) <= layer0_outputs(7492);
    layer1_outputs(1450) <= not(layer0_outputs(666)) or (layer0_outputs(4068));
    layer1_outputs(1451) <= (layer0_outputs(641)) or (layer0_outputs(523));
    layer1_outputs(1452) <= (layer0_outputs(6295)) and not (layer0_outputs(1891));
    layer1_outputs(1453) <= (layer0_outputs(4944)) and not (layer0_outputs(9227));
    layer1_outputs(1454) <= not(layer0_outputs(2101));
    layer1_outputs(1455) <= (layer0_outputs(1885)) xor (layer0_outputs(2888));
    layer1_outputs(1456) <= not(layer0_outputs(6833));
    layer1_outputs(1457) <= not(layer0_outputs(9473)) or (layer0_outputs(162));
    layer1_outputs(1458) <= (layer0_outputs(8501)) or (layer0_outputs(7895));
    layer1_outputs(1459) <= not(layer0_outputs(1105)) or (layer0_outputs(9258));
    layer1_outputs(1460) <= (layer0_outputs(4876)) and (layer0_outputs(3743));
    layer1_outputs(1461) <= '1';
    layer1_outputs(1462) <= not(layer0_outputs(4618)) or (layer0_outputs(9394));
    layer1_outputs(1463) <= (layer0_outputs(5900)) and (layer0_outputs(2292));
    layer1_outputs(1464) <= (layer0_outputs(4864)) or (layer0_outputs(6712));
    layer1_outputs(1465) <= not(layer0_outputs(5737));
    layer1_outputs(1466) <= (layer0_outputs(3651)) and not (layer0_outputs(473));
    layer1_outputs(1467) <= layer0_outputs(2497);
    layer1_outputs(1468) <= layer0_outputs(2564);
    layer1_outputs(1469) <= not(layer0_outputs(3157));
    layer1_outputs(1470) <= not(layer0_outputs(4172)) or (layer0_outputs(1084));
    layer1_outputs(1471) <= (layer0_outputs(297)) and not (layer0_outputs(8242));
    layer1_outputs(1472) <= (layer0_outputs(3244)) xor (layer0_outputs(2279));
    layer1_outputs(1473) <= (layer0_outputs(10014)) or (layer0_outputs(8138));
    layer1_outputs(1474) <= not((layer0_outputs(5329)) xor (layer0_outputs(4153)));
    layer1_outputs(1475) <= not(layer0_outputs(10075));
    layer1_outputs(1476) <= (layer0_outputs(1017)) and not (layer0_outputs(105));
    layer1_outputs(1477) <= not((layer0_outputs(8612)) or (layer0_outputs(6649)));
    layer1_outputs(1478) <= not(layer0_outputs(5335)) or (layer0_outputs(9481));
    layer1_outputs(1479) <= not(layer0_outputs(3089));
    layer1_outputs(1480) <= not((layer0_outputs(6076)) and (layer0_outputs(9518)));
    layer1_outputs(1481) <= layer0_outputs(6898);
    layer1_outputs(1482) <= not(layer0_outputs(1964)) or (layer0_outputs(5800));
    layer1_outputs(1483) <= not((layer0_outputs(3483)) or (layer0_outputs(9660)));
    layer1_outputs(1484) <= not((layer0_outputs(6902)) or (layer0_outputs(8847)));
    layer1_outputs(1485) <= not(layer0_outputs(1040));
    layer1_outputs(1486) <= '1';
    layer1_outputs(1487) <= not(layer0_outputs(1037)) or (layer0_outputs(5855));
    layer1_outputs(1488) <= (layer0_outputs(3807)) or (layer0_outputs(6519));
    layer1_outputs(1489) <= '0';
    layer1_outputs(1490) <= (layer0_outputs(7012)) and not (layer0_outputs(8033));
    layer1_outputs(1491) <= (layer0_outputs(5331)) and (layer0_outputs(2079));
    layer1_outputs(1492) <= (layer0_outputs(1647)) and not (layer0_outputs(2703));
    layer1_outputs(1493) <= (layer0_outputs(388)) and not (layer0_outputs(684));
    layer1_outputs(1494) <= '0';
    layer1_outputs(1495) <= (layer0_outputs(6591)) and not (layer0_outputs(8761));
    layer1_outputs(1496) <= not(layer0_outputs(6483));
    layer1_outputs(1497) <= (layer0_outputs(4414)) and not (layer0_outputs(4457));
    layer1_outputs(1498) <= not(layer0_outputs(3594));
    layer1_outputs(1499) <= not(layer0_outputs(2609)) or (layer0_outputs(1483));
    layer1_outputs(1500) <= not(layer0_outputs(6374));
    layer1_outputs(1501) <= (layer0_outputs(2477)) and (layer0_outputs(4422));
    layer1_outputs(1502) <= not(layer0_outputs(1605));
    layer1_outputs(1503) <= not(layer0_outputs(1207));
    layer1_outputs(1504) <= not((layer0_outputs(7275)) xor (layer0_outputs(8439)));
    layer1_outputs(1505) <= layer0_outputs(6320);
    layer1_outputs(1506) <= (layer0_outputs(5779)) and not (layer0_outputs(7227));
    layer1_outputs(1507) <= layer0_outputs(1561);
    layer1_outputs(1508) <= not((layer0_outputs(9787)) and (layer0_outputs(9589)));
    layer1_outputs(1509) <= not((layer0_outputs(8768)) xor (layer0_outputs(9134)));
    layer1_outputs(1510) <= not(layer0_outputs(5794));
    layer1_outputs(1511) <= not(layer0_outputs(2824));
    layer1_outputs(1512) <= not((layer0_outputs(6956)) or (layer0_outputs(6405)));
    layer1_outputs(1513) <= layer0_outputs(8203);
    layer1_outputs(1514) <= layer0_outputs(6704);
    layer1_outputs(1515) <= not(layer0_outputs(1979)) or (layer0_outputs(4885));
    layer1_outputs(1516) <= (layer0_outputs(2457)) and not (layer0_outputs(8654));
    layer1_outputs(1517) <= not((layer0_outputs(2994)) and (layer0_outputs(1236)));
    layer1_outputs(1518) <= layer0_outputs(8525);
    layer1_outputs(1519) <= not((layer0_outputs(4699)) and (layer0_outputs(5009)));
    layer1_outputs(1520) <= layer0_outputs(2602);
    layer1_outputs(1521) <= not(layer0_outputs(9396));
    layer1_outputs(1522) <= layer0_outputs(2894);
    layer1_outputs(1523) <= not(layer0_outputs(5485)) or (layer0_outputs(565));
    layer1_outputs(1524) <= (layer0_outputs(7019)) xor (layer0_outputs(649));
    layer1_outputs(1525) <= (layer0_outputs(2276)) or (layer0_outputs(5248));
    layer1_outputs(1526) <= not((layer0_outputs(1055)) and (layer0_outputs(6492)));
    layer1_outputs(1527) <= layer0_outputs(6535);
    layer1_outputs(1528) <= (layer0_outputs(8874)) and not (layer0_outputs(1783));
    layer1_outputs(1529) <= layer0_outputs(7632);
    layer1_outputs(1530) <= (layer0_outputs(8247)) and not (layer0_outputs(3722));
    layer1_outputs(1531) <= not(layer0_outputs(8101));
    layer1_outputs(1532) <= not((layer0_outputs(5222)) xor (layer0_outputs(4402)));
    layer1_outputs(1533) <= (layer0_outputs(9788)) or (layer0_outputs(7330));
    layer1_outputs(1534) <= not(layer0_outputs(2939));
    layer1_outputs(1535) <= (layer0_outputs(4433)) and not (layer0_outputs(2087));
    layer1_outputs(1536) <= (layer0_outputs(4657)) and not (layer0_outputs(2546));
    layer1_outputs(1537) <= '1';
    layer1_outputs(1538) <= not((layer0_outputs(4674)) or (layer0_outputs(111)));
    layer1_outputs(1539) <= not(layer0_outputs(2226));
    layer1_outputs(1540) <= not(layer0_outputs(4935)) or (layer0_outputs(7496));
    layer1_outputs(1541) <= not((layer0_outputs(9600)) or (layer0_outputs(8522)));
    layer1_outputs(1542) <= not(layer0_outputs(1253));
    layer1_outputs(1543) <= not(layer0_outputs(3036));
    layer1_outputs(1544) <= not((layer0_outputs(2619)) and (layer0_outputs(9696)));
    layer1_outputs(1545) <= not(layer0_outputs(33));
    layer1_outputs(1546) <= layer0_outputs(2157);
    layer1_outputs(1547) <= (layer0_outputs(1689)) and (layer0_outputs(6306));
    layer1_outputs(1548) <= not((layer0_outputs(958)) or (layer0_outputs(8647)));
    layer1_outputs(1549) <= not((layer0_outputs(2063)) or (layer0_outputs(8820)));
    layer1_outputs(1550) <= not(layer0_outputs(7937));
    layer1_outputs(1551) <= not((layer0_outputs(1127)) xor (layer0_outputs(5197)));
    layer1_outputs(1552) <= (layer0_outputs(469)) and not (layer0_outputs(50));
    layer1_outputs(1553) <= not(layer0_outputs(4079));
    layer1_outputs(1554) <= not((layer0_outputs(7779)) or (layer0_outputs(6091)));
    layer1_outputs(1555) <= not(layer0_outputs(1108)) or (layer0_outputs(3511));
    layer1_outputs(1556) <= not((layer0_outputs(3784)) and (layer0_outputs(1682)));
    layer1_outputs(1557) <= not(layer0_outputs(6453));
    layer1_outputs(1558) <= layer0_outputs(2242);
    layer1_outputs(1559) <= '1';
    layer1_outputs(1560) <= (layer0_outputs(9007)) xor (layer0_outputs(669));
    layer1_outputs(1561) <= not((layer0_outputs(9976)) or (layer0_outputs(4448)));
    layer1_outputs(1562) <= not((layer0_outputs(735)) xor (layer0_outputs(9543)));
    layer1_outputs(1563) <= layer0_outputs(1450);
    layer1_outputs(1564) <= layer0_outputs(1378);
    layer1_outputs(1565) <= not((layer0_outputs(8771)) and (layer0_outputs(5514)));
    layer1_outputs(1566) <= (layer0_outputs(4584)) and not (layer0_outputs(3803));
    layer1_outputs(1567) <= layer0_outputs(1788);
    layer1_outputs(1568) <= (layer0_outputs(6447)) xor (layer0_outputs(9255));
    layer1_outputs(1569) <= (layer0_outputs(8420)) or (layer0_outputs(4884));
    layer1_outputs(1570) <= (layer0_outputs(5839)) and not (layer0_outputs(8720));
    layer1_outputs(1571) <= layer0_outputs(4222);
    layer1_outputs(1572) <= layer0_outputs(10197);
    layer1_outputs(1573) <= not(layer0_outputs(8600)) or (layer0_outputs(10215));
    layer1_outputs(1574) <= not((layer0_outputs(9538)) and (layer0_outputs(8178)));
    layer1_outputs(1575) <= layer0_outputs(5178);
    layer1_outputs(1576) <= not((layer0_outputs(2767)) xor (layer0_outputs(9373)));
    layer1_outputs(1577) <= not(layer0_outputs(1405)) or (layer0_outputs(5130));
    layer1_outputs(1578) <= not((layer0_outputs(9364)) and (layer0_outputs(578)));
    layer1_outputs(1579) <= not(layer0_outputs(6376));
    layer1_outputs(1580) <= '1';
    layer1_outputs(1581) <= '1';
    layer1_outputs(1582) <= not(layer0_outputs(4209));
    layer1_outputs(1583) <= (layer0_outputs(1784)) and (layer0_outputs(9774));
    layer1_outputs(1584) <= not((layer0_outputs(9726)) xor (layer0_outputs(7526)));
    layer1_outputs(1585) <= not((layer0_outputs(9835)) xor (layer0_outputs(8232)));
    layer1_outputs(1586) <= (layer0_outputs(5398)) and not (layer0_outputs(3225));
    layer1_outputs(1587) <= not(layer0_outputs(8929));
    layer1_outputs(1588) <= '0';
    layer1_outputs(1589) <= not(layer0_outputs(10204));
    layer1_outputs(1590) <= not(layer0_outputs(5834)) or (layer0_outputs(1473));
    layer1_outputs(1591) <= (layer0_outputs(8204)) and not (layer0_outputs(3341));
    layer1_outputs(1592) <= not(layer0_outputs(8140)) or (layer0_outputs(4506));
    layer1_outputs(1593) <= layer0_outputs(7122);
    layer1_outputs(1594) <= not((layer0_outputs(9456)) and (layer0_outputs(3199)));
    layer1_outputs(1595) <= (layer0_outputs(9030)) or (layer0_outputs(365));
    layer1_outputs(1596) <= not((layer0_outputs(6665)) or (layer0_outputs(7092)));
    layer1_outputs(1597) <= (layer0_outputs(3463)) or (layer0_outputs(8713));
    layer1_outputs(1598) <= not((layer0_outputs(5592)) or (layer0_outputs(2072)));
    layer1_outputs(1599) <= (layer0_outputs(3167)) or (layer0_outputs(3118));
    layer1_outputs(1600) <= '1';
    layer1_outputs(1601) <= (layer0_outputs(5943)) and (layer0_outputs(3169));
    layer1_outputs(1602) <= (layer0_outputs(9176)) and not (layer0_outputs(3377));
    layer1_outputs(1603) <= not(layer0_outputs(6969)) or (layer0_outputs(9599));
    layer1_outputs(1604) <= (layer0_outputs(9962)) and (layer0_outputs(592));
    layer1_outputs(1605) <= layer0_outputs(4650);
    layer1_outputs(1606) <= not(layer0_outputs(227)) or (layer0_outputs(4379));
    layer1_outputs(1607) <= not((layer0_outputs(3569)) and (layer0_outputs(0)));
    layer1_outputs(1608) <= (layer0_outputs(8578)) xor (layer0_outputs(10232));
    layer1_outputs(1609) <= not((layer0_outputs(5928)) or (layer0_outputs(2023)));
    layer1_outputs(1610) <= not(layer0_outputs(2929));
    layer1_outputs(1611) <= layer0_outputs(1140);
    layer1_outputs(1612) <= layer0_outputs(5573);
    layer1_outputs(1613) <= not(layer0_outputs(10028)) or (layer0_outputs(10192));
    layer1_outputs(1614) <= not(layer0_outputs(2191));
    layer1_outputs(1615) <= layer0_outputs(4751);
    layer1_outputs(1616) <= layer0_outputs(3108);
    layer1_outputs(1617) <= not((layer0_outputs(4673)) or (layer0_outputs(10052)));
    layer1_outputs(1618) <= (layer0_outputs(1927)) or (layer0_outputs(4145));
    layer1_outputs(1619) <= (layer0_outputs(3117)) and (layer0_outputs(9340));
    layer1_outputs(1620) <= not(layer0_outputs(5231));
    layer1_outputs(1621) <= '1';
    layer1_outputs(1622) <= (layer0_outputs(6400)) or (layer0_outputs(5875));
    layer1_outputs(1623) <= not(layer0_outputs(6087));
    layer1_outputs(1624) <= (layer0_outputs(9615)) and (layer0_outputs(3871));
    layer1_outputs(1625) <= not(layer0_outputs(4992)) or (layer0_outputs(7864));
    layer1_outputs(1626) <= not(layer0_outputs(9516));
    layer1_outputs(1627) <= not(layer0_outputs(2492));
    layer1_outputs(1628) <= not(layer0_outputs(8504)) or (layer0_outputs(3362));
    layer1_outputs(1629) <= (layer0_outputs(1693)) and not (layer0_outputs(278));
    layer1_outputs(1630) <= layer0_outputs(2179);
    layer1_outputs(1631) <= layer0_outputs(9863);
    layer1_outputs(1632) <= layer0_outputs(6986);
    layer1_outputs(1633) <= not(layer0_outputs(3670));
    layer1_outputs(1634) <= (layer0_outputs(10103)) and not (layer0_outputs(8327));
    layer1_outputs(1635) <= '0';
    layer1_outputs(1636) <= not(layer0_outputs(5061)) or (layer0_outputs(5995));
    layer1_outputs(1637) <= not(layer0_outputs(3973));
    layer1_outputs(1638) <= (layer0_outputs(6912)) or (layer0_outputs(2354));
    layer1_outputs(1639) <= (layer0_outputs(7252)) and (layer0_outputs(1803));
    layer1_outputs(1640) <= (layer0_outputs(135)) and not (layer0_outputs(550));
    layer1_outputs(1641) <= not(layer0_outputs(2976));
    layer1_outputs(1642) <= (layer0_outputs(8859)) and not (layer0_outputs(10237));
    layer1_outputs(1643) <= not(layer0_outputs(4788));
    layer1_outputs(1644) <= (layer0_outputs(7141)) and not (layer0_outputs(3398));
    layer1_outputs(1645) <= not(layer0_outputs(2935));
    layer1_outputs(1646) <= not((layer0_outputs(5593)) or (layer0_outputs(9321)));
    layer1_outputs(1647) <= not((layer0_outputs(7909)) or (layer0_outputs(2884)));
    layer1_outputs(1648) <= layer0_outputs(3668);
    layer1_outputs(1649) <= (layer0_outputs(3075)) and not (layer0_outputs(7685));
    layer1_outputs(1650) <= '1';
    layer1_outputs(1651) <= (layer0_outputs(1989)) or (layer0_outputs(402));
    layer1_outputs(1652) <= (layer0_outputs(634)) and not (layer0_outputs(5822));
    layer1_outputs(1653) <= layer0_outputs(6972);
    layer1_outputs(1654) <= not(layer0_outputs(1975));
    layer1_outputs(1655) <= not(layer0_outputs(3411));
    layer1_outputs(1656) <= (layer0_outputs(10045)) and (layer0_outputs(10193));
    layer1_outputs(1657) <= layer0_outputs(4581);
    layer1_outputs(1658) <= not((layer0_outputs(158)) or (layer0_outputs(1950)));
    layer1_outputs(1659) <= '1';
    layer1_outputs(1660) <= layer0_outputs(1298);
    layer1_outputs(1661) <= not(layer0_outputs(3356));
    layer1_outputs(1662) <= layer0_outputs(7196);
    layer1_outputs(1663) <= layer0_outputs(2013);
    layer1_outputs(1664) <= (layer0_outputs(6260)) or (layer0_outputs(3592));
    layer1_outputs(1665) <= (layer0_outputs(6375)) and (layer0_outputs(69));
    layer1_outputs(1666) <= not(layer0_outputs(9802));
    layer1_outputs(1667) <= (layer0_outputs(8565)) and not (layer0_outputs(9745));
    layer1_outputs(1668) <= not((layer0_outputs(9163)) and (layer0_outputs(7867)));
    layer1_outputs(1669) <= not((layer0_outputs(1091)) xor (layer0_outputs(66)));
    layer1_outputs(1670) <= (layer0_outputs(791)) and not (layer0_outputs(7105));
    layer1_outputs(1671) <= not((layer0_outputs(6779)) or (layer0_outputs(9121)));
    layer1_outputs(1672) <= not(layer0_outputs(1821));
    layer1_outputs(1673) <= (layer0_outputs(459)) and not (layer0_outputs(6457));
    layer1_outputs(1674) <= '0';
    layer1_outputs(1675) <= '0';
    layer1_outputs(1676) <= layer0_outputs(5939);
    layer1_outputs(1677) <= not(layer0_outputs(4996)) or (layer0_outputs(5590));
    layer1_outputs(1678) <= not(layer0_outputs(4749)) or (layer0_outputs(758));
    layer1_outputs(1679) <= '0';
    layer1_outputs(1680) <= '0';
    layer1_outputs(1681) <= not((layer0_outputs(2785)) or (layer0_outputs(10210)));
    layer1_outputs(1682) <= layer0_outputs(6175);
    layer1_outputs(1683) <= not((layer0_outputs(9542)) or (layer0_outputs(10127)));
    layer1_outputs(1684) <= layer0_outputs(9725);
    layer1_outputs(1685) <= (layer0_outputs(3372)) and not (layer0_outputs(4454));
    layer1_outputs(1686) <= not((layer0_outputs(4675)) xor (layer0_outputs(3404)));
    layer1_outputs(1687) <= not((layer0_outputs(5041)) or (layer0_outputs(5677)));
    layer1_outputs(1688) <= (layer0_outputs(8068)) xor (layer0_outputs(10231));
    layer1_outputs(1689) <= '0';
    layer1_outputs(1690) <= layer0_outputs(6456);
    layer1_outputs(1691) <= (layer0_outputs(42)) and (layer0_outputs(7068));
    layer1_outputs(1692) <= layer0_outputs(9801);
    layer1_outputs(1693) <= '1';
    layer1_outputs(1694) <= (layer0_outputs(589)) xor (layer0_outputs(5346));
    layer1_outputs(1695) <= layer0_outputs(6968);
    layer1_outputs(1696) <= (layer0_outputs(3814)) and not (layer0_outputs(7853));
    layer1_outputs(1697) <= (layer0_outputs(510)) and not (layer0_outputs(5127));
    layer1_outputs(1698) <= layer0_outputs(2189);
    layer1_outputs(1699) <= (layer0_outputs(1744)) or (layer0_outputs(7694));
    layer1_outputs(1700) <= '1';
    layer1_outputs(1701) <= '1';
    layer1_outputs(1702) <= '0';
    layer1_outputs(1703) <= layer0_outputs(5784);
    layer1_outputs(1704) <= layer0_outputs(560);
    layer1_outputs(1705) <= not(layer0_outputs(1272));
    layer1_outputs(1706) <= layer0_outputs(788);
    layer1_outputs(1707) <= not(layer0_outputs(9497));
    layer1_outputs(1708) <= layer0_outputs(1296);
    layer1_outputs(1709) <= (layer0_outputs(1852)) and not (layer0_outputs(4328));
    layer1_outputs(1710) <= layer0_outputs(5387);
    layer1_outputs(1711) <= '1';
    layer1_outputs(1712) <= '1';
    layer1_outputs(1713) <= not(layer0_outputs(194));
    layer1_outputs(1714) <= (layer0_outputs(1275)) and not (layer0_outputs(625));
    layer1_outputs(1715) <= not(layer0_outputs(6552));
    layer1_outputs(1716) <= layer0_outputs(9850);
    layer1_outputs(1717) <= (layer0_outputs(1975)) and (layer0_outputs(4134));
    layer1_outputs(1718) <= not(layer0_outputs(78));
    layer1_outputs(1719) <= layer0_outputs(10003);
    layer1_outputs(1720) <= not((layer0_outputs(6476)) xor (layer0_outputs(670)));
    layer1_outputs(1721) <= not(layer0_outputs(1242));
    layer1_outputs(1722) <= layer0_outputs(295);
    layer1_outputs(1723) <= not(layer0_outputs(6624)) or (layer0_outputs(2730));
    layer1_outputs(1724) <= layer0_outputs(5147);
    layer1_outputs(1725) <= not((layer0_outputs(1671)) and (layer0_outputs(704)));
    layer1_outputs(1726) <= not(layer0_outputs(8557)) or (layer0_outputs(547));
    layer1_outputs(1727) <= layer0_outputs(9170);
    layer1_outputs(1728) <= (layer0_outputs(4210)) and not (layer0_outputs(2465));
    layer1_outputs(1729) <= layer0_outputs(4504);
    layer1_outputs(1730) <= not(layer0_outputs(5918));
    layer1_outputs(1731) <= layer0_outputs(6545);
    layer1_outputs(1732) <= '0';
    layer1_outputs(1733) <= (layer0_outputs(8037)) xor (layer0_outputs(4436));
    layer1_outputs(1734) <= not(layer0_outputs(5690));
    layer1_outputs(1735) <= (layer0_outputs(9248)) and not (layer0_outputs(3001));
    layer1_outputs(1736) <= not(layer0_outputs(4490));
    layer1_outputs(1737) <= (layer0_outputs(388)) xor (layer0_outputs(2059));
    layer1_outputs(1738) <= (layer0_outputs(1596)) and not (layer0_outputs(6756));
    layer1_outputs(1739) <= not((layer0_outputs(363)) and (layer0_outputs(5845)));
    layer1_outputs(1740) <= not(layer0_outputs(5668));
    layer1_outputs(1741) <= layer0_outputs(6242);
    layer1_outputs(1742) <= (layer0_outputs(4690)) and not (layer0_outputs(4290));
    layer1_outputs(1743) <= not((layer0_outputs(6318)) and (layer0_outputs(4501)));
    layer1_outputs(1744) <= layer0_outputs(4768);
    layer1_outputs(1745) <= '1';
    layer1_outputs(1746) <= (layer0_outputs(3288)) and (layer0_outputs(3092));
    layer1_outputs(1747) <= layer0_outputs(3413);
    layer1_outputs(1748) <= '1';
    layer1_outputs(1749) <= (layer0_outputs(9421)) and not (layer0_outputs(8701));
    layer1_outputs(1750) <= (layer0_outputs(4158)) and (layer0_outputs(4432));
    layer1_outputs(1751) <= (layer0_outputs(6121)) and not (layer0_outputs(3795));
    layer1_outputs(1752) <= (layer0_outputs(6380)) or (layer0_outputs(2601));
    layer1_outputs(1753) <= not(layer0_outputs(1235));
    layer1_outputs(1754) <= '0';
    layer1_outputs(1755) <= not(layer0_outputs(2214));
    layer1_outputs(1756) <= not(layer0_outputs(7075)) or (layer0_outputs(1554));
    layer1_outputs(1757) <= (layer0_outputs(1913)) or (layer0_outputs(4350));
    layer1_outputs(1758) <= not(layer0_outputs(7675));
    layer1_outputs(1759) <= not(layer0_outputs(4241));
    layer1_outputs(1760) <= not((layer0_outputs(6005)) and (layer0_outputs(5522)));
    layer1_outputs(1761) <= not(layer0_outputs(1915));
    layer1_outputs(1762) <= not((layer0_outputs(589)) xor (layer0_outputs(4180)));
    layer1_outputs(1763) <= not((layer0_outputs(3385)) and (layer0_outputs(7795)));
    layer1_outputs(1764) <= '1';
    layer1_outputs(1765) <= (layer0_outputs(2159)) or (layer0_outputs(1260));
    layer1_outputs(1766) <= not(layer0_outputs(1837)) or (layer0_outputs(9874));
    layer1_outputs(1767) <= not(layer0_outputs(9022)) or (layer0_outputs(6664));
    layer1_outputs(1768) <= '0';
    layer1_outputs(1769) <= (layer0_outputs(8034)) xor (layer0_outputs(2948));
    layer1_outputs(1770) <= not(layer0_outputs(123)) or (layer0_outputs(344));
    layer1_outputs(1771) <= not((layer0_outputs(9902)) and (layer0_outputs(6191)));
    layer1_outputs(1772) <= not((layer0_outputs(7546)) and (layer0_outputs(215)));
    layer1_outputs(1773) <= layer0_outputs(6880);
    layer1_outputs(1774) <= (layer0_outputs(3481)) and not (layer0_outputs(1854));
    layer1_outputs(1775) <= '0';
    layer1_outputs(1776) <= not((layer0_outputs(6766)) xor (layer0_outputs(7612)));
    layer1_outputs(1777) <= (layer0_outputs(7570)) and (layer0_outputs(7197));
    layer1_outputs(1778) <= layer0_outputs(5868);
    layer1_outputs(1779) <= not((layer0_outputs(5403)) or (layer0_outputs(4900)));
    layer1_outputs(1780) <= not(layer0_outputs(6092)) or (layer0_outputs(535));
    layer1_outputs(1781) <= (layer0_outputs(9293)) and (layer0_outputs(8328));
    layer1_outputs(1782) <= not((layer0_outputs(7482)) or (layer0_outputs(7278)));
    layer1_outputs(1783) <= not((layer0_outputs(2820)) xor (layer0_outputs(5064)));
    layer1_outputs(1784) <= '1';
    layer1_outputs(1785) <= not(layer0_outputs(939)) or (layer0_outputs(7722));
    layer1_outputs(1786) <= not(layer0_outputs(7972));
    layer1_outputs(1787) <= layer0_outputs(7781);
    layer1_outputs(1788) <= not(layer0_outputs(2012)) or (layer0_outputs(2153));
    layer1_outputs(1789) <= (layer0_outputs(2214)) and not (layer0_outputs(2534));
    layer1_outputs(1790) <= not(layer0_outputs(6976));
    layer1_outputs(1791) <= not(layer0_outputs(3321));
    layer1_outputs(1792) <= (layer0_outputs(552)) and not (layer0_outputs(8125));
    layer1_outputs(1793) <= not((layer0_outputs(6391)) and (layer0_outputs(5639)));
    layer1_outputs(1794) <= layer0_outputs(8284);
    layer1_outputs(1795) <= not((layer0_outputs(8601)) and (layer0_outputs(2238)));
    layer1_outputs(1796) <= not((layer0_outputs(9960)) xor (layer0_outputs(6855)));
    layer1_outputs(1797) <= not((layer0_outputs(7846)) and (layer0_outputs(5701)));
    layer1_outputs(1798) <= not(layer0_outputs(3765));
    layer1_outputs(1799) <= (layer0_outputs(748)) and not (layer0_outputs(6095));
    layer1_outputs(1800) <= not(layer0_outputs(8176)) or (layer0_outputs(9813));
    layer1_outputs(1801) <= (layer0_outputs(4428)) and not (layer0_outputs(729));
    layer1_outputs(1802) <= not((layer0_outputs(6083)) or (layer0_outputs(7748)));
    layer1_outputs(1803) <= not(layer0_outputs(7921)) or (layer0_outputs(370));
    layer1_outputs(1804) <= not(layer0_outputs(9920)) or (layer0_outputs(7747));
    layer1_outputs(1805) <= layer0_outputs(8992);
    layer1_outputs(1806) <= (layer0_outputs(2607)) xor (layer0_outputs(6517));
    layer1_outputs(1807) <= layer0_outputs(9076);
    layer1_outputs(1808) <= not(layer0_outputs(1728));
    layer1_outputs(1809) <= layer0_outputs(5857);
    layer1_outputs(1810) <= (layer0_outputs(8072)) and not (layer0_outputs(6939));
    layer1_outputs(1811) <= not((layer0_outputs(4336)) and (layer0_outputs(6697)));
    layer1_outputs(1812) <= not(layer0_outputs(5388));
    layer1_outputs(1813) <= '0';
    layer1_outputs(1814) <= not(layer0_outputs(9458));
    layer1_outputs(1815) <= (layer0_outputs(1845)) and not (layer0_outputs(9298));
    layer1_outputs(1816) <= not(layer0_outputs(7775)) or (layer0_outputs(7714));
    layer1_outputs(1817) <= (layer0_outputs(1001)) or (layer0_outputs(851));
    layer1_outputs(1818) <= not((layer0_outputs(3488)) and (layer0_outputs(10033)));
    layer1_outputs(1819) <= not(layer0_outputs(3638)) or (layer0_outputs(4723));
    layer1_outputs(1820) <= not((layer0_outputs(6092)) and (layer0_outputs(2641)));
    layer1_outputs(1821) <= not(layer0_outputs(3289)) or (layer0_outputs(1607));
    layer1_outputs(1822) <= (layer0_outputs(8154)) or (layer0_outputs(4075));
    layer1_outputs(1823) <= not((layer0_outputs(3901)) or (layer0_outputs(1640)));
    layer1_outputs(1824) <= layer0_outputs(6180);
    layer1_outputs(1825) <= (layer0_outputs(2557)) and (layer0_outputs(272));
    layer1_outputs(1826) <= (layer0_outputs(3576)) and (layer0_outputs(1817));
    layer1_outputs(1827) <= layer0_outputs(4593);
    layer1_outputs(1828) <= (layer0_outputs(8642)) or (layer0_outputs(136));
    layer1_outputs(1829) <= (layer0_outputs(3698)) or (layer0_outputs(299));
    layer1_outputs(1830) <= (layer0_outputs(624)) and not (layer0_outputs(4813));
    layer1_outputs(1831) <= (layer0_outputs(2717)) or (layer0_outputs(4145));
    layer1_outputs(1832) <= (layer0_outputs(19)) and not (layer0_outputs(5049));
    layer1_outputs(1833) <= '1';
    layer1_outputs(1834) <= layer0_outputs(1933);
    layer1_outputs(1835) <= not(layer0_outputs(3286)) or (layer0_outputs(372));
    layer1_outputs(1836) <= layer0_outputs(76);
    layer1_outputs(1837) <= not(layer0_outputs(2185));
    layer1_outputs(1838) <= (layer0_outputs(4924)) and (layer0_outputs(6882));
    layer1_outputs(1839) <= not((layer0_outputs(7994)) xor (layer0_outputs(443)));
    layer1_outputs(1840) <= (layer0_outputs(979)) or (layer0_outputs(3712));
    layer1_outputs(1841) <= (layer0_outputs(63)) and not (layer0_outputs(4319));
    layer1_outputs(1842) <= '1';
    layer1_outputs(1843) <= layer0_outputs(6668);
    layer1_outputs(1844) <= not((layer0_outputs(8229)) or (layer0_outputs(8307)));
    layer1_outputs(1845) <= not(layer0_outputs(5695)) or (layer0_outputs(2501));
    layer1_outputs(1846) <= not(layer0_outputs(5183));
    layer1_outputs(1847) <= (layer0_outputs(2997)) or (layer0_outputs(3124));
    layer1_outputs(1848) <= (layer0_outputs(189)) xor (layer0_outputs(5805));
    layer1_outputs(1849) <= layer0_outputs(1154);
    layer1_outputs(1850) <= not(layer0_outputs(9276));
    layer1_outputs(1851) <= layer0_outputs(1211);
    layer1_outputs(1852) <= not(layer0_outputs(182)) or (layer0_outputs(380));
    layer1_outputs(1853) <= layer0_outputs(1212);
    layer1_outputs(1854) <= not((layer0_outputs(2151)) and (layer0_outputs(947)));
    layer1_outputs(1855) <= (layer0_outputs(9401)) and (layer0_outputs(2126));
    layer1_outputs(1856) <= (layer0_outputs(667)) or (layer0_outputs(1312));
    layer1_outputs(1857) <= (layer0_outputs(8082)) and not (layer0_outputs(1688));
    layer1_outputs(1858) <= (layer0_outputs(1616)) or (layer0_outputs(9148));
    layer1_outputs(1859) <= layer0_outputs(8207);
    layer1_outputs(1860) <= not(layer0_outputs(5238));
    layer1_outputs(1861) <= (layer0_outputs(6430)) or (layer0_outputs(4715));
    layer1_outputs(1862) <= layer0_outputs(4767);
    layer1_outputs(1863) <= not(layer0_outputs(9483)) or (layer0_outputs(1283));
    layer1_outputs(1864) <= not((layer0_outputs(4661)) xor (layer0_outputs(4146)));
    layer1_outputs(1865) <= (layer0_outputs(9362)) or (layer0_outputs(2740));
    layer1_outputs(1866) <= '1';
    layer1_outputs(1867) <= not(layer0_outputs(4363));
    layer1_outputs(1868) <= not(layer0_outputs(1659));
    layer1_outputs(1869) <= (layer0_outputs(7438)) and not (layer0_outputs(431));
    layer1_outputs(1870) <= not((layer0_outputs(10163)) xor (layer0_outputs(8018)));
    layer1_outputs(1871) <= layer0_outputs(569);
    layer1_outputs(1872) <= layer0_outputs(7019);
    layer1_outputs(1873) <= (layer0_outputs(5592)) and not (layer0_outputs(9384));
    layer1_outputs(1874) <= not(layer0_outputs(2323));
    layer1_outputs(1875) <= not(layer0_outputs(5025));
    layer1_outputs(1876) <= (layer0_outputs(3095)) or (layer0_outputs(5579));
    layer1_outputs(1877) <= not(layer0_outputs(8702)) or (layer0_outputs(4251));
    layer1_outputs(1878) <= (layer0_outputs(2689)) xor (layer0_outputs(9019));
    layer1_outputs(1879) <= not(layer0_outputs(2258));
    layer1_outputs(1880) <= (layer0_outputs(1278)) and not (layer0_outputs(1609));
    layer1_outputs(1881) <= not(layer0_outputs(6781)) or (layer0_outputs(1113));
    layer1_outputs(1882) <= not((layer0_outputs(8007)) xor (layer0_outputs(921)));
    layer1_outputs(1883) <= not((layer0_outputs(2025)) xor (layer0_outputs(9660)));
    layer1_outputs(1884) <= layer0_outputs(7178);
    layer1_outputs(1885) <= layer0_outputs(2468);
    layer1_outputs(1886) <= not((layer0_outputs(2850)) and (layer0_outputs(3577)));
    layer1_outputs(1887) <= (layer0_outputs(6592)) and not (layer0_outputs(7883));
    layer1_outputs(1888) <= (layer0_outputs(9908)) and (layer0_outputs(113));
    layer1_outputs(1889) <= (layer0_outputs(9090)) xor (layer0_outputs(6951));
    layer1_outputs(1890) <= not((layer0_outputs(8184)) xor (layer0_outputs(9701)));
    layer1_outputs(1891) <= not(layer0_outputs(10202));
    layer1_outputs(1892) <= (layer0_outputs(9893)) or (layer0_outputs(430));
    layer1_outputs(1893) <= (layer0_outputs(8324)) or (layer0_outputs(3298));
    layer1_outputs(1894) <= not(layer0_outputs(5733)) or (layer0_outputs(2660));
    layer1_outputs(1895) <= (layer0_outputs(8221)) and not (layer0_outputs(1466));
    layer1_outputs(1896) <= not(layer0_outputs(6506)) or (layer0_outputs(922));
    layer1_outputs(1897) <= (layer0_outputs(5897)) or (layer0_outputs(1786));
    layer1_outputs(1898) <= (layer0_outputs(52)) and not (layer0_outputs(5047));
    layer1_outputs(1899) <= not(layer0_outputs(1113)) or (layer0_outputs(7171));
    layer1_outputs(1900) <= (layer0_outputs(850)) and (layer0_outputs(7058));
    layer1_outputs(1901) <= not(layer0_outputs(1641));
    layer1_outputs(1902) <= not((layer0_outputs(9950)) xor (layer0_outputs(10152)));
    layer1_outputs(1903) <= not(layer0_outputs(179));
    layer1_outputs(1904) <= (layer0_outputs(10100)) or (layer0_outputs(2745));
    layer1_outputs(1905) <= not((layer0_outputs(3981)) or (layer0_outputs(2696)));
    layer1_outputs(1906) <= not(layer0_outputs(2489));
    layer1_outputs(1907) <= layer0_outputs(854);
    layer1_outputs(1908) <= (layer0_outputs(4619)) and (layer0_outputs(8895));
    layer1_outputs(1909) <= not(layer0_outputs(4192));
    layer1_outputs(1910) <= not((layer0_outputs(7990)) xor (layer0_outputs(8717)));
    layer1_outputs(1911) <= not(layer0_outputs(3563));
    layer1_outputs(1912) <= not(layer0_outputs(3754)) or (layer0_outputs(2519));
    layer1_outputs(1913) <= not((layer0_outputs(2544)) and (layer0_outputs(8370)));
    layer1_outputs(1914) <= not(layer0_outputs(8754)) or (layer0_outputs(2410));
    layer1_outputs(1915) <= '0';
    layer1_outputs(1916) <= (layer0_outputs(6481)) and not (layer0_outputs(2985));
    layer1_outputs(1917) <= (layer0_outputs(9986)) and (layer0_outputs(8939));
    layer1_outputs(1918) <= (layer0_outputs(10160)) and (layer0_outputs(878));
    layer1_outputs(1919) <= not(layer0_outputs(6267));
    layer1_outputs(1920) <= '0';
    layer1_outputs(1921) <= not(layer0_outputs(4149));
    layer1_outputs(1922) <= layer0_outputs(4853);
    layer1_outputs(1923) <= layer0_outputs(1262);
    layer1_outputs(1924) <= not(layer0_outputs(4043)) or (layer0_outputs(7593));
    layer1_outputs(1925) <= not(layer0_outputs(893));
    layer1_outputs(1926) <= '0';
    layer1_outputs(1927) <= not(layer0_outputs(5805)) or (layer0_outputs(5258));
    layer1_outputs(1928) <= layer0_outputs(3476);
    layer1_outputs(1929) <= (layer0_outputs(1502)) and not (layer0_outputs(947));
    layer1_outputs(1930) <= not((layer0_outputs(9947)) and (layer0_outputs(7199)));
    layer1_outputs(1931) <= layer0_outputs(7080);
    layer1_outputs(1932) <= (layer0_outputs(5842)) and not (layer0_outputs(769));
    layer1_outputs(1933) <= not(layer0_outputs(2221)) or (layer0_outputs(9884));
    layer1_outputs(1934) <= (layer0_outputs(9729)) and not (layer0_outputs(2767));
    layer1_outputs(1935) <= layer0_outputs(7794);
    layer1_outputs(1936) <= not(layer0_outputs(34)) or (layer0_outputs(1034));
    layer1_outputs(1937) <= not(layer0_outputs(2661)) or (layer0_outputs(7607));
    layer1_outputs(1938) <= layer0_outputs(856);
    layer1_outputs(1939) <= not((layer0_outputs(1944)) and (layer0_outputs(317)));
    layer1_outputs(1940) <= not(layer0_outputs(8159)) or (layer0_outputs(497));
    layer1_outputs(1941) <= '1';
    layer1_outputs(1942) <= (layer0_outputs(8170)) or (layer0_outputs(8167));
    layer1_outputs(1943) <= layer0_outputs(1421);
    layer1_outputs(1944) <= not(layer0_outputs(4235));
    layer1_outputs(1945) <= layer0_outputs(5062);
    layer1_outputs(1946) <= not(layer0_outputs(3135)) or (layer0_outputs(3959));
    layer1_outputs(1947) <= layer0_outputs(3755);
    layer1_outputs(1948) <= (layer0_outputs(9316)) and (layer0_outputs(8481));
    layer1_outputs(1949) <= '1';
    layer1_outputs(1950) <= not((layer0_outputs(1832)) or (layer0_outputs(1644)));
    layer1_outputs(1951) <= not(layer0_outputs(3825));
    layer1_outputs(1952) <= layer0_outputs(2528);
    layer1_outputs(1953) <= not(layer0_outputs(747));
    layer1_outputs(1954) <= not((layer0_outputs(6450)) or (layer0_outputs(7975)));
    layer1_outputs(1955) <= '0';
    layer1_outputs(1956) <= not(layer0_outputs(6001));
    layer1_outputs(1957) <= not(layer0_outputs(6920));
    layer1_outputs(1958) <= layer0_outputs(715);
    layer1_outputs(1959) <= layer0_outputs(6495);
    layer1_outputs(1960) <= not(layer0_outputs(690)) or (layer0_outputs(8412));
    layer1_outputs(1961) <= not((layer0_outputs(6689)) and (layer0_outputs(8747)));
    layer1_outputs(1962) <= not(layer0_outputs(3440));
    layer1_outputs(1963) <= not((layer0_outputs(21)) or (layer0_outputs(8471)));
    layer1_outputs(1964) <= not((layer0_outputs(1374)) and (layer0_outputs(2992)));
    layer1_outputs(1965) <= (layer0_outputs(5322)) and not (layer0_outputs(3184));
    layer1_outputs(1966) <= not(layer0_outputs(7460)) or (layer0_outputs(2083));
    layer1_outputs(1967) <= not(layer0_outputs(608)) or (layer0_outputs(4600));
    layer1_outputs(1968) <= not(layer0_outputs(2572)) or (layer0_outputs(9536));
    layer1_outputs(1969) <= not(layer0_outputs(945));
    layer1_outputs(1970) <= layer0_outputs(3781);
    layer1_outputs(1971) <= (layer0_outputs(2030)) or (layer0_outputs(7274));
    layer1_outputs(1972) <= not(layer0_outputs(10104)) or (layer0_outputs(9717));
    layer1_outputs(1973) <= not((layer0_outputs(2138)) or (layer0_outputs(2522)));
    layer1_outputs(1974) <= (layer0_outputs(191)) and (layer0_outputs(2679));
    layer1_outputs(1975) <= (layer0_outputs(7301)) and (layer0_outputs(4560));
    layer1_outputs(1976) <= layer0_outputs(9877);
    layer1_outputs(1977) <= layer0_outputs(7636);
    layer1_outputs(1978) <= (layer0_outputs(7947)) xor (layer0_outputs(949));
    layer1_outputs(1979) <= '1';
    layer1_outputs(1980) <= (layer0_outputs(9843)) and not (layer0_outputs(8025));
    layer1_outputs(1981) <= not(layer0_outputs(263)) or (layer0_outputs(3058));
    layer1_outputs(1982) <= not(layer0_outputs(9375));
    layer1_outputs(1983) <= not(layer0_outputs(5950)) or (layer0_outputs(1262));
    layer1_outputs(1984) <= '1';
    layer1_outputs(1985) <= layer0_outputs(1808);
    layer1_outputs(1986) <= not(layer0_outputs(7074)) or (layer0_outputs(1851));
    layer1_outputs(1987) <= not((layer0_outputs(2777)) xor (layer0_outputs(8073)));
    layer1_outputs(1988) <= layer0_outputs(2299);
    layer1_outputs(1989) <= not((layer0_outputs(4142)) or (layer0_outputs(5143)));
    layer1_outputs(1990) <= layer0_outputs(9504);
    layer1_outputs(1991) <= not(layer0_outputs(4102)) or (layer0_outputs(3671));
    layer1_outputs(1992) <= (layer0_outputs(6199)) or (layer0_outputs(4665));
    layer1_outputs(1993) <= '0';
    layer1_outputs(1994) <= layer0_outputs(4720);
    layer1_outputs(1995) <= not(layer0_outputs(8383)) or (layer0_outputs(7082));
    layer1_outputs(1996) <= not(layer0_outputs(7515)) or (layer0_outputs(9174));
    layer1_outputs(1997) <= (layer0_outputs(7243)) or (layer0_outputs(671));
    layer1_outputs(1998) <= layer0_outputs(858);
    layer1_outputs(1999) <= layer0_outputs(1176);
    layer1_outputs(2000) <= layer0_outputs(4407);
    layer1_outputs(2001) <= (layer0_outputs(7821)) or (layer0_outputs(10145));
    layer1_outputs(2002) <= not((layer0_outputs(8922)) xor (layer0_outputs(8195)));
    layer1_outputs(2003) <= (layer0_outputs(842)) and not (layer0_outputs(5105));
    layer1_outputs(2004) <= layer0_outputs(7812);
    layer1_outputs(2005) <= not((layer0_outputs(4794)) or (layer0_outputs(8142)));
    layer1_outputs(2006) <= not(layer0_outputs(159)) or (layer0_outputs(9437));
    layer1_outputs(2007) <= not(layer0_outputs(8427)) or (layer0_outputs(3912));
    layer1_outputs(2008) <= layer0_outputs(9930);
    layer1_outputs(2009) <= not(layer0_outputs(5202));
    layer1_outputs(2010) <= '1';
    layer1_outputs(2011) <= layer0_outputs(7635);
    layer1_outputs(2012) <= not((layer0_outputs(3310)) or (layer0_outputs(2968)));
    layer1_outputs(2013) <= not(layer0_outputs(6589));
    layer1_outputs(2014) <= (layer0_outputs(9604)) xor (layer0_outputs(3924));
    layer1_outputs(2015) <= layer0_outputs(3577);
    layer1_outputs(2016) <= not((layer0_outputs(1372)) xor (layer0_outputs(4748)));
    layer1_outputs(2017) <= layer0_outputs(8886);
    layer1_outputs(2018) <= not(layer0_outputs(4558)) or (layer0_outputs(5523));
    layer1_outputs(2019) <= (layer0_outputs(2122)) and not (layer0_outputs(5505));
    layer1_outputs(2020) <= (layer0_outputs(7498)) or (layer0_outputs(8530));
    layer1_outputs(2021) <= (layer0_outputs(1027)) and (layer0_outputs(5091));
    layer1_outputs(2022) <= layer0_outputs(4107);
    layer1_outputs(2023) <= layer0_outputs(9143);
    layer1_outputs(2024) <= (layer0_outputs(4480)) and not (layer0_outputs(154));
    layer1_outputs(2025) <= (layer0_outputs(3416)) and not (layer0_outputs(200));
    layer1_outputs(2026) <= '0';
    layer1_outputs(2027) <= '0';
    layer1_outputs(2028) <= not((layer0_outputs(2792)) or (layer0_outputs(6262)));
    layer1_outputs(2029) <= layer0_outputs(855);
    layer1_outputs(2030) <= not((layer0_outputs(5567)) or (layer0_outputs(5195)));
    layer1_outputs(2031) <= not(layer0_outputs(646));
    layer1_outputs(2032) <= '1';
    layer1_outputs(2033) <= not(layer0_outputs(7844));
    layer1_outputs(2034) <= (layer0_outputs(9841)) xor (layer0_outputs(3019));
    layer1_outputs(2035) <= layer0_outputs(118);
    layer1_outputs(2036) <= (layer0_outputs(2021)) and not (layer0_outputs(7791));
    layer1_outputs(2037) <= not((layer0_outputs(1495)) and (layer0_outputs(238)));
    layer1_outputs(2038) <= (layer0_outputs(3656)) and (layer0_outputs(2110));
    layer1_outputs(2039) <= (layer0_outputs(1009)) and not (layer0_outputs(6594));
    layer1_outputs(2040) <= layer0_outputs(10118);
    layer1_outputs(2041) <= not(layer0_outputs(8790)) or (layer0_outputs(3817));
    layer1_outputs(2042) <= (layer0_outputs(9520)) xor (layer0_outputs(9432));
    layer1_outputs(2043) <= (layer0_outputs(7695)) and not (layer0_outputs(8844));
    layer1_outputs(2044) <= (layer0_outputs(7101)) xor (layer0_outputs(1303));
    layer1_outputs(2045) <= not(layer0_outputs(3109));
    layer1_outputs(2046) <= '0';
    layer1_outputs(2047) <= not(layer0_outputs(6867));
    layer1_outputs(2048) <= (layer0_outputs(2278)) and (layer0_outputs(5810));
    layer1_outputs(2049) <= not(layer0_outputs(3112));
    layer1_outputs(2050) <= layer0_outputs(595);
    layer1_outputs(2051) <= layer0_outputs(1579);
    layer1_outputs(2052) <= (layer0_outputs(183)) and not (layer0_outputs(10142));
    layer1_outputs(2053) <= layer0_outputs(2293);
    layer1_outputs(2054) <= '0';
    layer1_outputs(2055) <= layer0_outputs(3697);
    layer1_outputs(2056) <= (layer0_outputs(3821)) and not (layer0_outputs(559));
    layer1_outputs(2057) <= not((layer0_outputs(8952)) or (layer0_outputs(8312)));
    layer1_outputs(2058) <= layer0_outputs(6310);
    layer1_outputs(2059) <= not(layer0_outputs(89));
    layer1_outputs(2060) <= not(layer0_outputs(9342)) or (layer0_outputs(244));
    layer1_outputs(2061) <= '1';
    layer1_outputs(2062) <= (layer0_outputs(6507)) and not (layer0_outputs(4047));
    layer1_outputs(2063) <= not(layer0_outputs(4014));
    layer1_outputs(2064) <= layer0_outputs(4647);
    layer1_outputs(2065) <= not((layer0_outputs(1074)) xor (layer0_outputs(4849)));
    layer1_outputs(2066) <= not((layer0_outputs(6554)) or (layer0_outputs(9979)));
    layer1_outputs(2067) <= (layer0_outputs(7013)) and (layer0_outputs(7003));
    layer1_outputs(2068) <= not((layer0_outputs(8073)) and (layer0_outputs(4116)));
    layer1_outputs(2069) <= not((layer0_outputs(8992)) and (layer0_outputs(7686)));
    layer1_outputs(2070) <= '0';
    layer1_outputs(2071) <= (layer0_outputs(2326)) and (layer0_outputs(4947));
    layer1_outputs(2072) <= layer0_outputs(2427);
    layer1_outputs(2073) <= not(layer0_outputs(2077)) or (layer0_outputs(7512));
    layer1_outputs(2074) <= not((layer0_outputs(10229)) or (layer0_outputs(326)));
    layer1_outputs(2075) <= not((layer0_outputs(8260)) and (layer0_outputs(1311)));
    layer1_outputs(2076) <= layer0_outputs(2762);
    layer1_outputs(2077) <= (layer0_outputs(2299)) and not (layer0_outputs(9021));
    layer1_outputs(2078) <= '0';
    layer1_outputs(2079) <= '0';
    layer1_outputs(2080) <= (layer0_outputs(9101)) or (layer0_outputs(1541));
    layer1_outputs(2081) <= layer0_outputs(4697);
    layer1_outputs(2082) <= not(layer0_outputs(4541));
    layer1_outputs(2083) <= not(layer0_outputs(6134)) or (layer0_outputs(4211));
    layer1_outputs(2084) <= (layer0_outputs(1527)) or (layer0_outputs(5551));
    layer1_outputs(2085) <= '0';
    layer1_outputs(2086) <= (layer0_outputs(735)) and not (layer0_outputs(7057));
    layer1_outputs(2087) <= layer0_outputs(9526);
    layer1_outputs(2088) <= (layer0_outputs(5787)) and not (layer0_outputs(870));
    layer1_outputs(2089) <= not(layer0_outputs(3235));
    layer1_outputs(2090) <= '1';
    layer1_outputs(2091) <= (layer0_outputs(6117)) and not (layer0_outputs(4836));
    layer1_outputs(2092) <= layer0_outputs(3729);
    layer1_outputs(2093) <= '0';
    layer1_outputs(2094) <= layer0_outputs(4764);
    layer1_outputs(2095) <= not(layer0_outputs(6662));
    layer1_outputs(2096) <= not(layer0_outputs(2761)) or (layer0_outputs(6616));
    layer1_outputs(2097) <= layer0_outputs(2090);
    layer1_outputs(2098) <= not((layer0_outputs(6333)) and (layer0_outputs(1603)));
    layer1_outputs(2099) <= not(layer0_outputs(8693)) or (layer0_outputs(4222));
    layer1_outputs(2100) <= not((layer0_outputs(6874)) xor (layer0_outputs(9373)));
    layer1_outputs(2101) <= '0';
    layer1_outputs(2102) <= not(layer0_outputs(577));
    layer1_outputs(2103) <= (layer0_outputs(8856)) and (layer0_outputs(412));
    layer1_outputs(2104) <= layer0_outputs(5144);
    layer1_outputs(2105) <= not(layer0_outputs(6111));
    layer1_outputs(2106) <= '1';
    layer1_outputs(2107) <= not(layer0_outputs(7624)) or (layer0_outputs(1840));
    layer1_outputs(2108) <= (layer0_outputs(8408)) xor (layer0_outputs(8732));
    layer1_outputs(2109) <= not((layer0_outputs(4345)) xor (layer0_outputs(2598)));
    layer1_outputs(2110) <= '0';
    layer1_outputs(2111) <= (layer0_outputs(9907)) and (layer0_outputs(4220));
    layer1_outputs(2112) <= not((layer0_outputs(1834)) or (layer0_outputs(2158)));
    layer1_outputs(2113) <= '1';
    layer1_outputs(2114) <= (layer0_outputs(1110)) and not (layer0_outputs(7941));
    layer1_outputs(2115) <= '0';
    layer1_outputs(2116) <= (layer0_outputs(2340)) and (layer0_outputs(2849));
    layer1_outputs(2117) <= layer0_outputs(8344);
    layer1_outputs(2118) <= not(layer0_outputs(4574));
    layer1_outputs(2119) <= not(layer0_outputs(8009)) or (layer0_outputs(5402));
    layer1_outputs(2120) <= (layer0_outputs(3530)) or (layer0_outputs(6200));
    layer1_outputs(2121) <= not(layer0_outputs(8582));
    layer1_outputs(2122) <= (layer0_outputs(786)) and not (layer0_outputs(691));
    layer1_outputs(2123) <= not(layer0_outputs(1872)) or (layer0_outputs(2419));
    layer1_outputs(2124) <= layer0_outputs(3879);
    layer1_outputs(2125) <= layer0_outputs(4285);
    layer1_outputs(2126) <= (layer0_outputs(6640)) xor (layer0_outputs(1309));
    layer1_outputs(2127) <= not((layer0_outputs(10201)) and (layer0_outputs(820)));
    layer1_outputs(2128) <= layer0_outputs(6675);
    layer1_outputs(2129) <= not(layer0_outputs(4198));
    layer1_outputs(2130) <= layer0_outputs(835);
    layer1_outputs(2131) <= (layer0_outputs(3658)) and not (layer0_outputs(541));
    layer1_outputs(2132) <= '0';
    layer1_outputs(2133) <= not((layer0_outputs(342)) or (layer0_outputs(5296)));
    layer1_outputs(2134) <= (layer0_outputs(6775)) and (layer0_outputs(7531));
    layer1_outputs(2135) <= layer0_outputs(5168);
    layer1_outputs(2136) <= (layer0_outputs(4940)) or (layer0_outputs(3549));
    layer1_outputs(2137) <= (layer0_outputs(5487)) and not (layer0_outputs(1467));
    layer1_outputs(2138) <= layer0_outputs(6268);
    layer1_outputs(2139) <= '1';
    layer1_outputs(2140) <= layer0_outputs(255);
    layer1_outputs(2141) <= (layer0_outputs(3951)) and (layer0_outputs(8513));
    layer1_outputs(2142) <= (layer0_outputs(4496)) xor (layer0_outputs(4889));
    layer1_outputs(2143) <= layer0_outputs(2819);
    layer1_outputs(2144) <= not((layer0_outputs(6755)) or (layer0_outputs(6094)));
    layer1_outputs(2145) <= (layer0_outputs(1472)) and (layer0_outputs(5854));
    layer1_outputs(2146) <= (layer0_outputs(2372)) xor (layer0_outputs(524));
    layer1_outputs(2147) <= not(layer0_outputs(543));
    layer1_outputs(2148) <= not(layer0_outputs(3534)) or (layer0_outputs(6499));
    layer1_outputs(2149) <= not((layer0_outputs(1048)) or (layer0_outputs(5688)));
    layer1_outputs(2150) <= layer0_outputs(8358);
    layer1_outputs(2151) <= not(layer0_outputs(7959));
    layer1_outputs(2152) <= (layer0_outputs(8894)) or (layer0_outputs(2981));
    layer1_outputs(2153) <= (layer0_outputs(767)) and not (layer0_outputs(1725));
    layer1_outputs(2154) <= '0';
    layer1_outputs(2155) <= (layer0_outputs(554)) and not (layer0_outputs(542));
    layer1_outputs(2156) <= layer0_outputs(6988);
    layer1_outputs(2157) <= (layer0_outputs(4576)) and not (layer0_outputs(6611));
    layer1_outputs(2158) <= not((layer0_outputs(7766)) and (layer0_outputs(1413)));
    layer1_outputs(2159) <= not(layer0_outputs(2636));
    layer1_outputs(2160) <= not((layer0_outputs(9868)) xor (layer0_outputs(10126)));
    layer1_outputs(2161) <= layer0_outputs(5842);
    layer1_outputs(2162) <= (layer0_outputs(607)) and not (layer0_outputs(3323));
    layer1_outputs(2163) <= not(layer0_outputs(7170));
    layer1_outputs(2164) <= (layer0_outputs(9957)) and not (layer0_outputs(5809));
    layer1_outputs(2165) <= not(layer0_outputs(3055)) or (layer0_outputs(5929));
    layer1_outputs(2166) <= (layer0_outputs(2822)) or (layer0_outputs(2627));
    layer1_outputs(2167) <= layer0_outputs(8855);
    layer1_outputs(2168) <= not(layer0_outputs(4143)) or (layer0_outputs(2240));
    layer1_outputs(2169) <= (layer0_outputs(2697)) and (layer0_outputs(124));
    layer1_outputs(2170) <= (layer0_outputs(2596)) and not (layer0_outputs(3669));
    layer1_outputs(2171) <= not((layer0_outputs(1654)) or (layer0_outputs(3683)));
    layer1_outputs(2172) <= (layer0_outputs(7916)) or (layer0_outputs(3470));
    layer1_outputs(2173) <= not(layer0_outputs(4659)) or (layer0_outputs(5913));
    layer1_outputs(2174) <= (layer0_outputs(5394)) and not (layer0_outputs(8337));
    layer1_outputs(2175) <= '1';
    layer1_outputs(2176) <= (layer0_outputs(8252)) and not (layer0_outputs(974));
    layer1_outputs(2177) <= layer0_outputs(7993);
    layer1_outputs(2178) <= layer0_outputs(766);
    layer1_outputs(2179) <= '0';
    layer1_outputs(2180) <= layer0_outputs(8017);
    layer1_outputs(2181) <= (layer0_outputs(8921)) and not (layer0_outputs(5439));
    layer1_outputs(2182) <= (layer0_outputs(1179)) and (layer0_outputs(812));
    layer1_outputs(2183) <= '1';
    layer1_outputs(2184) <= (layer0_outputs(5993)) and (layer0_outputs(2549));
    layer1_outputs(2185) <= (layer0_outputs(389)) and not (layer0_outputs(1174));
    layer1_outputs(2186) <= (layer0_outputs(4317)) or (layer0_outputs(5211));
    layer1_outputs(2187) <= not(layer0_outputs(3567));
    layer1_outputs(2188) <= not((layer0_outputs(2399)) and (layer0_outputs(4268)));
    layer1_outputs(2189) <= not(layer0_outputs(1325));
    layer1_outputs(2190) <= (layer0_outputs(1968)) and (layer0_outputs(6903));
    layer1_outputs(2191) <= not((layer0_outputs(4041)) or (layer0_outputs(3900)));
    layer1_outputs(2192) <= (layer0_outputs(3585)) and (layer0_outputs(9383));
    layer1_outputs(2193) <= (layer0_outputs(1738)) and not (layer0_outputs(9376));
    layer1_outputs(2194) <= '1';
    layer1_outputs(2195) <= '1';
    layer1_outputs(2196) <= not(layer0_outputs(3330));
    layer1_outputs(2197) <= not(layer0_outputs(1324));
    layer1_outputs(2198) <= layer0_outputs(3417);
    layer1_outputs(2199) <= not(layer0_outputs(5845));
    layer1_outputs(2200) <= (layer0_outputs(4352)) and not (layer0_outputs(3828));
    layer1_outputs(2201) <= not(layer0_outputs(9703)) or (layer0_outputs(3879));
    layer1_outputs(2202) <= layer0_outputs(1118);
    layer1_outputs(2203) <= not(layer0_outputs(3953)) or (layer0_outputs(615));
    layer1_outputs(2204) <= not(layer0_outputs(8518)) or (layer0_outputs(5347));
    layer1_outputs(2205) <= not(layer0_outputs(3375));
    layer1_outputs(2206) <= layer0_outputs(5815);
    layer1_outputs(2207) <= not((layer0_outputs(6562)) or (layer0_outputs(3335)));
    layer1_outputs(2208) <= layer0_outputs(7796);
    layer1_outputs(2209) <= (layer0_outputs(6163)) and (layer0_outputs(2994));
    layer1_outputs(2210) <= (layer0_outputs(7754)) and (layer0_outputs(37));
    layer1_outputs(2211) <= not((layer0_outputs(6365)) and (layer0_outputs(2280)));
    layer1_outputs(2212) <= not(layer0_outputs(5754));
    layer1_outputs(2213) <= '0';
    layer1_outputs(2214) <= not(layer0_outputs(8465));
    layer1_outputs(2215) <= not(layer0_outputs(6194)) or (layer0_outputs(2266));
    layer1_outputs(2216) <= not(layer0_outputs(4949)) or (layer0_outputs(3600));
    layer1_outputs(2217) <= not(layer0_outputs(6614)) or (layer0_outputs(9293));
    layer1_outputs(2218) <= '1';
    layer1_outputs(2219) <= (layer0_outputs(1203)) and (layer0_outputs(8360));
    layer1_outputs(2220) <= '0';
    layer1_outputs(2221) <= '0';
    layer1_outputs(2222) <= (layer0_outputs(4692)) or (layer0_outputs(963));
    layer1_outputs(2223) <= '1';
    layer1_outputs(2224) <= (layer0_outputs(2391)) xor (layer0_outputs(269));
    layer1_outputs(2225) <= not(layer0_outputs(9539)) or (layer0_outputs(3312));
    layer1_outputs(2226) <= not(layer0_outputs(3087)) or (layer0_outputs(7509));
    layer1_outputs(2227) <= not((layer0_outputs(6611)) or (layer0_outputs(3727)));
    layer1_outputs(2228) <= not(layer0_outputs(2241));
    layer1_outputs(2229) <= '0';
    layer1_outputs(2230) <= not(layer0_outputs(8738));
    layer1_outputs(2231) <= (layer0_outputs(10146)) and not (layer0_outputs(3818));
    layer1_outputs(2232) <= (layer0_outputs(7629)) or (layer0_outputs(4608));
    layer1_outputs(2233) <= not(layer0_outputs(984));
    layer1_outputs(2234) <= not((layer0_outputs(2246)) and (layer0_outputs(8448)));
    layer1_outputs(2235) <= '0';
    layer1_outputs(2236) <= not((layer0_outputs(3104)) and (layer0_outputs(8967)));
    layer1_outputs(2237) <= not(layer0_outputs(2333));
    layer1_outputs(2238) <= not((layer0_outputs(8706)) and (layer0_outputs(2294)));
    layer1_outputs(2239) <= not(layer0_outputs(9758)) or (layer0_outputs(479));
    layer1_outputs(2240) <= not(layer0_outputs(7670));
    layer1_outputs(2241) <= '1';
    layer1_outputs(2242) <= not(layer0_outputs(7391));
    layer1_outputs(2243) <= (layer0_outputs(4274)) and not (layer0_outputs(2364));
    layer1_outputs(2244) <= not(layer0_outputs(1773));
    layer1_outputs(2245) <= layer0_outputs(2441);
    layer1_outputs(2246) <= (layer0_outputs(8711)) and not (layer0_outputs(3856));
    layer1_outputs(2247) <= (layer0_outputs(6915)) xor (layer0_outputs(4276));
    layer1_outputs(2248) <= not(layer0_outputs(6313));
    layer1_outputs(2249) <= not(layer0_outputs(3918)) or (layer0_outputs(940));
    layer1_outputs(2250) <= (layer0_outputs(3309)) and not (layer0_outputs(274));
    layer1_outputs(2251) <= not((layer0_outputs(4510)) and (layer0_outputs(1358)));
    layer1_outputs(2252) <= not(layer0_outputs(9986));
    layer1_outputs(2253) <= not(layer0_outputs(3664));
    layer1_outputs(2254) <= (layer0_outputs(1838)) or (layer0_outputs(6853));
    layer1_outputs(2255) <= not((layer0_outputs(7952)) and (layer0_outputs(6301)));
    layer1_outputs(2256) <= (layer0_outputs(5612)) and not (layer0_outputs(6399));
    layer1_outputs(2257) <= not((layer0_outputs(2317)) xor (layer0_outputs(2089)));
    layer1_outputs(2258) <= not((layer0_outputs(591)) and (layer0_outputs(7857)));
    layer1_outputs(2259) <= not(layer0_outputs(9980));
    layer1_outputs(2260) <= (layer0_outputs(60)) and not (layer0_outputs(9958));
    layer1_outputs(2261) <= not(layer0_outputs(5468));
    layer1_outputs(2262) <= not(layer0_outputs(2203)) or (layer0_outputs(3629));
    layer1_outputs(2263) <= not((layer0_outputs(9443)) and (layer0_outputs(1745)));
    layer1_outputs(2264) <= not((layer0_outputs(834)) and (layer0_outputs(4201)));
    layer1_outputs(2265) <= layer0_outputs(2523);
    layer1_outputs(2266) <= (layer0_outputs(686)) and not (layer0_outputs(3533));
    layer1_outputs(2267) <= layer0_outputs(409);
    layer1_outputs(2268) <= layer0_outputs(5048);
    layer1_outputs(2269) <= (layer0_outputs(9266)) or (layer0_outputs(4997));
    layer1_outputs(2270) <= '1';
    layer1_outputs(2271) <= not(layer0_outputs(1357));
    layer1_outputs(2272) <= not((layer0_outputs(8228)) and (layer0_outputs(6504)));
    layer1_outputs(2273) <= not(layer0_outputs(2610)) or (layer0_outputs(8050));
    layer1_outputs(2274) <= (layer0_outputs(3780)) and not (layer0_outputs(9288));
    layer1_outputs(2275) <= not(layer0_outputs(6857)) or (layer0_outputs(5927));
    layer1_outputs(2276) <= not(layer0_outputs(4477)) or (layer0_outputs(6622));
    layer1_outputs(2277) <= layer0_outputs(6208);
    layer1_outputs(2278) <= (layer0_outputs(1775)) and not (layer0_outputs(2057));
    layer1_outputs(2279) <= (layer0_outputs(7403)) and (layer0_outputs(8200));
    layer1_outputs(2280) <= not(layer0_outputs(975));
    layer1_outputs(2281) <= '0';
    layer1_outputs(2282) <= (layer0_outputs(4775)) xor (layer0_outputs(7861));
    layer1_outputs(2283) <= not(layer0_outputs(6323)) or (layer0_outputs(3474));
    layer1_outputs(2284) <= not(layer0_outputs(2175)) or (layer0_outputs(5841));
    layer1_outputs(2285) <= layer0_outputs(6002);
    layer1_outputs(2286) <= not((layer0_outputs(4505)) and (layer0_outputs(5756)));
    layer1_outputs(2287) <= (layer0_outputs(5816)) and not (layer0_outputs(5717));
    layer1_outputs(2288) <= not(layer0_outputs(2452));
    layer1_outputs(2289) <= not((layer0_outputs(6539)) and (layer0_outputs(1081)));
    layer1_outputs(2290) <= layer0_outputs(1651);
    layer1_outputs(2291) <= not((layer0_outputs(5549)) or (layer0_outputs(5633)));
    layer1_outputs(2292) <= not((layer0_outputs(4250)) and (layer0_outputs(6661)));
    layer1_outputs(2293) <= not(layer0_outputs(4777));
    layer1_outputs(2294) <= (layer0_outputs(1591)) and (layer0_outputs(3314));
    layer1_outputs(2295) <= not((layer0_outputs(4740)) or (layer0_outputs(10182)));
    layer1_outputs(2296) <= layer0_outputs(8922);
    layer1_outputs(2297) <= (layer0_outputs(2673)) or (layer0_outputs(4591));
    layer1_outputs(2298) <= not((layer0_outputs(7091)) and (layer0_outputs(1008)));
    layer1_outputs(2299) <= '1';
    layer1_outputs(2300) <= not((layer0_outputs(9537)) and (layer0_outputs(4333)));
    layer1_outputs(2301) <= (layer0_outputs(1992)) and (layer0_outputs(8635));
    layer1_outputs(2302) <= (layer0_outputs(3340)) and not (layer0_outputs(10125));
    layer1_outputs(2303) <= (layer0_outputs(8612)) and (layer0_outputs(872));
    layer1_outputs(2304) <= not((layer0_outputs(1256)) xor (layer0_outputs(7657)));
    layer1_outputs(2305) <= layer0_outputs(2216);
    layer1_outputs(2306) <= (layer0_outputs(1936)) xor (layer0_outputs(8308));
    layer1_outputs(2307) <= (layer0_outputs(4437)) and not (layer0_outputs(2191));
    layer1_outputs(2308) <= not(layer0_outputs(3747));
    layer1_outputs(2309) <= '0';
    layer1_outputs(2310) <= not((layer0_outputs(3488)) xor (layer0_outputs(5085)));
    layer1_outputs(2311) <= not(layer0_outputs(6723));
    layer1_outputs(2312) <= layer0_outputs(6074);
    layer1_outputs(2313) <= (layer0_outputs(3721)) and (layer0_outputs(1816));
    layer1_outputs(2314) <= (layer0_outputs(9230)) or (layer0_outputs(3074));
    layer1_outputs(2315) <= (layer0_outputs(1766)) and not (layer0_outputs(2236));
    layer1_outputs(2316) <= '1';
    layer1_outputs(2317) <= not(layer0_outputs(8319)) or (layer0_outputs(6298));
    layer1_outputs(2318) <= not(layer0_outputs(3175));
    layer1_outputs(2319) <= not((layer0_outputs(4582)) or (layer0_outputs(1310)));
    layer1_outputs(2320) <= not((layer0_outputs(9511)) and (layer0_outputs(5436)));
    layer1_outputs(2321) <= not(layer0_outputs(8713)) or (layer0_outputs(2583));
    layer1_outputs(2322) <= not(layer0_outputs(8459)) or (layer0_outputs(1978));
    layer1_outputs(2323) <= layer0_outputs(9889);
    layer1_outputs(2324) <= not((layer0_outputs(6035)) xor (layer0_outputs(2298)));
    layer1_outputs(2325) <= not((layer0_outputs(2368)) xor (layer0_outputs(1237)));
    layer1_outputs(2326) <= not(layer0_outputs(9922));
    layer1_outputs(2327) <= (layer0_outputs(1522)) and not (layer0_outputs(8580));
    layer1_outputs(2328) <= (layer0_outputs(4097)) and not (layer0_outputs(432));
    layer1_outputs(2329) <= not((layer0_outputs(6583)) and (layer0_outputs(172)));
    layer1_outputs(2330) <= not(layer0_outputs(2951));
    layer1_outputs(2331) <= not(layer0_outputs(3071));
    layer1_outputs(2332) <= not(layer0_outputs(6029));
    layer1_outputs(2333) <= not(layer0_outputs(1791)) or (layer0_outputs(10038));
    layer1_outputs(2334) <= (layer0_outputs(5163)) and (layer0_outputs(2749));
    layer1_outputs(2335) <= (layer0_outputs(7938)) and (layer0_outputs(7830));
    layer1_outputs(2336) <= '1';
    layer1_outputs(2337) <= not(layer0_outputs(9975));
    layer1_outputs(2338) <= layer0_outputs(1349);
    layer1_outputs(2339) <= not(layer0_outputs(6152));
    layer1_outputs(2340) <= '1';
    layer1_outputs(2341) <= layer0_outputs(8807);
    layer1_outputs(2342) <= not(layer0_outputs(9063)) or (layer0_outputs(4665));
    layer1_outputs(2343) <= (layer0_outputs(72)) or (layer0_outputs(7996));
    layer1_outputs(2344) <= not((layer0_outputs(9461)) or (layer0_outputs(5896)));
    layer1_outputs(2345) <= not((layer0_outputs(6022)) and (layer0_outputs(4292)));
    layer1_outputs(2346) <= (layer0_outputs(8420)) and not (layer0_outputs(2338));
    layer1_outputs(2347) <= not(layer0_outputs(2027));
    layer1_outputs(2348) <= layer0_outputs(7998);
    layer1_outputs(2349) <= not(layer0_outputs(3081)) or (layer0_outputs(7301));
    layer1_outputs(2350) <= (layer0_outputs(1946)) and (layer0_outputs(2378));
    layer1_outputs(2351) <= '1';
    layer1_outputs(2352) <= not((layer0_outputs(3073)) xor (layer0_outputs(4509)));
    layer1_outputs(2353) <= layer0_outputs(8124);
    layer1_outputs(2354) <= not((layer0_outputs(10081)) and (layer0_outputs(6824)));
    layer1_outputs(2355) <= '0';
    layer1_outputs(2356) <= '0';
    layer1_outputs(2357) <= (layer0_outputs(4332)) and not (layer0_outputs(3931));
    layer1_outputs(2358) <= '0';
    layer1_outputs(2359) <= layer0_outputs(2127);
    layer1_outputs(2360) <= (layer0_outputs(564)) and not (layer0_outputs(8389));
    layer1_outputs(2361) <= not(layer0_outputs(4812));
    layer1_outputs(2362) <= layer0_outputs(3662);
    layer1_outputs(2363) <= not((layer0_outputs(4000)) and (layer0_outputs(2340)));
    layer1_outputs(2364) <= '0';
    layer1_outputs(2365) <= not(layer0_outputs(9252));
    layer1_outputs(2366) <= not(layer0_outputs(4189));
    layer1_outputs(2367) <= (layer0_outputs(1145)) and (layer0_outputs(7088));
    layer1_outputs(2368) <= not((layer0_outputs(4230)) xor (layer0_outputs(4141)));
    layer1_outputs(2369) <= (layer0_outputs(2410)) and not (layer0_outputs(8603));
    layer1_outputs(2370) <= '0';
    layer1_outputs(2371) <= not((layer0_outputs(4568)) and (layer0_outputs(8644)));
    layer1_outputs(2372) <= not(layer0_outputs(122));
    layer1_outputs(2373) <= (layer0_outputs(3865)) and not (layer0_outputs(2682));
    layer1_outputs(2374) <= (layer0_outputs(5927)) and (layer0_outputs(1805));
    layer1_outputs(2375) <= (layer0_outputs(7482)) and not (layer0_outputs(3720));
    layer1_outputs(2376) <= not(layer0_outputs(5270));
    layer1_outputs(2377) <= layer0_outputs(4451);
    layer1_outputs(2378) <= not(layer0_outputs(6103));
    layer1_outputs(2379) <= layer0_outputs(6326);
    layer1_outputs(2380) <= not(layer0_outputs(2353)) or (layer0_outputs(3523));
    layer1_outputs(2381) <= (layer0_outputs(7784)) xor (layer0_outputs(8000));
    layer1_outputs(2382) <= not((layer0_outputs(449)) and (layer0_outputs(9891)));
    layer1_outputs(2383) <= layer0_outputs(196);
    layer1_outputs(2384) <= not((layer0_outputs(1004)) xor (layer0_outputs(4808)));
    layer1_outputs(2385) <= not((layer0_outputs(8396)) xor (layer0_outputs(9793)));
    layer1_outputs(2386) <= not(layer0_outputs(6851));
    layer1_outputs(2387) <= layer0_outputs(6393);
    layer1_outputs(2388) <= '1';
    layer1_outputs(2389) <= (layer0_outputs(4056)) and not (layer0_outputs(8627));
    layer1_outputs(2390) <= '0';
    layer1_outputs(2391) <= not(layer0_outputs(3563));
    layer1_outputs(2392) <= not(layer0_outputs(8054));
    layer1_outputs(2393) <= layer0_outputs(2616);
    layer1_outputs(2394) <= layer0_outputs(478);
    layer1_outputs(2395) <= not(layer0_outputs(3627));
    layer1_outputs(2396) <= layer0_outputs(7175);
    layer1_outputs(2397) <= (layer0_outputs(10113)) or (layer0_outputs(6246));
    layer1_outputs(2398) <= not(layer0_outputs(8253));
    layer1_outputs(2399) <= (layer0_outputs(1032)) and not (layer0_outputs(7546));
    layer1_outputs(2400) <= not(layer0_outputs(8318));
    layer1_outputs(2401) <= layer0_outputs(8775);
    layer1_outputs(2402) <= layer0_outputs(3309);
    layer1_outputs(2403) <= not(layer0_outputs(9596)) or (layer0_outputs(1734));
    layer1_outputs(2404) <= not(layer0_outputs(3971));
    layer1_outputs(2405) <= layer0_outputs(3836);
    layer1_outputs(2406) <= not((layer0_outputs(6713)) and (layer0_outputs(2193)));
    layer1_outputs(2407) <= '1';
    layer1_outputs(2408) <= layer0_outputs(6068);
    layer1_outputs(2409) <= not(layer0_outputs(636)) or (layer0_outputs(77));
    layer1_outputs(2410) <= layer0_outputs(316);
    layer1_outputs(2411) <= not((layer0_outputs(2969)) and (layer0_outputs(3210)));
    layer1_outputs(2412) <= not((layer0_outputs(4609)) and (layer0_outputs(4457)));
    layer1_outputs(2413) <= (layer0_outputs(9039)) and not (layer0_outputs(4804));
    layer1_outputs(2414) <= layer0_outputs(8161);
    layer1_outputs(2415) <= (layer0_outputs(356)) and not (layer0_outputs(5107));
    layer1_outputs(2416) <= (layer0_outputs(2265)) or (layer0_outputs(834));
    layer1_outputs(2417) <= not((layer0_outputs(4806)) xor (layer0_outputs(6255)));
    layer1_outputs(2418) <= layer0_outputs(4738);
    layer1_outputs(2419) <= (layer0_outputs(3923)) and (layer0_outputs(4112));
    layer1_outputs(2420) <= (layer0_outputs(906)) and not (layer0_outputs(9536));
    layer1_outputs(2421) <= layer0_outputs(4947);
    layer1_outputs(2422) <= layer0_outputs(7980);
    layer1_outputs(2423) <= not(layer0_outputs(5998)) or (layer0_outputs(6696));
    layer1_outputs(2424) <= not((layer0_outputs(8646)) and (layer0_outputs(4858)));
    layer1_outputs(2425) <= layer0_outputs(9990);
    layer1_outputs(2426) <= not(layer0_outputs(5558));
    layer1_outputs(2427) <= not(layer0_outputs(730)) or (layer0_outputs(10129));
    layer1_outputs(2428) <= (layer0_outputs(2886)) xor (layer0_outputs(1075));
    layer1_outputs(2429) <= layer0_outputs(5841);
    layer1_outputs(2430) <= '0';
    layer1_outputs(2431) <= not((layer0_outputs(8722)) xor (layer0_outputs(4917)));
    layer1_outputs(2432) <= layer0_outputs(1007);
    layer1_outputs(2433) <= (layer0_outputs(9400)) and not (layer0_outputs(4722));
    layer1_outputs(2434) <= (layer0_outputs(1933)) and not (layer0_outputs(3196));
    layer1_outputs(2435) <= not((layer0_outputs(1937)) xor (layer0_outputs(3967)));
    layer1_outputs(2436) <= layer0_outputs(3308);
    layer1_outputs(2437) <= '1';
    layer1_outputs(2438) <= not((layer0_outputs(9285)) or (layer0_outputs(9885)));
    layer1_outputs(2439) <= not(layer0_outputs(4424));
    layer1_outputs(2440) <= not((layer0_outputs(7914)) or (layer0_outputs(5474)));
    layer1_outputs(2441) <= not((layer0_outputs(1870)) and (layer0_outputs(488)));
    layer1_outputs(2442) <= layer0_outputs(3140);
    layer1_outputs(2443) <= (layer0_outputs(7740)) or (layer0_outputs(9217));
    layer1_outputs(2444) <= (layer0_outputs(1171)) and not (layer0_outputs(4756));
    layer1_outputs(2445) <= (layer0_outputs(9175)) xor (layer0_outputs(8834));
    layer1_outputs(2446) <= (layer0_outputs(2170)) xor (layer0_outputs(5683));
    layer1_outputs(2447) <= not((layer0_outputs(6821)) xor (layer0_outputs(8399)));
    layer1_outputs(2448) <= (layer0_outputs(8190)) and (layer0_outputs(3861));
    layer1_outputs(2449) <= not(layer0_outputs(7692)) or (layer0_outputs(2541));
    layer1_outputs(2450) <= not((layer0_outputs(7193)) or (layer0_outputs(4825)));
    layer1_outputs(2451) <= (layer0_outputs(9010)) xor (layer0_outputs(551));
    layer1_outputs(2452) <= not((layer0_outputs(420)) or (layer0_outputs(7583)));
    layer1_outputs(2453) <= (layer0_outputs(2341)) and not (layer0_outputs(5351));
    layer1_outputs(2454) <= layer0_outputs(106);
    layer1_outputs(2455) <= layer0_outputs(343);
    layer1_outputs(2456) <= layer0_outputs(6236);
    layer1_outputs(2457) <= not(layer0_outputs(9996));
    layer1_outputs(2458) <= not(layer0_outputs(1814));
    layer1_outputs(2459) <= '0';
    layer1_outputs(2460) <= not((layer0_outputs(7877)) or (layer0_outputs(9108)));
    layer1_outputs(2461) <= layer0_outputs(8081);
    layer1_outputs(2462) <= not(layer0_outputs(1551));
    layer1_outputs(2463) <= layer0_outputs(3393);
    layer1_outputs(2464) <= (layer0_outputs(2768)) and not (layer0_outputs(9069));
    layer1_outputs(2465) <= '1';
    layer1_outputs(2466) <= not(layer0_outputs(6790));
    layer1_outputs(2467) <= not((layer0_outputs(1138)) or (layer0_outputs(2097)));
    layer1_outputs(2468) <= layer0_outputs(7379);
    layer1_outputs(2469) <= layer0_outputs(7808);
    layer1_outputs(2470) <= not(layer0_outputs(6900));
    layer1_outputs(2471) <= not(layer0_outputs(212));
    layer1_outputs(2472) <= (layer0_outputs(4574)) and not (layer0_outputs(968));
    layer1_outputs(2473) <= not((layer0_outputs(2167)) and (layer0_outputs(3880)));
    layer1_outputs(2474) <= not(layer0_outputs(6183));
    layer1_outputs(2475) <= not(layer0_outputs(2106));
    layer1_outputs(2476) <= not(layer0_outputs(974)) or (layer0_outputs(5050));
    layer1_outputs(2477) <= layer0_outputs(6605);
    layer1_outputs(2478) <= not(layer0_outputs(3213)) or (layer0_outputs(708));
    layer1_outputs(2479) <= not(layer0_outputs(1152));
    layer1_outputs(2480) <= not(layer0_outputs(6149)) or (layer0_outputs(810));
    layer1_outputs(2481) <= layer0_outputs(10129);
    layer1_outputs(2482) <= '0';
    layer1_outputs(2483) <= not(layer0_outputs(8533)) or (layer0_outputs(170));
    layer1_outputs(2484) <= not(layer0_outputs(9440));
    layer1_outputs(2485) <= (layer0_outputs(6883)) and (layer0_outputs(5462));
    layer1_outputs(2486) <= (layer0_outputs(7136)) and (layer0_outputs(4733));
    layer1_outputs(2487) <= layer0_outputs(904);
    layer1_outputs(2488) <= not(layer0_outputs(1879));
    layer1_outputs(2489) <= (layer0_outputs(2115)) and (layer0_outputs(7910));
    layer1_outputs(2490) <= not(layer0_outputs(291)) or (layer0_outputs(1243));
    layer1_outputs(2491) <= layer0_outputs(3083);
    layer1_outputs(2492) <= layer0_outputs(642);
    layer1_outputs(2493) <= (layer0_outputs(3496)) or (layer0_outputs(3957));
    layer1_outputs(2494) <= '1';
    layer1_outputs(2495) <= '0';
    layer1_outputs(2496) <= (layer0_outputs(239)) or (layer0_outputs(6243));
    layer1_outputs(2497) <= not(layer0_outputs(7115));
    layer1_outputs(2498) <= '0';
    layer1_outputs(2499) <= not((layer0_outputs(3023)) and (layer0_outputs(212)));
    layer1_outputs(2500) <= layer0_outputs(4542);
    layer1_outputs(2501) <= not(layer0_outputs(5390)) or (layer0_outputs(1071));
    layer1_outputs(2502) <= not(layer0_outputs(2332));
    layer1_outputs(2503) <= not((layer0_outputs(6782)) or (layer0_outputs(6761)));
    layer1_outputs(2504) <= not(layer0_outputs(9067));
    layer1_outputs(2505) <= not(layer0_outputs(3010)) or (layer0_outputs(4477));
    layer1_outputs(2506) <= not(layer0_outputs(4586)) or (layer0_outputs(1462));
    layer1_outputs(2507) <= not(layer0_outputs(304)) or (layer0_outputs(8886));
    layer1_outputs(2508) <= layer0_outputs(9512);
    layer1_outputs(2509) <= (layer0_outputs(4946)) xor (layer0_outputs(9379));
    layer1_outputs(2510) <= not(layer0_outputs(8567));
    layer1_outputs(2511) <= (layer0_outputs(45)) and not (layer0_outputs(378));
    layer1_outputs(2512) <= not(layer0_outputs(2402)) or (layer0_outputs(6935));
    layer1_outputs(2513) <= not(layer0_outputs(4384));
    layer1_outputs(2514) <= not((layer0_outputs(8399)) and (layer0_outputs(2866)));
    layer1_outputs(2515) <= not(layer0_outputs(334)) or (layer0_outputs(8435));
    layer1_outputs(2516) <= (layer0_outputs(5731)) or (layer0_outputs(7710));
    layer1_outputs(2517) <= not(layer0_outputs(5196)) or (layer0_outputs(1591));
    layer1_outputs(2518) <= (layer0_outputs(8485)) or (layer0_outputs(5191));
    layer1_outputs(2519) <= layer0_outputs(7352);
    layer1_outputs(2520) <= layer0_outputs(3014);
    layer1_outputs(2521) <= layer0_outputs(8324);
    layer1_outputs(2522) <= not(layer0_outputs(8335));
    layer1_outputs(2523) <= not((layer0_outputs(2300)) and (layer0_outputs(1422)));
    layer1_outputs(2524) <= not(layer0_outputs(7282));
    layer1_outputs(2525) <= '1';
    layer1_outputs(2526) <= layer0_outputs(8305);
    layer1_outputs(2527) <= not(layer0_outputs(6321)) or (layer0_outputs(1556));
    layer1_outputs(2528) <= layer0_outputs(3753);
    layer1_outputs(2529) <= (layer0_outputs(6515)) and (layer0_outputs(6106));
    layer1_outputs(2530) <= not(layer0_outputs(5948));
    layer1_outputs(2531) <= layer0_outputs(3000);
    layer1_outputs(2532) <= '0';
    layer1_outputs(2533) <= layer0_outputs(8337);
    layer1_outputs(2534) <= layer0_outputs(9491);
    layer1_outputs(2535) <= not(layer0_outputs(8108)) or (layer0_outputs(8016));
    layer1_outputs(2536) <= not(layer0_outputs(338));
    layer1_outputs(2537) <= (layer0_outputs(6502)) and not (layer0_outputs(9256));
    layer1_outputs(2538) <= (layer0_outputs(7239)) or (layer0_outputs(5345));
    layer1_outputs(2539) <= '0';
    layer1_outputs(2540) <= layer0_outputs(3293);
    layer1_outputs(2541) <= (layer0_outputs(8043)) and not (layer0_outputs(5342));
    layer1_outputs(2542) <= not((layer0_outputs(5218)) and (layer0_outputs(3374)));
    layer1_outputs(2543) <= not((layer0_outputs(9830)) and (layer0_outputs(3704)));
    layer1_outputs(2544) <= (layer0_outputs(7704)) xor (layer0_outputs(8142));
    layer1_outputs(2545) <= (layer0_outputs(6262)) and not (layer0_outputs(5571));
    layer1_outputs(2546) <= layer0_outputs(6754);
    layer1_outputs(2547) <= not(layer0_outputs(7095)) or (layer0_outputs(1577));
    layer1_outputs(2548) <= (layer0_outputs(2965)) and (layer0_outputs(9301));
    layer1_outputs(2549) <= (layer0_outputs(9623)) and (layer0_outputs(734));
    layer1_outputs(2550) <= not(layer0_outputs(5108));
    layer1_outputs(2551) <= (layer0_outputs(6340)) or (layer0_outputs(6774));
    layer1_outputs(2552) <= not((layer0_outputs(9604)) xor (layer0_outputs(598)));
    layer1_outputs(2553) <= (layer0_outputs(9823)) and (layer0_outputs(1455));
    layer1_outputs(2554) <= (layer0_outputs(3077)) or (layer0_outputs(4291));
    layer1_outputs(2555) <= (layer0_outputs(9631)) and (layer0_outputs(283));
    layer1_outputs(2556) <= not(layer0_outputs(1265));
    layer1_outputs(2557) <= not((layer0_outputs(5897)) or (layer0_outputs(3139)));
    layer1_outputs(2558) <= not(layer0_outputs(9618)) or (layer0_outputs(3911));
    layer1_outputs(2559) <= (layer0_outputs(6802)) and not (layer0_outputs(1446));
    layer1_outputs(2560) <= layer0_outputs(5545);
    layer1_outputs(2561) <= not((layer0_outputs(4233)) and (layer0_outputs(3042)));
    layer1_outputs(2562) <= not(layer0_outputs(9772));
    layer1_outputs(2563) <= not(layer0_outputs(6209)) or (layer0_outputs(8971));
    layer1_outputs(2564) <= not(layer0_outputs(9257));
    layer1_outputs(2565) <= not((layer0_outputs(163)) and (layer0_outputs(4615)));
    layer1_outputs(2566) <= layer0_outputs(7090);
    layer1_outputs(2567) <= (layer0_outputs(2403)) and not (layer0_outputs(89));
    layer1_outputs(2568) <= '0';
    layer1_outputs(2569) <= '1';
    layer1_outputs(2570) <= not((layer0_outputs(9277)) and (layer0_outputs(7574)));
    layer1_outputs(2571) <= not(layer0_outputs(613));
    layer1_outputs(2572) <= not(layer0_outputs(2325));
    layer1_outputs(2573) <= not(layer0_outputs(6716));
    layer1_outputs(2574) <= (layer0_outputs(1102)) xor (layer0_outputs(6369));
    layer1_outputs(2575) <= layer0_outputs(5016);
    layer1_outputs(2576) <= (layer0_outputs(6691)) or (layer0_outputs(148));
    layer1_outputs(2577) <= not(layer0_outputs(363));
    layer1_outputs(2578) <= (layer0_outputs(4635)) and (layer0_outputs(2906));
    layer1_outputs(2579) <= not(layer0_outputs(3277));
    layer1_outputs(2580) <= not(layer0_outputs(624)) or (layer0_outputs(3520));
    layer1_outputs(2581) <= (layer0_outputs(4338)) xor (layer0_outputs(6388));
    layer1_outputs(2582) <= not(layer0_outputs(9563));
    layer1_outputs(2583) <= not((layer0_outputs(602)) xor (layer0_outputs(186)));
    layer1_outputs(2584) <= (layer0_outputs(2897)) xor (layer0_outputs(8555));
    layer1_outputs(2585) <= not(layer0_outputs(1280));
    layer1_outputs(2586) <= not((layer0_outputs(9567)) and (layer0_outputs(5412)));
    layer1_outputs(2587) <= not(layer0_outputs(1451));
    layer1_outputs(2588) <= not((layer0_outputs(6831)) xor (layer0_outputs(3734)));
    layer1_outputs(2589) <= (layer0_outputs(2714)) and (layer0_outputs(7550));
    layer1_outputs(2590) <= layer0_outputs(949);
    layer1_outputs(2591) <= not((layer0_outputs(3940)) or (layer0_outputs(137)));
    layer1_outputs(2592) <= (layer0_outputs(1614)) or (layer0_outputs(8809));
    layer1_outputs(2593) <= layer0_outputs(2148);
    layer1_outputs(2594) <= layer0_outputs(1161);
    layer1_outputs(2595) <= layer0_outputs(1437);
    layer1_outputs(2596) <= not((layer0_outputs(6333)) and (layer0_outputs(7500)));
    layer1_outputs(2597) <= not(layer0_outputs(7486)) or (layer0_outputs(5284));
    layer1_outputs(2598) <= not(layer0_outputs(9446));
    layer1_outputs(2599) <= layer0_outputs(4060);
    layer1_outputs(2600) <= not((layer0_outputs(4494)) xor (layer0_outputs(5394)));
    layer1_outputs(2601) <= not(layer0_outputs(8756)) or (layer0_outputs(9862));
    layer1_outputs(2602) <= not((layer0_outputs(9583)) or (layer0_outputs(9014)));
    layer1_outputs(2603) <= not(layer0_outputs(836));
    layer1_outputs(2604) <= layer0_outputs(4408);
    layer1_outputs(2605) <= (layer0_outputs(5443)) and (layer0_outputs(1410));
    layer1_outputs(2606) <= not(layer0_outputs(4683)) or (layer0_outputs(2582));
    layer1_outputs(2607) <= (layer0_outputs(1877)) and not (layer0_outputs(2837));
    layer1_outputs(2608) <= (layer0_outputs(7295)) and (layer0_outputs(10149));
    layer1_outputs(2609) <= (layer0_outputs(5835)) or (layer0_outputs(1329));
    layer1_outputs(2610) <= not(layer0_outputs(769));
    layer1_outputs(2611) <= not(layer0_outputs(512));
    layer1_outputs(2612) <= not(layer0_outputs(4402)) or (layer0_outputs(2037));
    layer1_outputs(2613) <= (layer0_outputs(8836)) xor (layer0_outputs(6114));
    layer1_outputs(2614) <= '1';
    layer1_outputs(2615) <= not(layer0_outputs(2823));
    layer1_outputs(2616) <= (layer0_outputs(1560)) and not (layer0_outputs(4232));
    layer1_outputs(2617) <= not(layer0_outputs(3146)) or (layer0_outputs(5850));
    layer1_outputs(2618) <= not(layer0_outputs(4697)) or (layer0_outputs(8609));
    layer1_outputs(2619) <= (layer0_outputs(2357)) xor (layer0_outputs(6877));
    layer1_outputs(2620) <= not((layer0_outputs(5342)) xor (layer0_outputs(1188)));
    layer1_outputs(2621) <= layer0_outputs(177);
    layer1_outputs(2622) <= layer0_outputs(6816);
    layer1_outputs(2623) <= (layer0_outputs(5949)) or (layer0_outputs(1158));
    layer1_outputs(2624) <= layer0_outputs(6844);
    layer1_outputs(2625) <= layer0_outputs(3926);
    layer1_outputs(2626) <= not((layer0_outputs(5738)) and (layer0_outputs(1678)));
    layer1_outputs(2627) <= layer0_outputs(5534);
    layer1_outputs(2628) <= not(layer0_outputs(7851)) or (layer0_outputs(668));
    layer1_outputs(2629) <= (layer0_outputs(9628)) and not (layer0_outputs(9249));
    layer1_outputs(2630) <= (layer0_outputs(6617)) and not (layer0_outputs(3521));
    layer1_outputs(2631) <= layer0_outputs(5450);
    layer1_outputs(2632) <= not(layer0_outputs(2371));
    layer1_outputs(2633) <= '1';
    layer1_outputs(2634) <= (layer0_outputs(397)) and not (layer0_outputs(8264));
    layer1_outputs(2635) <= layer0_outputs(7612);
    layer1_outputs(2636) <= not(layer0_outputs(6943));
    layer1_outputs(2637) <= not(layer0_outputs(4283)) or (layer0_outputs(5476));
    layer1_outputs(2638) <= layer0_outputs(6783);
    layer1_outputs(2639) <= (layer0_outputs(4445)) and (layer0_outputs(6293));
    layer1_outputs(2640) <= layer0_outputs(6809);
    layer1_outputs(2641) <= not((layer0_outputs(3981)) xor (layer0_outputs(7369)));
    layer1_outputs(2642) <= layer0_outputs(9124);
    layer1_outputs(2643) <= not((layer0_outputs(4102)) or (layer0_outputs(5670)));
    layer1_outputs(2644) <= (layer0_outputs(2311)) or (layer0_outputs(9553));
    layer1_outputs(2645) <= (layer0_outputs(1737)) and not (layer0_outputs(2488));
    layer1_outputs(2646) <= (layer0_outputs(8264)) and not (layer0_outputs(9407));
    layer1_outputs(2647) <= not((layer0_outputs(9522)) and (layer0_outputs(3258)));
    layer1_outputs(2648) <= layer0_outputs(818);
    layer1_outputs(2649) <= '0';
    layer1_outputs(2650) <= not(layer0_outputs(9128)) or (layer0_outputs(3774));
    layer1_outputs(2651) <= not(layer0_outputs(4344)) or (layer0_outputs(8493));
    layer1_outputs(2652) <= layer0_outputs(6109);
    layer1_outputs(2653) <= (layer0_outputs(10153)) and (layer0_outputs(7549));
    layer1_outputs(2654) <= layer0_outputs(2246);
    layer1_outputs(2655) <= not(layer0_outputs(9317));
    layer1_outputs(2656) <= (layer0_outputs(4939)) or (layer0_outputs(9147));
    layer1_outputs(2657) <= not((layer0_outputs(6632)) or (layer0_outputs(8261)));
    layer1_outputs(2658) <= (layer0_outputs(3100)) and (layer0_outputs(10047));
    layer1_outputs(2659) <= layer0_outputs(5136);
    layer1_outputs(2660) <= not(layer0_outputs(4646));
    layer1_outputs(2661) <= '1';
    layer1_outputs(2662) <= (layer0_outputs(7321)) and not (layer0_outputs(8293));
    layer1_outputs(2663) <= layer0_outputs(2380);
    layer1_outputs(2664) <= layer0_outputs(4841);
    layer1_outputs(2665) <= '0';
    layer1_outputs(2666) <= not(layer0_outputs(7606));
    layer1_outputs(2667) <= not(layer0_outputs(3983));
    layer1_outputs(2668) <= (layer0_outputs(8499)) and (layer0_outputs(7942));
    layer1_outputs(2669) <= not(layer0_outputs(57));
    layer1_outputs(2670) <= (layer0_outputs(8428)) and (layer0_outputs(10058));
    layer1_outputs(2671) <= (layer0_outputs(610)) and not (layer0_outputs(258));
    layer1_outputs(2672) <= (layer0_outputs(9155)) or (layer0_outputs(30));
    layer1_outputs(2673) <= not(layer0_outputs(7774)) or (layer0_outputs(2448));
    layer1_outputs(2674) <= not(layer0_outputs(8414));
    layer1_outputs(2675) <= not((layer0_outputs(8068)) and (layer0_outputs(7386)));
    layer1_outputs(2676) <= layer0_outputs(3201);
    layer1_outputs(2677) <= not(layer0_outputs(3509));
    layer1_outputs(2678) <= (layer0_outputs(9753)) and (layer0_outputs(9038));
    layer1_outputs(2679) <= not(layer0_outputs(1969));
    layer1_outputs(2680) <= layer0_outputs(9338);
    layer1_outputs(2681) <= not((layer0_outputs(5608)) and (layer0_outputs(7619)));
    layer1_outputs(2682) <= (layer0_outputs(10131)) and not (layer0_outputs(5631));
    layer1_outputs(2683) <= not((layer0_outputs(5883)) and (layer0_outputs(9366)));
    layer1_outputs(2684) <= layer0_outputs(1153);
    layer1_outputs(2685) <= layer0_outputs(2221);
    layer1_outputs(2686) <= not((layer0_outputs(3937)) and (layer0_outputs(2448)));
    layer1_outputs(2687) <= not((layer0_outputs(8825)) or (layer0_outputs(661)));
    layer1_outputs(2688) <= (layer0_outputs(5377)) or (layer0_outputs(4533));
    layer1_outputs(2689) <= layer0_outputs(7568);
    layer1_outputs(2690) <= layer0_outputs(5697);
    layer1_outputs(2691) <= not(layer0_outputs(9857)) or (layer0_outputs(6646));
    layer1_outputs(2692) <= (layer0_outputs(7618)) and not (layer0_outputs(6957));
    layer1_outputs(2693) <= (layer0_outputs(4318)) and not (layer0_outputs(429));
    layer1_outputs(2694) <= (layer0_outputs(948)) or (layer0_outputs(1471));
    layer1_outputs(2695) <= (layer0_outputs(2563)) and not (layer0_outputs(4444));
    layer1_outputs(2696) <= not(layer0_outputs(6958));
    layer1_outputs(2697) <= not(layer0_outputs(3861));
    layer1_outputs(2698) <= (layer0_outputs(8184)) xor (layer0_outputs(985));
    layer1_outputs(2699) <= (layer0_outputs(5405)) and not (layer0_outputs(2096));
    layer1_outputs(2700) <= not(layer0_outputs(9425));
    layer1_outputs(2701) <= (layer0_outputs(7083)) and (layer0_outputs(7149));
    layer1_outputs(2702) <= (layer0_outputs(5093)) or (layer0_outputs(1291));
    layer1_outputs(2703) <= (layer0_outputs(934)) xor (layer0_outputs(10236));
    layer1_outputs(2704) <= (layer0_outputs(5869)) and not (layer0_outputs(4891));
    layer1_outputs(2705) <= not((layer0_outputs(3750)) or (layer0_outputs(6269)));
    layer1_outputs(2706) <= not(layer0_outputs(5964));
    layer1_outputs(2707) <= (layer0_outputs(7453)) and not (layer0_outputs(8544));
    layer1_outputs(2708) <= layer0_outputs(1846);
    layer1_outputs(2709) <= not((layer0_outputs(8653)) and (layer0_outputs(2202)));
    layer1_outputs(2710) <= (layer0_outputs(201)) and not (layer0_outputs(1496));
    layer1_outputs(2711) <= (layer0_outputs(3155)) and (layer0_outputs(5399));
    layer1_outputs(2712) <= not(layer0_outputs(6537)) or (layer0_outputs(4185));
    layer1_outputs(2713) <= '0';
    layer1_outputs(2714) <= not(layer0_outputs(5809)) or (layer0_outputs(8266));
    layer1_outputs(2715) <= not(layer0_outputs(2257));
    layer1_outputs(2716) <= '0';
    layer1_outputs(2717) <= not(layer0_outputs(6501)) or (layer0_outputs(7878));
    layer1_outputs(2718) <= (layer0_outputs(2290)) and not (layer0_outputs(9495));
    layer1_outputs(2719) <= (layer0_outputs(8552)) and (layer0_outputs(7021));
    layer1_outputs(2720) <= not(layer0_outputs(9682));
    layer1_outputs(2721) <= not((layer0_outputs(4571)) or (layer0_outputs(9110)));
    layer1_outputs(2722) <= '1';
    layer1_outputs(2723) <= layer0_outputs(1550);
    layer1_outputs(2724) <= (layer0_outputs(4401)) and (layer0_outputs(707));
    layer1_outputs(2725) <= (layer0_outputs(8268)) and (layer0_outputs(7932));
    layer1_outputs(2726) <= (layer0_outputs(5648)) and not (layer0_outputs(4843));
    layer1_outputs(2727) <= not((layer0_outputs(3944)) and (layer0_outputs(6186)));
    layer1_outputs(2728) <= not(layer0_outputs(5992));
    layer1_outputs(2729) <= '1';
    layer1_outputs(2730) <= '0';
    layer1_outputs(2731) <= (layer0_outputs(4223)) or (layer0_outputs(9420));
    layer1_outputs(2732) <= '0';
    layer1_outputs(2733) <= not(layer0_outputs(4349));
    layer1_outputs(2734) <= (layer0_outputs(3917)) and not (layer0_outputs(1815));
    layer1_outputs(2735) <= not((layer0_outputs(1555)) or (layer0_outputs(3800)));
    layer1_outputs(2736) <= not((layer0_outputs(1286)) xor (layer0_outputs(1426)));
    layer1_outputs(2737) <= (layer0_outputs(1608)) and not (layer0_outputs(1628));
    layer1_outputs(2738) <= (layer0_outputs(6413)) and not (layer0_outputs(7644));
    layer1_outputs(2739) <= not(layer0_outputs(4017));
    layer1_outputs(2740) <= not(layer0_outputs(4614));
    layer1_outputs(2741) <= not(layer0_outputs(4468)) or (layer0_outputs(5556));
    layer1_outputs(2742) <= (layer0_outputs(3153)) and not (layer0_outputs(8560));
    layer1_outputs(2743) <= layer0_outputs(3608);
    layer1_outputs(2744) <= not(layer0_outputs(7735));
    layer1_outputs(2745) <= not(layer0_outputs(3143)) or (layer0_outputs(3229));
    layer1_outputs(2746) <= layer0_outputs(5942);
    layer1_outputs(2747) <= not((layer0_outputs(9418)) and (layer0_outputs(3368)));
    layer1_outputs(2748) <= (layer0_outputs(7016)) and (layer0_outputs(7145));
    layer1_outputs(2749) <= not(layer0_outputs(1600));
    layer1_outputs(2750) <= not((layer0_outputs(7268)) and (layer0_outputs(8480)));
    layer1_outputs(2751) <= not(layer0_outputs(3241)) or (layer0_outputs(5530));
    layer1_outputs(2752) <= (layer0_outputs(10090)) or (layer0_outputs(6296));
    layer1_outputs(2753) <= not(layer0_outputs(8664));
    layer1_outputs(2754) <= layer0_outputs(7423);
    layer1_outputs(2755) <= not(layer0_outputs(5655));
    layer1_outputs(2756) <= not((layer0_outputs(4804)) or (layer0_outputs(3633)));
    layer1_outputs(2757) <= layer0_outputs(9399);
    layer1_outputs(2758) <= not(layer0_outputs(5521)) or (layer0_outputs(182));
    layer1_outputs(2759) <= not(layer0_outputs(7882));
    layer1_outputs(2760) <= (layer0_outputs(4364)) or (layer0_outputs(9108));
    layer1_outputs(2761) <= layer0_outputs(5123);
    layer1_outputs(2762) <= '1';
    layer1_outputs(2763) <= not(layer0_outputs(2079));
    layer1_outputs(2764) <= (layer0_outputs(5542)) and not (layer0_outputs(892));
    layer1_outputs(2765) <= layer0_outputs(876);
    layer1_outputs(2766) <= layer0_outputs(10085);
    layer1_outputs(2767) <= not((layer0_outputs(8424)) and (layer0_outputs(4907)));
    layer1_outputs(2768) <= '1';
    layer1_outputs(2769) <= not((layer0_outputs(7538)) and (layer0_outputs(3848)));
    layer1_outputs(2770) <= layer0_outputs(5107);
    layer1_outputs(2771) <= layer0_outputs(1666);
    layer1_outputs(2772) <= not(layer0_outputs(9477));
    layer1_outputs(2773) <= layer0_outputs(2319);
    layer1_outputs(2774) <= not(layer0_outputs(7751));
    layer1_outputs(2775) <= not(layer0_outputs(6122));
    layer1_outputs(2776) <= (layer0_outputs(4904)) and not (layer0_outputs(9488));
    layer1_outputs(2777) <= '1';
    layer1_outputs(2778) <= (layer0_outputs(8663)) or (layer0_outputs(883));
    layer1_outputs(2779) <= (layer0_outputs(3972)) and (layer0_outputs(2080));
    layer1_outputs(2780) <= (layer0_outputs(6844)) and (layer0_outputs(5015));
    layer1_outputs(2781) <= (layer0_outputs(2554)) and not (layer0_outputs(8768));
    layer1_outputs(2782) <= (layer0_outputs(4522)) or (layer0_outputs(2962));
    layer1_outputs(2783) <= layer0_outputs(10164);
    layer1_outputs(2784) <= (layer0_outputs(7974)) or (layer0_outputs(2594));
    layer1_outputs(2785) <= not((layer0_outputs(1363)) and (layer0_outputs(2756)));
    layer1_outputs(2786) <= layer0_outputs(588);
    layer1_outputs(2787) <= not(layer0_outputs(4311)) or (layer0_outputs(2530));
    layer1_outputs(2788) <= layer0_outputs(9221);
    layer1_outputs(2789) <= not(layer0_outputs(6097)) or (layer0_outputs(9979));
    layer1_outputs(2790) <= (layer0_outputs(4623)) and not (layer0_outputs(5625));
    layer1_outputs(2791) <= not(layer0_outputs(7493)) or (layer0_outputs(5217));
    layer1_outputs(2792) <= not(layer0_outputs(5864));
    layer1_outputs(2793) <= layer0_outputs(8128);
    layer1_outputs(2794) <= not((layer0_outputs(5750)) or (layer0_outputs(169)));
    layer1_outputs(2795) <= not(layer0_outputs(2166));
    layer1_outputs(2796) <= layer0_outputs(9049);
    layer1_outputs(2797) <= (layer0_outputs(9820)) xor (layer0_outputs(4441));
    layer1_outputs(2798) <= not(layer0_outputs(7124)) or (layer0_outputs(59));
    layer1_outputs(2799) <= (layer0_outputs(8542)) and not (layer0_outputs(2865));
    layer1_outputs(2800) <= (layer0_outputs(5431)) xor (layer0_outputs(1389));
    layer1_outputs(2801) <= not(layer0_outputs(2684)) or (layer0_outputs(9137));
    layer1_outputs(2802) <= not(layer0_outputs(5279));
    layer1_outputs(2803) <= '0';
    layer1_outputs(2804) <= not((layer0_outputs(579)) and (layer0_outputs(8432)));
    layer1_outputs(2805) <= layer0_outputs(3973);
    layer1_outputs(2806) <= (layer0_outputs(6749)) and (layer0_outputs(9992));
    layer1_outputs(2807) <= layer0_outputs(1474);
    layer1_outputs(2808) <= (layer0_outputs(8297)) and not (layer0_outputs(2200));
    layer1_outputs(2809) <= (layer0_outputs(86)) and (layer0_outputs(2871));
    layer1_outputs(2810) <= not(layer0_outputs(9156));
    layer1_outputs(2811) <= not(layer0_outputs(4820));
    layer1_outputs(2812) <= (layer0_outputs(3625)) or (layer0_outputs(3016));
    layer1_outputs(2813) <= not(layer0_outputs(9043));
    layer1_outputs(2814) <= not(layer0_outputs(67));
    layer1_outputs(2815) <= not(layer0_outputs(1313));
    layer1_outputs(2816) <= (layer0_outputs(5361)) and not (layer0_outputs(2503));
    layer1_outputs(2817) <= not((layer0_outputs(1174)) or (layer0_outputs(8357)));
    layer1_outputs(2818) <= '1';
    layer1_outputs(2819) <= not(layer0_outputs(7007)) or (layer0_outputs(7976));
    layer1_outputs(2820) <= (layer0_outputs(7191)) and not (layer0_outputs(8411));
    layer1_outputs(2821) <= (layer0_outputs(1521)) and not (layer0_outputs(7780));
    layer1_outputs(2822) <= not(layer0_outputs(9204));
    layer1_outputs(2823) <= not(layer0_outputs(5239));
    layer1_outputs(2824) <= not(layer0_outputs(8270));
    layer1_outputs(2825) <= not(layer0_outputs(7165)) or (layer0_outputs(3614));
    layer1_outputs(2826) <= layer0_outputs(8856);
    layer1_outputs(2827) <= not(layer0_outputs(2923)) or (layer0_outputs(7487));
    layer1_outputs(2828) <= '1';
    layer1_outputs(2829) <= (layer0_outputs(3413)) and not (layer0_outputs(587));
    layer1_outputs(2830) <= not((layer0_outputs(7034)) or (layer0_outputs(3992)));
    layer1_outputs(2831) <= (layer0_outputs(7690)) and (layer0_outputs(4459));
    layer1_outputs(2832) <= not(layer0_outputs(7904)) or (layer0_outputs(9060));
    layer1_outputs(2833) <= layer0_outputs(581);
    layer1_outputs(2834) <= not(layer0_outputs(4856));
    layer1_outputs(2835) <= not(layer0_outputs(7762));
    layer1_outputs(2836) <= not(layer0_outputs(9377)) or (layer0_outputs(1224));
    layer1_outputs(2837) <= not(layer0_outputs(7989));
    layer1_outputs(2838) <= not(layer0_outputs(98));
    layer1_outputs(2839) <= not(layer0_outputs(6169)) or (layer0_outputs(9686));
    layer1_outputs(2840) <= not(layer0_outputs(3523));
    layer1_outputs(2841) <= '1';
    layer1_outputs(2842) <= not(layer0_outputs(5348)) or (layer0_outputs(1742));
    layer1_outputs(2843) <= (layer0_outputs(9167)) or (layer0_outputs(5116));
    layer1_outputs(2844) <= (layer0_outputs(259)) or (layer0_outputs(4329));
    layer1_outputs(2845) <= not(layer0_outputs(7384));
    layer1_outputs(2846) <= (layer0_outputs(3237)) or (layer0_outputs(6963));
    layer1_outputs(2847) <= not((layer0_outputs(5153)) and (layer0_outputs(627)));
    layer1_outputs(2848) <= '0';
    layer1_outputs(2849) <= not(layer0_outputs(8799));
    layer1_outputs(2850) <= layer0_outputs(6229);
    layer1_outputs(2851) <= layer0_outputs(4272);
    layer1_outputs(2852) <= (layer0_outputs(9097)) and (layer0_outputs(7499));
    layer1_outputs(2853) <= layer0_outputs(1185);
    layer1_outputs(2854) <= (layer0_outputs(2134)) or (layer0_outputs(2889));
    layer1_outputs(2855) <= not((layer0_outputs(3443)) and (layer0_outputs(3896)));
    layer1_outputs(2856) <= (layer0_outputs(8457)) and not (layer0_outputs(5623));
    layer1_outputs(2857) <= not(layer0_outputs(8920));
    layer1_outputs(2858) <= not((layer0_outputs(10221)) and (layer0_outputs(2819)));
    layer1_outputs(2859) <= not(layer0_outputs(3320));
    layer1_outputs(2860) <= '1';
    layer1_outputs(2861) <= layer0_outputs(2998);
    layer1_outputs(2862) <= not((layer0_outputs(3183)) and (layer0_outputs(9314)));
    layer1_outputs(2863) <= not((layer0_outputs(1493)) and (layer0_outputs(2902)));
    layer1_outputs(2864) <= (layer0_outputs(5682)) or (layer0_outputs(8595));
    layer1_outputs(2865) <= '0';
    layer1_outputs(2866) <= layer0_outputs(7540);
    layer1_outputs(2867) <= not(layer0_outputs(5337));
    layer1_outputs(2868) <= layer0_outputs(315);
    layer1_outputs(2869) <= '0';
    layer1_outputs(2870) <= not(layer0_outputs(3835)) or (layer0_outputs(4695));
    layer1_outputs(2871) <= (layer0_outputs(4085)) and not (layer0_outputs(984));
    layer1_outputs(2872) <= not(layer0_outputs(5642));
    layer1_outputs(2873) <= (layer0_outputs(6739)) xor (layer0_outputs(797));
    layer1_outputs(2874) <= not(layer0_outputs(7284));
    layer1_outputs(2875) <= layer0_outputs(3896);
    layer1_outputs(2876) <= layer0_outputs(5367);
    layer1_outputs(2877) <= not(layer0_outputs(3539));
    layer1_outputs(2878) <= not((layer0_outputs(3905)) and (layer0_outputs(6027)));
    layer1_outputs(2879) <= (layer0_outputs(9055)) and (layer0_outputs(7803));
    layer1_outputs(2880) <= not(layer0_outputs(10008));
    layer1_outputs(2881) <= not((layer0_outputs(3063)) and (layer0_outputs(4782)));
    layer1_outputs(2882) <= not(layer0_outputs(3770)) or (layer0_outputs(6015));
    layer1_outputs(2883) <= not(layer0_outputs(9149));
    layer1_outputs(2884) <= not(layer0_outputs(644));
    layer1_outputs(2885) <= not(layer0_outputs(5344));
    layer1_outputs(2886) <= not((layer0_outputs(9283)) and (layer0_outputs(9169)));
    layer1_outputs(2887) <= not((layer0_outputs(2100)) and (layer0_outputs(8521)));
    layer1_outputs(2888) <= not(layer0_outputs(9429)) or (layer0_outputs(3925));
    layer1_outputs(2889) <= not(layer0_outputs(3052));
    layer1_outputs(2890) <= not((layer0_outputs(1617)) and (layer0_outputs(6311)));
    layer1_outputs(2891) <= not(layer0_outputs(1116));
    layer1_outputs(2892) <= layer0_outputs(10141);
    layer1_outputs(2893) <= not(layer0_outputs(6633));
    layer1_outputs(2894) <= not((layer0_outputs(2627)) xor (layer0_outputs(5429)));
    layer1_outputs(2895) <= not(layer0_outputs(3162));
    layer1_outputs(2896) <= layer0_outputs(8645);
    layer1_outputs(2897) <= (layer0_outputs(5340)) xor (layer0_outputs(4249));
    layer1_outputs(2898) <= not((layer0_outputs(2606)) or (layer0_outputs(6582)));
    layer1_outputs(2899) <= (layer0_outputs(4540)) and (layer0_outputs(6891));
    layer1_outputs(2900) <= not(layer0_outputs(7506));
    layer1_outputs(2901) <= (layer0_outputs(2881)) xor (layer0_outputs(1817));
    layer1_outputs(2902) <= (layer0_outputs(7347)) and (layer0_outputs(5563));
    layer1_outputs(2903) <= '1';
    layer1_outputs(2904) <= (layer0_outputs(4760)) and (layer0_outputs(4655));
    layer1_outputs(2905) <= (layer0_outputs(778)) xor (layer0_outputs(1265));
    layer1_outputs(2906) <= (layer0_outputs(3873)) xor (layer0_outputs(4047));
    layer1_outputs(2907) <= (layer0_outputs(3209)) and not (layer0_outputs(9449));
    layer1_outputs(2908) <= layer0_outputs(1321);
    layer1_outputs(2909) <= not((layer0_outputs(9919)) or (layer0_outputs(253)));
    layer1_outputs(2910) <= (layer0_outputs(6402)) and not (layer0_outputs(9466));
    layer1_outputs(2911) <= not((layer0_outputs(1771)) and (layer0_outputs(1340)));
    layer1_outputs(2912) <= not(layer0_outputs(8763)) or (layer0_outputs(8463));
    layer1_outputs(2913) <= (layer0_outputs(5778)) and not (layer0_outputs(9858));
    layer1_outputs(2914) <= not(layer0_outputs(3189)) or (layer0_outputs(6782));
    layer1_outputs(2915) <= not(layer0_outputs(5719));
    layer1_outputs(2916) <= (layer0_outputs(1667)) xor (layer0_outputs(4254));
    layer1_outputs(2917) <= (layer0_outputs(627)) or (layer0_outputs(4114));
    layer1_outputs(2918) <= (layer0_outputs(2169)) and (layer0_outputs(3528));
    layer1_outputs(2919) <= (layer0_outputs(10069)) or (layer0_outputs(2321));
    layer1_outputs(2920) <= not((layer0_outputs(9963)) or (layer0_outputs(9764)));
    layer1_outputs(2921) <= '1';
    layer1_outputs(2922) <= (layer0_outputs(6612)) or (layer0_outputs(9066));
    layer1_outputs(2923) <= not(layer0_outputs(1613)) or (layer0_outputs(261));
    layer1_outputs(2924) <= not((layer0_outputs(8862)) or (layer0_outputs(7185)));
    layer1_outputs(2925) <= not((layer0_outputs(5267)) or (layer0_outputs(8038)));
    layer1_outputs(2926) <= layer0_outputs(4488);
    layer1_outputs(2927) <= not(layer0_outputs(4716)) or (layer0_outputs(4989));
    layer1_outputs(2928) <= (layer0_outputs(1899)) and (layer0_outputs(1212));
    layer1_outputs(2929) <= (layer0_outputs(3170)) xor (layer0_outputs(246));
    layer1_outputs(2930) <= layer0_outputs(4322);
    layer1_outputs(2931) <= not((layer0_outputs(7033)) and (layer0_outputs(204)));
    layer1_outputs(2932) <= (layer0_outputs(4709)) and not (layer0_outputs(8938));
    layer1_outputs(2933) <= not(layer0_outputs(4325)) or (layer0_outputs(10053));
    layer1_outputs(2934) <= (layer0_outputs(1360)) or (layer0_outputs(5514));
    layer1_outputs(2935) <= '0';
    layer1_outputs(2936) <= not((layer0_outputs(9481)) xor (layer0_outputs(6421)));
    layer1_outputs(2937) <= (layer0_outputs(2093)) and (layer0_outputs(9725));
    layer1_outputs(2938) <= not(layer0_outputs(4552)) or (layer0_outputs(3217));
    layer1_outputs(2939) <= layer0_outputs(10035);
    layer1_outputs(2940) <= not(layer0_outputs(3150));
    layer1_outputs(2941) <= not((layer0_outputs(1888)) or (layer0_outputs(2726)));
    layer1_outputs(2942) <= (layer0_outputs(7383)) xor (layer0_outputs(8999));
    layer1_outputs(2943) <= (layer0_outputs(7237)) and not (layer0_outputs(3663));
    layer1_outputs(2944) <= not((layer0_outputs(9084)) and (layer0_outputs(8983)));
    layer1_outputs(2945) <= (layer0_outputs(9515)) and not (layer0_outputs(1618));
    layer1_outputs(2946) <= not(layer0_outputs(3573));
    layer1_outputs(2947) <= not(layer0_outputs(2249));
    layer1_outputs(2948) <= not(layer0_outputs(6860));
    layer1_outputs(2949) <= (layer0_outputs(1655)) xor (layer0_outputs(8519));
    layer1_outputs(2950) <= layer0_outputs(3288);
    layer1_outputs(2951) <= '1';
    layer1_outputs(2952) <= (layer0_outputs(453)) and not (layer0_outputs(36));
    layer1_outputs(2953) <= not(layer0_outputs(444));
    layer1_outputs(2954) <= '0';
    layer1_outputs(2955) <= not(layer0_outputs(5949)) or (layer0_outputs(9506));
    layer1_outputs(2956) <= not(layer0_outputs(583)) or (layer0_outputs(6431));
    layer1_outputs(2957) <= not((layer0_outputs(7838)) and (layer0_outputs(7873)));
    layer1_outputs(2958) <= (layer0_outputs(7688)) or (layer0_outputs(2964));
    layer1_outputs(2959) <= not(layer0_outputs(2954));
    layer1_outputs(2960) <= not(layer0_outputs(8813));
    layer1_outputs(2961) <= (layer0_outputs(7)) and (layer0_outputs(1537));
    layer1_outputs(2962) <= (layer0_outputs(7790)) or (layer0_outputs(9731));
    layer1_outputs(2963) <= not(layer0_outputs(270)) or (layer0_outputs(8055));
    layer1_outputs(2964) <= not((layer0_outputs(9305)) or (layer0_outputs(8875)));
    layer1_outputs(2965) <= not(layer0_outputs(2662)) or (layer0_outputs(3265));
    layer1_outputs(2966) <= not(layer0_outputs(687));
    layer1_outputs(2967) <= (layer0_outputs(7621)) and not (layer0_outputs(6124));
    layer1_outputs(2968) <= not((layer0_outputs(6868)) xor (layer0_outputs(5426)));
    layer1_outputs(2969) <= not(layer0_outputs(1407));
    layer1_outputs(2970) <= (layer0_outputs(8246)) and not (layer0_outputs(8737));
    layer1_outputs(2971) <= not((layer0_outputs(10200)) xor (layer0_outputs(5456)));
    layer1_outputs(2972) <= (layer0_outputs(408)) and not (layer0_outputs(8174));
    layer1_outputs(2973) <= not(layer0_outputs(1069));
    layer1_outputs(2974) <= layer0_outputs(7360);
    layer1_outputs(2975) <= '1';
    layer1_outputs(2976) <= not(layer0_outputs(9281)) or (layer0_outputs(96));
    layer1_outputs(2977) <= not((layer0_outputs(8113)) and (layer0_outputs(3334)));
    layer1_outputs(2978) <= layer0_outputs(2268);
    layer1_outputs(2979) <= not(layer0_outputs(3548)) or (layer0_outputs(10195));
    layer1_outputs(2980) <= (layer0_outputs(2684)) and not (layer0_outputs(5111));
    layer1_outputs(2981) <= layer0_outputs(4798);
    layer1_outputs(2982) <= not((layer0_outputs(7349)) or (layer0_outputs(5091)));
    layer1_outputs(2983) <= (layer0_outputs(713)) or (layer0_outputs(8694));
    layer1_outputs(2984) <= (layer0_outputs(5705)) and not (layer0_outputs(3137));
    layer1_outputs(2985) <= not(layer0_outputs(4551));
    layer1_outputs(2986) <= '1';
    layer1_outputs(2987) <= '1';
    layer1_outputs(2988) <= '1';
    layer1_outputs(2989) <= layer0_outputs(4147);
    layer1_outputs(2990) <= (layer0_outputs(5713)) and (layer0_outputs(8339));
    layer1_outputs(2991) <= (layer0_outputs(9437)) and (layer0_outputs(9163));
    layer1_outputs(2992) <= not(layer0_outputs(6575)) or (layer0_outputs(3406));
    layer1_outputs(2993) <= (layer0_outputs(8320)) or (layer0_outputs(6475));
    layer1_outputs(2994) <= layer0_outputs(7794);
    layer1_outputs(2995) <= not(layer0_outputs(2707));
    layer1_outputs(2996) <= not(layer0_outputs(2818));
    layer1_outputs(2997) <= (layer0_outputs(6511)) and not (layer0_outputs(5862));
    layer1_outputs(2998) <= layer0_outputs(9338);
    layer1_outputs(2999) <= (layer0_outputs(6044)) and (layer0_outputs(6469));
    layer1_outputs(3000) <= not(layer0_outputs(2379));
    layer1_outputs(3001) <= (layer0_outputs(3038)) and not (layer0_outputs(6418));
    layer1_outputs(3002) <= '0';
    layer1_outputs(3003) <= not(layer0_outputs(4391)) or (layer0_outputs(6311));
    layer1_outputs(3004) <= (layer0_outputs(9785)) and not (layer0_outputs(3141));
    layer1_outputs(3005) <= '1';
    layer1_outputs(3006) <= (layer0_outputs(5912)) xor (layer0_outputs(7613));
    layer1_outputs(3007) <= not(layer0_outputs(4971)) or (layer0_outputs(8362));
    layer1_outputs(3008) <= not((layer0_outputs(7119)) or (layer0_outputs(9500)));
    layer1_outputs(3009) <= not(layer0_outputs(2641)) or (layer0_outputs(10120));
    layer1_outputs(3010) <= not((layer0_outputs(10169)) or (layer0_outputs(1593)));
    layer1_outputs(3011) <= not((layer0_outputs(6865)) xor (layer0_outputs(8928)));
    layer1_outputs(3012) <= not(layer0_outputs(9873));
    layer1_outputs(3013) <= layer0_outputs(6598);
    layer1_outputs(3014) <= (layer0_outputs(4316)) and (layer0_outputs(8218));
    layer1_outputs(3015) <= (layer0_outputs(3030)) and not (layer0_outputs(6315));
    layer1_outputs(3016) <= (layer0_outputs(557)) and (layer0_outputs(4892));
    layer1_outputs(3017) <= (layer0_outputs(10086)) xor (layer0_outputs(3414));
    layer1_outputs(3018) <= not(layer0_outputs(2060));
    layer1_outputs(3019) <= not(layer0_outputs(7954)) or (layer0_outputs(5066));
    layer1_outputs(3020) <= layer0_outputs(424);
    layer1_outputs(3021) <= not((layer0_outputs(1218)) and (layer0_outputs(7351)));
    layer1_outputs(3022) <= layer0_outputs(8988);
    layer1_outputs(3023) <= not((layer0_outputs(8953)) and (layer0_outputs(1754)));
    layer1_outputs(3024) <= not(layer0_outputs(1210)) or (layer0_outputs(3483));
    layer1_outputs(3025) <= '0';
    layer1_outputs(3026) <= (layer0_outputs(3245)) and (layer0_outputs(2425));
    layer1_outputs(3027) <= layer0_outputs(9855);
    layer1_outputs(3028) <= layer0_outputs(5078);
    layer1_outputs(3029) <= (layer0_outputs(436)) and (layer0_outputs(8353));
    layer1_outputs(3030) <= not((layer0_outputs(6266)) and (layer0_outputs(7269)));
    layer1_outputs(3031) <= layer0_outputs(9557);
    layer1_outputs(3032) <= not(layer0_outputs(3837));
    layer1_outputs(3033) <= not(layer0_outputs(10079)) or (layer0_outputs(3380));
    layer1_outputs(3034) <= '1';
    layer1_outputs(3035) <= not((layer0_outputs(9569)) and (layer0_outputs(8061)));
    layer1_outputs(3036) <= layer0_outputs(8660);
    layer1_outputs(3037) <= not(layer0_outputs(7886)) or (layer0_outputs(5127));
    layer1_outputs(3038) <= (layer0_outputs(1373)) or (layer0_outputs(3651));
    layer1_outputs(3039) <= not((layer0_outputs(5767)) and (layer0_outputs(6485)));
    layer1_outputs(3040) <= not((layer0_outputs(936)) and (layer0_outputs(8137)));
    layer1_outputs(3041) <= '0';
    layer1_outputs(3042) <= not((layer0_outputs(6284)) or (layer0_outputs(9194)));
    layer1_outputs(3043) <= not(layer0_outputs(7832));
    layer1_outputs(3044) <= '1';
    layer1_outputs(3045) <= (layer0_outputs(1926)) and (layer0_outputs(2082));
    layer1_outputs(3046) <= not((layer0_outputs(4564)) or (layer0_outputs(5296)));
    layer1_outputs(3047) <= not(layer0_outputs(9991));
    layer1_outputs(3048) <= layer0_outputs(3572);
    layer1_outputs(3049) <= not(layer0_outputs(9287)) or (layer0_outputs(6937));
    layer1_outputs(3050) <= (layer0_outputs(2055)) xor (layer0_outputs(2734));
    layer1_outputs(3051) <= not(layer0_outputs(6868));
    layer1_outputs(3052) <= not(layer0_outputs(2855));
    layer1_outputs(3053) <= layer0_outputs(5584);
    layer1_outputs(3054) <= not((layer0_outputs(8819)) and (layer0_outputs(8288)));
    layer1_outputs(3055) <= not(layer0_outputs(2377));
    layer1_outputs(3056) <= (layer0_outputs(3111)) and not (layer0_outputs(5931));
    layer1_outputs(3057) <= not((layer0_outputs(1259)) xor (layer0_outputs(3616)));
    layer1_outputs(3058) <= (layer0_outputs(1687)) xor (layer0_outputs(5994));
    layer1_outputs(3059) <= not(layer0_outputs(8194));
    layer1_outputs(3060) <= (layer0_outputs(5866)) and not (layer0_outputs(2731));
    layer1_outputs(3061) <= layer0_outputs(8962);
    layer1_outputs(3062) <= not((layer0_outputs(5960)) or (layer0_outputs(6458)));
    layer1_outputs(3063) <= not((layer0_outputs(9735)) and (layer0_outputs(5518)));
    layer1_outputs(3064) <= (layer0_outputs(1368)) and not (layer0_outputs(7224));
    layer1_outputs(3065) <= '0';
    layer1_outputs(3066) <= (layer0_outputs(5918)) and not (layer0_outputs(7085));
    layer1_outputs(3067) <= layer0_outputs(5293);
    layer1_outputs(3068) <= not((layer0_outputs(1202)) and (layer0_outputs(9218)));
    layer1_outputs(3069) <= '1';
    layer1_outputs(3070) <= not((layer0_outputs(1850)) and (layer0_outputs(2914)));
    layer1_outputs(3071) <= (layer0_outputs(942)) and not (layer0_outputs(4104));
    layer1_outputs(3072) <= not(layer0_outputs(9742));
    layer1_outputs(3073) <= '1';
    layer1_outputs(3074) <= not((layer0_outputs(931)) and (layer0_outputs(5071)));
    layer1_outputs(3075) <= not(layer0_outputs(8150));
    layer1_outputs(3076) <= (layer0_outputs(2335)) and not (layer0_outputs(3869));
    layer1_outputs(3077) <= (layer0_outputs(1610)) and not (layer0_outputs(5097));
    layer1_outputs(3078) <= '0';
    layer1_outputs(3079) <= (layer0_outputs(1383)) xor (layer0_outputs(6717));
    layer1_outputs(3080) <= not(layer0_outputs(1980));
    layer1_outputs(3081) <= not(layer0_outputs(6222)) or (layer0_outputs(5343));
    layer1_outputs(3082) <= '0';
    layer1_outputs(3083) <= (layer0_outputs(7717)) and (layer0_outputs(4959));
    layer1_outputs(3084) <= layer0_outputs(2490);
    layer1_outputs(3085) <= '1';
    layer1_outputs(3086) <= (layer0_outputs(249)) and not (layer0_outputs(6549));
    layer1_outputs(3087) <= '1';
    layer1_outputs(3088) <= layer0_outputs(6503);
    layer1_outputs(3089) <= not(layer0_outputs(9054)) or (layer0_outputs(3065));
    layer1_outputs(3090) <= '0';
    layer1_outputs(3091) <= not((layer0_outputs(9612)) and (layer0_outputs(2612)));
    layer1_outputs(3092) <= layer0_outputs(5171);
    layer1_outputs(3093) <= not(layer0_outputs(7257)) or (layer0_outputs(3440));
    layer1_outputs(3094) <= not((layer0_outputs(3387)) and (layer0_outputs(112)));
    layer1_outputs(3095) <= (layer0_outputs(5205)) and not (layer0_outputs(7307));
    layer1_outputs(3096) <= layer0_outputs(8193);
    layer1_outputs(3097) <= '1';
    layer1_outputs(3098) <= (layer0_outputs(1423)) xor (layer0_outputs(3835));
    layer1_outputs(3099) <= (layer0_outputs(6096)) and not (layer0_outputs(5691));
    layer1_outputs(3100) <= (layer0_outputs(849)) and not (layer0_outputs(6316));
    layer1_outputs(3101) <= not(layer0_outputs(4911));
    layer1_outputs(3102) <= not(layer0_outputs(6991)) or (layer0_outputs(6982));
    layer1_outputs(3103) <= layer0_outputs(147);
    layer1_outputs(3104) <= (layer0_outputs(4811)) and (layer0_outputs(2799));
    layer1_outputs(3105) <= layer0_outputs(10140);
    layer1_outputs(3106) <= layer0_outputs(726);
    layer1_outputs(3107) <= layer0_outputs(7953);
    layer1_outputs(3108) <= not(layer0_outputs(96));
    layer1_outputs(3109) <= not(layer0_outputs(647));
    layer1_outputs(3110) <= (layer0_outputs(1361)) or (layer0_outputs(3228));
    layer1_outputs(3111) <= '1';
    layer1_outputs(3112) <= not((layer0_outputs(823)) and (layer0_outputs(6428)));
    layer1_outputs(3113) <= not(layer0_outputs(3484));
    layer1_outputs(3114) <= not(layer0_outputs(3026)) or (layer0_outputs(4062));
    layer1_outputs(3115) <= (layer0_outputs(5042)) and not (layer0_outputs(5961));
    layer1_outputs(3116) <= (layer0_outputs(4721)) and (layer0_outputs(5917));
    layer1_outputs(3117) <= '1';
    layer1_outputs(3118) <= layer0_outputs(4135);
    layer1_outputs(3119) <= not(layer0_outputs(8961)) or (layer0_outputs(5840));
    layer1_outputs(3120) <= not((layer0_outputs(8896)) and (layer0_outputs(3739)));
    layer1_outputs(3121) <= not((layer0_outputs(2390)) xor (layer0_outputs(9172)));
    layer1_outputs(3122) <= layer0_outputs(6856);
    layer1_outputs(3123) <= not(layer0_outputs(3888));
    layer1_outputs(3124) <= layer0_outputs(3024);
    layer1_outputs(3125) <= not(layer0_outputs(3916));
    layer1_outputs(3126) <= not(layer0_outputs(4465));
    layer1_outputs(3127) <= not((layer0_outputs(4176)) and (layer0_outputs(482)));
    layer1_outputs(3128) <= not((layer0_outputs(1623)) xor (layer0_outputs(4650)));
    layer1_outputs(3129) <= not((layer0_outputs(3420)) and (layer0_outputs(1506)));
    layer1_outputs(3130) <= (layer0_outputs(401)) or (layer0_outputs(3919));
    layer1_outputs(3131) <= '1';
    layer1_outputs(3132) <= '1';
    layer1_outputs(3133) <= layer0_outputs(6173);
    layer1_outputs(3134) <= not((layer0_outputs(4907)) xor (layer0_outputs(252)));
    layer1_outputs(3135) <= not(layer0_outputs(9799));
    layer1_outputs(3136) <= layer0_outputs(8002);
    layer1_outputs(3137) <= (layer0_outputs(888)) xor (layer0_outputs(6362));
    layer1_outputs(3138) <= (layer0_outputs(2437)) or (layer0_outputs(2916));
    layer1_outputs(3139) <= not((layer0_outputs(8078)) or (layer0_outputs(2570)));
    layer1_outputs(3140) <= '0';
    layer1_outputs(3141) <= not(layer0_outputs(3588));
    layer1_outputs(3142) <= (layer0_outputs(5033)) and not (layer0_outputs(4184));
    layer1_outputs(3143) <= not((layer0_outputs(10069)) xor (layer0_outputs(9250)));
    layer1_outputs(3144) <= (layer0_outputs(7456)) and not (layer0_outputs(7193));
    layer1_outputs(3145) <= not(layer0_outputs(7204));
    layer1_outputs(3146) <= layer0_outputs(5008);
    layer1_outputs(3147) <= not(layer0_outputs(1049)) or (layer0_outputs(9909));
    layer1_outputs(3148) <= not(layer0_outputs(4518));
    layer1_outputs(3149) <= not(layer0_outputs(1749)) or (layer0_outputs(4256));
    layer1_outputs(3150) <= layer0_outputs(4923);
    layer1_outputs(3151) <= (layer0_outputs(5894)) and not (layer0_outputs(9406));
    layer1_outputs(3152) <= not(layer0_outputs(1048));
    layer1_outputs(3153) <= (layer0_outputs(2954)) and not (layer0_outputs(4915));
    layer1_outputs(3154) <= '0';
    layer1_outputs(3155) <= not((layer0_outputs(5753)) and (layer0_outputs(7630)));
    layer1_outputs(3156) <= not(layer0_outputs(275));
    layer1_outputs(3157) <= layer0_outputs(3623);
    layer1_outputs(3158) <= '1';
    layer1_outputs(3159) <= layer0_outputs(3993);
    layer1_outputs(3160) <= (layer0_outputs(4846)) and not (layer0_outputs(9283));
    layer1_outputs(3161) <= not((layer0_outputs(8987)) or (layer0_outputs(7061)));
    layer1_outputs(3162) <= (layer0_outputs(5463)) and (layer0_outputs(9828));
    layer1_outputs(3163) <= not(layer0_outputs(9041)) or (layer0_outputs(3095));
    layer1_outputs(3164) <= (layer0_outputs(7350)) and (layer0_outputs(3988));
    layer1_outputs(3165) <= '0';
    layer1_outputs(3166) <= '0';
    layer1_outputs(3167) <= not(layer0_outputs(1599));
    layer1_outputs(3168) <= (layer0_outputs(6531)) and not (layer0_outputs(775));
    layer1_outputs(3169) <= not((layer0_outputs(7520)) xor (layer0_outputs(6573)));
    layer1_outputs(3170) <= layer0_outputs(1313);
    layer1_outputs(3171) <= layer0_outputs(2552);
    layer1_outputs(3172) <= not(layer0_outputs(3201));
    layer1_outputs(3173) <= not(layer0_outputs(2446));
    layer1_outputs(3174) <= not((layer0_outputs(4919)) and (layer0_outputs(3197)));
    layer1_outputs(3175) <= layer0_outputs(800);
    layer1_outputs(3176) <= (layer0_outputs(4619)) and not (layer0_outputs(134));
    layer1_outputs(3177) <= not(layer0_outputs(6036));
    layer1_outputs(3178) <= (layer0_outputs(4271)) and not (layer0_outputs(9819));
    layer1_outputs(3179) <= (layer0_outputs(4593)) and not (layer0_outputs(2776));
    layer1_outputs(3180) <= '0';
    layer1_outputs(3181) <= layer0_outputs(6966);
    layer1_outputs(3182) <= not(layer0_outputs(8692)) or (layer0_outputs(9669));
    layer1_outputs(3183) <= (layer0_outputs(6955)) or (layer0_outputs(7150));
    layer1_outputs(3184) <= not(layer0_outputs(2070)) or (layer0_outputs(6859));
    layer1_outputs(3185) <= layer0_outputs(2630);
    layer1_outputs(3186) <= not(layer0_outputs(2600));
    layer1_outputs(3187) <= (layer0_outputs(4302)) and not (layer0_outputs(7985));
    layer1_outputs(3188) <= (layer0_outputs(10018)) and not (layer0_outputs(4367));
    layer1_outputs(3189) <= not(layer0_outputs(6308));
    layer1_outputs(3190) <= not((layer0_outputs(6777)) and (layer0_outputs(8669)));
    layer1_outputs(3191) <= (layer0_outputs(4329)) xor (layer0_outputs(267));
    layer1_outputs(3192) <= not(layer0_outputs(2814));
    layer1_outputs(3193) <= layer0_outputs(3009);
    layer1_outputs(3194) <= layer0_outputs(9376);
    layer1_outputs(3195) <= '1';
    layer1_outputs(3196) <= not(layer0_outputs(1146)) or (layer0_outputs(4054));
    layer1_outputs(3197) <= (layer0_outputs(231)) and not (layer0_outputs(1585));
    layer1_outputs(3198) <= (layer0_outputs(9916)) and not (layer0_outputs(5786));
    layer1_outputs(3199) <= not(layer0_outputs(2890)) or (layer0_outputs(9307));
    layer1_outputs(3200) <= layer0_outputs(8192);
    layer1_outputs(3201) <= (layer0_outputs(9736)) and not (layer0_outputs(5435));
    layer1_outputs(3202) <= not(layer0_outputs(4251));
    layer1_outputs(3203) <= layer0_outputs(1587);
    layer1_outputs(3204) <= not(layer0_outputs(862)) or (layer0_outputs(10017));
    layer1_outputs(3205) <= (layer0_outputs(1486)) and (layer0_outputs(3547));
    layer1_outputs(3206) <= (layer0_outputs(4810)) and (layer0_outputs(9246));
    layer1_outputs(3207) <= not((layer0_outputs(68)) and (layer0_outputs(2861)));
    layer1_outputs(3208) <= not(layer0_outputs(3039)) or (layer0_outputs(8949));
    layer1_outputs(3209) <= (layer0_outputs(1097)) xor (layer0_outputs(1643));
    layer1_outputs(3210) <= not(layer0_outputs(9379)) or (layer0_outputs(675));
    layer1_outputs(3211) <= (layer0_outputs(6381)) and not (layer0_outputs(2412));
    layer1_outputs(3212) <= not((layer0_outputs(670)) or (layer0_outputs(3771)));
    layer1_outputs(3213) <= not(layer0_outputs(7695)) or (layer0_outputs(7050));
    layer1_outputs(3214) <= not(layer0_outputs(1247));
    layer1_outputs(3215) <= (layer0_outputs(7498)) and not (layer0_outputs(1908));
    layer1_outputs(3216) <= (layer0_outputs(8121)) or (layer0_outputs(1934));
    layer1_outputs(3217) <= not(layer0_outputs(7715));
    layer1_outputs(3218) <= (layer0_outputs(7045)) or (layer0_outputs(6382));
    layer1_outputs(3219) <= (layer0_outputs(7282)) and (layer0_outputs(1811));
    layer1_outputs(3220) <= not(layer0_outputs(5250));
    layer1_outputs(3221) <= layer0_outputs(976);
    layer1_outputs(3222) <= (layer0_outputs(7254)) and (layer0_outputs(8060));
    layer1_outputs(3223) <= not(layer0_outputs(9210));
    layer1_outputs(3224) <= not(layer0_outputs(4648));
    layer1_outputs(3225) <= (layer0_outputs(4548)) and not (layer0_outputs(3253));
    layer1_outputs(3226) <= not(layer0_outputs(3)) or (layer0_outputs(1182));
    layer1_outputs(3227) <= (layer0_outputs(7402)) and (layer0_outputs(3826));
    layer1_outputs(3228) <= not((layer0_outputs(7199)) and (layer0_outputs(7104)));
    layer1_outputs(3229) <= layer0_outputs(1271);
    layer1_outputs(3230) <= (layer0_outputs(1776)) and not (layer0_outputs(1905));
    layer1_outputs(3231) <= (layer0_outputs(5600)) xor (layer0_outputs(3675));
    layer1_outputs(3232) <= not(layer0_outputs(5448)) or (layer0_outputs(4944));
    layer1_outputs(3233) <= layer0_outputs(9193);
    layer1_outputs(3234) <= not((layer0_outputs(1279)) and (layer0_outputs(9792)));
    layer1_outputs(3235) <= (layer0_outputs(8009)) and not (layer0_outputs(6814));
    layer1_outputs(3236) <= not(layer0_outputs(7957));
    layer1_outputs(3237) <= (layer0_outputs(6245)) xor (layer0_outputs(7728));
    layer1_outputs(3238) <= not((layer0_outputs(328)) and (layer0_outputs(5594)));
    layer1_outputs(3239) <= (layer0_outputs(7464)) and not (layer0_outputs(3280));
    layer1_outputs(3240) <= (layer0_outputs(157)) and not (layer0_outputs(537));
    layer1_outputs(3241) <= not((layer0_outputs(785)) xor (layer0_outputs(3777)));
    layer1_outputs(3242) <= not((layer0_outputs(3378)) or (layer0_outputs(8028)));
    layer1_outputs(3243) <= (layer0_outputs(289)) and (layer0_outputs(8535));
    layer1_outputs(3244) <= (layer0_outputs(152)) and not (layer0_outputs(9046));
    layer1_outputs(3245) <= layer0_outputs(3500);
    layer1_outputs(3246) <= not(layer0_outputs(6182));
    layer1_outputs(3247) <= not(layer0_outputs(1103));
    layer1_outputs(3248) <= (layer0_outputs(3968)) or (layer0_outputs(6157));
    layer1_outputs(3249) <= not(layer0_outputs(9080)) or (layer0_outputs(2863));
    layer1_outputs(3250) <= not(layer0_outputs(866)) or (layer0_outputs(9601));
    layer1_outputs(3251) <= not((layer0_outputs(2797)) xor (layer0_outputs(6480)));
    layer1_outputs(3252) <= (layer0_outputs(1698)) or (layer0_outputs(9117));
    layer1_outputs(3253) <= layer0_outputs(6886);
    layer1_outputs(3254) <= layer0_outputs(6112);
    layer1_outputs(3255) <= layer0_outputs(4272);
    layer1_outputs(3256) <= not((layer0_outputs(3131)) or (layer0_outputs(10124)));
    layer1_outputs(3257) <= (layer0_outputs(7012)) and (layer0_outputs(4333));
    layer1_outputs(3258) <= not(layer0_outputs(2546));
    layer1_outputs(3259) <= not(layer0_outputs(334));
    layer1_outputs(3260) <= (layer0_outputs(7189)) and not (layer0_outputs(4083));
    layer1_outputs(3261) <= (layer0_outputs(5244)) xor (layer0_outputs(6210));
    layer1_outputs(3262) <= '0';
    layer1_outputs(3263) <= layer0_outputs(6619);
    layer1_outputs(3264) <= '1';
    layer1_outputs(3265) <= (layer0_outputs(9354)) and (layer0_outputs(1665));
    layer1_outputs(3266) <= '1';
    layer1_outputs(3267) <= not((layer0_outputs(4734)) or (layer0_outputs(1904)));
    layer1_outputs(3268) <= not((layer0_outputs(4531)) and (layer0_outputs(3353)));
    layer1_outputs(3269) <= not((layer0_outputs(3168)) and (layer0_outputs(4988)));
    layer1_outputs(3270) <= (layer0_outputs(1317)) and (layer0_outputs(7899));
    layer1_outputs(3271) <= (layer0_outputs(6937)) and (layer0_outputs(8728));
    layer1_outputs(3272) <= layer0_outputs(2830);
    layer1_outputs(3273) <= not(layer0_outputs(2227));
    layer1_outputs(3274) <= (layer0_outputs(2017)) and (layer0_outputs(2630));
    layer1_outputs(3275) <= '0';
    layer1_outputs(3276) <= not(layer0_outputs(9267));
    layer1_outputs(3277) <= not(layer0_outputs(1457)) or (layer0_outputs(4933));
    layer1_outputs(3278) <= not(layer0_outputs(9048));
    layer1_outputs(3279) <= not(layer0_outputs(7230));
    layer1_outputs(3280) <= '0';
    layer1_outputs(3281) <= '1';
    layer1_outputs(3282) <= not(layer0_outputs(4687)) or (layer0_outputs(6239));
    layer1_outputs(3283) <= not((layer0_outputs(782)) and (layer0_outputs(9851)));
    layer1_outputs(3284) <= (layer0_outputs(1562)) and not (layer0_outputs(1860));
    layer1_outputs(3285) <= not(layer0_outputs(8369)) or (layer0_outputs(8804));
    layer1_outputs(3286) <= not(layer0_outputs(3205));
    layer1_outputs(3287) <= not(layer0_outputs(9022)) or (layer0_outputs(10162));
    layer1_outputs(3288) <= layer0_outputs(2205);
    layer1_outputs(3289) <= layer0_outputs(1732);
    layer1_outputs(3290) <= not(layer0_outputs(3407));
    layer1_outputs(3291) <= layer0_outputs(5442);
    layer1_outputs(3292) <= layer0_outputs(8156);
    layer1_outputs(3293) <= not((layer0_outputs(5453)) and (layer0_outputs(2666)));
    layer1_outputs(3294) <= not(layer0_outputs(649)) or (layer0_outputs(4120));
    layer1_outputs(3295) <= not(layer0_outputs(4046)) or (layer0_outputs(9252));
    layer1_outputs(3296) <= not(layer0_outputs(276)) or (layer0_outputs(1489));
    layer1_outputs(3297) <= '1';
    layer1_outputs(3298) <= layer0_outputs(8761);
    layer1_outputs(3299) <= (layer0_outputs(7677)) or (layer0_outputs(1783));
    layer1_outputs(3300) <= (layer0_outputs(7807)) and (layer0_outputs(6392));
    layer1_outputs(3301) <= not((layer0_outputs(4046)) or (layer0_outputs(7918)));
    layer1_outputs(3302) <= (layer0_outputs(2303)) and not (layer0_outputs(7291));
    layer1_outputs(3303) <= (layer0_outputs(2644)) and (layer0_outputs(83));
    layer1_outputs(3304) <= not((layer0_outputs(6317)) and (layer0_outputs(856)));
    layer1_outputs(3305) <= '0';
    layer1_outputs(3306) <= '1';
    layer1_outputs(3307) <= not((layer0_outputs(7481)) or (layer0_outputs(471)));
    layer1_outputs(3308) <= (layer0_outputs(4240)) and not (layer0_outputs(3475));
    layer1_outputs(3309) <= (layer0_outputs(5917)) and not (layer0_outputs(776));
    layer1_outputs(3310) <= (layer0_outputs(6849)) and not (layer0_outputs(7171));
    layer1_outputs(3311) <= not(layer0_outputs(5083)) or (layer0_outputs(10034));
    layer1_outputs(3312) <= not(layer0_outputs(3281));
    layer1_outputs(3313) <= not((layer0_outputs(9441)) or (layer0_outputs(2313)));
    layer1_outputs(3314) <= layer0_outputs(10072);
    layer1_outputs(3315) <= not((layer0_outputs(4725)) and (layer0_outputs(1196)));
    layer1_outputs(3316) <= layer0_outputs(7696);
    layer1_outputs(3317) <= not(layer0_outputs(6866));
    layer1_outputs(3318) <= (layer0_outputs(5183)) and not (layer0_outputs(5244));
    layer1_outputs(3319) <= layer0_outputs(7120);
    layer1_outputs(3320) <= layer0_outputs(1020);
    layer1_outputs(3321) <= not(layer0_outputs(5733)) or (layer0_outputs(2888));
    layer1_outputs(3322) <= not((layer0_outputs(8255)) xor (layer0_outputs(8883)));
    layer1_outputs(3323) <= layer0_outputs(8673);
    layer1_outputs(3324) <= not(layer0_outputs(6994)) or (layer0_outputs(1977));
    layer1_outputs(3325) <= not(layer0_outputs(1250)) or (layer0_outputs(4214));
    layer1_outputs(3326) <= '1';
    layer1_outputs(3327) <= layer0_outputs(6551);
    layer1_outputs(3328) <= not((layer0_outputs(6783)) and (layer0_outputs(7854)));
    layer1_outputs(3329) <= (layer0_outputs(4374)) and not (layer0_outputs(3675));
    layer1_outputs(3330) <= layer0_outputs(6449);
    layer1_outputs(3331) <= not(layer0_outputs(8605));
    layer1_outputs(3332) <= layer0_outputs(5026);
    layer1_outputs(3333) <= not(layer0_outputs(6948));
    layer1_outputs(3334) <= not(layer0_outputs(8304));
    layer1_outputs(3335) <= (layer0_outputs(3648)) and not (layer0_outputs(3970));
    layer1_outputs(3336) <= not(layer0_outputs(4372));
    layer1_outputs(3337) <= not((layer0_outputs(4189)) xor (layer0_outputs(8164)));
    layer1_outputs(3338) <= layer0_outputs(6621);
    layer1_outputs(3339) <= (layer0_outputs(8504)) and not (layer0_outputs(2233));
    layer1_outputs(3340) <= (layer0_outputs(8718)) or (layer0_outputs(3470));
    layer1_outputs(3341) <= (layer0_outputs(376)) xor (layer0_outputs(4030));
    layer1_outputs(3342) <= '1';
    layer1_outputs(3343) <= not(layer0_outputs(7457)) or (layer0_outputs(5555));
    layer1_outputs(3344) <= not(layer0_outputs(4188));
    layer1_outputs(3345) <= not((layer0_outputs(5989)) xor (layer0_outputs(2495)));
    layer1_outputs(3346) <= (layer0_outputs(9036)) xor (layer0_outputs(4548));
    layer1_outputs(3347) <= not(layer0_outputs(2774));
    layer1_outputs(3348) <= layer0_outputs(8604);
    layer1_outputs(3349) <= not(layer0_outputs(875)) or (layer0_outputs(1970));
    layer1_outputs(3350) <= not(layer0_outputs(7464)) or (layer0_outputs(3145));
    layer1_outputs(3351) <= not((layer0_outputs(7355)) or (layer0_outputs(5230)));
    layer1_outputs(3352) <= '1';
    layer1_outputs(3353) <= layer0_outputs(4737);
    layer1_outputs(3354) <= layer0_outputs(5347);
    layer1_outputs(3355) <= not((layer0_outputs(1796)) or (layer0_outputs(5934)));
    layer1_outputs(3356) <= not(layer0_outputs(3976)) or (layer0_outputs(10149));
    layer1_outputs(3357) <= (layer0_outputs(1534)) and (layer0_outputs(3565));
    layer1_outputs(3358) <= (layer0_outputs(7317)) and not (layer0_outputs(1309));
    layer1_outputs(3359) <= (layer0_outputs(238)) xor (layer0_outputs(5976));
    layer1_outputs(3360) <= (layer0_outputs(375)) and (layer0_outputs(8686));
    layer1_outputs(3361) <= not((layer0_outputs(3868)) and (layer0_outputs(3485)));
    layer1_outputs(3362) <= layer0_outputs(9783);
    layer1_outputs(3363) <= not(layer0_outputs(4799));
    layer1_outputs(3364) <= not(layer0_outputs(1124));
    layer1_outputs(3365) <= (layer0_outputs(20)) and not (layer0_outputs(77));
    layer1_outputs(3366) <= '0';
    layer1_outputs(3367) <= not(layer0_outputs(2640)) or (layer0_outputs(2181));
    layer1_outputs(3368) <= not(layer0_outputs(4309));
    layer1_outputs(3369) <= '0';
    layer1_outputs(3370) <= not((layer0_outputs(855)) or (layer0_outputs(8996)));
    layer1_outputs(3371) <= not(layer0_outputs(3874));
    layer1_outputs(3372) <= not((layer0_outputs(3688)) xor (layer0_outputs(3273)));
    layer1_outputs(3373) <= layer0_outputs(2457);
    layer1_outputs(3374) <= (layer0_outputs(6980)) and (layer0_outputs(6493));
    layer1_outputs(3375) <= not(layer0_outputs(5447));
    layer1_outputs(3376) <= (layer0_outputs(673)) and not (layer0_outputs(8546));
    layer1_outputs(3377) <= layer0_outputs(7098);
    layer1_outputs(3378) <= layer0_outputs(8602);
    layer1_outputs(3379) <= (layer0_outputs(4701)) xor (layer0_outputs(8339));
    layer1_outputs(3380) <= (layer0_outputs(9447)) xor (layer0_outputs(7723));
    layer1_outputs(3381) <= '0';
    layer1_outputs(3382) <= layer0_outputs(2061);
    layer1_outputs(3383) <= (layer0_outputs(8982)) and not (layer0_outputs(3766));
    layer1_outputs(3384) <= layer0_outputs(1321);
    layer1_outputs(3385) <= not((layer0_outputs(90)) and (layer0_outputs(1092)));
    layer1_outputs(3386) <= not(layer0_outputs(8734));
    layer1_outputs(3387) <= layer0_outputs(4215);
    layer1_outputs(3388) <= (layer0_outputs(4159)) or (layer0_outputs(2898));
    layer1_outputs(3389) <= not((layer0_outputs(8259)) or (layer0_outputs(313)));
    layer1_outputs(3390) <= not(layer0_outputs(1637));
    layer1_outputs(3391) <= not((layer0_outputs(2922)) or (layer0_outputs(3456)));
    layer1_outputs(3392) <= (layer0_outputs(9728)) and not (layer0_outputs(3757));
    layer1_outputs(3393) <= not(layer0_outputs(1656));
    layer1_outputs(3394) <= not(layer0_outputs(7310));
    layer1_outputs(3395) <= (layer0_outputs(6438)) and not (layer0_outputs(3227));
    layer1_outputs(3396) <= (layer0_outputs(6339)) or (layer0_outputs(5290));
    layer1_outputs(3397) <= not((layer0_outputs(1063)) xor (layer0_outputs(4766)));
    layer1_outputs(3398) <= '0';
    layer1_outputs(3399) <= (layer0_outputs(7142)) and not (layer0_outputs(8422));
    layer1_outputs(3400) <= not(layer0_outputs(6407)) or (layer0_outputs(1703));
    layer1_outputs(3401) <= '1';
    layer1_outputs(3402) <= not(layer0_outputs(6397)) or (layer0_outputs(5059));
    layer1_outputs(3403) <= not((layer0_outputs(1868)) or (layer0_outputs(7917)));
    layer1_outputs(3404) <= (layer0_outputs(1078)) or (layer0_outputs(1022));
    layer1_outputs(3405) <= (layer0_outputs(3450)) and (layer0_outputs(10064));
    layer1_outputs(3406) <= not((layer0_outputs(2232)) xor (layer0_outputs(10145)));
    layer1_outputs(3407) <= not(layer0_outputs(2879));
    layer1_outputs(3408) <= not(layer0_outputs(9248)) or (layer0_outputs(1072));
    layer1_outputs(3409) <= (layer0_outputs(768)) or (layer0_outputs(3945));
    layer1_outputs(3410) <= not(layer0_outputs(4962)) or (layer0_outputs(1439));
    layer1_outputs(3411) <= not(layer0_outputs(9977));
    layer1_outputs(3412) <= '0';
    layer1_outputs(3413) <= (layer0_outputs(1824)) and not (layer0_outputs(7570));
    layer1_outputs(3414) <= (layer0_outputs(8126)) and not (layer0_outputs(3905));
    layer1_outputs(3415) <= not((layer0_outputs(1577)) and (layer0_outputs(2020)));
    layer1_outputs(3416) <= (layer0_outputs(1217)) and not (layer0_outputs(5459));
    layer1_outputs(3417) <= layer0_outputs(5264);
    layer1_outputs(3418) <= (layer0_outputs(6793)) or (layer0_outputs(9328));
    layer1_outputs(3419) <= not((layer0_outputs(6163)) and (layer0_outputs(5131)));
    layer1_outputs(3420) <= layer0_outputs(9408);
    layer1_outputs(3421) <= not(layer0_outputs(6196));
    layer1_outputs(3422) <= not((layer0_outputs(6842)) and (layer0_outputs(3685)));
    layer1_outputs(3423) <= not(layer0_outputs(5315)) or (layer0_outputs(2807));
    layer1_outputs(3424) <= not(layer0_outputs(8536)) or (layer0_outputs(9796));
    layer1_outputs(3425) <= layer0_outputs(393);
    layer1_outputs(3426) <= (layer0_outputs(1882)) and (layer0_outputs(5021));
    layer1_outputs(3427) <= '0';
    layer1_outputs(3428) <= not(layer0_outputs(3799)) or (layer0_outputs(1237));
    layer1_outputs(3429) <= not(layer0_outputs(9693));
    layer1_outputs(3430) <= (layer0_outputs(7346)) or (layer0_outputs(2201));
    layer1_outputs(3431) <= '0';
    layer1_outputs(3432) <= layer0_outputs(1461);
    layer1_outputs(3433) <= layer0_outputs(1954);
    layer1_outputs(3434) <= layer0_outputs(3806);
    layer1_outputs(3435) <= not(layer0_outputs(1564)) or (layer0_outputs(9743));
    layer1_outputs(3436) <= not((layer0_outputs(1014)) xor (layer0_outputs(6930)));
    layer1_outputs(3437) <= (layer0_outputs(7429)) or (layer0_outputs(208));
    layer1_outputs(3438) <= '0';
    layer1_outputs(3439) <= layer0_outputs(2873);
    layer1_outputs(3440) <= not(layer0_outputs(620));
    layer1_outputs(3441) <= not(layer0_outputs(5452)) or (layer0_outputs(9618));
    layer1_outputs(3442) <= layer0_outputs(7785);
    layer1_outputs(3443) <= not((layer0_outputs(6099)) and (layer0_outputs(9150)));
    layer1_outputs(3444) <= not(layer0_outputs(2144));
    layer1_outputs(3445) <= not(layer0_outputs(8637));
    layer1_outputs(3446) <= (layer0_outputs(3969)) xor (layer0_outputs(1694));
    layer1_outputs(3447) <= not(layer0_outputs(9550));
    layer1_outputs(3448) <= '1';
    layer1_outputs(3449) <= layer0_outputs(1823);
    layer1_outputs(3450) <= (layer0_outputs(5681)) and not (layer0_outputs(5298));
    layer1_outputs(3451) <= not(layer0_outputs(2029)) or (layer0_outputs(4936));
    layer1_outputs(3452) <= not(layer0_outputs(4707));
    layer1_outputs(3453) <= '1';
    layer1_outputs(3454) <= layer0_outputs(5510);
    layer1_outputs(3455) <= (layer0_outputs(8252)) or (layer0_outputs(6354));
    layer1_outputs(3456) <= not(layer0_outputs(7028));
    layer1_outputs(3457) <= not(layer0_outputs(3257)) or (layer0_outputs(2823));
    layer1_outputs(3458) <= '1';
    layer1_outputs(3459) <= not((layer0_outputs(3552)) or (layer0_outputs(5939)));
    layer1_outputs(3460) <= not(layer0_outputs(7511));
    layer1_outputs(3461) <= not(layer0_outputs(8812));
    layer1_outputs(3462) <= layer0_outputs(5305);
    layer1_outputs(3463) <= not(layer0_outputs(7430)) or (layer0_outputs(5332));
    layer1_outputs(3464) <= layer0_outputs(1632);
    layer1_outputs(3465) <= layer0_outputs(6862);
    layer1_outputs(3466) <= not(layer0_outputs(8020));
    layer1_outputs(3467) <= not(layer0_outputs(5004));
    layer1_outputs(3468) <= layer0_outputs(5046);
    layer1_outputs(3469) <= not(layer0_outputs(3591)) or (layer0_outputs(4605));
    layer1_outputs(3470) <= (layer0_outputs(7984)) and not (layer0_outputs(4203));
    layer1_outputs(3471) <= (layer0_outputs(10024)) xor (layer0_outputs(4979));
    layer1_outputs(3472) <= (layer0_outputs(10043)) or (layer0_outputs(9646));
    layer1_outputs(3473) <= not((layer0_outputs(9700)) or (layer0_outputs(7840)));
    layer1_outputs(3474) <= not((layer0_outputs(8096)) xor (layer0_outputs(5606)));
    layer1_outputs(3475) <= not(layer0_outputs(3302)) or (layer0_outputs(356));
    layer1_outputs(3476) <= '1';
    layer1_outputs(3477) <= not(layer0_outputs(3724));
    layer1_outputs(3478) <= (layer0_outputs(599)) xor (layer0_outputs(9900));
    layer1_outputs(3479) <= not((layer0_outputs(8797)) and (layer0_outputs(4243)));
    layer1_outputs(3480) <= not((layer0_outputs(5786)) or (layer0_outputs(2897)));
    layer1_outputs(3481) <= (layer0_outputs(3160)) and (layer0_outputs(9154));
    layer1_outputs(3482) <= (layer0_outputs(195)) and (layer0_outputs(8904));
    layer1_outputs(3483) <= not(layer0_outputs(9984)) or (layer0_outputs(6720));
    layer1_outputs(3484) <= layer0_outputs(1574);
    layer1_outputs(3485) <= layer0_outputs(4760);
    layer1_outputs(3486) <= not((layer0_outputs(2438)) and (layer0_outputs(6437)));
    layer1_outputs(3487) <= not(layer0_outputs(8503)) or (layer0_outputs(9873));
    layer1_outputs(3488) <= not(layer0_outputs(7505));
    layer1_outputs(3489) <= not(layer0_outputs(7636));
    layer1_outputs(3490) <= (layer0_outputs(9697)) or (layer0_outputs(9542));
    layer1_outputs(3491) <= not(layer0_outputs(8827));
    layer1_outputs(3492) <= (layer0_outputs(2958)) or (layer0_outputs(2417));
    layer1_outputs(3493) <= layer0_outputs(5947);
    layer1_outputs(3494) <= not(layer0_outputs(10002));
    layer1_outputs(3495) <= (layer0_outputs(6759)) and not (layer0_outputs(4359));
    layer1_outputs(3496) <= layer0_outputs(5650);
    layer1_outputs(3497) <= not((layer0_outputs(821)) and (layer0_outputs(6792)));
    layer1_outputs(3498) <= not(layer0_outputs(6325)) or (layer0_outputs(5885));
    layer1_outputs(3499) <= (layer0_outputs(453)) and (layer0_outputs(9450));
    layer1_outputs(3500) <= not(layer0_outputs(8765));
    layer1_outputs(3501) <= '1';
    layer1_outputs(3502) <= not(layer0_outputs(11));
    layer1_outputs(3503) <= not(layer0_outputs(6771)) or (layer0_outputs(8523));
    layer1_outputs(3504) <= layer0_outputs(8630);
    layer1_outputs(3505) <= '1';
    layer1_outputs(3506) <= layer0_outputs(2013);
    layer1_outputs(3507) <= not(layer0_outputs(1304));
    layer1_outputs(3508) <= (layer0_outputs(4592)) and (layer0_outputs(6994));
    layer1_outputs(3509) <= not((layer0_outputs(9483)) and (layer0_outputs(1254)));
    layer1_outputs(3510) <= not((layer0_outputs(3461)) xor (layer0_outputs(8955)));
    layer1_outputs(3511) <= (layer0_outputs(5028)) and not (layer0_outputs(9465));
    layer1_outputs(3512) <= not((layer0_outputs(8403)) or (layer0_outputs(8865)));
    layer1_outputs(3513) <= layer0_outputs(5292);
    layer1_outputs(3514) <= (layer0_outputs(3593)) and not (layer0_outputs(4168));
    layer1_outputs(3515) <= layer0_outputs(9932);
    layer1_outputs(3516) <= not((layer0_outputs(3269)) or (layer0_outputs(4561)));
    layer1_outputs(3517) <= (layer0_outputs(1307)) and (layer0_outputs(5432));
    layer1_outputs(3518) <= (layer0_outputs(5505)) and not (layer0_outputs(1359));
    layer1_outputs(3519) <= not((layer0_outputs(2903)) and (layer0_outputs(5564)));
    layer1_outputs(3520) <= not(layer0_outputs(1538)) or (layer0_outputs(9476));
    layer1_outputs(3521) <= (layer0_outputs(9477)) and (layer0_outputs(7785));
    layer1_outputs(3522) <= not(layer0_outputs(2400)) or (layer0_outputs(8697));
    layer1_outputs(3523) <= not(layer0_outputs(1370));
    layer1_outputs(3524) <= not((layer0_outputs(9336)) and (layer0_outputs(4539)));
    layer1_outputs(3525) <= not(layer0_outputs(82)) or (layer0_outputs(5262));
    layer1_outputs(3526) <= '0';
    layer1_outputs(3527) <= (layer0_outputs(2076)) and (layer0_outputs(4487));
    layer1_outputs(3528) <= (layer0_outputs(4381)) or (layer0_outputs(1658));
    layer1_outputs(3529) <= (layer0_outputs(651)) or (layer0_outputs(90));
    layer1_outputs(3530) <= not(layer0_outputs(8502)) or (layer0_outputs(5830));
    layer1_outputs(3531) <= layer0_outputs(6953);
    layer1_outputs(3532) <= '0';
    layer1_outputs(3533) <= not((layer0_outputs(4293)) or (layer0_outputs(3740)));
    layer1_outputs(3534) <= (layer0_outputs(10150)) and not (layer0_outputs(807));
    layer1_outputs(3535) <= '1';
    layer1_outputs(3536) <= (layer0_outputs(626)) and not (layer0_outputs(7059));
    layer1_outputs(3537) <= layer0_outputs(6046);
    layer1_outputs(3538) <= (layer0_outputs(6614)) and (layer0_outputs(7826));
    layer1_outputs(3539) <= not(layer0_outputs(5547));
    layer1_outputs(3540) <= layer0_outputs(2997);
    layer1_outputs(3541) <= not((layer0_outputs(8909)) xor (layer0_outputs(2593)));
    layer1_outputs(3542) <= not(layer0_outputs(5530)) or (layer0_outputs(4019));
    layer1_outputs(3543) <= not((layer0_outputs(8817)) or (layer0_outputs(8120)));
    layer1_outputs(3544) <= '0';
    layer1_outputs(3545) <= (layer0_outputs(5582)) and not (layer0_outputs(6423));
    layer1_outputs(3546) <= not(layer0_outputs(9556));
    layer1_outputs(3547) <= (layer0_outputs(7924)) or (layer0_outputs(3859));
    layer1_outputs(3548) <= layer0_outputs(3847);
    layer1_outputs(3549) <= (layer0_outputs(220)) or (layer0_outputs(2059));
    layer1_outputs(3550) <= (layer0_outputs(4867)) or (layer0_outputs(4066));
    layer1_outputs(3551) <= layer0_outputs(9854);
    layer1_outputs(3552) <= not(layer0_outputs(7327));
    layer1_outputs(3553) <= not((layer0_outputs(772)) and (layer0_outputs(3460)));
    layer1_outputs(3554) <= layer0_outputs(3843);
    layer1_outputs(3555) <= (layer0_outputs(164)) and not (layer0_outputs(7832));
    layer1_outputs(3556) <= not((layer0_outputs(2717)) or (layer0_outputs(6117)));
    layer1_outputs(3557) <= layer0_outputs(516);
    layer1_outputs(3558) <= not((layer0_outputs(9346)) or (layer0_outputs(5861)));
    layer1_outputs(3559) <= not(layer0_outputs(10061));
    layer1_outputs(3560) <= not((layer0_outputs(7896)) and (layer0_outputs(2128)));
    layer1_outputs(3561) <= not((layer0_outputs(7128)) and (layer0_outputs(3009)));
    layer1_outputs(3562) <= not((layer0_outputs(6744)) xor (layer0_outputs(8890)));
    layer1_outputs(3563) <= layer0_outputs(2201);
    layer1_outputs(3564) <= layer0_outputs(5583);
    layer1_outputs(3565) <= not(layer0_outputs(7504)) or (layer0_outputs(6444));
    layer1_outputs(3566) <= layer0_outputs(7879);
    layer1_outputs(3567) <= '0';
    layer1_outputs(3568) <= not(layer0_outputs(6835));
    layer1_outputs(3569) <= not(layer0_outputs(3774));
    layer1_outputs(3570) <= (layer0_outputs(5038)) and not (layer0_outputs(3923));
    layer1_outputs(3571) <= not(layer0_outputs(8657));
    layer1_outputs(3572) <= layer0_outputs(7280);
    layer1_outputs(3573) <= (layer0_outputs(9934)) and not (layer0_outputs(329));
    layer1_outputs(3574) <= (layer0_outputs(6845)) and not (layer0_outputs(1645));
    layer1_outputs(3575) <= not(layer0_outputs(1634)) or (layer0_outputs(8975));
    layer1_outputs(3576) <= (layer0_outputs(8417)) or (layer0_outputs(8562));
    layer1_outputs(3577) <= '1';
    layer1_outputs(3578) <= not(layer0_outputs(7688));
    layer1_outputs(3579) <= (layer0_outputs(4128)) and not (layer0_outputs(4218));
    layer1_outputs(3580) <= not(layer0_outputs(1896));
    layer1_outputs(3581) <= layer0_outputs(6026);
    layer1_outputs(3582) <= layer0_outputs(7815);
    layer1_outputs(3583) <= not(layer0_outputs(8566)) or (layer0_outputs(6653));
    layer1_outputs(3584) <= layer0_outputs(394);
    layer1_outputs(3585) <= (layer0_outputs(1639)) or (layer0_outputs(293));
    layer1_outputs(3586) <= '1';
    layer1_outputs(3587) <= (layer0_outputs(2297)) and not (layer0_outputs(2328));
    layer1_outputs(3588) <= not(layer0_outputs(8460));
    layer1_outputs(3589) <= layer0_outputs(7303);
    layer1_outputs(3590) <= '1';
    layer1_outputs(3591) <= not(layer0_outputs(8689));
    layer1_outputs(3592) <= not((layer0_outputs(1921)) xor (layer0_outputs(1623)));
    layer1_outputs(3593) <= not(layer0_outputs(3142)) or (layer0_outputs(7682));
    layer1_outputs(3594) <= (layer0_outputs(5694)) xor (layer0_outputs(4059));
    layer1_outputs(3595) <= not((layer0_outputs(7693)) or (layer0_outputs(9847)));
    layer1_outputs(3596) <= not(layer0_outputs(8551));
    layer1_outputs(3597) <= not((layer0_outputs(6154)) and (layer0_outputs(9170)));
    layer1_outputs(3598) <= not((layer0_outputs(3844)) or (layer0_outputs(2459)));
    layer1_outputs(3599) <= (layer0_outputs(3457)) and not (layer0_outputs(2849));
    layer1_outputs(3600) <= not(layer0_outputs(7881));
    layer1_outputs(3601) <= (layer0_outputs(2657)) or (layer0_outputs(3428));
    layer1_outputs(3602) <= not(layer0_outputs(1826));
    layer1_outputs(3603) <= not((layer0_outputs(933)) and (layer0_outputs(4732)));
    layer1_outputs(3604) <= not((layer0_outputs(2663)) and (layer0_outputs(10041)));
    layer1_outputs(3605) <= (layer0_outputs(6331)) or (layer0_outputs(8248));
    layer1_outputs(3606) <= layer0_outputs(824);
    layer1_outputs(3607) <= not(layer0_outputs(4727)) or (layer0_outputs(2926));
    layer1_outputs(3608) <= (layer0_outputs(9734)) and (layer0_outputs(4813));
    layer1_outputs(3609) <= (layer0_outputs(6249)) xor (layer0_outputs(2620));
    layer1_outputs(3610) <= layer0_outputs(3052);
    layer1_outputs(3611) <= not(layer0_outputs(2316));
    layer1_outputs(3612) <= (layer0_outputs(6688)) and not (layer0_outputs(5241));
    layer1_outputs(3613) <= not(layer0_outputs(2676));
    layer1_outputs(3614) <= (layer0_outputs(3790)) and not (layer0_outputs(8970));
    layer1_outputs(3615) <= not(layer0_outputs(916)) or (layer0_outputs(944));
    layer1_outputs(3616) <= (layer0_outputs(4213)) or (layer0_outputs(2011));
    layer1_outputs(3617) <= not((layer0_outputs(4917)) or (layer0_outputs(4388)));
    layer1_outputs(3618) <= not((layer0_outputs(7973)) and (layer0_outputs(8044)));
    layer1_outputs(3619) <= not((layer0_outputs(877)) xor (layer0_outputs(8106)));
    layer1_outputs(3620) <= not(layer0_outputs(6181));
    layer1_outputs(3621) <= not(layer0_outputs(5378));
    layer1_outputs(3622) <= not(layer0_outputs(180));
    layer1_outputs(3623) <= not(layer0_outputs(1811)) or (layer0_outputs(3666));
    layer1_outputs(3624) <= layer0_outputs(9722);
    layer1_outputs(3625) <= (layer0_outputs(32)) and not (layer0_outputs(9334));
    layer1_outputs(3626) <= layer0_outputs(1204);
    layer1_outputs(3627) <= (layer0_outputs(10020)) or (layer0_outputs(2840));
    layer1_outputs(3628) <= '0';
    layer1_outputs(3629) <= (layer0_outputs(958)) and not (layer0_outputs(2208));
    layer1_outputs(3630) <= not(layer0_outputs(1499));
    layer1_outputs(3631) <= not((layer0_outputs(6584)) or (layer0_outputs(4777)));
    layer1_outputs(3632) <= not((layer0_outputs(6896)) or (layer0_outputs(3247)));
    layer1_outputs(3633) <= not(layer0_outputs(1997)) or (layer0_outputs(6364));
    layer1_outputs(3634) <= (layer0_outputs(10154)) xor (layer0_outputs(71));
    layer1_outputs(3635) <= (layer0_outputs(8364)) or (layer0_outputs(723));
    layer1_outputs(3636) <= not(layer0_outputs(5436)) or (layer0_outputs(58));
    layer1_outputs(3637) <= not((layer0_outputs(7456)) or (layer0_outputs(1352)));
    layer1_outputs(3638) <= not(layer0_outputs(5616)) or (layer0_outputs(2642));
    layer1_outputs(3639) <= (layer0_outputs(5816)) and not (layer0_outputs(4916));
    layer1_outputs(3640) <= (layer0_outputs(8837)) and not (layer0_outputs(1779));
    layer1_outputs(3641) <= (layer0_outputs(5961)) xor (layer0_outputs(6628));
    layer1_outputs(3642) <= not((layer0_outputs(7906)) and (layer0_outputs(9122)));
    layer1_outputs(3643) <= layer0_outputs(9031);
    layer1_outputs(3644) <= (layer0_outputs(7988)) or (layer0_outputs(1244));
    layer1_outputs(3645) <= not((layer0_outputs(777)) xor (layer0_outputs(4649)));
    layer1_outputs(3646) <= not((layer0_outputs(6199)) and (layer0_outputs(6055)));
    layer1_outputs(3647) <= (layer0_outputs(7602)) and not (layer0_outputs(6856));
    layer1_outputs(3648) <= layer0_outputs(6463);
    layer1_outputs(3649) <= not(layer0_outputs(1746)) or (layer0_outputs(6916));
    layer1_outputs(3650) <= layer0_outputs(5963);
    layer1_outputs(3651) <= not(layer0_outputs(5266)) or (layer0_outputs(3381));
    layer1_outputs(3652) <= (layer0_outputs(1626)) or (layer0_outputs(7540));
    layer1_outputs(3653) <= (layer0_outputs(8273)) and not (layer0_outputs(4870));
    layer1_outputs(3654) <= not((layer0_outputs(4101)) xor (layer0_outputs(8608)));
    layer1_outputs(3655) <= not(layer0_outputs(8330));
    layer1_outputs(3656) <= not((layer0_outputs(5152)) xor (layer0_outputs(5180)));
    layer1_outputs(3657) <= layer0_outputs(6046);
    layer1_outputs(3658) <= (layer0_outputs(8780)) and not (layer0_outputs(5426));
    layer1_outputs(3659) <= not(layer0_outputs(6327));
    layer1_outputs(3660) <= not(layer0_outputs(9731)) or (layer0_outputs(43));
    layer1_outputs(3661) <= not(layer0_outputs(2526));
    layer1_outputs(3662) <= layer0_outputs(2395);
    layer1_outputs(3663) <= not(layer0_outputs(7187));
    layer1_outputs(3664) <= layer0_outputs(7665);
    layer1_outputs(3665) <= layer0_outputs(9706);
    layer1_outputs(3666) <= layer0_outputs(9688);
    layer1_outputs(3667) <= not(layer0_outputs(1881));
    layer1_outputs(3668) <= '0';
    layer1_outputs(3669) <= not((layer0_outputs(4505)) xor (layer0_outputs(2243)));
    layer1_outputs(3670) <= '1';
    layer1_outputs(3671) <= layer0_outputs(8676);
    layer1_outputs(3672) <= (layer0_outputs(6685)) and (layer0_outputs(2083));
    layer1_outputs(3673) <= not(layer0_outputs(3091)) or (layer0_outputs(4671));
    layer1_outputs(3674) <= not(layer0_outputs(414)) or (layer0_outputs(7876));
    layer1_outputs(3675) <= not((layer0_outputs(8689)) xor (layer0_outputs(5468)));
    layer1_outputs(3676) <= not(layer0_outputs(10002));
    layer1_outputs(3677) <= not(layer0_outputs(2277)) or (layer0_outputs(5773));
    layer1_outputs(3678) <= (layer0_outputs(4400)) or (layer0_outputs(724));
    layer1_outputs(3679) <= layer0_outputs(9994);
    layer1_outputs(3680) <= layer0_outputs(4204);
    layer1_outputs(3681) <= '0';
    layer1_outputs(3682) <= not(layer0_outputs(3612)) or (layer0_outputs(3787));
    layer1_outputs(3683) <= not(layer0_outputs(2961));
    layer1_outputs(3684) <= (layer0_outputs(8078)) or (layer0_outputs(8613));
    layer1_outputs(3685) <= (layer0_outputs(5103)) and (layer0_outputs(3323));
    layer1_outputs(3686) <= not(layer0_outputs(4515));
    layer1_outputs(3687) <= (layer0_outputs(6031)) and not (layer0_outputs(2566));
    layer1_outputs(3688) <= (layer0_outputs(6571)) xor (layer0_outputs(1373));
    layer1_outputs(3689) <= not(layer0_outputs(9926)) or (layer0_outputs(5219));
    layer1_outputs(3690) <= not(layer0_outputs(4081));
    layer1_outputs(3691) <= not((layer0_outputs(10117)) xor (layer0_outputs(9829)));
    layer1_outputs(3692) <= not(layer0_outputs(3156));
    layer1_outputs(3693) <= (layer0_outputs(5299)) or (layer0_outputs(3530));
    layer1_outputs(3694) <= (layer0_outputs(5382)) and not (layer0_outputs(4621));
    layer1_outputs(3695) <= (layer0_outputs(7073)) and not (layer0_outputs(9219));
    layer1_outputs(3696) <= (layer0_outputs(9620)) and (layer0_outputs(6365));
    layer1_outputs(3697) <= not(layer0_outputs(7276));
    layer1_outputs(3698) <= (layer0_outputs(5660)) and not (layer0_outputs(3757));
    layer1_outputs(3699) <= not(layer0_outputs(7439));
    layer1_outputs(3700) <= (layer0_outputs(8291)) or (layer0_outputs(4861));
    layer1_outputs(3701) <= not(layer0_outputs(3100));
    layer1_outputs(3702) <= not(layer0_outputs(9457)) or (layer0_outputs(5159));
    layer1_outputs(3703) <= not(layer0_outputs(4634)) or (layer0_outputs(1951));
    layer1_outputs(3704) <= not(layer0_outputs(2860)) or (layer0_outputs(2038));
    layer1_outputs(3705) <= '0';
    layer1_outputs(3706) <= (layer0_outputs(5302)) or (layer0_outputs(3246));
    layer1_outputs(3707) <= (layer0_outputs(1261)) and not (layer0_outputs(5092));
    layer1_outputs(3708) <= (layer0_outputs(5931)) and not (layer0_outputs(8968));
    layer1_outputs(3709) <= (layer0_outputs(1059)) or (layer0_outputs(5018));
    layer1_outputs(3710) <= (layer0_outputs(7751)) and not (layer0_outputs(2342));
    layer1_outputs(3711) <= (layer0_outputs(6698)) and (layer0_outputs(2675));
    layer1_outputs(3712) <= not(layer0_outputs(4100)) or (layer0_outputs(6612));
    layer1_outputs(3713) <= (layer0_outputs(2752)) and (layer0_outputs(5529));
    layer1_outputs(3714) <= layer0_outputs(2733);
    layer1_outputs(3715) <= '1';
    layer1_outputs(3716) <= not(layer0_outputs(6727)) or (layer0_outputs(2901));
    layer1_outputs(3717) <= (layer0_outputs(9299)) and (layer0_outputs(8199));
    layer1_outputs(3718) <= not(layer0_outputs(4638));
    layer1_outputs(3719) <= layer0_outputs(8393);
    layer1_outputs(3720) <= not(layer0_outputs(9061)) or (layer0_outputs(5400));
    layer1_outputs(3721) <= layer0_outputs(2847);
    layer1_outputs(3722) <= (layer0_outputs(7898)) and not (layer0_outputs(3793));
    layer1_outputs(3723) <= (layer0_outputs(6223)) xor (layer0_outputs(5281));
    layer1_outputs(3724) <= (layer0_outputs(9715)) and not (layer0_outputs(2439));
    layer1_outputs(3725) <= (layer0_outputs(8382)) or (layer0_outputs(7474));
    layer1_outputs(3726) <= layer0_outputs(7449);
    layer1_outputs(3727) <= layer0_outputs(4805);
    layer1_outputs(3728) <= not(layer0_outputs(8477)) or (layer0_outputs(6433));
    layer1_outputs(3729) <= layer0_outputs(2744);
    layer1_outputs(3730) <= not((layer0_outputs(9374)) or (layer0_outputs(4775)));
    layer1_outputs(3731) <= not(layer0_outputs(5093)) or (layer0_outputs(1135));
    layer1_outputs(3732) <= not(layer0_outputs(7663));
    layer1_outputs(3733) <= '0';
    layer1_outputs(3734) <= not(layer0_outputs(3126));
    layer1_outputs(3735) <= not((layer0_outputs(6012)) and (layer0_outputs(5273)));
    layer1_outputs(3736) <= '0';
    layer1_outputs(3737) <= not(layer0_outputs(4424));
    layer1_outputs(3738) <= not(layer0_outputs(3358)) or (layer0_outputs(6235));
    layer1_outputs(3739) <= not((layer0_outputs(9698)) xor (layer0_outputs(5131)));
    layer1_outputs(3740) <= (layer0_outputs(1514)) xor (layer0_outputs(353));
    layer1_outputs(3741) <= (layer0_outputs(630)) xor (layer0_outputs(2367));
    layer1_outputs(3742) <= not(layer0_outputs(3622));
    layer1_outputs(3743) <= (layer0_outputs(2409)) and (layer0_outputs(4727));
    layer1_outputs(3744) <= not(layer0_outputs(8012));
    layer1_outputs(3745) <= (layer0_outputs(1660)) xor (layer0_outputs(5015));
    layer1_outputs(3746) <= (layer0_outputs(1464)) xor (layer0_outputs(8152));
    layer1_outputs(3747) <= not(layer0_outputs(9229));
    layer1_outputs(3748) <= not(layer0_outputs(3305));
    layer1_outputs(3749) <= not(layer0_outputs(1476));
    layer1_outputs(3750) <= not(layer0_outputs(6336));
    layer1_outputs(3751) <= not((layer0_outputs(7297)) and (layer0_outputs(8112)));
    layer1_outputs(3752) <= not((layer0_outputs(5142)) or (layer0_outputs(4928)));
    layer1_outputs(3753) <= not(layer0_outputs(4888)) or (layer0_outputs(6308));
    layer1_outputs(3754) <= (layer0_outputs(10005)) and not (layer0_outputs(51));
    layer1_outputs(3755) <= layer0_outputs(6440);
    layer1_outputs(3756) <= (layer0_outputs(5616)) and not (layer0_outputs(2455));
    layer1_outputs(3757) <= '0';
    layer1_outputs(3758) <= layer0_outputs(5881);
    layer1_outputs(3759) <= layer0_outputs(3494);
    layer1_outputs(3760) <= '0';
    layer1_outputs(3761) <= '1';
    layer1_outputs(3762) <= not(layer0_outputs(370));
    layer1_outputs(3763) <= (layer0_outputs(1548)) and not (layer0_outputs(6848));
    layer1_outputs(3764) <= not((layer0_outputs(6042)) and (layer0_outputs(2375)));
    layer1_outputs(3765) <= '0';
    layer1_outputs(3766) <= not(layer0_outputs(266)) or (layer0_outputs(435));
    layer1_outputs(3767) <= '0';
    layer1_outputs(3768) <= not(layer0_outputs(5801)) or (layer0_outputs(946));
    layer1_outputs(3769) <= not(layer0_outputs(7944));
    layer1_outputs(3770) <= (layer0_outputs(6251)) and (layer0_outputs(437));
    layer1_outputs(3771) <= not(layer0_outputs(8745));
    layer1_outputs(3772) <= '1';
    layer1_outputs(3773) <= not((layer0_outputs(3984)) and (layer0_outputs(381)));
    layer1_outputs(3774) <= layer0_outputs(5424);
    layer1_outputs(3775) <= (layer0_outputs(3833)) and not (layer0_outputs(2461));
    layer1_outputs(3776) <= not((layer0_outputs(7393)) or (layer0_outputs(8088)));
    layer1_outputs(3777) <= not(layer0_outputs(7829));
    layer1_outputs(3778) <= not((layer0_outputs(7274)) xor (layer0_outputs(2310)));
    layer1_outputs(3779) <= '1';
    layer1_outputs(3780) <= (layer0_outputs(9676)) and (layer0_outputs(5401));
    layer1_outputs(3781) <= not(layer0_outputs(6228));
    layer1_outputs(3782) <= not(layer0_outputs(7300));
    layer1_outputs(3783) <= (layer0_outputs(1442)) and not (layer0_outputs(7555));
    layer1_outputs(3784) <= not(layer0_outputs(9689));
    layer1_outputs(3785) <= '1';
    layer1_outputs(3786) <= not((layer0_outputs(5016)) and (layer0_outputs(9818)));
    layer1_outputs(3787) <= (layer0_outputs(4938)) xor (layer0_outputs(9806));
    layer1_outputs(3788) <= (layer0_outputs(4250)) and (layer0_outputs(7363));
    layer1_outputs(3789) <= not((layer0_outputs(10227)) and (layer0_outputs(3621)));
    layer1_outputs(3790) <= (layer0_outputs(951)) and not (layer0_outputs(683));
    layer1_outputs(3791) <= not(layer0_outputs(5417));
    layer1_outputs(3792) <= not(layer0_outputs(1316)) or (layer0_outputs(7833));
    layer1_outputs(3793) <= not(layer0_outputs(999));
    layer1_outputs(3794) <= (layer0_outputs(5979)) xor (layer0_outputs(5987));
    layer1_outputs(3795) <= not(layer0_outputs(1003)) or (layer0_outputs(5523));
    layer1_outputs(3796) <= (layer0_outputs(1793)) and (layer0_outputs(4864));
    layer1_outputs(3797) <= not((layer0_outputs(9261)) xor (layer0_outputs(8869)));
    layer1_outputs(3798) <= not(layer0_outputs(1322)) or (layer0_outputs(3435));
    layer1_outputs(3799) <= (layer0_outputs(7868)) and (layer0_outputs(9963));
    layer1_outputs(3800) <= not((layer0_outputs(2562)) or (layer0_outputs(4915)));
    layer1_outputs(3801) <= (layer0_outputs(5116)) and not (layer0_outputs(3513));
    layer1_outputs(3802) <= not((layer0_outputs(7674)) and (layer0_outputs(8460)));
    layer1_outputs(3803) <= (layer0_outputs(2867)) and not (layer0_outputs(7123));
    layer1_outputs(3804) <= (layer0_outputs(679)) xor (layer0_outputs(8410));
    layer1_outputs(3805) <= (layer0_outputs(1427)) xor (layer0_outputs(4041));
    layer1_outputs(3806) <= layer0_outputs(9936);
    layer1_outputs(3807) <= (layer0_outputs(3260)) and not (layer0_outputs(9246));
    layer1_outputs(3808) <= '0';
    layer1_outputs(3809) <= not((layer0_outputs(1481)) xor (layer0_outputs(3025)));
    layer1_outputs(3810) <= not(layer0_outputs(6679));
    layer1_outputs(3811) <= not((layer0_outputs(5561)) and (layer0_outputs(2024)));
    layer1_outputs(3812) <= not(layer0_outputs(8667));
    layer1_outputs(3813) <= layer0_outputs(3645);
    layer1_outputs(3814) <= layer0_outputs(8317);
    layer1_outputs(3815) <= (layer0_outputs(1736)) and not (layer0_outputs(5121));
    layer1_outputs(3816) <= layer0_outputs(1487);
    layer1_outputs(3817) <= not((layer0_outputs(78)) and (layer0_outputs(6745)));
    layer1_outputs(3818) <= not(layer0_outputs(5205)) or (layer0_outputs(6367));
    layer1_outputs(3819) <= (layer0_outputs(1875)) and not (layer0_outputs(6315));
    layer1_outputs(3820) <= layer0_outputs(7560);
    layer1_outputs(3821) <= not(layer0_outputs(2067)) or (layer0_outputs(8574));
    layer1_outputs(3822) <= (layer0_outputs(6887)) and not (layer0_outputs(9651));
    layer1_outputs(3823) <= not((layer0_outputs(7405)) and (layer0_outputs(8829)));
    layer1_outputs(3824) <= layer0_outputs(10026);
    layer1_outputs(3825) <= layer0_outputs(2257);
    layer1_outputs(3826) <= not(layer0_outputs(6545)) or (layer0_outputs(8035));
    layer1_outputs(3827) <= not(layer0_outputs(5409));
    layer1_outputs(3828) <= layer0_outputs(8416);
    layer1_outputs(3829) <= not(layer0_outputs(5433));
    layer1_outputs(3830) <= (layer0_outputs(7214)) and not (layer0_outputs(10018));
    layer1_outputs(3831) <= (layer0_outputs(2982)) and not (layer0_outputs(3813));
    layer1_outputs(3832) <= (layer0_outputs(3489)) and not (layer0_outputs(8201));
    layer1_outputs(3833) <= not(layer0_outputs(4378));
    layer1_outputs(3834) <= layer0_outputs(2058);
    layer1_outputs(3835) <= not(layer0_outputs(3360)) or (layer0_outputs(8054));
    layer1_outputs(3836) <= not((layer0_outputs(6885)) or (layer0_outputs(2154)));
    layer1_outputs(3837) <= '1';
    layer1_outputs(3838) <= layer0_outputs(82);
    layer1_outputs(3839) <= (layer0_outputs(3690)) and (layer0_outputs(1936));
    layer1_outputs(3840) <= not(layer0_outputs(6320));
    layer1_outputs(3841) <= not(layer0_outputs(3768));
    layer1_outputs(3842) <= not(layer0_outputs(6305));
    layer1_outputs(3843) <= not(layer0_outputs(8224)) or (layer0_outputs(1816));
    layer1_outputs(3844) <= '0';
    layer1_outputs(3845) <= '0';
    layer1_outputs(3846) <= not((layer0_outputs(10238)) or (layer0_outputs(8336)));
    layer1_outputs(3847) <= (layer0_outputs(8453)) and (layer0_outputs(3699));
    layer1_outputs(3848) <= layer0_outputs(5983);
    layer1_outputs(3849) <= not(layer0_outputs(4807));
    layer1_outputs(3850) <= not(layer0_outputs(2600));
    layer1_outputs(3851) <= not(layer0_outputs(215));
    layer1_outputs(3852) <= not((layer0_outputs(6725)) or (layer0_outputs(5827)));
    layer1_outputs(3853) <= (layer0_outputs(7279)) or (layer0_outputs(5405));
    layer1_outputs(3854) <= (layer0_outputs(3448)) and not (layer0_outputs(1481));
    layer1_outputs(3855) <= not(layer0_outputs(1));
    layer1_outputs(3856) <= layer0_outputs(2547);
    layer1_outputs(3857) <= (layer0_outputs(5628)) and (layer0_outputs(4343));
    layer1_outputs(3858) <= (layer0_outputs(9995)) and not (layer0_outputs(9173));
    layer1_outputs(3859) <= layer0_outputs(9);
    layer1_outputs(3860) <= layer0_outputs(943);
    layer1_outputs(3861) <= layer0_outputs(3512);
    layer1_outputs(3862) <= not(layer0_outputs(10162));
    layer1_outputs(3863) <= (layer0_outputs(3820)) and (layer0_outputs(2507));
    layer1_outputs(3864) <= (layer0_outputs(7873)) or (layer0_outputs(4608));
    layer1_outputs(3865) <= (layer0_outputs(884)) and (layer0_outputs(246));
    layer1_outputs(3866) <= not(layer0_outputs(2001)) or (layer0_outputs(360));
    layer1_outputs(3867) <= '1';
    layer1_outputs(3868) <= not(layer0_outputs(6283)) or (layer0_outputs(469));
    layer1_outputs(3869) <= not((layer0_outputs(4894)) or (layer0_outputs(343)));
    layer1_outputs(3870) <= not(layer0_outputs(6473));
    layer1_outputs(3871) <= layer0_outputs(9392);
    layer1_outputs(3872) <= '1';
    layer1_outputs(3873) <= layer0_outputs(7703);
    layer1_outputs(3874) <= not((layer0_outputs(8280)) xor (layer0_outputs(6020)));
    layer1_outputs(3875) <= not(layer0_outputs(4051));
    layer1_outputs(3876) <= not(layer0_outputs(3415)) or (layer0_outputs(1830));
    layer1_outputs(3877) <= (layer0_outputs(5238)) or (layer0_outputs(3321));
    layer1_outputs(3878) <= layer0_outputs(2127);
    layer1_outputs(3879) <= not((layer0_outputs(40)) or (layer0_outputs(8169)));
    layer1_outputs(3880) <= not((layer0_outputs(6536)) and (layer0_outputs(1266)));
    layer1_outputs(3881) <= (layer0_outputs(10191)) and not (layer0_outputs(3538));
    layer1_outputs(3882) <= (layer0_outputs(907)) and (layer0_outputs(6513));
    layer1_outputs(3883) <= '0';
    layer1_outputs(3884) <= (layer0_outputs(6486)) and (layer0_outputs(8685));
    layer1_outputs(3885) <= '1';
    layer1_outputs(3886) <= not(layer0_outputs(1165));
    layer1_outputs(3887) <= (layer0_outputs(5073)) and (layer0_outputs(7284));
    layer1_outputs(3888) <= not(layer0_outputs(8738)) or (layer0_outputs(5220));
    layer1_outputs(3889) <= '0';
    layer1_outputs(3890) <= '1';
    layer1_outputs(3891) <= not((layer0_outputs(6992)) or (layer0_outputs(563)));
    layer1_outputs(3892) <= layer0_outputs(1707);
    layer1_outputs(3893) <= not(layer0_outputs(3550));
    layer1_outputs(3894) <= not(layer0_outputs(8804));
    layer1_outputs(3895) <= not((layer0_outputs(4121)) xor (layer0_outputs(147)));
    layer1_outputs(3896) <= (layer0_outputs(4737)) and not (layer0_outputs(1344));
    layer1_outputs(3897) <= (layer0_outputs(2358)) and not (layer0_outputs(1084));
    layer1_outputs(3898) <= layer0_outputs(6827);
    layer1_outputs(3899) <= (layer0_outputs(9923)) and (layer0_outputs(4931));
    layer1_outputs(3900) <= not(layer0_outputs(9308));
    layer1_outputs(3901) <= (layer0_outputs(6909)) xor (layer0_outputs(2108));
    layer1_outputs(3902) <= not(layer0_outputs(6499));
    layer1_outputs(3903) <= (layer0_outputs(7929)) and not (layer0_outputs(2049));
    layer1_outputs(3904) <= not(layer0_outputs(4717));
    layer1_outputs(3905) <= layer0_outputs(7124);
    layer1_outputs(3906) <= not((layer0_outputs(9768)) or (layer0_outputs(1542)));
    layer1_outputs(3907) <= not(layer0_outputs(2402));
    layer1_outputs(3908) <= '0';
    layer1_outputs(3909) <= not(layer0_outputs(868)) or (layer0_outputs(6428));
    layer1_outputs(3910) <= not(layer0_outputs(8633));
    layer1_outputs(3911) <= (layer0_outputs(1859)) and (layer0_outputs(5919));
    layer1_outputs(3912) <= (layer0_outputs(8334)) or (layer0_outputs(674));
    layer1_outputs(3913) <= not(layer0_outputs(5120));
    layer1_outputs(3914) <= (layer0_outputs(2795)) and not (layer0_outputs(10219));
    layer1_outputs(3915) <= not((layer0_outputs(1957)) or (layer0_outputs(4498)));
    layer1_outputs(3916) <= layer0_outputs(4696);
    layer1_outputs(3917) <= layer0_outputs(8997);
    layer1_outputs(3918) <= (layer0_outputs(2655)) and not (layer0_outputs(699));
    layer1_outputs(3919) <= (layer0_outputs(9284)) and not (layer0_outputs(7236));
    layer1_outputs(3920) <= layer0_outputs(9464);
    layer1_outputs(3921) <= not(layer0_outputs(8863));
    layer1_outputs(3922) <= not(layer0_outputs(2047));
    layer1_outputs(3923) <= not(layer0_outputs(7089)) or (layer0_outputs(8206));
    layer1_outputs(3924) <= not((layer0_outputs(6525)) and (layer0_outputs(7789)));
    layer1_outputs(3925) <= (layer0_outputs(118)) and (layer0_outputs(7111));
    layer1_outputs(3926) <= '0';
    layer1_outputs(3927) <= not(layer0_outputs(9189)) or (layer0_outputs(7732));
    layer1_outputs(3928) <= not(layer0_outputs(8942)) or (layer0_outputs(259));
    layer1_outputs(3929) <= (layer0_outputs(1641)) or (layer0_outputs(4328));
    layer1_outputs(3930) <= not((layer0_outputs(7182)) or (layer0_outputs(9012)));
    layer1_outputs(3931) <= '0';
    layer1_outputs(3932) <= (layer0_outputs(4920)) or (layer0_outputs(9551));
    layer1_outputs(3933) <= not((layer0_outputs(2496)) and (layer0_outputs(6484)));
    layer1_outputs(3934) <= not((layer0_outputs(7249)) and (layer0_outputs(2474)));
    layer1_outputs(3935) <= '0';
    layer1_outputs(3936) <= not(layer0_outputs(4765));
    layer1_outputs(3937) <= not((layer0_outputs(4300)) or (layer0_outputs(5458)));
    layer1_outputs(3938) <= not((layer0_outputs(7235)) or (layer0_outputs(4050)));
    layer1_outputs(3939) <= (layer0_outputs(4248)) and not (layer0_outputs(10025));
    layer1_outputs(3940) <= not(layer0_outputs(1353));
    layer1_outputs(3941) <= not((layer0_outputs(314)) and (layer0_outputs(9595)));
    layer1_outputs(3942) <= '0';
    layer1_outputs(3943) <= not((layer0_outputs(6816)) or (layer0_outputs(0)));
    layer1_outputs(3944) <= layer0_outputs(1114);
    layer1_outputs(3945) <= (layer0_outputs(3676)) and (layer0_outputs(2914));
    layer1_outputs(3946) <= (layer0_outputs(5559)) or (layer0_outputs(2422));
    layer1_outputs(3947) <= not(layer0_outputs(2339)) or (layer0_outputs(3002));
    layer1_outputs(3948) <= not(layer0_outputs(7599));
    layer1_outputs(3949) <= not(layer0_outputs(4615)) or (layer0_outputs(9086));
    layer1_outputs(3950) <= (layer0_outputs(286)) or (layer0_outputs(1994));
    layer1_outputs(3951) <= '0';
    layer1_outputs(3952) <= layer0_outputs(6500);
    layer1_outputs(3953) <= not((layer0_outputs(3066)) or (layer0_outputs(5892)));
    layer1_outputs(3954) <= not(layer0_outputs(10214));
    layer1_outputs(3955) <= not(layer0_outputs(6482));
    layer1_outputs(3956) <= '1';
    layer1_outputs(3957) <= (layer0_outputs(5226)) and not (layer0_outputs(5190));
    layer1_outputs(3958) <= not((layer0_outputs(9425)) xor (layer0_outputs(972)));
    layer1_outputs(3959) <= '1';
    layer1_outputs(3960) <= (layer0_outputs(4899)) or (layer0_outputs(1515));
    layer1_outputs(3961) <= (layer0_outputs(6860)) and not (layer0_outputs(7730));
    layer1_outputs(3962) <= not(layer0_outputs(7594));
    layer1_outputs(3963) <= (layer0_outputs(6019)) and (layer0_outputs(3417));
    layer1_outputs(3964) <= not(layer0_outputs(9513)) or (layer0_outputs(1692));
    layer1_outputs(3965) <= (layer0_outputs(2943)) and not (layer0_outputs(7125));
    layer1_outputs(3966) <= not((layer0_outputs(6646)) or (layer0_outputs(1)));
    layer1_outputs(3967) <= layer0_outputs(8839);
    layer1_outputs(3968) <= layer0_outputs(6504);
    layer1_outputs(3969) <= (layer0_outputs(6404)) xor (layer0_outputs(1642));
    layer1_outputs(3970) <= layer0_outputs(6193);
    layer1_outputs(3971) <= (layer0_outputs(5165)) or (layer0_outputs(8826));
    layer1_outputs(3972) <= layer0_outputs(4856);
    layer1_outputs(3973) <= not(layer0_outputs(1488));
    layer1_outputs(3974) <= not((layer0_outputs(3704)) and (layer0_outputs(2816)));
    layer1_outputs(3975) <= not(layer0_outputs(6362)) or (layer0_outputs(37));
    layer1_outputs(3976) <= not(layer0_outputs(3929)) or (layer0_outputs(3256));
    layer1_outputs(3977) <= not((layer0_outputs(7920)) or (layer0_outputs(61)));
    layer1_outputs(3978) <= layer0_outputs(5502);
    layer1_outputs(3979) <= layer0_outputs(4010);
    layer1_outputs(3980) <= '1';
    layer1_outputs(3981) <= '1';
    layer1_outputs(3982) <= layer0_outputs(1902);
    layer1_outputs(3983) <= '0';
    layer1_outputs(3984) <= not(layer0_outputs(4525));
    layer1_outputs(3985) <= '0';
    layer1_outputs(3986) <= (layer0_outputs(2007)) and not (layer0_outputs(10109));
    layer1_outputs(3987) <= (layer0_outputs(3903)) xor (layer0_outputs(3236));
    layer1_outputs(3988) <= not((layer0_outputs(4795)) or (layer0_outputs(6631)));
    layer1_outputs(3989) <= (layer0_outputs(744)) and not (layer0_outputs(9571));
    layer1_outputs(3990) <= not((layer0_outputs(274)) and (layer0_outputs(9809)));
    layer1_outputs(3991) <= '1';
    layer1_outputs(3992) <= (layer0_outputs(8803)) and not (layer0_outputs(3314));
    layer1_outputs(3993) <= not((layer0_outputs(10179)) or (layer0_outputs(4005)));
    layer1_outputs(3994) <= layer0_outputs(796);
    layer1_outputs(3995) <= not(layer0_outputs(7700));
    layer1_outputs(3996) <= not(layer0_outputs(1293)) or (layer0_outputs(6329));
    layer1_outputs(3997) <= not(layer0_outputs(2074)) or (layer0_outputs(7862));
    layer1_outputs(3998) <= layer0_outputs(9296);
    layer1_outputs(3999) <= not(layer0_outputs(7412));
    layer1_outputs(4000) <= not(layer0_outputs(8916));
    layer1_outputs(4001) <= not((layer0_outputs(2581)) and (layer0_outputs(2495)));
    layer1_outputs(4002) <= layer0_outputs(4898);
    layer1_outputs(4003) <= '1';
    layer1_outputs(4004) <= '0';
    layer1_outputs(4005) <= (layer0_outputs(4247)) and not (layer0_outputs(2759));
    layer1_outputs(4006) <= layer0_outputs(6156);
    layer1_outputs(4007) <= (layer0_outputs(6074)) and (layer0_outputs(3194));
    layer1_outputs(4008) <= not((layer0_outputs(5040)) or (layer0_outputs(6710)));
    layer1_outputs(4009) <= (layer0_outputs(924)) or (layer0_outputs(10116));
    layer1_outputs(4010) <= not((layer0_outputs(8650)) and (layer0_outputs(3979)));
    layer1_outputs(4011) <= not((layer0_outputs(3779)) or (layer0_outputs(2407)));
    layer1_outputs(4012) <= (layer0_outputs(2245)) and not (layer0_outputs(8406));
    layer1_outputs(4013) <= not(layer0_outputs(5374));
    layer1_outputs(4014) <= (layer0_outputs(3694)) and not (layer0_outputs(6988));
    layer1_outputs(4015) <= '1';
    layer1_outputs(4016) <= not((layer0_outputs(8403)) xor (layer0_outputs(8681)));
    layer1_outputs(4017) <= (layer0_outputs(1987)) and not (layer0_outputs(2144));
    layer1_outputs(4018) <= not((layer0_outputs(6197)) xor (layer0_outputs(4637)));
    layer1_outputs(4019) <= not((layer0_outputs(4334)) or (layer0_outputs(4036)));
    layer1_outputs(4020) <= not(layer0_outputs(3087));
    layer1_outputs(4021) <= layer0_outputs(9485);
    layer1_outputs(4022) <= (layer0_outputs(6245)) and not (layer0_outputs(2112));
    layer1_outputs(4023) <= (layer0_outputs(4534)) and not (layer0_outputs(7592));
    layer1_outputs(4024) <= not(layer0_outputs(5508)) or (layer0_outputs(3503));
    layer1_outputs(4025) <= (layer0_outputs(9319)) and not (layer0_outputs(5665));
    layer1_outputs(4026) <= layer0_outputs(3767);
    layer1_outputs(4027) <= not(layer0_outputs(10080));
    layer1_outputs(4028) <= (layer0_outputs(5078)) and not (layer0_outputs(2755));
    layer1_outputs(4029) <= not((layer0_outputs(4439)) xor (layer0_outputs(759)));
    layer1_outputs(4030) <= '1';
    layer1_outputs(4031) <= not((layer0_outputs(5585)) or (layer0_outputs(5308)));
    layer1_outputs(4032) <= not(layer0_outputs(1912)) or (layer0_outputs(2162));
    layer1_outputs(4033) <= not(layer0_outputs(8)) or (layer0_outputs(9970));
    layer1_outputs(4034) <= not(layer0_outputs(8345));
    layer1_outputs(4035) <= layer0_outputs(10128);
    layer1_outputs(4036) <= '0';
    layer1_outputs(4037) <= '0';
    layer1_outputs(4038) <= not(layer0_outputs(4073)) or (layer0_outputs(7138));
    layer1_outputs(4039) <= not(layer0_outputs(778)) or (layer0_outputs(816));
    layer1_outputs(4040) <= not((layer0_outputs(1394)) and (layer0_outputs(2227)));
    layer1_outputs(4041) <= layer0_outputs(2934);
    layer1_outputs(4042) <= not(layer0_outputs(9479)) or (layer0_outputs(269));
    layer1_outputs(4043) <= layer0_outputs(9045);
    layer1_outputs(4044) <= layer0_outputs(9142);
    layer1_outputs(4045) <= not((layer0_outputs(7761)) xor (layer0_outputs(3295)));
    layer1_outputs(4046) <= not((layer0_outputs(1122)) or (layer0_outputs(1614)));
    layer1_outputs(4047) <= not(layer0_outputs(7030));
    layer1_outputs(4048) <= (layer0_outputs(9918)) and not (layer0_outputs(4691));
    layer1_outputs(4049) <= (layer0_outputs(7322)) and (layer0_outputs(7789));
    layer1_outputs(4050) <= '0';
    layer1_outputs(4051) <= (layer0_outputs(6352)) and not (layer0_outputs(8249));
    layer1_outputs(4052) <= layer0_outputs(7819);
    layer1_outputs(4053) <= '0';
    layer1_outputs(4054) <= layer0_outputs(5610);
    layer1_outputs(4055) <= not(layer0_outputs(1335));
    layer1_outputs(4056) <= not(layer0_outputs(7639));
    layer1_outputs(4057) <= not(layer0_outputs(6032));
    layer1_outputs(4058) <= not((layer0_outputs(9294)) or (layer0_outputs(9302)));
    layer1_outputs(4059) <= not(layer0_outputs(9747));
    layer1_outputs(4060) <= (layer0_outputs(2610)) or (layer0_outputs(8127));
    layer1_outputs(4061) <= (layer0_outputs(9385)) and not (layer0_outputs(5225));
    layer1_outputs(4062) <= '0';
    layer1_outputs(4063) <= (layer0_outputs(8013)) and (layer0_outputs(8197));
    layer1_outputs(4064) <= not((layer0_outputs(8227)) and (layer0_outputs(1762)));
    layer1_outputs(4065) <= (layer0_outputs(3646)) or (layer0_outputs(9106));
    layer1_outputs(4066) <= not((layer0_outputs(9306)) or (layer0_outputs(5483)));
    layer1_outputs(4067) <= layer0_outputs(6585);
    layer1_outputs(4068) <= (layer0_outputs(9945)) xor (layer0_outputs(839));
    layer1_outputs(4069) <= not(layer0_outputs(4645)) or (layer0_outputs(307));
    layer1_outputs(4070) <= layer0_outputs(1051);
    layer1_outputs(4071) <= layer0_outputs(4967);
    layer1_outputs(4072) <= layer0_outputs(418);
    layer1_outputs(4073) <= (layer0_outputs(2210)) and (layer0_outputs(3429));
    layer1_outputs(4074) <= (layer0_outputs(6290)) or (layer0_outputs(1225));
    layer1_outputs(4075) <= (layer0_outputs(1385)) and not (layer0_outputs(5027));
    layer1_outputs(4076) <= not(layer0_outputs(6677)) or (layer0_outputs(6560));
    layer1_outputs(4077) <= (layer0_outputs(8902)) or (layer0_outputs(3479));
    layer1_outputs(4078) <= not(layer0_outputs(6290));
    layer1_outputs(4079) <= layer0_outputs(8250);
    layer1_outputs(4080) <= '1';
    layer1_outputs(4081) <= (layer0_outputs(2978)) and not (layer0_outputs(1534));
    layer1_outputs(4082) <= (layer0_outputs(3583)) and not (layer0_outputs(2608));
    layer1_outputs(4083) <= layer0_outputs(3920);
    layer1_outputs(4084) <= not((layer0_outputs(4242)) and (layer0_outputs(9747)));
    layer1_outputs(4085) <= not(layer0_outputs(3681)) or (layer0_outputs(7737));
    layer1_outputs(4086) <= (layer0_outputs(3904)) and not (layer0_outputs(908));
    layer1_outputs(4087) <= (layer0_outputs(7311)) and (layer0_outputs(7169));
    layer1_outputs(4088) <= not(layer0_outputs(8037)) or (layer0_outputs(7474));
    layer1_outputs(4089) <= layer0_outputs(7245);
    layer1_outputs(4090) <= layer0_outputs(4719);
    layer1_outputs(4091) <= '0';
    layer1_outputs(4092) <= (layer0_outputs(2983)) and (layer0_outputs(5525));
    layer1_outputs(4093) <= (layer0_outputs(7601)) and not (layer0_outputs(6721));
    layer1_outputs(4094) <= not(layer0_outputs(8017));
    layer1_outputs(4095) <= not((layer0_outputs(1447)) xor (layer0_outputs(425)));
    layer1_outputs(4096) <= not((layer0_outputs(9704)) xor (layer0_outputs(6678)));
    layer1_outputs(4097) <= not(layer0_outputs(5220));
    layer1_outputs(4098) <= not((layer0_outputs(1818)) and (layer0_outputs(3727)));
    layer1_outputs(4099) <= not(layer0_outputs(3119));
    layer1_outputs(4100) <= '1';
    layer1_outputs(4101) <= not(layer0_outputs(8812));
    layer1_outputs(4102) <= not(layer0_outputs(7017));
    layer1_outputs(4103) <= layer0_outputs(5526);
    layer1_outputs(4104) <= not(layer0_outputs(3020)) or (layer0_outputs(4604));
    layer1_outputs(4105) <= not(layer0_outputs(2907)) or (layer0_outputs(6663));
    layer1_outputs(4106) <= (layer0_outputs(3271)) and not (layer0_outputs(1428));
    layer1_outputs(4107) <= not((layer0_outputs(371)) or (layer0_outputs(4761)));
    layer1_outputs(4108) <= not(layer0_outputs(6557)) or (layer0_outputs(7788));
    layer1_outputs(4109) <= not(layer0_outputs(5893));
    layer1_outputs(4110) <= not((layer0_outputs(5983)) and (layer0_outputs(10165)));
    layer1_outputs(4111) <= layer0_outputs(8081);
    layer1_outputs(4112) <= '0';
    layer1_outputs(4113) <= layer0_outputs(1645);
    layer1_outputs(4114) <= '1';
    layer1_outputs(4115) <= not(layer0_outputs(9882)) or (layer0_outputs(508));
    layer1_outputs(4116) <= '0';
    layer1_outputs(4117) <= not(layer0_outputs(6455));
    layer1_outputs(4118) <= not(layer0_outputs(4868));
    layer1_outputs(4119) <= '1';
    layer1_outputs(4120) <= (layer0_outputs(502)) and not (layer0_outputs(3174));
    layer1_outputs(4121) <= not((layer0_outputs(4063)) and (layer0_outputs(4099)));
    layer1_outputs(4122) <= not((layer0_outputs(3984)) or (layer0_outputs(7341)));
    layer1_outputs(4123) <= not(layer0_outputs(6858));
    layer1_outputs(4124) <= layer0_outputs(4151);
    layer1_outputs(4125) <= not(layer0_outputs(1684));
    layer1_outputs(4126) <= not(layer0_outputs(3132)) or (layer0_outputs(8815));
    layer1_outputs(4127) <= '0';
    layer1_outputs(4128) <= (layer0_outputs(8925)) and (layer0_outputs(7948));
    layer1_outputs(4129) <= not(layer0_outputs(4530)) or (layer0_outputs(564));
    layer1_outputs(4130) <= not(layer0_outputs(8109));
    layer1_outputs(4131) <= not(layer0_outputs(8212)) or (layer0_outputs(5600));
    layer1_outputs(4132) <= not((layer0_outputs(3750)) and (layer0_outputs(4603)));
    layer1_outputs(4133) <= layer0_outputs(6760);
    layer1_outputs(4134) <= (layer0_outputs(2693)) and not (layer0_outputs(9767));
    layer1_outputs(4135) <= (layer0_outputs(8621)) and not (layer0_outputs(4194));
    layer1_outputs(4136) <= not((layer0_outputs(2107)) xor (layer0_outputs(4830)));
    layer1_outputs(4137) <= (layer0_outputs(4417)) and not (layer0_outputs(705));
    layer1_outputs(4138) <= not((layer0_outputs(4138)) and (layer0_outputs(9031)));
    layer1_outputs(4139) <= not(layer0_outputs(6842)) or (layer0_outputs(6836));
    layer1_outputs(4140) <= not(layer0_outputs(9275)) or (layer0_outputs(6596));
    layer1_outputs(4141) <= not(layer0_outputs(5231)) or (layer0_outputs(2587));
    layer1_outputs(4142) <= layer0_outputs(2555);
    layer1_outputs(4143) <= layer0_outputs(7568);
    layer1_outputs(4144) <= not(layer0_outputs(6478)) or (layer0_outputs(1625));
    layer1_outputs(4145) <= '0';
    layer1_outputs(4146) <= '1';
    layer1_outputs(4147) <= not((layer0_outputs(1117)) or (layer0_outputs(6295)));
    layer1_outputs(4148) <= (layer0_outputs(298)) and (layer0_outputs(2840));
    layer1_outputs(4149) <= not(layer0_outputs(6082));
    layer1_outputs(4150) <= not((layer0_outputs(4258)) or (layer0_outputs(8458)));
    layer1_outputs(4151) <= not(layer0_outputs(10102)) or (layer0_outputs(7929));
    layer1_outputs(4152) <= not((layer0_outputs(3756)) and (layer0_outputs(4707)));
    layer1_outputs(4153) <= not(layer0_outputs(5672));
    layer1_outputs(4154) <= (layer0_outputs(4837)) and not (layer0_outputs(8208));
    layer1_outputs(4155) <= (layer0_outputs(9837)) or (layer0_outputs(448));
    layer1_outputs(4156) <= '0';
    layer1_outputs(4157) <= layer0_outputs(695);
    layer1_outputs(4158) <= '1';
    layer1_outputs(4159) <= '1';
    layer1_outputs(4160) <= layer0_outputs(9760);
    layer1_outputs(4161) <= not(layer0_outputs(2713)) or (layer0_outputs(637));
    layer1_outputs(4162) <= layer0_outputs(4863);
    layer1_outputs(4163) <= (layer0_outputs(461)) and not (layer0_outputs(9978));
    layer1_outputs(4164) <= (layer0_outputs(8305)) and (layer0_outputs(869));
    layer1_outputs(4165) <= layer0_outputs(6152);
    layer1_outputs(4166) <= not(layer0_outputs(4472));
    layer1_outputs(4167) <= (layer0_outputs(9017)) or (layer0_outputs(243));
    layer1_outputs(4168) <= not(layer0_outputs(2594));
    layer1_outputs(4169) <= (layer0_outputs(3776)) xor (layer0_outputs(4954));
    layer1_outputs(4170) <= not(layer0_outputs(10105));
    layer1_outputs(4171) <= not(layer0_outputs(9423)) or (layer0_outputs(2618));
    layer1_outputs(4172) <= not((layer0_outputs(5466)) or (layer0_outputs(175)));
    layer1_outputs(4173) <= (layer0_outputs(9900)) xor (layer0_outputs(7559));
    layer1_outputs(4174) <= layer0_outputs(3396);
    layer1_outputs(4175) <= not((layer0_outputs(3922)) or (layer0_outputs(1510)));
    layer1_outputs(4176) <= layer0_outputs(1465);
    layer1_outputs(4177) <= not((layer0_outputs(8474)) or (layer0_outputs(6673)));
    layer1_outputs(4178) <= not(layer0_outputs(6422)) or (layer0_outputs(4451));
    layer1_outputs(4179) <= layer0_outputs(3238);
    layer1_outputs(4180) <= not(layer0_outputs(4121));
    layer1_outputs(4181) <= not(layer0_outputs(7806));
    layer1_outputs(4182) <= layer0_outputs(2116);
    layer1_outputs(4183) <= layer0_outputs(4993);
    layer1_outputs(4184) <= (layer0_outputs(6339)) and not (layer0_outputs(7129));
    layer1_outputs(4185) <= (layer0_outputs(4851)) and not (layer0_outputs(3788));
    layer1_outputs(4186) <= (layer0_outputs(8536)) or (layer0_outputs(8643));
    layer1_outputs(4187) <= (layer0_outputs(2743)) and (layer0_outputs(2245));
    layer1_outputs(4188) <= not((layer0_outputs(409)) and (layer0_outputs(10212)));
    layer1_outputs(4189) <= not((layer0_outputs(8605)) xor (layer0_outputs(6216)));
    layer1_outputs(4190) <= not(layer0_outputs(9972)) or (layer0_outputs(7906));
    layer1_outputs(4191) <= '1';
    layer1_outputs(4192) <= (layer0_outputs(8529)) and (layer0_outputs(5306));
    layer1_outputs(4193) <= not((layer0_outputs(8915)) and (layer0_outputs(1269)));
    layer1_outputs(4194) <= layer0_outputs(65);
    layer1_outputs(4195) <= (layer0_outputs(4122)) and not (layer0_outputs(7672));
    layer1_outputs(4196) <= '1';
    layer1_outputs(4197) <= '1';
    layer1_outputs(4198) <= layer0_outputs(2040);
    layer1_outputs(4199) <= not(layer0_outputs(375));
    layer1_outputs(4200) <= layer0_outputs(1002);
    layer1_outputs(4201) <= (layer0_outputs(684)) and (layer0_outputs(9967));
    layer1_outputs(4202) <= (layer0_outputs(6073)) xor (layer0_outputs(6076));
    layer1_outputs(4203) <= not(layer0_outputs(9193));
    layer1_outputs(4204) <= '1';
    layer1_outputs(4205) <= '1';
    layer1_outputs(4206) <= (layer0_outputs(7782)) or (layer0_outputs(10089));
    layer1_outputs(4207) <= '0';
    layer1_outputs(4208) <= (layer0_outputs(5336)) or (layer0_outputs(4583));
    layer1_outputs(4209) <= not((layer0_outputs(914)) or (layer0_outputs(5020)));
    layer1_outputs(4210) <= (layer0_outputs(536)) and not (layer0_outputs(9708));
    layer1_outputs(4211) <= not((layer0_outputs(5565)) or (layer0_outputs(6342)));
    layer1_outputs(4212) <= not(layer0_outputs(6300)) or (layer0_outputs(3716));
    layer1_outputs(4213) <= not(layer0_outputs(9419));
    layer1_outputs(4214) <= not(layer0_outputs(9626)) or (layer0_outputs(1379));
    layer1_outputs(4215) <= layer0_outputs(8438);
    layer1_outputs(4216) <= (layer0_outputs(2870)) and (layer0_outputs(4093));
    layer1_outputs(4217) <= (layer0_outputs(9386)) and (layer0_outputs(3170));
    layer1_outputs(4218) <= not(layer0_outputs(9450)) or (layer0_outputs(5072));
    layer1_outputs(4219) <= not((layer0_outputs(4651)) or (layer0_outputs(2388)));
    layer1_outputs(4220) <= layer0_outputs(4776);
    layer1_outputs(4221) <= (layer0_outputs(3178)) and (layer0_outputs(9052));
    layer1_outputs(4222) <= not(layer0_outputs(901));
    layer1_outputs(4223) <= not(layer0_outputs(5681)) or (layer0_outputs(3736));
    layer1_outputs(4224) <= (layer0_outputs(7828)) and not (layer0_outputs(8741));
    layer1_outputs(4225) <= (layer0_outputs(6913)) and not (layer0_outputs(5571));
    layer1_outputs(4226) <= '1';
    layer1_outputs(4227) <= (layer0_outputs(1576)) and (layer0_outputs(4950));
    layer1_outputs(4228) <= not(layer0_outputs(8814)) or (layer0_outputs(1712));
    layer1_outputs(4229) <= not(layer0_outputs(10235)) or (layer0_outputs(9198));
    layer1_outputs(4230) <= layer0_outputs(7556);
    layer1_outputs(4231) <= layer0_outputs(7376);
    layer1_outputs(4232) <= (layer0_outputs(6041)) and (layer0_outputs(2922));
    layer1_outputs(4233) <= not(layer0_outputs(9187));
    layer1_outputs(4234) <= (layer0_outputs(1498)) or (layer0_outputs(2926));
    layer1_outputs(4235) <= layer0_outputs(8684);
    layer1_outputs(4236) <= (layer0_outputs(231)) and not (layer0_outputs(8709));
    layer1_outputs(4237) <= not((layer0_outputs(8934)) and (layer0_outputs(8235)));
    layer1_outputs(4238) <= not(layer0_outputs(982)) or (layer0_outputs(1574));
    layer1_outputs(4239) <= layer0_outputs(3225);
    layer1_outputs(4240) <= (layer0_outputs(8163)) and not (layer0_outputs(795));
    layer1_outputs(4241) <= not(layer0_outputs(8907));
    layer1_outputs(4242) <= (layer0_outputs(9215)) xor (layer0_outputs(8967));
    layer1_outputs(4243) <= layer0_outputs(9489);
    layer1_outputs(4244) <= not(layer0_outputs(1352));
    layer1_outputs(4245) <= not(layer0_outputs(9003));
    layer1_outputs(4246) <= not(layer0_outputs(10203));
    layer1_outputs(4247) <= layer0_outputs(10206);
    layer1_outputs(4248) <= layer0_outputs(4460);
    layer1_outputs(4249) <= (layer0_outputs(4981)) and not (layer0_outputs(9555));
    layer1_outputs(4250) <= not(layer0_outputs(9709)) or (layer0_outputs(9995));
    layer1_outputs(4251) <= '1';
    layer1_outputs(4252) <= not(layer0_outputs(9474)) or (layer0_outputs(1543));
    layer1_outputs(4253) <= not(layer0_outputs(2085));
    layer1_outputs(4254) <= not(layer0_outputs(3820));
    layer1_outputs(4255) <= (layer0_outputs(8371)) and not (layer0_outputs(8495));
    layer1_outputs(4256) <= '0';
    layer1_outputs(4257) <= '0';
    layer1_outputs(4258) <= not(layer0_outputs(1827));
    layer1_outputs(4259) <= layer0_outputs(6493);
    layer1_outputs(4260) <= (layer0_outputs(2502)) and (layer0_outputs(8416));
    layer1_outputs(4261) <= not(layer0_outputs(3860));
    layer1_outputs(4262) <= not(layer0_outputs(7344));
    layer1_outputs(4263) <= not(layer0_outputs(3047)) or (layer0_outputs(8540));
    layer1_outputs(4264) <= (layer0_outputs(8402)) and not (layer0_outputs(2937));
    layer1_outputs(4265) <= layer0_outputs(6220);
    layer1_outputs(4266) <= not(layer0_outputs(8258));
    layer1_outputs(4267) <= not(layer0_outputs(8383)) or (layer0_outputs(4824));
    layer1_outputs(4268) <= not(layer0_outputs(8028)) or (layer0_outputs(9401));
    layer1_outputs(4269) <= not(layer0_outputs(701)) or (layer0_outputs(8292));
    layer1_outputs(4270) <= (layer0_outputs(7069)) and (layer0_outputs(5467));
    layer1_outputs(4271) <= (layer0_outputs(7424)) and not (layer0_outputs(6703));
    layer1_outputs(4272) <= layer0_outputs(4690);
    layer1_outputs(4273) <= (layer0_outputs(6894)) and (layer0_outputs(7932));
    layer1_outputs(4274) <= layer0_outputs(2951);
    layer1_outputs(4275) <= not((layer0_outputs(1681)) and (layer0_outputs(3884)));
    layer1_outputs(4276) <= (layer0_outputs(448)) or (layer0_outputs(9864));
    layer1_outputs(4277) <= (layer0_outputs(694)) and (layer0_outputs(919));
    layer1_outputs(4278) <= layer0_outputs(5987);
    layer1_outputs(4279) <= (layer0_outputs(5570)) or (layer0_outputs(1138));
    layer1_outputs(4280) <= (layer0_outputs(1633)) and not (layer0_outputs(9399));
    layer1_outputs(4281) <= (layer0_outputs(2196)) and not (layer0_outputs(603));
    layer1_outputs(4282) <= layer0_outputs(8283);
    layer1_outputs(4283) <= (layer0_outputs(3716)) and (layer0_outputs(5605));
    layer1_outputs(4284) <= (layer0_outputs(4190)) and not (layer0_outputs(2634));
    layer1_outputs(4285) <= (layer0_outputs(7675)) and not (layer0_outputs(25));
    layer1_outputs(4286) <= not((layer0_outputs(2826)) xor (layer0_outputs(6251)));
    layer1_outputs(4287) <= not(layer0_outputs(9178));
    layer1_outputs(4288) <= layer0_outputs(7534);
    layer1_outputs(4289) <= (layer0_outputs(942)) and (layer0_outputs(9270));
    layer1_outputs(4290) <= '0';
    layer1_outputs(4291) <= '1';
    layer1_outputs(4292) <= not(layer0_outputs(4525));
    layer1_outputs(4293) <= not((layer0_outputs(7667)) xor (layer0_outputs(8733)));
    layer1_outputs(4294) <= not(layer0_outputs(5624));
    layer1_outputs(4295) <= (layer0_outputs(5397)) and not (layer0_outputs(3962));
    layer1_outputs(4296) <= not(layer0_outputs(580)) or (layer0_outputs(9904));
    layer1_outputs(4297) <= not((layer0_outputs(10133)) or (layer0_outputs(6363)));
    layer1_outputs(4298) <= (layer0_outputs(3080)) xor (layer0_outputs(3438));
    layer1_outputs(4299) <= not((layer0_outputs(4284)) or (layer0_outputs(1799)));
    layer1_outputs(4300) <= not((layer0_outputs(4173)) xor (layer0_outputs(6889)));
    layer1_outputs(4301) <= (layer0_outputs(1326)) or (layer0_outputs(4714));
    layer1_outputs(4302) <= layer0_outputs(4115);
    layer1_outputs(4303) <= not(layer0_outputs(4197));
    layer1_outputs(4304) <= (layer0_outputs(7870)) or (layer0_outputs(7240));
    layer1_outputs(4305) <= not(layer0_outputs(6227));
    layer1_outputs(4306) <= not(layer0_outputs(7898));
    layer1_outputs(4307) <= not(layer0_outputs(5166));
    layer1_outputs(4308) <= not((layer0_outputs(9956)) xor (layer0_outputs(9622)));
    layer1_outputs(4309) <= not(layer0_outputs(742));
    layer1_outputs(4310) <= (layer0_outputs(6019)) or (layer0_outputs(3077));
    layer1_outputs(4311) <= not(layer0_outputs(7865)) or (layer0_outputs(7777));
    layer1_outputs(4312) <= (layer0_outputs(7529)) and (layer0_outputs(4834));
    layer1_outputs(4313) <= not((layer0_outputs(941)) and (layer0_outputs(4621)));
    layer1_outputs(4314) <= not((layer0_outputs(1336)) or (layer0_outputs(770)));
    layer1_outputs(4315) <= (layer0_outputs(10033)) and not (layer0_outputs(1348));
    layer1_outputs(4316) <= not(layer0_outputs(4156)) or (layer0_outputs(9645));
    layer1_outputs(4317) <= layer0_outputs(5537);
    layer1_outputs(4318) <= not(layer0_outputs(5856)) or (layer0_outputs(7725));
    layer1_outputs(4319) <= (layer0_outputs(4119)) or (layer0_outputs(7207));
    layer1_outputs(4320) <= layer0_outputs(5168);
    layer1_outputs(4321) <= (layer0_outputs(5256)) or (layer0_outputs(4609));
    layer1_outputs(4322) <= (layer0_outputs(6105)) and not (layer0_outputs(1263));
    layer1_outputs(4323) <= (layer0_outputs(3395)) and not (layer0_outputs(7905));
    layer1_outputs(4324) <= '0';
    layer1_outputs(4325) <= not(layer0_outputs(944));
    layer1_outputs(4326) <= (layer0_outputs(900)) or (layer0_outputs(1935));
    layer1_outputs(4327) <= layer0_outputs(6658);
    layer1_outputs(4328) <= not(layer0_outputs(9449)) or (layer0_outputs(7071));
    layer1_outputs(4329) <= (layer0_outputs(8972)) and not (layer0_outputs(458));
    layer1_outputs(4330) <= not(layer0_outputs(1188));
    layer1_outputs(4331) <= not(layer0_outputs(5874)) or (layer0_outputs(3516));
    layer1_outputs(4332) <= layer0_outputs(5566);
    layer1_outputs(4333) <= (layer0_outputs(1867)) and (layer0_outputs(2156));
    layer1_outputs(4334) <= not((layer0_outputs(2966)) or (layer0_outputs(6010)));
    layer1_outputs(4335) <= not(layer0_outputs(7812));
    layer1_outputs(4336) <= layer0_outputs(4573);
    layer1_outputs(4337) <= layer0_outputs(6528);
    layer1_outputs(4338) <= not(layer0_outputs(4244)) or (layer0_outputs(4750));
    layer1_outputs(4339) <= layer0_outputs(7951);
    layer1_outputs(4340) <= not(layer0_outputs(1331)) or (layer0_outputs(5667));
    layer1_outputs(4341) <= not((layer0_outputs(4686)) or (layer0_outputs(5188)));
    layer1_outputs(4342) <= not((layer0_outputs(368)) and (layer0_outputs(8833)));
    layer1_outputs(4343) <= (layer0_outputs(4147)) xor (layer0_outputs(5332));
    layer1_outputs(4344) <= '0';
    layer1_outputs(4345) <= layer0_outputs(4119);
    layer1_outputs(4346) <= layer0_outputs(531);
    layer1_outputs(4347) <= layer0_outputs(8367);
    layer1_outputs(4348) <= not(layer0_outputs(2857));
    layer1_outputs(4349) <= not(layer0_outputs(4207));
    layer1_outputs(4350) <= (layer0_outputs(3805)) or (layer0_outputs(10105));
    layer1_outputs(4351) <= not(layer0_outputs(899));
    layer1_outputs(4352) <= layer0_outputs(1492);
    layer1_outputs(4353) <= not(layer0_outputs(4892));
    layer1_outputs(4354) <= layer0_outputs(6348);
    layer1_outputs(4355) <= not(layer0_outputs(996)) or (layer0_outputs(8220));
    layer1_outputs(4356) <= (layer0_outputs(2039)) and not (layer0_outputs(9989));
    layer1_outputs(4357) <= layer0_outputs(386);
    layer1_outputs(4358) <= (layer0_outputs(3315)) or (layer0_outputs(1637));
    layer1_outputs(4359) <= layer0_outputs(5314);
    layer1_outputs(4360) <= (layer0_outputs(9208)) and (layer0_outputs(4506));
    layer1_outputs(4361) <= not(layer0_outputs(4517));
    layer1_outputs(4362) <= not(layer0_outputs(3147)) or (layer0_outputs(7512));
    layer1_outputs(4363) <= (layer0_outputs(2474)) and (layer0_outputs(5799));
    layer1_outputs(4364) <= (layer0_outputs(9642)) and not (layer0_outputs(8873));
    layer1_outputs(4365) <= layer0_outputs(9205);
    layer1_outputs(4366) <= (layer0_outputs(6083)) and not (layer0_outputs(5879));
    layer1_outputs(4367) <= not(layer0_outputs(5170));
    layer1_outputs(4368) <= layer0_outputs(3732);
    layer1_outputs(4369) <= not(layer0_outputs(3695));
    layer1_outputs(4370) <= (layer0_outputs(1372)) and not (layer0_outputs(7888));
    layer1_outputs(4371) <= layer0_outputs(7614);
    layer1_outputs(4372) <= not((layer0_outputs(6942)) or (layer0_outputs(5984)));
    layer1_outputs(4373) <= not((layer0_outputs(7082)) or (layer0_outputs(115)));
    layer1_outputs(4374) <= not((layer0_outputs(1205)) and (layer0_outputs(5843)));
    layer1_outputs(4375) <= not((layer0_outputs(3194)) xor (layer0_outputs(2365)));
    layer1_outputs(4376) <= not(layer0_outputs(3097));
    layer1_outputs(4377) <= (layer0_outputs(9622)) or (layer0_outputs(1430));
    layer1_outputs(4378) <= not((layer0_outputs(787)) xor (layer0_outputs(2860)));
    layer1_outputs(4379) <= not((layer0_outputs(5012)) and (layer0_outputs(962)));
    layer1_outputs(4380) <= layer0_outputs(1112);
    layer1_outputs(4381) <= (layer0_outputs(3989)) and not (layer0_outputs(1653));
    layer1_outputs(4382) <= (layer0_outputs(6748)) or (layer0_outputs(4188));
    layer1_outputs(4383) <= not(layer0_outputs(4323)) or (layer0_outputs(3522));
    layer1_outputs(4384) <= layer0_outputs(1369);
    layer1_outputs(4385) <= (layer0_outputs(1058)) xor (layer0_outputs(8705));
    layer1_outputs(4386) <= not(layer0_outputs(3874)) or (layer0_outputs(3717));
    layer1_outputs(4387) <= layer0_outputs(4790);
    layer1_outputs(4388) <= (layer0_outputs(364)) and not (layer0_outputs(2677));
    layer1_outputs(4389) <= not((layer0_outputs(917)) xor (layer0_outputs(7727)));
    layer1_outputs(4390) <= (layer0_outputs(4006)) and not (layer0_outputs(2804));
    layer1_outputs(4391) <= layer0_outputs(6358);
    layer1_outputs(4392) <= layer0_outputs(8728);
    layer1_outputs(4393) <= (layer0_outputs(5697)) xor (layer0_outputs(6112));
    layer1_outputs(4394) <= layer0_outputs(2760);
    layer1_outputs(4395) <= (layer0_outputs(3218)) and not (layer0_outputs(1034));
    layer1_outputs(4396) <= not((layer0_outputs(7531)) or (layer0_outputs(951)));
    layer1_outputs(4397) <= not((layer0_outputs(1027)) and (layer0_outputs(10181)));
    layer1_outputs(4398) <= not((layer0_outputs(5509)) and (layer0_outputs(4822)));
    layer1_outputs(4399) <= (layer0_outputs(189)) and (layer0_outputs(10062));
    layer1_outputs(4400) <= not((layer0_outputs(7802)) or (layer0_outputs(7604)));
    layer1_outputs(4401) <= (layer0_outputs(3096)) and not (layer0_outputs(260));
    layer1_outputs(4402) <= (layer0_outputs(7160)) and not (layer0_outputs(7671));
    layer1_outputs(4403) <= layer0_outputs(5798);
    layer1_outputs(4404) <= not((layer0_outputs(7448)) or (layer0_outputs(4157)));
    layer1_outputs(4405) <= (layer0_outputs(7547)) or (layer0_outputs(8665));
    layer1_outputs(4406) <= not((layer0_outputs(1221)) and (layer0_outputs(1159)));
    layer1_outputs(4407) <= (layer0_outputs(5909)) and (layer0_outputs(8296));
    layer1_outputs(4408) <= not(layer0_outputs(2022)) or (layer0_outputs(9985));
    layer1_outputs(4409) <= (layer0_outputs(441)) and not (layer0_outputs(521));
    layer1_outputs(4410) <= (layer0_outputs(4981)) and not (layer0_outputs(2350));
    layer1_outputs(4411) <= not(layer0_outputs(4458));
    layer1_outputs(4412) <= not((layer0_outputs(10230)) or (layer0_outputs(4355)));
    layer1_outputs(4413) <= not(layer0_outputs(3346));
    layer1_outputs(4414) <= not(layer0_outputs(4288));
    layer1_outputs(4415) <= not(layer0_outputs(9988)) or (layer0_outputs(9251));
    layer1_outputs(4416) <= layer0_outputs(9562);
    layer1_outputs(4417) <= (layer0_outputs(8892)) xor (layer0_outputs(6366));
    layer1_outputs(4418) <= (layer0_outputs(1784)) xor (layer0_outputs(2801));
    layer1_outputs(4419) <= not(layer0_outputs(1590)) or (layer0_outputs(1151));
    layer1_outputs(4420) <= (layer0_outputs(4284)) or (layer0_outputs(6223));
    layer1_outputs(4421) <= (layer0_outputs(5283)) or (layer0_outputs(2773));
    layer1_outputs(4422) <= (layer0_outputs(9843)) xor (layer0_outputs(10137));
    layer1_outputs(4423) <= (layer0_outputs(2381)) and not (layer0_outputs(5423));
    layer1_outputs(4424) <= (layer0_outputs(8130)) and (layer0_outputs(23));
    layer1_outputs(4425) <= (layer0_outputs(6626)) and (layer0_outputs(2498));
    layer1_outputs(4426) <= not(layer0_outputs(979)) or (layer0_outputs(5399));
    layer1_outputs(4427) <= '1';
    layer1_outputs(4428) <= layer0_outputs(8538);
    layer1_outputs(4429) <= (layer0_outputs(9578)) and not (layer0_outputs(1327));
    layer1_outputs(4430) <= not(layer0_outputs(7465));
    layer1_outputs(4431) <= (layer0_outputs(7588)) and (layer0_outputs(2224));
    layer1_outputs(4432) <= (layer0_outputs(5212)) and not (layer0_outputs(785));
    layer1_outputs(4433) <= layer0_outputs(7550);
    layer1_outputs(4434) <= not(layer0_outputs(3996));
    layer1_outputs(4435) <= (layer0_outputs(8119)) or (layer0_outputs(9358));
    layer1_outputs(4436) <= layer0_outputs(980);
    layer1_outputs(4437) <= (layer0_outputs(6869)) xor (layer0_outputs(9023));
    layer1_outputs(4438) <= not(layer0_outputs(6654));
    layer1_outputs(4439) <= not((layer0_outputs(8412)) xor (layer0_outputs(6706)));
    layer1_outputs(4440) <= not((layer0_outputs(8467)) and (layer0_outputs(5811)));
    layer1_outputs(4441) <= layer0_outputs(7328);
    layer1_outputs(4442) <= not(layer0_outputs(1838)) or (layer0_outputs(439));
    layer1_outputs(4443) <= not((layer0_outputs(1607)) and (layer0_outputs(6373)));
    layer1_outputs(4444) <= '1';
    layer1_outputs(4445) <= layer0_outputs(9888);
    layer1_outputs(4446) <= (layer0_outputs(7132)) and not (layer0_outputs(933));
    layer1_outputs(4447) <= not(layer0_outputs(1451)) or (layer0_outputs(331));
    layer1_outputs(4448) <= (layer0_outputs(3366)) and not (layer0_outputs(1471));
    layer1_outputs(4449) <= not(layer0_outputs(9720));
    layer1_outputs(4450) <= (layer0_outputs(4850)) or (layer0_outputs(2304));
    layer1_outputs(4451) <= not(layer0_outputs(1436));
    layer1_outputs(4452) <= not(layer0_outputs(640)) or (layer0_outputs(6765));
    layer1_outputs(4453) <= not((layer0_outputs(3796)) or (layer0_outputs(5538)));
    layer1_outputs(4454) <= (layer0_outputs(2748)) xor (layer0_outputs(2489));
    layer1_outputs(4455) <= layer0_outputs(62);
    layer1_outputs(4456) <= not(layer0_outputs(4260));
    layer1_outputs(4457) <= (layer0_outputs(7004)) and (layer0_outputs(9931));
    layer1_outputs(4458) <= (layer0_outputs(1966)) and (layer0_outputs(6648));
    layer1_outputs(4459) <= not(layer0_outputs(5819)) or (layer0_outputs(9390));
    layer1_outputs(4460) <= not(layer0_outputs(3324)) or (layer0_outputs(3173));
    layer1_outputs(4461) <= not((layer0_outputs(7495)) and (layer0_outputs(5353)));
    layer1_outputs(4462) <= not((layer0_outputs(3839)) xor (layer0_outputs(8312)));
    layer1_outputs(4463) <= not(layer0_outputs(2846));
    layer1_outputs(4464) <= not((layer0_outputs(9341)) and (layer0_outputs(4554)));
    layer1_outputs(4465) <= layer0_outputs(995);
    layer1_outputs(4466) <= not(layer0_outputs(7339)) or (layer0_outputs(5155));
    layer1_outputs(4467) <= '1';
    layer1_outputs(4468) <= not(layer0_outputs(1052));
    layer1_outputs(4469) <= not(layer0_outputs(5812)) or (layer0_outputs(28));
    layer1_outputs(4470) <= not(layer0_outputs(7155));
    layer1_outputs(4471) <= layer0_outputs(7255);
    layer1_outputs(4472) <= not((layer0_outputs(2846)) and (layer0_outputs(2778)));
    layer1_outputs(4473) <= not(layer0_outputs(5392));
    layer1_outputs(4474) <= not((layer0_outputs(2336)) and (layer0_outputs(567)));
    layer1_outputs(4475) <= not(layer0_outputs(4881));
    layer1_outputs(4476) <= layer0_outputs(6875);
    layer1_outputs(4477) <= (layer0_outputs(10136)) and (layer0_outputs(8046));
    layer1_outputs(4478) <= not((layer0_outputs(56)) or (layer0_outputs(2133)));
    layer1_outputs(4479) <= layer0_outputs(5176);
    layer1_outputs(4480) <= layer0_outputs(1555);
    layer1_outputs(4481) <= (layer0_outputs(10163)) and (layer0_outputs(5768));
    layer1_outputs(4482) <= not(layer0_outputs(9410)) or (layer0_outputs(2099));
    layer1_outputs(4483) <= '1';
    layer1_outputs(4484) <= '1';
    layer1_outputs(4485) <= (layer0_outputs(9194)) or (layer0_outputs(6862));
    layer1_outputs(4486) <= (layer0_outputs(8650)) and not (layer0_outputs(1963));
    layer1_outputs(4487) <= not(layer0_outputs(1526)) or (layer0_outputs(7338));
    layer1_outputs(4488) <= layer0_outputs(7249);
    layer1_outputs(4489) <= (layer0_outputs(6510)) and not (layer0_outputs(3993));
    layer1_outputs(4490) <= (layer0_outputs(4880)) and not (layer0_outputs(7763));
    layer1_outputs(4491) <= not((layer0_outputs(500)) or (layer0_outputs(8940)));
    layer1_outputs(4492) <= (layer0_outputs(2984)) and not (layer0_outputs(925));
    layer1_outputs(4493) <= not(layer0_outputs(2061)) or (layer0_outputs(2983));
    layer1_outputs(4494) <= not(layer0_outputs(6062));
    layer1_outputs(4495) <= '0';
    layer1_outputs(4496) <= not(layer0_outputs(5329));
    layer1_outputs(4497) <= (layer0_outputs(4710)) and not (layer0_outputs(6940));
    layer1_outputs(4498) <= layer0_outputs(4946);
    layer1_outputs(4499) <= (layer0_outputs(4270)) xor (layer0_outputs(8109));
    layer1_outputs(4500) <= '1';
    layer1_outputs(4501) <= not(layer0_outputs(2622)) or (layer0_outputs(9674));
    layer1_outputs(4502) <= '1';
    layer1_outputs(4503) <= not((layer0_outputs(2469)) or (layer0_outputs(1106)));
    layer1_outputs(4504) <= not(layer0_outputs(9803)) or (layer0_outputs(7940));
    layer1_outputs(4505) <= (layer0_outputs(7160)) or (layer0_outputs(7729));
    layer1_outputs(4506) <= not(layer0_outputs(9369));
    layer1_outputs(4507) <= (layer0_outputs(2355)) and not (layer0_outputs(8032));
    layer1_outputs(4508) <= not((layer0_outputs(5378)) or (layer0_outputs(6824)));
    layer1_outputs(4509) <= (layer0_outputs(4393)) and not (layer0_outputs(5139));
    layer1_outputs(4510) <= not(layer0_outputs(5916));
    layer1_outputs(4511) <= layer0_outputs(9834);
    layer1_outputs(4512) <= not(layer0_outputs(9504));
    layer1_outputs(4513) <= not(layer0_outputs(433));
    layer1_outputs(4514) <= (layer0_outputs(9238)) and not (layer0_outputs(9367));
    layer1_outputs(4515) <= layer0_outputs(9103);
    layer1_outputs(4516) <= (layer0_outputs(1810)) and not (layer0_outputs(4970));
    layer1_outputs(4517) <= layer0_outputs(1906);
    layer1_outputs(4518) <= '1';
    layer1_outputs(4519) <= not(layer0_outputs(9971));
    layer1_outputs(4520) <= not(layer0_outputs(8554)) or (layer0_outputs(7913));
    layer1_outputs(4521) <= not(layer0_outputs(3371));
    layer1_outputs(4522) <= (layer0_outputs(7662)) xor (layer0_outputs(7063));
    layer1_outputs(4523) <= not((layer0_outputs(2206)) xor (layer0_outputs(5787)));
    layer1_outputs(4524) <= '1';
    layer1_outputs(4525) <= not(layer0_outputs(6249));
    layer1_outputs(4526) <= not(layer0_outputs(3296));
    layer1_outputs(4527) <= not((layer0_outputs(1720)) and (layer0_outputs(4961)));
    layer1_outputs(4528) <= not(layer0_outputs(9075)) or (layer0_outputs(2839));
    layer1_outputs(4529) <= not(layer0_outputs(9882)) or (layer0_outputs(8319));
    layer1_outputs(4530) <= (layer0_outputs(6284)) and not (layer0_outputs(304));
    layer1_outputs(4531) <= (layer0_outputs(6403)) and (layer0_outputs(4862));
    layer1_outputs(4532) <= (layer0_outputs(8045)) xor (layer0_outputs(2699));
    layer1_outputs(4533) <= layer0_outputs(6459);
    layer1_outputs(4534) <= not((layer0_outputs(1663)) and (layer0_outputs(903)));
    layer1_outputs(4535) <= not((layer0_outputs(8348)) or (layer0_outputs(8995)));
    layer1_outputs(4536) <= not((layer0_outputs(3844)) or (layer0_outputs(1204)));
    layer1_outputs(4537) <= not(layer0_outputs(6056)) or (layer0_outputs(5940));
    layer1_outputs(4538) <= not(layer0_outputs(9631));
    layer1_outputs(4539) <= not(layer0_outputs(8716)) or (layer0_outputs(3197));
    layer1_outputs(4540) <= '1';
    layer1_outputs(4541) <= layer0_outputs(5430);
    layer1_outputs(4542) <= not((layer0_outputs(2140)) or (layer0_outputs(3693)));
    layer1_outputs(4543) <= layer0_outputs(9800);
    layer1_outputs(4544) <= not(layer0_outputs(1461)) or (layer0_outputs(10210));
    layer1_outputs(4545) <= layer0_outputs(1055);
    layer1_outputs(4546) <= not((layer0_outputs(5221)) and (layer0_outputs(5642)));
    layer1_outputs(4547) <= (layer0_outputs(3329)) or (layer0_outputs(456));
    layer1_outputs(4548) <= layer0_outputs(8576);
    layer1_outputs(4549) <= not(layer0_outputs(3099)) or (layer0_outputs(3086));
    layer1_outputs(4550) <= (layer0_outputs(630)) or (layer0_outputs(2262));
    layer1_outputs(4551) <= not(layer0_outputs(8375)) or (layer0_outputs(2344));
    layer1_outputs(4552) <= not(layer0_outputs(4772)) or (layer0_outputs(3841));
    layer1_outputs(4553) <= (layer0_outputs(8964)) xor (layer0_outputs(7607));
    layer1_outputs(4554) <= not(layer0_outputs(1909)) or (layer0_outputs(1983));
    layer1_outputs(4555) <= layer0_outputs(4583);
    layer1_outputs(4556) <= '1';
    layer1_outputs(4557) <= layer0_outputs(4106);
    layer1_outputs(4558) <= not(layer0_outputs(7047));
    layer1_outputs(4559) <= (layer0_outputs(7045)) and (layer0_outputs(7238));
    layer1_outputs(4560) <= not(layer0_outputs(8483));
    layer1_outputs(4561) <= layer0_outputs(2288);
    layer1_outputs(4562) <= not(layer0_outputs(8935));
    layer1_outputs(4563) <= not((layer0_outputs(578)) and (layer0_outputs(1812)));
    layer1_outputs(4564) <= (layer0_outputs(4059)) and (layer0_outputs(9435));
    layer1_outputs(4565) <= (layer0_outputs(1153)) and not (layer0_outputs(5550));
    layer1_outputs(4566) <= (layer0_outputs(7764)) or (layer0_outputs(2442));
    layer1_outputs(4567) <= not((layer0_outputs(7625)) or (layer0_outputs(5895)));
    layer1_outputs(4568) <= layer0_outputs(10207);
    layer1_outputs(4569) <= (layer0_outputs(7720)) and (layer0_outputs(2366));
    layer1_outputs(4570) <= not(layer0_outputs(2596));
    layer1_outputs(4571) <= not(layer0_outputs(9382)) or (layer0_outputs(1583));
    layer1_outputs(4572) <= (layer0_outputs(8018)) and not (layer0_outputs(8215));
    layer1_outputs(4573) <= not(layer0_outputs(7666)) or (layer0_outputs(400));
    layer1_outputs(4574) <= '0';
    layer1_outputs(4575) <= (layer0_outputs(6157)) or (layer0_outputs(8998));
    layer1_outputs(4576) <= (layer0_outputs(7283)) xor (layer0_outputs(3397));
    layer1_outputs(4577) <= '1';
    layer1_outputs(4578) <= not(layer0_outputs(4751));
    layer1_outputs(4579) <= not(layer0_outputs(6305));
    layer1_outputs(4580) <= not(layer0_outputs(1657));
    layer1_outputs(4581) <= (layer0_outputs(604)) and not (layer0_outputs(419));
    layer1_outputs(4582) <= not((layer0_outputs(6081)) xor (layer0_outputs(3457)));
    layer1_outputs(4583) <= not(layer0_outputs(4598));
    layer1_outputs(4584) <= not((layer0_outputs(3695)) xor (layer0_outputs(2943)));
    layer1_outputs(4585) <= (layer0_outputs(3493)) and not (layer0_outputs(1154));
    layer1_outputs(4586) <= (layer0_outputs(7056)) xor (layer0_outputs(1890));
    layer1_outputs(4587) <= '0';
    layer1_outputs(4588) <= not(layer0_outputs(5520));
    layer1_outputs(4589) <= (layer0_outputs(349)) and not (layer0_outputs(5123));
    layer1_outputs(4590) <= (layer0_outputs(5915)) and not (layer0_outputs(5387));
    layer1_outputs(4591) <= '1';
    layer1_outputs(4592) <= (layer0_outputs(5443)) and (layer0_outputs(3159));
    layer1_outputs(4593) <= layer0_outputs(2714);
    layer1_outputs(4594) <= not(layer0_outputs(3216));
    layer1_outputs(4595) <= (layer0_outputs(7356)) and not (layer0_outputs(782));
    layer1_outputs(4596) <= not(layer0_outputs(7542));
    layer1_outputs(4597) <= not(layer0_outputs(5429));
    layer1_outputs(4598) <= not(layer0_outputs(1250));
    layer1_outputs(4599) <= not(layer0_outputs(8085));
    layer1_outputs(4600) <= not((layer0_outputs(622)) and (layer0_outputs(9633)));
    layer1_outputs(4601) <= '0';
    layer1_outputs(4602) <= (layer0_outputs(1961)) and not (layer0_outputs(2758));
    layer1_outputs(4603) <= layer0_outputs(2460);
    layer1_outputs(4604) <= not((layer0_outputs(8953)) or (layer0_outputs(1871)));
    layer1_outputs(4605) <= (layer0_outputs(2426)) and not (layer0_outputs(2140));
    layer1_outputs(4606) <= (layer0_outputs(2894)) or (layer0_outputs(2344));
    layer1_outputs(4607) <= (layer0_outputs(5080)) and not (layer0_outputs(354));
    layer1_outputs(4608) <= layer0_outputs(4360);
    layer1_outputs(4609) <= not(layer0_outputs(8661)) or (layer0_outputs(9096));
    layer1_outputs(4610) <= not((layer0_outputs(3914)) or (layer0_outputs(6201)));
    layer1_outputs(4611) <= (layer0_outputs(7269)) or (layer0_outputs(7153));
    layer1_outputs(4612) <= not(layer0_outputs(4113));
    layer1_outputs(4613) <= (layer0_outputs(1769)) and not (layer0_outputs(2687));
    layer1_outputs(4614) <= not((layer0_outputs(9591)) or (layer0_outputs(1454)));
    layer1_outputs(4615) <= not((layer0_outputs(9643)) or (layer0_outputs(2310)));
    layer1_outputs(4616) <= (layer0_outputs(7188)) and (layer0_outputs(1268));
    layer1_outputs(4617) <= not((layer0_outputs(5471)) xor (layer0_outputs(1491)));
    layer1_outputs(4618) <= layer0_outputs(523);
    layer1_outputs(4619) <= layer0_outputs(185);
    layer1_outputs(4620) <= not(layer0_outputs(512));
    layer1_outputs(4621) <= not(layer0_outputs(9791)) or (layer0_outputs(5447));
    layer1_outputs(4622) <= not(layer0_outputs(1468));
    layer1_outputs(4623) <= layer0_outputs(4363);
    layer1_outputs(4624) <= (layer0_outputs(6796)) and not (layer0_outputs(549));
    layer1_outputs(4625) <= (layer0_outputs(6670)) and not (layer0_outputs(791));
    layer1_outputs(4626) <= not((layer0_outputs(396)) and (layer0_outputs(191)));
    layer1_outputs(4627) <= not(layer0_outputs(167)) or (layer0_outputs(1525));
    layer1_outputs(4628) <= not(layer0_outputs(8531));
    layer1_outputs(4629) <= (layer0_outputs(9654)) xor (layer0_outputs(10072));
    layer1_outputs(4630) <= '0';
    layer1_outputs(4631) <= not((layer0_outputs(4673)) and (layer0_outputs(7692)));
    layer1_outputs(4632) <= layer0_outputs(9519);
    layer1_outputs(4633) <= (layer0_outputs(6468)) and not (layer0_outputs(6704));
    layer1_outputs(4634) <= (layer0_outputs(7491)) or (layer0_outputs(8294));
    layer1_outputs(4635) <= (layer0_outputs(8083)) or (layer0_outputs(4144));
    layer1_outputs(4636) <= not((layer0_outputs(1512)) or (layer0_outputs(2656)));
    layer1_outputs(4637) <= layer0_outputs(8632);
    layer1_outputs(4638) <= layer0_outputs(9555);
    layer1_outputs(4639) <= not(layer0_outputs(4031));
    layer1_outputs(4640) <= (layer0_outputs(9998)) and (layer0_outputs(8917));
    layer1_outputs(4641) <= not(layer0_outputs(1433)) or (layer0_outputs(3610));
    layer1_outputs(4642) <= not(layer0_outputs(9468));
    layer1_outputs(4643) <= not(layer0_outputs(6053));
    layer1_outputs(4644) <= not(layer0_outputs(4984));
    layer1_outputs(4645) <= (layer0_outputs(8095)) xor (layer0_outputs(5985));
    layer1_outputs(4646) <= '0';
    layer1_outputs(4647) <= (layer0_outputs(4543)) and not (layer0_outputs(5393));
    layer1_outputs(4648) <= not((layer0_outputs(646)) and (layer0_outputs(4617)));
    layer1_outputs(4649) <= not((layer0_outputs(2895)) or (layer0_outputs(9396)));
    layer1_outputs(4650) <= '0';
    layer1_outputs(4651) <= (layer0_outputs(5837)) or (layer0_outputs(6817));
    layer1_outputs(4652) <= '0';
    layer1_outputs(4653) <= not((layer0_outputs(4067)) xor (layer0_outputs(9068)));
    layer1_outputs(4654) <= not(layer0_outputs(5323));
    layer1_outputs(4655) <= layer0_outputs(7584);
    layer1_outputs(4656) <= '1';
    layer1_outputs(4657) <= (layer0_outputs(6218)) and not (layer0_outputs(4918));
    layer1_outputs(4658) <= not(layer0_outputs(4629)) or (layer0_outputs(6145));
    layer1_outputs(4659) <= not(layer0_outputs(5565)) or (layer0_outputs(7259));
    layer1_outputs(4660) <= (layer0_outputs(4074)) and not (layer0_outputs(6714));
    layer1_outputs(4661) <= '1';
    layer1_outputs(4662) <= not(layer0_outputs(6750)) or (layer0_outputs(5821));
    layer1_outputs(4663) <= layer0_outputs(6587);
    layer1_outputs(4664) <= (layer0_outputs(6861)) and (layer0_outputs(1050));
    layer1_outputs(4665) <= layer0_outputs(10188);
    layer1_outputs(4666) <= not(layer0_outputs(5913)) or (layer0_outputs(4356));
    layer1_outputs(4667) <= (layer0_outputs(929)) xor (layer0_outputs(7055));
    layer1_outputs(4668) <= not((layer0_outputs(3584)) xor (layer0_outputs(6505)));
    layer1_outputs(4669) <= not(layer0_outputs(5066));
    layer1_outputs(4670) <= layer0_outputs(1921);
    layer1_outputs(4671) <= not((layer0_outputs(8991)) or (layer0_outputs(8780)));
    layer1_outputs(4672) <= (layer0_outputs(1239)) or (layer0_outputs(9012));
    layer1_outputs(4673) <= not(layer0_outputs(3482));
    layer1_outputs(4674) <= not(layer0_outputs(697));
    layer1_outputs(4675) <= (layer0_outputs(4866)) and not (layer0_outputs(9107));
    layer1_outputs(4676) <= (layer0_outputs(460)) and not (layer0_outputs(6622));
    layer1_outputs(4677) <= not(layer0_outputs(5867)) or (layer0_outputs(4011));
    layer1_outputs(4678) <= (layer0_outputs(3502)) and not (layer0_outputs(8008));
    layer1_outputs(4679) <= layer0_outputs(10054);
    layer1_outputs(4680) <= layer0_outputs(9232);
    layer1_outputs(4681) <= not(layer0_outputs(5598));
    layer1_outputs(4682) <= layer0_outputs(505);
    layer1_outputs(4683) <= (layer0_outputs(4151)) and not (layer0_outputs(7336));
    layer1_outputs(4684) <= not((layer0_outputs(8814)) xor (layer0_outputs(410)));
    layer1_outputs(4685) <= (layer0_outputs(4647)) and not (layer0_outputs(4611));
    layer1_outputs(4686) <= (layer0_outputs(5995)) and (layer0_outputs(2327));
    layer1_outputs(4687) <= not((layer0_outputs(6796)) xor (layer0_outputs(3892)));
    layer1_outputs(4688) <= not(layer0_outputs(5795));
    layer1_outputs(4689) <= layer0_outputs(4899);
    layer1_outputs(4690) <= (layer0_outputs(8311)) xor (layer0_outputs(3889));
    layer1_outputs(4691) <= '1';
    layer1_outputs(4692) <= (layer0_outputs(3003)) and (layer0_outputs(8986));
    layer1_outputs(4693) <= not(layer0_outputs(5695)) or (layer0_outputs(7106));
    layer1_outputs(4694) <= not((layer0_outputs(2520)) xor (layer0_outputs(7315)));
    layer1_outputs(4695) <= '1';
    layer1_outputs(4696) <= not((layer0_outputs(6202)) and (layer0_outputs(2569)));
    layer1_outputs(4697) <= '0';
    layer1_outputs(4698) <= not(layer0_outputs(2721));
    layer1_outputs(4699) <= layer0_outputs(7158);
    layer1_outputs(4700) <= not(layer0_outputs(8141)) or (layer0_outputs(7835));
    layer1_outputs(4701) <= not((layer0_outputs(5566)) xor (layer0_outputs(8979)));
    layer1_outputs(4702) <= not(layer0_outputs(6618));
    layer1_outputs(4703) <= not(layer0_outputs(114));
    layer1_outputs(4704) <= not(layer0_outputs(2927)) or (layer0_outputs(3581));
    layer1_outputs(4705) <= not(layer0_outputs(6231)) or (layer0_outputs(1482));
    layer1_outputs(4706) <= (layer0_outputs(7608)) and (layer0_outputs(6327));
    layer1_outputs(4707) <= (layer0_outputs(1729)) and not (layer0_outputs(4083));
    layer1_outputs(4708) <= layer0_outputs(7085);
    layer1_outputs(4709) <= layer0_outputs(8848);
    layer1_outputs(4710) <= (layer0_outputs(4551)) and (layer0_outputs(4881));
    layer1_outputs(4711) <= (layer0_outputs(6610)) xor (layer0_outputs(1480));
    layer1_outputs(4712) <= not(layer0_outputs(2760));
    layer1_outputs(4713) <= (layer0_outputs(6579)) and not (layer0_outputs(3072));
    layer1_outputs(4714) <= not(layer0_outputs(7478)) or (layer0_outputs(6911));
    layer1_outputs(4715) <= layer0_outputs(8241);
    layer1_outputs(4716) <= (layer0_outputs(9484)) and not (layer0_outputs(5343));
    layer1_outputs(4717) <= (layer0_outputs(1294)) and (layer0_outputs(3349));
    layer1_outputs(4718) <= (layer0_outputs(9016)) and (layer0_outputs(9961));
    layer1_outputs(4719) <= not((layer0_outputs(5914)) and (layer0_outputs(3867)));
    layer1_outputs(4720) <= not(layer0_outputs(8566));
    layer1_outputs(4721) <= not((layer0_outputs(3121)) or (layer0_outputs(2190)));
    layer1_outputs(4722) <= (layer0_outputs(6544)) and not (layer0_outputs(4594));
    layer1_outputs(4723) <= not(layer0_outputs(8586));
    layer1_outputs(4724) <= not(layer0_outputs(879)) or (layer0_outputs(3208));
    layer1_outputs(4725) <= not(layer0_outputs(3445)) or (layer0_outputs(2314));
    layer1_outputs(4726) <= (layer0_outputs(1305)) xor (layer0_outputs(9345));
    layer1_outputs(4727) <= '1';
    layer1_outputs(4728) <= layer0_outputs(1273);
    layer1_outputs(4729) <= not(layer0_outputs(1740));
    layer1_outputs(4730) <= (layer0_outputs(3649)) and (layer0_outputs(3150));
    layer1_outputs(4731) <= (layer0_outputs(9870)) or (layer0_outputs(2920));
    layer1_outputs(4732) <= not(layer0_outputs(6638)) or (layer0_outputs(7510));
    layer1_outputs(4733) <= (layer0_outputs(911)) or (layer0_outputs(7673));
    layer1_outputs(4734) <= not(layer0_outputs(8946));
    layer1_outputs(4735) <= not(layer0_outputs(4087)) or (layer0_outputs(4745));
    layer1_outputs(4736) <= not(layer0_outputs(3409));
    layer1_outputs(4737) <= not(layer0_outputs(6372)) or (layer0_outputs(8));
    layer1_outputs(4738) <= layer0_outputs(3188);
    layer1_outputs(4739) <= '0';
    layer1_outputs(4740) <= (layer0_outputs(4153)) and not (layer0_outputs(5216));
    layer1_outputs(4741) <= layer0_outputs(5500);
    layer1_outputs(4742) <= (layer0_outputs(6136)) and not (layer0_outputs(7051));
    layer1_outputs(4743) <= not(layer0_outputs(1986));
    layer1_outputs(4744) <= layer0_outputs(9969);
    layer1_outputs(4745) <= not(layer0_outputs(6178)) or (layer0_outputs(3357));
    layer1_outputs(4746) <= not(layer0_outputs(3142));
    layer1_outputs(4747) <= '0';
    layer1_outputs(4748) <= (layer0_outputs(461)) and not (layer0_outputs(5375));
    layer1_outputs(4749) <= (layer0_outputs(5887)) or (layer0_outputs(6217));
    layer1_outputs(4750) <= '0';
    layer1_outputs(4751) <= (layer0_outputs(3265)) xor (layer0_outputs(1176));
    layer1_outputs(4752) <= layer0_outputs(1054);
    layer1_outputs(4753) <= not(layer0_outputs(2305)) or (layer0_outputs(5357));
    layer1_outputs(4754) <= layer0_outputs(5484);
    layer1_outputs(4755) <= not(layer0_outputs(8624)) or (layer0_outputs(7697));
    layer1_outputs(4756) <= layer0_outputs(3047);
    layer1_outputs(4757) <= not((layer0_outputs(4055)) and (layer0_outputs(528)));
    layer1_outputs(4758) <= (layer0_outputs(482)) and not (layer0_outputs(7130));
    layer1_outputs(4759) <= (layer0_outputs(8115)) and (layer0_outputs(3499));
    layer1_outputs(4760) <= (layer0_outputs(9276)) and not (layer0_outputs(7044));
    layer1_outputs(4761) <= not(layer0_outputs(9377)) or (layer0_outputs(511));
    layer1_outputs(4762) <= not((layer0_outputs(4169)) xor (layer0_outputs(2880)));
    layer1_outputs(4763) <= layer0_outputs(6066);
    layer1_outputs(4764) <= not((layer0_outputs(10232)) and (layer0_outputs(446)));
    layer1_outputs(4765) <= (layer0_outputs(4865)) and (layer0_outputs(2910));
    layer1_outputs(4766) <= (layer0_outputs(2238)) and not (layer0_outputs(4966));
    layer1_outputs(4767) <= not((layer0_outputs(3599)) and (layer0_outputs(7616)));
    layer1_outputs(4768) <= not((layer0_outputs(9330)) or (layer0_outputs(6980)));
    layer1_outputs(4769) <= not(layer0_outputs(6919));
    layer1_outputs(4770) <= '1';
    layer1_outputs(4771) <= (layer0_outputs(716)) and (layer0_outputs(92));
    layer1_outputs(4772) <= not(layer0_outputs(6719)) or (layer0_outputs(6434));
    layer1_outputs(4773) <= layer0_outputs(134);
    layer1_outputs(4774) <= not(layer0_outputs(4463)) or (layer0_outputs(3749));
    layer1_outputs(4775) <= not(layer0_outputs(6417));
    layer1_outputs(4776) <= not(layer0_outputs(9637));
    layer1_outputs(4777) <= (layer0_outputs(4423)) or (layer0_outputs(8413));
    layer1_outputs(4778) <= layer0_outputs(9505);
    layer1_outputs(4779) <= (layer0_outputs(1767)) and not (layer0_outputs(6387));
    layer1_outputs(4780) <= (layer0_outputs(10227)) and not (layer0_outputs(264));
    layer1_outputs(4781) <= (layer0_outputs(7798)) and (layer0_outputs(3696));
    layer1_outputs(4782) <= not(layer0_outputs(7524)) or (layer0_outputs(39));
    layer1_outputs(4783) <= '1';
    layer1_outputs(4784) <= (layer0_outputs(2916)) or (layer0_outputs(1260));
    layer1_outputs(4785) <= not((layer0_outputs(1193)) or (layer0_outputs(3270)));
    layer1_outputs(4786) <= layer0_outputs(373);
    layer1_outputs(4787) <= (layer0_outputs(8860)) xor (layer0_outputs(6650));
    layer1_outputs(4788) <= not(layer0_outputs(2480));
    layer1_outputs(4789) <= (layer0_outputs(64)) xor (layer0_outputs(5233));
    layer1_outputs(4790) <= (layer0_outputs(6637)) and (layer0_outputs(4281));
    layer1_outputs(4791) <= (layer0_outputs(3001)) or (layer0_outputs(4028));
    layer1_outputs(4792) <= not((layer0_outputs(1393)) and (layer0_outputs(972)));
    layer1_outputs(4793) <= not((layer0_outputs(4685)) and (layer0_outputs(7904)));
    layer1_outputs(4794) <= (layer0_outputs(413)) or (layer0_outputs(10091));
    layer1_outputs(4795) <= (layer0_outputs(2054)) and not (layer0_outputs(9649));
    layer1_outputs(4796) <= '1';
    layer1_outputs(4797) <= '1';
    layer1_outputs(4798) <= (layer0_outputs(3711)) or (layer0_outputs(4497));
    layer1_outputs(4799) <= not((layer0_outputs(6455)) xor (layer0_outputs(3025)));
    layer1_outputs(4800) <= not(layer0_outputs(8062)) or (layer0_outputs(10134));
    layer1_outputs(4801) <= not(layer0_outputs(463));
    layer1_outputs(4802) <= not(layer0_outputs(7836));
    layer1_outputs(4803) <= not(layer0_outputs(7288));
    layer1_outputs(4804) <= layer0_outputs(284);
    layer1_outputs(4805) <= (layer0_outputs(5729)) xor (layer0_outputs(7551));
    layer1_outputs(4806) <= not(layer0_outputs(6079));
    layer1_outputs(4807) <= not(layer0_outputs(6752));
    layer1_outputs(4808) <= not(layer0_outputs(302));
    layer1_outputs(4809) <= layer0_outputs(5400);
    layer1_outputs(4810) <= not(layer0_outputs(8283)) or (layer0_outputs(6212));
    layer1_outputs(4811) <= layer0_outputs(9941);
    layer1_outputs(4812) <= not((layer0_outputs(4801)) xor (layer0_outputs(9440)));
    layer1_outputs(4813) <= layer0_outputs(3965);
    layer1_outputs(4814) <= '1';
    layer1_outputs(4815) <= (layer0_outputs(7964)) or (layer0_outputs(3916));
    layer1_outputs(4816) <= not(layer0_outputs(8213)) or (layer0_outputs(6265));
    layer1_outputs(4817) <= not(layer0_outputs(1337));
    layer1_outputs(4818) <= not(layer0_outputs(4071));
    layer1_outputs(4819) <= (layer0_outputs(3713)) and (layer0_outputs(4103));
    layer1_outputs(4820) <= not((layer0_outputs(8323)) and (layer0_outputs(3700)));
    layer1_outputs(4821) <= (layer0_outputs(8831)) or (layer0_outputs(1077));
    layer1_outputs(4822) <= (layer0_outputs(101)) and not (layer0_outputs(4898));
    layer1_outputs(4823) <= '1';
    layer1_outputs(4824) <= not((layer0_outputs(9937)) and (layer0_outputs(7265)));
    layer1_outputs(4825) <= not((layer0_outputs(8051)) and (layer0_outputs(2327)));
    layer1_outputs(4826) <= not((layer0_outputs(6935)) or (layer0_outputs(9274)));
    layer1_outputs(4827) <= (layer0_outputs(2780)) and not (layer0_outputs(1764));
    layer1_outputs(4828) <= '0';
    layer1_outputs(4829) <= (layer0_outputs(571)) or (layer0_outputs(1483));
    layer1_outputs(4830) <= (layer0_outputs(7461)) or (layer0_outputs(648));
    layer1_outputs(4831) <= not((layer0_outputs(8119)) and (layer0_outputs(3070)));
    layer1_outputs(4832) <= (layer0_outputs(7450)) and not (layer0_outputs(8896));
    layer1_outputs(4833) <= '1';
    layer1_outputs(4834) <= (layer0_outputs(8461)) and not (layer0_outputs(5144));
    layer1_outputs(4835) <= not((layer0_outputs(905)) or (layer0_outputs(5620)));
    layer1_outputs(4836) <= (layer0_outputs(7141)) and not (layer0_outputs(9315));
    layer1_outputs(4837) <= (layer0_outputs(389)) xor (layer0_outputs(1448));
    layer1_outputs(4838) <= '1';
    layer1_outputs(4839) <= not((layer0_outputs(74)) and (layer0_outputs(1427)));
    layer1_outputs(4840) <= not((layer0_outputs(485)) and (layer0_outputs(6738)));
    layer1_outputs(4841) <= (layer0_outputs(4639)) or (layer0_outputs(6850));
    layer1_outputs(4842) <= not((layer0_outputs(7452)) or (layer0_outputs(7441)));
    layer1_outputs(4843) <= (layer0_outputs(8062)) or (layer0_outputs(10063));
    layer1_outputs(4844) <= not(layer0_outputs(7522));
    layer1_outputs(4845) <= (layer0_outputs(10151)) or (layer0_outputs(9982));
    layer1_outputs(4846) <= (layer0_outputs(4840)) and (layer0_outputs(1835));
    layer1_outputs(4847) <= (layer0_outputs(5886)) and not (layer0_outputs(7787));
    layer1_outputs(4848) <= not((layer0_outputs(1382)) or (layer0_outputs(3839)));
    layer1_outputs(4849) <= (layer0_outputs(7988)) and not (layer0_outputs(5053));
    layer1_outputs(4850) <= (layer0_outputs(7770)) and not (layer0_outputs(7035));
    layer1_outputs(4851) <= layer0_outputs(6314);
    layer1_outputs(4852) <= (layer0_outputs(1075)) and (layer0_outputs(9815));
    layer1_outputs(4853) <= (layer0_outputs(4835)) and not (layer0_outputs(6125));
    layer1_outputs(4854) <= '0';
    layer1_outputs(4855) <= not(layer0_outputs(8662)) or (layer0_outputs(5070));
    layer1_outputs(4856) <= not(layer0_outputs(579)) or (layer0_outputs(7781));
    layer1_outputs(4857) <= not(layer0_outputs(194));
    layer1_outputs(4858) <= layer0_outputs(3446);
    layer1_outputs(4859) <= layer0_outputs(8387);
    layer1_outputs(4860) <= layer0_outputs(7234);
    layer1_outputs(4861) <= not((layer0_outputs(5104)) and (layer0_outputs(406)));
    layer1_outputs(4862) <= not((layer0_outputs(5496)) and (layer0_outputs(903)));
    layer1_outputs(4863) <= (layer0_outputs(9800)) and (layer0_outputs(8499));
    layer1_outputs(4864) <= not(layer0_outputs(2291));
    layer1_outputs(4865) <= (layer0_outputs(916)) and not (layer0_outputs(4231));
    layer1_outputs(4866) <= (layer0_outputs(9868)) and (layer0_outputs(7009));
    layer1_outputs(4867) <= layer0_outputs(1751);
    layer1_outputs(4868) <= '0';
    layer1_outputs(4869) <= not(layer0_outputs(2702)) or (layer0_outputs(7411));
    layer1_outputs(4870) <= layer0_outputs(6632);
    layer1_outputs(4871) <= layer0_outputs(62);
    layer1_outputs(4872) <= layer0_outputs(143);
    layer1_outputs(4873) <= not(layer0_outputs(2576));
    layer1_outputs(4874) <= layer0_outputs(7671);
    layer1_outputs(4875) <= not((layer0_outputs(2621)) xor (layer0_outputs(8750)));
    layer1_outputs(4876) <= not(layer0_outputs(1863));
    layer1_outputs(4877) <= '1';
    layer1_outputs(4878) <= (layer0_outputs(2573)) and not (layer0_outputs(9033));
    layer1_outputs(4879) <= (layer0_outputs(7036)) and not (layer0_outputs(5137));
    layer1_outputs(4880) <= not(layer0_outputs(980));
    layer1_outputs(4881) <= not((layer0_outputs(2345)) xor (layer0_outputs(3445)));
    layer1_outputs(4882) <= not((layer0_outputs(6247)) and (layer0_outputs(9104)));
    layer1_outputs(4883) <= layer0_outputs(2404);
    layer1_outputs(4884) <= not(layer0_outputs(4199)) or (layer0_outputs(8588));
    layer1_outputs(4885) <= (layer0_outputs(542)) or (layer0_outputs(1255));
    layer1_outputs(4886) <= not((layer0_outputs(7209)) and (layer0_outputs(6460)));
    layer1_outputs(4887) <= (layer0_outputs(9057)) or (layer0_outputs(1452));
    layer1_outputs(4888) <= layer0_outputs(6487);
    layer1_outputs(4889) <= not(layer0_outputs(4134));
    layer1_outputs(4890) <= not((layer0_outputs(5273)) or (layer0_outputs(2592)));
    layer1_outputs(4891) <= (layer0_outputs(7490)) or (layer0_outputs(6599));
    layer1_outputs(4892) <= (layer0_outputs(7492)) and not (layer0_outputs(4238));
    layer1_outputs(4893) <= not((layer0_outputs(5368)) and (layer0_outputs(2690)));
    layer1_outputs(4894) <= (layer0_outputs(5886)) or (layer0_outputs(7245));
    layer1_outputs(4895) <= layer0_outputs(6606);
    layer1_outputs(4896) <= (layer0_outputs(2732)) or (layer0_outputs(1508));
    layer1_outputs(4897) <= (layer0_outputs(1039)) xor (layer0_outputs(8461));
    layer1_outputs(4898) <= not(layer0_outputs(6637)) or (layer0_outputs(1570));
    layer1_outputs(4899) <= not((layer0_outputs(5103)) and (layer0_outputs(7676)));
    layer1_outputs(4900) <= not((layer0_outputs(9292)) or (layer0_outputs(9316)));
    layer1_outputs(4901) <= (layer0_outputs(1226)) and not (layer0_outputs(8155));
    layer1_outputs(4902) <= (layer0_outputs(2565)) and not (layer0_outputs(6656));
    layer1_outputs(4903) <= not((layer0_outputs(7399)) or (layer0_outputs(9676)));
    layer1_outputs(4904) <= '0';
    layer1_outputs(4905) <= (layer0_outputs(3885)) or (layer0_outputs(2363));
    layer1_outputs(4906) <= layer0_outputs(3433);
    layer1_outputs(4907) <= not(layer0_outputs(9607));
    layer1_outputs(4908) <= not(layer0_outputs(8279)) or (layer0_outputs(9527));
    layer1_outputs(4909) <= not(layer0_outputs(9321));
    layer1_outputs(4910) <= (layer0_outputs(3831)) and (layer0_outputs(3443));
    layer1_outputs(4911) <= not(layer0_outputs(5254)) or (layer0_outputs(2290));
    layer1_outputs(4912) <= layer0_outputs(262);
    layer1_outputs(4913) <= (layer0_outputs(2632)) xor (layer0_outputs(5409));
    layer1_outputs(4914) <= not((layer0_outputs(3899)) or (layer0_outputs(237)));
    layer1_outputs(4915) <= (layer0_outputs(9181)) and not (layer0_outputs(9853));
    layer1_outputs(4916) <= '0';
    layer1_outputs(4917) <= not((layer0_outputs(1581)) and (layer0_outputs(1552)));
    layer1_outputs(4918) <= not((layer0_outputs(5075)) and (layer0_outputs(8565)));
    layer1_outputs(4919) <= layer0_outputs(9068);
    layer1_outputs(4920) <= not((layer0_outputs(2815)) and (layer0_outputs(6660)));
    layer1_outputs(4921) <= not((layer0_outputs(6513)) xor (layer0_outputs(8792)));
    layer1_outputs(4922) <= not(layer0_outputs(7016));
    layer1_outputs(4923) <= layer0_outputs(1273);
    layer1_outputs(4924) <= not(layer0_outputs(3171)) or (layer0_outputs(4450));
    layer1_outputs(4925) <= (layer0_outputs(3692)) or (layer0_outputs(5770));
    layer1_outputs(4926) <= not(layer0_outputs(4977));
    layer1_outputs(4927) <= (layer0_outputs(10089)) and (layer0_outputs(5287));
    layer1_outputs(4928) <= '0';
    layer1_outputs(4929) <= not((layer0_outputs(3044)) and (layer0_outputs(7084)));
    layer1_outputs(4930) <= not((layer0_outputs(5802)) and (layer0_outputs(5808)));
    layer1_outputs(4931) <= not(layer0_outputs(6649));
    layer1_outputs(4932) <= (layer0_outputs(9634)) and (layer0_outputs(324));
    layer1_outputs(4933) <= not((layer0_outputs(6077)) and (layer0_outputs(7334)));
    layer1_outputs(4934) <= (layer0_outputs(9834)) and not (layer0_outputs(5261));
    layer1_outputs(4935) <= not((layer0_outputs(2841)) or (layer0_outputs(6941)));
    layer1_outputs(4936) <= not(layer0_outputs(9773)) or (layer0_outputs(9010));
    layer1_outputs(4937) <= '0';
    layer1_outputs(4938) <= not(layer0_outputs(5331));
    layer1_outputs(4939) <= not(layer0_outputs(8512));
    layer1_outputs(4940) <= (layer0_outputs(6542)) xor (layer0_outputs(4569));
    layer1_outputs(4941) <= not((layer0_outputs(5781)) or (layer0_outputs(7142)));
    layer1_outputs(4942) <= (layer0_outputs(9209)) and (layer0_outputs(235));
    layer1_outputs(4943) <= '0';
    layer1_outputs(4944) <= layer0_outputs(9624);
    layer1_outputs(4945) <= layer0_outputs(8986);
    layer1_outputs(4946) <= (layer0_outputs(6929)) and not (layer0_outputs(5114));
    layer1_outputs(4947) <= layer0_outputs(7318);
    layer1_outputs(4948) <= (layer0_outputs(3524)) and not (layer0_outputs(5479));
    layer1_outputs(4949) <= not(layer0_outputs(8752)) or (layer0_outputs(9939));
    layer1_outputs(4950) <= (layer0_outputs(5513)) and not (layer0_outputs(8309));
    layer1_outputs(4951) <= (layer0_outputs(4862)) xor (layer0_outputs(4412));
    layer1_outputs(4952) <= layer0_outputs(9785);
    layer1_outputs(4953) <= not(layer0_outputs(1627));
    layer1_outputs(4954) <= not(layer0_outputs(2094));
    layer1_outputs(4955) <= '1';
    layer1_outputs(4956) <= (layer0_outputs(4385)) and not (layer0_outputs(6863));
    layer1_outputs(4957) <= (layer0_outputs(9490)) and not (layer0_outputs(2862));
    layer1_outputs(4958) <= layer0_outputs(8223);
    layer1_outputs(4959) <= not(layer0_outputs(1768)) or (layer0_outputs(2481));
    layer1_outputs(4960) <= not((layer0_outputs(4683)) or (layer0_outputs(6354)));
    layer1_outputs(4961) <= not((layer0_outputs(8854)) or (layer0_outputs(2439)));
    layer1_outputs(4962) <= '1';
    layer1_outputs(4963) <= (layer0_outputs(2517)) or (layer0_outputs(5055));
    layer1_outputs(4964) <= (layer0_outputs(7767)) or (layer0_outputs(8726));
    layer1_outputs(4965) <= not((layer0_outputs(517)) or (layer0_outputs(2679)));
    layer1_outputs(4966) <= not(layer0_outputs(3465));
    layer1_outputs(4967) <= '1';
    layer1_outputs(4968) <= layer0_outputs(5133);
    layer1_outputs(4969) <= layer0_outputs(7946);
    layer1_outputs(4970) <= not(layer0_outputs(838));
    layer1_outputs(4971) <= (layer0_outputs(3752)) or (layer0_outputs(4752));
    layer1_outputs(4972) <= (layer0_outputs(1940)) or (layer0_outputs(124));
    layer1_outputs(4973) <= not(layer0_outputs(3699));
    layer1_outputs(4974) <= (layer0_outputs(677)) and not (layer0_outputs(2281));
    layer1_outputs(4975) <= not(layer0_outputs(9563)) or (layer0_outputs(1564));
    layer1_outputs(4976) <= layer0_outputs(4920);
    layer1_outputs(4977) <= not((layer0_outputs(2500)) and (layer0_outputs(4415)));
    layer1_outputs(4978) <= (layer0_outputs(9580)) and not (layer0_outputs(6512));
    layer1_outputs(4979) <= (layer0_outputs(3846)) and not (layer0_outputs(9225));
    layer1_outputs(4980) <= not((layer0_outputs(6951)) or (layer0_outputs(4693)));
    layer1_outputs(4981) <= (layer0_outputs(7368)) and (layer0_outputs(5503));
    layer1_outputs(4982) <= layer0_outputs(8651);
    layer1_outputs(4983) <= '0';
    layer1_outputs(4984) <= (layer0_outputs(57)) xor (layer0_outputs(1185));
    layer1_outputs(4985) <= not(layer0_outputs(9889));
    layer1_outputs(4986) <= not(layer0_outputs(4340));
    layer1_outputs(4987) <= not(layer0_outputs(4365));
    layer1_outputs(4988) <= not(layer0_outputs(4410)) or (layer0_outputs(9439));
    layer1_outputs(4989) <= (layer0_outputs(7925)) and (layer0_outputs(1520));
    layer1_outputs(4990) <= '0';
    layer1_outputs(4991) <= not(layer0_outputs(2058)) or (layer0_outputs(16));
    layer1_outputs(4992) <= not(layer0_outputs(1270)) or (layer0_outputs(3277));
    layer1_outputs(4993) <= (layer0_outputs(3854)) xor (layer0_outputs(4528));
    layer1_outputs(4994) <= (layer0_outputs(1691)) and not (layer0_outputs(616));
    layer1_outputs(4995) <= layer0_outputs(1743);
    layer1_outputs(4996) <= not(layer0_outputs(5167)) or (layer0_outputs(7669));
    layer1_outputs(4997) <= not(layer0_outputs(1460));
    layer1_outputs(4998) <= not(layer0_outputs(1781));
    layer1_outputs(4999) <= (layer0_outputs(3573)) or (layer0_outputs(7377));
    layer1_outputs(5000) <= not((layer0_outputs(8003)) xor (layer0_outputs(8610)));
    layer1_outputs(5001) <= '0';
    layer1_outputs(5002) <= not((layer0_outputs(5899)) xor (layer0_outputs(3278)));
    layer1_outputs(5003) <= (layer0_outputs(1332)) and not (layer0_outputs(9326));
    layer1_outputs(5004) <= not(layer0_outputs(4331)) or (layer0_outputs(10231));
    layer1_outputs(5005) <= (layer0_outputs(10217)) xor (layer0_outputs(4622));
    layer1_outputs(5006) <= not(layer0_outputs(4485));
    layer1_outputs(5007) <= (layer0_outputs(9281)) and not (layer0_outputs(4023));
    layer1_outputs(5008) <= not(layer0_outputs(2467));
    layer1_outputs(5009) <= not(layer0_outputs(9914)) or (layer0_outputs(5848));
    layer1_outputs(5010) <= layer0_outputs(9487);
    layer1_outputs(5011) <= not((layer0_outputs(8316)) and (layer0_outputs(7881)));
    layer1_outputs(5012) <= layer0_outputs(10116);
    layer1_outputs(5013) <= not((layer0_outputs(5508)) and (layer0_outputs(7247)));
    layer1_outputs(5014) <= not(layer0_outputs(9492));
    layer1_outputs(5015) <= not(layer0_outputs(1714)) or (layer0_outputs(6979));
    layer1_outputs(5016) <= (layer0_outputs(3237)) or (layer0_outputs(8425));
    layer1_outputs(5017) <= not((layer0_outputs(3500)) or (layer0_outputs(9133)));
    layer1_outputs(5018) <= not(layer0_outputs(1118)) or (layer0_outputs(9574));
    layer1_outputs(5019) <= layer0_outputs(6763);
    layer1_outputs(5020) <= '1';
    layer1_outputs(5021) <= layer0_outputs(6032);
    layer1_outputs(5022) <= layer0_outputs(739);
    layer1_outputs(5023) <= '0';
    layer1_outputs(5024) <= (layer0_outputs(2623)) and not (layer0_outputs(3367));
    layer1_outputs(5025) <= not(layer0_outputs(5755)) or (layer0_outputs(3071));
    layer1_outputs(5026) <= not(layer0_outputs(6498)) or (layer0_outputs(3622));
    layer1_outputs(5027) <= (layer0_outputs(2761)) and (layer0_outputs(9354));
    layer1_outputs(5028) <= not(layer0_outputs(9199));
    layer1_outputs(5029) <= (layer0_outputs(8785)) or (layer0_outputs(4255));
    layer1_outputs(5030) <= not(layer0_outputs(7090)) or (layer0_outputs(911));
    layer1_outputs(5031) <= not(layer0_outputs(5407)) or (layer0_outputs(3798));
    layer1_outputs(5032) <= layer0_outputs(9564);
    layer1_outputs(5033) <= not(layer0_outputs(2646));
    layer1_outputs(5034) <= (layer0_outputs(8070)) and not (layer0_outputs(6433));
    layer1_outputs(5035) <= (layer0_outputs(2628)) xor (layer0_outputs(9197));
    layer1_outputs(5036) <= '1';
    layer1_outputs(5037) <= not(layer0_outputs(6497));
    layer1_outputs(5038) <= '0';
    layer1_outputs(5039) <= layer0_outputs(3410);
    layer1_outputs(5040) <= not(layer0_outputs(2164)) or (layer0_outputs(9499));
    layer1_outputs(5041) <= layer0_outputs(1359);
    layer1_outputs(5042) <= (layer0_outputs(5269)) and (layer0_outputs(5814));
    layer1_outputs(5043) <= not(layer0_outputs(3307)) or (layer0_outputs(2917));
    layer1_outputs(5044) <= not((layer0_outputs(736)) xor (layer0_outputs(8036)));
    layer1_outputs(5045) <= layer0_outputs(3527);
    layer1_outputs(5046) <= '0';
    layer1_outputs(5047) <= (layer0_outputs(1103)) and not (layer0_outputs(2064));
    layer1_outputs(5048) <= (layer0_outputs(5943)) and not (layer0_outputs(8067));
    layer1_outputs(5049) <= '0';
    layer1_outputs(5050) <= (layer0_outputs(8370)) and not (layer0_outputs(1350));
    layer1_outputs(5051) <= not((layer0_outputs(10067)) or (layer0_outputs(2405)));
    layer1_outputs(5052) <= layer0_outputs(1612);
    layer1_outputs(5053) <= not(layer0_outputs(1536));
    layer1_outputs(5054) <= layer0_outputs(2111);
    layer1_outputs(5055) <= not(layer0_outputs(8354));
    layer1_outputs(5056) <= (layer0_outputs(4140)) xor (layer0_outputs(9475));
    layer1_outputs(5057) <= layer0_outputs(1215);
    layer1_outputs(5058) <= (layer0_outputs(110)) or (layer0_outputs(1983));
    layer1_outputs(5059) <= layer0_outputs(8881);
    layer1_outputs(5060) <= (layer0_outputs(2588)) and not (layer0_outputs(108));
    layer1_outputs(5061) <= not(layer0_outputs(1338)) or (layer0_outputs(9946));
    layer1_outputs(5062) <= not(layer0_outputs(3950));
    layer1_outputs(5063) <= not(layer0_outputs(6204)) or (layer0_outputs(4090));
    layer1_outputs(5064) <= not(layer0_outputs(8490));
    layer1_outputs(5065) <= not((layer0_outputs(3553)) xor (layer0_outputs(1873)));
    layer1_outputs(5066) <= '1';
    layer1_outputs(5067) <= (layer0_outputs(3217)) and (layer0_outputs(7211));
    layer1_outputs(5068) <= (layer0_outputs(7545)) and not (layer0_outputs(9493));
    layer1_outputs(5069) <= not(layer0_outputs(965)) or (layer0_outputs(2053));
    layer1_outputs(5070) <= not(layer0_outputs(8409)) or (layer0_outputs(10198));
    layer1_outputs(5071) <= (layer0_outputs(3400)) and not (layer0_outputs(6038));
    layer1_outputs(5072) <= not(layer0_outputs(1158));
    layer1_outputs(5073) <= (layer0_outputs(1768)) and not (layer0_outputs(1513));
    layer1_outputs(5074) <= (layer0_outputs(7220)) and (layer0_outputs(7848));
    layer1_outputs(5075) <= not(layer0_outputs(8316));
    layer1_outputs(5076) <= (layer0_outputs(8361)) or (layer0_outputs(1014));
    layer1_outputs(5077) <= not(layer0_outputs(6530));
    layer1_outputs(5078) <= layer0_outputs(223);
    layer1_outputs(5079) <= (layer0_outputs(1028)) or (layer0_outputs(1278));
    layer1_outputs(5080) <= not((layer0_outputs(3773)) or (layer0_outputs(9740)));
    layer1_outputs(5081) <= (layer0_outputs(5140)) or (layer0_outputs(8825));
    layer1_outputs(5082) <= (layer0_outputs(9682)) xor (layer0_outputs(4641));
    layer1_outputs(5083) <= layer0_outputs(1763);
    layer1_outputs(5084) <= (layer0_outputs(6985)) and not (layer0_outputs(1891));
    layer1_outputs(5085) <= not(layer0_outputs(3964));
    layer1_outputs(5086) <= not(layer0_outputs(2521));
    layer1_outputs(5087) <= (layer0_outputs(4498)) xor (layer0_outputs(7814));
    layer1_outputs(5088) <= (layer0_outputs(9277)) and not (layer0_outputs(5707));
    layer1_outputs(5089) <= layer0_outputs(1343);
    layer1_outputs(5090) <= (layer0_outputs(3744)) or (layer0_outputs(2453));
    layer1_outputs(5091) <= '0';
    layer1_outputs(5092) <= layer0_outputs(2434);
    layer1_outputs(5093) <= (layer0_outputs(815)) or (layer0_outputs(1849));
    layer1_outputs(5094) <= layer0_outputs(21);
    layer1_outputs(5095) <= '0';
    layer1_outputs(5096) <= (layer0_outputs(4421)) or (layer0_outputs(9878));
    layer1_outputs(5097) <= not(layer0_outputs(10114));
    layer1_outputs(5098) <= (layer0_outputs(3064)) or (layer0_outputs(1967));
    layer1_outputs(5099) <= (layer0_outputs(7331)) and (layer0_outputs(772));
    layer1_outputs(5100) <= '1';
    layer1_outputs(5101) <= not((layer0_outputs(3943)) or (layer0_outputs(1336)));
    layer1_outputs(5102) <= layer0_outputs(2725);
    layer1_outputs(5103) <= layer0_outputs(1680);
    layer1_outputs(5104) <= not(layer0_outputs(171));
    layer1_outputs(5105) <= not(layer0_outputs(2737));
    layer1_outputs(5106) <= (layer0_outputs(9228)) and (layer0_outputs(8122));
    layer1_outputs(5107) <= not(layer0_outputs(9565));
    layer1_outputs(5108) <= (layer0_outputs(10181)) xor (layer0_outputs(4029));
    layer1_outputs(5109) <= (layer0_outputs(9877)) and not (layer0_outputs(2948));
    layer1_outputs(5110) <= not(layer0_outputs(8257));
    layer1_outputs(5111) <= not(layer0_outputs(3188)) or (layer0_outputs(8180));
    layer1_outputs(5112) <= not(layer0_outputs(7279));
    layer1_outputs(5113) <= layer0_outputs(9799);
    layer1_outputs(5114) <= (layer0_outputs(8668)) and (layer0_outputs(5746));
    layer1_outputs(5115) <= (layer0_outputs(5587)) and not (layer0_outputs(2506));
    layer1_outputs(5116) <= layer0_outputs(5149);
    layer1_outputs(5117) <= not(layer0_outputs(5420)) or (layer0_outputs(2154));
    layer1_outputs(5118) <= (layer0_outputs(5719)) and not (layer0_outputs(8840));
    layer1_outputs(5119) <= (layer0_outputs(9836)) or (layer0_outputs(1963));
    layer1_outputs(5120) <= layer0_outputs(9266);
    layer1_outputs(5121) <= not((layer0_outputs(6211)) xor (layer0_outputs(5907)));
    layer1_outputs(5122) <= layer0_outputs(2961);
    layer1_outputs(5123) <= layer0_outputs(9043);
    layer1_outputs(5124) <= not((layer0_outputs(1556)) or (layer0_outputs(5457)));
    layer1_outputs(5125) <= layer0_outputs(8108);
    layer1_outputs(5126) <= not(layer0_outputs(7166));
    layer1_outputs(5127) <= not(layer0_outputs(6048));
    layer1_outputs(5128) <= (layer0_outputs(1774)) xor (layer0_outputs(1697));
    layer1_outputs(5129) <= not(layer0_outputs(6282)) or (layer0_outputs(2931));
    layer1_outputs(5130) <= not((layer0_outputs(6267)) or (layer0_outputs(8670)));
    layer1_outputs(5131) <= not((layer0_outputs(4552)) or (layer0_outputs(7700)));
    layer1_outputs(5132) <= not((layer0_outputs(2491)) and (layer0_outputs(6953)));
    layer1_outputs(5133) <= not(layer0_outputs(4893)) or (layer0_outputs(6751));
    layer1_outputs(5134) <= not(layer0_outputs(5291));
    layer1_outputs(5135) <= layer0_outputs(5964);
    layer1_outputs(5136) <= not((layer0_outputs(2374)) or (layer0_outputs(4688)));
    layer1_outputs(5137) <= layer0_outputs(3261);
    layer1_outputs(5138) <= (layer0_outputs(9391)) and not (layer0_outputs(9486));
    layer1_outputs(5139) <= not(layer0_outputs(9592));
    layer1_outputs(5140) <= layer0_outputs(9482);
    layer1_outputs(5141) <= '0';
    layer1_outputs(5142) <= not(layer0_outputs(5820));
    layer1_outputs(5143) <= layer0_outputs(7501);
    layer1_outputs(5144) <= not(layer0_outputs(3535));
    layer1_outputs(5145) <= not((layer0_outputs(1719)) and (layer0_outputs(234)));
    layer1_outputs(5146) <= (layer0_outputs(6384)) and not (layer0_outputs(4115));
    layer1_outputs(5147) <= (layer0_outputs(6432)) and not (layer0_outputs(4279));
    layer1_outputs(5148) <= not(layer0_outputs(6574));
    layer1_outputs(5149) <= not(layer0_outputs(6425));
    layer1_outputs(5150) <= (layer0_outputs(5139)) and (layer0_outputs(8788));
    layer1_outputs(5151) <= layer0_outputs(4524);
    layer1_outputs(5152) <= not((layer0_outputs(1182)) and (layer0_outputs(5445)));
    layer1_outputs(5153) <= not((layer0_outputs(6903)) xor (layer0_outputs(455)));
    layer1_outputs(5154) <= not(layer0_outputs(2892));
    layer1_outputs(5155) <= not((layer0_outputs(8138)) or (layer0_outputs(4356)));
    layer1_outputs(5156) <= layer0_outputs(1540);
    layer1_outputs(5157) <= not(layer0_outputs(3018));
    layer1_outputs(5158) <= (layer0_outputs(7829)) or (layer0_outputs(3724));
    layer1_outputs(5159) <= layer0_outputs(9300);
    layer1_outputs(5160) <= layer0_outputs(4932);
    layer1_outputs(5161) <= not(layer0_outputs(51)) or (layer0_outputs(7445));
    layer1_outputs(5162) <= not(layer0_outputs(2434)) or (layer0_outputs(2222));
    layer1_outputs(5163) <= not(layer0_outputs(5439));
    layer1_outputs(5164) <= not((layer0_outputs(6097)) and (layer0_outputs(6723)));
    layer1_outputs(5165) <= layer0_outputs(7166);
    layer1_outputs(5166) <= (layer0_outputs(573)) and not (layer0_outputs(890));
    layer1_outputs(5167) <= (layer0_outputs(2464)) or (layer0_outputs(1594));
    layer1_outputs(5168) <= layer0_outputs(8772);
    layer1_outputs(5169) <= layer0_outputs(5657);
    layer1_outputs(5170) <= not(layer0_outputs(4183));
    layer1_outputs(5171) <= (layer0_outputs(6177)) and (layer0_outputs(8684));
    layer1_outputs(5172) <= not(layer0_outputs(9038)) or (layer0_outputs(9641));
    layer1_outputs(5173) <= layer0_outputs(7336);
    layer1_outputs(5174) <= not(layer0_outputs(398));
    layer1_outputs(5175) <= '1';
    layer1_outputs(5176) <= not(layer0_outputs(3074));
    layer1_outputs(5177) <= not(layer0_outputs(2199)) or (layer0_outputs(746));
    layer1_outputs(5178) <= (layer0_outputs(2414)) or (layer0_outputs(5532));
    layer1_outputs(5179) <= not(layer0_outputs(2255));
    layer1_outputs(5180) <= not(layer0_outputs(3781));
    layer1_outputs(5181) <= not(layer0_outputs(4936)) or (layer0_outputs(4557));
    layer1_outputs(5182) <= not((layer0_outputs(8520)) and (layer0_outputs(392)));
    layer1_outputs(5183) <= not(layer0_outputs(7706));
    layer1_outputs(5184) <= '1';
    layer1_outputs(5185) <= '1';
    layer1_outputs(5186) <= not(layer0_outputs(2999));
    layer1_outputs(5187) <= (layer0_outputs(3432)) and not (layer0_outputs(8898));
    layer1_outputs(5188) <= (layer0_outputs(8341)) and not (layer0_outputs(10095));
    layer1_outputs(5189) <= not((layer0_outputs(8301)) or (layer0_outputs(7267)));
    layer1_outputs(5190) <= not(layer0_outputs(7476)) or (layer0_outputs(2129));
    layer1_outputs(5191) <= not((layer0_outputs(6370)) or (layer0_outputs(5307)));
    layer1_outputs(5192) <= (layer0_outputs(5352)) and not (layer0_outputs(2194));
    layer1_outputs(5193) <= (layer0_outputs(3119)) and not (layer0_outputs(2950));
    layer1_outputs(5194) <= not(layer0_outputs(4916));
    layer1_outputs(5195) <= layer0_outputs(8863);
    layer1_outputs(5196) <= layer0_outputs(9046);
    layer1_outputs(5197) <= not(layer0_outputs(4094)) or (layer0_outputs(6776));
    layer1_outputs(5198) <= not(layer0_outputs(7959));
    layer1_outputs(5199) <= not((layer0_outputs(686)) and (layer0_outputs(5662)));
    layer1_outputs(5200) <= (layer0_outputs(9411)) or (layer0_outputs(6675));
    layer1_outputs(5201) <= (layer0_outputs(2379)) or (layer0_outputs(9659));
    layer1_outputs(5202) <= not(layer0_outputs(1621)) or (layer0_outputs(6788));
    layer1_outputs(5203) <= not(layer0_outputs(6221));
    layer1_outputs(5204) <= (layer0_outputs(530)) and not (layer0_outputs(2668));
    layer1_outputs(5205) <= layer0_outputs(2107);
    layer1_outputs(5206) <= not(layer0_outputs(27)) or (layer0_outputs(2072));
    layer1_outputs(5207) <= not((layer0_outputs(333)) and (layer0_outputs(9773)));
    layer1_outputs(5208) <= not(layer0_outputs(116)) or (layer0_outputs(9409));
    layer1_outputs(5209) <= layer0_outputs(8811);
    layer1_outputs(5210) <= '0';
    layer1_outputs(5211) <= not((layer0_outputs(9923)) and (layer0_outputs(6349)));
    layer1_outputs(5212) <= (layer0_outputs(6665)) or (layer0_outputs(10219));
    layer1_outputs(5213) <= (layer0_outputs(2478)) and not (layer0_outputs(817));
    layer1_outputs(5214) <= (layer0_outputs(7316)) and not (layer0_outputs(8939));
    layer1_outputs(5215) <= (layer0_outputs(7759)) and not (layer0_outputs(3524));
    layer1_outputs(5216) <= '1';
    layer1_outputs(5217) <= (layer0_outputs(1617)) and (layer0_outputs(6383));
    layer1_outputs(5218) <= (layer0_outputs(5020)) or (layer0_outputs(2642));
    layer1_outputs(5219) <= layer0_outputs(9071);
    layer1_outputs(5220) <= not(layer0_outputs(3655));
    layer1_outputs(5221) <= layer0_outputs(9003);
    layer1_outputs(5222) <= not(layer0_outputs(9770));
    layer1_outputs(5223) <= not(layer0_outputs(6137));
    layer1_outputs(5224) <= (layer0_outputs(4278)) and not (layer0_outputs(950));
    layer1_outputs(5225) <= not(layer0_outputs(4216));
    layer1_outputs(5226) <= layer0_outputs(1504);
    layer1_outputs(5227) <= not((layer0_outputs(9363)) and (layer0_outputs(144)));
    layer1_outputs(5228) <= not(layer0_outputs(9245)) or (layer0_outputs(5076));
    layer1_outputs(5229) <= not(layer0_outputs(8373)) or (layer0_outputs(187));
    layer1_outputs(5230) <= (layer0_outputs(54)) or (layer0_outputs(3812));
    layer1_outputs(5231) <= (layer0_outputs(6900)) and not (layer0_outputs(723));
    layer1_outputs(5232) <= not((layer0_outputs(9908)) or (layer0_outputs(2669)));
    layer1_outputs(5233) <= (layer0_outputs(3865)) or (layer0_outputs(5898));
    layer1_outputs(5234) <= (layer0_outputs(4479)) or (layer0_outputs(9263));
    layer1_outputs(5235) <= (layer0_outputs(413)) or (layer0_outputs(9360));
    layer1_outputs(5236) <= layer0_outputs(1381);
    layer1_outputs(5237) <= layer0_outputs(6299);
    layer1_outputs(5238) <= not(layer0_outputs(7470));
    layer1_outputs(5239) <= (layer0_outputs(3777)) and not (layer0_outputs(199));
    layer1_outputs(5240) <= not(layer0_outputs(9630)) or (layer0_outputs(5380));
    layer1_outputs(5241) <= layer0_outputs(793);
    layer1_outputs(5242) <= (layer0_outputs(6728)) or (layer0_outputs(2742));
    layer1_outputs(5243) <= '0';
    layer1_outputs(5244) <= not(layer0_outputs(3801));
    layer1_outputs(5245) <= (layer0_outputs(5269)) and (layer0_outputs(10059));
    layer1_outputs(5246) <= not((layer0_outputs(6742)) xor (layer0_outputs(4207)));
    layer1_outputs(5247) <= (layer0_outputs(3422)) or (layer0_outputs(5904));
    layer1_outputs(5248) <= (layer0_outputs(6841)) or (layer0_outputs(7135));
    layer1_outputs(5249) <= layer0_outputs(2557);
    layer1_outputs(5250) <= (layer0_outputs(6561)) and not (layer0_outputs(1568));
    layer1_outputs(5251) <= (layer0_outputs(4514)) and not (layer0_outputs(8107));
    layer1_outputs(5252) <= not(layer0_outputs(7733)) or (layer0_outputs(1544));
    layer1_outputs(5253) <= (layer0_outputs(7608)) or (layer0_outputs(7407));
    layer1_outputs(5254) <= not((layer0_outputs(3606)) xor (layer0_outputs(7244)));
    layer1_outputs(5255) <= layer0_outputs(128);
    layer1_outputs(5256) <= layer0_outputs(9740);
    layer1_outputs(5257) <= not(layer0_outputs(1884));
    layer1_outputs(5258) <= not((layer0_outputs(7913)) or (layer0_outputs(9558)));
    layer1_outputs(5259) <= (layer0_outputs(4475)) and not (layer0_outputs(792));
    layer1_outputs(5260) <= (layer0_outputs(9968)) and not (layer0_outputs(4069));
    layer1_outputs(5261) <= '0';
    layer1_outputs(5262) <= not((layer0_outputs(5793)) xor (layer0_outputs(4716)));
    layer1_outputs(5263) <= (layer0_outputs(8075)) xor (layer0_outputs(2524));
    layer1_outputs(5264) <= (layer0_outputs(3504)) xor (layer0_outputs(2385));
    layer1_outputs(5265) <= not((layer0_outputs(4026)) and (layer0_outputs(2556)));
    layer1_outputs(5266) <= not((layer0_outputs(1953)) and (layer0_outputs(9851)));
    layer1_outputs(5267) <= '0';
    layer1_outputs(5268) <= (layer0_outputs(7799)) xor (layer0_outputs(6026));
    layer1_outputs(5269) <= (layer0_outputs(2902)) and not (layer0_outputs(6313));
    layer1_outputs(5270) <= layer0_outputs(1543);
    layer1_outputs(5271) <= (layer0_outputs(3569)) and (layer0_outputs(6123));
    layer1_outputs(5272) <= layer0_outputs(4335);
    layer1_outputs(5273) <= not(layer0_outputs(4591)) or (layer0_outputs(8212));
    layer1_outputs(5274) <= not((layer0_outputs(8608)) or (layer0_outputs(8454)));
    layer1_outputs(5275) <= not(layer0_outputs(9662));
    layer1_outputs(5276) <= (layer0_outputs(3152)) and (layer0_outputs(1500));
    layer1_outputs(5277) <= not(layer0_outputs(5859)) or (layer0_outputs(1660));
    layer1_outputs(5278) <= '0';
    layer1_outputs(5279) <= not(layer0_outputs(3939)) or (layer0_outputs(8966));
    layer1_outputs(5280) <= not((layer0_outputs(2575)) or (layer0_outputs(8913)));
    layer1_outputs(5281) <= layer0_outputs(4455);
    layer1_outputs(5282) <= (layer0_outputs(3701)) and not (layer0_outputs(7036));
    layer1_outputs(5283) <= '0';
    layer1_outputs(5284) <= layer0_outputs(1469);
    layer1_outputs(5285) <= not((layer0_outputs(1651)) xor (layer0_outputs(1213)));
    layer1_outputs(5286) <= not(layer0_outputs(150));
    layer1_outputs(5287) <= not(layer0_outputs(10112)) or (layer0_outputs(1470));
    layer1_outputs(5288) <= (layer0_outputs(7406)) and (layer0_outputs(47));
    layer1_outputs(5289) <= (layer0_outputs(1606)) and not (layer0_outputs(10108));
    layer1_outputs(5290) <= not(layer0_outputs(7919));
    layer1_outputs(5291) <= (layer0_outputs(5006)) and not (layer0_outputs(141));
    layer1_outputs(5292) <= '1';
    layer1_outputs(5293) <= (layer0_outputs(1792)) xor (layer0_outputs(1594));
    layer1_outputs(5294) <= layer0_outputs(2873);
    layer1_outputs(5295) <= (layer0_outputs(4705)) and not (layer0_outputs(6089));
    layer1_outputs(5296) <= not(layer0_outputs(6068));
    layer1_outputs(5297) <= (layer0_outputs(4396)) or (layer0_outputs(6910));
    layer1_outputs(5298) <= not(layer0_outputs(7508));
    layer1_outputs(5299) <= layer0_outputs(9840);
    layer1_outputs(5300) <= not((layer0_outputs(9782)) and (layer0_outputs(7852)));
    layer1_outputs(5301) <= (layer0_outputs(3562)) and (layer0_outputs(5225));
    layer1_outputs(5302) <= (layer0_outputs(8838)) and not (layer0_outputs(1012));
    layer1_outputs(5303) <= not((layer0_outputs(7767)) xor (layer0_outputs(5492)));
    layer1_outputs(5304) <= not((layer0_outputs(3231)) or (layer0_outputs(4785)));
    layer1_outputs(5305) <= (layer0_outputs(6933)) or (layer0_outputs(8235));
    layer1_outputs(5306) <= not((layer0_outputs(6979)) and (layer0_outputs(6348)));
    layer1_outputs(5307) <= (layer0_outputs(3021)) and (layer0_outputs(7541));
    layer1_outputs(5308) <= (layer0_outputs(9226)) and not (layer0_outputs(3169));
    layer1_outputs(5309) <= (layer0_outputs(6996)) xor (layer0_outputs(2598));
    layer1_outputs(5310) <= not((layer0_outputs(359)) xor (layer0_outputs(4774)));
    layer1_outputs(5311) <= not((layer0_outputs(204)) xor (layer0_outputs(5756)));
    layer1_outputs(5312) <= layer0_outputs(7743);
    layer1_outputs(5313) <= not((layer0_outputs(6596)) and (layer0_outputs(5312)));
    layer1_outputs(5314) <= (layer0_outputs(5645)) and not (layer0_outputs(9220));
    layer1_outputs(5315) <= (layer0_outputs(9152)) xor (layer0_outputs(2959));
    layer1_outputs(5316) <= (layer0_outputs(2412)) and (layer0_outputs(48));
    layer1_outputs(5317) <= not(layer0_outputs(4480));
    layer1_outputs(5318) <= layer0_outputs(9932);
    layer1_outputs(5319) <= '1';
    layer1_outputs(5320) <= not((layer0_outputs(451)) xor (layer0_outputs(8591)));
    layer1_outputs(5321) <= (layer0_outputs(9635)) and not (layer0_outputs(7684));
    layer1_outputs(5322) <= layer0_outputs(3595);
    layer1_outputs(5323) <= not((layer0_outputs(1147)) or (layer0_outputs(7903)));
    layer1_outputs(5324) <= not((layer0_outputs(6863)) or (layer0_outputs(2921)));
    layer1_outputs(5325) <= (layer0_outputs(1724)) or (layer0_outputs(1447));
    layer1_outputs(5326) <= not((layer0_outputs(7747)) and (layer0_outputs(9796)));
    layer1_outputs(5327) <= not(layer0_outputs(6872));
    layer1_outputs(5328) <= not(layer0_outputs(8478)) or (layer0_outputs(4841));
    layer1_outputs(5329) <= (layer0_outputs(2180)) or (layer0_outputs(3371));
    layer1_outputs(5330) <= layer0_outputs(7315);
    layer1_outputs(5331) <= '1';
    layer1_outputs(5332) <= not((layer0_outputs(8575)) or (layer0_outputs(5075)));
    layer1_outputs(5333) <= not(layer0_outputs(5198));
    layer1_outputs(5334) <= not(layer0_outputs(2183)) or (layer0_outputs(7916));
    layer1_outputs(5335) <= layer0_outputs(1592);
    layer1_outputs(5336) <= not(layer0_outputs(9098));
    layer1_outputs(5337) <= '1';
    layer1_outputs(5338) <= (layer0_outputs(9865)) and (layer0_outputs(3635));
    layer1_outputs(5339) <= '1';
    layer1_outputs(5340) <= not(layer0_outputs(1661)) or (layer0_outputs(5154));
    layer1_outputs(5341) <= not((layer0_outputs(5268)) and (layer0_outputs(2062)));
    layer1_outputs(5342) <= not((layer0_outputs(9581)) and (layer0_outputs(7337)));
    layer1_outputs(5343) <= not((layer0_outputs(7347)) or (layer0_outputs(166)));
    layer1_outputs(5344) <= not((layer0_outputs(5096)) and (layer0_outputs(9427)));
    layer1_outputs(5345) <= '0';
    layer1_outputs(5346) <= not(layer0_outputs(5483));
    layer1_outputs(5347) <= layer0_outputs(7646);
    layer1_outputs(5348) <= layer0_outputs(4682);
    layer1_outputs(5349) <= layer0_outputs(1717);
    layer1_outputs(5350) <= '1';
    layer1_outputs(5351) <= (layer0_outputs(4453)) and not (layer0_outputs(6406));
    layer1_outputs(5352) <= '1';
    layer1_outputs(5353) <= not((layer0_outputs(6085)) or (layer0_outputs(5476)));
    layer1_outputs(5354) <= not(layer0_outputs(2051)) or (layer0_outputs(10120));
    layer1_outputs(5355) <= not((layer0_outputs(6224)) or (layer0_outputs(279)));
    layer1_outputs(5356) <= not(layer0_outputs(232)) or (layer0_outputs(321));
    layer1_outputs(5357) <= not((layer0_outputs(3386)) or (layer0_outputs(1406)));
    layer1_outputs(5358) <= not((layer0_outputs(4759)) xor (layer0_outputs(2877)));
    layer1_outputs(5359) <= (layer0_outputs(2367)) xor (layer0_outputs(7979));
    layer1_outputs(5360) <= not(layer0_outputs(4976)) or (layer0_outputs(8832));
    layer1_outputs(5361) <= (layer0_outputs(6586)) and not (layer0_outputs(1761));
    layer1_outputs(5362) <= not(layer0_outputs(5583)) or (layer0_outputs(8783));
    layer1_outputs(5363) <= layer0_outputs(5062);
    layer1_outputs(5364) <= not(layer0_outputs(9455)) or (layer0_outputs(1271));
    layer1_outputs(5365) <= not(layer0_outputs(6550));
    layer1_outputs(5366) <= layer0_outputs(1725);
    layer1_outputs(5367) <= not(layer0_outputs(7402));
    layer1_outputs(5368) <= not((layer0_outputs(534)) or (layer0_outputs(8394)));
    layer1_outputs(5369) <= not(layer0_outputs(6826));
    layer1_outputs(5370) <= (layer0_outputs(4400)) and (layer0_outputs(2683));
    layer1_outputs(5371) <= layer0_outputs(7362);
    layer1_outputs(5372) <= not((layer0_outputs(1755)) and (layer0_outputs(9145)));
    layer1_outputs(5373) <= (layer0_outputs(906)) and (layer0_outputs(5788));
    layer1_outputs(5374) <= (layer0_outputs(79)) and not (layer0_outputs(2967));
    layer1_outputs(5375) <= (layer0_outputs(6514)) and not (layer0_outputs(3679));
    layer1_outputs(5376) <= not((layer0_outputs(1411)) or (layer0_outputs(3308)));
    layer1_outputs(5377) <= layer0_outputs(8484);
    layer1_outputs(5378) <= (layer0_outputs(9387)) xor (layer0_outputs(1507));
    layer1_outputs(5379) <= layer0_outputs(256);
    layer1_outputs(5380) <= not(layer0_outputs(7817)) or (layer0_outputs(2378));
    layer1_outputs(5381) <= '0';
    layer1_outputs(5382) <= not(layer0_outputs(7823)) or (layer0_outputs(7392));
    layer1_outputs(5383) <= not(layer0_outputs(4156)) or (layer0_outputs(2769));
    layer1_outputs(5384) <= not(layer0_outputs(8463));
    layer1_outputs(5385) <= '1';
    layer1_outputs(5386) <= not(layer0_outputs(2628)) or (layer0_outputs(3351));
    layer1_outputs(5387) <= (layer0_outputs(3302)) or (layer0_outputs(8376));
    layer1_outputs(5388) <= not(layer0_outputs(9811));
    layer1_outputs(5389) <= not(layer0_outputs(2031));
    layer1_outputs(5390) <= layer0_outputs(9789);
    layer1_outputs(5391) <= not((layer0_outputs(6509)) and (layer0_outputs(3612)));
    layer1_outputs(5392) <= not((layer0_outputs(2209)) xor (layer0_outputs(2889)));
    layer1_outputs(5393) <= not((layer0_outputs(2695)) and (layer0_outputs(7159)));
    layer1_outputs(5394) <= layer0_outputs(4049);
    layer1_outputs(5395) <= not(layer0_outputs(5156));
    layer1_outputs(5396) <= (layer0_outputs(3384)) and not (layer0_outputs(5552));
    layer1_outputs(5397) <= not(layer0_outputs(2959)) or (layer0_outputs(1779));
    layer1_outputs(5398) <= not((layer0_outputs(1189)) xor (layer0_outputs(3144)));
    layer1_outputs(5399) <= '0';
    layer1_outputs(5400) <= not(layer0_outputs(2260)) or (layer0_outputs(6174));
    layer1_outputs(5401) <= not((layer0_outputs(8785)) xor (layer0_outputs(4631)));
    layer1_outputs(5402) <= not((layer0_outputs(8564)) or (layer0_outputs(3707)));
    layer1_outputs(5403) <= not(layer0_outputs(4823));
    layer1_outputs(5404) <= (layer0_outputs(5834)) and (layer0_outputs(5453));
    layer1_outputs(5405) <= not(layer0_outputs(758));
    layer1_outputs(5406) <= (layer0_outputs(3579)) and (layer0_outputs(3643));
    layer1_outputs(5407) <= not((layer0_outputs(7238)) and (layer0_outputs(6907)));
    layer1_outputs(5408) <= not((layer0_outputs(8340)) and (layer0_outputs(5541)));
    layer1_outputs(5409) <= not((layer0_outputs(3705)) xor (layer0_outputs(3414)));
    layer1_outputs(5410) <= (layer0_outputs(2455)) and not (layer0_outputs(5262));
    layer1_outputs(5411) <= not(layer0_outputs(7656));
    layer1_outputs(5412) <= (layer0_outputs(5122)) and (layer0_outputs(3730));
    layer1_outputs(5413) <= (layer0_outputs(1657)) and not (layer0_outputs(6941));
    layer1_outputs(5414) <= not(layer0_outputs(5130));
    layer1_outputs(5415) <= layer0_outputs(6582);
    layer1_outputs(5416) <= not((layer0_outputs(3566)) or (layer0_outputs(2671)));
    layer1_outputs(5417) <= (layer0_outputs(4289)) and not (layer0_outputs(4312));
    layer1_outputs(5418) <= not((layer0_outputs(2850)) and (layer0_outputs(3007)));
    layer1_outputs(5419) <= not(layer0_outputs(1744)) or (layer0_outputs(8569));
    layer1_outputs(5420) <= layer0_outputs(8693);
    layer1_outputs(5421) <= not((layer0_outputs(6760)) and (layer0_outputs(1238)));
    layer1_outputs(5422) <= (layer0_outputs(7027)) and (layer0_outputs(2105));
    layer1_outputs(5423) <= layer0_outputs(3350);
    layer1_outputs(5424) <= (layer0_outputs(10027)) or (layer0_outputs(3388));
    layer1_outputs(5425) <= not(layer0_outputs(703));
    layer1_outputs(5426) <= not(layer0_outputs(6122)) or (layer0_outputs(5831));
    layer1_outputs(5427) <= '1';
    layer1_outputs(5428) <= layer0_outputs(9738);
    layer1_outputs(5429) <= layer0_outputs(6470);
    layer1_outputs(5430) <= (layer0_outputs(5965)) and (layer0_outputs(5201));
    layer1_outputs(5431) <= not(layer0_outputs(1059));
    layer1_outputs(5432) <= (layer0_outputs(2124)) xor (layer0_outputs(6510));
    layer1_outputs(5433) <= (layer0_outputs(9357)) and (layer0_outputs(10196));
    layer1_outputs(5434) <= (layer0_outputs(3297)) or (layer0_outputs(1020));
    layer1_outputs(5435) <= layer0_outputs(9640);
    layer1_outputs(5436) <= (layer0_outputs(9693)) and (layer0_outputs(8082));
    layer1_outputs(5437) <= not(layer0_outputs(963)) or (layer0_outputs(8671));
    layer1_outputs(5438) <= '1';
    layer1_outputs(5439) <= not((layer0_outputs(1810)) and (layer0_outputs(1606)));
    layer1_outputs(5440) <= not(layer0_outputs(4767));
    layer1_outputs(5441) <= layer0_outputs(4355);
    layer1_outputs(5442) <= not((layer0_outputs(2397)) and (layer0_outputs(2905)));
    layer1_outputs(5443) <= (layer0_outputs(3597)) or (layer0_outputs(9224));
    layer1_outputs(5444) <= '0';
    layer1_outputs(5445) <= layer0_outputs(3209);
    layer1_outputs(5446) <= layer0_outputs(3137);
    layer1_outputs(5447) <= not(layer0_outputs(2712)) or (layer0_outputs(3236));
    layer1_outputs(5448) <= not(layer0_outputs(6297)) or (layer0_outputs(2137));
    layer1_outputs(5449) <= (layer0_outputs(1195)) and not (layer0_outputs(7426));
    layer1_outputs(5450) <= '0';
    layer1_outputs(5451) <= (layer0_outputs(5209)) or (layer0_outputs(6625));
    layer1_outputs(5452) <= (layer0_outputs(2384)) and not (layer0_outputs(9285));
    layer1_outputs(5453) <= not(layer0_outputs(9304));
    layer1_outputs(5454) <= layer0_outputs(2765);
    layer1_outputs(5455) <= not((layer0_outputs(5766)) or (layer0_outputs(1468)));
    layer1_outputs(5456) <= (layer0_outputs(5276)) and (layer0_outputs(9066));
    layer1_outputs(5457) <= (layer0_outputs(8470)) and not (layer0_outputs(6130));
    layer1_outputs(5458) <= not((layer0_outputs(5327)) or (layer0_outputs(5169)));
    layer1_outputs(5459) <= layer0_outputs(6531);
    layer1_outputs(5460) <= layer0_outputs(6713);
    layer1_outputs(5461) <= not(layer0_outputs(9619)) or (layer0_outputs(7875));
    layer1_outputs(5462) <= not((layer0_outputs(4736)) or (layer0_outputs(2376)));
    layer1_outputs(5463) <= not((layer0_outputs(8744)) or (layer0_outputs(9582)));
    layer1_outputs(5464) <= not(layer0_outputs(7048));
    layer1_outputs(5465) <= '1';
    layer1_outputs(5466) <= (layer0_outputs(6670)) xor (layer0_outputs(4567));
    layer1_outputs(5467) <= layer0_outputs(5865);
    layer1_outputs(5468) <= not(layer0_outputs(9689));
    layer1_outputs(5469) <= not(layer0_outputs(8147)) or (layer0_outputs(2807));
    layer1_outputs(5470) <= '1';
    layer1_outputs(5471) <= not((layer0_outputs(1708)) or (layer0_outputs(8881)));
    layer1_outputs(5472) <= not(layer0_outputs(6572)) or (layer0_outputs(938));
    layer1_outputs(5473) <= not(layer0_outputs(7573)) or (layer0_outputs(9463));
    layer1_outputs(5474) <= (layer0_outputs(554)) or (layer0_outputs(2930));
    layer1_outputs(5475) <= not((layer0_outputs(5360)) xor (layer0_outputs(3402)));
    layer1_outputs(5476) <= (layer0_outputs(5792)) and (layer0_outputs(2893));
    layer1_outputs(5477) <= (layer0_outputs(5622)) and not (layer0_outputs(1862));
    layer1_outputs(5478) <= layer0_outputs(1519);
    layer1_outputs(5479) <= layer0_outputs(710);
    layer1_outputs(5480) <= not((layer0_outputs(6656)) and (layer0_outputs(4460)));
    layer1_outputs(5481) <= (layer0_outputs(2020)) xor (layer0_outputs(1386));
    layer1_outputs(5482) <= (layer0_outputs(1172)) and not (layer0_outputs(5953));
    layer1_outputs(5483) <= (layer0_outputs(4757)) or (layer0_outputs(6377));
    layer1_outputs(5484) <= (layer0_outputs(617)) and not (layer0_outputs(6179));
    layer1_outputs(5485) <= not(layer0_outputs(8105)) or (layer0_outputs(10062));
    layer1_outputs(5486) <= '0';
    layer1_outputs(5487) <= (layer0_outputs(6264)) and not (layer0_outputs(7052));
    layer1_outputs(5488) <= (layer0_outputs(9325)) or (layer0_outputs(5574));
    layer1_outputs(5489) <= (layer0_outputs(7557)) and not (layer0_outputs(1147));
    layer1_outputs(5490) <= (layer0_outputs(440)) xor (layer0_outputs(8835));
    layer1_outputs(5491) <= not(layer0_outputs(1046)) or (layer0_outputs(9484));
    layer1_outputs(5492) <= layer0_outputs(9335);
    layer1_outputs(5493) <= layer0_outputs(7066);
    layer1_outputs(5494) <= not(layer0_outputs(7155));
    layer1_outputs(5495) <= '0';
    layer1_outputs(5496) <= layer0_outputs(3036);
    layer1_outputs(5497) <= (layer0_outputs(187)) and not (layer0_outputs(7662));
    layer1_outputs(5498) <= layer0_outputs(4014);
    layer1_outputs(5499) <= (layer0_outputs(3832)) and not (layer0_outputs(2114));
    layer1_outputs(5500) <= not(layer0_outputs(9060));
    layer1_outputs(5501) <= not(layer0_outputs(983));
    layer1_outputs(5502) <= '1';
    layer1_outputs(5503) <= (layer0_outputs(7590)) and not (layer0_outputs(6899));
    layer1_outputs(5504) <= not(layer0_outputs(5053)) or (layer0_outputs(3326));
    layer1_outputs(5505) <= not((layer0_outputs(4596)) and (layer0_outputs(2551)));
    layer1_outputs(5506) <= (layer0_outputs(8481)) xor (layer0_outputs(10207));
    layer1_outputs(5507) <= not(layer0_outputs(3094)) or (layer0_outputs(9789));
    layer1_outputs(5508) <= (layer0_outputs(6416)) or (layer0_outputs(635));
    layer1_outputs(5509) <= not((layer0_outputs(8638)) and (layer0_outputs(372)));
    layer1_outputs(5510) <= (layer0_outputs(4857)) and not (layer0_outputs(410));
    layer1_outputs(5511) <= not(layer0_outputs(9774)) or (layer0_outputs(5200));
    layer1_outputs(5512) <= layer0_outputs(577);
    layer1_outputs(5513) <= layer0_outputs(7406);
    layer1_outputs(5514) <= layer0_outputs(4365);
    layer1_outputs(5515) <= (layer0_outputs(5578)) and (layer0_outputs(6189));
    layer1_outputs(5516) <= '1';
    layer1_outputs(5517) <= (layer0_outputs(4202)) and not (layer0_outputs(801));
    layer1_outputs(5518) <= not(layer0_outputs(8748)) or (layer0_outputs(5079));
    layer1_outputs(5519) <= not(layer0_outputs(1156)) or (layer0_outputs(2267));
    layer1_outputs(5520) <= (layer0_outputs(4234)) and not (layer0_outputs(7591));
    layer1_outputs(5521) <= (layer0_outputs(1823)) and not (layer0_outputs(4088));
    layer1_outputs(5522) <= (layer0_outputs(225)) or (layer0_outputs(4794));
    layer1_outputs(5523) <= (layer0_outputs(7118)) and not (layer0_outputs(2543));
    layer1_outputs(5524) <= (layer0_outputs(7332)) and (layer0_outputs(6164));
    layer1_outputs(5525) <= not((layer0_outputs(1415)) or (layer0_outputs(7431)));
    layer1_outputs(5526) <= not(layer0_outputs(5415));
    layer1_outputs(5527) <= not(layer0_outputs(237)) or (layer0_outputs(8070));
    layer1_outputs(5528) <= not(layer0_outputs(2272)) or (layer0_outputs(3051));
    layer1_outputs(5529) <= not((layer0_outputs(8272)) and (layer0_outputs(9410)));
    layer1_outputs(5530) <= (layer0_outputs(5473)) or (layer0_outputs(9762));
    layer1_outputs(5531) <= '1';
    layer1_outputs(5532) <= '0';
    layer1_outputs(5533) <= not(layer0_outputs(8315)) or (layer0_outputs(3082));
    layer1_outputs(5534) <= not(layer0_outputs(4037));
    layer1_outputs(5535) <= '1';
    layer1_outputs(5536) <= not(layer0_outputs(2171));
    layer1_outputs(5537) <= layer0_outputs(3995);
    layer1_outputs(5538) <= not(layer0_outputs(226)) or (layer0_outputs(8436));
    layer1_outputs(5539) <= not(layer0_outputs(7907));
    layer1_outputs(5540) <= '0';
    layer1_outputs(5541) <= (layer0_outputs(4877)) and not (layer0_outputs(58));
    layer1_outputs(5542) <= (layer0_outputs(4550)) and not (layer0_outputs(8616));
    layer1_outputs(5543) <= not(layer0_outputs(7900));
    layer1_outputs(5544) <= not((layer0_outputs(9744)) and (layer0_outputs(1426)));
    layer1_outputs(5545) <= '1';
    layer1_outputs(5546) <= layer0_outputs(2609);
    layer1_outputs(5547) <= (layer0_outputs(654)) xor (layer0_outputs(2471));
    layer1_outputs(5548) <= not(layer0_outputs(6094));
    layer1_outputs(5549) <= (layer0_outputs(5264)) and not (layer0_outputs(7418));
    layer1_outputs(5550) <= (layer0_outputs(4413)) or (layer0_outputs(5095));
    layer1_outputs(5551) <= layer0_outputs(9662);
    layer1_outputs(5552) <= (layer0_outputs(8734)) or (layer0_outputs(3809));
    layer1_outputs(5553) <= not((layer0_outputs(7518)) xor (layer0_outputs(9234)));
    layer1_outputs(5554) <= (layer0_outputs(6436)) and (layer0_outputs(4913));
    layer1_outputs(5555) <= (layer0_outputs(1197)) and (layer0_outputs(6962));
    layer1_outputs(5556) <= (layer0_outputs(5771)) or (layer0_outputs(4492));
    layer1_outputs(5557) <= (layer0_outputs(4882)) xor (layer0_outputs(7669));
    layer1_outputs(5558) <= (layer0_outputs(1957)) and (layer0_outputs(1943));
    layer1_outputs(5559) <= (layer0_outputs(6920)) and not (layer0_outputs(756));
    layer1_outputs(5560) <= not((layer0_outputs(2801)) and (layer0_outputs(2661)));
    layer1_outputs(5561) <= (layer0_outputs(9237)) and not (layer0_outputs(2638));
    layer1_outputs(5562) <= not(layer0_outputs(8375));
    layer1_outputs(5563) <= not((layer0_outputs(8110)) or (layer0_outputs(457)));
    layer1_outputs(5564) <= layer0_outputs(4729);
    layer1_outputs(5565) <= (layer0_outputs(4310)) or (layer0_outputs(7984));
    layer1_outputs(5566) <= not(layer0_outputs(7808));
    layer1_outputs(5567) <= '0';
    layer1_outputs(5568) <= (layer0_outputs(3372)) and (layer0_outputs(7317));
    layer1_outputs(5569) <= not(layer0_outputs(8597));
    layer1_outputs(5570) <= not(layer0_outputs(7101));
    layer1_outputs(5571) <= '1';
    layer1_outputs(5572) <= (layer0_outputs(6911)) xor (layer0_outputs(7046));
    layer1_outputs(5573) <= layer0_outputs(1517);
    layer1_outputs(5574) <= layer0_outputs(8878);
    layer1_outputs(5575) <= not(layer0_outputs(2213));
    layer1_outputs(5576) <= '0';
    layer1_outputs(5577) <= (layer0_outputs(310)) xor (layer0_outputs(549));
    layer1_outputs(5578) <= not(layer0_outputs(2406));
    layer1_outputs(5579) <= '0';
    layer1_outputs(5580) <= layer0_outputs(8334);
    layer1_outputs(5581) <= not(layer0_outputs(9803));
    layer1_outputs(5582) <= not(layer0_outputs(5057));
    layer1_outputs(5583) <= not(layer0_outputs(3929));
    layer1_outputs(5584) <= (layer0_outputs(7374)) and not (layer0_outputs(8545));
    layer1_outputs(5585) <= (layer0_outputs(6556)) xor (layer0_outputs(2978));
    layer1_outputs(5586) <= '1';
    layer1_outputs(5587) <= '1';
    layer1_outputs(5588) <= (layer0_outputs(5683)) and not (layer0_outputs(6439));
    layer1_outputs(5589) <= not(layer0_outputs(8325)) or (layer0_outputs(5855));
    layer1_outputs(5590) <= (layer0_outputs(5084)) or (layer0_outputs(9540));
    layer1_outputs(5591) <= '0';
    layer1_outputs(5592) <= (layer0_outputs(715)) and not (layer0_outputs(2567));
    layer1_outputs(5593) <= (layer0_outputs(9677)) xor (layer0_outputs(2048));
    layer1_outputs(5594) <= not(layer0_outputs(8503)) or (layer0_outputs(5465));
    layer1_outputs(5595) <= layer0_outputs(6461);
    layer1_outputs(5596) <= (layer0_outputs(4373)) xor (layer0_outputs(9389));
    layer1_outputs(5597) <= not((layer0_outputs(1442)) xor (layer0_outputs(2045)));
    layer1_outputs(5598) <= not((layer0_outputs(1487)) and (layer0_outputs(6415)));
    layer1_outputs(5599) <= not((layer0_outputs(720)) or (layer0_outputs(6049)));
    layer1_outputs(5600) <= '0';
    layer1_outputs(5601) <= not(layer0_outputs(1847));
    layer1_outputs(5602) <= not(layer0_outputs(2824));
    layer1_outputs(5603) <= not(layer0_outputs(6234));
    layer1_outputs(5604) <= (layer0_outputs(1929)) and not (layer0_outputs(6411));
    layer1_outputs(5605) <= '1';
    layer1_outputs(5606) <= (layer0_outputs(9498)) or (layer0_outputs(2602));
    layer1_outputs(5607) <= not(layer0_outputs(6078));
    layer1_outputs(5608) <= not(layer0_outputs(9349)) or (layer0_outputs(907));
    layer1_outputs(5609) <= not(layer0_outputs(2250)) or (layer0_outputs(6977));
    layer1_outputs(5610) <= layer0_outputs(4049);
    layer1_outputs(5611) <= '1';
    layer1_outputs(5612) <= not(layer0_outputs(6709));
    layer1_outputs(5613) <= (layer0_outputs(7810)) and (layer0_outputs(9130));
    layer1_outputs(5614) <= (layer0_outputs(9185)) and not (layer0_outputs(6690));
    layer1_outputs(5615) <= not((layer0_outputs(4961)) xor (layer0_outputs(5836)));
    layer1_outputs(5616) <= (layer0_outputs(2531)) and not (layer0_outputs(5852));
    layer1_outputs(5617) <= '0';
    layer1_outputs(5618) <= not((layer0_outputs(8906)) xor (layer0_outputs(3156)));
    layer1_outputs(5619) <= '0';
    layer1_outputs(5620) <= not(layer0_outputs(10228));
    layer1_outputs(5621) <= not(layer0_outputs(3681)) or (layer0_outputs(8630));
    layer1_outputs(5622) <= not(layer0_outputs(3891)) or (layer0_outputs(7581));
    layer1_outputs(5623) <= '1';
    layer1_outputs(5624) <= not(layer0_outputs(3578));
    layer1_outputs(5625) <= (layer0_outputs(5962)) or (layer0_outputs(3059));
    layer1_outputs(5626) <= (layer0_outputs(6853)) and (layer0_outputs(1700));
    layer1_outputs(5627) <= (layer0_outputs(794)) and (layer0_outputs(8071));
    layer1_outputs(5628) <= (layer0_outputs(8899)) and not (layer0_outputs(8210));
    layer1_outputs(5629) <= not((layer0_outputs(2331)) xor (layer0_outputs(9595)));
    layer1_outputs(5630) <= '1';
    layer1_outputs(5631) <= not((layer0_outputs(421)) and (layer0_outputs(9959)));
    layer1_outputs(5632) <= '0';
    layer1_outputs(5633) <= (layer0_outputs(4166)) and not (layer0_outputs(426));
    layer1_outputs(5634) <= not((layer0_outputs(1002)) xor (layer0_outputs(7778)));
    layer1_outputs(5635) <= (layer0_outputs(8343)) or (layer0_outputs(7373));
    layer1_outputs(5636) <= (layer0_outputs(8484)) and (layer0_outputs(9924));
    layer1_outputs(5637) <= not(layer0_outputs(9295)) or (layer0_outputs(5520));
    layer1_outputs(5638) <= layer0_outputs(273);
    layer1_outputs(5639) <= (layer0_outputs(570)) and not (layer0_outputs(7760));
    layer1_outputs(5640) <= not((layer0_outputs(2380)) or (layer0_outputs(9782)));
    layer1_outputs(5641) <= layer0_outputs(6474);
    layer1_outputs(5642) <= (layer0_outputs(7177)) and (layer0_outputs(7858));
    layer1_outputs(5643) <= '0';
    layer1_outputs(5644) <= not(layer0_outputs(10090));
    layer1_outputs(5645) <= not((layer0_outputs(3957)) xor (layer0_outputs(628)));
    layer1_outputs(5646) <= layer0_outputs(7015);
    layer1_outputs(5647) <= not(layer0_outputs(6961)) or (layer0_outputs(333));
    layer1_outputs(5648) <= not(layer0_outputs(1629)) or (layer0_outputs(403));
    layer1_outputs(5649) <= (layer0_outputs(4711)) xor (layer0_outputs(3034));
    layer1_outputs(5650) <= not(layer0_outputs(1520));
    layer1_outputs(5651) <= layer0_outputs(6402);
    layer1_outputs(5652) <= not((layer0_outputs(4341)) or (layer0_outputs(3816)));
    layer1_outputs(5653) <= not((layer0_outputs(7112)) xor (layer0_outputs(3034)));
    layer1_outputs(5654) <= (layer0_outputs(7915)) or (layer0_outputs(2337));
    layer1_outputs(5655) <= (layer0_outputs(8791)) and not (layer0_outputs(5680));
    layer1_outputs(5656) <= not(layer0_outputs(4510)) or (layer0_outputs(1739));
    layer1_outputs(5657) <= (layer0_outputs(9871)) and (layer0_outputs(4006));
    layer1_outputs(5658) <= not(layer0_outputs(4162)) or (layer0_outputs(3677));
    layer1_outputs(5659) <= not((layer0_outputs(2136)) and (layer0_outputs(7053)));
    layer1_outputs(5660) <= (layer0_outputs(7102)) xor (layer0_outputs(7509));
    layer1_outputs(5661) <= layer0_outputs(10021);
    layer1_outputs(5662) <= not((layer0_outputs(6438)) and (layer0_outputs(3785)));
    layer1_outputs(5663) <= '1';
    layer1_outputs(5664) <= (layer0_outputs(9523)) and (layer0_outputs(4617));
    layer1_outputs(5665) <= not(layer0_outputs(9818));
    layer1_outputs(5666) <= not((layer0_outputs(8923)) xor (layer0_outputs(5172)));
    layer1_outputs(5667) <= not(layer0_outputs(2724)) or (layer0_outputs(8695));
    layer1_outputs(5668) <= '0';
    layer1_outputs(5669) <= (layer0_outputs(1808)) and not (layer0_outputs(340));
    layer1_outputs(5670) <= (layer0_outputs(6062)) and not (layer0_outputs(9777));
    layer1_outputs(5671) <= not(layer0_outputs(3591));
    layer1_outputs(5672) <= layer0_outputs(7388);
    layer1_outputs(5673) <= not((layer0_outputs(2789)) or (layer0_outputs(3974)));
    layer1_outputs(5674) <= not(layer0_outputs(3421)) or (layer0_outputs(7572));
    layer1_outputs(5675) <= layer0_outputs(7704);
    layer1_outputs(5676) <= not(layer0_outputs(4240));
    layer1_outputs(5677) <= not(layer0_outputs(7410));
    layer1_outputs(5678) <= (layer0_outputs(4914)) and not (layer0_outputs(3778));
    layer1_outputs(5679) <= (layer0_outputs(2125)) and not (layer0_outputs(2852));
    layer1_outputs(5680) <= not((layer0_outputs(9730)) xor (layer0_outputs(9612)));
    layer1_outputs(5681) <= not(layer0_outputs(1066)) or (layer0_outputs(9545));
    layer1_outputs(5682) <= not((layer0_outputs(9081)) or (layer0_outputs(7665)));
    layer1_outputs(5683) <= (layer0_outputs(8902)) and not (layer0_outputs(41));
    layer1_outputs(5684) <= layer0_outputs(5440);
    layer1_outputs(5685) <= not(layer0_outputs(1562));
    layer1_outputs(5686) <= not((layer0_outputs(4984)) and (layer0_outputs(2691)));
    layer1_outputs(5687) <= not(layer0_outputs(5120));
    layer1_outputs(5688) <= not((layer0_outputs(7708)) and (layer0_outputs(153)));
    layer1_outputs(5689) <= (layer0_outputs(3702)) or (layer0_outputs(6136));
    layer1_outputs(5690) <= not((layer0_outputs(1377)) and (layer0_outputs(8625)));
    layer1_outputs(5691) <= layer0_outputs(5304);
    layer1_outputs(5692) <= not(layer0_outputs(5923)) or (layer0_outputs(6065));
    layer1_outputs(5693) <= not((layer0_outputs(6730)) and (layer0_outputs(1186)));
    layer1_outputs(5694) <= not(layer0_outputs(6188));
    layer1_outputs(5695) <= '1';
    layer1_outputs(5696) <= (layer0_outputs(3340)) and (layer0_outputs(7231));
    layer1_outputs(5697) <= (layer0_outputs(1306)) or (layer0_outputs(8243));
    layer1_outputs(5698) <= (layer0_outputs(5080)) and (layer0_outputs(8926));
    layer1_outputs(5699) <= not(layer0_outputs(6205));
    layer1_outputs(5700) <= not(layer0_outputs(7167));
    layer1_outputs(5701) <= not(layer0_outputs(7248));
    layer1_outputs(5702) <= layer0_outputs(3319);
    layer1_outputs(5703) <= not((layer0_outputs(4977)) or (layer0_outputs(5007)));
    layer1_outputs(5704) <= not(layer0_outputs(7272)) or (layer0_outputs(5789));
    layer1_outputs(5705) <= '0';
    layer1_outputs(5706) <= not(layer0_outputs(6677));
    layer1_outputs(5707) <= layer0_outputs(7748);
    layer1_outputs(5708) <= not((layer0_outputs(2791)) xor (layer0_outputs(1795)));
    layer1_outputs(5709) <= (layer0_outputs(7887)) and not (layer0_outputs(5449));
    layer1_outputs(5710) <= (layer0_outputs(2076)) and not (layer0_outputs(5774));
    layer1_outputs(5711) <= not(layer0_outputs(3910)) or (layer0_outputs(2523));
    layer1_outputs(5712) <= (layer0_outputs(5635)) and not (layer0_outputs(7146));
    layer1_outputs(5713) <= not((layer0_outputs(2296)) xor (layer0_outputs(248)));
    layer1_outputs(5714) <= not(layer0_outputs(8905)) or (layer0_outputs(1413));
    layer1_outputs(5715) <= (layer0_outputs(8372)) or (layer0_outputs(5627));
    layer1_outputs(5716) <= (layer0_outputs(7892)) and (layer0_outputs(8242));
    layer1_outputs(5717) <= not(layer0_outputs(7871));
    layer1_outputs(5718) <= (layer0_outputs(1177)) and not (layer0_outputs(7437));
    layer1_outputs(5719) <= not((layer0_outputs(2359)) or (layer0_outputs(181)));
    layer1_outputs(5720) <= (layer0_outputs(7316)) or (layer0_outputs(6888));
    layer1_outputs(5721) <= not(layer0_outputs(8458)) or (layer0_outputs(2805));
    layer1_outputs(5722) <= (layer0_outputs(4127)) and not (layer0_outputs(2682));
    layer1_outputs(5723) <= not((layer0_outputs(3583)) xor (layer0_outputs(9492)));
    layer1_outputs(5724) <= (layer0_outputs(3531)) and not (layer0_outputs(7992));
    layer1_outputs(5725) <= not(layer0_outputs(8871));
    layer1_outputs(5726) <= layer0_outputs(1897);
    layer1_outputs(5727) <= not(layer0_outputs(4164));
    layer1_outputs(5728) <= (layer0_outputs(5044)) or (layer0_outputs(5711));
    layer1_outputs(5729) <= not(layer0_outputs(5350)) or (layer0_outputs(7366));
    layer1_outputs(5730) <= '1';
    layer1_outputs(5731) <= not((layer0_outputs(8328)) or (layer0_outputs(10094)));
    layer1_outputs(5732) <= (layer0_outputs(4594)) and not (layer0_outputs(5538));
    layer1_outputs(5733) <= not(layer0_outputs(9638)) or (layer0_outputs(8289));
    layer1_outputs(5734) <= layer0_outputs(4149);
    layer1_outputs(5735) <= layer0_outputs(1281);
    layer1_outputs(5736) <= layer0_outputs(8954);
    layer1_outputs(5737) <= not((layer0_outputs(2035)) or (layer0_outputs(2582)));
    layer1_outputs(5738) <= '1';
    layer1_outputs(5739) <= not(layer0_outputs(5265)) or (layer0_outputs(7047));
    layer1_outputs(5740) <= layer0_outputs(845);
    layer1_outputs(5741) <= not((layer0_outputs(1679)) and (layer0_outputs(913)));
    layer1_outputs(5742) <= (layer0_outputs(582)) and (layer0_outputs(5656));
    layer1_outputs(5743) <= not(layer0_outputs(4698));
    layer1_outputs(5744) <= not(layer0_outputs(9558));
    layer1_outputs(5745) <= not(layer0_outputs(6573));
    layer1_outputs(5746) <= not(layer0_outputs(1346));
    layer1_outputs(5747) <= not(layer0_outputs(6636));
    layer1_outputs(5748) <= not((layer0_outputs(5755)) or (layer0_outputs(1733)));
    layer1_outputs(5749) <= (layer0_outputs(5502)) or (layer0_outputs(8571));
    layer1_outputs(5750) <= '1';
    layer1_outputs(5751) <= not((layer0_outputs(3385)) xor (layer0_outputs(573)));
    layer1_outputs(5752) <= layer0_outputs(4031);
    layer1_outputs(5753) <= (layer0_outputs(2231)) or (layer0_outputs(7837));
    layer1_outputs(5754) <= not(layer0_outputs(5576));
    layer1_outputs(5755) <= not((layer0_outputs(7326)) and (layer0_outputs(6395)));
    layer1_outputs(5756) <= (layer0_outputs(1824)) or (layer0_outputs(6541));
    layer1_outputs(5757) <= layer0_outputs(7643);
    layer1_outputs(5758) <= (layer0_outputs(6797)) and (layer0_outputs(5761));
    layer1_outputs(5759) <= (layer0_outputs(6344)) xor (layer0_outputs(832));
    layer1_outputs(5760) <= not(layer0_outputs(8327));
    layer1_outputs(5761) <= not(layer0_outputs(4434));
    layer1_outputs(5762) <= not(layer0_outputs(4428)) or (layer0_outputs(3075));
    layer1_outputs(5763) <= not(layer0_outputs(8036));
    layer1_outputs(5764) <= '1';
    layer1_outputs(5765) <= layer0_outputs(8281);
    layer1_outputs(5766) <= not(layer0_outputs(901)) or (layer0_outputs(4353));
    layer1_outputs(5767) <= not(layer0_outputs(6025)) or (layer0_outputs(3618));
    layer1_outputs(5768) <= layer0_outputs(5428);
    layer1_outputs(5769) <= layer0_outputs(2222);
    layer1_outputs(5770) <= not(layer0_outputs(9881));
    layer1_outputs(5771) <= (layer0_outputs(6662)) and not (layer0_outputs(3300));
    layer1_outputs(5772) <= not((layer0_outputs(1361)) or (layer0_outputs(1151)));
    layer1_outputs(5773) <= layer0_outputs(3014);
    layer1_outputs(5774) <= not(layer0_outputs(1205));
    layer1_outputs(5775) <= (layer0_outputs(1246)) xor (layer0_outputs(8039));
    layer1_outputs(5776) <= (layer0_outputs(9714)) and (layer0_outputs(5373));
    layer1_outputs(5777) <= not(layer0_outputs(846)) or (layer0_outputs(5667));
    layer1_outputs(5778) <= layer0_outputs(352);
    layer1_outputs(5779) <= layer0_outputs(2862);
    layer1_outputs(5780) <= not(layer0_outputs(8178)) or (layer0_outputs(9404));
    layer1_outputs(5781) <= (layer0_outputs(5074)) and (layer0_outputs(1380));
    layer1_outputs(5782) <= '0';
    layer1_outputs(5783) <= '1';
    layer1_outputs(5784) <= (layer0_outputs(1378)) xor (layer0_outputs(8960));
    layer1_outputs(5785) <= not(layer0_outputs(6054));
    layer1_outputs(5786) <= not(layer0_outputs(5873));
    layer1_outputs(5787) <= not((layer0_outputs(3898)) and (layer0_outputs(4702)));
    layer1_outputs(5788) <= (layer0_outputs(2950)) or (layer0_outputs(8841));
    layer1_outputs(5789) <= not((layer0_outputs(1728)) and (layer0_outputs(3964)));
    layer1_outputs(5790) <= layer0_outputs(7362);
    layer1_outputs(5791) <= not((layer0_outputs(2859)) or (layer0_outputs(6958)));
    layer1_outputs(5792) <= (layer0_outputs(9723)) and not (layer0_outputs(5854));
    layer1_outputs(5793) <= not(layer0_outputs(8154)) or (layer0_outputs(2078));
    layer1_outputs(5794) <= not((layer0_outputs(5322)) xor (layer0_outputs(1440)));
    layer1_outputs(5795) <= (layer0_outputs(2016)) and (layer0_outputs(1566));
    layer1_outputs(5796) <= layer0_outputs(4817);
    layer1_outputs(5797) <= not(layer0_outputs(1790));
    layer1_outputs(5798) <= not(layer0_outputs(2883));
    layer1_outputs(5799) <= '0';
    layer1_outputs(5800) <= not(layer0_outputs(4726));
    layer1_outputs(5801) <= (layer0_outputs(6684)) and (layer0_outputs(4334));
    layer1_outputs(5802) <= not(layer0_outputs(4117));
    layer1_outputs(5803) <= (layer0_outputs(556)) and not (layer0_outputs(6291));
    layer1_outputs(5804) <= not(layer0_outputs(9109)) or (layer0_outputs(2830));
    layer1_outputs(5805) <= not(layer0_outputs(7810)) or (layer0_outputs(1676));
    layer1_outputs(5806) <= not(layer0_outputs(8558)) or (layer0_outputs(3725));
    layer1_outputs(5807) <= not(layer0_outputs(1407)) or (layer0_outputs(7227));
    layer1_outputs(5808) <= layer0_outputs(3792);
    layer1_outputs(5809) <= (layer0_outputs(9013)) and not (layer0_outputs(6815));
    layer1_outputs(5810) <= (layer0_outputs(2973)) or (layer0_outputs(1511));
    layer1_outputs(5811) <= (layer0_outputs(9025)) and (layer0_outputs(1022));
    layer1_outputs(5812) <= (layer0_outputs(9368)) and not (layer0_outputs(5179));
    layer1_outputs(5813) <= not(layer0_outputs(2710));
    layer1_outputs(5814) <= not((layer0_outputs(6984)) xor (layer0_outputs(1061)));
    layer1_outputs(5815) <= layer0_outputs(9999);
    layer1_outputs(5816) <= layer0_outputs(3147);
    layer1_outputs(5817) <= (layer0_outputs(2325)) xor (layer0_outputs(5924));
    layer1_outputs(5818) <= not((layer0_outputs(7797)) and (layer0_outputs(6271)));
    layer1_outputs(5819) <= '1';
    layer1_outputs(5820) <= not(layer0_outputs(2088));
    layer1_outputs(5821) <= layer0_outputs(9183);
    layer1_outputs(5822) <= '1';
    layer1_outputs(5823) <= layer0_outputs(4809);
    layer1_outputs(5824) <= not(layer0_outputs(6040));
    layer1_outputs(5825) <= (layer0_outputs(10070)) xor (layer0_outputs(9617));
    layer1_outputs(5826) <= not(layer0_outputs(8784));
    layer1_outputs(5827) <= not(layer0_outputs(5194)) or (layer0_outputs(4666));
    layer1_outputs(5828) <= layer0_outputs(5603);
    layer1_outputs(5829) <= (layer0_outputs(7221)) and not (layer0_outputs(5266));
    layer1_outputs(5830) <= not(layer0_outputs(6884));
    layer1_outputs(5831) <= (layer0_outputs(7566)) xor (layer0_outputs(9007));
    layer1_outputs(5832) <= (layer0_outputs(5664)) xor (layer0_outputs(9638));
    layer1_outputs(5833) <= not(layer0_outputs(5652)) or (layer0_outputs(3529));
    layer1_outputs(5834) <= not(layer0_outputs(4680));
    layer1_outputs(5835) <= not(layer0_outputs(3157)) or (layer0_outputs(5477));
    layer1_outputs(5836) <= not(layer0_outputs(197)) or (layer0_outputs(1085));
    layer1_outputs(5837) <= '1';
    layer1_outputs(5838) <= layer0_outputs(8808);
    layer1_outputs(5839) <= layer0_outputs(7966);
    layer1_outputs(5840) <= layer0_outputs(5058);
    layer1_outputs(5841) <= layer0_outputs(521);
    layer1_outputs(5842) <= not(layer0_outputs(3719)) or (layer0_outputs(5119));
    layer1_outputs(5843) <= not((layer0_outputs(5625)) and (layer0_outputs(7176)));
    layer1_outputs(5844) <= not((layer0_outputs(5226)) xor (layer0_outputs(4702)));
    layer1_outputs(5845) <= not(layer0_outputs(5920));
    layer1_outputs(5846) <= (layer0_outputs(5676)) and (layer0_outputs(4797));
    layer1_outputs(5847) <= layer0_outputs(87);
    layer1_outputs(5848) <= not(layer0_outputs(3453));
    layer1_outputs(5849) <= (layer0_outputs(814)) or (layer0_outputs(5032));
    layer1_outputs(5850) <= layer0_outputs(1991);
    layer1_outputs(5851) <= (layer0_outputs(902)) or (layer0_outputs(6446));
    layer1_outputs(5852) <= not(layer0_outputs(7291)) or (layer0_outputs(7885));
    layer1_outputs(5853) <= (layer0_outputs(3069)) and not (layer0_outputs(3090));
    layer1_outputs(5854) <= not((layer0_outputs(2420)) or (layer0_outputs(1795)));
    layer1_outputs(5855) <= not(layer0_outputs(4669));
    layer1_outputs(5856) <= (layer0_outputs(6807)) and not (layer0_outputs(805));
    layer1_outputs(5857) <= not((layer0_outputs(2828)) or (layer0_outputs(5363)));
    layer1_outputs(5858) <= (layer0_outputs(2071)) or (layer0_outputs(9091));
    layer1_outputs(5859) <= (layer0_outputs(7584)) and not (layer0_outputs(6099));
    layer1_outputs(5860) <= not(layer0_outputs(9160));
    layer1_outputs(5861) <= not(layer0_outputs(6718));
    layer1_outputs(5862) <= layer0_outputs(9239);
    layer1_outputs(5863) <= layer0_outputs(102);
    layer1_outputs(5864) <= '1';
    layer1_outputs(5865) <= (layer0_outputs(9603)) xor (layer0_outputs(2510));
    layer1_outputs(5866) <= not((layer0_outputs(6740)) or (layer0_outputs(7380)));
    layer1_outputs(5867) <= (layer0_outputs(9138)) and (layer0_outputs(9641));
    layer1_outputs(5868) <= (layer0_outputs(5689)) and not (layer0_outputs(5137));
    layer1_outputs(5869) <= not(layer0_outputs(6183)) or (layer0_outputs(9201));
    layer1_outputs(5870) <= not(layer0_outputs(9997)) or (layer0_outputs(2230));
    layer1_outputs(5871) <= not((layer0_outputs(3496)) xor (layer0_outputs(9609)));
    layer1_outputs(5872) <= layer0_outputs(8568);
    layer1_outputs(5873) <= (layer0_outputs(3221)) and not (layer0_outputs(6090));
    layer1_outputs(5874) <= not(layer0_outputs(1045));
    layer1_outputs(5875) <= (layer0_outputs(4632)) or (layer0_outputs(7170));
    layer1_outputs(5876) <= not(layer0_outputs(1807)) or (layer0_outputs(4931));
    layer1_outputs(5877) <= '0';
    layer1_outputs(5878) <= not((layer0_outputs(3101)) xor (layer0_outputs(3200)));
    layer1_outputs(5879) <= not((layer0_outputs(7720)) and (layer0_outputs(8251)));
    layer1_outputs(5880) <= layer0_outputs(4039);
    layer1_outputs(5881) <= (layer0_outputs(5684)) xor (layer0_outputs(3055));
    layer1_outputs(5882) <= layer0_outputs(3315);
    layer1_outputs(5883) <= not((layer0_outputs(720)) and (layer0_outputs(242)));
    layer1_outputs(5884) <= not(layer0_outputs(2280));
    layer1_outputs(5885) <= not(layer0_outputs(897));
    layer1_outputs(5886) <= not(layer0_outputs(8904)) or (layer0_outputs(8796));
    layer1_outputs(5887) <= (layer0_outputs(6874)) and not (layer0_outputs(4012));
    layer1_outputs(5888) <= layer0_outputs(4781);
    layer1_outputs(5889) <= layer0_outputs(1395);
    layer1_outputs(5890) <= not((layer0_outputs(9568)) or (layer0_outputs(7087)));
    layer1_outputs(5891) <= (layer0_outputs(5495)) xor (layer0_outputs(3860));
    layer1_outputs(5892) <= not(layer0_outputs(4038));
    layer1_outputs(5893) <= not(layer0_outputs(6439)) or (layer0_outputs(10040));
    layer1_outputs(5894) <= not((layer0_outputs(4162)) xor (layer0_outputs(9991)));
    layer1_outputs(5895) <= (layer0_outputs(3096)) and not (layer0_outputs(6050));
    layer1_outputs(5896) <= not(layer0_outputs(8021)) or (layer0_outputs(594));
    layer1_outputs(5897) <= not((layer0_outputs(5758)) and (layer0_outputs(6748)));
    layer1_outputs(5898) <= not(layer0_outputs(9353)) or (layer0_outputs(2104));
    layer1_outputs(5899) <= not((layer0_outputs(10168)) or (layer0_outputs(351)));
    layer1_outputs(5900) <= layer0_outputs(8940);
    layer1_outputs(5901) <= not(layer0_outputs(7288));
    layer1_outputs(5902) <= layer0_outputs(5789);
    layer1_outputs(5903) <= (layer0_outputs(4758)) and not (layer0_outputs(4535));
    layer1_outputs(5904) <= '0';
    layer1_outputs(5905) <= layer0_outputs(629);
    layer1_outputs(5906) <= '1';
    layer1_outputs(5907) <= layer0_outputs(3823);
    layer1_outputs(5908) <= not((layer0_outputs(4788)) xor (layer0_outputs(4843)));
    layer1_outputs(5909) <= (layer0_outputs(3056)) or (layer0_outputs(3213));
    layer1_outputs(5910) <= (layer0_outputs(7475)) and not (layer0_outputs(9428));
    layer1_outputs(5911) <= (layer0_outputs(3127)) and (layer0_outputs(18));
    layer1_outputs(5912) <= (layer0_outputs(9455)) or (layer0_outputs(1947));
    layer1_outputs(5913) <= not(layer0_outputs(6115));
    layer1_outputs(5914) <= (layer0_outputs(5136)) and (layer0_outputs(6590));
    layer1_outputs(5915) <= not((layer0_outputs(3263)) and (layer0_outputs(1216)));
    layer1_outputs(5916) <= '1';
    layer1_outputs(5917) <= (layer0_outputs(3570)) or (layer0_outputs(9917));
    layer1_outputs(5918) <= layer0_outputs(7289);
    layer1_outputs(5919) <= (layer0_outputs(2044)) and not (layer0_outputs(1991));
    layer1_outputs(5920) <= (layer0_outputs(1384)) and not (layer0_outputs(2202));
    layer1_outputs(5921) <= '0';
    layer1_outputs(5922) <= not(layer0_outputs(937));
    layer1_outputs(5923) <= layer0_outputs(3306);
    layer1_outputs(5924) <= (layer0_outputs(8731)) and not (layer0_outputs(168));
    layer1_outputs(5925) <= layer0_outputs(6232);
    layer1_outputs(5926) <= not((layer0_outputs(1485)) or (layer0_outputs(9806)));
    layer1_outputs(5927) <= (layer0_outputs(8822)) xor (layer0_outputs(5685));
    layer1_outputs(5928) <= '1';
    layer1_outputs(5929) <= (layer0_outputs(2225)) xor (layer0_outputs(7637));
    layer1_outputs(5930) <= not(layer0_outputs(1942)) or (layer0_outputs(3183));
    layer1_outputs(5931) <= (layer0_outputs(4763)) xor (layer0_outputs(7335));
    layer1_outputs(5932) <= '0';
    layer1_outputs(5933) <= '1';
    layer1_outputs(5934) <= not(layer0_outputs(1203)) or (layer0_outputs(7392));
    layer1_outputs(5935) <= layer0_outputs(6676);
    layer1_outputs(5936) <= layer0_outputs(1246);
    layer1_outputs(5937) <= not((layer0_outputs(6410)) or (layer0_outputs(4381)));
    layer1_outputs(5938) <= not(layer0_outputs(2561)) or (layer0_outputs(9339));
    layer1_outputs(5939) <= (layer0_outputs(3444)) and (layer0_outputs(5359));
    layer1_outputs(5940) <= (layer0_outputs(6454)) or (layer0_outputs(2753));
    layer1_outputs(5941) <= not(layer0_outputs(8392)) or (layer0_outputs(7049));
    layer1_outputs(5942) <= not(layer0_outputs(8936));
    layer1_outputs(5943) <= not((layer0_outputs(2883)) or (layer0_outputs(1652)));
    layer1_outputs(5944) <= layer0_outputs(3897);
    layer1_outputs(5945) <= (layer0_outputs(1183)) and (layer0_outputs(1030));
    layer1_outputs(5946) <= not((layer0_outputs(6119)) and (layer0_outputs(4021)));
    layer1_outputs(5947) <= not((layer0_outputs(1051)) and (layer0_outputs(4139)));
    layer1_outputs(5948) <= (layer0_outputs(807)) or (layer0_outputs(3107));
    layer1_outputs(5949) <= not((layer0_outputs(801)) xor (layer0_outputs(9982)));
    layer1_outputs(5950) <= (layer0_outputs(1719)) and (layer0_outputs(2418));
    layer1_outputs(5951) <= not(layer0_outputs(717));
    layer1_outputs(5952) <= not(layer0_outputs(8331)) or (layer0_outputs(8603));
    layer1_outputs(5953) <= not((layer0_outputs(1399)) xor (layer0_outputs(5349)));
    layer1_outputs(5954) <= layer0_outputs(8682);
    layer1_outputs(5955) <= layer0_outputs(9842);
    layer1_outputs(5956) <= not((layer0_outputs(8894)) xor (layer0_outputs(10190)));
    layer1_outputs(5957) <= (layer0_outputs(2749)) and not (layer0_outputs(9836));
    layer1_outputs(5958) <= layer0_outputs(6780);
    layer1_outputs(5959) <= (layer0_outputs(7745)) xor (layer0_outputs(6965));
    layer1_outputs(5960) <= (layer0_outputs(9766)) or (layer0_outputs(8354));
    layer1_outputs(5961) <= '0';
    layer1_outputs(5962) <= not(layer0_outputs(3338));
    layer1_outputs(5963) <= (layer0_outputs(5668)) and (layer0_outputs(6945));
    layer1_outputs(5964) <= not((layer0_outputs(5977)) and (layer0_outputs(6906)));
    layer1_outputs(5965) <= layer0_outputs(5933);
    layer1_outputs(5966) <= not((layer0_outputs(3232)) xor (layer0_outputs(84)));
    layer1_outputs(5967) <= (layer0_outputs(10119)) and not (layer0_outputs(616));
    layer1_outputs(5968) <= not(layer0_outputs(5185));
    layer1_outputs(5969) <= not(layer0_outputs(8563));
    layer1_outputs(5970) <= '0';
    layer1_outputs(5971) <= layer0_outputs(7493);
    layer1_outputs(5972) <= not(layer0_outputs(9244));
    layer1_outputs(5973) <= not(layer0_outputs(2009)) or (layer0_outputs(3453));
    layer1_outputs(5974) <= not(layer0_outputs(5960));
    layer1_outputs(5975) <= (layer0_outputs(9980)) xor (layer0_outputs(5602));
    layer1_outputs(5976) <= not(layer0_outputs(6753)) or (layer0_outputs(3498));
    layer1_outputs(5977) <= not(layer0_outputs(2169));
    layer1_outputs(5978) <= not((layer0_outputs(6012)) and (layer0_outputs(5274)));
    layer1_outputs(5979) <= not((layer0_outputs(3665)) or (layer0_outputs(33)));
    layer1_outputs(5980) <= not((layer0_outputs(6260)) and (layer0_outputs(4473)));
    layer1_outputs(5981) <= not(layer0_outputs(2386)) or (layer0_outputs(7064));
    layer1_outputs(5982) <= not(layer0_outputs(4717)) or (layer0_outputs(1857));
    layer1_outputs(5983) <= not((layer0_outputs(4018)) xor (layer0_outputs(332)));
    layer1_outputs(5984) <= layer0_outputs(3882);
    layer1_outputs(5985) <= layer0_outputs(9921);
    layer1_outputs(5986) <= not(layer0_outputs(4001));
    layer1_outputs(5987) <= not((layer0_outputs(9062)) or (layer0_outputs(2868)));
    layer1_outputs(5988) <= layer0_outputs(1017);
    layer1_outputs(5989) <= not(layer0_outputs(8793));
    layer1_outputs(5990) <= not((layer0_outputs(8407)) xor (layer0_outputs(2466)));
    layer1_outputs(5991) <= not((layer0_outputs(7769)) or (layer0_outputs(8990)));
    layer1_outputs(5992) <= (layer0_outputs(9371)) and not (layer0_outputs(9297));
    layer1_outputs(5993) <= (layer0_outputs(3387)) and (layer0_outputs(1464));
    layer1_outputs(5994) <= not(layer0_outputs(6263));
    layer1_outputs(5995) <= (layer0_outputs(7856)) or (layer0_outputs(1196));
    layer1_outputs(5996) <= not(layer0_outputs(2620)) or (layer0_outputs(9759));
    layer1_outputs(5997) <= not(layer0_outputs(5829)) or (layer0_outputs(9039));
    layer1_outputs(5998) <= (layer0_outputs(9696)) and not (layer0_outputs(3251));
    layer1_outputs(5999) <= (layer0_outputs(6364)) and not (layer0_outputs(3215));
    layer1_outputs(6000) <= not(layer0_outputs(1828));
    layer1_outputs(6001) <= not(layer0_outputs(3080)) or (layer0_outputs(3073));
    layer1_outputs(6002) <= layer0_outputs(2313);
    layer1_outputs(6003) <= not(layer0_outputs(853)) or (layer0_outputs(2117));
    layer1_outputs(6004) <= (layer0_outputs(1680)) xor (layer0_outputs(1208));
    layer1_outputs(6005) <= '1';
    layer1_outputs(6006) <= (layer0_outputs(672)) and not (layer0_outputs(1218));
    layer1_outputs(6007) <= (layer0_outputs(4492)) or (layer0_outputs(4270));
    layer1_outputs(6008) <= (layer0_outputs(3801)) and (layer0_outputs(527));
    layer1_outputs(6009) <= not((layer0_outputs(3468)) and (layer0_outputs(1993)));
    layer1_outputs(6010) <= '0';
    layer1_outputs(6011) <= layer0_outputs(9815);
    layer1_outputs(6012) <= not((layer0_outputs(5420)) xor (layer0_outputs(8670)));
    layer1_outputs(6013) <= not((layer0_outputs(625)) xor (layer0_outputs(7495)));
    layer1_outputs(6014) <= (layer0_outputs(8958)) xor (layer0_outputs(8957));
    layer1_outputs(6015) <= layer0_outputs(7585);
    layer1_outputs(6016) <= not((layer0_outputs(8786)) and (layer0_outputs(6007)));
    layer1_outputs(6017) <= layer0_outputs(6837);
    layer1_outputs(6018) <= (layer0_outputs(9495)) xor (layer0_outputs(1702));
    layer1_outputs(6019) <= not(layer0_outputs(5475));
    layer1_outputs(6020) <= not(layer0_outputs(9324));
    layer1_outputs(6021) <= layer0_outputs(8092);
    layer1_outputs(6022) <= (layer0_outputs(2349)) or (layer0_outputs(7312));
    layer1_outputs(6023) <= not(layer0_outputs(7707)) or (layer0_outputs(9969));
    layer1_outputs(6024) <= (layer0_outputs(3684)) and not (layer0_outputs(966));
    layer1_outputs(6025) <= not(layer0_outputs(5524));
    layer1_outputs(6026) <= not(layer0_outputs(9462)) or (layer0_outputs(3858));
    layer1_outputs(6027) <= not(layer0_outputs(2015));
    layer1_outputs(6028) <= not((layer0_outputs(234)) xor (layer0_outputs(473)));
    layer1_outputs(6029) <= not(layer0_outputs(4789)) or (layer0_outputs(227));
    layer1_outputs(6030) <= '0';
    layer1_outputs(6031) <= layer0_outputs(6011);
    layer1_outputs(6032) <= not(layer0_outputs(3042)) or (layer0_outputs(9825));
    layer1_outputs(6033) <= (layer0_outputs(5337)) and (layer0_outputs(900));
    layer1_outputs(6034) <= not((layer0_outputs(1244)) or (layer0_outputs(5654)));
    layer1_outputs(6035) <= not((layer0_outputs(1671)) xor (layer0_outputs(1859)));
    layer1_outputs(6036) <= not((layer0_outputs(1421)) and (layer0_outputs(3399)));
    layer1_outputs(6037) <= not(layer0_outputs(2718));
    layer1_outputs(6038) <= (layer0_outputs(2263)) xor (layer0_outputs(5034));
    layer1_outputs(6039) <= (layer0_outputs(3514)) xor (layer0_outputs(557));
    layer1_outputs(6040) <= (layer0_outputs(3313)) and not (layer0_outputs(6360));
    layer1_outputs(6041) <= not((layer0_outputs(8431)) and (layer0_outputs(5014)));
    layer1_outputs(6042) <= not(layer0_outputs(4280));
    layer1_outputs(6043) <= not((layer0_outputs(6803)) xor (layer0_outputs(595)));
    layer1_outputs(6044) <= (layer0_outputs(3894)) or (layer0_outputs(7960));
    layer1_outputs(6045) <= not((layer0_outputs(7869)) or (layer0_outputs(6719)));
    layer1_outputs(6046) <= not((layer0_outputs(9133)) or (layer0_outputs(5095)));
    layer1_outputs(6047) <= not(layer0_outputs(9320));
    layer1_outputs(6048) <= not(layer0_outputs(831));
    layer1_outputs(6049) <= not((layer0_outputs(7060)) and (layer0_outputs(1370)));
    layer1_outputs(6050) <= layer0_outputs(1330);
    layer1_outputs(6051) <= not(layer0_outputs(2268));
    layer1_outputs(6052) <= not((layer0_outputs(6495)) xor (layer0_outputs(7689)));
    layer1_outputs(6053) <= not(layer0_outputs(9097)) or (layer0_outputs(2724));
    layer1_outputs(6054) <= (layer0_outputs(2932)) xor (layer0_outputs(4597));
    layer1_outputs(6055) <= (layer0_outputs(3873)) xor (layer0_outputs(9534));
    layer1_outputs(6056) <= '1';
    layer1_outputs(6057) <= (layer0_outputs(4822)) or (layer0_outputs(5039));
    layer1_outputs(6058) <= (layer0_outputs(9222)) and (layer0_outputs(12));
    layer1_outputs(6059) <= (layer0_outputs(10158)) and not (layer0_outputs(10128));
    layer1_outputs(6060) <= not((layer0_outputs(8496)) and (layer0_outputs(8774)));
    layer1_outputs(6061) <= (layer0_outputs(9429)) and not (layer0_outputs(4126));
    layer1_outputs(6062) <= not(layer0_outputs(2042));
    layer1_outputs(6063) <= (layer0_outputs(4487)) and (layer0_outputs(5030));
    layer1_outputs(6064) <= not((layer0_outputs(5516)) xor (layer0_outputs(8773)));
    layer1_outputs(6065) <= layer0_outputs(32);
    layer1_outputs(6066) <= not(layer0_outputs(1760));
    layer1_outputs(6067) <= not((layer0_outputs(2037)) xor (layer0_outputs(663)));
    layer1_outputs(6068) <= '0';
    layer1_outputs(6069) <= layer0_outputs(5905);
    layer1_outputs(6070) <= (layer0_outputs(2911)) or (layer0_outputs(6487));
    layer1_outputs(6071) <= (layer0_outputs(5866)) xor (layer0_outputs(3178));
    layer1_outputs(6072) <= not(layer0_outputs(6475)) or (layer0_outputs(6430));
    layer1_outputs(6073) <= layer0_outputs(2255);
    layer1_outputs(6074) <= layer0_outputs(702);
    layer1_outputs(6075) <= not((layer0_outputs(7395)) xor (layer0_outputs(4221)));
    layer1_outputs(6076) <= not(layer0_outputs(4954));
    layer1_outputs(6077) <= (layer0_outputs(750)) or (layer0_outputs(1368));
    layer1_outputs(6078) <= not((layer0_outputs(7628)) or (layer0_outputs(9161)));
    layer1_outputs(6079) <= not(layer0_outputs(6942));
    layer1_outputs(6080) <= '1';
    layer1_outputs(6081) <= (layer0_outputs(7157)) and (layer0_outputs(7353));
    layer1_outputs(6082) <= not((layer0_outputs(9859)) xor (layer0_outputs(398)));
    layer1_outputs(6083) <= not(layer0_outputs(2786)) or (layer0_outputs(6800));
    layer1_outputs(6084) <= layer0_outputs(8188);
    layer1_outputs(6085) <= (layer0_outputs(1932)) and not (layer0_outputs(4462));
    layer1_outputs(6086) <= (layer0_outputs(760)) xor (layer0_outputs(6520));
    layer1_outputs(6087) <= not((layer0_outputs(9539)) or (layer0_outputs(7000)));
    layer1_outputs(6088) <= not(layer0_outputs(3045));
    layer1_outputs(6089) <= not(layer0_outputs(3438)) or (layer0_outputs(8459));
    layer1_outputs(6090) <= not((layer0_outputs(9560)) and (layer0_outputs(2018)));
    layer1_outputs(6091) <= (layer0_outputs(4077)) and not (layer0_outputs(7032));
    layer1_outputs(6092) <= (layer0_outputs(174)) and (layer0_outputs(9665));
    layer1_outputs(6093) <= layer0_outputs(2720);
    layer1_outputs(6094) <= not(layer0_outputs(7955)) or (layer0_outputs(8837));
    layer1_outputs(6095) <= not(layer0_outputs(7066)) or (layer0_outputs(2376));
    layer1_outputs(6096) <= (layer0_outputs(9557)) or (layer0_outputs(8400));
    layer1_outputs(6097) <= not(layer0_outputs(3045)) or (layer0_outputs(8272));
    layer1_outputs(6098) <= (layer0_outputs(7801)) and not (layer0_outputs(4987));
    layer1_outputs(6099) <= (layer0_outputs(5732)) or (layer0_outputs(6279));
    layer1_outputs(6100) <= not(layer0_outputs(6682));
    layer1_outputs(6101) <= layer0_outputs(5925);
    layer1_outputs(6102) <= not(layer0_outputs(2111));
    layer1_outputs(6103) <= not(layer0_outputs(493));
    layer1_outputs(6104) <= not(layer0_outputs(7253)) or (layer0_outputs(3402));
    layer1_outputs(6105) <= (layer0_outputs(1673)) or (layer0_outputs(913));
    layer1_outputs(6106) <= (layer0_outputs(7548)) and (layer0_outputs(7157));
    layer1_outputs(6107) <= (layer0_outputs(7887)) and not (layer0_outputs(9508));
    layer1_outputs(6108) <= not(layer0_outputs(7519));
    layer1_outputs(6109) <= (layer0_outputs(6203)) and (layer0_outputs(480));
    layer1_outputs(6110) <= (layer0_outputs(6532)) and not (layer0_outputs(4366));
    layer1_outputs(6111) <= (layer0_outputs(3466)) xor (layer0_outputs(841));
    layer1_outputs(6112) <= layer0_outputs(3928);
    layer1_outputs(6113) <= layer0_outputs(272);
    layer1_outputs(6114) <= layer0_outputs(9632);
    layer1_outputs(6115) <= not(layer0_outputs(4941)) or (layer0_outputs(4544));
    layer1_outputs(6116) <= (layer0_outputs(197)) xor (layer0_outputs(3836));
    layer1_outputs(6117) <= layer0_outputs(5396);
    layer1_outputs(6118) <= (layer0_outputs(5853)) or (layer0_outputs(3291));
    layer1_outputs(6119) <= '1';
    layer1_outputs(6120) <= not(layer0_outputs(10226));
    layer1_outputs(6121) <= not((layer0_outputs(2818)) or (layer0_outputs(3660)));
    layer1_outputs(6122) <= not(layer0_outputs(7220));
    layer1_outputs(6123) <= (layer0_outputs(1763)) or (layer0_outputs(7312));
    layer1_outputs(6124) <= '1';
    layer1_outputs(6125) <= (layer0_outputs(3132)) and not (layer0_outputs(8122));
    layer1_outputs(6126) <= not(layer0_outputs(2386));
    layer1_outputs(6127) <= not(layer0_outputs(599)) or (layer0_outputs(7403));
    layer1_outputs(6128) <= (layer0_outputs(6207)) and not (layer0_outputs(3909));
    layer1_outputs(6129) <= not(layer0_outputs(6957)) or (layer0_outputs(9566));
    layer1_outputs(6130) <= layer0_outputs(7442);
    layer1_outputs(6131) <= not(layer0_outputs(7272));
    layer1_outputs(6132) <= (layer0_outputs(712)) and (layer0_outputs(229));
    layer1_outputs(6133) <= (layer0_outputs(799)) and (layer0_outputs(7427));
    layer1_outputs(6134) <= (layer0_outputs(5813)) xor (layer0_outputs(8909));
    layer1_outputs(6135) <= not(layer0_outputs(4654));
    layer1_outputs(6136) <= (layer0_outputs(7382)) xor (layer0_outputs(4040));
    layer1_outputs(6137) <= (layer0_outputs(771)) or (layer0_outputs(6391));
    layer1_outputs(6138) <= layer0_outputs(9195);
    layer1_outputs(6139) <= (layer0_outputs(4536)) xor (layer0_outputs(6442));
    layer1_outputs(6140) <= layer0_outputs(4262);
    layer1_outputs(6141) <= not(layer0_outputs(5189));
    layer1_outputs(6142) <= not(layer0_outputs(1362));
    layer1_outputs(6143) <= not((layer0_outputs(5460)) or (layer0_outputs(3180)));
    layer1_outputs(6144) <= not(layer0_outputs(4193)) or (layer0_outputs(4513));
    layer1_outputs(6145) <= not(layer0_outputs(1351)) or (layer0_outputs(5611));
    layer1_outputs(6146) <= not(layer0_outputs(5298));
    layer1_outputs(6147) <= not(layer0_outputs(6409));
    layer1_outputs(6148) <= not((layer0_outputs(6522)) or (layer0_outputs(5308)));
    layer1_outputs(6149) <= not((layer0_outputs(9414)) xor (layer0_outputs(1254)));
    layer1_outputs(6150) <= not((layer0_outputs(6644)) and (layer0_outputs(7357)));
    layer1_outputs(6151) <= (layer0_outputs(6963)) and (layer0_outputs(3186));
    layer1_outputs(6152) <= not(layer0_outputs(829));
    layer1_outputs(6153) <= not(layer0_outputs(1274));
    layer1_outputs(6154) <= not((layer0_outputs(836)) and (layer0_outputs(3968)));
    layer1_outputs(6155) <= not(layer0_outputs(935));
    layer1_outputs(6156) <= '1';
    layer1_outputs(6157) <= not(layer0_outputs(273));
    layer1_outputs(6158) <= (layer0_outputs(1713)) and (layer0_outputs(1173));
    layer1_outputs(6159) <= (layer0_outputs(9027)) and not (layer0_outputs(5628));
    layer1_outputs(6160) <= layer0_outputs(9945);
    layer1_outputs(6161) <= (layer0_outputs(3869)) or (layer0_outputs(224));
    layer1_outputs(6162) <= (layer0_outputs(8238)) and (layer0_outputs(2569));
    layer1_outputs(6163) <= not(layer0_outputs(22)) or (layer0_outputs(4953));
    layer1_outputs(6164) <= layer0_outputs(1966);
    layer1_outputs(6165) <= (layer0_outputs(2284)) and not (layer0_outputs(5441));
    layer1_outputs(6166) <= (layer0_outputs(3667)) and (layer0_outputs(6225));
    layer1_outputs(6167) <= (layer0_outputs(1624)) or (layer0_outputs(7853));
    layer1_outputs(6168) <= not(layer0_outputs(4902)) or (layer0_outputs(10039));
    layer1_outputs(6169) <= not(layer0_outputs(7603));
    layer1_outputs(6170) <= not((layer0_outputs(9506)) or (layer0_outputs(7252)));
    layer1_outputs(6171) <= not((layer0_outputs(5479)) and (layer0_outputs(9575)));
    layer1_outputs(6172) <= not(layer0_outputs(3688)) or (layer0_outputs(6692));
    layer1_outputs(6173) <= (layer0_outputs(4137)) and not (layer0_outputs(6248));
    layer1_outputs(6174) <= (layer0_outputs(3240)) or (layer0_outputs(1206));
    layer1_outputs(6175) <= (layer0_outputs(3412)) and not (layer0_outputs(3320));
    layer1_outputs(6176) <= not((layer0_outputs(2259)) or (layer0_outputs(619)));
    layer1_outputs(6177) <= not(layer0_outputs(8537)) or (layer0_outputs(2419));
    layer1_outputs(6178) <= not((layer0_outputs(4256)) and (layer0_outputs(8261)));
    layer1_outputs(6179) <= not(layer0_outputs(1081));
    layer1_outputs(6180) <= layer0_outputs(4471);
    layer1_outputs(6181) <= not((layer0_outputs(2114)) and (layer0_outputs(31)));
    layer1_outputs(6182) <= not((layer0_outputs(3161)) xor (layer0_outputs(8799)));
    layer1_outputs(6183) <= not((layer0_outputs(1251)) or (layer0_outputs(3276)));
    layer1_outputs(6184) <= not(layer0_outputs(6372)) or (layer0_outputs(2651));
    layer1_outputs(6185) <= '0';
    layer1_outputs(6186) <= '1';
    layer1_outputs(6187) <= not(layer0_outputs(3543)) or (layer0_outputs(8202));
    layer1_outputs(6188) <= (layer0_outputs(9726)) and not (layer0_outputs(7385));
    layer1_outputs(6189) <= layer0_outputs(4914);
    layer1_outputs(6190) <= '1';
    layer1_outputs(6191) <= not(layer0_outputs(7945));
    layer1_outputs(6192) <= layer0_outputs(8086);
    layer1_outputs(6193) <= not((layer0_outputs(7818)) xor (layer0_outputs(5870)));
    layer1_outputs(6194) <= not((layer0_outputs(3845)) xor (layer0_outputs(9279)));
    layer1_outputs(6195) <= layer0_outputs(3535);
    layer1_outputs(6196) <= not((layer0_outputs(6581)) or (layer0_outputs(41)));
    layer1_outputs(6197) <= not(layer0_outputs(414));
    layer1_outputs(6198) <= (layer0_outputs(996)) and (layer0_outputs(3900));
    layer1_outputs(6199) <= (layer0_outputs(4186)) and not (layer0_outputs(2102));
    layer1_outputs(6200) <= not((layer0_outputs(84)) and (layer0_outputs(1537)));
    layer1_outputs(6201) <= (layer0_outputs(918)) and not (layer0_outputs(2652));
    layer1_outputs(6202) <= not(layer0_outputs(4861));
    layer1_outputs(6203) <= (layer0_outputs(7766)) or (layer0_outputs(7987));
    layer1_outputs(6204) <= '1';
    layer1_outputs(6205) <= layer0_outputs(8437);
    layer1_outputs(6206) <= not(layer0_outputs(9332));
    layer1_outputs(6207) <= not(layer0_outputs(6716)) or (layer0_outputs(8928));
    layer1_outputs(6208) <= '0';
    layer1_outputs(6209) <= (layer0_outputs(4263)) or (layer0_outputs(2271));
    layer1_outputs(6210) <= not(layer0_outputs(6301));
    layer1_outputs(6211) <= (layer0_outputs(5304)) and not (layer0_outputs(8843));
    layer1_outputs(6212) <= layer0_outputs(9331);
    layer1_outputs(6213) <= layer0_outputs(3435);
    layer1_outputs(6214) <= not(layer0_outputs(1663));
    layer1_outputs(6215) <= layer0_outputs(897);
    layer1_outputs(6216) <= (layer0_outputs(4818)) and (layer0_outputs(9485));
    layer1_outputs(6217) <= not(layer0_outputs(6745)) or (layer0_outputs(8065));
    layer1_outputs(6218) <= (layer0_outputs(7590)) or (layer0_outputs(7705));
    layer1_outputs(6219) <= not(layer0_outputs(3599));
    layer1_outputs(6220) <= (layer0_outputs(7799)) and not (layer0_outputs(10066));
    layer1_outputs(6221) <= not((layer0_outputs(9271)) and (layer0_outputs(3400)));
    layer1_outputs(6222) <= not(layer0_outputs(8027));
    layer1_outputs(6223) <= (layer0_outputs(7927)) xor (layer0_outputs(9808));
    layer1_outputs(6224) <= not(layer0_outputs(160));
    layer1_outputs(6225) <= not(layer0_outputs(251)) or (layer0_outputs(5623));
    layer1_outputs(6226) <= layer0_outputs(9606);
    layer1_outputs(6227) <= layer0_outputs(912);
    layer1_outputs(6228) <= layer0_outputs(2811);
    layer1_outputs(6229) <= layer0_outputs(1753);
    layer1_outputs(6230) <= not(layer0_outputs(4471));
    layer1_outputs(6231) <= not((layer0_outputs(1886)) and (layer0_outputs(9821)));
    layer1_outputs(6232) <= not(layer0_outputs(5935)) or (layer0_outputs(3223));
    layer1_outputs(6233) <= not(layer0_outputs(726));
    layer1_outputs(6234) <= not(layer0_outputs(8314)) or (layer0_outputs(8313));
    layer1_outputs(6235) <= (layer0_outputs(5176)) and not (layer0_outputs(3301));
    layer1_outputs(6236) <= (layer0_outputs(7924)) and not (layer0_outputs(9981));
    layer1_outputs(6237) <= (layer0_outputs(8360)) and not (layer0_outputs(3335));
    layer1_outputs(6238) <= not(layer0_outputs(9467)) or (layer0_outputs(4313));
    layer1_outputs(6239) <= layer0_outputs(7522);
    layer1_outputs(6240) <= layer0_outputs(7828);
    layer1_outputs(6241) <= not(layer0_outputs(354));
    layer1_outputs(6242) <= not(layer0_outputs(5864)) or (layer0_outputs(1866));
    layer1_outputs(6243) <= not((layer0_outputs(7218)) and (layer0_outputs(3143)));
    layer1_outputs(6244) <= not((layer0_outputs(1545)) or (layer0_outputs(1282)));
    layer1_outputs(6245) <= layer0_outputs(1381);
    layer1_outputs(6246) <= not(layer0_outputs(2803)) or (layer0_outputs(4623));
    layer1_outputs(6247) <= '0';
    layer1_outputs(6248) <= not(layer0_outputs(7295)) or (layer0_outputs(3870));
    layer1_outputs(6249) <= (layer0_outputs(5967)) and (layer0_outputs(5389));
    layer1_outputs(6250) <= layer0_outputs(5019);
    layer1_outputs(6251) <= layer0_outputs(3536);
    layer1_outputs(6252) <= not((layer0_outputs(5509)) and (layer0_outputs(64)));
    layer1_outputs(6253) <= (layer0_outputs(7404)) or (layer0_outputs(4926));
    layer1_outputs(6254) <= layer0_outputs(6326);
    layer1_outputs(6255) <= not((layer0_outputs(2871)) and (layer0_outputs(386)));
    layer1_outputs(6256) <= not(layer0_outputs(10205)) or (layer0_outputs(2911));
    layer1_outputs(6257) <= layer0_outputs(4179);
    layer1_outputs(6258) <= not((layer0_outputs(5162)) or (layer0_outputs(9840)));
    layer1_outputs(6259) <= not(layer0_outputs(4764));
    layer1_outputs(6260) <= not((layer0_outputs(1864)) or (layer0_outputs(2120)));
    layer1_outputs(6261) <= (layer0_outputs(377)) xor (layer0_outputs(1257));
    layer1_outputs(6262) <= not(layer0_outputs(8374)) or (layer0_outputs(4901));
    layer1_outputs(6263) <= not(layer0_outputs(8245)) or (layer0_outputs(8826));
    layer1_outputs(6264) <= '1';
    layer1_outputs(6265) <= not((layer0_outputs(1423)) and (layer0_outputs(5641)));
    layer1_outputs(6266) <= '0';
    layer1_outputs(6267) <= layer0_outputs(9308);
    layer1_outputs(6268) <= layer0_outputs(3436);
    layer1_outputs(6269) <= '0';
    layer1_outputs(6270) <= not((layer0_outputs(8469)) and (layer0_outputs(4613)));
    layer1_outputs(6271) <= not(layer0_outputs(9778));
    layer1_outputs(6272) <= not(layer0_outputs(416));
    layer1_outputs(6273) <= not((layer0_outputs(4731)) and (layer0_outputs(6013)));
    layer1_outputs(6274) <= not((layer0_outputs(3769)) xor (layer0_outputs(7965)));
    layer1_outputs(6275) <= not((layer0_outputs(6609)) xor (layer0_outputs(8766)));
    layer1_outputs(6276) <= not(layer0_outputs(9874));
    layer1_outputs(6277) <= not(layer0_outputs(2735)) or (layer0_outputs(3960));
    layer1_outputs(6278) <= not(layer0_outputs(4055));
    layer1_outputs(6279) <= not(layer0_outputs(9888));
    layer1_outputs(6280) <= (layer0_outputs(2793)) or (layer0_outputs(2318));
    layer1_outputs(6281) <= '0';
    layer1_outputs(6282) <= (layer0_outputs(9459)) and not (layer0_outputs(1497));
    layer1_outputs(6283) <= (layer0_outputs(3648)) and (layer0_outputs(10106));
    layer1_outputs(6284) <= (layer0_outputs(3322)) and not (layer0_outputs(1379));
    layer1_outputs(6285) <= not(layer0_outputs(5890)) or (layer0_outputs(5318));
    layer1_outputs(6286) <= not((layer0_outputs(2113)) and (layer0_outputs(8374)));
    layer1_outputs(6287) <= not((layer0_outputs(7241)) or (layer0_outputs(1563)));
    layer1_outputs(6288) <= not(layer0_outputs(7265));
    layer1_outputs(6289) <= '1';
    layer1_outputs(6290) <= layer0_outputs(4516);
    layer1_outputs(6291) <= not(layer0_outputs(4234)) or (layer0_outputs(7597));
    layer1_outputs(6292) <= not((layer0_outputs(5218)) and (layer0_outputs(6209)));
    layer1_outputs(6293) <= not(layer0_outputs(4582)) or (layer0_outputs(811));
    layer1_outputs(6294) <= not((layer0_outputs(5749)) or (layer0_outputs(5904)));
    layer1_outputs(6295) <= not((layer0_outputs(2073)) and (layer0_outputs(4109)));
    layer1_outputs(6296) <= (layer0_outputs(4678)) or (layer0_outputs(3909));
    layer1_outputs(6297) <= not((layer0_outputs(1731)) and (layer0_outputs(5958)));
    layer1_outputs(6298) <= not(layer0_outputs(2005)) or (layer0_outputs(930));
    layer1_outputs(6299) <= not((layer0_outputs(2637)) or (layer0_outputs(2646)));
    layer1_outputs(6300) <= not(layer0_outputs(9510)) or (layer0_outputs(9826));
    layer1_outputs(6301) <= (layer0_outputs(8912)) and not (layer0_outputs(2105));
    layer1_outputs(6302) <= (layer0_outputs(623)) or (layer0_outputs(3966));
    layer1_outputs(6303) <= (layer0_outputs(1799)) and not (layer0_outputs(8948));
    layer1_outputs(6304) <= not(layer0_outputs(7638)) or (layer0_outputs(10186));
    layer1_outputs(6305) <= layer0_outputs(1497);
    layer1_outputs(6306) <= (layer0_outputs(956)) xor (layer0_outputs(447));
    layer1_outputs(6307) <= (layer0_outputs(4038)) xor (layer0_outputs(8590));
    layer1_outputs(6308) <= not(layer0_outputs(1042));
    layer1_outputs(6309) <= not(layer0_outputs(9627));
    layer1_outputs(6310) <= (layer0_outputs(9131)) xor (layer0_outputs(6705));
    layer1_outputs(6311) <= not(layer0_outputs(7190));
    layer1_outputs(6312) <= '1';
    layer1_outputs(6313) <= layer0_outputs(9976);
    layer1_outputs(6314) <= (layer0_outputs(9058)) and (layer0_outputs(8031));
    layer1_outputs(6315) <= '1';
    layer1_outputs(6316) <= not((layer0_outputs(3287)) or (layer0_outputs(2405)));
    layer1_outputs(6317) <= layer0_outputs(6341);
    layer1_outputs(6318) <= '0';
    layer1_outputs(6319) <= not(layer0_outputs(5408)) or (layer0_outputs(1345));
    layer1_outputs(6320) <= not(layer0_outputs(8517)) or (layer0_outputs(4840));
    layer1_outputs(6321) <= (layer0_outputs(6422)) or (layer0_outputs(5235));
    layer1_outputs(6322) <= not(layer0_outputs(10127));
    layer1_outputs(6323) <= (layer0_outputs(7405)) and not (layer0_outputs(6072));
    layer1_outputs(6324) <= not(layer0_outputs(7709));
    layer1_outputs(6325) <= layer0_outputs(1722);
    layer1_outputs(6326) <= '0';
    layer1_outputs(6327) <= not(layer0_outputs(3422));
    layer1_outputs(6328) <= (layer0_outputs(8853)) and not (layer0_outputs(3463));
    layer1_outputs(6329) <= not(layer0_outputs(4106));
    layer1_outputs(6330) <= '0';
    layer1_outputs(6331) <= not(layer0_outputs(5878));
    layer1_outputs(6332) <= not((layer0_outputs(6123)) or (layer0_outputs(7176)));
    layer1_outputs(6333) <= not(layer0_outputs(4973));
    layer1_outputs(6334) <= (layer0_outputs(5891)) and not (layer0_outputs(1688));
    layer1_outputs(6335) <= not((layer0_outputs(4390)) and (layer0_outputs(8551)));
    layer1_outputs(6336) <= not(layer0_outputs(748));
    layer1_outputs(6337) <= not((layer0_outputs(4874)) or (layer0_outputs(2532)));
    layer1_outputs(6338) <= not(layer0_outputs(1504));
    layer1_outputs(6339) <= (layer0_outputs(6795)) or (layer0_outputs(8197));
    layer1_outputs(6340) <= not(layer0_outputs(264)) or (layer0_outputs(9000));
    layer1_outputs(6341) <= not(layer0_outputs(5729));
    layer1_outputs(6342) <= not(layer0_outputs(9340));
    layer1_outputs(6343) <= layer0_outputs(3635);
    layer1_outputs(6344) <= (layer0_outputs(2235)) xor (layer0_outputs(4883));
    layer1_outputs(6345) <= layer0_outputs(662);
    layer1_outputs(6346) <= not((layer0_outputs(5991)) xor (layer0_outputs(4504)));
    layer1_outputs(6347) <= (layer0_outputs(2361)) xor (layer0_outputs(8847));
    layer1_outputs(6348) <= not((layer0_outputs(4332)) and (layer0_outputs(1630)));
    layer1_outputs(6349) <= not((layer0_outputs(9101)) and (layer0_outputs(2350)));
    layer1_outputs(6350) <= not(layer0_outputs(131));
    layer1_outputs(6351) <= (layer0_outputs(8712)) and (layer0_outputs(2855));
    layer1_outputs(6352) <= '0';
    layer1_outputs(6353) <= not((layer0_outputs(2134)) and (layer0_outputs(1307)));
    layer1_outputs(6354) <= layer0_outputs(310);
    layer1_outputs(6355) <= not(layer0_outputs(9072)) or (layer0_outputs(146));
    layer1_outputs(6356) <= (layer0_outputs(5922)) and not (layer0_outputs(1731));
    layer1_outputs(6357) <= not(layer0_outputs(2516));
    layer1_outputs(6358) <= not(layer0_outputs(7513));
    layer1_outputs(6359) <= (layer0_outputs(863)) and (layer0_outputs(1175));
    layer1_outputs(6360) <= not((layer0_outputs(7664)) and (layer0_outputs(3723)));
    layer1_outputs(6361) <= not((layer0_outputs(1971)) and (layer0_outputs(479)));
    layer1_outputs(6362) <= not(layer0_outputs(2043)) or (layer0_outputs(9461));
    layer1_outputs(6363) <= (layer0_outputs(7548)) and not (layer0_outputs(6580));
    layer1_outputs(6364) <= (layer0_outputs(415)) xor (layer0_outputs(2931));
    layer1_outputs(6365) <= layer0_outputs(5590);
    layer1_outputs(6366) <= not(layer0_outputs(7745));
    layer1_outputs(6367) <= layer0_outputs(7733);
    layer1_outputs(6368) <= not(layer0_outputs(8677));
    layer1_outputs(6369) <= layer0_outputs(8384);
    layer1_outputs(6370) <= layer0_outputs(7814);
    layer1_outputs(6371) <= layer0_outputs(4446);
    layer1_outputs(6372) <= (layer0_outputs(6090)) or (layer0_outputs(1365));
    layer1_outputs(6373) <= not(layer0_outputs(5128)) or (layer0_outputs(2563));
    layer1_outputs(6374) <= not(layer0_outputs(3554)) or (layer0_outputs(9226));
    layer1_outputs(6375) <= layer0_outputs(7015);
    layer1_outputs(6376) <= (layer0_outputs(7382)) and not (layer0_outputs(7094));
    layer1_outputs(6377) <= not(layer0_outputs(4839)) or (layer0_outputs(6744));
    layer1_outputs(6378) <= '0';
    layer1_outputs(6379) <= not(layer0_outputs(4273));
    layer1_outputs(6380) <= not(layer0_outputs(6840));
    layer1_outputs(6381) <= not(layer0_outputs(764));
    layer1_outputs(6382) <= not((layer0_outputs(9378)) or (layer0_outputs(4522)));
    layer1_outputs(6383) <= layer0_outputs(5932);
    layer1_outputs(6384) <= (layer0_outputs(5969)) and not (layer0_outputs(3921));
    layer1_outputs(6385) <= layer0_outputs(10215);
    layer1_outputs(6386) <= (layer0_outputs(9655)) xor (layer0_outputs(9644));
    layer1_outputs(6387) <= (layer0_outputs(5554)) xor (layer0_outputs(8472));
    layer1_outputs(6388) <= not(layer0_outputs(9390)) or (layer0_outputs(7511));
    layer1_outputs(6389) <= not(layer0_outputs(5065)) or (layer0_outputs(971));
    layer1_outputs(6390) <= (layer0_outputs(7436)) and not (layer0_outputs(1782));
    layer1_outputs(6391) <= layer0_outputs(6947);
    layer1_outputs(6392) <= (layer0_outputs(7148)) and not (layer0_outputs(1757));
    layer1_outputs(6393) <= not(layer0_outputs(7302));
    layer1_outputs(6394) <= not((layer0_outputs(2476)) or (layer0_outputs(3497)));
    layer1_outputs(6395) <= '1';
    layer1_outputs(6396) <= (layer0_outputs(2022)) or (layer0_outputs(6217));
    layer1_outputs(6397) <= '0';
    layer1_outputs(6398) <= layer0_outputs(1833);
    layer1_outputs(6399) <= not(layer0_outputs(4998));
    layer1_outputs(6400) <= not(layer0_outputs(3446));
    layer1_outputs(6401) <= layer0_outputs(4874);
    layer1_outputs(6402) <= layer0_outputs(8104);
    layer1_outputs(6403) <= not(layer0_outputs(8408));
    layer1_outputs(6404) <= '0';
    layer1_outputs(6405) <= not(layer0_outputs(6444));
    layer1_outputs(6406) <= not((layer0_outputs(4502)) and (layer0_outputs(597)));
    layer1_outputs(6407) <= not((layer0_outputs(1162)) or (layer0_outputs(5372)));
    layer1_outputs(6408) <= (layer0_outputs(1285)) xor (layer0_outputs(3848));
    layer1_outputs(6409) <= not((layer0_outputs(5872)) or (layer0_outputs(1049)));
    layer1_outputs(6410) <= not(layer0_outputs(762));
    layer1_outputs(6411) <= (layer0_outputs(9627)) or (layer0_outputs(9050));
    layer1_outputs(6412) <= not((layer0_outputs(1038)) or (layer0_outputs(2)));
    layer1_outputs(6413) <= not(layer0_outputs(7246)) or (layer0_outputs(6465));
    layer1_outputs(6414) <= not(layer0_outputs(4128)) or (layer0_outputs(2553));
    layer1_outputs(6415) <= (layer0_outputs(5769)) xor (layer0_outputs(5696));
    layer1_outputs(6416) <= layer0_outputs(9208);
    layer1_outputs(6417) <= not(layer0_outputs(7600)) or (layer0_outputs(695));
    layer1_outputs(6418) <= layer0_outputs(5481);
    layer1_outputs(6419) <= (layer0_outputs(9605)) or (layer0_outputs(2542));
    layer1_outputs(6420) <= '1';
    layer1_outputs(6421) <= layer0_outputs(5596);
    layer1_outputs(6422) <= (layer0_outputs(6833)) or (layer0_outputs(1729));
    layer1_outputs(6423) <= (layer0_outputs(572)) and not (layer0_outputs(693));
    layer1_outputs(6424) <= not(layer0_outputs(7216)) or (layer0_outputs(7354));
    layer1_outputs(6425) <= layer0_outputs(9118);
    layer1_outputs(6426) <= not(layer0_outputs(6543)) or (layer0_outputs(6421));
    layer1_outputs(6427) <= (layer0_outputs(1201)) and not (layer0_outputs(5577));
    layer1_outputs(6428) <= (layer0_outputs(8769)) xor (layer0_outputs(6534));
    layer1_outputs(6429) <= not(layer0_outputs(509));
    layer1_outputs(6430) <= '1';
    layer1_outputs(6431) <= (layer0_outputs(6279)) and not (layer0_outputs(9915));
    layer1_outputs(6432) <= not((layer0_outputs(2872)) or (layer0_outputs(3701)));
    layer1_outputs(6433) <= not(layer0_outputs(804)) or (layer0_outputs(4605));
    layer1_outputs(6434) <= layer0_outputs(4015);
    layer1_outputs(6435) <= not(layer0_outputs(4820)) or (layer0_outputs(4079));
    layer1_outputs(6436) <= (layer0_outputs(765)) or (layer0_outputs(9330));
    layer1_outputs(6437) <= (layer0_outputs(5753)) and not (layer0_outputs(6414));
    layer1_outputs(6438) <= not(layer0_outputs(8236));
    layer1_outputs(6439) <= (layer0_outputs(3515)) and not (layer0_outputs(4762));
    layer1_outputs(6440) <= not(layer0_outputs(7555));
    layer1_outputs(6441) <= not(layer0_outputs(9422));
    layer1_outputs(6442) <= layer0_outputs(8662);
    layer1_outputs(6443) <= not(layer0_outputs(7340));
    layer1_outputs(6444) <= '0';
    layer1_outputs(6445) <= not(layer0_outputs(1319)) or (layer0_outputs(8660));
    layer1_outputs(6446) <= not((layer0_outputs(10068)) and (layer0_outputs(407)));
    layer1_outputs(6447) <= (layer0_outputs(8678)) and (layer0_outputs(236));
    layer1_outputs(6448) <= not(layer0_outputs(210));
    layer1_outputs(6449) <= '1';
    layer1_outputs(6450) <= not(layer0_outputs(1396)) or (layer0_outputs(1978));
    layer1_outputs(6451) <= (layer0_outputs(120)) and (layer0_outputs(3249));
    layer1_outputs(6452) <= layer0_outputs(2748);
    layer1_outputs(6453) <= (layer0_outputs(2806)) or (layer0_outputs(5242));
    layer1_outputs(6454) <= (layer0_outputs(5204)) and not (layer0_outputs(3855));
    layer1_outputs(6455) <= (layer0_outputs(4876)) and not (layer0_outputs(1095));
    layer1_outputs(6456) <= not(layer0_outputs(8686));
    layer1_outputs(6457) <= (layer0_outputs(1077)) and (layer0_outputs(7122));
    layer1_outputs(6458) <= not((layer0_outputs(3823)) and (layer0_outputs(4868)));
    layer1_outputs(6459) <= layer0_outputs(6550);
    layer1_outputs(6460) <= not(layer0_outputs(4816)) or (layer0_outputs(2740));
    layer1_outputs(6461) <= (layer0_outputs(9781)) and (layer0_outputs(2942));
    layer1_outputs(6462) <= not(layer0_outputs(845)) or (layer0_outputs(2236));
    layer1_outputs(6463) <= not(layer0_outputs(75));
    layer1_outputs(6464) <= layer0_outputs(7572);
    layer1_outputs(6465) <= not(layer0_outputs(9289));
    layer1_outputs(6466) <= not(layer0_outputs(8895));
    layer1_outputs(6467) <= (layer0_outputs(4571)) xor (layer0_outputs(2659));
    layer1_outputs(6468) <= not((layer0_outputs(6702)) or (layer0_outputs(2670)));
    layer1_outputs(6469) <= not(layer0_outputs(9446)) or (layer0_outputs(4118));
    layer1_outputs(6470) <= layer0_outputs(308);
    layer1_outputs(6471) <= (layer0_outputs(10233)) or (layer0_outputs(3269));
    layer1_outputs(6472) <= not(layer0_outputs(4562));
    layer1_outputs(6473) <= (layer0_outputs(7432)) and not (layer0_outputs(7024));
    layer1_outputs(6474) <= (layer0_outputs(679)) and not (layer0_outputs(1857));
    layer1_outputs(6475) <= not(layer0_outputs(335));
    layer1_outputs(6476) <= not(layer0_outputs(4964));
    layer1_outputs(6477) <= not((layer0_outputs(8336)) and (layer0_outputs(3574)));
    layer1_outputs(6478) <= '0';
    layer1_outputs(6479) <= layer0_outputs(4044);
    layer1_outputs(6480) <= not(layer0_outputs(101)) or (layer0_outputs(9594));
    layer1_outputs(6481) <= not(layer0_outputs(6044)) or (layer0_outputs(7637));
    layer1_outputs(6482) <= not(layer0_outputs(3027));
    layer1_outputs(6483) <= (layer0_outputs(4664)) and (layer0_outputs(2617));
    layer1_outputs(6484) <= (layer0_outputs(4839)) and not (layer0_outputs(173));
    layer1_outputs(6485) <= (layer0_outputs(10084)) xor (layer0_outputs(5010));
    layer1_outputs(6486) <= (layer0_outputs(5544)) or (layer0_outputs(6175));
    layer1_outputs(6487) <= '1';
    layer1_outputs(6488) <= not((layer0_outputs(2086)) xor (layer0_outputs(203)));
    layer1_outputs(6489) <= not(layer0_outputs(4204));
    layer1_outputs(6490) <= layer0_outputs(6566);
    layer1_outputs(6491) <= (layer0_outputs(10107)) and (layer0_outputs(10060));
    layer1_outputs(6492) <= (layer0_outputs(7744)) xor (layer0_outputs(5037));
    layer1_outputs(6493) <= not(layer0_outputs(3765));
    layer1_outputs(6494) <= '0';
    layer1_outputs(6495) <= (layer0_outputs(9304)) and not (layer0_outputs(7417));
    layer1_outputs(6496) <= not(layer0_outputs(2772)) or (layer0_outputs(4976));
    layer1_outputs(6497) <= not(layer0_outputs(9331));
    layer1_outputs(6498) <= layer0_outputs(9630);
    layer1_outputs(6499) <= not(layer0_outputs(4957));
    layer1_outputs(6500) <= not(layer0_outputs(997));
    layer1_outputs(6501) <= (layer0_outputs(1699)) and (layer0_outputs(8782));
    layer1_outputs(6502) <= (layer0_outputs(1088)) and not (layer0_outputs(1602));
    layer1_outputs(6503) <= (layer0_outputs(7846)) xor (layer0_outputs(2189));
    layer1_outputs(6504) <= not(layer0_outputs(266)) or (layer0_outputs(2315));
    layer1_outputs(6505) <= (layer0_outputs(6274)) and (layer0_outputs(6624));
    layer1_outputs(6506) <= not(layer0_outputs(3355)) or (layer0_outputs(7551));
    layer1_outputs(6507) <= not(layer0_outputs(849));
    layer1_outputs(6508) <= '0';
    layer1_outputs(6509) <= not(layer0_outputs(5089));
    layer1_outputs(6510) <= (layer0_outputs(9702)) and not (layer0_outputs(2319));
    layer1_outputs(6511) <= '1';
    layer1_outputs(6512) <= not((layer0_outputs(9828)) xor (layer0_outputs(3670)));
    layer1_outputs(6513) <= not(layer0_outputs(6709)) or (layer0_outputs(10037));
    layer1_outputs(6514) <= (layer0_outputs(6302)) and (layer0_outputs(221));
    layer1_outputs(6515) <= not((layer0_outputs(2851)) and (layer0_outputs(5650)));
    layer1_outputs(6516) <= layer0_outputs(10212);
    layer1_outputs(6517) <= (layer0_outputs(2794)) and not (layer0_outputs(6441));
    layer1_outputs(6518) <= not(layer0_outputs(4652));
    layer1_outputs(6519) <= (layer0_outputs(8562)) and (layer0_outputs(313));
    layer1_outputs(6520) <= (layer0_outputs(7061)) and not (layer0_outputs(10146));
    layer1_outputs(6521) <= not(layer0_outputs(5981));
    layer1_outputs(6522) <= not(layer0_outputs(3761));
    layer1_outputs(6523) <= '1';
    layer1_outputs(6524) <= not(layer0_outputs(6919));
    layer1_outputs(6525) <= layer0_outputs(1366);
    layer1_outputs(6526) <= (layer0_outputs(2521)) and (layer0_outputs(1432));
    layer1_outputs(6527) <= not(layer0_outputs(5160));
    layer1_outputs(6528) <= not(layer0_outputs(3887)) or (layer0_outputs(3305));
    layer1_outputs(6529) <= not((layer0_outputs(7631)) and (layer0_outputs(4982)));
    layer1_outputs(6530) <= layer0_outputs(2043);
    layer1_outputs(6531) <= not((layer0_outputs(5126)) and (layer0_outputs(8819)));
    layer1_outputs(6532) <= not((layer0_outputs(1972)) or (layer0_outputs(1860)));
    layer1_outputs(6533) <= (layer0_outputs(5024)) xor (layer0_outputs(9233));
    layer1_outputs(6534) <= (layer0_outputs(10091)) and not (layer0_outputs(4403));
    layer1_outputs(6535) <= not((layer0_outputs(95)) and (layer0_outputs(3102)));
    layer1_outputs(6536) <= not(layer0_outputs(1959));
    layer1_outputs(6537) <= not(layer0_outputs(3424));
    layer1_outputs(6538) <= (layer0_outputs(4244)) and not (layer0_outputs(7856));
    layer1_outputs(6539) <= '0';
    layer1_outputs(6540) <= '1';
    layer1_outputs(6541) <= not(layer0_outputs(9565)) or (layer0_outputs(42));
    layer1_outputs(6542) <= not(layer0_outputs(202));
    layer1_outputs(6543) <= layer0_outputs(2125);
    layer1_outputs(6544) <= layer0_outputs(9430);
    layer1_outputs(6545) <= (layer0_outputs(4653)) and not (layer0_outputs(9509));
    layer1_outputs(6546) <= not((layer0_outputs(4964)) and (layer0_outputs(4521)));
    layer1_outputs(6547) <= '0';
    layer1_outputs(6548) <= (layer0_outputs(5088)) or (layer0_outputs(4808));
    layer1_outputs(6549) <= (layer0_outputs(5316)) xor (layer0_outputs(4243));
    layer1_outputs(6550) <= not((layer0_outputs(3379)) xor (layer0_outputs(1831)));
    layer1_outputs(6551) <= not((layer0_outputs(5198)) and (layer0_outputs(3690)));
    layer1_outputs(6552) <= not((layer0_outputs(1042)) or (layer0_outputs(3437)));
    layer1_outputs(6553) <= not((layer0_outputs(4095)) and (layer0_outputs(10173)));
    layer1_outputs(6554) <= not(layer0_outputs(10220)) or (layer0_outputs(1656));
    layer1_outputs(6555) <= layer0_outputs(5539);
    layer1_outputs(6556) <= not(layer0_outputs(2218));
    layer1_outputs(6557) <= not((layer0_outputs(432)) xor (layer0_outputs(7476)));
    layer1_outputs(6558) <= layer0_outputs(5630);
    layer1_outputs(6559) <= (layer0_outputs(2453)) and (layer0_outputs(8961));
    layer1_outputs(6560) <= not((layer0_outputs(967)) xor (layer0_outputs(10087)));
    layer1_outputs(6561) <= not(layer0_outputs(7335));
    layer1_outputs(6562) <= not(layer0_outputs(7921));
    layer1_outputs(6563) <= layer0_outputs(653);
    layer1_outputs(6564) <= not((layer0_outputs(6608)) and (layer0_outputs(8582)));
    layer1_outputs(6565) <= not((layer0_outputs(1691)) or (layer0_outputs(3876)));
    layer1_outputs(6566) <= (layer0_outputs(4660)) and not (layer0_outputs(2400));
    layer1_outputs(6567) <= not(layer0_outputs(9438));
    layer1_outputs(6568) <= (layer0_outputs(2825)) and (layer0_outputs(4520));
    layer1_outputs(6569) <= '1';
    layer1_outputs(6570) <= not(layer0_outputs(419));
    layer1_outputs(6571) <= not(layer0_outputs(5185));
    layer1_outputs(6572) <= (layer0_outputs(4576)) or (layer0_outputs(1223));
    layer1_outputs(6573) <= (layer0_outputs(8129)) and not (layer0_outputs(9435));
    layer1_outputs(6574) <= layer0_outputs(8748);
    layer1_outputs(6575) <= not((layer0_outputs(9077)) or (layer0_outputs(6602)));
    layer1_outputs(6576) <= not((layer0_outputs(3586)) and (layer0_outputs(9082)));
    layer1_outputs(6577) <= layer0_outputs(8376);
    layer1_outputs(6578) <= not(layer0_outputs(3579));
    layer1_outputs(6579) <= (layer0_outputs(4483)) and (layer0_outputs(2832));
    layer1_outputs(6580) <= not(layer0_outputs(9402));
    layer1_outputs(6581) <= not(layer0_outputs(9811));
    layer1_outputs(6582) <= (layer0_outputs(4869)) and (layer0_outputs(1686));
    layer1_outputs(6583) <= not((layer0_outputs(1899)) and (layer0_outputs(98)));
    layer1_outputs(6584) <= not(layer0_outputs(6143)) or (layer0_outputs(2046));
    layer1_outputs(6585) <= (layer0_outputs(1257)) and not (layer0_outputs(5102));
    layer1_outputs(6586) <= layer0_outputs(10172);
    layer1_outputs(6587) <= not(layer0_outputs(3914));
    layer1_outputs(6588) <= layer0_outputs(6399);
    layer1_outputs(6589) <= '1';
    layer1_outputs(6590) <= layer0_outputs(8642);
    layer1_outputs(6591) <= layer0_outputs(8845);
    layer1_outputs(6592) <= not(layer0_outputs(4658)) or (layer0_outputs(5701));
    layer1_outputs(6593) <= (layer0_outputs(2981)) and (layer0_outputs(847));
    layer1_outputs(6594) <= layer0_outputs(2311);
    layer1_outputs(6595) <= not(layer0_outputs(6129));
    layer1_outputs(6596) <= (layer0_outputs(5832)) or (layer0_outputs(6929));
    layer1_outputs(6597) <= not((layer0_outputs(5010)) or (layer0_outputs(2188)));
    layer1_outputs(6598) <= not((layer0_outputs(9562)) and (layer0_outputs(3821)));
    layer1_outputs(6599) <= not((layer0_outputs(5970)) and (layer0_outputs(9223)));
    layer1_outputs(6600) <= not(layer0_outputs(10012)) or (layer0_outputs(1300));
    layer1_outputs(6601) <= not((layer0_outputs(7023)) xor (layer0_outputs(6623)));
    layer1_outputs(6602) <= not(layer0_outputs(5189));
    layer1_outputs(6603) <= not(layer0_outputs(3447)) or (layer0_outputs(148));
    layer1_outputs(6604) <= not((layer0_outputs(4036)) or (layer0_outputs(1297)));
    layer1_outputs(6605) <= not((layer0_outputs(2398)) and (layer0_outputs(7319)));
    layer1_outputs(6606) <= not((layer0_outputs(8767)) and (layer0_outputs(2197)));
    layer1_outputs(6607) <= not((layer0_outputs(9784)) and (layer0_outputs(5064)));
    layer1_outputs(6608) <= (layer0_outputs(6447)) and not (layer0_outputs(2204));
    layer1_outputs(6609) <= not((layer0_outputs(3638)) xor (layer0_outputs(4125)));
    layer1_outputs(6610) <= not(layer0_outputs(6673)) or (layer0_outputs(8500));
    layer1_outputs(6611) <= (layer0_outputs(1064)) and not (layer0_outputs(8497));
    layer1_outputs(6612) <= (layer0_outputs(3977)) and not (layer0_outputs(6998));
    layer1_outputs(6613) <= not(layer0_outputs(1376)) or (layer0_outputs(1037));
    layer1_outputs(6614) <= '1';
    layer1_outputs(6615) <= not((layer0_outputs(7114)) xor (layer0_outputs(9136)));
    layer1_outputs(6616) <= not((layer0_outputs(6880)) xor (layer0_outputs(1896)));
    layer1_outputs(6617) <= not((layer0_outputs(5938)) and (layer0_outputs(1853)));
    layer1_outputs(6618) <= (layer0_outputs(9685)) and not (layer0_outputs(548));
    layer1_outputs(6619) <= (layer0_outputs(9123)) or (layer0_outputs(1227));
    layer1_outputs(6620) <= layer0_outputs(4203);
    layer1_outputs(6621) <= not((layer0_outputs(939)) and (layer0_outputs(9768)));
    layer1_outputs(6622) <= not(layer0_outputs(9332));
    layer1_outputs(6623) <= not(layer0_outputs(282));
    layer1_outputs(6624) <= (layer0_outputs(2771)) and not (layer0_outputs(5948));
    layer1_outputs(6625) <= not(layer0_outputs(3182)) or (layer0_outputs(1337));
    layer1_outputs(6626) <= not(layer0_outputs(3561));
    layer1_outputs(6627) <= layer0_outputs(7140);
    layer1_outputs(6628) <= (layer0_outputs(1149)) xor (layer0_outputs(9228));
    layer1_outputs(6629) <= not(layer0_outputs(9451));
    layer1_outputs(6630) <= (layer0_outputs(1873)) and not (layer0_outputs(5812));
    layer1_outputs(6631) <= '1';
    layer1_outputs(6632) <= not((layer0_outputs(6558)) and (layer0_outputs(1759)));
    layer1_outputs(6633) <= not(layer0_outputs(926)) or (layer0_outputs(1065));
    layer1_outputs(6634) <= not(layer0_outputs(8769));
    layer1_outputs(6635) <= layer0_outputs(667);
    layer1_outputs(6636) <= not(layer0_outputs(3847));
    layer1_outputs(6637) <= (layer0_outputs(2586)) and (layer0_outputs(6018));
    layer1_outputs(6638) <= not(layer0_outputs(4431));
    layer1_outputs(6639) <= not(layer0_outputs(7968)) or (layer0_outputs(7778));
    layer1_outputs(6640) <= layer0_outputs(383);
    layer1_outputs(6641) <= not((layer0_outputs(8749)) or (layer0_outputs(337)));
    layer1_outputs(6642) <= not((layer0_outputs(5601)) and (layer0_outputs(5003)));
    layer1_outputs(6643) <= layer0_outputs(6718);
    layer1_outputs(6644) <= (layer0_outputs(4994)) and not (layer0_outputs(5181));
    layer1_outputs(6645) <= (layer0_outputs(4572)) and not (layer0_outputs(5356));
    layer1_outputs(6646) <= (layer0_outputs(4173)) or (layer0_outputs(6389));
    layer1_outputs(6647) <= (layer0_outputs(8462)) and (layer0_outputs(5303));
    layer1_outputs(6648) <= layer0_outputs(7419);
    layer1_outputs(6649) <= (layer0_outputs(3961)) or (layer0_outputs(6400));
    layer1_outputs(6650) <= layer0_outputs(3418);
    layer1_outputs(6651) <= not(layer0_outputs(10122)) or (layer0_outputs(3589));
    layer1_outputs(6652) <= not((layer0_outputs(8066)) and (layer0_outputs(8053)));
    layer1_outputs(6653) <= not(layer0_outputs(9883));
    layer1_outputs(6654) <= not((layer0_outputs(6472)) and (layer0_outputs(590)));
    layer1_outputs(6655) <= (layer0_outputs(10082)) or (layer0_outputs(9053));
    layer1_outputs(6656) <= not(layer0_outputs(6337)) or (layer0_outputs(1323));
    layer1_outputs(6657) <= (layer0_outputs(6530)) and not (layer0_outputs(3830));
    layer1_outputs(6658) <= layer0_outputs(2326);
    layer1_outputs(6659) <= (layer0_outputs(6506)) or (layer0_outputs(4180));
    layer1_outputs(6660) <= (layer0_outputs(8183)) and not (layer0_outputs(4503));
    layer1_outputs(6661) <= (layer0_outputs(2915)) or (layer0_outputs(2723));
    layer1_outputs(6662) <= (layer0_outputs(7528)) and not (layer0_outputs(7530));
    layer1_outputs(6663) <= '0';
    layer1_outputs(6664) <= not(layer0_outputs(8698));
    layer1_outputs(6665) <= layer0_outputs(3745);
    layer1_outputs(6666) <= not((layer0_outputs(7480)) or (layer0_outputs(8233)));
    layer1_outputs(6667) <= (layer0_outputs(9587)) xor (layer0_outputs(734));
    layer1_outputs(6668) <= not((layer0_outputs(921)) and (layer0_outputs(5311)));
    layer1_outputs(6669) <= not(layer0_outputs(6458));
    layer1_outputs(6670) <= '0';
    layer1_outputs(6671) <= layer0_outputs(2335);
    layer1_outputs(6672) <= '0';
    layer1_outputs(6673) <= layer0_outputs(8861);
    layer1_outputs(6674) <= '0';
    layer1_outputs(6675) <= not(layer0_outputs(7201)) or (layer0_outputs(63));
    layer1_outputs(6676) <= layer0_outputs(2034);
    layer1_outputs(6677) <= layer0_outputs(1180);
    layer1_outputs(6678) <= (layer0_outputs(6981)) and not (layer0_outputs(655));
    layer1_outputs(6679) <= not(layer0_outputs(3219)) or (layer0_outputs(2551));
    layer1_outputs(6680) <= not(layer0_outputs(8549)) or (layer0_outputs(7065));
    layer1_outputs(6681) <= layer0_outputs(6241);
    layer1_outputs(6682) <= not(layer0_outputs(9407));
    layer1_outputs(6683) <= not(layer0_outputs(5197));
    layer1_outputs(6684) <= not(layer0_outputs(4590)) or (layer0_outputs(9073));
    layer1_outputs(6685) <= not(layer0_outputs(6787));
    layer1_outputs(6686) <= (layer0_outputs(7807)) or (layer0_outputs(1245));
    layer1_outputs(6687) <= layer0_outputs(2371);
    layer1_outputs(6688) <= not(layer0_outputs(8382)) or (layer0_outputs(3192));
    layer1_outputs(6689) <= not(layer0_outputs(3161)) or (layer0_outputs(3460));
    layer1_outputs(6690) <= layer0_outputs(3976);
    layer1_outputs(6691) <= not(layer0_outputs(4581));
    layer1_outputs(6692) <= '1';
    layer1_outputs(6693) <= not((layer0_outputs(1492)) and (layer0_outputs(2445)));
    layer1_outputs(6694) <= (layer0_outputs(4194)) and not (layer0_outputs(9741));
    layer1_outputs(6695) <= '0';
    layer1_outputs(6696) <= not(layer0_outputs(2433)) or (layer0_outputs(552));
    layer1_outputs(6697) <= '1';
    layer1_outputs(6698) <= not((layer0_outputs(5451)) xor (layer0_outputs(8275)));
    layer1_outputs(6699) <= (layer0_outputs(3324)) and not (layer0_outputs(3986));
    layer1_outputs(6700) <= layer0_outputs(3057);
    layer1_outputs(6701) <= not(layer0_outputs(2240));
    layer1_outputs(6702) <= layer0_outputs(710);
    layer1_outputs(6703) <= not((layer0_outputs(4000)) or (layer0_outputs(10121)));
    layer1_outputs(6704) <= (layer0_outputs(3035)) or (layer0_outputs(1375));
    layer1_outputs(6705) <= (layer0_outputs(3158)) and not (layer0_outputs(819));
    layer1_outputs(6706) <= (layer0_outputs(2692)) and (layer0_outputs(6459));
    layer1_outputs(6707) <= not(layer0_outputs(9916));
    layer1_outputs(6708) <= not((layer0_outputs(5275)) or (layer0_outputs(5634)));
    layer1_outputs(6709) <= (layer0_outputs(7559)) xor (layer0_outputs(4007));
    layer1_outputs(6710) <= (layer0_outputs(5208)) and not (layer0_outputs(1682));
    layer1_outputs(6711) <= (layer0_outputs(5099)) and (layer0_outputs(6801));
    layer1_outputs(6712) <= not(layer0_outputs(2813)) or (layer0_outputs(1758));
    layer1_outputs(6713) <= (layer0_outputs(4152)) or (layer0_outputs(9219));
    layer1_outputs(6714) <= not((layer0_outputs(10100)) and (layer0_outputs(5056)));
    layer1_outputs(6715) <= not(layer0_outputs(8806));
    layer1_outputs(6716) <= not(layer0_outputs(6879)) or (layer0_outputs(5865));
    layer1_outputs(6717) <= not(layer0_outputs(8208));
    layer1_outputs(6718) <= not(layer0_outputs(4891)) or (layer0_outputs(3366));
    layer1_outputs(6719) <= not((layer0_outputs(2292)) or (layer0_outputs(9131)));
    layer1_outputs(6720) <= layer0_outputs(8587);
    layer1_outputs(6721) <= not(layer0_outputs(6989));
    layer1_outputs(6722) <= not(layer0_outputs(753));
    layer1_outputs(6723) <= not((layer0_outputs(3049)) xor (layer0_outputs(347)));
    layer1_outputs(6724) <= not((layer0_outputs(1935)) and (layer0_outputs(1798)));
    layer1_outputs(6725) <= '0';
    layer1_outputs(6726) <= not(layer0_outputs(8253));
    layer1_outputs(6727) <= layer0_outputs(139);
    layer1_outputs(6728) <= not((layer0_outputs(8507)) or (layer0_outputs(3361)));
    layer1_outputs(6729) <= (layer0_outputs(6756)) and (layer0_outputs(162));
    layer1_outputs(6730) <= '0';
    layer1_outputs(6731) <= not((layer0_outputs(8424)) or (layer0_outputs(8246)));
    layer1_outputs(6732) <= (layer0_outputs(442)) and not (layer0_outputs(5823));
    layer1_outputs(6733) <= layer0_outputs(1168);
    layer1_outputs(6734) <= '0';
    layer1_outputs(6735) <= not(layer0_outputs(6946));
    layer1_outputs(6736) <= layer0_outputs(2073);
    layer1_outputs(6737) <= (layer0_outputs(4463)) xor (layer0_outputs(7894));
    layer1_outputs(6738) <= not((layer0_outputs(4765)) and (layer0_outputs(4682)));
    layer1_outputs(6739) <= not((layer0_outputs(9583)) or (layer0_outputs(4474)));
    layer1_outputs(6740) <= (layer0_outputs(4904)) xor (layer0_outputs(7792));
    layer1_outputs(6741) <= not(layer0_outputs(7842)) or (layer0_outputs(2147));
    layer1_outputs(6742) <= not((layer0_outputs(7685)) or (layer0_outputs(1930)));
    layer1_outputs(6743) <= (layer0_outputs(1470)) and (layer0_outputs(3822));
    layer1_outputs(6744) <= not(layer0_outputs(4501));
    layer1_outputs(6745) <= not(layer0_outputs(9182));
    layer1_outputs(6746) <= not(layer0_outputs(4039));
    layer1_outputs(6747) <= '1';
    layer1_outputs(6748) <= not(layer0_outputs(3088));
    layer1_outputs(6749) <= not(layer0_outputs(2375));
    layer1_outputs(6750) <= layer0_outputs(1119);
    layer1_outputs(6751) <= layer0_outputs(2710);
    layer1_outputs(6752) <= not(layer0_outputs(9486));
    layer1_outputs(6753) <= not((layer0_outputs(9538)) or (layer0_outputs(3886)));
    layer1_outputs(6754) <= not((layer0_outputs(3766)) or (layer0_outputs(9690)));
    layer1_outputs(6755) <= (layer0_outputs(813)) and (layer0_outputs(6641));
    layer1_outputs(6756) <= (layer0_outputs(7804)) and not (layer0_outputs(9077));
    layer1_outputs(6757) <= not((layer0_outputs(6127)) and (layer0_outputs(3467)));
    layer1_outputs(6758) <= not((layer0_outputs(3076)) and (layer0_outputs(3937)));
    layer1_outputs(6759) <= (layer0_outputs(7205)) or (layer0_outputs(8787));
    layer1_outputs(6760) <= (layer0_outputs(2542)) and (layer0_outputs(2461));
    layer1_outputs(6761) <= (layer0_outputs(2775)) and (layer0_outputs(4809));
    layer1_outputs(6762) <= (layer0_outputs(9855)) and (layer0_outputs(5406));
    layer1_outputs(6763) <= (layer0_outputs(3081)) and (layer0_outputs(10019));
    layer1_outputs(6764) <= not(layer0_outputs(4798)) or (layer0_outputs(2929));
    layer1_outputs(6765) <= not((layer0_outputs(3571)) xor (layer0_outputs(1593)));
    layer1_outputs(6766) <= not(layer0_outputs(3285));
    layer1_outputs(6767) <= (layer0_outputs(2980)) and (layer0_outputs(8507));
    layer1_outputs(6768) <= layer0_outputs(5032);
    layer1_outputs(6769) <= layer0_outputs(7163);
    layer1_outputs(6770) <= (layer0_outputs(7331)) and not (layer0_outputs(1579));
    layer1_outputs(6771) <= not(layer0_outputs(4486)) or (layer0_outputs(1652));
    layer1_outputs(6772) <= (layer0_outputs(4090)) or (layer0_outputs(2160));
    layer1_outputs(6773) <= not((layer0_outputs(8659)) and (layer0_outputs(6021)));
    layer1_outputs(6774) <= '0';
    layer1_outputs(6775) <= layer0_outputs(4101);
    layer1_outputs(6776) <= not((layer0_outputs(4748)) xor (layer0_outputs(4741)));
    layer1_outputs(6777) <= not(layer0_outputs(5833)) or (layer0_outputs(528));
    layer1_outputs(6778) <= not(layer0_outputs(3490));
    layer1_outputs(6779) <= (layer0_outputs(8639)) or (layer0_outputs(8347));
    layer1_outputs(6780) <= not((layer0_outputs(2479)) or (layer0_outputs(8394)));
    layer1_outputs(6781) <= not(layer0_outputs(3944)) or (layer0_outputs(4528));
    layer1_outputs(6782) <= not((layer0_outputs(8602)) and (layer0_outputs(2901)));
    layer1_outputs(6783) <= not((layer0_outputs(8100)) xor (layer0_outputs(8010)));
    layer1_outputs(6784) <= not(layer0_outputs(3345));
    layer1_outputs(6785) <= not((layer0_outputs(3532)) or (layer0_outputs(8413)));
    layer1_outputs(6786) <= layer0_outputs(438);
    layer1_outputs(6787) <= not((layer0_outputs(6481)) or (layer0_outputs(3085)));
    layer1_outputs(6788) <= not(layer0_outputs(6159));
    layer1_outputs(6789) <= (layer0_outputs(6877)) xor (layer0_outputs(5281));
    layer1_outputs(6790) <= (layer0_outputs(4385)) and (layer0_outputs(5574));
    layer1_outputs(6791) <= layer0_outputs(1292);
    layer1_outputs(6792) <= not((layer0_outputs(3066)) xor (layer0_outputs(10218)));
    layer1_outputs(6793) <= '1';
    layer1_outputs(6794) <= layer0_outputs(4461);
    layer1_outputs(6795) <= layer0_outputs(5054);
    layer1_outputs(6796) <= not(layer0_outputs(5310)) or (layer0_outputs(6033));
    layer1_outputs(6797) <= (layer0_outputs(7760)) or (layer0_outputs(729));
    layer1_outputs(6798) <= (layer0_outputs(306)) or (layer0_outputs(1064));
    layer1_outputs(6799) <= (layer0_outputs(10164)) and not (layer0_outputs(1169));
    layer1_outputs(6800) <= not((layer0_outputs(7712)) or (layer0_outputs(2098)));
    layer1_outputs(6801) <= not((layer0_outputs(308)) and (layer0_outputs(6030)));
    layer1_outputs(6802) <= layer0_outputs(494);
    layer1_outputs(6803) <= (layer0_outputs(5446)) and (layer0_outputs(4730));
    layer1_outputs(6804) <= not(layer0_outputs(8782));
    layer1_outputs(6805) <= (layer0_outputs(8580)) and not (layer0_outputs(6312));
    layer1_outputs(6806) <= not((layer0_outputs(2444)) or (layer0_outputs(1878)));
    layer1_outputs(6807) <= not(layer0_outputs(7469));
    layer1_outputs(6808) <= '0';
    layer1_outputs(6809) <= '0';
    layer1_outputs(6810) <= not(layer0_outputs(854)) or (layer0_outputs(6905));
    layer1_outputs(6811) <= '1';
    layer1_outputs(6812) <= not((layer0_outputs(4694)) xor (layer0_outputs(4844)));
    layer1_outputs(6813) <= (layer0_outputs(1512)) and (layer0_outputs(6538));
    layer1_outputs(6814) <= not((layer0_outputs(4178)) or (layer0_outputs(8434)));
    layer1_outputs(6815) <= not(layer0_outputs(2746));
    layer1_outputs(6816) <= not(layer0_outputs(10197)) or (layer0_outputs(326));
    layer1_outputs(6817) <= not(layer0_outputs(1366)) or (layer0_outputs(2398));
    layer1_outputs(6818) <= (layer0_outputs(6016)) and not (layer0_outputs(1415));
    layer1_outputs(6819) <= layer0_outputs(9921);
    layer1_outputs(6820) <= (layer0_outputs(4632)) or (layer0_outputs(7389));
    layer1_outputs(6821) <= (layer0_outputs(6691)) and not (layer0_outputs(5283));
    layer1_outputs(6822) <= layer0_outputs(893);
    layer1_outputs(6823) <= (layer0_outputs(2535)) and (layer0_outputs(3833));
    layer1_outputs(6824) <= '0';
    layer1_outputs(6825) <= not((layer0_outputs(7968)) or (layer0_outputs(4805)));
    layer1_outputs(6826) <= not(layer0_outputs(6137));
    layer1_outputs(6827) <= not((layer0_outputs(5957)) and (layer0_outputs(9)));
    layer1_outputs(6828) <= layer0_outputs(740);
    layer1_outputs(6829) <= layer0_outputs(1851);
    layer1_outputs(6830) <= layer0_outputs(2956);
    layer1_outputs(6831) <= not(layer0_outputs(2839)) or (layer0_outputs(3221));
    layer1_outputs(6832) <= (layer0_outputs(5862)) and not (layer0_outputs(8219));
    layer1_outputs(6833) <= not(layer0_outputs(7433)) or (layer0_outputs(4354));
    layer1_outputs(6834) <= not(layer0_outputs(9054));
    layer1_outputs(6835) <= not((layer0_outputs(9278)) or (layer0_outputs(10045)));
    layer1_outputs(6836) <= (layer0_outputs(8529)) and not (layer0_outputs(1143));
    layer1_outputs(6837) <= layer0_outputs(2343);
    layer1_outputs(6838) <= layer0_outputs(3735);
    layer1_outputs(6839) <= (layer0_outputs(9361)) and (layer0_outputs(1119));
    layer1_outputs(6840) <= not(layer0_outputs(8204)) or (layer0_outputs(7836));
    layer1_outputs(6841) <= (layer0_outputs(4136)) and not (layer0_outputs(9675));
    layer1_outputs(6842) <= (layer0_outputs(1786)) xor (layer0_outputs(7834));
    layer1_outputs(6843) <= not(layer0_outputs(3273));
    layer1_outputs(6844) <= (layer0_outputs(117)) and (layer0_outputs(3041));
    layer1_outputs(6845) <= layer0_outputs(7603);
    layer1_outputs(6846) <= (layer0_outputs(724)) xor (layer0_outputs(7037));
    layer1_outputs(6847) <= not(layer0_outputs(5356));
    layer1_outputs(6848) <= not(layer0_outputs(9135));
    layer1_outputs(6849) <= (layer0_outputs(9742)) and (layer0_outputs(7431));
    layer1_outputs(6850) <= (layer0_outputs(6544)) or (layer0_outputs(7254));
    layer1_outputs(6851) <= not(layer0_outputs(7051));
    layer1_outputs(6852) <= (layer0_outputs(3029)) or (layer0_outputs(4803));
    layer1_outputs(6853) <= (layer0_outputs(2393)) and (layer0_outputs(1599));
    layer1_outputs(6854) <= layer0_outputs(4770);
    layer1_outputs(6855) <= (layer0_outputs(8455)) and not (layer0_outputs(638));
    layer1_outputs(6856) <= not(layer0_outputs(3692));
    layer1_outputs(6857) <= (layer0_outputs(2675)) and (layer0_outputs(1740));
    layer1_outputs(6858) <= not(layer0_outputs(6)) or (layer0_outputs(7035));
    layer1_outputs(6859) <= not(layer0_outputs(3711)) or (layer0_outputs(9765));
    layer1_outputs(6860) <= (layer0_outputs(3737)) and not (layer0_outputs(2007));
    layer1_outputs(6861) <= not((layer0_outputs(9236)) or (layer0_outputs(8021)));
    layer1_outputs(6862) <= (layer0_outputs(8102)) and not (layer0_outputs(29));
    layer1_outputs(6863) <= not(layer0_outputs(5588)) or (layer0_outputs(8893));
    layer1_outputs(6864) <= not(layer0_outputs(1367)) or (layer0_outputs(8440));
    layer1_outputs(6865) <= (layer0_outputs(9198)) and not (layer0_outputs(4426));
    layer1_outputs(6866) <= (layer0_outputs(44)) and not (layer0_outputs(7860));
    layer1_outputs(6867) <= not(layer0_outputs(8874)) or (layer0_outputs(2648));
    layer1_outputs(6868) <= (layer0_outputs(1214)) xor (layer0_outputs(2595));
    layer1_outputs(6869) <= not(layer0_outputs(390));
    layer1_outputs(6870) <= '1';
    layer1_outputs(6871) <= layer0_outputs(7714);
    layer1_outputs(6872) <= '1';
    layer1_outputs(6873) <= layer0_outputs(8594);
    layer1_outputs(6874) <= (layer0_outputs(1715)) and (layer0_outputs(8216));
    layer1_outputs(6875) <= (layer0_outputs(4698)) and (layer0_outputs(8834));
    layer1_outputs(6876) <= not((layer0_outputs(7611)) xor (layer0_outputs(2213)));
    layer1_outputs(6877) <= not(layer0_outputs(6934));
    layer1_outputs(6878) <= (layer0_outputs(1301)) and not (layer0_outputs(6467));
    layer1_outputs(6879) <= (layer0_outputs(6822)) and (layer0_outputs(1830));
    layer1_outputs(6880) <= layer0_outputs(5946);
    layer1_outputs(6881) <= layer0_outputs(8880);
    layer1_outputs(6882) <= not(layer0_outputs(4949));
    layer1_outputs(6883) <= '1';
    layer1_outputs(6884) <= (layer0_outputs(2023)) and not (layer0_outputs(9070));
    layer1_outputs(6885) <= (layer0_outputs(9960)) and (layer0_outputs(4175));
    layer1_outputs(6886) <= not(layer0_outputs(6488));
    layer1_outputs(6887) <= (layer0_outputs(3199)) xor (layer0_outputs(8299));
    layer1_outputs(6888) <= layer0_outputs(7121);
    layer1_outputs(6889) <= not((layer0_outputs(4906)) and (layer0_outputs(243)));
    layer1_outputs(6890) <= not(layer0_outputs(8347));
    layer1_outputs(6891) <= (layer0_outputs(2436)) and not (layer0_outputs(2157));
    layer1_outputs(6892) <= layer0_outputs(230);
    layer1_outputs(6893) <= not((layer0_outputs(4965)) or (layer0_outputs(7054)));
    layer1_outputs(6894) <= '0';
    layer1_outputs(6895) <= (layer0_outputs(3965)) and not (layer0_outputs(8831));
    layer1_outputs(6896) <= (layer0_outputs(4943)) or (layer0_outputs(8085));
    layer1_outputs(6897) <= (layer0_outputs(636)) and (layer0_outputs(6861));
    layer1_outputs(6898) <= not(layer0_outputs(8314));
    layer1_outputs(6899) <= not((layer0_outputs(1096)) or (layer0_outputs(9129)));
    layer1_outputs(6900) <= not((layer0_outputs(1653)) xor (layer0_outputs(5098)));
    layer1_outputs(6901) <= layer0_outputs(10049);
    layer1_outputs(6902) <= not(layer0_outputs(3933)) or (layer0_outputs(6037));
    layer1_outputs(6903) <= layer0_outputs(9057);
    layer1_outputs(6904) <= layer0_outputs(9174);
    layer1_outputs(6905) <= (layer0_outputs(2009)) xor (layer0_outputs(1181));
    layer1_outputs(6906) <= (layer0_outputs(655)) xor (layer0_outputs(3195));
    layer1_outputs(6907) <= (layer0_outputs(5863)) and (layer0_outputs(4779));
    layer1_outputs(6908) <= '1';
    layer1_outputs(6909) <= (layer0_outputs(10198)) and not (layer0_outputs(8794));
    layer1_outputs(6910) <= (layer0_outputs(6674)) xor (layer0_outputs(3644));
    layer1_outputs(6911) <= layer0_outputs(8371);
    layer1_outputs(6912) <= '1';
    layer1_outputs(6913) <= not(layer0_outputs(2081));
    layer1_outputs(6914) <= '0';
    layer1_outputs(6915) <= not(layer0_outputs(9899));
    layer1_outputs(6916) <= (layer0_outputs(8530)) and not (layer0_outputs(570));
    layer1_outputs(6917) <= not(layer0_outputs(2662));
    layer1_outputs(6918) <= not(layer0_outputs(6794));
    layer1_outputs(6919) <= not((layer0_outputs(1879)) or (layer0_outputs(732)));
    layer1_outputs(6920) <= (layer0_outputs(7605)) and not (layer0_outputs(574));
    layer1_outputs(6921) <= (layer0_outputs(7292)) and not (layer0_outputs(8221));
    layer1_outputs(6922) <= (layer0_outputs(8014)) and not (layer0_outputs(6641));
    layer1_outputs(6923) <= (layer0_outputs(8962)) or (layer0_outputs(4903));
    layer1_outputs(6924) <= not(layer0_outputs(7537)) or (layer0_outputs(8296));
    layer1_outputs(6925) <= not(layer0_outputs(9259)) or (layer0_outputs(9783));
    layer1_outputs(6926) <= (layer0_outputs(5354)) xor (layer0_outputs(3631));
    layer1_outputs(6927) <= layer0_outputs(8214);
    layer1_outputs(6928) <= '0';
    layer1_outputs(6929) <= not((layer0_outputs(3179)) or (layer0_outputs(7229)));
    layer1_outputs(6930) <= not(layer0_outputs(301)) or (layer0_outputs(7622));
    layer1_outputs(6931) <= layer0_outputs(3452);
    layer1_outputs(6932) <= not(layer0_outputs(4266)) or (layer0_outputs(1328));
    layer1_outputs(6933) <= '0';
    layer1_outputs(6934) <= not((layer0_outputs(3432)) xor (layer0_outputs(7112)));
    layer1_outputs(6935) <= not(layer0_outputs(8661)) or (layer0_outputs(1971));
    layer1_outputs(6936) <= not(layer0_outputs(8586));
    layer1_outputs(6937) <= (layer0_outputs(9824)) and not (layer0_outputs(698));
    layer1_outputs(6938) <= layer0_outputs(8875);
    layer1_outputs(6939) <= not(layer0_outputs(9343)) or (layer0_outputs(5749));
    layer1_outputs(6940) <= (layer0_outputs(3958)) and not (layer0_outputs(5498));
    layer1_outputs(6941) <= not(layer0_outputs(9411));
    layer1_outputs(6942) <= layer0_outputs(9047);
    layer1_outputs(6943) <= (layer0_outputs(1922)) or (layer0_outputs(9024));
    layer1_outputs(6944) <= not(layer0_outputs(5206)) or (layer0_outputs(7615));
    layer1_outputs(6945) <= not(layer0_outputs(8541));
    layer1_outputs(6946) <= layer0_outputs(876);
    layer1_outputs(6947) <= not(layer0_outputs(3284)) or (layer0_outputs(2218));
    layer1_outputs(6948) <= (layer0_outputs(9162)) and (layer0_outputs(2372));
    layer1_outputs(6949) <= layer0_outputs(1952);
    layer1_outputs(6950) <= not((layer0_outputs(6563)) or (layer0_outputs(5626)));
    layer1_outputs(6951) <= '0';
    layer1_outputs(6952) <= (layer0_outputs(5614)) and not (layer0_outputs(5058));
    layer1_outputs(6953) <= layer0_outputs(9944);
    layer1_outputs(6954) <= layer0_outputs(985);
    layer1_outputs(6955) <= (layer0_outputs(5916)) xor (layer0_outputs(5174));
    layer1_outputs(6956) <= layer0_outputs(5610);
    layer1_outputs(6957) <= (layer0_outputs(884)) and not (layer0_outputs(6133));
    layer1_outputs(6958) <= (layer0_outputs(2999)) or (layer0_outputs(399));
    layer1_outputs(6959) <= not(layer0_outputs(4968)) or (layer0_outputs(9052));
    layer1_outputs(6960) <= '1';
    layer1_outputs(6961) <= not((layer0_outputs(9831)) and (layer0_outputs(8697)));
    layer1_outputs(6962) <= (layer0_outputs(1462)) xor (layer0_outputs(9822));
    layer1_outputs(6963) <= (layer0_outputs(1996)) and (layer0_outputs(5493));
    layer1_outputs(6964) <= not((layer0_outputs(4587)) or (layer0_outputs(2677)));
    layer1_outputs(6965) <= (layer0_outputs(7582)) and not (layer0_outputs(5397));
    layer1_outputs(6966) <= layer0_outputs(299);
    layer1_outputs(6967) <= layer0_outputs(3015);
    layer1_outputs(6968) <= not(layer0_outputs(5026)) or (layer0_outputs(1721));
    layer1_outputs(6969) <= '0';
    layer1_outputs(6970) <= layer0_outputs(7167);
    layer1_outputs(6971) <= not(layer0_outputs(3684)) or (layer0_outputs(8405));
    layer1_outputs(6972) <= (layer0_outputs(1598)) or (layer0_outputs(1806));
    layer1_outputs(6973) <= not(layer0_outputs(3203));
    layer1_outputs(6974) <= '1';
    layer1_outputs(6975) <= layer0_outputs(3254);
    layer1_outputs(6976) <= (layer0_outputs(2763)) xor (layer0_outputs(815));
    layer1_outputs(6977) <= (layer0_outputs(2520)) and not (layer0_outputs(47));
    layer1_outputs(6978) <= layer0_outputs(9265);
    layer1_outputs(6979) <= layer0_outputs(8647);
    layer1_outputs(6980) <= not(layer0_outputs(4490));
    layer1_outputs(6981) <= layer0_outputs(2892);
    layer1_outputs(6982) <= not(layer0_outputs(7534));
    layer1_outputs(6983) <= layer0_outputs(8700);
    layer1_outputs(6984) <= (layer0_outputs(8727)) and not (layer0_outputs(1647));
    layer1_outputs(6985) <= (layer0_outputs(8519)) and (layer0_outputs(3639));
    layer1_outputs(6986) <= not(layer0_outputs(7370));
    layer1_outputs(6987) <= not(layer0_outputs(8011)) or (layer0_outputs(8568));
    layer1_outputs(6988) <= (layer0_outputs(3317)) and not (layer0_outputs(1726));
    layer1_outputs(6989) <= not((layer0_outputs(5604)) xor (layer0_outputs(5641)));
    layer1_outputs(6990) <= not(layer0_outputs(7966)) or (layer0_outputs(8133));
    layer1_outputs(6991) <= layer0_outputs(2560);
    layer1_outputs(6992) <= (layer0_outputs(1886)) and not (layer0_outputs(9561));
    layer1_outputs(6993) <= (layer0_outputs(5339)) xor (layer0_outputs(9213));
    layer1_outputs(6994) <= (layer0_outputs(2800)) and not (layer0_outputs(9913));
    layer1_outputs(6995) <= not(layer0_outputs(2885)) or (layer0_outputs(5585));
    layer1_outputs(6996) <= not(layer0_outputs(5184)) or (layer0_outputs(1281));
    layer1_outputs(6997) <= layer0_outputs(8401);
    layer1_outputs(6998) <= not(layer0_outputs(8984));
    layer1_outputs(6999) <= not((layer0_outputs(5384)) or (layer0_outputs(8333)));
    layer1_outputs(7000) <= (layer0_outputs(22)) and not (layer0_outputs(8914));
    layer1_outputs(7001) <= not((layer0_outputs(8631)) or (layer0_outputs(6206)));
    layer1_outputs(7002) <= layer0_outputs(9645);
    layer1_outputs(7003) <= layer0_outputs(6896);
    layer1_outputs(7004) <= layer0_outputs(5425);
    layer1_outputs(7005) <= not(layer0_outputs(2446));
    layer1_outputs(7006) <= layer0_outputs(5676);
    layer1_outputs(7007) <= not((layer0_outputs(3325)) and (layer0_outputs(6445)));
    layer1_outputs(7008) <= (layer0_outputs(6959)) and (layer0_outputs(2782));
    layer1_outputs(7009) <= not(layer0_outputs(6247)) or (layer0_outputs(4327));
    layer1_outputs(7010) <= not(layer0_outputs(478)) or (layer0_outputs(1769));
    layer1_outputs(7011) <= not((layer0_outputs(2987)) or (layer0_outputs(8040)));
    layer1_outputs(7012) <= (layer0_outputs(10139)) and not (layer0_outputs(562));
    layer1_outputs(7013) <= (layer0_outputs(9516)) and (layer0_outputs(4177));
    layer1_outputs(7014) <= not(layer0_outputs(6057));
    layer1_outputs(7015) <= layer0_outputs(7687);
    layer1_outputs(7016) <= (layer0_outputs(10143)) or (layer0_outputs(5525));
    layer1_outputs(7017) <= layer0_outputs(8251);
    layer1_outputs(7018) <= (layer0_outputs(10082)) and not (layer0_outputs(676));
    layer1_outputs(7019) <= (layer0_outputs(4686)) and not (layer0_outputs(4437));
    layer1_outputs(7020) <= '0';
    layer1_outputs(7021) <= layer0_outputs(7620);
    layer1_outputs(7022) <= not(layer0_outputs(8238));
    layer1_outputs(7023) <= '0';
    layer1_outputs(7024) <= not((layer0_outputs(6272)) and (layer0_outputs(7355)));
    layer1_outputs(7025) <= not((layer0_outputs(8729)) xor (layer0_outputs(6849)));
    layer1_outputs(7026) <= (layer0_outputs(4974)) and not (layer0_outputs(8175));
    layer1_outputs(7027) <= (layer0_outputs(5041)) and not (layer0_outputs(486));
    layer1_outputs(7028) <= '0';
    layer1_outputs(7029) <= (layer0_outputs(5201)) and not (layer0_outputs(7151));
    layer1_outputs(7030) <= not(layer0_outputs(384));
    layer1_outputs(7031) <= layer0_outputs(5655);
    layer1_outputs(7032) <= not((layer0_outputs(6056)) or (layer0_outputs(2415)));
    layer1_outputs(7033) <= not(layer0_outputs(6303)) or (layer0_outputs(6100));
    layer1_outputs(7034) <= not(layer0_outputs(8979));
    layer1_outputs(7035) <= '0';
    layer1_outputs(7036) <= layer0_outputs(2869);
    layer1_outputs(7037) <= (layer0_outputs(3605)) and (layer0_outputs(4167));
    layer1_outputs(7038) <= not(layer0_outputs(7055)) or (layer0_outputs(2265));
    layer1_outputs(7039) <= (layer0_outputs(4236)) and (layer0_outputs(29));
    layer1_outputs(7040) <= (layer0_outputs(5994)) and (layer0_outputs(584));
    layer1_outputs(7041) <= not(layer0_outputs(1240));
    layer1_outputs(7042) <= (layer0_outputs(4514)) and not (layer0_outputs(8617));
    layer1_outputs(7043) <= not((layer0_outputs(3434)) xor (layer0_outputs(9532)));
    layer1_outputs(7044) <= not((layer0_outputs(2014)) or (layer0_outputs(2019)));
    layer1_outputs(7045) <= not((layer0_outputs(4271)) xor (layer0_outputs(1919)));
    layer1_outputs(7046) <= layer0_outputs(404);
    layer1_outputs(7047) <= not((layer0_outputs(5315)) and (layer0_outputs(4893)));
    layer1_outputs(7048) <= not(layer0_outputs(1996)) or (layer0_outputs(1788));
    layer1_outputs(7049) <= layer0_outputs(5653);
    layer1_outputs(7050) <= layer0_outputs(1258);
    layer1_outputs(7051) <= not(layer0_outputs(2592));
    layer1_outputs(7052) <= not(layer0_outputs(2003));
    layer1_outputs(7053) <= not((layer0_outputs(7536)) xor (layer0_outputs(4945)));
    layer1_outputs(7054) <= (layer0_outputs(430)) and not (layer0_outputs(3940));
    layer1_outputs(7055) <= (layer0_outputs(5069)) or (layer0_outputs(4392));
    layer1_outputs(7056) <= not(layer0_outputs(10077)) or (layer0_outputs(793));
    layer1_outputs(7057) <= not(layer0_outputs(2750)) or (layer0_outputs(6142));
    layer1_outputs(7058) <= '0';
    layer1_outputs(7059) <= (layer0_outputs(9176)) and not (layer0_outputs(404));
    layer1_outputs(7060) <= not((layer0_outputs(8286)) or (layer0_outputs(6)));
    layer1_outputs(7061) <= (layer0_outputs(3601)) and not (layer0_outputs(7446));
    layer1_outputs(7062) <= '1';
    layer1_outputs(7063) <= layer0_outputs(3495);
    layer1_outputs(7064) <= not(layer0_outputs(5301)) or (layer0_outputs(2603));
    layer1_outputs(7065) <= not(layer0_outputs(5858)) or (layer0_outputs(471));
    layer1_outputs(7066) <= not(layer0_outputs(5278));
    layer1_outputs(7067) <= (layer0_outputs(6714)) xor (layer0_outputs(4022));
    layer1_outputs(7068) <= not(layer0_outputs(3492));
    layer1_outputs(7069) <= '0';
    layer1_outputs(7070) <= layer0_outputs(7478);
    layer1_outputs(7071) <= not(layer0_outputs(3084));
    layer1_outputs(7072) <= not(layer0_outputs(7285));
    layer1_outputs(7073) <= (layer0_outputs(4429)) xor (layer0_outputs(2152));
    layer1_outputs(7074) <= not(layer0_outputs(5442)) or (layer0_outputs(3084));
    layer1_outputs(7075) <= (layer0_outputs(3481)) or (layer0_outputs(9456));
    layer1_outputs(7076) <= layer0_outputs(6240);
    layer1_outputs(7077) <= not(layer0_outputs(2613)) or (layer0_outputs(6156));
    layer1_outputs(7078) <= '1';
    layer1_outputs(7079) <= '0';
    layer1_outputs(7080) <= layer0_outputs(3452);
    layer1_outputs(7081) <= not((layer0_outputs(7862)) xor (layer0_outputs(9909)));
    layer1_outputs(7082) <= not((layer0_outputs(175)) or (layer0_outputs(2481)));
    layer1_outputs(7083) <= not((layer0_outputs(7361)) or (layer0_outputs(1827)));
    layer1_outputs(7084) <= not(layer0_outputs(6037));
    layer1_outputs(7085) <= not((layer0_outputs(826)) xor (layer0_outputs(1072)));
    layer1_outputs(7086) <= not((layer0_outputs(9549)) or (layer0_outputs(8575)));
    layer1_outputs(7087) <= not((layer0_outputs(1809)) xor (layer0_outputs(5774)));
    layer1_outputs(7088) <= not((layer0_outputs(3840)) xor (layer0_outputs(2177)));
    layer1_outputs(7089) <= not((layer0_outputs(5381)) and (layer0_outputs(2135)));
    layer1_outputs(7090) <= '0';
    layer1_outputs(7091) <= '1';
    layer1_outputs(7092) <= not((layer0_outputs(1958)) or (layer0_outputs(9625)));
    layer1_outputs(7093) <= not(layer0_outputs(8658)) or (layer0_outputs(1026));
    layer1_outputs(7094) <= (layer0_outputs(5235)) and (layer0_outputs(8343));
    layer1_outputs(7095) <= '0';
    layer1_outputs(7096) <= not((layer0_outputs(9132)) and (layer0_outputs(9553)));
    layer1_outputs(7097) <= (layer0_outputs(152)) and not (layer0_outputs(4849));
    layer1_outputs(7098) <= not(layer0_outputs(8265)) or (layer0_outputs(2496));
    layer1_outputs(7099) <= not(layer0_outputs(2129)) or (layer0_outputs(5609));
    layer1_outputs(7100) <= not(layer0_outputs(7169)) or (layer0_outputs(8941));
    layer1_outputs(7101) <= '0';
    layer1_outputs(7102) <= not(layer0_outputs(6154));
    layer1_outputs(7103) <= not(layer0_outputs(7280)) or (layer0_outputs(3206));
    layer1_outputs(7104) <= not(layer0_outputs(4573));
    layer1_outputs(7105) <= not(layer0_outputs(5217));
    layer1_outputs(7106) <= not(layer0_outputs(9755));
    layer1_outputs(7107) <= layer0_outputs(2989);
    layer1_outputs(7108) <= (layer0_outputs(8051)) or (layer0_outputs(3374));
    layer1_outputs(7109) <= not(layer0_outputs(1360)) or (layer0_outputs(3739));
    layer1_outputs(7110) <= (layer0_outputs(9896)) xor (layer0_outputs(9844));
    layer1_outputs(7111) <= (layer0_outputs(2387)) xor (layer0_outputs(746));
    layer1_outputs(7112) <= not(layer0_outputs(6751));
    layer1_outputs(7113) <= '1';
    layer1_outputs(7114) <= not(layer0_outputs(8631)) or (layer0_outputs(3110));
    layer1_outputs(7115) <= layer0_outputs(2119);
    layer1_outputs(7116) <= layer0_outputs(1516);
    layer1_outputs(7117) <= not((layer0_outputs(2686)) and (layer0_outputs(9498)));
    layer1_outputs(7118) <= '1';
    layer1_outputs(7119) <= (layer0_outputs(2701)) and not (layer0_outputs(7707));
    layer1_outputs(7120) <= not((layer0_outputs(7451)) or (layer0_outputs(7800)));
    layer1_outputs(7121) <= '1';
    layer1_outputs(7122) <= layer0_outputs(5146);
    layer1_outputs(7123) <= layer0_outputs(9112);
    layer1_outputs(7124) <= not(layer0_outputs(1031));
    layer1_outputs(7125) <= layer0_outputs(9853);
    layer1_outputs(7126) <= not((layer0_outputs(8364)) xor (layer0_outputs(9860)));
    layer1_outputs(7127) <= not(layer0_outputs(10191));
    layer1_outputs(7128) <= (layer0_outputs(7375)) and not (layer0_outputs(1029));
    layer1_outputs(7129) <= not(layer0_outputs(4695)) or (layer0_outputs(4429));
    layer1_outputs(7130) <= not(layer0_outputs(9852));
    layer1_outputs(7131) <= layer0_outputs(775);
    layer1_outputs(7132) <= not(layer0_outputs(5002));
    layer1_outputs(7133) <= not(layer0_outputs(8524));
    layer1_outputs(7134) <= layer0_outputs(9241);
    layer1_outputs(7135) <= (layer0_outputs(10223)) and (layer0_outputs(3000));
    layer1_outputs(7136) <= not(layer0_outputs(3011)) or (layer0_outputs(493));
    layer1_outputs(7137) <= layer0_outputs(8032);
    layer1_outputs(7138) <= (layer0_outputs(5210)) and not (layer0_outputs(131));
    layer1_outputs(7139) <= layer0_outputs(888);
    layer1_outputs(7140) <= (layer0_outputs(7987)) or (layer0_outputs(738));
    layer1_outputs(7141) <= not((layer0_outputs(6936)) or (layer0_outputs(3526)));
    layer1_outputs(7142) <= not((layer0_outputs(7258)) or (layer0_outputs(2282)));
    layer1_outputs(7143) <= (layer0_outputs(1217)) xor (layer0_outputs(1582));
    layer1_outputs(7144) <= (layer0_outputs(5544)) xor (layer0_outputs(2148));
    layer1_outputs(7145) <= not(layer0_outputs(3890));
    layer1_outputs(7146) <= not((layer0_outputs(1369)) and (layer0_outputs(8084)));
    layer1_outputs(7147) <= not((layer0_outputs(3261)) or (layer0_outputs(1589)));
    layer1_outputs(7148) <= not(layer0_outputs(5783)) or (layer0_outputs(7102));
    layer1_outputs(7149) <= layer0_outputs(6934);
    layer1_outputs(7150) <= (layer0_outputs(9956)) and (layer0_outputs(8049));
    layer1_outputs(7151) <= not(layer0_outputs(2971)) or (layer0_outputs(4901));
    layer1_outputs(7152) <= not(layer0_outputs(1320)) or (layer0_outputs(1584));
    layer1_outputs(7153) <= '0';
    layer1_outputs(7154) <= (layer0_outputs(480)) xor (layer0_outputs(5169));
    layer1_outputs(7155) <= '1';
    layer1_outputs(7156) <= not((layer0_outputs(5)) or (layer0_outputs(5151)));
    layer1_outputs(7157) <= layer0_outputs(5459);
    layer1_outputs(7158) <= not(layer0_outputs(1686)) or (layer0_outputs(2347));
    layer1_outputs(7159) <= (layer0_outputs(1766)) or (layer0_outputs(2091));
    layer1_outputs(7160) <= layer0_outputs(1480);
    layer1_outputs(7161) <= '0';
    layer1_outputs(7162) <= not(layer0_outputs(3610));
    layer1_outputs(7163) <= (layer0_outputs(3850)) xor (layer0_outputs(7454));
    layer1_outputs(7164) <= not(layer0_outputs(6057));
    layer1_outputs(7165) <= not(layer0_outputs(6359)) or (layer0_outputs(380));
    layer1_outputs(7166) <= not((layer0_outputs(3581)) or (layer0_outputs(9144)));
    layer1_outputs(7167) <= layer0_outputs(5117);
    layer1_outputs(7168) <= not(layer0_outputs(1486));
    layer1_outputs(7169) <= not(layer0_outputs(5280)) or (layer0_outputs(9906));
    layer1_outputs(7170) <= (layer0_outputs(586)) and not (layer0_outputs(8501));
    layer1_outputs(7171) <= '1';
    layer1_outputs(7172) <= (layer0_outputs(4780)) and not (layer0_outputs(1523));
    layer1_outputs(7173) <= not(layer0_outputs(6376));
    layer1_outputs(7174) <= not(layer0_outputs(7385)) or (layer0_outputs(2731));
    layer1_outputs(7175) <= not(layer0_outputs(3419)) or (layer0_outputs(4299));
    layer1_outputs(7176) <= '1';
    layer1_outputs(7177) <= layer0_outputs(8123);
    layer1_outputs(7178) <= not(layer0_outputs(3397));
    layer1_outputs(7179) <= not((layer0_outputs(1226)) or (layer0_outputs(8648)));
    layer1_outputs(7180) <= not(layer0_outputs(2065));
    layer1_outputs(7181) <= (layer0_outputs(1995)) and not (layer0_outputs(7900));
    layer1_outputs(7182) <= (layer0_outputs(7940)) or (layer0_outputs(4613));
    layer1_outputs(7183) <= (layer0_outputs(3193)) or (layer0_outputs(5005));
    layer1_outputs(7184) <= not(layer0_outputs(9794));
    layer1_outputs(7185) <= (layer0_outputs(8215)) xor (layer0_outputs(7646));
    layer1_outputs(7186) <= layer0_outputs(6954);
    layer1_outputs(7187) <= (layer0_outputs(8969)) or (layer0_outputs(6809));
    layer1_outputs(7188) <= not((layer0_outputs(3642)) xor (layer0_outputs(3004)));
    layer1_outputs(7189) <= not(layer0_outputs(7943));
    layer1_outputs(7190) <= not(layer0_outputs(2772)) or (layer0_outputs(1292));
    layer1_outputs(7191) <= '1';
    layer1_outputs(7192) <= not(layer0_outputs(8674)) or (layer0_outputs(1585));
    layer1_outputs(7193) <= not(layer0_outputs(2284));
    layer1_outputs(7194) <= layer0_outputs(5314);
    layer1_outputs(7195) <= layer0_outputs(2864);
    layer1_outputs(7196) <= not(layer0_outputs(6834));
    layer1_outputs(7197) <= layer0_outputs(2621);
    layer1_outputs(7198) <= (layer0_outputs(9552)) and (layer0_outputs(7487));
    layer1_outputs(7199) <= '0';
    layer1_outputs(7200) <= not(layer0_outputs(9083)) or (layer0_outputs(870));
    layer1_outputs(7201) <= layer0_outputs(265);
    layer1_outputs(7202) <= not((layer0_outputs(8931)) and (layer0_outputs(9268)));
    layer1_outputs(7203) <= (layer0_outputs(6390)) and not (layer0_outputs(10132));
    layer1_outputs(7204) <= (layer0_outputs(4435)) or (layer0_outputs(3292));
    layer1_outputs(7205) <= layer0_outputs(3687);
    layer1_outputs(7206) <= not(layer0_outputs(606));
    layer1_outputs(7207) <= not((layer0_outputs(8858)) xor (layer0_outputs(1202)));
    layer1_outputs(7208) <= not((layer0_outputs(5112)) xor (layer0_outputs(3628)));
    layer1_outputs(7209) <= not(layer0_outputs(4138));
    layer1_outputs(7210) <= layer0_outputs(5427);
    layer1_outputs(7211) <= not((layer0_outputs(5791)) and (layer0_outputs(9016)));
    layer1_outputs(7212) <= (layer0_outputs(4972)) and not (layer0_outputs(5938));
    layer1_outputs(7213) <= not(layer0_outputs(8800));
    layer1_outputs(7214) <= (layer0_outputs(8451)) and (layer0_outputs(9561));
    layer1_outputs(7215) <= (layer0_outputs(7256)) and (layer0_outputs(7524));
    layer1_outputs(7216) <= layer0_outputs(7497);
    layer1_outputs(7217) <= (layer0_outputs(843)) and (layer0_outputs(7918));
    layer1_outputs(7218) <= not(layer0_outputs(323));
    layer1_outputs(7219) <= (layer0_outputs(7752)) and not (layer0_outputs(3490));
    layer1_outputs(7220) <= not(layer0_outputs(7872)) or (layer0_outputs(7835));
    layer1_outputs(7221) <= not(layer0_outputs(8800));
    layer1_outputs(7222) <= not(layer0_outputs(7721));
    layer1_outputs(7223) <= (layer0_outputs(7715)) and (layer0_outputs(8555));
    layer1_outputs(7224) <= (layer0_outputs(2050)) xor (layer0_outputs(3748));
    layer1_outputs(7225) <= layer0_outputs(4965);
    layer1_outputs(7226) <= '1';
    layer1_outputs(7227) <= not((layer0_outputs(4884)) or (layer0_outputs(5744)));
    layer1_outputs(7228) <= not(layer0_outputs(9444));
    layer1_outputs(7229) <= not((layer0_outputs(3653)) or (layer0_outputs(3999)));
    layer1_outputs(7230) <= not(layer0_outputs(5003));
    layer1_outputs(7231) <= not((layer0_outputs(4942)) xor (layer0_outputs(9917)));
    layer1_outputs(7232) <= layer0_outputs(7574);
    layer1_outputs(7233) <= not((layer0_outputs(9169)) and (layer0_outputs(5497)));
    layer1_outputs(7234) <= not((layer0_outputs(6472)) xor (layer0_outputs(8024)));
    layer1_outputs(7235) <= (layer0_outputs(4975)) and not (layer0_outputs(8310));
    layer1_outputs(7236) <= (layer0_outputs(6850)) or (layer0_outputs(8980));
    layer1_outputs(7237) <= not(layer0_outputs(2112)) or (layer0_outputs(6682));
    layer1_outputs(7238) <= '1';
    layer1_outputs(7239) <= not(layer0_outputs(8269));
    layer1_outputs(7240) <= not(layer0_outputs(38)) or (layer0_outputs(3632));
    layer1_outputs(7241) <= '0';
    layer1_outputs(7242) <= not(layer0_outputs(5926));
    layer1_outputs(7243) <= layer0_outputs(5268);
    layer1_outputs(7244) <= layer0_outputs(7270);
    layer1_outputs(7245) <= (layer0_outputs(10006)) and not (layer0_outputs(9820));
    layer1_outputs(7246) <= not(layer0_outputs(6451));
    layer1_outputs(7247) <= not(layer0_outputs(5996));
    layer1_outputs(7248) <= not(layer0_outputs(5785));
    layer1_outputs(7249) <= not(layer0_outputs(4937));
    layer1_outputs(7250) <= (layer0_outputs(9414)) and not (layer0_outputs(9268));
    layer1_outputs(7251) <= (layer0_outputs(2471)) or (layer0_outputs(8357));
    layer1_outputs(7252) <= (layer0_outputs(8307)) and not (layer0_outputs(10236));
    layer1_outputs(7253) <= '0';
    layer1_outputs(7254) <= layer0_outputs(1928);
    layer1_outputs(7255) <= not(layer0_outputs(1298)) or (layer0_outputs(1759));
    layer1_outputs(7256) <= '0';
    layer1_outputs(7257) <= layer0_outputs(6514);
    layer1_outputs(7258) <= layer0_outputs(6727);
    layer1_outputs(7259) <= not((layer0_outputs(288)) or (layer0_outputs(4610)));
    layer1_outputs(7260) <= layer0_outputs(10209);
    layer1_outputs(7261) <= (layer0_outputs(7576)) and not (layer0_outputs(5180));
    layer1_outputs(7262) <= (layer0_outputs(4599)) or (layer0_outputs(7865));
    layer1_outputs(7263) <= (layer0_outputs(10125)) or (layer0_outputs(7912));
    layer1_outputs(7264) <= (layer0_outputs(5007)) or (layer0_outputs(7391));
    layer1_outputs(7265) <= not((layer0_outputs(252)) or (layer0_outputs(5272)));
    layer1_outputs(7266) <= layer0_outputs(761);
    layer1_outputs(7267) <= not(layer0_outputs(7005));
    layer1_outputs(7268) <= layer0_outputs(6413);
    layer1_outputs(7269) <= not(layer0_outputs(1723));
    layer1_outputs(7270) <= not(layer0_outputs(1234));
    layer1_outputs(7271) <= '1';
    layer1_outputs(7272) <= (layer0_outputs(6576)) and (layer0_outputs(743));
    layer1_outputs(7273) <= '0';
    layer1_outputs(7274) <= not(layer0_outputs(8760));
    layer1_outputs(7275) <= (layer0_outputs(7222)) and not (layer0_outputs(6105));
    layer1_outputs(7276) <= not(layer0_outputs(3027));
    layer1_outputs(7277) <= (layer0_outputs(1962)) and not (layer0_outputs(2789));
    layer1_outputs(7278) <= not(layer0_outputs(5776));
    layer1_outputs(7279) <= not(layer0_outputs(7298));
    layer1_outputs(7280) <= not((layer0_outputs(3656)) or (layer0_outputs(5294)));
    layer1_outputs(7281) <= '0';
    layer1_outputs(7282) <= not(layer0_outputs(510)) or (layer0_outputs(4704));
    layer1_outputs(7283) <= (layer0_outputs(1191)) or (layer0_outputs(6895));
    layer1_outputs(7284) <= (layer0_outputs(868)) and not (layer0_outputs(315));
    layer1_outputs(7285) <= not((layer0_outputs(2550)) and (layer0_outputs(2635)));
    layer1_outputs(7286) <= not(layer0_outputs(4382));
    layer1_outputs(7287) <= not(layer0_outputs(518));
    layer1_outputs(7288) <= not((layer0_outputs(2729)) xor (layer0_outputs(8162)));
    layer1_outputs(7289) <= (layer0_outputs(6273)) xor (layer0_outputs(6600));
    layer1_outputs(7290) <= not((layer0_outputs(9955)) or (layer0_outputs(2581)));
    layer1_outputs(7291) <= (layer0_outputs(7415)) or (layer0_outputs(4549));
    layer1_outputs(7292) <= (layer0_outputs(7641)) and not (layer0_outputs(2852));
    layer1_outputs(7293) <= not(layer0_outputs(2753));
    layer1_outputs(7294) <= (layer0_outputs(2462)) and not (layer0_outputs(8719));
    layer1_outputs(7295) <= not(layer0_outputs(1840)) or (layer0_outputs(216));
    layer1_outputs(7296) <= not(layer0_outputs(4080));
    layer1_outputs(7297) <= '1';
    layer1_outputs(7298) <= (layer0_outputs(7410)) and not (layer0_outputs(9770));
    layer1_outputs(7299) <= not((layer0_outputs(8593)) xor (layer0_outputs(6772)));
    layer1_outputs(7300) <= '1';
    layer1_outputs(7301) <= (layer0_outputs(5237)) and (layer0_outputs(2177));
    layer1_outputs(7302) <= not(layer0_outputs(5194)) or (layer0_outputs(780));
    layer1_outputs(7303) <= '1';
    layer1_outputs(7304) <= layer0_outputs(4067);
    layer1_outputs(7305) <= not(layer0_outputs(4811)) or (layer0_outputs(7309));
    layer1_outputs(7306) <= not(layer0_outputs(5572)) or (layer0_outputs(4664));
    layer1_outputs(7307) <= not(layer0_outputs(10187)) or (layer0_outputs(4922));
    layer1_outputs(7308) <= (layer0_outputs(1215)) or (layer0_outputs(5236));
    layer1_outputs(7309) <= not(layer0_outputs(8466));
    layer1_outputs(7310) <= not((layer0_outputs(6367)) xor (layer0_outputs(481)));
    layer1_outputs(7311) <= layer0_outputs(1393);
    layer1_outputs(7312) <= not((layer0_outputs(4095)) and (layer0_outputs(8833)));
    layer1_outputs(7313) <= not(layer0_outputs(3698)) or (layer0_outputs(2571));
    layer1_outputs(7314) <= '0';
    layer1_outputs(7315) <= (layer0_outputs(9754)) and not (layer0_outputs(1912));
    layer1_outputs(7316) <= '1';
    layer1_outputs(7317) <= '0';
    layer1_outputs(7318) <= not((layer0_outputs(5101)) and (layer0_outputs(2795)));
    layer1_outputs(7319) <= not((layer0_outputs(3707)) or (layer0_outputs(6795)));
    layer1_outputs(7320) <= '1';
    layer1_outputs(7321) <= (layer0_outputs(3532)) or (layer0_outputs(9035));
    layer1_outputs(7322) <= not((layer0_outputs(7311)) or (layer0_outputs(6568)));
    layer1_outputs(7323) <= (layer0_outputs(10030)) or (layer0_outputs(3791));
    layer1_outputs(7324) <= (layer0_outputs(1602)) and (layer0_outputs(1992));
    layer1_outputs(7325) <= not(layer0_outputs(2428)) or (layer0_outputs(8131));
    layer1_outputs(7326) <= not(layer0_outputs(1186));
    layer1_outputs(7327) <= not((layer0_outputs(8934)) or (layer0_outputs(9573)));
    layer1_outputs(7328) <= not((layer0_outputs(4940)) and (layer0_outputs(6658)));
    layer1_outputs(7329) <= not(layer0_outputs(10064));
    layer1_outputs(7330) <= '0';
    layer1_outputs(7331) <= (layer0_outputs(2579)) and (layer0_outputs(3313));
    layer1_outputs(7332) <= (layer0_outputs(2087)) or (layer0_outputs(4452));
    layer1_outputs(7333) <= (layer0_outputs(6876)) and not (layer0_outputs(3615));
    layer1_outputs(7334) <= not(layer0_outputs(454)) or (layer0_outputs(1402));
    layer1_outputs(7335) <= (layer0_outputs(1052)) and not (layer0_outputs(7123));
    layer1_outputs(7336) <= (layer0_outputs(67)) and not (layer0_outputs(5981));
    layer1_outputs(7337) <= '0';
    layer1_outputs(7338) <= not(layer0_outputs(2933)) or (layer0_outputs(5286));
    layer1_outputs(7339) <= not((layer0_outputs(3211)) or (layer0_outputs(639)));
    layer1_outputs(7340) <= (layer0_outputs(6974)) or (layer0_outputs(4405));
    layer1_outputs(7341) <= layer0_outputs(287);
    layer1_outputs(7342) <= (layer0_outputs(3245)) and (layer0_outputs(4758));
    layer1_outputs(7343) <= not((layer0_outputs(9448)) or (layer0_outputs(250)));
    layer1_outputs(7344) <= not((layer0_outputs(3758)) xor (layer0_outputs(6798)));
    layer1_outputs(7345) <= layer0_outputs(4246);
    layer1_outputs(7346) <= (layer0_outputs(3607)) and not (layer0_outputs(3461));
    layer1_outputs(7347) <= not(layer0_outputs(3705)) or (layer0_outputs(2199));
    layer1_outputs(7348) <= not((layer0_outputs(2273)) or (layer0_outputs(4423)));
    layer1_outputs(7349) <= not(layer0_outputs(1324));
    layer1_outputs(7350) <= not((layer0_outputs(657)) and (layer0_outputs(9757)));
    layer1_outputs(7351) <= layer0_outputs(1767);
    layer1_outputs(7352) <= not(layer0_outputs(7659)) or (layer0_outputs(7467));
    layer1_outputs(7353) <= layer0_outputs(3239);
    layer1_outputs(7354) <= not((layer0_outputs(8716)) or (layer0_outputs(6258)));
    layer1_outputs(7355) <= not(layer0_outputs(1706));
    layer1_outputs(7356) <= not(layer0_outputs(9905));
    layer1_outputs(7357) <= not((layer0_outputs(2534)) or (layer0_outputs(294)));
    layer1_outputs(7358) <= not(layer0_outputs(9402));
    layer1_outputs(7359) <= not(layer0_outputs(4600));
    layer1_outputs(7360) <= (layer0_outputs(3304)) and (layer0_outputs(5849));
    layer1_outputs(7361) <= (layer0_outputs(9556)) or (layer0_outputs(267));
    layer1_outputs(7362) <= (layer0_outputs(8653)) or (layer0_outputs(4835));
    layer1_outputs(7363) <= (layer0_outputs(1844)) or (layer0_outputs(4321));
    layer1_outputs(7364) <= not(layer0_outputs(8513));
    layer1_outputs(7365) <= (layer0_outputs(5940)) xor (layer0_outputs(322));
    layer1_outputs(7366) <= not(layer0_outputs(1960)) or (layer0_outputs(8443));
    layer1_outputs(7367) <= not((layer0_outputs(4577)) and (layer0_outputs(5974)));
    layer1_outputs(7368) <= not((layer0_outputs(2936)) and (layer0_outputs(1087)));
    layer1_outputs(7369) <= not(layer0_outputs(4348));
    layer1_outputs(7370) <= (layer0_outputs(9086)) and not (layer0_outputs(85));
    layer1_outputs(7371) <= '0';
    layer1_outputs(7372) <= not((layer0_outputs(5791)) and (layer0_outputs(8097)));
    layer1_outputs(7373) <= not((layer0_outputs(5345)) or (layer0_outputs(2715)));
    layer1_outputs(7374) <= '0';
    layer1_outputs(7375) <= not(layer0_outputs(9675));
    layer1_outputs(7376) <= layer0_outputs(3947);
    layer1_outputs(7377) <= not(layer0_outputs(1478)) or (layer0_outputs(9829));
    layer1_outputs(7378) <= not(layer0_outputs(2483));
    layer1_outputs(7379) <= layer0_outputs(3522);
    layer1_outputs(7380) <= (layer0_outputs(5256)) and (layer0_outputs(5348));
    layer1_outputs(7381) <= (layer0_outputs(3093)) and (layer0_outputs(4088));
    layer1_outputs(7382) <= not(layer0_outputs(2842)) or (layer0_outputs(7931));
    layer1_outputs(7383) <= (layer0_outputs(2665)) and not (layer0_outputs(6058));
    layer1_outputs(7384) <= not(layer0_outputs(6396));
    layer1_outputs(7385) <= (layer0_outputs(1193)) and (layer0_outputs(2900));
    layer1_outputs(7386) <= '0';
    layer1_outputs(7387) <= (layer0_outputs(9337)) xor (layer0_outputs(5840));
    layer1_outputs(7388) <= (layer0_outputs(10042)) and not (layer0_outputs(7022));
    layer1_outputs(7389) <= layer0_outputs(8943);
    layer1_outputs(7390) <= (layer0_outputs(1456)) and not (layer0_outputs(7909));
    layer1_outputs(7391) <= layer0_outputs(8290);
    layer1_outputs(7392) <= (layer0_outputs(9985)) or (layer0_outputs(7243));
    layer1_outputs(7393) <= layer0_outputs(1726);
    layer1_outputs(7394) <= not((layer0_outputs(497)) or (layer0_outputs(10175)));
    layer1_outputs(7395) <= layer0_outputs(1227);
    layer1_outputs(7396) <= layer0_outputs(9253);
    layer1_outputs(7397) <= (layer0_outputs(111)) and not (layer0_outputs(4070));
    layer1_outputs(7398) <= (layer0_outputs(4467)) and not (layer0_outputs(4733));
    layer1_outputs(7399) <= not(layer0_outputs(38)) or (layer0_outputs(7499));
    layer1_outputs(7400) <= '0';
    layer1_outputs(7401) <= '1';
    layer1_outputs(7402) <= layer0_outputs(796);
    layer1_outputs(7403) <= not(layer0_outputs(1939));
    layer1_outputs(7404) <= not((layer0_outputs(3586)) or (layer0_outputs(5737)));
    layer1_outputs(7405) <= not((layer0_outputs(706)) xor (layer0_outputs(4499)));
    layer1_outputs(7406) <= not(layer0_outputs(8868)) or (layer0_outputs(1493));
    layer1_outputs(7407) <= not((layer0_outputs(8880)) and (layer0_outputs(2250)));
    layer1_outputs(7408) <= '0';
    layer1_outputs(7409) <= (layer0_outputs(4857)) and not (layer0_outputs(5161));
    layer1_outputs(7410) <= layer0_outputs(5321);
    layer1_outputs(7411) <= '0';
    layer1_outputs(7412) <= not(layer0_outputs(10174));
    layer1_outputs(7413) <= (layer0_outputs(3682)) or (layer0_outputs(4034));
    layer1_outputs(7414) <= (layer0_outputs(226)) xor (layer0_outputs(305));
    layer1_outputs(7415) <= layer0_outputs(8128);
    layer1_outputs(7416) <= layer0_outputs(8899);
    layer1_outputs(7417) <= (layer0_outputs(8274)) and (layer0_outputs(6187));
    layer1_outputs(7418) <= not(layer0_outputs(5484));
    layer1_outputs(7419) <= (layer0_outputs(1367)) and (layer0_outputs(10178));
    layer1_outputs(7420) <= (layer0_outputs(514)) and not (layer0_outputs(3592));
    layer1_outputs(7421) <= not((layer0_outputs(4630)) and (layer0_outputs(5640)));
    layer1_outputs(7422) <= not(layer0_outputs(9530));
    layer1_outputs(7423) <= (layer0_outputs(607)) and (layer0_outputs(4956));
    layer1_outputs(7424) <= not((layer0_outputs(3945)) xor (layer0_outputs(2395)));
    layer1_outputs(7425) <= (layer0_outputs(6629)) and (layer0_outputs(7840));
    layer1_outputs(7426) <= not((layer0_outputs(1190)) or (layer0_outputs(9895)));
    layer1_outputs(7427) <= not(layer0_outputs(9323)) or (layer0_outputs(938));
    layer1_outputs(7428) <= '0';
    layer1_outputs(7429) <= (layer0_outputs(1404)) and not (layer0_outputs(1333));
    layer1_outputs(7430) <= not(layer0_outputs(8263)) or (layer0_outputs(1137));
    layer1_outputs(7431) <= not(layer0_outputs(4662));
    layer1_outputs(7432) <= not(layer0_outputs(9680));
    layer1_outputs(7433) <= not(layer0_outputs(9006)) or (layer0_outputs(1582));
    layer1_outputs(7434) <= '1';
    layer1_outputs(7435) <= not(layer0_outputs(9791)) or (layer0_outputs(8779));
    layer1_outputs(7436) <= not((layer0_outputs(1385)) or (layer0_outputs(7562)));
    layer1_outputs(7437) <= not(layer0_outputs(6427));
    layer1_outputs(7438) <= layer0_outputs(4736);
    layer1_outputs(7439) <= (layer0_outputs(1578)) or (layer0_outputs(3141));
    layer1_outputs(7440) <= not((layer0_outputs(4693)) or (layer0_outputs(3198)));
    layer1_outputs(7441) <= not(layer0_outputs(4384)) or (layer0_outputs(7516));
    layer1_outputs(7442) <= layer0_outputs(6757);
    layer1_outputs(7443) <= (layer0_outputs(10088)) and (layer0_outputs(7571));
    layer1_outputs(7444) <= not((layer0_outputs(8611)) or (layer0_outputs(5229)));
    layer1_outputs(7445) <= not(layer0_outputs(8405));
    layer1_outputs(7446) <= layer0_outputs(6978);
    layer1_outputs(7447) <= (layer0_outputs(4261)) and (layer0_outputs(4021));
    layer1_outputs(7448) <= layer0_outputs(7908);
    layer1_outputs(7449) <= (layer0_outputs(878)) and not (layer0_outputs(7328));
    layer1_outputs(7450) <= not((layer0_outputs(4942)) and (layer0_outputs(7755)));
    layer1_outputs(7451) <= (layer0_outputs(8136)) and (layer0_outputs(754));
    layer1_outputs(7452) <= layer0_outputs(4179);
    layer1_outputs(7453) <= not(layer0_outputs(5391));
    layer1_outputs(7454) <= (layer0_outputs(6882)) and not (layer0_outputs(1752));
    layer1_outputs(7455) <= not((layer0_outputs(1169)) or (layer0_outputs(3650)));
    layer1_outputs(7456) <= (layer0_outputs(5022)) xor (layer0_outputs(1964));
    layer1_outputs(7457) <= not(layer0_outputs(5825));
    layer1_outputs(7458) <= layer0_outputs(5832);
    layer1_outputs(7459) <= not(layer0_outputs(4051)) or (layer0_outputs(6414));
    layer1_outputs(7460) <= not(layer0_outputs(5685));
    layer1_outputs(7461) <= (layer0_outputs(467)) xor (layer0_outputs(819));
    layer1_outputs(7462) <= layer0_outputs(2047);
    layer1_outputs(7463) <= not((layer0_outputs(8279)) or (layer0_outputs(5313)));
    layer1_outputs(7464) <= not((layer0_outputs(8189)) and (layer0_outputs(9261)));
    layer1_outputs(7465) <= not(layer0_outputs(1086)) or (layer0_outputs(1718));
    layer1_outputs(7466) <= not((layer0_outputs(7566)) or (layer0_outputs(2165)));
    layer1_outputs(7467) <= not((layer0_outputs(9042)) and (layer0_outputs(1412)));
    layer1_outputs(7468) <= layer0_outputs(7387);
    layer1_outputs(7469) <= layer0_outputs(4020);
    layer1_outputs(7470) <= (layer0_outputs(3352)) and (layer0_outputs(9393));
    layer1_outputs(7471) <= not(layer0_outputs(1501)) or (layer0_outputs(2702));
    layer1_outputs(7472) <= not((layer0_outputs(3613)) and (layer0_outputs(2277)));
    layer1_outputs(7473) <= not(layer0_outputs(8022)) or (layer0_outputs(6987));
    layer1_outputs(7474) <= not((layer0_outputs(1294)) and (layer0_outputs(4142)));
    layer1_outputs(7475) <= not(layer0_outputs(1021));
    layer1_outputs(7476) <= layer0_outputs(6864);
    layer1_outputs(7477) <= not(layer0_outputs(8545));
    layer1_outputs(7478) <= not(layer0_outputs(481));
    layer1_outputs(7479) <= (layer0_outputs(4056)) and (layer0_outputs(5060));
    layer1_outputs(7480) <= layer0_outputs(9678);
    layer1_outputs(7481) <= layer0_outputs(184);
    layer1_outputs(7482) <= not(layer0_outputs(1080));
    layer1_outputs(7483) <= (layer0_outputs(8209)) xor (layer0_outputs(835));
    layer1_outputs(7484) <= (layer0_outputs(6169)) and not (layer0_outputs(4443));
    layer1_outputs(7485) <= layer0_outputs(10147);
    layer1_outputs(7486) <= not(layer0_outputs(9990)) or (layer0_outputs(9371));
    layer1_outputs(7487) <= (layer0_outputs(3553)) and not (layer0_outputs(8381));
    layer1_outputs(7488) <= (layer0_outputs(6484)) and (layer0_outputs(1864));
    layer1_outputs(7489) <= not(layer0_outputs(5562));
    layer1_outputs(7490) <= (layer0_outputs(4399)) xor (layer0_outputs(5135));
    layer1_outputs(7491) <= not((layer0_outputs(5234)) and (layer0_outputs(4473)));
    layer1_outputs(7492) <= not(layer0_outputs(4336)) or (layer0_outputs(3122));
    layer1_outputs(7493) <= '1';
    layer1_outputs(7494) <= '0';
    layer1_outputs(7495) <= not(layer0_outputs(7727));
    layer1_outputs(7496) <= not(layer0_outputs(2936));
    layer1_outputs(7497) <= (layer0_outputs(6648)) and (layer0_outputs(3722));
    layer1_outputs(7498) <= not((layer0_outputs(9186)) or (layer0_outputs(3250)));
    layer1_outputs(7499) <= not((layer0_outputs(9199)) and (layer0_outputs(390)));
    layer1_outputs(7500) <= not((layer0_outputs(5861)) and (layer0_outputs(100)));
    layer1_outputs(7501) <= not(layer0_outputs(5174));
    layer1_outputs(7502) <= (layer0_outputs(6379)) and not (layer0_outputs(781));
    layer1_outputs(7503) <= not(layer0_outputs(5979)) or (layer0_outputs(1690));
    layer1_outputs(7504) <= (layer0_outputs(6093)) or (layer0_outputs(4370));
    layer1_outputs(7505) <= (layer0_outputs(3098)) xor (layer0_outputs(5001));
    layer1_outputs(7506) <= not(layer0_outputs(9746)) or (layer0_outputs(6165));
    layer1_outputs(7507) <= not(layer0_outputs(3849)) or (layer0_outputs(4233));
    layer1_outputs(7508) <= not((layer0_outputs(9691)) or (layer0_outputs(3505)));
    layer1_outputs(7509) <= not((layer0_outputs(3617)) and (layer0_outputs(5711)));
    layer1_outputs(7510) <= not(layer0_outputs(5309));
    layer1_outputs(7511) <= not((layer0_outputs(7479)) or (layer0_outputs(4303)));
    layer1_outputs(7512) <= not(layer0_outputs(9381));
    layer1_outputs(7513) <= not((layer0_outputs(8202)) or (layer0_outputs(10121)));
    layer1_outputs(7514) <= not(layer0_outputs(6489));
    layer1_outputs(7515) <= '1';
    layer1_outputs(7516) <= '1';
    layer1_outputs(7517) <= layer0_outputs(3877);
    layer1_outputs(7518) <= (layer0_outputs(9065)) and (layer0_outputs(2035));
    layer1_outputs(7519) <= (layer0_outputs(6195)) and not (layer0_outputs(121));
    layer1_outputs(7520) <= not(layer0_outputs(1611)) or (layer0_outputs(8752));
    layer1_outputs(7521) <= '0';
    layer1_outputs(7522) <= '0';
    layer1_outputs(7523) <= not(layer0_outputs(3858));
    layer1_outputs(7524) <= not((layer0_outputs(1679)) or (layer0_outputs(6891)));
    layer1_outputs(7525) <= layer0_outputs(808);
    layer1_outputs(7526) <= not((layer0_outputs(4265)) xor (layer0_outputs(2188)));
    layer1_outputs(7527) <= not(layer0_outputs(2844)) or (layer0_outputs(280));
    layer1_outputs(7528) <= not(layer0_outputs(2568)) or (layer0_outputs(5271));
    layer1_outputs(7529) <= layer0_outputs(6395);
    layer1_outputs(7530) <= (layer0_outputs(4499)) and not (layer0_outputs(3715));
    layer1_outputs(7531) <= not((layer0_outputs(2219)) and (layer0_outputs(6235)));
    layer1_outputs(7532) <= not(layer0_outputs(10030));
    layer1_outputs(7533) <= not(layer0_outputs(3878)) or (layer0_outputs(1705));
    layer1_outputs(7534) <= not(layer0_outputs(6187)) or (layer0_outputs(8727));
    layer1_outputs(7535) <= layer0_outputs(6230);
    layer1_outputs(7536) <= not((layer0_outputs(4527)) xor (layer0_outputs(1067)));
    layer1_outputs(7537) <= (layer0_outputs(6794)) and not (layer0_outputs(9790));
    layer1_outputs(7538) <= (layer0_outputs(8112)) and not (layer0_outputs(5823));
    layer1_outputs(7539) <= not(layer0_outputs(7596)) or (layer0_outputs(417));
    layer1_outputs(7540) <= not(layer0_outputs(475)) or (layer0_outputs(9656));
    layer1_outputs(7541) <= (layer0_outputs(5604)) and (layer0_outputs(5504));
    layer1_outputs(7542) <= layer0_outputs(5163);
    layer1_outputs(7543) <= (layer0_outputs(2658)) or (layer0_outputs(452));
    layer1_outputs(7544) <= not((layer0_outputs(2878)) and (layer0_outputs(1099)));
    layer1_outputs(7545) <= (layer0_outputs(2538)) and not (layer0_outputs(8254));
    layer1_outputs(7546) <= not(layer0_outputs(6808));
    layer1_outputs(7547) <= (layer0_outputs(2369)) and not (layer0_outputs(9085));
    layer1_outputs(7548) <= (layer0_outputs(5488)) or (layer0_outputs(5415));
    layer1_outputs(7549) <= not((layer0_outputs(5125)) and (layer0_outputs(277)));
    layer1_outputs(7550) <= '0';
    layer1_outputs(7551) <= not(layer0_outputs(2093));
    layer1_outputs(7552) <= layer0_outputs(53);
    layer1_outputs(7553) <= not(layer0_outputs(8479));
    layer1_outputs(7554) <= layer0_outputs(7388);
    layer1_outputs(7555) <= '0';
    layer1_outputs(7556) <= not(layer0_outputs(9034));
    layer1_outputs(7557) <= '0';
    layer1_outputs(7558) <= not(layer0_outputs(4607));
    layer1_outputs(7559) <= (layer0_outputs(7343)) and not (layer0_outputs(6733));
    layer1_outputs(7560) <= not(layer0_outputs(3893));
    layer1_outputs(7561) <= not(layer0_outputs(9934));
    layer1_outputs(7562) <= (layer0_outputs(1733)) xor (layer0_outputs(5517));
    layer1_outputs(7563) <= not(layer0_outputs(8987));
    layer1_outputs(7564) <= layer0_outputs(5712);
    layer1_outputs(7565) <= layer0_outputs(8052);
    layer1_outputs(7566) <= not(layer0_outputs(9626)) or (layer0_outputs(4241));
    layer1_outputs(7567) <= (layer0_outputs(1509)) and not (layer0_outputs(4503));
    layer1_outputs(7568) <= not(layer0_outputs(1636));
    layer1_outputs(7569) <= (layer0_outputs(7202)) and not (layer0_outputs(8256));
    layer1_outputs(7570) <= (layer0_outputs(8351)) or (layer0_outputs(2356));
    layer1_outputs(7571) <= not(layer0_outputs(1949));
    layer1_outputs(7572) <= not((layer0_outputs(2908)) and (layer0_outputs(4263)));
    layer1_outputs(7573) <= (layer0_outputs(2507)) and not (layer0_outputs(7951));
    layer1_outputs(7574) <= '1';
    layer1_outputs(7575) <= not(layer0_outputs(3542)) or (layer0_outputs(2034));
    layer1_outputs(7576) <= not(layer0_outputs(511)) or (layer0_outputs(8722));
    layer1_outputs(7577) <= not(layer0_outputs(5599)) or (layer0_outputs(1775));
    layer1_outputs(7578) <= not((layer0_outputs(2067)) and (layer0_outputs(8510)));
    layer1_outputs(7579) <= not(layer0_outputs(5499)) or (layer0_outputs(2707));
    layer1_outputs(7580) <= not((layer0_outputs(2401)) xor (layer0_outputs(621)));
    layer1_outputs(7581) <= '0';
    layer1_outputs(7582) <= (layer0_outputs(9367)) or (layer0_outputs(4177));
    layer1_outputs(7583) <= not(layer0_outputs(3006)) or (layer0_outputs(7037));
    layer1_outputs(7584) <= not((layer0_outputs(9642)) and (layer0_outputs(8822)));
    layer1_outputs(7585) <= not(layer0_outputs(7796));
    layer1_outputs(7586) <= not(layer0_outputs(4578));
    layer1_outputs(7587) <= (layer0_outputs(257)) and (layer0_outputs(846));
    layer1_outputs(7588) <= (layer0_outputs(880)) and (layer0_outputs(6695));
    layer1_outputs(7589) <= (layer0_outputs(8981)) or (layer0_outputs(2469));
    layer1_outputs(7590) <= not(layer0_outputs(7236)) or (layer0_outputs(2776));
    layer1_outputs(7591) <= (layer0_outputs(9309)) and not (layer0_outputs(374));
    layer1_outputs(7592) <= not(layer0_outputs(4983)) or (layer0_outputs(3228));
    layer1_outputs(7593) <= not(layer0_outputs(2321));
    layer1_outputs(7594) <= (layer0_outputs(5636)) or (layer0_outputs(5006));
    layer1_outputs(7595) <= '1';
    layer1_outputs(7596) <= not(layer0_outputs(605)) or (layer0_outputs(6897));
    layer1_outputs(7597) <= (layer0_outputs(5522)) or (layer0_outputs(8956));
    layer1_outputs(7598) <= not((layer0_outputs(7108)) and (layer0_outputs(2339)));
    layer1_outputs(7599) <= (layer0_outputs(1476)) and not (layer0_outputs(5746));
    layer1_outputs(7600) <= not((layer0_outputs(251)) and (layer0_outputs(3677)));
    layer1_outputs(7601) <= not((layer0_outputs(7131)) and (layer0_outputs(2440)));
    layer1_outputs(7602) <= (layer0_outputs(8889)) and (layer0_outputs(4872));
    layer1_outputs(7603) <= not(layer0_outputs(8303)) or (layer0_outputs(9412));
    layer1_outputs(7604) <= not((layer0_outputs(8309)) or (layer0_outputs(6855)));
    layer1_outputs(7605) <= '0';
    layer1_outputs(7606) <= not(layer0_outputs(5243));
    layer1_outputs(7607) <= layer0_outputs(8267);
    layer1_outputs(7608) <= not(layer0_outputs(7698));
    layer1_outputs(7609) <= layer0_outputs(9134);
    layer1_outputs(7610) <= (layer0_outputs(5977)) and (layer0_outputs(9184));
    layer1_outputs(7611) <= not(layer0_outputs(8129));
    layer1_outputs(7612) <= '1';
    layer1_outputs(7613) <= not((layer0_outputs(7459)) and (layer0_outputs(3125)));
    layer1_outputs(7614) <= layer0_outputs(7213);
    layer1_outputs(7615) <= '0';
    layer1_outputs(7616) <= '1';
    layer1_outputs(7617) <= not((layer0_outputs(6686)) and (layer0_outputs(955)));
    layer1_outputs(7618) <= (layer0_outputs(1650)) and not (layer0_outputs(4324));
    layer1_outputs(7619) <= '0';
    layer1_outputs(7620) <= not((layer0_outputs(598)) or (layer0_outputs(9699)));
    layer1_outputs(7621) <= not((layer0_outputs(10228)) xor (layer0_outputs(9325)));
    layer1_outputs(7622) <= not(layer0_outputs(1968)) or (layer0_outputs(6473));
    layer1_outputs(7623) <= not((layer0_outputs(6899)) and (layer0_outputs(3493)));
    layer1_outputs(7624) <= not(layer0_outputs(7165));
    layer1_outputs(7625) <= (layer0_outputs(3281)) xor (layer0_outputs(9211));
    layer1_outputs(7626) <= layer0_outputs(1517);
    layer1_outputs(7627) <= not((layer0_outputs(4724)) or (layer0_outputs(6746)));
    layer1_outputs(7628) <= not(layer0_outputs(2885));
    layer1_outputs(7629) <= (layer0_outputs(1013)) and (layer0_outputs(5004));
    layer1_outputs(7630) <= not(layer0_outputs(3051)) or (layer0_outputs(5519));
    layer1_outputs(7631) <= (layer0_outputs(9223)) or (layer0_outputs(5166));
    layer1_outputs(7632) <= (layer0_outputs(7880)) or (layer0_outputs(7451));
    layer1_outputs(7633) <= not(layer0_outputs(7500)) or (layer0_outputs(2867));
    layer1_outputs(7634) <= '1';
    layer1_outputs(7635) <= '0';
    layer1_outputs(7636) <= (layer0_outputs(4307)) and not (layer0_outputs(3906));
    layer1_outputs(7637) <= not((layer0_outputs(6657)) or (layer0_outputs(2139)));
    layer1_outputs(7638) <= not(layer0_outputs(3409));
    layer1_outputs(7639) <= not(layer0_outputs(6948));
    layer1_outputs(7640) <= (layer0_outputs(8224)) or (layer0_outputs(2077));
    layer1_outputs(7641) <= (layer0_outputs(7701)) xor (layer0_outputs(10048));
    layer1_outputs(7642) <= not((layer0_outputs(2179)) xor (layer0_outputs(7903)));
    layer1_outputs(7643) <= '0';
    layer1_outputs(7644) <= not(layer0_outputs(5804));
    layer1_outputs(7645) <= layer0_outputs(4704);
    layer1_outputs(7646) <= '0';
    layer1_outputs(7647) <= '1';
    layer1_outputs(7648) <= layer0_outputs(8559);
    layer1_outputs(7649) <= not(layer0_outputs(7298));
    layer1_outputs(7650) <= not(layer0_outputs(5945)) or (layer0_outputs(7884));
    layer1_outputs(7651) <= (layer0_outputs(9119)) and not (layer0_outputs(8759));
    layer1_outputs(7652) <= layer0_outputs(8527);
    layer1_outputs(7653) <= not((layer0_outputs(7719)) or (layer0_outputs(1107)));
    layer1_outputs(7654) <= (layer0_outputs(8029)) or (layer0_outputs(6722));
    layer1_outputs(7655) <= not(layer0_outputs(9173)) or (layer0_outputs(9609));
    layer1_outputs(7656) <= not(layer0_outputs(6173));
    layer1_outputs(7657) <= (layer0_outputs(7043)) and not (layer0_outputs(5682));
    layer1_outputs(7658) <= not((layer0_outputs(3420)) or (layer0_outputs(2944)));
    layer1_outputs(7659) <= (layer0_outputs(3054)) and (layer0_outputs(3316));
    layer1_outputs(7660) <= '1';
    layer1_outputs(7661) <= not((layer0_outputs(4390)) and (layer0_outputs(5118)));
    layer1_outputs(7662) <= (layer0_outputs(1457)) and not (layer0_outputs(6607));
    layer1_outputs(7663) <= (layer0_outputs(4420)) and (layer0_outputs(6060));
    layer1_outputs(7664) <= not(layer0_outputs(9588)) or (layer0_outputs(2515));
    layer1_outputs(7665) <= not(layer0_outputs(2186));
    layer1_outputs(7666) <= layer0_outputs(7137);
    layer1_outputs(7667) <= '1';
    layer1_outputs(7668) <= not((layer0_outputs(7377)) xor (layer0_outputs(700)));
    layer1_outputs(7669) <= not((layer0_outputs(8280)) xor (layer0_outputs(7554)));
    layer1_outputs(7670) <= not(layer0_outputs(93)) or (layer0_outputs(7661));
    layer1_outputs(7671) <= layer0_outputs(4960);
    layer1_outputs(7672) <= (layer0_outputs(6746)) and (layer0_outputs(8805));
    layer1_outputs(7673) <= '0';
    layer1_outputs(7674) <= not(layer0_outputs(4872));
    layer1_outputs(7675) <= (layer0_outputs(1293)) and not (layer0_outputs(9973));
    layer1_outputs(7676) <= not(layer0_outputs(2930));
    layer1_outputs(7677) <= not((layer0_outputs(9091)) xor (layer0_outputs(1888)));
    layer1_outputs(7678) <= not(layer0_outputs(9125));
    layer1_outputs(7679) <= '0';
    layer1_outputs(7680) <= layer0_outputs(2934);
    layer1_outputs(7681) <= layer0_outputs(5632);
    layer1_outputs(7682) <= not(layer0_outputs(10224));
    layer1_outputs(7683) <= not((layer0_outputs(8121)) xor (layer0_outputs(1804)));
    layer1_outputs(7684) <= (layer0_outputs(7543)) and not (layer0_outputs(4375));
    layer1_outputs(7685) <= '0';
    layer1_outputs(7686) <= layer0_outputs(588);
    layer1_outputs(7687) <= not(layer0_outputs(4708));
    layer1_outputs(7688) <= '0';
    layer1_outputs(7689) <= layer0_outputs(312);
    layer1_outputs(7690) <= not((layer0_outputs(5593)) or (layer0_outputs(6186)));
    layer1_outputs(7691) <= (layer0_outputs(4670)) or (layer0_outputs(8244));
    layer1_outputs(7692) <= (layer0_outputs(7942)) and (layer0_outputs(6103));
    layer1_outputs(7693) <= (layer0_outputs(4098)) or (layer0_outputs(4395));
    layer1_outputs(7694) <= not(layer0_outputs(6592));
    layer1_outputs(7695) <= not((layer0_outputs(5411)) and (layer0_outputs(4488)));
    layer1_outputs(7696) <= not(layer0_outputs(1184));
    layer1_outputs(7697) <= not((layer0_outputs(6322)) or (layer0_outputs(745)));
    layer1_outputs(7698) <= layer0_outputs(2316);
    layer1_outputs(7699) <= (layer0_outputs(3580)) or (layer0_outputs(9380));
    layer1_outputs(7700) <= not(layer0_outputs(6432)) or (layer0_outputs(7583));
    layer1_outputs(7701) <= not(layer0_outputs(7969)) or (layer0_outputs(1276));
    layer1_outputs(7702) <= not(layer0_outputs(7444));
    layer1_outputs(7703) <= (layer0_outputs(1675)) or (layer0_outputs(3620));
    layer1_outputs(7704) <= (layer0_outputs(4076)) or (layer0_outputs(5128));
    layer1_outputs(7705) <= layer0_outputs(2301);
    layer1_outputs(7706) <= '0';
    layer1_outputs(7707) <= (layer0_outputs(7660)) and (layer0_outputs(1231));
    layer1_outputs(7708) <= not(layer0_outputs(8872)) or (layer0_outputs(5926));
    layer1_outputs(7709) <= not(layer0_outputs(8345));
    layer1_outputs(7710) <= not((layer0_outputs(7397)) and (layer0_outputs(954)));
    layer1_outputs(7711) <= (layer0_outputs(2738)) and (layer0_outputs(3908));
    layer1_outputs(7712) <= not(layer0_outputs(6815));
    layer1_outputs(7713) <= (layer0_outputs(8964)) and not (layer0_outputs(6289));
    layer1_outputs(7714) <= '1';
    layer1_outputs(7715) <= (layer0_outputs(10050)) or (layer0_outputs(4305));
    layer1_outputs(7716) <= not(layer0_outputs(7883));
    layer1_outputs(7717) <= layer0_outputs(4198);
    layer1_outputs(7718) <= layer0_outputs(4889);
    layer1_outputs(7719) <= '0';
    layer1_outputs(7720) <= not(layer0_outputs(6615)) or (layer0_outputs(3510));
    layer1_outputs(7721) <= layer0_outputs(8139);
    layer1_outputs(7722) <= not((layer0_outputs(4442)) or (layer0_outputs(7210)));
    layer1_outputs(7723) <= layer0_outputs(7139);
    layer1_outputs(7724) <= not((layer0_outputs(9164)) xor (layer0_outputs(8492)));
    layer1_outputs(7725) <= not(layer0_outputs(3478));
    layer1_outputs(7726) <= (layer0_outputs(296)) xor (layer0_outputs(60));
    layer1_outputs(7727) <= not(layer0_outputs(2389));
    layer1_outputs(7728) <= '0';
    layer1_outputs(7729) <= not(layer0_outputs(5689));
    layer1_outputs(7730) <= not((layer0_outputs(7095)) xor (layer0_outputs(4918)));
    layer1_outputs(7731) <= not(layer0_outputs(154));
    layer1_outputs(7732) <= not((layer0_outputs(2030)) or (layer0_outputs(10234)));
    layer1_outputs(7733) <= layer0_outputs(9690);
    layer1_outputs(7734) <= not(layer0_outputs(6424));
    layer1_outputs(7735) <= not(layer0_outputs(2666)) or (layer0_outputs(2080));
    layer1_outputs(7736) <= not(layer0_outputs(5607)) or (layer0_outputs(6832));
    layer1_outputs(7737) <= not(layer0_outputs(4470)) or (layer0_outputs(8755));
    layer1_outputs(7738) <= not((layer0_outputs(3862)) xor (layer0_outputs(7587)));
    layer1_outputs(7739) <= layer0_outputs(1730);
    layer1_outputs(7740) <= (layer0_outputs(993)) and not (layer0_outputs(8430));
    layer1_outputs(7741) <= (layer0_outputs(6275)) xor (layer0_outputs(3565));
    layer1_outputs(7742) <= not(layer0_outputs(9442));
    layer1_outputs(7743) <= not((layer0_outputs(357)) or (layer0_outputs(7507)));
    layer1_outputs(7744) <= not(layer0_outputs(5435));
    layer1_outputs(7745) <= (layer0_outputs(2445)) or (layer0_outputs(3819));
    layer1_outputs(7746) <= not((layer0_outputs(601)) xor (layer0_outputs(4086)));
    layer1_outputs(7747) <= '1';
    layer1_outputs(7748) <= not(layer0_outputs(9395)) or (layer0_outputs(7132));
    layer1_outputs(7749) <= (layer0_outputs(1911)) or (layer0_outputs(6569));
    layer1_outputs(7750) <= layer0_outputs(5533);
    layer1_outputs(7751) <= not(layer0_outputs(8146));
    layer1_outputs(7752) <= '1';
    layer1_outputs(7753) <= not(layer0_outputs(2778));
    layer1_outputs(7754) <= '0';
    layer1_outputs(7755) <= layer0_outputs(8350);
    layer1_outputs(7756) <= '0';
    layer1_outputs(7757) <= layer0_outputs(2704);
    layer1_outputs(7758) <= not(layer0_outputs(5410));
    layer1_outputs(7759) <= not(layer0_outputs(9247)) or (layer0_outputs(4444));
    layer1_outputs(7760) <= not(layer0_outputs(1420));
    layer1_outputs(7761) <= layer0_outputs(5868);
    layer1_outputs(7762) <= not((layer0_outputs(9661)) and (layer0_outputs(9844)));
    layer1_outputs(7763) <= not(layer0_outputs(3026));
    layer1_outputs(7764) <= not(layer0_outputs(3176));
    layer1_outputs(7765) <= (layer0_outputs(6259)) xor (layer0_outputs(1111));
    layer1_outputs(7766) <= not(layer0_outputs(2365)) or (layer0_outputs(957));
    layer1_outputs(7767) <= not(layer0_outputs(9817)) or (layer0_outputs(1672));
    layer1_outputs(7768) <= layer0_outputs(8764);
    layer1_outputs(7769) <= (layer0_outputs(7525)) or (layer0_outputs(5290));
    layer1_outputs(7770) <= not(layer0_outputs(8552)) or (layer0_outputs(6583));
    layer1_outputs(7771) <= not(layer0_outputs(2421));
    layer1_outputs(7772) <= '1';
    layer1_outputs(7773) <= not((layer0_outputs(10138)) or (layer0_outputs(8640)));
    layer1_outputs(7774) <= layer0_outputs(4470);
    layer1_outputs(7775) <= layer0_outputs(484);
    layer1_outputs(7776) <= (layer0_outputs(7996)) or (layer0_outputs(344));
    layer1_outputs(7777) <= (layer0_outputs(443)) and not (layer0_outputs(1889));
    layer1_outputs(7778) <= not(layer0_outputs(2264));
    layer1_outputs(7779) <= layer0_outputs(6674);
    layer1_outputs(7780) <= not((layer0_outputs(7693)) and (layer0_outputs(415)));
    layer1_outputs(7781) <= (layer0_outputs(7151)) and (layer0_outputs(10239));
    layer1_outputs(7782) <= not((layer0_outputs(9093)) xor (layer0_outputs(5463)));
    layer1_outputs(7783) <= layer0_outputs(5646);
    layer1_outputs(7784) <= not(layer0_outputs(3464));
    layer1_outputs(7785) <= layer0_outputs(7237);
    layer1_outputs(7786) <= not(layer0_outputs(2289));
    layer1_outputs(7787) <= layer0_outputs(8340);
    layer1_outputs(7788) <= not((layer0_outputs(9586)) or (layer0_outputs(1741)));
    layer1_outputs(7789) <= not(layer0_outputs(4706)) or (layer0_outputs(6931));
    layer1_outputs(7790) <= (layer0_outputs(10134)) xor (layer0_outputs(5457));
    layer1_outputs(7791) <= not((layer0_outputs(9300)) and (layer0_outputs(9758)));
    layer1_outputs(7792) <= (layer0_outputs(6817)) or (layer0_outputs(10005));
    layer1_outputs(7793) <= layer0_outputs(4343);
    layer1_outputs(7794) <= not(layer0_outputs(8736));
    layer1_outputs(7795) <= not((layer0_outputs(9306)) and (layer0_outputs(1588)));
    layer1_outputs(7796) <= not(layer0_outputs(6735));
    layer1_outputs(7797) <= not(layer0_outputs(2528));
    layer1_outputs(7798) <= not((layer0_outputs(9920)) and (layer0_outputs(6597)));
    layer1_outputs(7799) <= layer0_outputs(5891);
    layer1_outputs(7800) <= (layer0_outputs(3960)) and not (layer0_outputs(4413));
    layer1_outputs(7801) <= layer0_outputs(3423);
    layer1_outputs(7802) <= not(layer0_outputs(8302));
    layer1_outputs(7803) <= '0';
    layer1_outputs(7804) <= '0';
    layer1_outputs(7805) <= not((layer0_outputs(4620)) and (layer0_outputs(4495)));
    layer1_outputs(7806) <= layer0_outputs(4656);
    layer1_outputs(7807) <= not(layer0_outputs(8976));
    layer1_outputs(7808) <= layer0_outputs(9113);
    layer1_outputs(7809) <= layer0_outputs(2097);
    layer1_outputs(7810) <= not((layer0_outputs(1698)) or (layer0_outputs(1490)));
    layer1_outputs(7811) <= (layer0_outputs(7983)) xor (layer0_outputs(1121));
    layer1_outputs(7812) <= (layer0_outputs(7756)) or (layer0_outputs(5528));
    layer1_outputs(7813) <= (layer0_outputs(170)) and (layer0_outputs(6680));
    layer1_outputs(7814) <= (layer0_outputs(3949)) and not (layer0_outputs(3437));
    layer1_outputs(7815) <= (layer0_outputs(3128)) or (layer0_outputs(3276));
    layer1_outputs(7816) <= (layer0_outputs(2848)) and not (layer0_outputs(7890));
    layer1_outputs(7817) <= not(layer0_outputs(5086));
    layer1_outputs(7818) <= layer0_outputs(7578);
    layer1_outputs(7819) <= layer0_outputs(1224);
    layer1_outputs(7820) <= not(layer0_outputs(2559));
    layer1_outputs(7821) <= layer0_outputs(4237);
    layer1_outputs(7822) <= not(layer0_outputs(5366)) or (layer0_outputs(5736));
    layer1_outputs(7823) <= (layer0_outputs(6388)) or (layer0_outputs(3574));
    layer1_outputs(7824) <= layer0_outputs(4262);
    layer1_outputs(7825) <= not(layer0_outputs(7523));
    layer1_outputs(7826) <= (layer0_outputs(161)) and (layer0_outputs(9259));
    layer1_outputs(7827) <= layer0_outputs(2802);
    layer1_outputs(7828) <= layer0_outputs(284);
    layer1_outputs(7829) <= (layer0_outputs(1161)) and (layer0_outputs(887));
    layer1_outputs(7830) <= not(layer0_outputs(9745)) or (layer0_outputs(520));
    layer1_outputs(7831) <= not((layer0_outputs(5710)) xor (layer0_outputs(6181)));
    layer1_outputs(7832) <= not((layer0_outputs(9257)) and (layer0_outputs(113)));
    layer1_outputs(7833) <= not(layer0_outputs(645));
    layer1_outputs(7834) <= (layer0_outputs(1592)) and not (layer0_outputs(5445));
    layer1_outputs(7835) <= layer0_outputs(8141);
    layer1_outputs(7836) <= layer0_outputs(3815);
    layer1_outputs(7837) <= layer0_outputs(3580);
    layer1_outputs(7838) <= not((layer0_outputs(9020)) xor (layer0_outputs(1820)));
    layer1_outputs(7839) <= (layer0_outputs(2858)) and not (layer0_outputs(6390));
    layer1_outputs(7840) <= (layer0_outputs(5141)) and not (layer0_outputs(5629));
    layer1_outputs(7841) <= '1';
    layer1_outputs(7842) <= not(layer0_outputs(946)) or (layer0_outputs(494));
    layer1_outputs(7843) <= layer0_outputs(4374);
    layer1_outputs(7844) <= not(layer0_outputs(10224));
    layer1_outputs(7845) <= not(layer0_outputs(1443)) or (layer0_outputs(4560));
    layer1_outputs(7846) <= not(layer0_outputs(2126));
    layer1_outputs(7847) <= (layer0_outputs(7256)) and not (layer0_outputs(7610));
    layer1_outputs(7848) <= layer0_outputs(8614);
    layer1_outputs(7849) <= not(layer0_outputs(4057));
    layer1_outputs(7850) <= '1';
    layer1_outputs(7851) <= '1';
    layer1_outputs(7852) <= not(layer0_outputs(2333));
    layer1_outputs(7853) <= (layer0_outputs(8724)) and not (layer0_outputs(7874));
    layer1_outputs(7854) <= not(layer0_outputs(9935)) or (layer0_outputs(5500));
    layer1_outputs(7855) <= not((layer0_outputs(9710)) or (layer0_outputs(9826)));
    layer1_outputs(7856) <= not(layer0_outputs(970));
    layer1_outputs(7857) <= not(layer0_outputs(4150));
    layer1_outputs(7858) <= (layer0_outputs(9415)) and not (layer0_outputs(4756));
    layer1_outputs(7859) <= not((layer0_outputs(8569)) xor (layer0_outputs(1747)));
    layer1_outputs(7860) <= not(layer0_outputs(848));
    layer1_outputs(7861) <= '0';
    layer1_outputs(7862) <= (layer0_outputs(5735)) and not (layer0_outputs(3190));
    layer1_outputs(7863) <= not(layer0_outputs(6408));
    layer1_outputs(7864) <= (layer0_outputs(7624)) or (layer0_outputs(355));
    layer1_outputs(7865) <= not((layer0_outputs(9051)) xor (layer0_outputs(2450)));
    layer1_outputs(7866) <= layer0_outputs(4308);
    layer1_outputs(7867) <= not(layer0_outputs(2352)) or (layer0_outputs(4315));
    layer1_outputs(7868) <= (layer0_outputs(7618)) and not (layer0_outputs(7033));
    layer1_outputs(7869) <= not((layer0_outputs(4626)) or (layer0_outputs(2827)));
    layer1_outputs(7870) <= (layer0_outputs(3267)) and (layer0_outputs(2615));
    layer1_outputs(7871) <= not(layer0_outputs(8326));
    layer1_outputs(7872) <= (layer0_outputs(2459)) and not (layer0_outputs(5254));
    layer1_outputs(7873) <= not(layer0_outputs(180)) or (layer0_outputs(6355));
    layer1_outputs(7874) <= not((layer0_outputs(1914)) and (layer0_outputs(5576)));
    layer1_outputs(7875) <= not(layer0_outputs(5797)) or (layer0_outputs(3216));
    layer1_outputs(7876) <= layer0_outputs(9215);
    layer1_outputs(7877) <= not(layer0_outputs(3894)) or (layer0_outputs(5553));
    layer1_outputs(7878) <= not((layer0_outputs(898)) and (layer0_outputs(6180)));
    layer1_outputs(7879) <= (layer0_outputs(2899)) and not (layer0_outputs(7651));
    layer1_outputs(7880) <= not(layer0_outputs(5470));
    layer1_outputs(7881) <= (layer0_outputs(2810)) and not (layer0_outputs(9212));
    layer1_outputs(7882) <= not((layer0_outputs(7496)) or (layer0_outputs(9333)));
    layer1_outputs(7883) <= not((layer0_outputs(2985)) and (layer0_outputs(7625)));
    layer1_outputs(7884) <= (layer0_outputs(3881)) xor (layer0_outputs(4540));
    layer1_outputs(7885) <= not(layer0_outputs(1918));
    layer1_outputs(7886) <= not(layer0_outputs(6840)) or (layer0_outputs(976));
    layer1_outputs(7887) <= '0';
    layer1_outputs(7888) <= not(layer0_outputs(10058));
    layer1_outputs(7889) <= not((layer0_outputs(183)) and (layer0_outputs(8515)));
    layer1_outputs(7890) <= layer0_outputs(455);
    layer1_outputs(7891) <= not(layer0_outputs(5106)) or (layer0_outputs(2996));
    layer1_outputs(7892) <= (layer0_outputs(1780)) or (layer0_outputs(7934));
    layer1_outputs(7893) <= (layer0_outputs(2370)) and (layer0_outputs(130));
    layer1_outputs(7894) <= not(layer0_outputs(2773));
    layer1_outputs(7895) <= not((layer0_outputs(759)) and (layer0_outputs(5152)));
    layer1_outputs(7896) <= layer0_outputs(6242);
    layer1_outputs(7897) <= layer0_outputs(1448);
    layer1_outputs(7898) <= not((layer0_outputs(9019)) xor (layer0_outputs(705)));
    layer1_outputs(7899) <= not(layer0_outputs(9639));
    layer1_outputs(7900) <= not(layer0_outputs(1922)) or (layer0_outputs(9375));
    layer1_outputs(7901) <= layer0_outputs(476);
    layer1_outputs(7902) <= (layer0_outputs(6363)) or (layer0_outputs(311));
    layer1_outputs(7903) <= not(layer0_outputs(4446));
    layer1_outputs(7904) <= not(layer0_outputs(546)) or (layer0_outputs(4562));
    layer1_outputs(7905) <= '1';
    layer1_outputs(7906) <= not(layer0_outputs(1765));
    layer1_outputs(7907) <= not(layer0_outputs(2669));
    layer1_outputs(7908) <= (layer0_outputs(8798)) and (layer0_outputs(2928));
    layer1_outputs(7909) <= (layer0_outputs(6453)) or (layer0_outputs(6234));
    layer1_outputs(7910) <= (layer0_outputs(9901)) and not (layer0_outputs(4456));
    layer1_outputs(7911) <= not((layer0_outputs(4799)) and (layer0_outputs(69)));
    layer1_outputs(7912) <= '0';
    layer1_outputs(7913) <= (layer0_outputs(8096)) or (layer0_outputs(526));
    layer1_outputs(7914) <= layer0_outputs(5243);
    layer1_outputs(7915) <= not(layer0_outputs(2166));
    layer1_outputs(7916) <= not((layer0_outputs(7780)) or (layer0_outputs(7813)));
    layer1_outputs(7917) <= '1';
    layer1_outputs(7918) <= not(layer0_outputs(3117));
    layer1_outputs(7919) <= not(layer0_outputs(2554)) or (layer0_outputs(3653));
    layer1_outputs(7920) <= layer0_outputs(1016);
    layer1_outputs(7921) <= (layer0_outputs(4352)) and not (layer0_outputs(1249));
    layer1_outputs(7922) <= not(layer0_outputs(9531));
    layer1_outputs(7923) <= not((layer0_outputs(7591)) or (layer0_outputs(3050)));
    layer1_outputs(7924) <= not(layer0_outputs(5925));
    layer1_outputs(7925) <= '0';
    layer1_outputs(7926) <= not((layer0_outputs(5478)) or (layer0_outputs(10167)));
    layer1_outputs(7927) <= (layer0_outputs(4455)) and (layer0_outputs(7204));
    layer1_outputs(7928) <= not(layer0_outputs(2437));
    layer1_outputs(7929) <= (layer0_outputs(8771)) xor (layer0_outputs(7421));
    layer1_outputs(7930) <= (layer0_outputs(3471)) and (layer0_outputs(6389));
    layer1_outputs(7931) <= not((layer0_outputs(1295)) or (layer0_outputs(2251)));
    layer1_outputs(7932) <= layer0_outputs(9342);
    layer1_outputs(7933) <= (layer0_outputs(2392)) xor (layer0_outputs(8801));
    layer1_outputs(7934) <= (layer0_outputs(9827)) and not (layer0_outputs(2938));
    layer1_outputs(7935) <= not(layer0_outputs(3311)) or (layer0_outputs(4001));
    layer1_outputs(7936) <= layer0_outputs(9927);
    layer1_outputs(7937) <= '1';
    layer1_outputs(7938) <= '0';
    layer1_outputs(7939) <= not((layer0_outputs(4476)) or (layer0_outputs(8325)));
    layer1_outputs(7940) <= (layer0_outputs(5242)) xor (layer0_outputs(8225));
    layer1_outputs(7941) <= layer0_outputs(3950);
    layer1_outputs(7942) <= not(layer0_outputs(5660));
    layer1_outputs(7943) <= not((layer0_outputs(10067)) or (layer0_outputs(8550)));
    layer1_outputs(7944) <= (layer0_outputs(10177)) and not (layer0_outputs(9146));
    layer1_outputs(7945) <= (layer0_outputs(8426)) and not (layer0_outputs(1940));
    layer1_outputs(7946) <= layer0_outputs(7737);
    layer1_outputs(7947) <= (layer0_outputs(2186)) and not (layer0_outputs(5042));
    layer1_outputs(7948) <= '0';
    layer1_outputs(7949) <= not(layer0_outputs(4224));
    layer1_outputs(7950) <= not(layer0_outputs(8572));
    layer1_outputs(7951) <= not(layer0_outputs(4330));
    layer1_outputs(7952) <= layer0_outputs(8985);
    layer1_outputs(7953) <= layer0_outputs(6533);
    layer1_outputs(7954) <= (layer0_outputs(9279)) and (layer0_outputs(9113));
    layer1_outputs(7955) <= (layer0_outputs(5158)) and (layer0_outputs(2424));
    layer1_outputs(7956) <= (layer0_outputs(4248)) or (layer0_outputs(2886));
    layer1_outputs(7957) <= (layer0_outputs(8956)) or (layer0_outputs(2160));
    layer1_outputs(7958) <= not(layer0_outputs(4590));
    layer1_outputs(7959) <= layer0_outputs(1674);
    layer1_outputs(7960) <= not(layer0_outputs(9756));
    layer1_outputs(7961) <= not(layer0_outputs(4409)) or (layer0_outputs(8681));
    layer1_outputs(7962) <= (layer0_outputs(4253)) and (layer0_outputs(5307));
    layer1_outputs(7963) <= '1';
    layer1_outputs(7964) <= (layer0_outputs(5687)) and not (layer0_outputs(7893));
    layer1_outputs(7965) <= (layer0_outputs(408)) or (layer0_outputs(1581));
    layer1_outputs(7966) <= (layer0_outputs(9584)) and not (layer0_outputs(2454));
    layer1_outputs(7967) <= not((layer0_outputs(4689)) and (layer0_outputs(1221)));
    layer1_outputs(7968) <= layer0_outputs(8538);
    layer1_outputs(7969) <= not((layer0_outputs(8509)) xor (layer0_outputs(7305)));
    layer1_outputs(7970) <= not(layer0_outputs(3857)) or (layer0_outputs(2219));
    layer1_outputs(7971) <= layer0_outputs(5187);
    layer1_outputs(7972) <= layer0_outputs(4634);
    layer1_outputs(7973) <= not(layer0_outputs(6065));
    layer1_outputs(7974) <= not(layer0_outputs(8655)) or (layer0_outputs(1453));
    layer1_outputs(7975) <= not(layer0_outputs(4667));
    layer1_outputs(7976) <= not(layer0_outputs(7115));
    layer1_outputs(7977) <= (layer0_outputs(325)) and not (layer0_outputs(1168));
    layer1_outputs(7978) <= '0';
    layer1_outputs(7979) <= '1';
    layer1_outputs(7980) <= not(layer0_outputs(9192)) or (layer0_outputs(4163));
    layer1_outputs(7981) <= not(layer0_outputs(5392)) or (layer0_outputs(8160));
    layer1_outputs(7982) <= not(layer0_outputs(2589)) or (layer0_outputs(665));
    layer1_outputs(7983) <= not(layer0_outputs(6974));
    layer1_outputs(7984) <= (layer0_outputs(6620)) or (layer0_outputs(7041));
    layer1_outputs(7985) <= '1';
    layer1_outputs(7986) <= layer0_outputs(4347);
    layer1_outputs(7987) <= layer0_outputs(4225);
    layer1_outputs(7988) <= not(layer0_outputs(1450)) or (layer0_outputs(4422));
    layer1_outputs(7989) <= (layer0_outputs(5557)) and (layer0_outputs(631));
    layer1_outputs(7990) <= (layer0_outputs(9875)) or (layer0_outputs(4301));
    layer1_outputs(7991) <= not(layer0_outputs(2856));
    layer1_outputs(7992) <= not(layer0_outputs(2006));
    layer1_outputs(7993) <= not(layer0_outputs(5512)) or (layer0_outputs(2918));
    layer1_outputs(7994) <= not((layer0_outputs(7752)) or (layer0_outputs(7809)));
    layer1_outputs(7995) <= not((layer0_outputs(8870)) and (layer0_outputs(820)));
    layer1_outputs(7996) <= (layer0_outputs(744)) and (layer0_outputs(1058));
    layer1_outputs(7997) <= (layer0_outputs(2124)) and not (layer0_outputs(8048));
    layer1_outputs(7998) <= not((layer0_outputs(6621)) or (layer0_outputs(46)));
    layer1_outputs(7999) <= not(layer0_outputs(6532));
    layer1_outputs(8000) <= layer0_outputs(1721);
    layer1_outputs(8001) <= layer0_outputs(3459);
    layer1_outputs(8002) <= not(layer0_outputs(7645));
    layer1_outputs(8003) <= (layer0_outputs(6524)) and not (layer0_outputs(9718));
    layer1_outputs(8004) <= (layer0_outputs(55)) and (layer0_outputs(7573));
    layer1_outputs(8005) <= (layer0_outputs(4867)) and (layer0_outputs(638));
    layer1_outputs(8006) <= (layer0_outputs(5369)) and (layer0_outputs(4909));
    layer1_outputs(8007) <= layer0_outputs(548);
    layer1_outputs(8008) <= '1';
    layer1_outputs(8009) <= not(layer0_outputs(10029)) or (layer0_outputs(8104));
    layer1_outputs(8010) <= layer0_outputs(8836);
    layer1_outputs(8011) <= layer0_outputs(6669);
    layer1_outputs(8012) <= not(layer0_outputs(9688));
    layer1_outputs(8013) <= not(layer0_outputs(7225)) or (layer0_outputs(7915));
    layer1_outputs(8014) <= (layer0_outputs(2843)) or (layer0_outputs(4545));
    layer1_outputs(8015) <= '1';
    layer1_outputs(8016) <= (layer0_outputs(8620)) and (layer0_outputs(7247));
    layer1_outputs(8017) <= not((layer0_outputs(1948)) or (layer0_outputs(1806)));
    layer1_outputs(8018) <= (layer0_outputs(9420)) or (layer0_outputs(5376));
    layer1_outputs(8019) <= not((layer0_outputs(3980)) and (layer0_outputs(1214)));
    layer1_outputs(8020) <= not((layer0_outputs(8511)) or (layer0_outputs(3966)));
    layer1_outputs(8021) <= not(layer0_outputs(9798)) or (layer0_outputs(1925));
    layer1_outputs(8022) <= (layer0_outputs(1259)) and not (layer0_outputs(8179));
    layer1_outputs(8023) <= (layer0_outputs(4130)) or (layer0_outputs(5330));
    layer1_outputs(8024) <= (layer0_outputs(7223)) xor (layer0_outputs(295));
    layer1_outputs(8025) <= layer0_outputs(4152);
    layer1_outputs(8026) <= (layer0_outputs(2095)) or (layer0_outputs(5557));
    layer1_outputs(8027) <= not(layer0_outputs(2946)) or (layer0_outputs(3338));
    layer1_outputs(8028) <= not((layer0_outputs(2171)) or (layer0_outputs(7000)));
    layer1_outputs(8029) <= '0';
    layer1_outputs(8030) <= layer0_outputs(4927);
    layer1_outputs(8031) <= not(layer0_outputs(7027)) or (layer0_outputs(6659));
    layer1_outputs(8032) <= not(layer0_outputs(1363)) or (layer0_outputs(2864));
    layer1_outputs(8033) <= '1';
    layer1_outputs(8034) <= (layer0_outputs(1892)) and not (layer0_outputs(613));
    layer1_outputs(8035) <= not(layer0_outputs(874));
    layer1_outputs(8036) <= not(layer0_outputs(2725));
    layer1_outputs(8037) <= not((layer0_outputs(3761)) or (layer0_outputs(2793)));
    layer1_outputs(8038) <= not((layer0_outputs(2699)) and (layer0_outputs(1848)));
    layer1_outputs(8039) <= not((layer0_outputs(5775)) or (layer0_outputs(349)));
    layer1_outputs(8040) <= not(layer0_outputs(5109));
    layer1_outputs(8041) <= not((layer0_outputs(9746)) and (layer0_outputs(7616)));
    layer1_outputs(8042) <= '1';
    layer1_outputs(8043) <= not(layer0_outputs(2882)) or (layer0_outputs(4937));
    layer1_outputs(8044) <= (layer0_outputs(8500)) and not (layer0_outputs(9166));
    layer1_outputs(8045) <= '1';
    layer1_outputs(8046) <= (layer0_outputs(8534)) and not (layer0_outputs(8781));
    layer1_outputs(8047) <= not((layer0_outputs(2526)) xor (layer0_outputs(8590)));
    layer1_outputs(8048) <= not((layer0_outputs(3782)) and (layer0_outputs(2695)));
    layer1_outputs(8049) <= layer0_outputs(5835);
    layer1_outputs(8050) <= not(layer0_outputs(4667)) or (layer0_outputs(5100));
    layer1_outputs(8051) <= not(layer0_outputs(3151)) or (layer0_outputs(4132));
    layer1_outputs(8052) <= not(layer0_outputs(4559));
    layer1_outputs(8053) <= not(layer0_outputs(6091));
    layer1_outputs(8054) <= not((layer0_outputs(2070)) and (layer0_outputs(7971)));
    layer1_outputs(8055) <= '1';
    layer1_outputs(8056) <= not(layer0_outputs(9490));
    layer1_outputs(8057) <= not(layer0_outputs(3419));
    layer1_outputs(8058) <= layer0_outputs(2158);
    layer1_outputs(8059) <= not((layer0_outputs(9151)) or (layer0_outputs(10057)));
    layer1_outputs(8060) <= (layer0_outputs(9989)) and (layer0_outputs(1612));
    layer1_outputs(8061) <= not(layer0_outputs(2728));
    layer1_outputs(8062) <= (layer0_outputs(2993)) and not (layer0_outputs(7533));
    layer1_outputs(8063) <= not(layer0_outputs(9717));
    layer1_outputs(8064) <= (layer0_outputs(9168)) and (layer0_outputs(8583));
    layer1_outputs(8065) <= '1';
    layer1_outputs(8066) <= not((layer0_outputs(6928)) xor (layer0_outputs(9254)));
    layer1_outputs(8067) <= '0';
    layer1_outputs(8068) <= not((layer0_outputs(9189)) or (layer0_outputs(3963)));
    layer1_outputs(8069) <= not((layer0_outputs(4908)) xor (layer0_outputs(1264)));
    layer1_outputs(8070) <= layer0_outputs(3948);
    layer1_outputs(8071) <= not(layer0_outputs(3165)) or (layer0_outputs(8682));
    layer1_outputs(8072) <= (layer0_outputs(7579)) or (layer0_outputs(2808));
    layer1_outputs(8073) <= not((layer0_outputs(441)) xor (layer0_outputs(7871)));
    layer1_outputs(8074) <= (layer0_outputs(561)) or (layer0_outputs(7513));
    layer1_outputs(8075) <= layer0_outputs(9153);
    layer1_outputs(8076) <= not(layer0_outputs(3587));
    layer1_outputs(8077) <= layer0_outputs(4481);
    layer1_outputs(8078) <= not((layer0_outputs(4980)) xor (layer0_outputs(9360)));
    layer1_outputs(8079) <= (layer0_outputs(1285)) and not (layer0_outputs(1854));
    layer1_outputs(8080) <= (layer0_outputs(10052)) and not (layer0_outputs(9473));
    layer1_outputs(8081) <= (layer0_outputs(5627)) and (layer0_outputs(5515));
    layer1_outputs(8082) <= '0';
    layer1_outputs(8083) <= layer0_outputs(1112);
    layer1_outputs(8084) <= not(layer0_outputs(5143));
    layer1_outputs(8085) <= (layer0_outputs(9175)) and not (layer0_outputs(8186));
    layer1_outputs(8086) <= not((layer0_outputs(7736)) and (layer0_outputs(1950)));
    layer1_outputs(8087) <= (layer0_outputs(4847)) and (layer0_outputs(8960));
    layer1_outputs(8088) <= not((layer0_outputs(3815)) xor (layer0_outputs(15)));
    layer1_outputs(8089) <= layer0_outputs(5540);
    layer1_outputs(8090) <= not((layer0_outputs(714)) or (layer0_outputs(5305)));
    layer1_outputs(8091) <= not((layer0_outputs(9564)) and (layer0_outputs(3938)));
    layer1_outputs(8092) <= not((layer0_outputs(3485)) or (layer0_outputs(9195)));
    layer1_outputs(8093) <= not(layer0_outputs(1157));
    layer1_outputs(8094) <= (layer0_outputs(983)) and not (layer0_outputs(489));
    layer1_outputs(8095) <= not((layer0_outputs(4508)) or (layer0_outputs(4618)));
    layer1_outputs(8096) <= not((layer0_outputs(3814)) or (layer0_outputs(8950)));
    layer1_outputs(8097) <= not(layer0_outputs(1546)) or (layer0_outputs(5489));
    layer1_outputs(8098) <= (layer0_outputs(8891)) and not (layer0_outputs(8396));
    layer1_outputs(8099) <= '0';
    layer1_outputs(8100) <= not(layer0_outputs(5651));
    layer1_outputs(8101) <= not(layer0_outputs(156));
    layer1_outputs(8102) <= layer0_outputs(9364);
    layer1_outputs(8103) <= layer0_outputs(2385);
    layer1_outputs(8104) <= (layer0_outputs(9356)) or (layer0_outputs(8061));
    layer1_outputs(8105) <= (layer0_outputs(9568)) and (layer0_outputs(2085));
    layer1_outputs(8106) <= layer0_outputs(8802);
    layer1_outputs(8107) <= not((layer0_outputs(5045)) or (layer0_outputs(2625)));
    layer1_outputs(8108) <= (layer0_outputs(6357)) and (layer0_outputs(4921));
    layer1_outputs(8109) <= (layer0_outputs(2708)) or (layer0_outputs(4231));
    layer1_outputs(8110) <= not((layer0_outputs(2636)) or (layer0_outputs(8743)));
    layer1_outputs(8111) <= layer0_outputs(7068);
    layer1_outputs(8112) <= not(layer0_outputs(8849));
    layer1_outputs(8113) <= not(layer0_outputs(4607));
    layer1_outputs(8114) <= layer0_outputs(2033);
    layer1_outputs(8115) <= (layer0_outputs(3298)) and (layer0_outputs(8377));
    layer1_outputs(8116) <= not((layer0_outputs(3634)) xor (layer0_outputs(3557)));
    layer1_outputs(8117) <= not(layer0_outputs(5806));
    layer1_outputs(8118) <= layer0_outputs(9831);
    layer1_outputs(8119) <= (layer0_outputs(5875)) and not (layer0_outputs(6790));
    layer1_outputs(8120) <= not(layer0_outputs(3449));
    layer1_outputs(8121) <= '1';
    layer1_outputs(8122) <= layer0_outputs(674);
    layer1_outputs(8123) <= (layer0_outputs(7739)) or (layer0_outputs(886));
    layer1_outputs(8124) <= not((layer0_outputs(3427)) xor (layer0_outputs(8308)));
    layer1_outputs(8125) <= not((layer0_outputs(9753)) and (layer0_outputs(9910)));
    layer1_outputs(8126) <= not((layer0_outputs(3431)) or (layer0_outputs(5543)));
    layer1_outputs(8127) <= (layer0_outputs(7667)) and not (layer0_outputs(156));
    layer1_outputs(8128) <= not((layer0_outputs(1802)) or (layer0_outputs(5496)));
    layer1_outputs(8129) <= not((layer0_outputs(292)) or (layer0_outputs(5425)));
    layer1_outputs(8130) <= not(layer0_outputs(3325)) or (layer0_outputs(3619));
    layer1_outputs(8131) <= not((layer0_outputs(6237)) or (layer0_outputs(2987)));
    layer1_outputs(8132) <= not(layer0_outputs(4827));
    layer1_outputs(8133) <= layer0_outputs(4150);
    layer1_outputs(8134) <= (layer0_outputs(8901)) or (layer0_outputs(8136));
    layer1_outputs(8135) <= (layer0_outputs(3274)) and not (layer0_outputs(555));
    layer1_outputs(8136) <= (layer0_outputs(1869)) and (layer0_outputs(4016));
    layer1_outputs(8137) <= (layer0_outputs(2473)) and not (layer0_outputs(7181));
    layer1_outputs(8138) <= layer0_outputs(3851);
    layer1_outputs(8139) <= not(layer0_outputs(5945));
    layer1_outputs(8140) <= not(layer0_outputs(4019));
    layer1_outputs(8141) <= '1';
    layer1_outputs(8142) <= '1';
    layer1_outputs(8143) <= (layer0_outputs(4814)) and not (layer0_outputs(2606));
    layer1_outputs(8144) <= not((layer0_outputs(4824)) or (layer0_outputs(6441)));
    layer1_outputs(8145) <= (layer0_outputs(6466)) and not (layer0_outputs(4780));
    layer1_outputs(8146) <= not(layer0_outputs(2431)) or (layer0_outputs(7028));
    layer1_outputs(8147) <= (layer0_outputs(634)) and not (layer0_outputs(6080));
    layer1_outputs(8148) <= (layer0_outputs(1856)) and (layer0_outputs(5339));
    layer1_outputs(8149) <= '1';
    layer1_outputs(8150) <= not(layer0_outputs(5721)) or (layer0_outputs(5034));
    layer1_outputs(8151) <= not(layer0_outputs(1620));
    layer1_outputs(8152) <= layer0_outputs(3401);
    layer1_outputs(8153) <= layer0_outputs(6548);
    layer1_outputs(8154) <= (layer0_outputs(8787)) and not (layer0_outputs(1902));
    layer1_outputs(8155) <= (layer0_outputs(8333)) xor (layer0_outputs(6483));
    layer1_outputs(8156) <= '1';
    layer1_outputs(8157) <= not(layer0_outputs(8080));
    layer1_outputs(8158) <= layer0_outputs(5545);
    layer1_outputs(8159) <= layer0_outputs(2451);
    layer1_outputs(8160) <= not((layer0_outputs(973)) and (layer0_outputs(9076)));
    layer1_outputs(8161) <= '0';
    layer1_outputs(8162) <= (layer0_outputs(8770)) and not (layer0_outputs(9239));
    layer1_outputs(8163) <= not(layer0_outputs(1580)) or (layer0_outputs(7955));
    layer1_outputs(8164) <= (layer0_outputs(5360)) and not (layer0_outputs(5653));
    layer1_outputs(8165) <= (layer0_outputs(7803)) and (layer0_outputs(524));
    layer1_outputs(8166) <= (layer0_outputs(3719)) or (layer0_outputs(9871));
    layer1_outputs(8167) <= (layer0_outputs(1099)) and (layer0_outputs(1231));
    layer1_outputs(8168) <= (layer0_outputs(7310)) and not (layer0_outputs(4140));
    layer1_outputs(8169) <= layer0_outputs(8072);
    layer1_outputs(8170) <= not((layer0_outputs(7995)) or (layer0_outputs(8181)));
    layer1_outputs(8171) <= (layer0_outputs(484)) and not (layer0_outputs(4527));
    layer1_outputs(8172) <= (layer0_outputs(3518)) and not (layer0_outputs(9894));
    layer1_outputs(8173) <= not(layer0_outputs(9928));
    layer1_outputs(8174) <= not(layer0_outputs(6627));
    layer1_outputs(8175) <= '0';
    layer1_outputs(8176) <= not((layer0_outputs(1171)) or (layer0_outputs(2256)));
    layer1_outputs(8177) <= not(layer0_outputs(9365));
    layer1_outputs(8178) <= '1';
    layer1_outputs(8179) <= layer0_outputs(312);
    layer1_outputs(8180) <= layer0_outputs(1089);
    layer1_outputs(8181) <= not((layer0_outputs(10217)) and (layer0_outputs(4226)));
    layer1_outputs(8182) <= (layer0_outputs(3809)) and not (layer0_outputs(7429));
    layer1_outputs(8183) <= (layer0_outputs(99)) xor (layer0_outputs(9723));
    layer1_outputs(8184) <= layer0_outputs(434);
    layer1_outputs(8185) <= not((layer0_outputs(8621)) or (layer0_outputs(2306)));
    layer1_outputs(8186) <= (layer0_outputs(9616)) and not (layer0_outputs(8278));
    layer1_outputs(8187) <= not(layer0_outputs(4324));
    layer1_outputs(8188) <= '0';
    layer1_outputs(8189) <= '0';
    layer1_outputs(8190) <= not((layer0_outputs(2347)) and (layer0_outputs(4139)));
    layer1_outputs(8191) <= not(layer0_outputs(6429));
    layer1_outputs(8192) <= not(layer0_outputs(9029)) or (layer0_outputs(4554));
    layer1_outputs(8193) <= not(layer0_outputs(3244));
    layer1_outputs(8194) <= not((layer0_outputs(6084)) xor (layer0_outputs(220)));
    layer1_outputs(8195) <= (layer0_outputs(1559)) or (layer0_outputs(5692));
    layer1_outputs(8196) <= '1';
    layer1_outputs(8197) <= layer0_outputs(2307);
    layer1_outputs(8198) <= not((layer0_outputs(7029)) or (layer0_outputs(1664)));
    layer1_outputs(8199) <= layer0_outputs(4092);
    layer1_outputs(8200) <= not(layer0_outputs(5908));
    layer1_outputs(8201) <= (layer0_outputs(1750)) and not (layer0_outputs(5013));
    layer1_outputs(8202) <= not((layer0_outputs(6490)) or (layer0_outputs(8024)));
    layer1_outputs(8203) <= layer0_outputs(4890);
    layer1_outputs(8204) <= (layer0_outputs(3998)) or (layer0_outputs(6465));
    layer1_outputs(8205) <= (layer0_outputs(10011)) and not (layer0_outputs(6802));
    layer1_outputs(8206) <= not(layer0_outputs(2135)) or (layer0_outputs(1343));
    layer1_outputs(8207) <= not(layer0_outputs(3041));
    layer1_outputs(8208) <= not((layer0_outputs(1905)) xor (layer0_outputs(5742)));
    layer1_outputs(8209) <= not(layer0_outputs(3421)) or (layer0_outputs(8419));
    layer1_outputs(8210) <= not(layer0_outputs(6553)) or (layer0_outputs(4285));
    layer1_outputs(8211) <= (layer0_outputs(2285)) xor (layer0_outputs(8789));
    layer1_outputs(8212) <= (layer0_outputs(311)) or (layer0_outputs(8883));
    layer1_outputs(8213) <= not((layer0_outputs(5827)) or (layer0_outputs(4668)));
    layer1_outputs(8214) <= (layer0_outputs(5803)) and not (layer0_outputs(8165));
    layer1_outputs(8215) <= not(layer0_outputs(6443));
    layer1_outputs(8216) <= layer0_outputs(3568);
    layer1_outputs(8217) <= (layer0_outputs(454)) and not (layer0_outputs(6683));
    layer1_outputs(8218) <= layer0_outputs(7593);
    layer1_outputs(8219) <= layer0_outputs(6149);
    layer1_outputs(8220) <= not((layer0_outputs(287)) or (layer0_outputs(805)));
    layer1_outputs(8221) <= (layer0_outputs(978)) and not (layer0_outputs(5069));
    layer1_outputs(8222) <= '1';
    layer1_outputs(8223) <= layer0_outputs(5358);
    layer1_outputs(8224) <= layer0_outputs(291);
    layer1_outputs(8225) <= not(layer0_outputs(7104));
    layer1_outputs(8226) <= layer0_outputs(6962);
    layer1_outputs(8227) <= '1';
    layer1_outputs(8228) <= not(layer0_outputs(302));
    layer1_outputs(8229) <= not((layer0_outputs(5423)) and (layer0_outputs(1926)));
    layer1_outputs(8230) <= not(layer0_outputs(8083)) or (layer0_outputs(6580));
    layer1_outputs(8231) <= not(layer0_outputs(8183));
    layer1_outputs(8232) <= (layer0_outputs(586)) and not (layer0_outputs(7609));
    layer1_outputs(8233) <= (layer0_outputs(1527)) and not (layer0_outputs(9154));
    layer1_outputs(8234) <= (layer0_outputs(2790)) and not (layer0_outputs(8679));
    layer1_outputs(8235) <= (layer0_outputs(8641)) or (layer0_outputs(9269));
    layer1_outputs(8236) <= (layer0_outputs(5402)) and (layer0_outputs(5888));
    layer1_outputs(8237) <= layer0_outputs(8816);
    layer1_outputs(8238) <= not((layer0_outputs(3064)) or (layer0_outputs(44)));
    layer1_outputs(8239) <= not(layer0_outputs(881)) or (layer0_outputs(2194));
    layer1_outputs(8240) <= (layer0_outputs(1459)) and not (layer0_outputs(4640));
    layer1_outputs(8241) <= (layer0_outputs(7229)) and (layer0_outputs(7981));
    layer1_outputs(8242) <= (layer0_outputs(8508)) and (layer0_outputs(3275));
    layer1_outputs(8243) <= not(layer0_outputs(9880));
    layer1_outputs(8244) <= not((layer0_outputs(7597)) or (layer0_outputs(10170)));
    layer1_outputs(8245) <= not((layer0_outputs(7926)) and (layer0_outputs(4217)));
    layer1_outputs(8246) <= '1';
    layer1_outputs(8247) <= not((layer0_outputs(6353)) and (layer0_outputs(7726)));
    layer1_outputs(8248) <= not(layer0_outputs(619)) or (layer0_outputs(9135));
    layer1_outputs(8249) <= layer0_outputs(3472);
    layer1_outputs(8250) <= not(layer0_outputs(1772));
    layer1_outputs(8251) <= layer0_outputs(2163);
    layer1_outputs(8252) <= layer0_outputs(8821);
    layer1_outputs(8253) <= not(layer0_outputs(7305));
    layer1_outputs(8254) <= (layer0_outputs(887)) and (layer0_outputs(10179));
    layer1_outputs(8255) <= (layer0_outputs(2306)) and not (layer0_outputs(150));
    layer1_outputs(8256) <= (layer0_outputs(5148)) xor (layer0_outputs(575));
    layer1_outputs(8257) <= not(layer0_outputs(4588)) or (layer0_outputs(9431));
    layer1_outputs(8258) <= layer0_outputs(5274);
    layer1_outputs(8259) <= not(layer0_outputs(8350));
    layer1_outputs(8260) <= (layer0_outputs(10026)) and (layer0_outputs(8451));
    layer1_outputs(8261) <= not((layer0_outputs(9670)) xor (layer0_outputs(1261)));
    layer1_outputs(8262) <= layer0_outputs(9004);
    layer1_outputs(8263) <= not((layer0_outputs(4769)) or (layer0_outputs(9110)));
    layer1_outputs(8264) <= layer0_outputs(6838);
    layer1_outputs(8265) <= (layer0_outputs(5534)) or (layer0_outputs(4378));
    layer1_outputs(8266) <= (layer0_outputs(8439)) and not (layer0_outputs(5764));
    layer1_outputs(8267) <= (layer0_outputs(5874)) xor (layer0_outputs(2396));
    layer1_outputs(8268) <= (layer0_outputs(10151)) and not (layer0_outputs(2614));
    layer1_outputs(8269) <= not(layer0_outputs(3202));
    layer1_outputs(8270) <= not((layer0_outputs(841)) and (layer0_outputs(2182)));
    layer1_outputs(8271) <= '1';
    layer1_outputs(8272) <= (layer0_outputs(8311)) and not (layer0_outputs(3995));
    layer1_outputs(8273) <= (layer0_outputs(691)) xor (layer0_outputs(1267));
    layer1_outputs(8274) <= layer0_outputs(5344);
    layer1_outputs(8275) <= not(layer0_outputs(7765)) or (layer0_outputs(7647));
    layer1_outputs(8276) <= (layer0_outputs(8640)) xor (layer0_outputs(3776));
    layer1_outputs(8277) <= (layer0_outputs(1303)) or (layer0_outputs(7663));
    layer1_outputs(8278) <= not(layer0_outputs(2903)) or (layer0_outputs(3643));
    layer1_outputs(8279) <= not(layer0_outputs(6071));
    layer1_outputs(8280) <= not(layer0_outputs(2244)) or (layer0_outputs(5843));
    layer1_outputs(8281) <= not((layer0_outputs(6165)) or (layer0_outputs(9812)));
    layer1_outputs(8282) <= (layer0_outputs(7847)) and not (layer0_outputs(5568));
    layer1_outputs(8283) <= not((layer0_outputs(6079)) or (layer0_outputs(7070)));
    layer1_outputs(8284) <= (layer0_outputs(3948)) and not (layer0_outputs(3782));
    layer1_outputs(8285) <= not(layer0_outputs(9936)) or (layer0_outputs(2904));
    layer1_outputs(8286) <= (layer0_outputs(5589)) and not (layer0_outputs(3056));
    layer1_outputs(8287) <= layer0_outputs(8143);
    layer1_outputs(8288) <= (layer0_outputs(4712)) and not (layer0_outputs(3060));
    layer1_outputs(8289) <= layer0_outputs(2039);
    layer1_outputs(8290) <= not(layer0_outputs(1143));
    layer1_outputs(8291) <= not(layer0_outputs(6821)) or (layer0_outputs(581));
    layer1_outputs(8292) <= '1';
    layer1_outputs(8293) <= (layer0_outputs(2745)) and not (layer0_outputs(8366));
    layer1_outputs(8294) <= not((layer0_outputs(5395)) or (layer0_outputs(4561)));
    layer1_outputs(8295) <= not((layer0_outputs(6777)) or (layer0_outputs(4100)));
    layer1_outputs(8296) <= layer0_outputs(422);
    layer1_outputs(8297) <= layer0_outputs(8074);
    layer1_outputs(8298) <= (layer0_outputs(7613)) and not (layer0_outputs(7542));
    layer1_outputs(8299) <= (layer0_outputs(437)) or (layer0_outputs(7864));
    layer1_outputs(8300) <= not((layer0_outputs(8300)) and (layer0_outputs(8972)));
    layer1_outputs(8301) <= layer0_outputs(337);
    layer1_outputs(8302) <= '0';
    layer1_outputs(8303) <= not(layer0_outputs(8676));
    layer1_outputs(8304) <= (layer0_outputs(593)) and not (layer0_outputs(3426));
    layer1_outputs(8305) <= not(layer0_outputs(9892));
    layer1_outputs(8306) <= layer0_outputs(7639);
    layer1_outputs(8307) <= not(layer0_outputs(8176));
    layer1_outputs(8308) <= (layer0_outputs(7369)) and not (layer0_outputs(8317));
    layer1_outputs(8309) <= (layer0_outputs(2204)) and not (layer0_outputs(4890));
    layer1_outputs(8310) <= not((layer0_outputs(5321)) or (layer0_outputs(8165)));
    layer1_outputs(8311) <= not(layer0_outputs(8579)) or (layer0_outputs(7535));
    layer1_outputs(8312) <= not(layer0_outputs(7595)) or (layer0_outputs(9274));
    layer1_outputs(8313) <= (layer0_outputs(774)) xor (layer0_outputs(4476));
    layer1_outputs(8314) <= (layer0_outputs(5422)) and not (layer0_outputs(2967));
    layer1_outputs(8315) <= (layer0_outputs(2062)) or (layer0_outputs(1716));
    layer1_outputs(8316) <= (layer0_outputs(5181)) or (layer0_outputs(2484));
    layer1_outputs(8317) <= not(layer0_outputs(718));
    layer1_outputs(8318) <= not(layer0_outputs(3501)) or (layer0_outputs(9138));
    layer1_outputs(8319) <= not((layer0_outputs(9244)) or (layer0_outputs(472)));
    layer1_outputs(8320) <= (layer0_outputs(6768)) and (layer0_outputs(307));
    layer1_outputs(8321) <= (layer0_outputs(8241)) and not (layer0_outputs(9329));
    layer1_outputs(8322) <= '1';
    layer1_outputs(8323) <= (layer0_outputs(4782)) or (layer0_outputs(7319));
    layer1_outputs(8324) <= layer0_outputs(7394);
    layer1_outputs(8325) <= not(layer0_outputs(1785)) or (layer0_outputs(1137));
    layer1_outputs(8326) <= not((layer0_outputs(7538)) and (layer0_outputs(10187)));
    layer1_outputs(8327) <= not((layer0_outputs(4550)) or (layer0_outputs(6238)));
    layer1_outputs(8328) <= layer0_outputs(6003);
    layer1_outputs(8329) <= layer0_outputs(2355);
    layer1_outputs(8330) <= (layer0_outputs(5227)) or (layer0_outputs(9028));
    layer1_outputs(8331) <= layer0_outputs(587);
    layer1_outputs(8332) <= not((layer0_outputs(1015)) and (layer0_outputs(1342)));
    layer1_outputs(8333) <= layer0_outputs(7186);
    layer1_outputs(8334) <= (layer0_outputs(4589)) and not (layer0_outputs(2132));
    layer1_outputs(8335) <= (layer0_outputs(2800)) or (layer0_outputs(3987));
    layer1_outputs(8336) <= layer0_outputs(3266);
    layer1_outputs(8337) <= not(layer0_outputs(8240));
    layer1_outputs(8338) <= not((layer0_outputs(5486)) and (layer0_outputs(1687)));
    layer1_outputs(8339) <= not(layer0_outputs(2004));
    layer1_outputs(8340) <= (layer0_outputs(5148)) and (layer0_outputs(3363));
    layer1_outputs(8341) <= (layer0_outputs(9078)) and not (layer0_outputs(9092));
    layer1_outputs(8342) <= not(layer0_outputs(5233)) or (layer0_outputs(6070));
    layer1_outputs(8343) <= not(layer0_outputs(3786)) or (layer0_outputs(198));
    layer1_outputs(8344) <= (layer0_outputs(9018)) and not (layer0_outputs(6417));
    layer1_outputs(8345) <= layer0_outputs(6317);
    layer1_outputs(8346) <= layer0_outputs(7634);
    layer1_outputs(8347) <= not((layer0_outputs(7875)) or (layer0_outputs(8056)));
    layer1_outputs(8348) <= not(layer0_outputs(7148)) or (layer0_outputs(4556));
    layer1_outputs(8349) <= not(layer0_outputs(8234)) or (layer0_outputs(1525));
    layer1_outputs(8350) <= (layer0_outputs(967)) or (layer0_outputs(7258));
    layer1_outputs(8351) <= not((layer0_outputs(385)) or (layer0_outputs(7042)));
    layer1_outputs(8352) <= not((layer0_outputs(4346)) and (layer0_outputs(8668)));
    layer1_outputs(8353) <= '1';
    layer1_outputs(8354) <= layer0_outputs(6922);
    layer1_outputs(8355) <= layer0_outputs(1233);
    layer1_outputs(8356) <= not(layer0_outputs(2861));
    layer1_outputs(8357) <= not(layer0_outputs(6378));
    layer1_outputs(8358) <= layer0_outputs(8794);
    layer1_outputs(8359) <= (layer0_outputs(6188)) and not (layer0_outputs(2654));
    layer1_outputs(8360) <= (layer0_outputs(7390)) and (layer0_outputs(7905));
    layer1_outputs(8361) <= (layer0_outputs(2831)) and not (layer0_outputs(8531));
    layer1_outputs(8362) <= not(layer0_outputs(4448));
    layer1_outputs(8363) <= not(layer0_outputs(2267));
    layer1_outputs(8364) <= not((layer0_outputs(6776)) and (layer0_outputs(8514)));
    layer1_outputs(8365) <= layer0_outputs(2809);
    layer1_outputs(8366) <= not(layer0_outputs(5203)) or (layer0_outputs(3851));
    layer1_outputs(8367) <= (layer0_outputs(8945)) and not (layer0_outputs(9684));
    layer1_outputs(8368) <= (layer0_outputs(9004)) xor (layer0_outputs(2788));
    layer1_outputs(8369) <= layer0_outputs(8951);
    layer1_outputs(8370) <= (layer0_outputs(1319)) and not (layer0_outputs(6276));
    layer1_outputs(8371) <= not(layer0_outputs(5721)) or (layer0_outputs(3068));
    layer1_outputs(8372) <= (layer0_outputs(8332)) or (layer0_outputs(490));
    layer1_outputs(8373) <= not(layer0_outputs(780));
    layer1_outputs(8374) <= layer0_outputs(6043);
    layer1_outputs(8375) <= (layer0_outputs(5190)) or (layer0_outputs(2893));
    layer1_outputs(8376) <= layer0_outputs(7623);
    layer1_outputs(8377) <= layer0_outputs(1133);
    layer1_outputs(8378) <= layer0_outputs(8715);
    layer1_outputs(8379) <= not(layer0_outputs(3368)) or (layer0_outputs(9541));
    layer1_outputs(8380) <= (layer0_outputs(5470)) and not (layer0_outputs(8363));
    layer1_outputs(8381) <= not((layer0_outputs(4466)) or (layer0_outputs(5873)));
    layer1_outputs(8382) <= '1';
    layer1_outputs(8383) <= not((layer0_outputs(6270)) or (layer0_outputs(1399)));
    layer1_outputs(8384) <= (layer0_outputs(5971)) and (layer0_outputs(9035));
    layer1_outputs(8385) <= not(layer0_outputs(5540)) or (layer0_outputs(5022));
    layer1_outputs(8386) <= not((layer0_outputs(3274)) and (layer0_outputs(9712)));
    layer1_outputs(8387) <= layer0_outputs(2494);
    layer1_outputs(8388) <= layer0_outputs(1436);
    layer1_outputs(8389) <= (layer0_outputs(8362)) or (layer0_outputs(4672));
    layer1_outputs(8390) <= layer0_outputs(4566);
    layer1_outputs(8391) <= '1';
    layer1_outputs(8392) <= (layer0_outputs(5471)) and not (layer0_outputs(2353));
    layer1_outputs(8393) <= not(layer0_outputs(9346)) or (layer0_outputs(2653));
    layer1_outputs(8394) <= '1';
    layer1_outputs(8395) <= not((layer0_outputs(4720)) xor (layer0_outputs(5519)));
    layer1_outputs(8396) <= (layer0_outputs(1453)) or (layer0_outputs(10176));
    layer1_outputs(8397) <= (layer0_outputs(5998)) and (layer0_outputs(9708));
    layer1_outputs(8398) <= not(layer0_outputs(4223)) or (layer0_outputs(1286));
    layer1_outputs(8399) <= '1';
    layer1_outputs(8400) <= not(layer0_outputs(8356));
    layer1_outputs(8401) <= not((layer0_outputs(7888)) and (layer0_outputs(5206)));
    layer1_outputs(8402) <= (layer0_outputs(2443)) xor (layer0_outputs(2964));
    layer1_outputs(8403) <= '0';
    layer1_outputs(8404) <= (layer0_outputs(3930)) and not (layer0_outputs(3741));
    layer1_outputs(8405) <= not((layer0_outputs(8446)) xor (layer0_outputs(6758)));
    layer1_outputs(8406) <= not((layer0_outputs(3755)) or (layer0_outputs(7261)));
    layer1_outputs(8407) <= layer0_outputs(35);
    layer1_outputs(8408) <= not(layer0_outputs(4399)) or (layer0_outputs(3732));
    layer1_outputs(8409) <= '1';
    layer1_outputs(8410) <= (layer0_outputs(1007)) and (layer0_outputs(2223));
    layer1_outputs(8411) <= layer0_outputs(2159);
    layer1_outputs(8412) <= (layer0_outputs(1083)) xor (layer0_outputs(7393));
    layer1_outputs(8413) <= layer0_outputs(2805);
    layer1_outputs(8414) <= not((layer0_outputs(293)) or (layer0_outputs(6729)));
    layer1_outputs(8415) <= layer0_outputs(6644);
    layer1_outputs(8416) <= (layer0_outputs(8600)) or (layer0_outputs(5763));
    layer1_outputs(8417) <= (layer0_outputs(4105)) and (layer0_outputs(1532));
    layer1_outputs(8418) <= '0';
    layer1_outputs(8419) <= (layer0_outputs(5227)) and not (layer0_outputs(3547));
    layer1_outputs(8420) <= not(layer0_outputs(6598)) or (layer0_outputs(6950));
    layer1_outputs(8421) <= not(layer0_outputs(7762));
    layer1_outputs(8422) <= (layer0_outputs(9805)) and not (layer0_outputs(3667));
    layer1_outputs(8423) <= not((layer0_outputs(5129)) or (layer0_outputs(4971)));
    layer1_outputs(8424) <= not((layer0_outputs(5434)) or (layer0_outputs(3928)));
    layer1_outputs(8425) <= not(layer0_outputs(4513)) or (layer0_outputs(1067));
    layer1_outputs(8426) <= not((layer0_outputs(7207)) or (layer0_outputs(6655)));
    layer1_outputs(8427) <= '0';
    layer1_outputs(8428) <= not(layer0_outputs(2492));
    layer1_outputs(8429) <= not(layer0_outputs(4491));
    layer1_outputs(8430) <= (layer0_outputs(9647)) and (layer0_outputs(4386));
    layer1_outputs(8431) <= not(layer0_outputs(1994)) or (layer0_outputs(1701));
    layer1_outputs(8432) <= not(layer0_outputs(8342)) or (layer0_outputs(5959));
    layer1_outputs(8433) <= (layer0_outputs(2295)) and (layer0_outputs(12));
    layer1_outputs(8434) <= not(layer0_outputs(8100));
    layer1_outputs(8435) <= not((layer0_outputs(7437)) or (layer0_outputs(6145)));
    layer1_outputs(8436) <= not(layer0_outputs(8111)) or (layer0_outputs(3279));
    layer1_outputs(8437) <= not((layer0_outputs(6603)) and (layer0_outputs(4277)));
    layer1_outputs(8438) <= (layer0_outputs(8509)) or (layer0_outputs(4370));
    layer1_outputs(8439) <= not((layer0_outputs(9993)) and (layer0_outputs(117)));
    layer1_outputs(8440) <= '1';
    layer1_outputs(8441) <= (layer0_outputs(1258)) and not (layer0_outputs(4986));
    layer1_outputs(8442) <= not(layer0_outputs(7179));
    layer1_outputs(8443) <= (layer0_outputs(2006)) xor (layer0_outputs(5098));
    layer1_outputs(8444) <= (layer0_outputs(1104)) xor (layer0_outputs(8335));
    layer1_outputs(8445) <= '1';
    layer1_outputs(8446) <= '1';
    layer1_outputs(8447) <= (layer0_outputs(629)) or (layer0_outputs(2890));
    layer1_outputs(8448) <= '1';
    layer1_outputs(8449) <= '0';
    layer1_outputs(8450) <= '1';
    layer1_outputs(8451) <= not(layer0_outputs(3920)) or (layer0_outputs(1867));
    layer1_outputs(8452) <= (layer0_outputs(777)) and not (layer0_outputs(5731));
    layer1_outputs(8453) <= not((layer0_outputs(9406)) xor (layer0_outputs(917)));
    layer1_outputs(8454) <= (layer0_outputs(7627)) or (layer0_outputs(5539));
    layer1_outputs(8455) <= (layer0_outputs(6936)) and not (layer0_outputs(10239));
    layer1_outputs(8456) <= not(layer0_outputs(8166));
    layer1_outputs(8457) <= (layer0_outputs(9588)) and not (layer0_outputs(4662));
    layer1_outputs(8458) <= not(layer0_outputs(5149));
    layer1_outputs(8459) <= layer0_outputs(6908);
    layer1_outputs(8460) <= not((layer0_outputs(937)) and (layer0_outputs(5947)));
    layer1_outputs(8461) <= not(layer0_outputs(4292)) or (layer0_outputs(121));
    layer1_outputs(8462) <= not(layer0_outputs(4298));
    layer1_outputs(8463) <= '0';
    layer1_outputs(8464) <= (layer0_outputs(4169)) and (layer0_outputs(5613));
    layer1_outputs(8465) <= layer0_outputs(3174);
    layer1_outputs(8466) <= not(layer0_outputs(5740));
    layer1_outputs(8467) <= (layer0_outputs(2485)) and not (layer0_outputs(1509));
    layer1_outputs(8468) <= not(layer0_outputs(8547)) or (layer0_outputs(127));
    layer1_outputs(8469) <= (layer0_outputs(5742)) or (layer0_outputs(129));
    layer1_outputs(8470) <= '0';
    layer1_outputs(8471) <= not((layer0_outputs(2363)) and (layer0_outputs(3290)));
    layer1_outputs(8472) <= layer0_outputs(7867);
    layer1_outputs(8473) <= not((layer0_outputs(2649)) xor (layer0_outputs(2970)));
    layer1_outputs(8474) <= layer0_outputs(6590);
    layer1_outputs(8475) <= (layer0_outputs(2049)) xor (layer0_outputs(3258));
    layer1_outputs(8476) <= (layer0_outputs(400)) and not (layer0_outputs(7218));
    layer1_outputs(8477) <= (layer0_outputs(9100)) xor (layer0_outputs(1903));
    layer1_outputs(8478) <= not(layer0_outputs(9524));
    layer1_outputs(8479) <= layer0_outputs(1267);
    layer1_outputs(8480) <= (layer0_outputs(5936)) and not (layer0_outputs(7341));
    layer1_outputs(8481) <= not((layer0_outputs(1843)) and (layer0_outputs(2467)));
    layer1_outputs(8482) <= (layer0_outputs(1791)) and not (layer0_outputs(6270));
    layer1_outputs(8483) <= not(layer0_outputs(727)) or (layer0_outputs(8397));
    layer1_outputs(8484) <= not(layer0_outputs(8687));
    layer1_outputs(8485) <= not(layer0_outputs(4205));
    layer1_outputs(8486) <= (layer0_outputs(7999)) xor (layer0_outputs(3991));
    layer1_outputs(8487) <= not((layer0_outputs(4033)) xor (layer0_outputs(6781)));
    layer1_outputs(8488) <= not((layer0_outputs(2891)) and (layer0_outputs(6063)));
    layer1_outputs(8489) <= (layer0_outputs(6540)) and (layer0_outputs(5740));
    layer1_outputs(8490) <= (layer0_outputs(9684)) and not (layer0_outputs(9132));
    layer1_outputs(8491) <= (layer0_outputs(6574)) and not (layer0_outputs(4738));
    layer1_outputs(8492) <= not((layer0_outputs(7770)) xor (layer0_outputs(8777)));
    layer1_outputs(8493) <= not((layer0_outputs(4629)) and (layer0_outputs(4842)));
    layer1_outputs(8494) <= not((layer0_outputs(7093)) or (layer0_outputs(9864)));
    layer1_outputs(8495) <= '0';
    layer1_outputs(8496) <= (layer0_outputs(8669)) xor (layer0_outputs(7407));
    layer1_outputs(8497) <= not(layer0_outputs(2687));
    layer1_outputs(8498) <= layer0_outputs(8256);
    layer1_outputs(8499) <= (layer0_outputs(4260)) or (layer0_outputs(6384));
    layer1_outputs(8500) <= not((layer0_outputs(4537)) or (layer0_outputs(3222)));
    layer1_outputs(8501) <= not(layer0_outputs(3284));
    layer1_outputs(8502) <= not(layer0_outputs(9021));
    layer1_outputs(8503) <= not((layer0_outputs(233)) xor (layer0_outputs(3571)));
    layer1_outputs(8504) <= layer0_outputs(7934);
    layer1_outputs(8505) <= not((layer0_outputs(9095)) or (layer0_outputs(9649)));
    layer1_outputs(8506) <= (layer0_outputs(5573)) or (layer0_outputs(7345));
    layer1_outputs(8507) <= (layer0_outputs(4905)) and not (layer0_outputs(2075));
    layer1_outputs(8508) <= not(layer0_outputs(7901));
    layer1_outputs(8509) <= not(layer0_outputs(1435)) or (layer0_outputs(5119));
    layer1_outputs(8510) <= not((layer0_outputs(8344)) or (layer0_outputs(8239)));
    layer1_outputs(8511) <= not((layer0_outputs(1801)) or (layer0_outputs(5709)));
    layer1_outputs(8512) <= (layer0_outputs(3941)) and (layer0_outputs(4181));
    layer1_outputs(8513) <= (layer0_outputs(2909)) or (layer0_outputs(7944));
    layer1_outputs(8514) <= not(layer0_outputs(1104));
    layer1_outputs(8515) <= not(layer0_outputs(9668));
    layer1_outputs(8516) <= layer0_outputs(8759);
    layer1_outputs(8517) <= not(layer0_outputs(2736)) or (layer0_outputs(9417));
    layer1_outputs(8518) <= not(layer0_outputs(7278));
    layer1_outputs(8519) <= '1';
    layer1_outputs(8520) <= not(layer0_outputs(4911));
    layer1_outputs(8521) <= not(layer0_outputs(4989)) or (layer0_outputs(6878));
    layer1_outputs(8522) <= (layer0_outputs(3649)) xor (layer0_outputs(5888));
    layer1_outputs(8523) <= (layer0_outputs(614)) or (layer0_outputs(1454));
    layer1_outputs(8524) <= not(layer0_outputs(1209));
    layer1_outputs(8525) <= not((layer0_outputs(9050)) or (layer0_outputs(10216)));
    layer1_outputs(8526) <= (layer0_outputs(2667)) or (layer0_outputs(1825));
    layer1_outputs(8527) <= (layer0_outputs(3030)) xor (layer0_outputs(1917));
    layer1_outputs(8528) <= not(layer0_outputs(8965));
    layer1_outputs(8529) <= (layer0_outputs(8367)) and (layer0_outputs(2733));
    layer1_outputs(8530) <= not(layer0_outputs(803));
    layer1_outputs(8531) <= layer0_outputs(5320);
    layer1_outputs(8532) <= not((layer0_outputs(8425)) xor (layer0_outputs(10009)));
    layer1_outputs(8533) <= layer0_outputs(4818);
    layer1_outputs(8534) <= not((layer0_outputs(7177)) or (layer0_outputs(2570)));
    layer1_outputs(8535) <= not(layer0_outputs(9438)) or (layer0_outputs(4269));
    layer1_outputs(8536) <= (layer0_outputs(1230)) and not (layer0_outputs(2529));
    layer1_outputs(8537) <= not(layer0_outputs(8757));
    layer1_outputs(8538) <= '0';
    layer1_outputs(8539) <= not(layer0_outputs(6110));
    layer1_outputs(8540) <= '0';
    layer1_outputs(8541) <= not(layer0_outputs(1954)) or (layer0_outputs(9933));
    layer1_outputs(8542) <= not(layer0_outputs(2161));
    layer1_outputs(8543) <= layer0_outputs(5419);
    layer1_outputs(8544) <= not(layer0_outputs(9045));
    layer1_outputs(8545) <= layer0_outputs(7763);
    layer1_outputs(8546) <= (layer0_outputs(1098)) and not (layer0_outputs(808));
    layer1_outputs(8547) <= not(layer0_outputs(7020));
    layer1_outputs(8548) <= not(layer0_outputs(2200));
    layer1_outputs(8549) <= not((layer0_outputs(6385)) and (layer0_outputs(5277)));
    layer1_outputs(8550) <= not(layer0_outputs(7308)) or (layer0_outputs(2165));
    layer1_outputs(8551) <= (layer0_outputs(1133)) and not (layer0_outputs(4002));
    layer1_outputs(8552) <= (layer0_outputs(9197)) and not (layer0_outputs(5455));
    layer1_outputs(8553) <= '0';
    layer1_outputs(8554) <= not((layer0_outputs(2312)) xor (layer0_outputs(9973)));
    layer1_outputs(8555) <= '1';
    layer1_outputs(8556) <= layer0_outputs(3572);
    layer1_outputs(8557) <= not((layer0_outputs(7001)) or (layer0_outputs(2791)));
    layer1_outputs(8558) <= (layer0_outputs(9582)) and not (layer0_outputs(10182));
    layer1_outputs(8559) <= not(layer0_outputs(346));
    layer1_outputs(8560) <= (layer0_outputs(9085)) and not (layer0_outputs(384));
    layer1_outputs(8561) <= not(layer0_outputs(8691));
    layer1_outputs(8562) <= not(layer0_outputs(3482)) or (layer0_outputs(5370));
    layer1_outputs(8563) <= (layer0_outputs(7649)) and not (layer0_outputs(6643));
    layer1_outputs(8564) <= not(layer0_outputs(6875));
    layer1_outputs(8565) <= not((layer0_outputs(3505)) and (layer0_outputs(362)));
    layer1_outputs(8566) <= layer0_outputs(4579);
    layer1_outputs(8567) <= layer0_outputs(5700);
    layer1_outputs(8568) <= not(layer0_outputs(8244));
    layer1_outputs(8569) <= not(layer0_outputs(3207)) or (layer0_outputs(5708));
    layer1_outputs(8570) <= not(layer0_outputs(4825)) or (layer0_outputs(8864));
    layer1_outputs(8571) <= (layer0_outputs(3552)) xor (layer0_outputs(5215));
    layer1_outputs(8572) <= (layer0_outputs(7408)) xor (layer0_outputs(7002));
    layer1_outputs(8573) <= (layer0_outputs(5967)) and not (layer0_outputs(8851));
    layer1_outputs(8574) <= '1';
    layer1_outputs(8575) <= not(layer0_outputs(2190));
    layer1_outputs(8576) <= not(layer0_outputs(7920));
    layer1_outputs(8577) <= not(layer0_outputs(1681));
    layer1_outputs(8578) <= (layer0_outputs(1557)) or (layer0_outputs(2766));
    layer1_outputs(8579) <= (layer0_outputs(7683)) and not (layer0_outputs(8026));
    layer1_outputs(8580) <= not((layer0_outputs(4833)) and (layer0_outputs(8046)));
    layer1_outputs(8581) <= (layer0_outputs(3791)) xor (layer0_outputs(8144));
    layer1_outputs(8582) <= not(layer0_outputs(1611)) or (layer0_outputs(4957));
    layer1_outputs(8583) <= not(layer0_outputs(6902)) or (layer0_outputs(3680));
    layer1_outputs(8584) <= (layer0_outputs(6952)) and not (layer0_outputs(4375));
    layer1_outputs(8585) <= not((layer0_outputs(1097)) and (layer0_outputs(5968)));
    layer1_outputs(8586) <= not((layer0_outputs(5818)) or (layer0_outputs(7348)));
    layer1_outputs(8587) <= not((layer0_outputs(2960)) xor (layer0_outputs(87)));
    layer1_outputs(8588) <= (layer0_outputs(2634)) xor (layer0_outputs(6294));
    layer1_outputs(8589) <= not(layer0_outputs(2804)) or (layer0_outputs(7455));
    layer1_outputs(8590) <= (layer0_outputs(218)) and not (layer0_outputs(7059));
    layer1_outputs(8591) <= not((layer0_outputs(7673)) and (layer0_outputs(9475)));
    layer1_outputs(8592) <= '0';
    layer1_outputs(8593) <= not((layer0_outputs(4990)) or (layer0_outputs(395)));
    layer1_outputs(8594) <= (layer0_outputs(8675)) xor (layer0_outputs(9291));
    layer1_outputs(8595) <= (layer0_outputs(562)) or (layer0_outputs(6167));
    layer1_outputs(8596) <= layer0_outputs(5341);
    layer1_outputs(8597) <= not(layer0_outputs(7857)) or (layer0_outputs(1247));
    layer1_outputs(8598) <= (layer0_outputs(8543)) xor (layer0_outputs(6689));
    layer1_outputs(8599) <= (layer0_outputs(6355)) xor (layer0_outputs(4902));
    layer1_outputs(8600) <= (layer0_outputs(9666)) and not (layer0_outputs(7755));
    layer1_outputs(8601) <= not(layer0_outputs(7324));
    layer1_outputs(8602) <= not(layer0_outputs(4580));
    layer1_outputs(8603) <= (layer0_outputs(7159)) and (layer0_outputs(6889));
    layer1_outputs(8604) <= not((layer0_outputs(3753)) or (layer0_outputs(5393)));
    layer1_outputs(8605) <= (layer0_outputs(733)) or (layer0_outputs(9972));
    layer1_outputs(8606) <= (layer0_outputs(8607)) and (layer0_outputs(128));
    layer1_outputs(8607) <= layer0_outputs(6358);
    layer1_outputs(8608) <= not(layer0_outputs(3262)) or (layer0_outputs(5309));
    layer1_outputs(8609) <= not((layer0_outputs(3260)) or (layer0_outputs(9965)));
    layer1_outputs(8610) <= not(layer0_outputs(8937));
    layer1_outputs(8611) <= (layer0_outputs(596)) and not (layer0_outputs(1665));
    layer1_outputs(8612) <= layer0_outputs(3433);
    layer1_outputs(8613) <= '0';
    layer1_outputs(8614) <= layer0_outputs(9733);
    layer1_outputs(8615) <= (layer0_outputs(9048)) and not (layer0_outputs(3582));
    layer1_outputs(8616) <= not((layer0_outputs(518)) or (layer0_outputs(7325)));
    layer1_outputs(8617) <= (layer0_outputs(545)) and (layer0_outputs(4530));
    layer1_outputs(8618) <= '0';
    layer1_outputs(8619) <= (layer0_outputs(2909)) and (layer0_outputs(2460));
    layer1_outputs(8620) <= (layer0_outputs(6505)) and (layer0_outputs(4526));
    layer1_outputs(8621) <= (layer0_outputs(7232)) and not (layer0_outputs(4075));
    layer1_outputs(8622) <= '1';
    layer1_outputs(8623) <= not((layer0_outputs(652)) or (layer0_outputs(4933)));
    layer1_outputs(8624) <= not(layer0_outputs(2512)) or (layer0_outputs(8158));
    layer1_outputs(8625) <= (layer0_outputs(3175)) and not (layer0_outputs(4110));
    layer1_outputs(8626) <= not((layer0_outputs(3811)) or (layer0_outputs(797)));
    layer1_outputs(8627) <= not(layer0_outputs(8388));
    layer1_outputs(8628) <= not(layer0_outputs(3467)) or (layer0_outputs(9584));
    layer1_outputs(8629) <= layer0_outputs(7183);
    layer1_outputs(8630) <= (layer0_outputs(722)) and (layer0_outputs(9441));
    layer1_outputs(8631) <= not((layer0_outputs(4148)) xor (layer0_outputs(6381)));
    layer1_outputs(8632) <= (layer0_outputs(2142)) and (layer0_outputs(1880));
    layer1_outputs(8633) <= layer0_outputs(8929);
    layer1_outputs(8634) <= (layer0_outputs(9597)) and not (layer0_outputs(1139));
    layer1_outputs(8635) <= not(layer0_outputs(1524));
    layer1_outputs(8636) <= '1';
    layer1_outputs(8637) <= not(layer0_outputs(8974));
    layer1_outputs(8638) <= not(layer0_outputs(2485));
    layer1_outputs(8639) <= '0';
    layer1_outputs(8640) <= not(layer0_outputs(1706)) or (layer0_outputs(10221));
    layer1_outputs(8641) <= (layer0_outputs(6552)) xor (layer0_outputs(7659));
    layer1_outputs(8642) <= (layer0_outputs(1356)) and not (layer0_outputs(2505));
    layer1_outputs(8643) <= not((layer0_outputs(1897)) xor (layer0_outputs(9621)));
    layer1_outputs(8644) <= '0';
    layer1_outputs(8645) <= (layer0_outputs(6392)) and (layer0_outputs(3090));
    layer1_outputs(8646) <= '0';
    layer1_outputs(8647) <= layer0_outputs(7648);
    layer1_outputs(8648) <= (layer0_outputs(8030)) or (layer0_outputs(9180));
    layer1_outputs(8649) <= (layer0_outputs(9088)) and not (layer0_outputs(10230));
    layer1_outputs(8650) <= layer0_outputs(9578);
    layer1_outputs(8651) <= not((layer0_outputs(2566)) or (layer0_outputs(5081)));
    layer1_outputs(8652) <= (layer0_outputs(2905)) or (layer0_outputs(9512));
    layer1_outputs(8653) <= (layer0_outputs(5930)) and not (layer0_outputs(9814));
    layer1_outputs(8654) <= (layer0_outputs(1073)) and not (layer0_outputs(9161));
    layer1_outputs(8655) <= layer0_outputs(335);
    layer1_outputs(8656) <= '0';
    layer1_outputs(8657) <= (layer0_outputs(3039)) and (layer0_outputs(8080));
    layer1_outputs(8658) <= (layer0_outputs(4419)) xor (layer0_outputs(8646));
    layer1_outputs(8659) <= (layer0_outputs(8478)) and not (layer0_outputs(4877));
    layer1_outputs(8660) <= layer0_outputs(8429);
    layer1_outputs(8661) <= not((layer0_outputs(2088)) and (layer0_outputs(7235)));
    layer1_outputs(8662) <= not(layer0_outputs(3718)) or (layer0_outputs(7652));
    layer1_outputs(8663) <= (layer0_outputs(9494)) and not (layer0_outputs(6585));
    layer1_outputs(8664) <= (layer0_outputs(3764)) and (layer0_outputs(5784));
    layer1_outputs(8665) <= not((layer0_outputs(6496)) and (layer0_outputs(5572)));
    layer1_outputs(8666) <= not(layer0_outputs(5748));
    layer1_outputs(8667) <= '1';
    layer1_outputs(8668) <= (layer0_outputs(8329)) and not (layer0_outputs(8753));
    layer1_outputs(8669) <= not(layer0_outputs(2504)) or (layer0_outputs(233));
    layer1_outputs(8670) <= '1';
    layer1_outputs(8671) <= (layer0_outputs(8438)) or (layer0_outputs(6819));
    layer1_outputs(8672) <= not(layer0_outputs(9460)) or (layer0_outputs(6490));
    layer1_outputs(8673) <= not(layer0_outputs(737));
    layer1_outputs(8674) <= not(layer0_outputs(10148)) or (layer0_outputs(7327));
    layer1_outputs(8675) <= layer0_outputs(8599);
    layer1_outputs(8676) <= (layer0_outputs(9887)) and (layer0_outputs(4325));
    layer1_outputs(8677) <= not(layer0_outputs(374)) or (layer0_outputs(4910));
    layer1_outputs(8678) <= not(layer0_outputs(590)) or (layer0_outputs(8321));
    layer1_outputs(8679) <= not(layer0_outputs(366));
    layer1_outputs(8680) <= (layer0_outputs(229)) and not (layer0_outputs(5614));
    layer1_outputs(8681) <= not(layer0_outputs(6419)) or (layer0_outputs(2514));
    layer1_outputs(8682) <= layer0_outputs(9157);
    layer1_outputs(8683) <= not((layer0_outputs(6155)) or (layer0_outputs(5087)));
    layer1_outputs(8684) <= not(layer0_outputs(9974));
    layer1_outputs(8685) <= not((layer0_outputs(882)) xor (layer0_outputs(1622)));
    layer1_outputs(8686) <= layer0_outputs(103);
    layer1_outputs(8687) <= not((layer0_outputs(10007)) xor (layer0_outputs(5260)));
    layer1_outputs(8688) <= not(layer0_outputs(1144));
    layer1_outputs(8689) <= (layer0_outputs(222)) and not (layer0_outputs(3088));
    layer1_outputs(8690) <= not((layer0_outputs(1624)) or (layer0_outputs(3091)));
    layer1_outputs(8691) <= not(layer0_outputs(9026)) or (layer0_outputs(25));
    layer1_outputs(8692) <= not(layer0_outputs(7416));
    layer1_outputs(8693) <= not((layer0_outputs(4534)) or (layer0_outputs(941)));
    layer1_outputs(8694) <= (layer0_outputs(6221)) and (layer0_outputs(3353));
    layer1_outputs(8695) <= not(layer0_outputs(1985));
    layer1_outputs(8696) <= not(layer0_outputs(359));
    layer1_outputs(8697) <= (layer0_outputs(7486)) and not (layer0_outputs(9143));
    layer1_outputs(8698) <= (layer0_outputs(4827)) xor (layer0_outputs(4111));
    layer1_outputs(8699) <= (layer0_outputs(3664)) or (layer0_outputs(7420));
    layer1_outputs(8700) <= not((layer0_outputs(1794)) xor (layer0_outputs(4133)));
    layer1_outputs(8701) <= not(layer0_outputs(5140)) or (layer0_outputs(7563));
    layer1_outputs(8702) <= layer0_outputs(6098);
    layer1_outputs(8703) <= not(layer0_outputs(3152)) or (layer0_outputs(6635));
    layer1_outputs(8704) <= not(layer0_outputs(132));
    layer1_outputs(8705) <= not(layer0_outputs(1984));
    layer1_outputs(8706) <= not(layer0_outputs(5501)) or (layer0_outputs(9646));
    layer1_outputs(8707) <= not(layer0_outputs(5726)) or (layer0_outputs(1901));
    layer1_outputs(8708) <= not(layer0_outputs(2869));
    layer1_outputs(8709) <= not(layer0_outputs(7957)) or (layer0_outputs(7497));
    layer1_outputs(8710) <= layer0_outputs(3021);
    layer1_outputs(8711) <= (layer0_outputs(8656)) or (layer0_outputs(3350));
    layer1_outputs(8712) <= (layer0_outputs(345)) and not (layer0_outputs(9639));
    layer1_outputs(8713) <= not(layer0_outputs(1458)) or (layer0_outputs(213));
    layer1_outputs(8714) <= (layer0_outputs(2552)) and (layer0_outputs(9721));
    layer1_outputs(8715) <= not(layer0_outputs(8472));
    layer1_outputs(8716) <= not(layer0_outputs(5978)) or (layer0_outputs(4793));
    layer1_outputs(8717) <= '1';
    layer1_outputs(8718) <= not(layer0_outputs(2665));
    layer1_outputs(8719) <= not((layer0_outputs(2019)) or (layer0_outputs(1172)));
    layer1_outputs(8720) <= layer0_outputs(8013);
    layer1_outputs(8721) <= (layer0_outputs(6731)) xor (layer0_outputs(8950));
    layer1_outputs(8722) <= not(layer0_outputs(1856)) or (layer0_outputs(1032));
    layer1_outputs(8723) <= not(layer0_outputs(6374)) or (layer0_outputs(1334));
    layer1_outputs(8724) <= layer0_outputs(7182);
    layer1_outputs(8725) <= (layer0_outputs(6509)) xor (layer0_outputs(1755));
    layer1_outputs(8726) <= '1';
    layer1_outputs(8727) <= not(layer0_outputs(8498));
    layer1_outputs(8728) <= (layer0_outputs(1586)) and not (layer0_outputs(3867));
    layer1_outputs(8729) <= not((layer0_outputs(787)) xor (layer0_outputs(5932)));
    layer1_outputs(8730) <= not(layer0_outputs(341));
    layer1_outputs(8731) <= not((layer0_outputs(5838)) xor (layer0_outputs(6536)));
    layer1_outputs(8732) <= (layer0_outputs(352)) xor (layer0_outputs(72));
    layer1_outputs(8733) <= layer0_outputs(5783);
    layer1_outputs(8734) <= '1';
    layer1_outputs(8735) <= not((layer0_outputs(5762)) and (layer0_outputs(8854)));
    layer1_outputs(8736) <= layer0_outputs(8944);
    layer1_outputs(8737) <= '1';
    layer1_outputs(8738) <= (layer0_outputs(9533)) xor (layer0_outputs(3065));
    layer1_outputs(8739) <= not(layer0_outputs(254)) or (layer0_outputs(3299));
    layer1_outputs(8740) <= layer0_outputs(3046);
    layer1_outputs(8741) <= (layer0_outputs(4838)) and not (layer0_outputs(961));
    layer1_outputs(8742) <= not(layer0_outputs(1958)) or (layer0_outputs(9115));
    layer1_outputs(8743) <= (layer0_outputs(4065)) and not (layer0_outputs(653));
    layer1_outputs(8744) <= layer0_outputs(4261);
    layer1_outputs(8745) <= not((layer0_outputs(6226)) and (layer0_outputs(10237)));
    layer1_outputs(8746) <= (layer0_outputs(7203)) and not (layer0_outputs(9238));
    layer1_outputs(8747) <= not((layer0_outputs(4999)) and (layer0_outputs(1472)));
    layer1_outputs(8748) <= '0';
    layer1_outputs(8749) <= not(layer0_outputs(8273));
    layer1_outputs(8750) <= (layer0_outputs(3596)) and not (layer0_outputs(6066));
    layer1_outputs(8751) <= (layer0_outputs(3754)) or (layer0_outputs(1130));
    layer1_outputs(8752) <= (layer0_outputs(9884)) and not (layer0_outputs(716));
    layer1_outputs(8753) <= layer0_outputs(1955);
    layer1_outputs(8754) <= '1';
    layer1_outputs(8755) <= not((layer0_outputs(6838)) or (layer0_outputs(9336)));
    layer1_outputs(8756) <= not(layer0_outputs(10042));
    layer1_outputs(8757) <= layer0_outputs(8528);
    layer1_outputs(8758) <= layer0_outputs(5618);
    layer1_outputs(8759) <= not((layer0_outputs(8195)) and (layer0_outputs(9694)));
    layer1_outputs(8760) <= not(layer0_outputs(1835)) or (layer0_outputs(6601));
    layer1_outputs(8761) <= (layer0_outputs(8680)) and not (layer0_outputs(4165));
    layer1_outputs(8762) <= not(layer0_outputs(129));
    layer1_outputs(8763) <= not((layer0_outputs(5803)) and (layer0_outputs(771)));
    layer1_outputs(8764) <= (layer0_outputs(5929)) and not (layer0_outputs(8724));
    layer1_outputs(8765) <= not((layer0_outputs(1658)) xor (layer0_outputs(4676)));
    layer1_outputs(8766) <= '1';
    layer1_outputs(8767) <= not((layer0_outputs(7046)) or (layer0_outputs(9664)));
    layer1_outputs(8768) <= (layer0_outputs(5748)) xor (layer0_outputs(2591));
    layer1_outputs(8769) <= (layer0_outputs(817)) and not (layer0_outputs(9352));
    layer1_outputs(8770) <= layer0_outputs(9385);
    layer1_outputs(8771) <= (layer0_outputs(844)) and not (layer0_outputs(7927));
    layer1_outputs(8772) <= not(layer0_outputs(2041));
    layer1_outputs(8773) <= '0';
    layer1_outputs(8774) <= layer0_outputs(6266);
    layer1_outputs(8775) <= not((layer0_outputs(8456)) or (layer0_outputs(8387)));
    layer1_outputs(8776) <= not((layer0_outputs(8421)) or (layer0_outputs(1283)));
    layer1_outputs(8777) <= (layer0_outputs(9548)) xor (layer0_outputs(9153));
    layer1_outputs(8778) <= (layer0_outputs(6671)) and not (layer0_outputs(1420));
    layer1_outputs(8779) <= not(layer0_outputs(9188));
    layer1_outputs(8780) <= not(layer0_outputs(2782));
    layer1_outputs(8781) <= (layer0_outputs(346)) xor (layer0_outputs(8231));
    layer1_outputs(8782) <= not((layer0_outputs(5936)) or (layer0_outputs(10222)));
    layer1_outputs(8783) <= not(layer0_outputs(6995));
    layer1_outputs(8784) <= not((layer0_outputs(355)) xor (layer0_outputs(1841)));
    layer1_outputs(8785) <= not(layer0_outputs(5374)) or (layer0_outputs(6741));
    layer1_outputs(8786) <= not(layer0_outputs(7208));
    layer1_outputs(8787) <= not(layer0_outputs(3394)) or (layer0_outputs(4300));
    layer1_outputs(8788) <= layer0_outputs(601);
    layer1_outputs(8789) <= layer0_outputs(1491);
    layer1_outputs(8790) <= (layer0_outputs(6265)) and not (layer0_outputs(4340));
    layer1_outputs(8791) <= not(layer0_outputs(6463));
    layer1_outputs(8792) <= (layer0_outputs(4703)) and not (layer0_outputs(1952));
    layer1_outputs(8793) <= not((layer0_outputs(6839)) xor (layer0_outputs(2366)));
    layer1_outputs(8794) <= layer0_outputs(3430);
    layer1_outputs(8795) <= not(layer0_outputs(4595));
    layer1_outputs(8796) <= not(layer0_outputs(4206));
    layer1_outputs(8797) <= (layer0_outputs(10111)) or (layer0_outputs(145));
    layer1_outputs(8798) <= not(layer0_outputs(7823));
    layer1_outputs(8799) <= not(layer0_outputs(7192));
    layer1_outputs(8800) <= not((layer0_outputs(8067)) and (layer0_outputs(2771)));
    layer1_outputs(8801) <= (layer0_outputs(7338)) and not (layer0_outputs(551));
    layer1_outputs(8802) <= not(layer0_outputs(3682));
    layer1_outputs(8803) <= (layer0_outputs(7783)) or (layer0_outputs(8678));
    layer1_outputs(8804) <= not((layer0_outputs(5856)) or (layer0_outputs(4202)));
    layer1_outputs(8805) <= (layer0_outputs(2723)) and not (layer0_outputs(7775));
    layer1_outputs(8806) <= not(layer0_outputs(3614)) or (layer0_outputs(4166));
    layer1_outputs(8807) <= '1';
    layer1_outputs(8808) <= layer0_outputs(9122);
    layer1_outputs(8809) <= not(layer0_outputs(9535)) or (layer0_outputs(7049));
    layer1_outputs(8810) <= not(layer0_outputs(9462)) or (layer0_outputs(989));
    layer1_outputs(8811) <= not(layer0_outputs(1757));
    layer1_outputs(8812) <= layer0_outputs(184);
    layer1_outputs(8813) <= layer0_outputs(8517);
    layer1_outputs(8814) <= (layer0_outputs(8498)) and not (layer0_outputs(2361));
    layer1_outputs(8815) <= (layer0_outputs(97)) or (layer0_outputs(4186));
    layer1_outputs(8816) <= '1';
    layer1_outputs(8817) <= (layer0_outputs(1005)) and not (layer0_outputs(3514));
    layer1_outputs(8818) <= not(layer0_outputs(8190)) or (layer0_outputs(1170));
    layer1_outputs(8819) <= '0';
    layer1_outputs(8820) <= not(layer0_outputs(7571));
    layer1_outputs(8821) <= (layer0_outputs(9459)) and not (layer0_outputs(7712));
    layer1_outputs(8822) <= (layer0_outputs(7756)) and not (layer0_outputs(6304));
    layer1_outputs(8823) <= layer0_outputs(142);
    layer1_outputs(8824) <= layer0_outputs(10168);
    layer1_outputs(8825) <= not((layer0_outputs(8310)) or (layer0_outputs(6332)));
    layer1_outputs(8826) <= '1';
    layer1_outputs(8827) <= not(layer0_outputs(1953));
    layer1_outputs(8828) <= not((layer0_outputs(3997)) or (layer0_outputs(1819)));
    layer1_outputs(8829) <= not(layer0_outputs(1609));
    layer1_outputs(8830) <= (layer0_outputs(2025)) xor (layer0_outputs(3800));
    layer1_outputs(8831) <= layer0_outputs(9126);
    layer1_outputs(8832) <= not(layer0_outputs(8712)) or (layer0_outputs(6604));
    layer1_outputs(8833) <= layer0_outputs(442);
    layer1_outputs(8834) <= not((layer0_outputs(9222)) or (layer0_outputs(6237)));
    layer1_outputs(8835) <= not((layer0_outputs(5472)) or (layer0_outputs(4071)));
    layer1_outputs(8836) <= layer0_outputs(1822);
    layer1_outputs(8837) <= (layer0_outputs(3907)) and (layer0_outputs(2286));
    layer1_outputs(8838) <= not(layer0_outputs(9089)) or (layer0_outputs(5647));
    layer1_outputs(8839) <= '1';
    layer1_outputs(8840) <= not((layer0_outputs(4425)) or (layer0_outputs(4768)));
    layer1_outputs(8841) <= layer0_outputs(6812);
    layer1_outputs(8842) <= not(layer0_outputs(2584));
    layer1_outputs(8843) <= '0';
    layer1_outputs(8844) <= not(layer0_outputs(620));
    layer1_outputs(8845) <= layer0_outputs(990);
    layer1_outputs(8846) <= (layer0_outputs(9394)) or (layer0_outputs(6058));
    layer1_outputs(8847) <= (layer0_outputs(8209)) and not (layer0_outputs(530));
    layer1_outputs(8848) <= (layer0_outputs(1398)) and (layer0_outputs(8745));
    layer1_outputs(8849) <= (layer0_outputs(757)) xor (layer0_outputs(8889));
    layer1_outputs(8850) <= not(layer0_outputs(9499)) or (layer0_outputs(10157));
    layer1_outputs(8851) <= not((layer0_outputs(8101)) and (layer0_outputs(8614)));
    layer1_outputs(8852) <= (layer0_outputs(8984)) and not (layer0_outputs(486));
    layer1_outputs(8853) <= not((layer0_outputs(2147)) and (layer0_outputs(3889)));
    layer1_outputs(8854) <= layer0_outputs(5450);
    layer1_outputs(8855) <= layer0_outputs(1463);
    layer1_outputs(8856) <= not(layer0_outputs(5464));
    layer1_outputs(8857) <= layer0_outputs(4114);
    layer1_outputs(8858) <= (layer0_outputs(10083)) and not (layer0_outputs(4712));
    layer1_outputs(8859) <= layer0_outputs(5009);
    layer1_outputs(8860) <= (layer0_outputs(3380)) and (layer0_outputs(8449));
    layer1_outputs(8861) <= layer0_outputs(8173);
    layer1_outputs(8862) <= '0';
    layer1_outputs(8863) <= (layer0_outputs(7467)) xor (layer0_outputs(10046));
    layer1_outputs(8864) <= not(layer0_outputs(3363)) or (layer0_outputs(635));
    layer1_outputs(8865) <= (layer0_outputs(8077)) xor (layer0_outputs(4830));
    layer1_outputs(8866) <= not(layer0_outputs(5621));
    layer1_outputs(8867) <= not(layer0_outputs(7440)) or (layer0_outputs(7866));
    layer1_outputs(8868) <= layer0_outputs(7050);
    layer1_outputs(8869) <= not(layer0_outputs(5876)) or (layer0_outputs(3863));
    layer1_outputs(8870) <= layer0_outputs(852);
    layer1_outputs(8871) <= (layer0_outputs(4110)) and not (layer0_outputs(7992));
    layer1_outputs(8872) <= '1';
    layer1_outputs(8873) <= layer0_outputs(3392);
    layer1_outputs(8874) <= not(layer0_outputs(5951));
    layer1_outputs(8875) <= (layer0_outputs(4543)) and not (layer0_outputs(3611));
    layer1_outputs(8876) <= '1';
    layer1_outputs(8877) <= not(layer0_outputs(7032)) or (layer0_outputs(7672));
    layer1_outputs(8878) <= layer0_outputs(8707);
    layer1_outputs(8879) <= '1';
    layer1_outputs(8880) <= (layer0_outputs(529)) xor (layer0_outputs(10013));
    layer1_outputs(8881) <= '0';
    layer1_outputs(8882) <= not((layer0_outputs(3694)) or (layer0_outputs(2974)));
    layer1_outputs(8883) <= not((layer0_outputs(9760)) or (layer0_outputs(2103)));
    layer1_outputs(8884) <= '0';
    layer1_outputs(8885) <= (layer0_outputs(3501)) or (layer0_outputs(8262));
    layer1_outputs(8886) <= layer0_outputs(4396);
    layer1_outputs(8887) <= (layer0_outputs(1065)) and (layer0_outputs(3424));
    layer1_outputs(8888) <= not((layer0_outputs(2113)) xor (layer0_outputs(5240)));
    layer1_outputs(8889) <= not(layer0_outputs(7293)) or (layer0_outputs(2693));
    layer1_outputs(8890) <= layer0_outputs(3316);
    layer1_outputs(8891) <= (layer0_outputs(9679)) and not (layer0_outputs(3805));
    layer1_outputs(8892) <= not((layer0_outputs(1876)) or (layer0_outputs(9471)));
    layer1_outputs(8893) <= (layer0_outputs(8733)) or (layer0_outputs(9707));
    layer1_outputs(8894) <= (layer0_outputs(5172)) or (layer0_outputs(6774));
    layer1_outputs(8895) <= not((layer0_outputs(3742)) and (layer0_outputs(2021)));
    layer1_outputs(8896) <= (layer0_outputs(9201)) and (layer0_outputs(507));
    layer1_outputs(8897) <= not((layer0_outputs(2933)) or (layer0_outputs(6587)));
    layer1_outputs(8898) <= not(layer0_outputs(8140));
    layer1_outputs(8899) <= (layer0_outputs(9971)) xor (layer0_outputs(240));
    layer1_outputs(8900) <= not(layer0_outputs(3172)) or (layer0_outputs(5299));
    layer1_outputs(8901) <= layer0_outputs(10133);
    layer1_outputs(8902) <= not(layer0_outputs(1191));
    layer1_outputs(8903) <= layer0_outputs(6785);
    layer1_outputs(8904) <= (layer0_outputs(3013)) and not (layer0_outputs(6616));
    layer1_outputs(8905) <= not(layer0_outputs(5722)) or (layer0_outputs(1761));
    layer1_outputs(8906) <= layer0_outputs(2991);
    layer1_outputs(8907) <= layer0_outputs(7446);
    layer1_outputs(8908) <= (layer0_outputs(8250)) xor (layer0_outputs(8471));
    layer1_outputs(8909) <= not((layer0_outputs(9856)) and (layer0_outputs(4357)));
    layer1_outputs(8910) <= layer0_outputs(5000);
    layer1_outputs(8911) <= (layer0_outputs(1925)) and not (layer0_outputs(1676));
    layer1_outputs(8912) <= '1';
    layer1_outputs(8913) <= (layer0_outputs(3357)) and not (layer0_outputs(8228));
    layer1_outputs(8914) <= layer0_outputs(8919);
    layer1_outputs(8915) <= not((layer0_outputs(358)) or (layer0_outputs(9419)));
    layer1_outputs(8916) <= layer0_outputs(2066);
    layer1_outputs(8917) <= layer0_outputs(879);
    layer1_outputs(8918) <= not(layer0_outputs(6420)) or (layer0_outputs(6403));
    layer1_outputs(8919) <= '0';
    layer1_outputs(8920) <= not(layer0_outputs(392));
    layer1_outputs(8921) <= (layer0_outputs(4397)) and (layer0_outputs(179));
    layer1_outputs(8922) <= (layer0_outputs(394)) and (layer0_outputs(102));
    layer1_outputs(8923) <= not((layer0_outputs(4157)) or (layer0_outputs(3996)));
    layer1_outputs(8924) <= (layer0_outputs(1843)) and not (layer0_outputs(4376));
    layer1_outputs(8925) <= (layer0_outputs(4246)) and not (layer0_outputs(1829));
    layer1_outputs(8926) <= layer0_outputs(9251);
    layer1_outputs(8927) <= (layer0_outputs(1243)) and not (layer0_outputs(3264));
    layer1_outputs(8928) <= not(layer0_outputs(3083));
    layer1_outputs(8929) <= not(layer0_outputs(628));
    layer1_outputs(8930) <= not(layer0_outputs(6121));
    layer1_outputs(8931) <= not(layer0_outputs(9220));
    layer1_outputs(8932) <= not(layer0_outputs(2431));
    layer1_outputs(8933) <= not(layer0_outputs(5609)) or (layer0_outputs(4897));
    layer1_outputs(8934) <= (layer0_outputs(3736)) and (layer0_outputs(2352));
    layer1_outputs(8935) <= not((layer0_outputs(6893)) or (layer0_outputs(732)));
    layer1_outputs(8936) <= (layer0_outputs(4227)) and not (layer0_outputs(5404));
    layer1_outputs(8937) <= not((layer0_outputs(9559)) xor (layer0_outputs(2750)));
    layer1_outputs(8938) <= (layer0_outputs(2001)) xor (layer0_outputs(9750));
    layer1_outputs(8939) <= not(layer0_outputs(5578));
    layer1_outputs(8940) <= not((layer0_outputs(7670)) and (layer0_outputs(3954)));
    layer1_outputs(8941) <= not(layer0_outputs(7196)) or (layer0_outputs(5145));
    layer1_outputs(8942) <= (layer0_outputs(3176)) or (layer0_outputs(3337));
    layer1_outputs(8943) <= not(layer0_outputs(5782)) or (layer0_outputs(3130));
    layer1_outputs(8944) <= (layer0_outputs(8217)) or (layer0_outputs(5802));
    layer1_outputs(8945) <= not(layer0_outputs(257));
    layer1_outputs(8946) <= not((layer0_outputs(8654)) and (layer0_outputs(7127)));
    layer1_outputs(8947) <= (layer0_outputs(3899)) and not (layer0_outputs(4082));
    layer1_outputs(8948) <= (layer0_outputs(2593)) or (layer0_outputs(811));
    layer1_outputs(8949) <= not((layer0_outputs(4626)) or (layer0_outputs(7521)));
    layer1_outputs(8950) <= (layer0_outputs(2053)) and not (layer0_outputs(3837));
    layer1_outputs(8951) <= not(layer0_outputs(3415)) or (layer0_outputs(1354));
    layer1_outputs(8952) <= (layer0_outputs(2228)) and not (layer0_outputs(1162));
    layer1_outputs(8953) <= (layer0_outputs(136)) and not (layer0_outputs(5780));
    layer1_outputs(8954) <= not(layer0_outputs(4731));
    layer1_outputs(8955) <= not((layer0_outputs(3868)) and (layer0_outputs(5624)));
    layer1_outputs(8956) <= not(layer0_outputs(6166));
    layer1_outputs(8957) <= '1';
    layer1_outputs(8958) <= not(layer0_outputs(6351));
    layer1_outputs(8959) <= not(layer0_outputs(7275));
    layer1_outputs(8960) <= not((layer0_outputs(825)) and (layer0_outputs(1410)));
    layer1_outputs(8961) <= layer0_outputs(2312);
    layer1_outputs(8962) <= not(layer0_outputs(3857));
    layer1_outputs(8963) <= layer0_outputs(4351);
    layer1_outputs(8964) <= (layer0_outputs(8378)) and not (layer0_outputs(7930));
    layer1_outputs(8965) <= not((layer0_outputs(7131)) and (layer0_outputs(5419)));
    layer1_outputs(8966) <= '0';
    layer1_outputs(8967) <= layer0_outputs(9809);
    layer1_outputs(8968) <= layer0_outputs(6927);
    layer1_outputs(8969) <= (layer0_outputs(7758)) and not (layer0_outputs(7649));
    layer1_outputs(8970) <= layer0_outputs(6947);
    layer1_outputs(8971) <= not(layer0_outputs(6471));
    layer1_outputs(8972) <= '0';
    layer1_outputs(8973) <= (layer0_outputs(871)) or (layer0_outputs(6236));
    layer1_outputs(8974) <= '0';
    layer1_outputs(8975) <= not(layer0_outputs(6437));
    layer1_outputs(8976) <= (layer0_outputs(5257)) and not (layer0_outputs(7998));
    layer1_outputs(8977) <= not(layer0_outputs(3451));
    layer1_outputs(8978) <= layer0_outputs(7304);
    layer1_outputs(8979) <= (layer0_outputs(10205)) or (layer0_outputs(9430));
    layer1_outputs(8980) <= not(layer0_outputs(8628));
    layer1_outputs(8981) <= not(layer0_outputs(8180)) or (layer0_outputs(3941));
    layer1_outputs(8982) <= layer0_outputs(1588);
    layer1_outputs(8983) <= not(layer0_outputs(6278));
    layer1_outputs(8984) <= (layer0_outputs(10012)) and not (layer0_outputs(7057));
    layer1_outputs(8985) <= not((layer0_outputs(4197)) or (layer0_outputs(2580)));
    layer1_outputs(8986) <= '1';
    layer1_outputs(8987) <= (layer0_outputs(7367)) and not (layer0_outputs(7184));
    layer1_outputs(8988) <= layer0_outputs(3304);
    layer1_outputs(8989) <= (layer0_outputs(4081)) and not (layer0_outputs(85));
    layer1_outputs(8990) <= not((layer0_outputs(2104)) and (layer0_outputs(8903)));
    layer1_outputs(8991) <= (layer0_outputs(4692)) or (layer0_outputs(8432));
    layer1_outputs(8992) <= not((layer0_outputs(9080)) or (layer0_outputs(2947)));
    layer1_outputs(8993) <= (layer0_outputs(779)) xor (layer0_outputs(2068));
    layer1_outputs(8994) <= not(layer0_outputs(1569));
    layer1_outputs(8995) <= not((layer0_outputs(4992)) and (layer0_outputs(2519)));
    layer1_outputs(8996) <= (layer0_outputs(3111)) xor (layer0_outputs(6926));
    layer1_outputs(8997) <= layer0_outputs(994);
    layer1_outputs(8998) <= (layer0_outputs(818)) and (layer0_outputs(7212));
    layer1_outputs(8999) <= not(layer0_outputs(9532)) or (layer0_outputs(10073));
    layer1_outputs(9000) <= layer0_outputs(2796);
    layer1_outputs(9001) <= (layer0_outputs(5839)) or (layer0_outputs(6559));
    layer1_outputs(9002) <= layer0_outputs(2220);
    layer1_outputs(9003) <= not(layer0_outputs(6162)) or (layer0_outputs(6323));
    layer1_outputs(9004) <= not((layer0_outputs(519)) or (layer0_outputs(6161)));
    layer1_outputs(9005) <= layer0_outputs(5333);
    layer1_outputs(9006) <= not(layer0_outputs(3659)) or (layer0_outputs(5090));
    layer1_outputs(9007) <= not((layer0_outputs(5300)) and (layer0_outputs(6554)));
    layer1_outputs(9008) <= not(layer0_outputs(485));
    layer1_outputs(9009) <= (layer0_outputs(8076)) and not (layer0_outputs(2632));
    layer1_outputs(9010) <= not((layer0_outputs(1727)) and (layer0_outputs(1836)));
    layer1_outputs(9011) <= not((layer0_outputs(3767)) or (layer0_outputs(3624)));
    layer1_outputs(9012) <= (layer0_outputs(7976)) and not (layer0_outputs(565));
    layer1_outputs(9013) <= not(layer0_outputs(966));
    layer1_outputs(9014) <= (layer0_outputs(7106)) and not (layer0_outputs(3769));
    layer1_outputs(9015) <= not(layer0_outputs(2414)) or (layer0_outputs(3205));
    layer1_outputs(9016) <= '0';
    layer1_outputs(9017) <= '0';
    layer1_outputs(9018) <= not(layer0_outputs(9339));
    layer1_outputs(9019) <= not(layer0_outputs(792)) or (layer0_outputs(4129));
    layer1_outputs(9020) <= not((layer0_outputs(232)) or (layer0_outputs(8652)));
    layer1_outputs(9021) <= (layer0_outputs(6288)) and (layer0_outputs(929));
    layer1_outputs(9022) <= not(layer0_outputs(8900));
    layer1_outputs(9023) <= not(layer0_outputs(2056)) or (layer0_outputs(2320));
    layer1_outputs(9024) <= '0';
    layer1_outputs(9025) <= not((layer0_outputs(2472)) xor (layer0_outputs(9409)));
    layer1_outputs(9026) <= not(layer0_outputs(9797));
    layer1_outputs(9027) <= layer0_outputs(8048);
    layer1_outputs(9028) <= layer0_outputs(873);
    layer1_outputs(9029) <= not(layer0_outputs(71));
    layer1_outputs(9030) <= not(layer0_outputs(8625));
    layer1_outputs(9031) <= (layer0_outputs(433)) and not (layer0_outputs(8098));
    layer1_outputs(9032) <= not(layer0_outputs(8278)) or (layer0_outputs(2979));
    layer1_outputs(9033) <= layer0_outputs(6210);
    layer1_outputs(9034) <= not(layer0_outputs(2337)) or (layer0_outputs(3428));
    layer1_outputs(9035) <= not((layer0_outputs(7841)) xor (layer0_outputs(5432)));
    layer1_outputs(9036) <= layer0_outputs(9837);
    layer1_outputs(9037) <= (layer0_outputs(36)) and not (layer0_outputs(412));
    layer1_outputs(9038) <= (layer0_outputs(9192)) and not (layer0_outputs(7855));
    layer1_outputs(9039) <= layer0_outputs(4641);
    layer1_outputs(9040) <= not(layer0_outputs(3404));
    layer1_outputs(9041) <= layer0_outputs(2248);
    layer1_outputs(9042) <= not((layer0_outputs(3735)) and (layer0_outputs(2872)));
    layer1_outputs(9043) <= (layer0_outputs(7842)) and not (layer0_outputs(6647));
    layer1_outputs(9044) <= (layer0_outputs(1120)) or (layer0_outputs(5581));
    layer1_outputs(9045) <= not(layer0_outputs(5884));
    layer1_outputs(9046) <= (layer0_outputs(5993)) and (layer0_outputs(8830));
    layer1_outputs(9047) <= not((layer0_outputs(5759)) and (layer0_outputs(9983)));
    layer1_outputs(9048) <= layer0_outputs(8709);
    layer1_outputs(9049) <= layer0_outputs(393);
    layer1_outputs(9050) <= not(layer0_outputs(8016)) or (layer0_outputs(9299));
    layer1_outputs(9051) <= layer0_outputs(2937);
    layer1_outputs(9052) <= not((layer0_outputs(2432)) and (layer0_outputs(622)));
    layer1_outputs(9053) <= not(layer0_outputs(7333));
    layer1_outputs(9054) <= not(layer0_outputs(2711));
    layer1_outputs(9055) <= not((layer0_outputs(3253)) and (layer0_outputs(9472)));
    layer1_outputs(9056) <= (layer0_outputs(4905)) and not (layer0_outputs(1894));
    layer1_outputs(9057) <= (layer0_outputs(6700)) or (layer0_outputs(3393));
    layer1_outputs(9058) <= not(layer0_outputs(3120)) or (layer0_outputs(6155));
    layer1_outputs(9059) <= (layer0_outputs(8134)) and not (layer0_outputs(8148));
    layer1_outputs(9060) <= not(layer0_outputs(9629));
    layer1_outputs(9061) <= '1';
    layer1_outputs(9062) <= layer0_outputs(8598);
    layer1_outputs(9063) <= (layer0_outputs(9480)) and (layer0_outputs(1146));
    layer1_outputs(9064) <= not(layer0_outputs(7440));
    layer1_outputs(9065) <= not((layer0_outputs(6930)) xor (layer0_outputs(7363)));
    layer1_outputs(9066) <= (layer0_outputs(8326)) xor (layer0_outputs(9464));
    layer1_outputs(9067) <= '0';
    layer1_outputs(9068) <= layer0_outputs(2637);
    layer1_outputs(9069) <= (layer0_outputs(7299)) xor (layer0_outputs(2096));
    layer1_outputs(9070) <= not((layer0_outputs(4298)) or (layer0_outputs(1541)));
    layer1_outputs(9071) <= (layer0_outputs(5872)) and not (layer0_outputs(2024));
    layer1_outputs(9072) <= not(layer0_outputs(8395));
    layer1_outputs(9073) <= not(layer0_outputs(1544));
    layer1_outputs(9074) <= not((layer0_outputs(7506)) or (layer0_outputs(5694)));
    layer1_outputs(9075) <= not((layer0_outputs(1441)) or (layer0_outputs(637)));
    layer1_outputs(9076) <= (layer0_outputs(149)) and not (layer0_outputs(5700));
    layer1_outputs(9077) <= (layer0_outputs(4159)) or (layer0_outputs(3389));
    layer1_outputs(9078) <= not((layer0_outputs(8091)) and (layer0_outputs(809)));
    layer1_outputs(9079) <= (layer0_outputs(8577)) and not (layer0_outputs(5652));
    layer1_outputs(9080) <= (layer0_outputs(2373)) and not (layer0_outputs(7802));
    layer1_outputs(9081) <= not((layer0_outputs(682)) or (layer0_outputs(6633)));
    layer1_outputs(9082) <= (layer0_outputs(4743)) and (layer0_outputs(5067));
    layer1_outputs(9083) <= (layer0_outputs(2826)) and not (layer0_outputs(5224));
    layer1_outputs(9084) <= (layer0_outputs(824)) and (layer0_outputs(6064));
    layer1_outputs(9085) <= not(layer0_outputs(7067));
    layer1_outputs(9086) <= not(layer0_outputs(4040));
    layer1_outputs(9087) <= layer0_outputs(1498);
    layer1_outputs(9088) <= not(layer0_outputs(285)) or (layer0_outputs(7804));
    layer1_outputs(9089) <= not((layer0_outputs(4275)) and (layer0_outputs(1433)));
    layer1_outputs(9090) <= '0';
    layer1_outputs(9091) <= not((layer0_outputs(3204)) or (layer0_outputs(7271)));
    layer1_outputs(9092) <= '0';
    layer1_outputs(9093) <= (layer0_outputs(9755)) or (layer0_outputs(9087));
    layer1_outputs(9094) <= layer0_outputs(3078);
    layer1_outputs(9095) <= not((layer0_outputs(3935)) or (layer0_outputs(5454)));
    layer1_outputs(9096) <= not(layer0_outputs(10144));
    layer1_outputs(9097) <= not((layer0_outputs(10068)) or (layer0_outputs(5819)));
    layer1_outputs(9098) <= (layer0_outputs(6287)) xor (layer0_outputs(5618));
    layer1_outputs(9099) <= not((layer0_outputs(7732)) and (layer0_outputs(4732)));
    layer1_outputs(9100) <= layer0_outputs(925);
    layer1_outputs(9101) <= (layer0_outputs(5773)) or (layer0_outputs(2845));
    layer1_outputs(9102) <= (layer0_outputs(3033)) xor (layer0_outputs(6426));
    layer1_outputs(9103) <= (layer0_outputs(10004)) and not (layer0_outputs(789));
    layer1_outputs(9104) <= '1';
    layer1_outputs(9105) <= (layer0_outputs(4657)) and not (layer0_outputs(4778));
    layer1_outputs(9106) <= not(layer0_outputs(7447)) or (layer0_outputs(7421));
    layer1_outputs(9107) <= (layer0_outputs(219)) or (layer0_outputs(8093));
    layer1_outputs(9108) <= layer0_outputs(3354);
    layer1_outputs(9109) <= not(layer0_outputs(8146)) or (layer0_outputs(190));
    layer1_outputs(9110) <= (layer0_outputs(4478)) xor (layer0_outputs(9987));
    layer1_outputs(9111) <= layer0_outputs(3751);
    layer1_outputs(9112) <= not(layer0_outputs(1126));
    layer1_outputs(9113) <= not(layer0_outputs(7462)) or (layer0_outputs(1044));
    layer1_outputs(9114) <= not(layer0_outputs(4567)) or (layer0_outputs(6488));
    layer1_outputs(9115) <= not(layer0_outputs(1570));
    layer1_outputs(9116) <= (layer0_outputs(31)) and (layer0_outputs(7427));
    layer1_outputs(9117) <= layer0_outputs(10110);
    layer1_outputs(9118) <= not(layer0_outputs(3351));
    layer1_outputs(9119) <= layer0_outputs(9521);
    layer1_outputs(9120) <= not(layer0_outputs(5556));
    layer1_outputs(9121) <= (layer0_outputs(10171)) xor (layer0_outputs(1758));
    layer1_outputs(9122) <= (layer0_outputs(858)) and (layer0_outputs(6075));
    layer1_outputs(9123) <= (layer0_outputs(5012)) and not (layer0_outputs(7519));
    layer1_outputs(9124) <= (layer0_outputs(3645)) xor (layer0_outputs(3961));
    layer1_outputs(9125) <= (layer0_outputs(10098)) and (layer0_outputs(6418));
    layer1_outputs(9126) <= not(layer0_outputs(9370));
    layer1_outputs(9127) <= (layer0_outputs(4361)) and (layer0_outputs(987));
    layer1_outputs(9128) <= not(layer0_outputs(9256));
    layer1_outputs(9129) <= not((layer0_outputs(9668)) and (layer0_outputs(2963)));
    layer1_outputs(9130) <= layer0_outputs(9526);
    layer1_outputs(9131) <= not((layer0_outputs(4468)) and (layer0_outputs(3396)));
    layer1_outputs(9132) <= (layer0_outputs(4578)) and (layer0_outputs(5735));
    layer1_outputs(9133) <= not(layer0_outputs(8468)) or (layer0_outputs(3103));
    layer1_outputs(9134) <= layer0_outputs(4449);
    layer1_outputs(9135) <= '0';
    layer1_outputs(9136) <= (layer0_outputs(5561)) or (layer0_outputs(8194));
    layer1_outputs(9137) <= not((layer0_outputs(489)) and (layer0_outputs(8743)));
    layer1_outputs(9138) <= layer0_outputs(2639);
    layer1_outputs(9139) <= (layer0_outputs(1965)) or (layer0_outputs(2968));
    layer1_outputs(9140) <= layer0_outputs(2360);
    layer1_outputs(9141) <= not(layer0_outputs(8356)) or (layer0_outputs(9451));
    layer1_outputs(9142) <= not(layer0_outputs(4903));
    layer1_outputs(9143) <= not(layer0_outputs(5884));
    layer1_outputs(9144) <= not(layer0_outputs(978)) or (layer0_outputs(178));
    layer1_outputs(9145) <= not(layer0_outputs(9030)) or (layer0_outputs(10059));
    layer1_outputs(9146) <= (layer0_outputs(4829)) and (layer0_outputs(998));
    layer1_outputs(9147) <= (layer0_outputs(5860)) xor (layer0_outputs(7401));
    layer1_outputs(9148) <= layer0_outputs(809);
    layer1_outputs(9149) <= (layer0_outputs(2351)) and (layer0_outputs(5113));
    layer1_outputs(9150) <= layer0_outputs(6602);
    layer1_outputs(9151) <= not((layer0_outputs(4044)) or (layer0_outputs(9258)));
    layer1_outputs(9152) <= not(layer0_outputs(2757));
    layer1_outputs(9153) <= layer0_outputs(4729);
    layer1_outputs(9154) <= not(layer0_outputs(1566));
    layer1_outputs(9155) <= (layer0_outputs(6873)) or (layer0_outputs(4317));
    layer1_outputs(9156) <= not(layer0_outputs(6347)) or (layer0_outputs(7438));
    layer1_outputs(9157) <= not(layer0_outputs(9357)) or (layer0_outputs(915));
    layer1_outputs(9158) <= layer0_outputs(2941);
    layer1_outputs(9159) <= not(layer0_outputs(8116)) or (layer0_outputs(3497));
    layer1_outputs(9160) <= not(layer0_outputs(5497)) or (layer0_outputs(5709));
    layer1_outputs(9161) <= not(layer0_outputs(754));
    layer1_outputs(9162) <= not(layer0_outputs(8778)) or (layer0_outputs(7078));
    layer1_outputs(9163) <= layer0_outputs(4082);
    layer1_outputs(9164) <= not((layer0_outputs(5017)) and (layer0_outputs(6445)));
    layer1_outputs(9165) <= layer0_outputs(9529);
    layer1_outputs(9166) <= '0';
    layer1_outputs(9167) <= not(layer0_outputs(8593)) or (layer0_outputs(4184));
    layer1_outputs(9168) <= not((layer0_outputs(6806)) xor (layer0_outputs(9705)));
    layer1_outputs(9169) <= '1';
    layer1_outputs(9170) <= not(layer0_outputs(7108)) or (layer0_outputs(8230));
    layer1_outputs(9171) <= not(layer0_outputs(932)) or (layer0_outputs(5535));
    layer1_outputs(9172) <= not((layer0_outputs(9547)) and (layer0_outputs(9952)));
    layer1_outputs(9173) <= not(layer0_outputs(4131)) or (layer0_outputs(1023));
    layer1_outputs(9174) <= '1';
    layer1_outputs(9175) <= (layer0_outputs(2084)) or (layer0_outputs(8673));
    layer1_outputs(9176) <= '1';
    layer1_outputs(9177) <= not(layer0_outputs(6216)) or (layer0_outputs(7761));
    layer1_outputs(9178) <= layer0_outputs(7400);
    layer1_outputs(9179) <= not((layer0_outputs(902)) xor (layer0_outputs(6720)));
    layer1_outputs(9180) <= (layer0_outputs(527)) or (layer0_outputs(9368));
    layer1_outputs(9181) <= not((layer0_outputs(3487)) or (layer0_outputs(6711)));
    layer1_outputs(9182) <= not((layer0_outputs(1477)) and (layer0_outputs(9891)));
    layer1_outputs(9183) <= not(layer0_outputs(6401)) or (layer0_outputs(1004));
    layer1_outputs(9184) <= not(layer0_outputs(1206)) or (layer0_outputs(9067));
    layer1_outputs(9185) <= (layer0_outputs(3725)) and not (layer0_outputs(4670));
    layer1_outputs(9186) <= (layer0_outputs(7034)) xor (layer0_outputs(2229));
    layer1_outputs(9187) <= layer0_outputs(5792);
    layer1_outputs(9188) <= '1';
    layer1_outputs(9189) <= (layer0_outputs(3311)) xor (layer0_outputs(7713));
    layer1_outputs(9190) <= layer0_outputs(9126);
    layer1_outputs(9191) <= not(layer0_outputs(6826));
    layer1_outputs(9192) <= not(layer0_outputs(8047)) or (layer0_outputs(10037));
    layer1_outputs(9193) <= layer0_outputs(8585);
    layer1_outputs(9194) <= layer0_outputs(7567);
    layer1_outputs(9195) <= not(layer0_outputs(4297));
    layer1_outputs(9196) <= not((layer0_outputs(3526)) or (layer0_outputs(4104)));
    layer1_outputs(9197) <= not((layer0_outputs(7396)) xor (layer0_outputs(1431)));
    layer1_outputs(9198) <= (layer0_outputs(8634)) and not (layer0_outputs(10160));
    layer1_outputs(9199) <= not((layer0_outputs(5876)) or (layer0_outputs(8434)));
    layer1_outputs(9200) <= '1';
    layer1_outputs(9201) <= (layer0_outputs(3046)) xor (layer0_outputs(7859));
    layer1_outputs(9202) <= (layer0_outputs(8957)) or (layer0_outputs(2452));
    layer1_outputs(9203) <= '0';
    layer1_outputs(9204) <= (layer0_outputs(9666)) xor (layer0_outputs(9744));
    layer1_outputs(9205) <= (layer0_outputs(10167)) and (layer0_outputs(6527));
    layer1_outputs(9206) <= layer0_outputs(7194);
    layer1_outputs(9207) <= (layer0_outputs(8379)) and not (layer0_outputs(4368));
    layer1_outputs(9208) <= (layer0_outputs(3231)) and not (layer0_outputs(9950));
    layer1_outputs(9209) <= (layer0_outputs(10189)) and not (layer0_outputs(1333));
    layer1_outputs(9210) <= (layer0_outputs(5852)) xor (layer0_outputs(1490));
    layer1_outputs(9211) <= layer0_outputs(3840);
    layer1_outputs(9212) <= layer0_outputs(1187);
    layer1_outputs(9213) <= not(layer0_outputs(3398));
    layer1_outputs(9214) <= (layer0_outputs(3870)) and (layer0_outputs(7026));
    layer1_outputs(9215) <= layer0_outputs(2302);
    layer1_outputs(9216) <= (layer0_outputs(7381)) and (layer0_outputs(3876));
    layer1_outputs(9217) <= (layer0_outputs(3097)) and not (layer0_outputs(6960));
    layer1_outputs(9218) <= not(layer0_outputs(6431)) or (layer0_outputs(3112));
    layer1_outputs(9219) <= not((layer0_outputs(7264)) and (layer0_outputs(2429)));
    layer1_outputs(9220) <= (layer0_outputs(1690)) and (layer0_outputs(6227));
    layer1_outputs(9221) <= (layer0_outputs(8042)) or (layer0_outputs(9171));
    layer1_outputs(9222) <= not(layer0_outputs(7537));
    layer1_outputs(9223) <= (layer0_outputs(4630)) and (layer0_outputs(6028));
    layer1_outputs(9224) <= (layer0_outputs(6753)) and (layer0_outputs(10170));
    layer1_outputs(9225) <= (layer0_outputs(1642)) and not (layer0_outputs(6804));
    layer1_outputs(9226) <= not((layer0_outputs(3085)) and (layer0_outputs(704)));
    layer1_outputs(9227) <= not((layer0_outputs(9109)) or (layer0_outputs(2896)));
    layer1_outputs(9228) <= not(layer0_outputs(8243));
    layer1_outputs(9229) <= not(layer0_outputs(2617));
    layer1_outputs(9230) <= (layer0_outputs(6793)) and not (layer0_outputs(4746));
    layer1_outputs(9231) <= layer0_outputs(6696);
    layer1_outputs(9232) <= not(layer0_outputs(4335));
    layer1_outputs(9233) <= (layer0_outputs(347)) or (layer0_outputs(4054));
    layer1_outputs(9234) <= (layer0_outputs(4802)) and (layer0_outputs(7387));
    layer1_outputs(9235) <= not(layer0_outputs(6710));
    layer1_outputs(9236) <= layer0_outputs(6178);
    layer1_outputs(9237) <= layer0_outputs(9511);
    layer1_outputs(9238) <= '0';
    layer1_outputs(9239) <= '1';
    layer1_outputs(9240) <= layer0_outputs(837);
    layer1_outputs(9241) <= not(layer0_outputs(7322)) or (layer0_outputs(4281));
    layer1_outputs(9242) <= not((layer0_outputs(55)) or (layer0_outputs(6738)));
    layer1_outputs(9243) <= layer0_outputs(3418);
    layer1_outputs(9244) <= '1';
    layer1_outputs(9245) <= layer0_outputs(699);
    layer1_outputs(9246) <= '0';
    layer1_outputs(9247) <= (layer0_outputs(323)) and not (layer0_outputs(2423));
    layer1_outputs(9248) <= (layer0_outputs(5031)) and (layer0_outputs(7253));
    layer1_outputs(9249) <= not(layer0_outputs(567));
    layer1_outputs(9250) <= '0';
    layer1_outputs(9251) <= not(layer0_outputs(4699));
    layer1_outputs(9252) <= not(layer0_outputs(2137)) or (layer0_outputs(2659));
    layer1_outputs(9253) <= not(layer0_outputs(4405));
    layer1_outputs(9254) <= not(layer0_outputs(1985));
    layer1_outputs(9255) <= not(layer0_outputs(5894)) or (layer0_outputs(6549));
    layer1_outputs(9256) <= not(layer0_outputs(4103));
    layer1_outputs(9257) <= (layer0_outputs(3541)) or (layer0_outputs(6070));
    layer1_outputs(9258) <= layer0_outputs(2170);
    layer1_outputs(9259) <= (layer0_outputs(420)) and not (layer0_outputs(4124));
    layer1_outputs(9260) <= '0';
    layer1_outputs(9261) <= not(layer0_outputs(1291));
    layer1_outputs(9262) <= (layer0_outputs(6479)) and not (layer0_outputs(3588));
    layer1_outputs(9263) <= not((layer0_outputs(3598)) or (layer0_outputs(242)));
    layer1_outputs(9264) <= not(layer0_outputs(3464));
    layer1_outputs(9265) <= '0';
    layer1_outputs(9266) <= (layer0_outputs(5191)) and (layer0_outputs(1678));
    layer1_outputs(9267) <= not(layer0_outputs(2920));
    layer1_outputs(9268) <= not((layer0_outputs(9714)) xor (layer0_outputs(3332)));
    layer1_outputs(9269) <= not((layer0_outputs(2016)) xor (layer0_outputs(2786)));
    layer1_outputs(9270) <= layer0_outputs(9571);
    layer1_outputs(9271) <= not(layer0_outputs(4724));
    layer1_outputs(9272) <= (layer0_outputs(8556)) and (layer0_outputs(3207));
    layer1_outputs(9273) <= not((layer0_outputs(3361)) or (layer0_outputs(6578)));
    layer1_outputs(9274) <= not(layer0_outputs(1529)) or (layer0_outputs(4364));
    layer1_outputs(9275) <= (layer0_outputs(2597)) or (layer0_outputs(7342));
    layer1_outputs(9276) <= layer0_outputs(8266);
    layer1_outputs(9277) <= layer0_outputs(765);
    layer1_outputs(9278) <= not((layer0_outputs(2195)) xor (layer0_outputs(10055)));
    layer1_outputs(9279) <= not((layer0_outputs(1220)) xor (layer0_outputs(5285)));
    layer1_outputs(9280) <= (layer0_outputs(6047)) and (layer0_outputs(5247));
    layer1_outputs(9281) <= (layer0_outputs(2286)) and not (layer0_outputs(8581));
    layer1_outputs(9282) <= layer0_outputs(5200);
    layer1_outputs(9283) <= not((layer0_outputs(7113)) and (layer0_outputs(4888)));
    layer1_outputs(9284) <= not((layer0_outputs(1026)) and (layer0_outputs(9271)));
    layer1_outputs(9285) <= (layer0_outputs(5422)) and not (layer0_outputs(2195));
    layer1_outputs(9286) <= not((layer0_outputs(2531)) xor (layer0_outputs(712)));
    layer1_outputs(9287) <= not(layer0_outputs(4500)) or (layer0_outputs(7863));
    layer1_outputs(9288) <= '1';
    layer1_outputs(9289) <= layer0_outputs(4687);
    layer1_outputs(9290) <= layer0_outputs(7248);
    layer1_outputs(9291) <= layer0_outputs(1082);
    layer1_outputs(9292) <= (layer0_outputs(7294)) or (layer0_outputs(8548));
    layer1_outputs(9293) <= not(layer0_outputs(9544));
    layer1_outputs(9294) <= not(layer0_outputs(1408));
    layer1_outputs(9295) <= (layer0_outputs(5698)) xor (layer0_outputs(6269));
    layer1_outputs(9296) <= (layer0_outputs(9926)) and not (layer0_outputs(7325));
    layer1_outputs(9297) <= (layer0_outputs(4948)) and not (layer0_outputs(3343));
    layer1_outputs(9298) <= (layer0_outputs(5966)) or (layer0_outputs(5334));
    layer1_outputs(9299) <= '1';
    layer1_outputs(9300) <= (layer0_outputs(2150)) and not (layer0_outputs(3499));
    layer1_outputs(9301) <= layer0_outputs(5021);
    layer1_outputs(9302) <= (layer0_outputs(5851)) and not (layer0_outputs(10011));
    layer1_outputs(9303) <= not(layer0_outputs(8878));
    layer1_outputs(9304) <= '0';
    layer1_outputs(9305) <= not(layer0_outputs(640)) or (layer0_outputs(4388));
    layer1_outputs(9306) <= layer0_outputs(6812);
    layer1_outputs(9307) <= layer0_outputs(2146);
    layer1_outputs(9308) <= (layer0_outputs(10063)) and (layer0_outputs(2413));
    layer1_outputs(9309) <= not((layer0_outputs(6179)) xor (layer0_outputs(1384)));
    layer1_outputs(9310) <= (layer0_outputs(2206)) xor (layer0_outputs(1449));
    layer1_outputs(9311) <= not(layer0_outputs(322)) or (layer0_outputs(6894));
    layer1_outputs(9312) <= not((layer0_outputs(6575)) and (layer0_outputs(4419)));
    layer1_outputs(9313) <= (layer0_outputs(4495)) and not (layer0_outputs(2360));
    layer1_outputs(9314) <= '0';
    layer1_outputs(9315) <= not(layer0_outputs(1362));
    layer1_outputs(9316) <= not(layer0_outputs(3094));
    layer1_outputs(9317) <= (layer0_outputs(6482)) and not (layer0_outputs(8044));
    layer1_outputs(9318) <= not(layer0_outputs(5214));
    layer1_outputs(9319) <= not(layer0_outputs(4182));
    layer1_outputs(9320) <= (layer0_outputs(8618)) xor (layer0_outputs(1515));
    layer1_outputs(9321) <= '1';
    layer1_outputs(9322) <= layer0_outputs(6134);
    layer1_outputs(9323) <= not((layer0_outputs(840)) or (layer0_outputs(6555)));
    layer1_outputs(9324) <= (layer0_outputs(3771)) or (layer0_outputs(2254));
    layer1_outputs(9325) <= (layer0_outputs(10019)) or (layer0_outputs(633));
    layer1_outputs(9326) <= (layer0_outputs(6132)) and (layer0_outputs(3931));
    layer1_outputs(9327) <= not(layer0_outputs(3220));
    layer1_outputs(9328) <= not(layer0_outputs(2482));
    layer1_outputs(9329) <= '0';
    layer1_outputs(9330) <= not(layer0_outputs(2549)) or (layer0_outputs(4755));
    layer1_outputs(9331) <= (layer0_outputs(8649)) and (layer0_outputs(4302));
    layer1_outputs(9332) <= not(layer0_outputs(3730)) or (layer0_outputs(8525));
    layer1_outputs(9333) <= not(layer0_outputs(7954)) or (layer0_outputs(2584));
    layer1_outputs(9334) <= not((layer0_outputs(7251)) or (layer0_outputs(5953)));
    layer1_outputs(9335) <= '1';
    layer1_outputs(9336) <= '0';
    layer1_outputs(9337) <= layer0_outputs(5493);
    layer1_outputs(9338) <= (layer0_outputs(7753)) and (layer0_outputs(1302));
    layer1_outputs(9339) <= (layer0_outputs(2692)) and (layer0_outputs(6956));
    layer1_outputs(9340) <= not(layer0_outputs(8570));
    layer1_outputs(9341) <= layer0_outputs(3626);
    layer1_outputs(9342) <= (layer0_outputs(644)) and not (layer0_outputs(7971));
    layer1_outputs(9343) <= not(layer0_outputs(10199)) or (layer0_outputs(2834));
    layer1_outputs(9344) <= (layer0_outputs(6492)) and (layer0_outputs(4819));
    layer1_outputs(9345) <= '1';
    layer1_outputs(9346) <= not((layer0_outputs(8470)) and (layer0_outputs(7213)));
    layer1_outputs(9347) <= not(layer0_outputs(411));
    layer1_outputs(9348) <= not(layer0_outputs(9825)) or (layer0_outputs(3487));
    layer1_outputs(9349) <= (layer0_outputs(3647)) and not (layer0_outputs(4026));
    layer1_outputs(9350) <= (layer0_outputs(6606)) and not (layer0_outputs(2995));
    layer1_outputs(9351) <= not((layer0_outputs(2513)) or (layer0_outputs(169)));
    layer1_outputs(9352) <= not((layer0_outputs(1629)) and (layer0_outputs(8871)));
    layer1_outputs(9353) <= not(layer0_outputs(4757)) or (layer0_outputs(8144));
    layer1_outputs(9354) <= not(layer0_outputs(1255)) or (layer0_outputs(5830));
    layer1_outputs(9355) <= not(layer0_outputs(8479)) or (layer0_outputs(7168));
    layer1_outputs(9356) <= not((layer0_outputs(4485)) and (layer0_outputs(6626)));
    layer1_outputs(9357) <= layer0_outputs(3972);
    layer1_outputs(9358) <= layer0_outputs(4034);
    layer1_outputs(9359) <= not(layer0_outputs(6128));
    layer1_outputs(9360) <= (layer0_outputs(10010)) and not (layer0_outputs(8365));
    layer1_outputs(9361) <= (layer0_outputs(8171)) and not (layer0_outputs(5341));
    layer1_outputs(9362) <= (layer0_outputs(4447)) and (layer0_outputs(6789));
    layer1_outputs(9363) <= (layer0_outputs(6588)) and (layer0_outputs(3816));
    layer1_outputs(9364) <= not(layer0_outputs(7739));
    layer1_outputs(9365) <= (layer0_outputs(1310)) and (layer0_outputs(9716));
    layer1_outputs(9366) <= not(layer0_outputs(2957));
    layer1_outputs(9367) <= layer0_outputs(5848);
    layer1_outputs(9368) <= layer0_outputs(3978);
    layer1_outputs(9369) <= not(layer0_outputs(5796)) or (layer0_outputs(5630));
    layer1_outputs(9370) <= not(layer0_outputs(6739));
    layer1_outputs(9371) <= (layer0_outputs(6561)) and (layer0_outputs(4020));
    layer1_outputs(9372) <= not((layer0_outputs(3187)) xor (layer0_outputs(9469)));
    layer1_outputs(9373) <= not(layer0_outputs(4966)) or (layer0_outputs(6907));
    layer1_outputs(9374) <= layer0_outputs(6975);
    layer1_outputs(9375) <= not(layer0_outputs(377));
    layer1_outputs(9376) <= '1';
    layer1_outputs(9377) <= not((layer0_outputs(3568)) xor (layer0_outputs(3642)));
    layer1_outputs(9378) <= layer0_outputs(612);
    layer1_outputs(9379) <= (layer0_outputs(9345)) xor (layer0_outputs(8559));
    layer1_outputs(9380) <= (layer0_outputs(7174)) xor (layer0_outputs(10001));
    layer1_outputs(9381) <= (layer0_outputs(1080)) and not (layer0_outputs(5282));
    layer1_outputs(9382) <= not((layer0_outputs(993)) or (layer0_outputs(8651)));
    layer1_outputs(9383) <= not(layer0_outputs(10073)) or (layer0_outputs(6589));
    layer1_outputs(9384) <= not(layer0_outputs(7077));
    layer1_outputs(9385) <= layer0_outputs(7058);
    layer1_outputs(9386) <= (layer0_outputs(3370)) or (layer0_outputs(9830));
    layer1_outputs(9387) <= layer0_outputs(8996);
    layer1_outputs(9388) <= not(layer0_outputs(1428)) or (layer0_outputs(8627));
    layer1_outputs(9389) <= layer0_outputs(4420);
    layer1_outputs(9390) <= layer0_outputs(3495);
    layer1_outputs(9391) <= layer0_outputs(9335);
    layer1_outputs(9392) <= (layer0_outputs(4688)) xor (layer0_outputs(677));
    layer1_outputs(9393) <= layer0_outputs(7592);
    layer1_outputs(9394) <= layer0_outputs(2564);
    layer1_outputs(9395) <= (layer0_outputs(7144)) and not (layer0_outputs(1431));
    layer1_outputs(9396) <= '1';
    layer1_outputs(9397) <= (layer0_outputs(8287)) and not (layer0_outputs(5171));
    layer1_outputs(9398) <= not(layer0_outputs(8002));
    layer1_outputs(9399) <= not((layer0_outputs(10080)) and (layer0_outputs(5564)));
    layer1_outputs(9400) <= not(layer0_outputs(7374)) or (layer0_outputs(2553));
    layer1_outputs(9401) <= (layer0_outputs(9593)) and (layer0_outputs(17));
    layer1_outputs(9402) <= (layer0_outputs(8407)) or (layer0_outputs(9075));
    layer1_outputs(9403) <= (layer0_outputs(9089)) xor (layer0_outputs(8753));
    layer1_outputs(9404) <= not(layer0_outputs(1981)) or (layer0_outputs(3623));
    layer1_outputs(9405) <= not(layer0_outputs(8772));
    layer1_outputs(9406) <= not(layer0_outputs(9366));
    layer1_outputs(9407) <= '1';
    layer1_outputs(9408) <= not(layer0_outputs(4045)) or (layer0_outputs(5023));
    layer1_outputs(9409) <= (layer0_outputs(1969)) and not (layer0_outputs(7472));
    layer1_outputs(9410) <= layer0_outputs(8879);
    layer1_outputs(9411) <= layer0_outputs(5605);
    layer1_outputs(9412) <= not(layer0_outputs(5002)) or (layer0_outputs(6319));
    layer1_outputs(9413) <= not((layer0_outputs(6639)) xor (layer0_outputs(4391)));
    layer1_outputs(9414) <= (layer0_outputs(3)) xor (layer0_outputs(1839));
    layer1_outputs(9415) <= layer0_outputs(8963);
    layer1_outputs(9416) <= (layer0_outputs(9865)) and not (layer0_outputs(7759));
    layer1_outputs(9417) <= not((layer0_outputs(9069)) xor (layer0_outputs(9099)));
    layer1_outputs(9418) <= not(layer0_outputs(2304));
    layer1_outputs(9419) <= not(layer0_outputs(4790));
    layer1_outputs(9420) <= (layer0_outputs(6960)) xor (layer0_outputs(10166));
    layer1_outputs(9421) <= '0';
    layer1_outputs(9422) <= not(layer0_outputs(3078)) or (layer0_outputs(2234));
    layer1_outputs(9423) <= layer0_outputs(303);
    layer1_outputs(9424) <= '0';
    layer1_outputs(9425) <= not(layer0_outputs(5421)) or (layer0_outputs(982));
    layer1_outputs(9426) <= not(layer0_outputs(7120)) or (layer0_outputs(5526));
    layer1_outputs(9427) <= (layer0_outputs(4923)) or (layer0_outputs(6832));
    layer1_outputs(9428) <= not((layer0_outputs(4926)) xor (layer0_outputs(4178)));
    layer1_outputs(9429) <= (layer0_outputs(5167)) and not (layer0_outputs(3411));
    layer1_outputs(9430) <= not((layer0_outputs(3609)) and (layer0_outputs(6292)));
    layer1_outputs(9431) <= not(layer0_outputs(9426)) or (layer0_outputs(5828));
    layer1_outputs(9432) <= layer0_outputs(4453);
    layer1_outputs(9433) <= '0';
    layer1_outputs(9434) <= (layer0_outputs(8869)) and not (layer0_outputs(9121));
    layer1_outputs(9435) <= (layer0_outputs(7970)) and not (layer0_outputs(2917));
    layer1_outputs(9436) <= not(layer0_outputs(3492));
    layer1_outputs(9437) <= '0';
    layer1_outputs(9438) <= layer0_outputs(8520);
    layer1_outputs(9439) <= (layer0_outputs(680)) or (layer0_outputs(8094));
    layer1_outputs(9440) <= not((layer0_outputs(6502)) and (layer0_outputs(2041)));
    layer1_outputs(9441) <= layer0_outputs(6464);
    layer1_outputs(9442) <= not(layer0_outputs(7945)) or (layer0_outputs(1248));
    layer1_outputs(9443) <= layer0_outputs(423);
    layer1_outputs(9444) <= not(layer0_outputs(6386)) or (layer0_outputs(1079));
    layer1_outputs(9445) <= not((layer0_outputs(7777)) or (layer0_outputs(930)));
    layer1_outputs(9446) <= not(layer0_outputs(4612)) or (layer0_outputs(4922));
    layer1_outputs(9447) <= layer0_outputs(2720);
    layer1_outputs(9448) <= (layer0_outputs(1009)) and not (layer0_outputs(4521));
    layer1_outputs(9449) <= not(layer0_outputs(7965));
    layer1_outputs(9450) <= not(layer0_outputs(2590));
    layer1_outputs(9451) <= (layer0_outputs(2464)) and (layer0_outputs(6508));
    layer1_outputs(9452) <= (layer0_outputs(6740)) and not (layer0_outputs(713));
    layer1_outputs(9453) <= (layer0_outputs(1863)) or (layer0_outputs(7893));
    layer1_outputs(9454) <= (layer0_outputs(5537)) and (layer0_outputs(9559));
    layer1_outputs(9455) <= (layer0_outputs(3392)) or (layer0_outputs(9327));
    layer1_outputs(9456) <= not((layer0_outputs(971)) and (layer0_outputs(4321)));
    layer1_outputs(9457) <= not(layer0_outputs(7587)) or (layer0_outputs(2988));
    layer1_outputs(9458) <= not(layer0_outputs(2722));
    layer1_outputs(9459) <= layer0_outputs(8601);
    layer1_outputs(9460) <= (layer0_outputs(1301)) or (layer0_outputs(3358));
    layer1_outputs(9461) <= '0';
    layer1_outputs(9462) <= not(layer0_outputs(3252)) or (layer0_outputs(3548));
    layer1_outputs(9463) <= layer0_outputs(3292);
    layer1_outputs(9464) <= (layer0_outputs(10043)) and not (layer0_outputs(2514));
    layer1_outputs(9465) <= (layer0_outputs(3880)) xor (layer0_outputs(5431));
    layer1_outputs(9466) <= layer0_outputs(8366);
    layer1_outputs(9467) <= (layer0_outputs(470)) and not (layer0_outputs(2728));
    layer1_outputs(9468) <= not((layer0_outputs(9681)) and (layer0_outputs(3412)));
    layer1_outputs(9469) <= (layer0_outputs(8361)) and not (layer0_outputs(4066));
    layer1_outputs(9470) <= layer0_outputs(5499);
    layer1_outputs(9471) <= not((layer0_outputs(3832)) or (layer0_outputs(2688)));
    layer1_outputs(9472) <= not(layer0_outputs(8315)) or (layer0_outputs(3939));
    layer1_outputs(9473) <= not(layer0_outputs(3295)) or (layer0_outputs(7514));
    layer1_outputs(9474) <= (layer0_outputs(5942)) and not (layer0_outputs(4980));
    layer1_outputs(9475) <= '1';
    layer1_outputs(9476) <= layer0_outputs(1956);
    layer1_outputs(9477) <= (layer0_outputs(783)) or (layer0_outputs(7460));
    layer1_outputs(9478) <= (layer0_outputs(1125)) xor (layer0_outputs(5030));
    layer1_outputs(9479) <= (layer0_outputs(7364)) and not (layer0_outputs(1236));
    layer1_outputs(9480) <= layer0_outputs(5688);
    layer1_outputs(9481) <= not(layer0_outputs(3341));
    layer1_outputs(9482) <= (layer0_outputs(6307)) and not (layer0_outputs(8995));
    layer1_outputs(9483) <= not(layer0_outputs(4694)) or (layer0_outputs(766));
    layer1_outputs(9484) <= (layer0_outputs(6604)) xor (layer0_outputs(9849));
    layer1_outputs(9485) <= (layer0_outputs(50)) and not (layer0_outputs(1417));
    layer1_outputs(9486) <= layer0_outputs(1358);
    layer1_outputs(9487) <= layer0_outputs(166);
    layer1_outputs(9488) <= '1';
    layer1_outputs(9489) <= '0';
    layer1_outputs(9490) <= (layer0_outputs(6843)) or (layer0_outputs(7118));
    layer1_outputs(9491) <= not((layer0_outputs(6789)) or (layer0_outputs(1539)));
    layer1_outputs(9492) <= not(layer0_outputs(7168));
    layer1_outputs(9493) <= (layer0_outputs(5196)) and (layer0_outputs(5745));
    layer1_outputs(9494) <= (layer0_outputs(8514)) or (layer0_outputs(8389));
    layer1_outputs(9495) <= (layer0_outputs(8968)) and not (layer0_outputs(9861));
    layer1_outputs(9496) <= layer0_outputs(4754);
    layer1_outputs(9497) <= not((layer0_outputs(3154)) xor (layer0_outputs(9105)));
    layer1_outputs(9498) <= '0';
    layer1_outputs(9499) <= layer0_outputs(4620);
    layer1_outputs(9500) <= not(layer0_outputs(776)) or (layer0_outputs(8368));
    layer1_outputs(9501) <= '0';
    layer1_outputs(9502) <= layer0_outputs(8040);
    layer1_outputs(9503) <= layer0_outputs(9416);
    layer1_outputs(9504) <= not(layer0_outputs(9070));
    layer1_outputs(9505) <= not((layer0_outputs(5336)) xor (layer0_outputs(8457)));
    layer1_outputs(9506) <= (layer0_outputs(9112)) or (layer0_outputs(1998));
    layer1_outputs(9507) <= not((layer0_outputs(3012)) xor (layer0_outputs(997)));
    layer1_outputs(9508) <= (layer0_outputs(9224)) and not (layer0_outputs(3383));
    layer1_outputs(9509) <= not(layer0_outputs(2518));
    layer1_outputs(9510) <= not(layer0_outputs(8622));
    layer1_outputs(9511) <= not(layer0_outputs(3878));
    layer1_outputs(9512) <= not(layer0_outputs(8516)) or (layer0_outputs(195));
    layer1_outputs(9513) <= '1';
    layer1_outputs(9514) <= not((layer0_outputs(5147)) or (layer0_outputs(7620)));
    layer1_outputs(9515) <= (layer0_outputs(4674)) and (layer0_outputs(7109));
    layer1_outputs(9516) <= (layer0_outputs(5693)) and not (layer0_outputs(8776));
    layer1_outputs(9517) <= layer0_outputs(1021);
    layer1_outputs(9518) <= layer0_outputs(8916);
    layer1_outputs(9519) <= (layer0_outputs(9692)) xor (layer0_outputs(1898));
    layer1_outputs(9520) <= not((layer0_outputs(2156)) xor (layer0_outputs(747)));
    layer1_outputs(9521) <= not((layer0_outputs(477)) and (layer0_outputs(8583)));
    layer1_outputs(9522) <= not(layer0_outputs(6082)) or (layer0_outputs(7081));
    layer1_outputs(9523) <= layer0_outputs(4414);
    layer1_outputs(9524) <= layer0_outputs(5323);
    layer1_outputs(9525) <= (layer0_outputs(2486)) xor (layer0_outputs(1762));
    layer1_outputs(9526) <= (layer0_outputs(8549)) xor (layer0_outputs(6630));
    layer1_outputs(9527) <= layer0_outputs(1513);
    layer1_outputs(9528) <= not((layer0_outputs(1167)) or (layer0_outputs(1737)));
    layer1_outputs(9529) <= not((layer0_outputs(9127)) xor (layer0_outputs(4643)));
    layer1_outputs(9530) <= (layer0_outputs(6813)) or (layer0_outputs(4224));
    layer1_outputs(9531) <= not(layer0_outputs(1388));
    layer1_outputs(9532) <= layer0_outputs(5472);
    layer1_outputs(9533) <= not(layer0_outputs(8401)) or (layer0_outputs(2262));
    layer1_outputs(9534) <= not((layer0_outputs(4635)) or (layer0_outputs(2175)));
    layer1_outputs(9535) <= (layer0_outputs(9242)) and (layer0_outputs(7711));
    layer1_outputs(9536) <= (layer0_outputs(3062)) and (layer0_outputs(7831));
    layer1_outputs(9537) <= not(layer0_outputs(6906));
    layer1_outputs(9538) <= (layer0_outputs(10041)) xor (layer0_outputs(3224));
    layer1_outputs(9539) <= not(layer0_outputs(8877));
    layer1_outputs(9540) <= '0';
    layer1_outputs(9541) <= (layer0_outputs(8816)) and not (layer0_outputs(2503));
    layer1_outputs(9542) <= layer0_outputs(7719);
    layer1_outputs(9543) <= (layer0_outputs(6546)) and not (layer0_outputs(3149));
    layer1_outputs(9544) <= (layer0_outputs(2226)) and not (layer0_outputs(6360));
    layer1_outputs(9545) <= (layer0_outputs(4555)) or (layer0_outputs(2269));
    layer1_outputs(9546) <= not(layer0_outputs(4286)) or (layer0_outputs(10016));
    layer1_outputs(9547) <= layer0_outputs(4387);
    layer1_outputs(9548) <= (layer0_outputs(23)) xor (layer0_outputs(4906));
    layer1_outputs(9549) <= layer0_outputs(8506);
    layer1_outputs(9550) <= layer0_outputs(6140);
    layer1_outputs(9551) <= not(layer0_outputs(861)) or (layer0_outputs(6102));
    layer1_outputs(9552) <= not(layer0_outputs(959));
    layer1_outputs(9553) <= (layer0_outputs(4185)) and (layer0_outputs(435));
    layer1_outputs(9554) <= layer0_outputs(3093);
    layer1_outputs(9555) <= not((layer0_outputs(2143)) and (layer0_outputs(1717)));
    layer1_outputs(9556) <= not(layer0_outputs(6967));
    layer1_outputs(9557) <= layer0_outputs(2821);
    layer1_outputs(9558) <= layer0_outputs(5051);
    layer1_outputs(9559) <= (layer0_outputs(10076)) or (layer0_outputs(6553));
    layer1_outputs(9560) <= layer0_outputs(1041);
    layer1_outputs(9561) <= '1';
    layer1_outputs(9562) <= not(layer0_outputs(5170)) or (layer0_outputs(7585));
    layer1_outputs(9563) <= (layer0_outputs(1600)) xor (layer0_outputs(543));
    layer1_outputs(9564) <= layer0_outputs(9763);
    layer1_outputs(9565) <= not((layer0_outputs(7653)) or (layer0_outputs(621)));
    layer1_outputs(9566) <= (layer0_outputs(9648)) and not (layer0_outputs(7679));
    layer1_outputs(9567) <= not(layer0_outputs(1150));
    layer1_outputs(9568) <= (layer0_outputs(7494)) and not (layer0_outputs(2389));
    layer1_outputs(9569) <= not(layer0_outputs(9983));
    layer1_outputs(9570) <= not(layer0_outputs(7970));
    layer1_outputs(9571) <= not((layer0_outputs(561)) or (layer0_outputs(8636)));
    layer1_outputs(9572) <= (layer0_outputs(6722)) or (layer0_outputs(10084));
    layer1_outputs(9573) <= not(layer0_outputs(5121));
    layer1_outputs(9574) <= (layer0_outputs(6617)) and not (layer0_outputs(6040));
    layer1_outputs(9575) <= not((layer0_outputs(7128)) or (layer0_outputs(3226)));
    layer1_outputs(9576) <= not(layer0_outputs(3070));
    layer1_outputs(9577) <= not((layer0_outputs(3597)) or (layer0_outputs(2109)));
    layer1_outputs(9578) <= layer0_outputs(6025);
    layer1_outputs(9579) <= not(layer0_outputs(9413));
    layer1_outputs(9580) <= (layer0_outputs(8877)) and not (layer0_outputs(9570));
    layer1_outputs(9581) <= not(layer0_outputs(7578));
    layer1_outputs(9582) <= not((layer0_outputs(7786)) and (layer0_outputs(9981)));
    layer1_outputs(9583) <= (layer0_outputs(9858)) and not (layer0_outputs(6456));
    layer1_outputs(9584) <= not(layer0_outputs(4656));
    layer1_outputs(9585) <= not(layer0_outputs(3480)) or (layer0_outputs(8859));
    layer1_outputs(9586) <= layer0_outputs(7485);
    layer1_outputs(9587) <= not(layer0_outputs(1580));
    layer1_outputs(9588) <= not(layer0_outputs(9090));
    layer1_outputs(9589) <= not((layer0_outputs(4373)) or (layer0_outputs(8714)));
    layer1_outputs(9590) <= '1';
    layer1_outputs(9591) <= '0';
    layer1_outputs(9592) <= layer0_outputs(6972);
    layer1_outputs(9593) <= (layer0_outputs(1455)) and not (layer0_outputs(5142));
    layer1_outputs(9594) <= layer0_outputs(1814);
    layer1_outputs(9595) <= (layer0_outputs(10013)) and not (layer0_outputs(5647));
    layer1_outputs(9596) <= (layer0_outputs(1797)) or (layer0_outputs(2403));
    layer1_outputs(9597) <= (layer0_outputs(3477)) or (layer0_outputs(5086));
    layer1_outputs(9598) <= not(layer0_outputs(8474)) or (layer0_outputs(1148));
    layer1_outputs(9599) <= not(layer0_outputs(4895)) or (layer0_outputs(9997));
    layer1_outputs(9600) <= not(layer0_outputs(5444));
    layer1_outputs(9601) <= (layer0_outputs(5974)) and not (layer0_outputs(1458));
    layer1_outputs(9602) <= not(layer0_outputs(350));
    layer1_outputs(9603) <= (layer0_outputs(2578)) and (layer0_outputs(3444));
    layer1_outputs(9604) <= layer0_outputs(6100);
    layer1_outputs(9605) <= not((layer0_outputs(5955)) and (layer0_outputs(4863)));
    layer1_outputs(9606) <= layer0_outputs(73);
    layer1_outputs(9607) <= '1';
    layer1_outputs(9608) <= not(layer0_outputs(6548)) or (layer0_outputs(4519));
    layer1_outputs(9609) <= not((layer0_outputs(1644)) and (layer0_outputs(8835)));
    layer1_outputs(9610) <= layer0_outputs(3598);
    layer1_outputs(9611) <= not(layer0_outputs(8486));
    layer1_outputs(9612) <= (layer0_outputs(9678)) and (layer0_outputs(9893));
    layer1_outputs(9613) <= (layer0_outputs(8423)) and not (layer0_outputs(6666));
    layer1_outputs(9614) <= not((layer0_outputs(9255)) and (layer0_outputs(5330)));
    layer1_outputs(9615) <= (layer0_outputs(5024)) xor (layer0_outputs(5084));
    layer1_outputs(9616) <= not((layer0_outputs(6150)) or (layer0_outputs(1418)));
    layer1_outputs(9617) <= not(layer0_outputs(6087));
    layer1_outputs(9618) <= (layer0_outputs(3747)) xor (layer0_outputs(202));
    layer1_outputs(9619) <= (layer0_outputs(8284)) and not (layer0_outputs(7963));
    layer1_outputs(9620) <= (layer0_outputs(6219)) and not (layer0_outputs(5365));
    layer1_outputs(9621) <= layer0_outputs(8285);
    layer1_outputs(9622) <= (layer0_outputs(5089)) and not (layer0_outputs(3257));
    layer1_outputs(9623) <= (layer0_outputs(5295)) and not (layer0_outputs(10074));
    layer1_outputs(9624) <= not(layer0_outputs(2010));
    layer1_outputs(9625) <= not(layer0_outputs(8990)) or (layer0_outputs(3550));
    layer1_outputs(9626) <= '1';
    layer1_outputs(9627) <= (layer0_outputs(4483)) and (layer0_outputs(80));
    layer1_outputs(9628) <= '1';
    layer1_outputs(9629) <= layer0_outputs(13);
    layer1_outputs(9630) <= not(layer0_outputs(1535));
    layer1_outputs(9631) <= (layer0_outputs(7296)) or (layer0_outputs(5772));
    layer1_outputs(9632) <= (layer0_outputs(3012)) and not (layer0_outputs(7086));
    layer1_outputs(9633) <= not(layer0_outputs(1625)) or (layer0_outputs(4406));
    layer1_outputs(9634) <= (layer0_outputs(5793)) and not (layer0_outputs(7896));
    layer1_outputs(9635) <= not(layer0_outputs(3344));
    layer1_outputs(9636) <= (layer0_outputs(994)) or (layer0_outputs(4595));
    layer1_outputs(9637) <= (layer0_outputs(3578)) and not (layer0_outputs(6285));
    layer1_outputs(9638) <= (layer0_outputs(803)) or (layer0_outputs(81));
    layer1_outputs(9639) <= not((layer0_outputs(1192)) and (layer0_outputs(7699)));
    layer1_outputs(9640) <= not(layer0_outputs(1604)) or (layer0_outputs(1959));
    layer1_outputs(9641) <= layer0_outputs(472);
    layer1_outputs(9642) <= layer0_outputs(9439);
    layer1_outputs(9643) <= (layer0_outputs(7064)) or (layer0_outputs(6338));
    layer1_outputs(9644) <= layer0_outputs(8058);
    layer1_outputs(9645) <= not(layer0_outputs(509));
    layer1_outputs(9646) <= layer0_outputs(6762);
    layer1_outputs(9647) <= not(layer0_outputs(4395)) or (layer0_outputs(606));
    layer1_outputs(9648) <= not((layer0_outputs(2797)) and (layer0_outputs(3866)));
    layer1_outputs(9649) <= (layer0_outputs(5481)) and not (layer0_outputs(7741));
    layer1_outputs(9650) <= not((layer0_outputs(9550)) or (layer0_outputs(5857)));
    layer1_outputs(9651) <= (layer0_outputs(6497)) or (layer0_outputs(9489));
    layer1_outputs(9652) <= (layer0_outputs(4614)) and (layer0_outputs(1338));
    layer1_outputs(9653) <= (layer0_outputs(1834)) xor (layer0_outputs(2421));
    layer1_outputs(9654) <= layer0_outputs(5390);
    layer1_outputs(9655) <= not(layer0_outputs(7449));
    layer1_outputs(9656) <= layer0_outputs(7831);
    layer1_outputs(9657) <= not(layer0_outputs(5764));
    layer1_outputs(9658) <= not(layer0_outputs(1109));
    layer1_outputs(9659) <= layer0_outputs(2258);
    layer1_outputs(9660) <= layer0_outputs(9434);
    layer1_outputs(9661) <= not(layer0_outputs(7445));
    layer1_outputs(9662) <= layer0_outputs(6312);
    layer1_outputs(9663) <= not((layer0_outputs(2558)) or (layer0_outputs(8806)));
    layer1_outputs(9664) <= layer0_outputs(1484);
    layer1_outputs(9665) <= not((layer0_outputs(7330)) and (layer0_outputs(9478)));
    layer1_outputs(9666) <= not((layer0_outputs(7300)) and (layer0_outputs(104)));
    layer1_outputs(9667) <= not(layer0_outputs(5999));
    layer1_outputs(9668) <= (layer0_outputs(10165)) and not (layer0_outputs(137));
    layer1_outputs(9669) <= not(layer0_outputs(5871));
    layer1_outputs(9670) <= (layer0_outputs(10006)) xor (layer0_outputs(1284));
    layer1_outputs(9671) <= not((layer0_outputs(7661)) xor (layer0_outputs(4772)));
    layer1_outputs(9672) <= (layer0_outputs(3768)) or (layer0_outputs(602));
    layer1_outputs(9673) <= '0';
    layer1_outputs(9674) <= (layer0_outputs(7885)) and not (layer0_outputs(221));
    layer1_outputs(9675) <= (layer0_outputs(5289)) and (layer0_outputs(4855));
    layer1_outputs(9676) <= layer0_outputs(894);
    layer1_outputs(9677) <= not(layer0_outputs(10126)) or (layer0_outputs(9517));
    layer1_outputs(9678) <= '0';
    layer1_outputs(9679) <= not(layer0_outputs(3403)) or (layer0_outputs(325));
    layer1_outputs(9680) <= '1';
    layer1_outputs(9681) <= (layer0_outputs(8793)) and (layer0_outputs(7734));
    layer1_outputs(9682) <= not((layer0_outputs(2568)) and (layer0_outputs(3634)));
    layer1_outputs(9683) <= (layer0_outputs(6275)) and not (layer0_outputs(8730));
    layer1_outputs(9684) <= (layer0_outputs(5363)) and not (layer0_outputs(3516));
    layer1_outputs(9685) <= '1';
    layer1_outputs(9686) <= layer0_outputs(8626);
    layer1_outputs(9687) <= not((layer0_outputs(2475)) or (layer0_outputs(7459)));
    layer1_outputs(9688) <= not((layer0_outputs(1764)) or (layer0_outputs(7321)));
    layer1_outputs(9689) <= layer0_outputs(2373);
    layer1_outputs(9690) <= layer0_outputs(6254);
    layer1_outputs(9691) <= layer0_outputs(2678);
    layer1_outputs(9692) <= layer0_outputs(5440);
    layer1_outputs(9693) <= (layer0_outputs(6371)) and not (layer0_outputs(105));
    layer1_outputs(9694) <= not((layer0_outputs(391)) or (layer0_outputs(8978)));
    layer1_outputs(9695) <= layer0_outputs(1673);
    layer1_outputs(9696) <= not(layer0_outputs(7044)) or (layer0_outputs(6164));
    layer1_outputs(9697) <= not(layer0_outputs(7329)) or (layer0_outputs(9749));
    layer1_outputs(9698) <= not((layer0_outputs(91)) and (layer0_outputs(3399)));
    layer1_outputs(9699) <= not((layer0_outputs(9812)) xor (layer0_outputs(8915)));
    layer1_outputs(9700) <= not(layer0_outputs(5988));
    layer1_outputs(9701) <= layer0_outputs(991);
    layer1_outputs(9702) <= not(layer0_outputs(4252));
    layer1_outputs(9703) <= (layer0_outputs(6539)) xor (layer0_outputs(271));
    layer1_outputs(9704) <= not(layer0_outputs(6035)) or (layer0_outputs(5448));
    layer1_outputs(9705) <= layer0_outputs(9445);
    layer1_outputs(9706) <= (layer0_outputs(7203)) or (layer0_outputs(8735));
    layer1_outputs(9707) <= layer0_outputs(5325);
    layer1_outputs(9708) <= not((layer0_outputs(9913)) or (layer0_outputs(4416)));
    layer1_outputs(9709) <= layer0_outputs(6603);
    layer1_outputs(9710) <= layer0_outputs(9547);
    layer1_outputs(9711) <= (layer0_outputs(9737)) and (layer0_outputs(5230));
    layer1_outputs(9712) <= not(layer0_outputs(4995));
    layer1_outputs(9713) <= (layer0_outputs(9958)) and not (layer0_outputs(719));
    layer1_outputs(9714) <= layer0_outputs(8672);
    layer1_outputs(9715) <= (layer0_outputs(891)) and (layer0_outputs(8074));
    layer1_outputs(9716) <= not(layer0_outputs(6052));
    layer1_outputs(9717) <= '0';
    layer1_outputs(9718) <= layer0_outputs(1683);
    layer1_outputs(9719) <= '1';
    layer1_outputs(9720) <= layer0_outputs(3788);
    layer1_outputs(9721) <= layer0_outputs(2882);
    layer1_outputs(9722) <= not(layer0_outputs(3955));
    layer1_outputs(9723) <= (layer0_outputs(6565)) or (layer0_outputs(9804));
    layer1_outputs(9724) <= not(layer0_outputs(6747));
    layer1_outputs(9725) <= (layer0_outputs(2346)) or (layer0_outputs(672));
    layer1_outputs(9726) <= (layer0_outputs(3668)) or (layer0_outputs(7329));
    layer1_outputs(9727) <= not((layer0_outputs(3479)) xor (layer0_outputs(5063)));
    layer1_outputs(9728) <= not(layer0_outputs(8533));
    layer1_outputs(9729) <= not(layer0_outputs(6501)) or (layer0_outputs(7890));
    layer1_outputs(9730) <= not(layer0_outputs(9856)) or (layer0_outputs(1028));
    layer1_outputs(9731) <= not(layer0_outputs(9214));
    layer1_outputs(9732) <= not(layer0_outputs(6498)) or (layer0_outputs(2556));
    layer1_outputs(9733) <= (layer0_outputs(6867)) and not (layer0_outputs(3980));
    layer1_outputs(9734) <= not(layer0_outputs(4569)) or (layer0_outputs(6923));
    layer1_outputs(9735) <= (layer0_outputs(4013)) xor (layer0_outputs(8739));
    layer1_outputs(9736) <= '1';
    layer1_outputs(9737) <= layer0_outputs(1289);
    layer1_outputs(9738) <= (layer0_outputs(6822)) or (layer0_outputs(7334));
    layer1_outputs(9739) <= not(layer0_outputs(362));
    layer1_outputs(9740) <= '0';
    layer1_outputs(9741) <= not((layer0_outputs(3386)) or (layer0_outputs(7749)));
    layer1_outputs(9742) <= not((layer0_outputs(1388)) and (layer0_outputs(5138)));
    layer1_outputs(9743) <= '1';
    layer1_outputs(9744) <= (layer0_outputs(948)) or (layer0_outputs(2430));
    layer1_outputs(9745) <= not(layer0_outputs(889));
    layer1_outputs(9746) <= (layer0_outputs(5760)) xor (layer0_outputs(1942));
    layer1_outputs(9747) <= '1';
    layer1_outputs(9748) <= layer0_outputs(2737);
    layer1_outputs(9749) <= not(layer0_outputs(6218)) or (layer0_outputs(9951));
    layer1_outputs(9750) <= not(layer0_outputs(2979)) or (layer0_outputs(3770));
    layer1_outputs(9751) <= '0';
    layer1_outputs(9752) <= (layer0_outputs(3997)) and (layer0_outputs(8599));
    layer1_outputs(9753) <= (layer0_outputs(2545)) or (layer0_outputs(6126));
    layer1_outputs(9754) <= '0';
    layer1_outputs(9755) <= not(layer0_outputs(403)) or (layer0_outputs(1159));
    layer1_outputs(9756) <= not(layer0_outputs(10057)) or (layer0_outputs(7535));
    layer1_outputs(9757) <= not(layer0_outputs(7710));
    layer1_outputs(9758) <= not((layer0_outputs(6038)) or (layer0_outputs(9064)));
    layer1_outputs(9759) <= not(layer0_outputs(6835));
    layer1_outputs(9760) <= layer0_outputs(9866);
    layer1_outputs(9761) <= not((layer0_outputs(10158)) and (layer0_outputs(3564)));
    layer1_outputs(9762) <= layer0_outputs(4249);
    layer1_outputs(9763) <= not(layer0_outputs(5047));
    layer1_outputs(9764) <= layer0_outputs(7286);
    layer1_outputs(9765) <= not(layer0_outputs(1101)) or (layer0_outputs(9854));
    layer1_outputs(9766) <= not(layer0_outputs(7458));
    layer1_outputs(9767) <= (layer0_outputs(2017)) and not (layer0_outputs(10036));
    layer1_outputs(9768) <= (layer0_outputs(5352)) and (layer0_outputs(4577));
    layer1_outputs(9769) <= (layer0_outputs(6651)) or (layer0_outputs(3285));
    layer1_outputs(9770) <= not((layer0_outputs(6971)) and (layer0_outputs(4226)));
    layer1_outputs(9771) <= layer0_outputs(2229);
    layer1_outputs(9772) <= not(layer0_outputs(8855));
    layer1_outputs(9773) <= not(layer0_outputs(10166));
    layer1_outputs(9774) <= (layer0_outputs(9652)) and (layer0_outputs(6901));
    layer1_outputs(9775) <= (layer0_outputs(9102)) and not (layer0_outputs(3322));
    layer1_outputs(9776) <= layer0_outputs(5973);
    layer1_outputs(9777) <= not(layer0_outputs(1910));
    layer1_outputs(9778) <= not(layer0_outputs(8803));
    layer1_outputs(9779) <= not((layer0_outputs(8026)) xor (layer0_outputs(9927)));
    layer1_outputs(9780) <= layer0_outputs(3200);
    layer1_outputs(9781) <= not(layer0_outputs(2002)) or (layer0_outputs(2029));
    layer1_outputs(9782) <= '0';
    layer1_outputs(9783) <= not((layer0_outputs(1229)) and (layer0_outputs(1213)));
    layer1_outputs(9784) <= layer0_outputs(8218);
    layer1_outputs(9785) <= not(layer0_outputs(3602));
    layer1_outputs(9786) <= (layer0_outputs(4938)) and not (layer0_outputs(7079));
    layer1_outputs(9787) <= not(layer0_outputs(8705)) or (layer0_outputs(9002));
    layer1_outputs(9788) <= '0';
    layer1_outputs(9789) <= not((layer0_outputs(1010)) and (layer0_outputs(5743)));
    layer1_outputs(9790) <= layer0_outputs(7569);
    layer1_outputs(9791) <= (layer0_outputs(4803)) or (layer0_outputs(8226));
    layer1_outputs(9792) <= (layer0_outputs(5134)) and not (layer0_outputs(2223));
    layer1_outputs(9793) <= not((layer0_outputs(799)) and (layer0_outputs(7273)));
    layer1_outputs(9794) <= (layer0_outputs(7738)) and (layer0_outputs(2856));
    layer1_outputs(9795) <= layer0_outputs(3145);
    layer1_outputs(9796) <= not((layer0_outputs(2317)) xor (layer0_outputs(8400)));
    layer1_outputs(9797) <= not(layer0_outputs(4741));
    layer1_outputs(9798) <= not(layer0_outputs(4616));
    layer1_outputs(9799) <= not(layer0_outputs(3714)) or (layer0_outputs(7937));
    layer1_outputs(9800) <= not(layer0_outputs(228)) or (layer0_outputs(2315));
    layer1_outputs(9801) <= layer0_outputs(1518);
    layer1_outputs(9802) <= not((layer0_outputs(9580)) xor (layer0_outputs(3331)));
    layer1_outputs(9803) <= (layer0_outputs(8185)) and not (layer0_outputs(3022));
    layer1_outputs(9804) <= not(layer0_outputs(405));
    layer1_outputs(9805) <= '1';
    layer1_outputs(9806) <= not((layer0_outputs(5017)) or (layer0_outputs(7668)));
    layer1_outputs(9807) <= not((layer0_outputs(1252)) xor (layer0_outputs(2686)));
    layer1_outputs(9808) <= not(layer0_outputs(6728));
    layer1_outputs(9809) <= layer0_outputs(4885);
    layer1_outputs(9810) <= not(layer0_outputs(4486)) or (layer0_outputs(2857));
    layer1_outputs(9811) <= (layer0_outputs(4167)) and not (layer0_outputs(9779));
    layer1_outputs(9812) <= (layer0_outputs(9787)) xor (layer0_outputs(2865));
    layer1_outputs(9813) <= not(layer0_outputs(2794)) or (layer0_outputs(7820));
    layer1_outputs(9814) <= (layer0_outputs(4963)) or (layer0_outputs(7491));
    layer1_outputs(9815) <= layer0_outputs(4924);
    layer1_outputs(9816) <= (layer0_outputs(9188)) and not (layer0_outputs(4280));
    layer1_outputs(9817) <= not(layer0_outputs(8620));
    layer1_outputs(9818) <= (layer0_outputs(3116)) and not (layer0_outputs(8882));
    layer1_outputs(9819) <= not(layer0_outputs(5467));
    layer1_outputs(9820) <= not((layer0_outputs(9648)) xor (layer0_outputs(3585)));
    layer1_outputs(9821) <= (layer0_outputs(1092)) or (layer0_outputs(276));
    layer1_outputs(9822) <= (layer0_outputs(9463)) and (layer0_outputs(6250));
    layer1_outputs(9823) <= not(layer0_outputs(3624));
    layer1_outputs(9824) <= not(layer0_outputs(7441));
    layer1_outputs(9825) <= (layer0_outputs(4828)) and not (layer0_outputs(5693));
    layer1_outputs(9826) <= not((layer0_outputs(6281)) and (layer0_outputs(6466)));
    layer1_outputs(9827) <= (layer0_outputs(8505)) and (layer0_outputs(6176));
    layer1_outputs(9828) <= not(layer0_outputs(4228));
    layer1_outputs(9829) <= not(layer0_outputs(1485));
    layer1_outputs(9830) <= layer0_outputs(718);
    layer1_outputs(9831) <= (layer0_outputs(7514)) and not (layer0_outputs(4858));
    layer1_outputs(9832) <= not(layer0_outputs(3864));
    layer1_outputs(9833) <= not(layer0_outputs(964)) or (layer0_outputs(10159));
    layer1_outputs(9834) <= not(layer0_outputs(2859));
    layer1_outputs(9835) <= '0';
    layer1_outputs(9836) <= not(layer0_outputs(2274));
    layer1_outputs(9837) <= layer0_outputs(6570);
    layer1_outputs(9838) <= layer0_outputs(9151);
    layer1_outputs(9839) <= not((layer0_outputs(6486)) or (layer0_outputs(1622)));
    layer1_outputs(9840) <= (layer0_outputs(6993)) or (layer0_outputs(1150));
    layer1_outputs(9841) <= not((layer0_outputs(2119)) or (layer0_outputs(5587)));
    layer1_outputs(9842) <= not(layer0_outputs(1589));
    layer1_outputs(9843) <= '1';
    layer1_outputs(9844) <= layer0_outputs(9967);
    layer1_outputs(9845) <= not((layer0_outputs(1650)) and (layer0_outputs(3319)));
    layer1_outputs(9846) <= not((layer0_outputs(9318)) and (layer0_outputs(8163)));
    layer1_outputs(9847) <= layer0_outputs(10208);
    layer1_outputs(9848) <= not(layer0_outputs(7901)) or (layer0_outputs(279));
    layer1_outputs(9849) <= not((layer0_outputs(6220)) or (layer0_outputs(798)));
    layer1_outputs(9850) <= (layer0_outputs(2996)) xor (layer0_outputs(4306));
    layer1_outputs(9851) <= (layer0_outputs(7411)) xor (layer0_outputs(1223));
    layer1_outputs(9852) <= not((layer0_outputs(9727)) or (layer0_outputs(5633)));
    layer1_outputs(9853) <= not((layer0_outputs(6031)) or (layer0_outputs(3462)));
    layer1_outputs(9854) <= not(layer0_outputs(7152));
    layer1_outputs(9855) <= not((layer0_outputs(2416)) and (layer0_outputs(1962)));
    layer1_outputs(9856) <= (layer0_outputs(3665)) and (layer0_outputs(8372));
    layer1_outputs(9857) <= not(layer0_outputs(2242));
    layer1_outputs(9858) <= layer0_outputs(1559);
    layer1_outputs(9859) <= (layer0_outputs(4710)) xor (layer0_outputs(4959));
    layer1_outputs(9860) <= (layer0_outputs(1938)) and (layer0_outputs(600));
    layer1_outputs(9861) <= not((layer0_outputs(5986)) and (layer0_outputs(6969)));
    layer1_outputs(9862) <= layer0_outputs(2342);
    layer1_outputs(9863) <= (layer0_outputs(9264)) and not (layer0_outputs(9650));
    layer1_outputs(9864) <= (layer0_outputs(8973)) and (layer0_outputs(10156));
    layer1_outputs(9865) <= not(layer0_outputs(7084)) or (layer0_outputs(2397));
    layer1_outputs(9866) <= not(layer0_outputs(928)) or (layer0_outputs(9105));
    layer1_outputs(9867) <= not(layer0_outputs(3793));
    layer1_outputs(9868) <= (layer0_outputs(4511)) and not (layer0_outputs(6729));
    layer1_outputs(9869) <= '1';
    layer1_outputs(9870) <= not(layer0_outputs(1662));
    layer1_outputs(9871) <= (layer0_outputs(7413)) and not (layer0_outputs(5706));
    layer1_outputs(9872) <= not(layer0_outputs(2982)) or (layer0_outputs(6335));
    layer1_outputs(9873) <= not(layer0_outputs(3631));
    layer1_outputs(9874) <= (layer0_outputs(721)) and not (layer0_outputs(623));
    layer1_outputs(9875) <= not(layer0_outputs(9314));
    layer1_outputs(9876) <= layer0_outputs(3127);
    layer1_outputs(9877) <= (layer0_outputs(125)) xor (layer0_outputs(3048));
    layer1_outputs(9878) <= not(layer0_outputs(193));
    layer1_outputs(9879) <= (layer0_outputs(4464)) xor (layer0_outputs(3458));
    layer1_outputs(9880) <= (layer0_outputs(5154)) and not (layer0_outputs(3712));
    layer1_outputs(9881) <= layer0_outputs(9890);
    layer1_outputs(9882) <= not((layer0_outputs(9573)) and (layer0_outputs(9544)));
    layer1_outputs(9883) <= '0';
    layer1_outputs(9884) <= layer0_outputs(331);
    layer1_outputs(9885) <= not(layer0_outputs(6420)) or (layer0_outputs(4575));
    layer1_outputs(9886) <= not((layer0_outputs(7502)) or (layer0_outputs(8696)));
    layer1_outputs(9887) <= not(layer0_outputs(5990));
    layer1_outputs(9888) <= not((layer0_outputs(2956)) and (layer0_outputs(8282)));
    layer1_outputs(9889) <= not((layer0_outputs(107)) xor (layer0_outputs(1643)));
    layer1_outputs(9890) <= not(layer0_outputs(9037));
    layer1_outputs(9891) <= (layer0_outputs(9633)) and (layer0_outputs(4369));
    layer1_outputs(9892) <= not(layer0_outputs(6160)) or (layer0_outputs(1692));
    layer1_outputs(9893) <= not(layer0_outputs(8116)) or (layer0_outputs(3604));
    layer1_outputs(9894) <= (layer0_outputs(8117)) and not (layer0_outputs(6528));
    layer1_outputs(9895) <= (layer0_outputs(2239)) xor (layer0_outputs(2382));
    layer1_outputs(9896) <= (layer0_outputs(6597)) and (layer0_outputs(2694));
    layer1_outputs(9897) <= not(layer0_outputs(5108));
    layer1_outputs(9898) <= not((layer0_outputs(6508)) xor (layer0_outputs(163)));
    layer1_outputs(9899) <= not((layer0_outputs(2579)) xor (layer0_outputs(9001)));
    layer1_outputs(9900) <= '0';
    layer1_outputs(9901) <= (layer0_outputs(1391)) or (layer0_outputs(8890));
    layer1_outputs(9902) <= (layer0_outputs(8098)) and (layer0_outputs(2294));
    layer1_outputs(9903) <= (layer0_outputs(2727)) and not (layer0_outputs(5349));
    layer1_outputs(9904) <= not((layer0_outputs(9975)) and (layer0_outputs(1449)));
    layer1_outputs(9905) <= not((layer0_outputs(3759)) and (layer0_outputs(3762)));
    layer1_outputs(9906) <= layer0_outputs(8341);
    layer1_outputs(9907) <= not(layer0_outputs(4042));
    layer1_outputs(9908) <= not(layer0_outputs(7097)) or (layer0_outputs(10180));
    layer1_outputs(9909) <= not(layer0_outputs(1438)) or (layer0_outputs(9128));
    layer1_outputs(9910) <= not(layer0_outputs(9899)) or (layer0_outputs(5941));
    layer1_outputs(9911) <= (layer0_outputs(5686)) or (layer0_outputs(3035));
    layer1_outputs(9912) <= layer0_outputs(4557);
    layer1_outputs(9913) <= not(layer0_outputs(4988));
    layer1_outputs(9914) <= '1';
    layer1_outputs(9915) <= not(layer0_outputs(11));
    layer1_outputs(9916) <= layer0_outputs(4648);
    layer1_outputs(9917) <= (layer0_outputs(7979)) and (layer0_outputs(1695));
    layer1_outputs(9918) <= layer0_outputs(1511);
    layer1_outputs(9919) <= layer0_outputs(9264);
    layer1_outputs(9920) <= not(layer0_outputs(2784)) or (layer0_outputs(538));
    layer1_outputs(9921) <= not((layer0_outputs(3864)) or (layer0_outputs(3118)));
    layer1_outputs(9922) <= not((layer0_outputs(6949)) or (layer0_outputs(9168)));
    layer1_outputs(9923) <= not((layer0_outputs(872)) xor (layer0_outputs(10095)));
    layer1_outputs(9924) <= (layer0_outputs(6005)) and not (layer0_outputs(294));
    layer1_outputs(9925) <= not(layer0_outputs(5253)) or (layer0_outputs(1495));
    layer1_outputs(9926) <= not(layer0_outputs(3508));
    layer1_outputs(9927) <= not(layer0_outputs(3749)) or (layer0_outputs(2225));
    layer1_outputs(9928) <= not((layer0_outputs(597)) and (layer0_outputs(6797)));
    layer1_outputs(9929) <= not(layer0_outputs(9643)) or (layer0_outputs(8265));
    layer1_outputs(9930) <= not(layer0_outputs(4948));
    layer1_outputs(9931) <= not(layer0_outputs(4478)) or (layer0_outputs(5644));
    layer1_outputs(9932) <= not((layer0_outputs(9732)) or (layer0_outputs(1166)));
    layer1_outputs(9933) <= layer0_outputs(5779);
    layer1_outputs(9934) <= not(layer0_outputs(3709));
    layer1_outputs(9935) <= not(layer0_outputs(9324));
    layer1_outputs(9936) <= not(layer0_outputs(4099)) or (layer0_outputs(9911));
    layer1_outputs(9937) <= not((layer0_outputs(8850)) or (layer0_outputs(6931)));
    layer1_outputs(9938) <= (layer0_outputs(6791)) and not (layer0_outputs(6938));
    layer1_outputs(9939) <= not(layer0_outputs(7586)) or (layer0_outputs(7031));
    layer1_outputs(9940) <= not((layer0_outputs(2940)) or (layer0_outputs(9303)));
    layer1_outputs(9941) <= (layer0_outputs(4035)) and (layer0_outputs(4666));
    layer1_outputs(9942) <= (layer0_outputs(3786)) and (layer0_outputs(9949));
    layer1_outputs(9943) <= not(layer0_outputs(9656)) or (layer0_outputs(4330));
    layer1_outputs(9944) <= layer0_outputs(9574);
    layer1_outputs(9945) <= layer0_outputs(7642);
    layer1_outputs(9946) <= (layer0_outputs(4091)) or (layer0_outputs(3136));
    layer1_outputs(9947) <= (layer0_outputs(14)) and not (layer0_outputs(7255));
    layer1_outputs(9948) <= not((layer0_outputs(1198)) xor (layer0_outputs(3842)));
    layer1_outputs(9949) <= '1';
    layer1_outputs(9950) <= (layer0_outputs(2249)) and (layer0_outputs(8557));
    layer1_outputs(9951) <= not(layer0_outputs(7600)) or (layer0_outputs(3289));
    layer1_outputs(9952) <= (layer0_outputs(2726)) and not (layer0_outputs(1961));
    layer1_outputs(9953) <= not(layer0_outputs(7219)) or (layer0_outputs(8628));
    layer1_outputs(9954) <= layer0_outputs(7006);
    layer1_outputs(9955) <= not((layer0_outputs(3303)) or (layer0_outputs(1973)));
    layer1_outputs(9956) <= (layer0_outputs(7386)) and not (layer0_outputs(800));
    layer1_outputs(9957) <= (layer0_outputs(2973)) or (layer0_outputs(5076));
    layer1_outputs(9958) <= not(layer0_outputs(109)) or (layer0_outputs(8629));
    layer1_outputs(9959) <= '1';
    layer1_outputs(9960) <= not(layer0_outputs(5418)) or (layer0_outputs(7501));
    layer1_outputs(9961) <= not((layer0_outputs(7200)) and (layer0_outputs(1090)));
    layer1_outputs(9962) <= not((layer0_outputs(4214)) or (layer0_outputs(10143)));
    layer1_outputs(9963) <= layer0_outputs(7723);
    layer1_outputs(9964) <= (layer0_outputs(666)) and (layer0_outputs(2318));
    layer1_outputs(9965) <= not(layer0_outputs(5777));
    layer1_outputs(9966) <= (layer0_outputs(7348)) xor (layer0_outputs(9683));
    layer1_outputs(9967) <= not((layer0_outputs(4144)) or (layer0_outputs(3296)));
    layer1_outputs(9968) <= not(layer0_outputs(6792));
    layer1_outputs(9969) <= layer0_outputs(6412);
    layer1_outputs(9970) <= not((layer0_outputs(1124)) xor (layer0_outputs(8059)));
    layer1_outputs(9971) <= not(layer0_outputs(3451));
    layer1_outputs(9972) <= (layer0_outputs(673)) xor (layer0_outputs(3113));
    layer1_outputs(9973) <= not(layer0_outputs(1730));
    layer1_outputs(9974) <= not(layer0_outputs(2887));
    layer1_outputs(9975) <= layer0_outputs(9423);
    layer1_outputs(9976) <= (layer0_outputs(1648)) or (layer0_outputs(10194));
    layer1_outputs(9977) <= layer0_outputs(6064);
    layer1_outputs(9978) <= '0';
    layer1_outputs(9979) <= not(layer0_outputs(3845)) or (layer0_outputs(7989));
    layer1_outputs(9980) <= layer0_outputs(7645);
    layer1_outputs(9981) <= (layer0_outputs(280)) and (layer0_outputs(9502));
    layer1_outputs(9982) <= not(layer0_outputs(6051));
    layer1_outputs(9983) <= layer0_outputs(3478);
    layer1_outputs(9984) <= layer0_outputs(9849);
    layer1_outputs(9985) <= not(layer0_outputs(387)) or (layer0_outputs(7520));
    layer1_outputs(9986) <= not((layer0_outputs(5569)) or (layer0_outputs(6681)));
    layer1_outputs(9987) <= not(layer0_outputs(1696)) or (layer0_outputs(6113));
    layer1_outputs(9988) <= not(layer0_outputs(211)) or (layer0_outputs(4278));
    layer1_outputs(9989) <= (layer0_outputs(2703)) and (layer0_outputs(5670));
    layer1_outputs(9990) <= not(layer0_outputs(3185));
    layer1_outputs(9991) <= layer0_outputs(2587);
    layer1_outputs(9992) <= (layer0_outputs(8263)) or (layer0_outputs(7417));
    layer1_outputs(9993) <= not(layer0_outputs(5403));
    layer1_outputs(9994) <= (layer0_outputs(2413)) and not (layer0_outputs(2044));
    layer1_outputs(9995) <= not((layer0_outputs(4482)) or (layer0_outputs(4005)));
    layer1_outputs(9996) <= layer0_outputs(4199);
    layer1_outputs(9997) <= (layer0_outputs(8131)) and not (layer0_outputs(5643));
    layer1_outputs(9998) <= not(layer0_outputs(7801)) or (layer0_outputs(6344));
    layer1_outputs(9999) <= '1';
    layer1_outputs(10000) <= not(layer0_outputs(4421));
    layer1_outputs(10001) <= (layer0_outputs(5134)) and (layer0_outputs(9359));
    layer1_outputs(10002) <= not((layer0_outputs(6336)) or (layer0_outputs(8558)));
    layer1_outputs(10003) <= not((layer0_outputs(6321)) or (layer0_outputs(8110)));
    layer1_outputs(10004) <= not(layer0_outputs(9064));
    layer1_outputs(10005) <= layer0_outputs(8409);
    layer1_outputs(10006) <= layer0_outputs(8528);
    layer1_outputs(10007) <= (layer0_outputs(3908)) and not (layer0_outputs(7544));
    layer1_outputs(10008) <= not((layer0_outputs(506)) xor (layer0_outputs(761)));
    layer1_outputs(10009) <= not(layer0_outputs(7302));
    layer1_outputs(10010) <= not((layer0_outputs(401)) and (layer0_outputs(2854)));
    layer1_outputs(10011) <= (layer0_outputs(6045)) or (layer0_outputs(5996));
    layer1_outputs(10012) <= not(layer0_outputs(1889));
    layer1_outputs(10013) <= not(layer0_outputs(3652));
    layer1_outputs(10014) <= '1';
    layer1_outputs(10015) <= not(layer0_outputs(1142));
    layer1_outputs(10016) <= layer0_outputs(7822);
    layer1_outputs(10017) <= not(layer0_outputs(411));
    layer1_outputs(10018) <= not(layer0_outputs(977));
    layer1_outputs(10019) <= not(layer0_outputs(8456)) or (layer0_outputs(9704));
    layer1_outputs(10020) <= not(layer0_outputs(891));
    layer1_outputs(10021) <= layer0_outputs(4063);
    layer1_outputs(10022) <= not(layer0_outputs(6469));
    layer1_outputs(10023) <= (layer0_outputs(1631)) or (layer0_outputs(7969));
    layer1_outputs(10024) <= not(layer0_outputs(3545));
    layer1_outputs(10025) <= (layer0_outputs(297)) xor (layer0_outputs(1847));
    layer1_outputs(10026) <= '1';
    layer1_outputs(10027) <= (layer0_outputs(2501)) or (layer0_outputs(4464));
    layer1_outputs(10028) <= not((layer0_outputs(10031)) or (layer0_outputs(2392)));
    layer1_outputs(10029) <= not(layer0_outputs(4745));
    layer1_outputs(10030) <= not((layer0_outputs(1123)) and (layer0_outputs(1268)));
    layer1_outputs(10031) <= not(layer0_outputs(8796));
    layer1_outputs(10032) <= not(layer0_outputs(9107));
    layer1_outputs(10033) <= not(layer0_outputs(1997));
    layer1_outputs(10034) <= layer0_outputs(7198);
    layer1_outputs(10035) <= layer0_outputs(379);
    layer1_outputs(10036) <= (layer0_outputs(40)) or (layer0_outputs(9886));
    layer1_outputs(10037) <= not(layer0_outputs(2506));
    layer1_outputs(10038) <= (layer0_outputs(10049)) or (layer0_outputs(6343));
    layer1_outputs(10039) <= (layer0_outputs(5416)) or (layer0_outputs(6194));
    layer1_outputs(10040) <= not(layer0_outputs(9733));
    layer1_outputs(10041) <= (layer0_outputs(1288)) and not (layer0_outputs(1135));
    layer1_outputs(10042) <= '0';
    layer1_outputs(10043) <= layer0_outputs(8641);
    layer1_outputs(10044) <= (layer0_outputs(2813)) and not (layer0_outputs(6024));
    layer1_outputs(10045) <= not((layer0_outputs(4958)) xor (layer0_outputs(9036)));
    layer1_outputs(10046) <= not(layer0_outputs(7010));
    layer1_outputs(10047) <= not(layer0_outputs(9756));
    layer1_outputs(10048) <= (layer0_outputs(6733)) and not (layer0_outputs(5575));
    layer1_outputs(10049) <= (layer0_outputs(6952)) and not (layer0_outputs(4472));
    layer1_outputs(10050) <= '1';
    layer1_outputs(10051) <= not(layer0_outputs(9344));
    layer1_outputs(10052) <= layer0_outputs(3886);
    layer1_outputs(10053) <= layer0_outputs(6010);
    layer1_outputs(10054) <= (layer0_outputs(4747)) or (layer0_outputs(952));
    layer1_outputs(10055) <= (layer0_outputs(2247)) and (layer0_outputs(3806));
    layer1_outputs(10056) <= not(layer0_outputs(5550)) or (layer0_outputs(5713));
    layer1_outputs(10057) <= not(layer0_outputs(2781)) or (layer0_outputs(376));
    layer1_outputs(10058) <= not(layer0_outputs(3243));
    layer1_outputs(10059) <= (layer0_outputs(1432)) and (layer0_outputs(8510));
    layer1_outputs(10060) <= layer0_outputs(8720);
    layer1_outputs(10061) <= layer0_outputs(3779);
    layer1_outputs(10062) <= not(layer0_outputs(9297)) or (layer0_outputs(4677));
    layer1_outputs(10063) <= '1';
    layer1_outputs(10064) <= (layer0_outputs(3673)) and not (layer0_outputs(2071));
    layer1_outputs(10065) <= (layer0_outputs(3602)) and not (layer0_outputs(176));
    layer1_outputs(10066) <= not(layer0_outputs(9262));
    layer1_outputs(10067) <= not(layer0_outputs(5902));
    layer1_outputs(10068) <= layer0_outputs(5906);
    layer1_outputs(10069) <= not(layer0_outputs(8166));
    layer1_outputs(10070) <= not(layer0_outputs(1627));
    layer1_outputs(10071) <= not(layer0_outputs(6407));
    layer1_outputs(10072) <= not((layer0_outputs(8505)) or (layer0_outputs(9613)));
    layer1_outputs(10073) <= not(layer0_outputs(4200));
    layer1_outputs(10074) <= not(layer0_outputs(7076)) or (layer0_outputs(8249));
    layer1_outputs(10075) <= layer0_outputs(999);
    layer1_outputs(10076) <= '1';
    layer1_outputs(10077) <= layer0_outputs(1474);
    layer1_outputs(10078) <= not(layer0_outputs(7426)) or (layer0_outputs(839));
    layer1_outputs(10079) <= '0';
    layer1_outputs(10080) <= layer0_outputs(515);
    layer1_outputs(10081) <= not(layer0_outputs(2060));
    layer1_outputs(10082) <= not(layer0_outputs(1716));
    layer1_outputs(10083) <= not(layer0_outputs(4320)) or (layer0_outputs(5071));
    layer1_outputs(10084) <= not(layer0_outputs(7455));
    layer1_outputs(10085) <= not(layer0_outputs(2878));
    layer1_outputs(10086) <= not((layer0_outputs(6257)) and (layer0_outputs(3822)));
    layer1_outputs(10087) <= layer0_outputs(4800);
    layer1_outputs(10088) <= not((layer0_outputs(5302)) xor (layer0_outputs(9444)));
    layer1_outputs(10089) <= '1';
    layer1_outputs(10090) <= not(layer0_outputs(5613));
    layer1_outputs(10091) <= not((layer0_outputs(4986)) or (layer0_outputs(5896)));
    layer1_outputs(10092) <= not(layer0_outputs(3517)) or (layer0_outputs(10122));
    layer1_outputs(10093) <= not(layer0_outputs(9653));
    layer1_outputs(10094) <= not((layer0_outputs(457)) or (layer0_outputs(9400)));
    layer1_outputs(10095) <= not((layer0_outputs(7978)) and (layer0_outputs(5094)));
    layer1_outputs(10096) <= (layer0_outputs(4774)) or (layer0_outputs(7228));
    layer1_outputs(10097) <= (layer0_outputs(6724)) and not (layer0_outputs(2132));
    layer1_outputs(10098) <= (layer0_outputs(6761)) or (layer0_outputs(4161));
    layer1_outputs(10099) <= (layer0_outputs(4711)) and not (layer0_outputs(3327));
    layer1_outputs(10100) <= layer0_outputs(8991);
    layer1_outputs(10101) <= not((layer0_outputs(8086)) xor (layer0_outputs(5968)));
    layer1_outputs(10102) <= (layer0_outputs(2109)) or (layer0_outputs(7444));
    layer1_outputs(10103) <= not(layer0_outputs(5338)) or (layer0_outputs(1073));
    layer1_outputs(10104) <= not(layer0_outputs(6098));
    layer1_outputs(10105) <= layer0_outputs(9211);
    layer1_outputs(10106) <= (layer0_outputs(6818)) and not (layer0_outputs(7133));
    layer1_outputs(10107) <= layer0_outputs(7339);
    layer1_outputs(10108) <= not(layer0_outputs(7641)) or (layer0_outputs(8798));
    layer1_outputs(10109) <= not(layer0_outputs(5326));
    layer1_outputs(10110) <= layer0_outputs(5081);
    layer1_outputs(10111) <= not(layer0_outputs(7420));
    layer1_outputs(10112) <= not(layer0_outputs(5607));
    layer1_outputs(10113) <= '1';
    layer1_outputs(10114) <= not((layer0_outputs(6039)) or (layer0_outputs(9632)));
    layer1_outputs(10115) <= layer0_outputs(1316);
    layer1_outputs(10116) <= not((layer0_outputs(1382)) and (layer0_outputs(541)));
    layer1_outputs(10117) <= not((layer0_outputs(5157)) or (layer0_outputs(3426)));
    layer1_outputs(10118) <= layer0_outputs(3040);
    layer1_outputs(10119) <= (layer0_outputs(5070)) and (layer0_outputs(4941));
    layer1_outputs(10120) <= not(layer0_outputs(2390));
    layer1_outputs(10121) <= (layer0_outputs(8030)) and not (layer0_outputs(8736));
    layer1_outputs(10122) <= layer0_outputs(1033);
    layer1_outputs(10123) <= (layer0_outputs(5914)) xor (layer0_outputs(9750));
    layer1_outputs(10124) <= (layer0_outputs(6280)) and (layer0_outputs(167));
    layer1_outputs(10125) <= '1';
    layer1_outputs(10126) <= (layer0_outputs(7119)) xor (layer0_outputs(8232));
    layer1_outputs(10127) <= layer0_outputs(5248);
    layer1_outputs(10128) <= (layer0_outputs(3195)) or (layer0_outputs(6904));
    layer1_outputs(10129) <= (layer0_outputs(1349)) and not (layer0_outputs(9938));
    layer1_outputs(10130) <= not((layer0_outputs(1809)) and (layer0_outputs(1488)));
    layer1_outputs(10131) <= not((layer0_outputs(2442)) and (layer0_outputs(3842)));
    layer1_outputs(10132) <= not(layer0_outputs(1429)) or (layer0_outputs(9687));
    layer1_outputs(10133) <= layer0_outputs(91);
    layer1_outputs(10134) <= (layer0_outputs(2231)) and not (layer0_outputs(8989));
    layer1_outputs(10135) <= not(layer0_outputs(8289)) or (layer0_outputs(6285));
    layer1_outputs(10136) <= (layer0_outputs(4158)) or (layer0_outputs(544));
    layer1_outputs(10137) <= layer0_outputs(6533);
    layer1_outputs(10138) <= not(layer0_outputs(3306)) or (layer0_outputs(9754));
    layer1_outputs(10139) <= layer0_outputs(3262);
    layer1_outputs(10140) <= not(layer0_outputs(6852)) or (layer0_outputs(8749));
    layer1_outputs(10141) <= (layer0_outputs(8223)) or (layer0_outputs(336));
    layer1_outputs(10142) <= layer0_outputs(7569);
    layer1_outputs(10143) <= not(layer0_outputs(3810));
    layer1_outputs(10144) <= not(layer0_outputs(5383));
    layer1_outputs(10145) <= (layer0_outputs(2820)) or (layer0_outputs(6208));
    layer1_outputs(10146) <= layer0_outputs(8910);
    layer1_outputs(10147) <= not((layer0_outputs(7532)) xor (layer0_outputs(8897)));
    layer1_outputs(10148) <= layer0_outputs(8935);
    layer1_outputs(10149) <= layer0_outputs(495);
    layer1_outputs(10150) <= '0';
    layer1_outputs(10151) <= not(layer0_outputs(10040)) or (layer0_outputs(8222));
    layer1_outputs(10152) <= not(layer0_outputs(5029)) or (layer0_outputs(4235));
    layer1_outputs(10153) <= not(layer0_outputs(7753)) or (layer0_outputs(7948));
    layer1_outputs(10154) <= '1';
    layer1_outputs(10155) <= (layer0_outputs(9954)) or (layer0_outputs(2765));
    layer1_outputs(10156) <= not((layer0_outputs(9141)) or (layer0_outputs(4016)));
    layer1_outputs(10157) <= not(layer0_outputs(873)) or (layer0_outputs(1184));
    layer1_outputs(10158) <= layer0_outputs(4654);
    layer1_outputs(10159) <= not(layer0_outputs(1701));
    layer1_outputs(10160) <= (layer0_outputs(4517)) and not (layer0_outputs(2198));
    layer1_outputs(10161) <= layer0_outputs(4852);
    layer1_outputs(10162) <= (layer0_outputs(1347)) and (layer0_outputs(1770));
    layer1_outputs(10163) <= layer0_outputs(1818);
    layer1_outputs(10164) <= not(layer0_outputs(7682)) or (layer0_outputs(97));
    layer1_outputs(10165) <= not(layer0_outputs(3235));
    layer1_outputs(10166) <= not(layer0_outputs(7443));
    layer1_outputs(10167) <= layer0_outputs(2145);
    layer1_outputs(10168) <= (layer0_outputs(4377)) and not (layer0_outputs(4201));
    layer1_outputs(10169) <= (layer0_outputs(4219)) and not (layer0_outputs(7078));
    layer1_outputs(10170) <= layer0_outputs(1530);
    layer1_outputs(10171) <= layer0_outputs(1885);
    layer1_outputs(10172) <= (layer0_outputs(9431)) xor (layer0_outputs(2155));
    layer1_outputs(10173) <= not(layer0_outputs(8526)) or (layer0_outputs(659));
    layer1_outputs(10174) <= '1';
    layer1_outputs(10175) <= not((layer0_outputs(9233)) xor (layer0_outputs(10074)));
    layer1_outputs(10176) <= (layer0_outputs(5615)) and not (layer0_outputs(126));
    layer1_outputs(10177) <= not(layer0_outputs(1383));
    layer1_outputs(10178) <= layer0_outputs(9701);
    layer1_outputs(10179) <= (layer0_outputs(986)) and not (layer0_outputs(3191));
    layer1_outputs(10180) <= (layer0_outputs(964)) xor (layer0_outputs(4025));
    layer1_outputs(10181) <= layer0_outputs(6409);
    layer1_outputs(10182) <= (layer0_outputs(8171)) and not (layer0_outputs(7395));
    layer1_outputs(10183) <= (layer0_outputs(3783)) and not (layer0_outputs(7005));
    layer1_outputs(10184) <= layer0_outputs(534);
    layer1_outputs(10185) <= not(layer0_outputs(4681)) or (layer0_outputs(2802));
    layer1_outputs(10186) <= (layer0_outputs(8386)) and not (layer0_outputs(3408));
    layer1_outputs(10187) <= not(layer0_outputs(228)) or (layer0_outputs(5100));
    layer1_outputs(10188) <= not(layer0_outputs(8064));
    layer1_outputs(10189) <= not(layer0_outputs(4125));
    layer1_outputs(10190) <= (layer0_outputs(6914)) and (layer0_outputs(4295));
    layer1_outputs(10191) <= not(layer0_outputs(3318));
    layer1_outputs(10192) <= not((layer0_outputs(5765)) or (layer0_outputs(5750)));
    layer1_outputs(10193) <= layer0_outputs(8926);
    layer1_outputs(10194) <= '0';
    layer1_outputs(10195) <= (layer0_outputs(1550)) and not (layer0_outputs(327));
    layer1_outputs(10196) <= not(layer0_outputs(7024)) or (layer0_outputs(953));
    layer1_outputs(10197) <= layer0_outputs(706);
    layer1_outputs(10198) <= not((layer0_outputs(2435)) and (layer0_outputs(4880)));
    layer1_outputs(10199) <= (layer0_outputs(81)) and not (layer0_outputs(5788));
    layer1_outputs(10200) <= (layer0_outputs(4084)) or (layer0_outputs(1446));
    layer1_outputs(10201) <= (layer0_outputs(934)) and not (layer0_outputs(8415));
    layer1_outputs(10202) <= (layer0_outputs(487)) xor (layer0_outputs(3525));
    layer1_outputs(10203) <= not(layer0_outputs(7838));
    layer1_outputs(10204) <= not(layer0_outputs(790)) or (layer0_outputs(1931));
    layer1_outputs(10205) <= '1';
    layer1_outputs(10206) <= not(layer0_outputs(7532)) or (layer0_outputs(822));
    layer1_outputs(10207) <= layer0_outputs(9918);
    layer1_outputs(10208) <= '0';
    layer1_outputs(10209) <= not(layer0_outputs(6567));
    layer1_outputs(10210) <= (layer0_outputs(424)) and (layer0_outputs(1710));
    layer1_outputs(10211) <= not((layer0_outputs(6721)) and (layer0_outputs(8285)));
    layer1_outputs(10212) <= layer0_outputs(6706);
    layer1_outputs(10213) <= (layer0_outputs(4417)) xor (layer0_outputs(1563));
    layer1_outputs(10214) <= (layer0_outputs(7681)) and not (layer0_outputs(3971));
    layer1_outputs(10215) <= (layer0_outputs(3942)) and not (layer0_outputs(6608));
    layer1_outputs(10216) <= not(layer0_outputs(3654));
    layer1_outputs(10217) <= not(layer0_outputs(1598)) or (layer0_outputs(8908));
    layer1_outputs(10218) <= '0';
    layer1_outputs(10219) <= not(layer0_outputs(10044)) or (layer0_outputs(8887));
    layer1_outputs(10220) <= layer0_outputs(66);
    layer1_outputs(10221) <= (layer0_outputs(2561)) and not (layer0_outputs(9832));
    layer1_outputs(10222) <= not((layer0_outputs(1720)) xor (layer0_outputs(6072)));
    layer1_outputs(10223) <= not(layer0_outputs(3123)) or (layer0_outputs(7251));
    layer1_outputs(10224) <= not(layer0_outputs(5487));
    layer1_outputs(10225) <= not(layer0_outputs(9892));
    layer1_outputs(10226) <= not(layer0_outputs(8363)) or (layer0_outputs(6356));
    layer1_outputs(10227) <= not((layer0_outputs(7378)) xor (layer0_outputs(378)));
    layer1_outputs(10228) <= (layer0_outputs(9040)) and not (layer0_outputs(6024));
    layer1_outputs(10229) <= not((layer0_outputs(9243)) xor (layer0_outputs(3537)));
    layer1_outputs(10230) <= layer0_outputs(9737);
    layer1_outputs(10231) <= layer0_outputs(1998);
    layer1_outputs(10232) <= not((layer0_outputs(3834)) or (layer0_outputs(5320)));
    layer1_outputs(10233) <= '1';
    layer1_outputs(10234) <= (layer0_outputs(4669)) and not (layer0_outputs(8755));
    layer1_outputs(10235) <= not(layer0_outputs(5591));
    layer1_outputs(10236) <= not(layer0_outputs(423));
    layer1_outputs(10237) <= not(layer0_outputs(3153));
    layer1_outputs(10238) <= layer0_outputs(5982);
    layer1_outputs(10239) <= not((layer0_outputs(8071)) and (layer0_outputs(5444)));
    layer2_outputs(0) <= not(layer1_outputs(8766));
    layer2_outputs(1) <= (layer1_outputs(1498)) or (layer1_outputs(8510));
    layer2_outputs(2) <= not(layer1_outputs(2656));
    layer2_outputs(3) <= layer1_outputs(9059);
    layer2_outputs(4) <= (layer1_outputs(2296)) and not (layer1_outputs(1705));
    layer2_outputs(5) <= layer1_outputs(6741);
    layer2_outputs(6) <= (layer1_outputs(2210)) and not (layer1_outputs(3746));
    layer2_outputs(7) <= layer1_outputs(3459);
    layer2_outputs(8) <= layer1_outputs(6102);
    layer2_outputs(9) <= layer1_outputs(7495);
    layer2_outputs(10) <= (layer1_outputs(8485)) or (layer1_outputs(3702));
    layer2_outputs(11) <= not(layer1_outputs(6093));
    layer2_outputs(12) <= not(layer1_outputs(3965)) or (layer1_outputs(2039));
    layer2_outputs(13) <= (layer1_outputs(8239)) or (layer1_outputs(1354));
    layer2_outputs(14) <= not(layer1_outputs(6396));
    layer2_outputs(15) <= not(layer1_outputs(398)) or (layer1_outputs(1929));
    layer2_outputs(16) <= not(layer1_outputs(8357)) or (layer1_outputs(5612));
    layer2_outputs(17) <= (layer1_outputs(1644)) and not (layer1_outputs(5111));
    layer2_outputs(18) <= '0';
    layer2_outputs(19) <= '1';
    layer2_outputs(20) <= layer1_outputs(5962);
    layer2_outputs(21) <= '0';
    layer2_outputs(22) <= layer1_outputs(8851);
    layer2_outputs(23) <= (layer1_outputs(4255)) and (layer1_outputs(1019));
    layer2_outputs(24) <= (layer1_outputs(6571)) and (layer1_outputs(6219));
    layer2_outputs(25) <= not(layer1_outputs(6372)) or (layer1_outputs(8125));
    layer2_outputs(26) <= (layer1_outputs(8152)) and not (layer1_outputs(4698));
    layer2_outputs(27) <= not(layer1_outputs(574));
    layer2_outputs(28) <= not((layer1_outputs(3549)) and (layer1_outputs(4258)));
    layer2_outputs(29) <= (layer1_outputs(848)) and not (layer1_outputs(9906));
    layer2_outputs(30) <= not((layer1_outputs(8253)) and (layer1_outputs(8229)));
    layer2_outputs(31) <= (layer1_outputs(4801)) and (layer1_outputs(3280));
    layer2_outputs(32) <= (layer1_outputs(3597)) and not (layer1_outputs(1618));
    layer2_outputs(33) <= not(layer1_outputs(2566));
    layer2_outputs(34) <= '0';
    layer2_outputs(35) <= not(layer1_outputs(4674)) or (layer1_outputs(9016));
    layer2_outputs(36) <= (layer1_outputs(4656)) or (layer1_outputs(6943));
    layer2_outputs(37) <= not(layer1_outputs(4432)) or (layer1_outputs(5095));
    layer2_outputs(38) <= not(layer1_outputs(777));
    layer2_outputs(39) <= (layer1_outputs(127)) and not (layer1_outputs(3254));
    layer2_outputs(40) <= not(layer1_outputs(4710));
    layer2_outputs(41) <= not((layer1_outputs(9413)) or (layer1_outputs(8511)));
    layer2_outputs(42) <= not(layer1_outputs(1583)) or (layer1_outputs(102));
    layer2_outputs(43) <= layer1_outputs(1102);
    layer2_outputs(44) <= not(layer1_outputs(4229));
    layer2_outputs(45) <= not((layer1_outputs(10186)) or (layer1_outputs(8353)));
    layer2_outputs(46) <= not(layer1_outputs(3559));
    layer2_outputs(47) <= not((layer1_outputs(5130)) xor (layer1_outputs(8501)));
    layer2_outputs(48) <= not(layer1_outputs(8062));
    layer2_outputs(49) <= not(layer1_outputs(7259));
    layer2_outputs(50) <= '1';
    layer2_outputs(51) <= layer1_outputs(9362);
    layer2_outputs(52) <= (layer1_outputs(2755)) and not (layer1_outputs(6152));
    layer2_outputs(53) <= not(layer1_outputs(7967));
    layer2_outputs(54) <= '0';
    layer2_outputs(55) <= layer1_outputs(8595);
    layer2_outputs(56) <= layer1_outputs(7123);
    layer2_outputs(57) <= layer1_outputs(3811);
    layer2_outputs(58) <= '0';
    layer2_outputs(59) <= not(layer1_outputs(2838));
    layer2_outputs(60) <= not(layer1_outputs(1698));
    layer2_outputs(61) <= '0';
    layer2_outputs(62) <= not(layer1_outputs(9645)) or (layer1_outputs(460));
    layer2_outputs(63) <= not((layer1_outputs(1773)) xor (layer1_outputs(368)));
    layer2_outputs(64) <= not(layer1_outputs(6194)) or (layer1_outputs(6684));
    layer2_outputs(65) <= (layer1_outputs(7815)) and not (layer1_outputs(8165));
    layer2_outputs(66) <= not(layer1_outputs(7348));
    layer2_outputs(67) <= layer1_outputs(7958);
    layer2_outputs(68) <= (layer1_outputs(5445)) and (layer1_outputs(2038));
    layer2_outputs(69) <= not(layer1_outputs(5687));
    layer2_outputs(70) <= not((layer1_outputs(828)) and (layer1_outputs(2375)));
    layer2_outputs(71) <= (layer1_outputs(2146)) and (layer1_outputs(1272));
    layer2_outputs(72) <= layer1_outputs(433);
    layer2_outputs(73) <= not(layer1_outputs(6393));
    layer2_outputs(74) <= layer1_outputs(9219);
    layer2_outputs(75) <= not(layer1_outputs(3513)) or (layer1_outputs(1172));
    layer2_outputs(76) <= (layer1_outputs(8429)) or (layer1_outputs(2557));
    layer2_outputs(77) <= (layer1_outputs(2592)) and not (layer1_outputs(9980));
    layer2_outputs(78) <= not((layer1_outputs(373)) and (layer1_outputs(5873)));
    layer2_outputs(79) <= (layer1_outputs(1419)) or (layer1_outputs(4778));
    layer2_outputs(80) <= layer1_outputs(6429);
    layer2_outputs(81) <= not(layer1_outputs(4598));
    layer2_outputs(82) <= not(layer1_outputs(2798));
    layer2_outputs(83) <= layer1_outputs(2128);
    layer2_outputs(84) <= not(layer1_outputs(3284)) or (layer1_outputs(8251));
    layer2_outputs(85) <= (layer1_outputs(7040)) and not (layer1_outputs(1562));
    layer2_outputs(86) <= layer1_outputs(7738);
    layer2_outputs(87) <= '0';
    layer2_outputs(88) <= layer1_outputs(4908);
    layer2_outputs(89) <= (layer1_outputs(5009)) and not (layer1_outputs(305));
    layer2_outputs(90) <= not(layer1_outputs(7783));
    layer2_outputs(91) <= not(layer1_outputs(4419));
    layer2_outputs(92) <= (layer1_outputs(6680)) and (layer1_outputs(3701));
    layer2_outputs(93) <= not((layer1_outputs(6600)) xor (layer1_outputs(7636)));
    layer2_outputs(94) <= layer1_outputs(7725);
    layer2_outputs(95) <= (layer1_outputs(2702)) or (layer1_outputs(9799));
    layer2_outputs(96) <= (layer1_outputs(7720)) or (layer1_outputs(6038));
    layer2_outputs(97) <= not(layer1_outputs(97));
    layer2_outputs(98) <= (layer1_outputs(5935)) and not (layer1_outputs(4365));
    layer2_outputs(99) <= not(layer1_outputs(1683));
    layer2_outputs(100) <= layer1_outputs(9704);
    layer2_outputs(101) <= layer1_outputs(74);
    layer2_outputs(102) <= (layer1_outputs(3710)) xor (layer1_outputs(1821));
    layer2_outputs(103) <= not(layer1_outputs(3714)) or (layer1_outputs(9890));
    layer2_outputs(104) <= (layer1_outputs(9432)) and not (layer1_outputs(3829));
    layer2_outputs(105) <= layer1_outputs(1811);
    layer2_outputs(106) <= '0';
    layer2_outputs(107) <= (layer1_outputs(7998)) and (layer1_outputs(9119));
    layer2_outputs(108) <= (layer1_outputs(742)) xor (layer1_outputs(11));
    layer2_outputs(109) <= not(layer1_outputs(2595));
    layer2_outputs(110) <= not(layer1_outputs(9287)) or (layer1_outputs(7212));
    layer2_outputs(111) <= not(layer1_outputs(7069)) or (layer1_outputs(2561));
    layer2_outputs(112) <= not((layer1_outputs(3691)) xor (layer1_outputs(1222)));
    layer2_outputs(113) <= not((layer1_outputs(1887)) or (layer1_outputs(3467)));
    layer2_outputs(114) <= layer1_outputs(1149);
    layer2_outputs(115) <= (layer1_outputs(2878)) and not (layer1_outputs(1524));
    layer2_outputs(116) <= not(layer1_outputs(7659));
    layer2_outputs(117) <= not(layer1_outputs(6267));
    layer2_outputs(118) <= layer1_outputs(2196);
    layer2_outputs(119) <= layer1_outputs(7389);
    layer2_outputs(120) <= layer1_outputs(9967);
    layer2_outputs(121) <= not(layer1_outputs(2520)) or (layer1_outputs(621));
    layer2_outputs(122) <= (layer1_outputs(5383)) and (layer1_outputs(6529));
    layer2_outputs(123) <= not(layer1_outputs(3706)) or (layer1_outputs(3968));
    layer2_outputs(124) <= not((layer1_outputs(2721)) or (layer1_outputs(4861)));
    layer2_outputs(125) <= not(layer1_outputs(5652));
    layer2_outputs(126) <= not(layer1_outputs(8248));
    layer2_outputs(127) <= (layer1_outputs(3418)) and not (layer1_outputs(2199));
    layer2_outputs(128) <= not(layer1_outputs(6705));
    layer2_outputs(129) <= layer1_outputs(3952);
    layer2_outputs(130) <= not(layer1_outputs(7827)) or (layer1_outputs(5683));
    layer2_outputs(131) <= not(layer1_outputs(6000));
    layer2_outputs(132) <= not(layer1_outputs(5851));
    layer2_outputs(133) <= not(layer1_outputs(6500));
    layer2_outputs(134) <= (layer1_outputs(1760)) and not (layer1_outputs(1373));
    layer2_outputs(135) <= not(layer1_outputs(5976));
    layer2_outputs(136) <= not((layer1_outputs(5114)) and (layer1_outputs(8099)));
    layer2_outputs(137) <= (layer1_outputs(76)) and (layer1_outputs(6157));
    layer2_outputs(138) <= not(layer1_outputs(8819)) or (layer1_outputs(8790));
    layer2_outputs(139) <= layer1_outputs(8040);
    layer2_outputs(140) <= not((layer1_outputs(8916)) xor (layer1_outputs(3870)));
    layer2_outputs(141) <= (layer1_outputs(7032)) and (layer1_outputs(9495));
    layer2_outputs(142) <= layer1_outputs(7840);
    layer2_outputs(143) <= (layer1_outputs(7205)) xor (layer1_outputs(2440));
    layer2_outputs(144) <= not(layer1_outputs(436));
    layer2_outputs(145) <= '0';
    layer2_outputs(146) <= not(layer1_outputs(4541)) or (layer1_outputs(389));
    layer2_outputs(147) <= not(layer1_outputs(4601));
    layer2_outputs(148) <= layer1_outputs(1453);
    layer2_outputs(149) <= layer1_outputs(1078);
    layer2_outputs(150) <= not(layer1_outputs(1321)) or (layer1_outputs(7681));
    layer2_outputs(151) <= layer1_outputs(6620);
    layer2_outputs(152) <= not(layer1_outputs(9538));
    layer2_outputs(153) <= layer1_outputs(6401);
    layer2_outputs(154) <= not(layer1_outputs(911));
    layer2_outputs(155) <= (layer1_outputs(8367)) and (layer1_outputs(9692));
    layer2_outputs(156) <= not(layer1_outputs(7170));
    layer2_outputs(157) <= not(layer1_outputs(5355));
    layer2_outputs(158) <= not(layer1_outputs(7879)) or (layer1_outputs(8010));
    layer2_outputs(159) <= (layer1_outputs(5240)) and (layer1_outputs(10226));
    layer2_outputs(160) <= layer1_outputs(6317);
    layer2_outputs(161) <= not(layer1_outputs(9576));
    layer2_outputs(162) <= not((layer1_outputs(4923)) and (layer1_outputs(920)));
    layer2_outputs(163) <= not(layer1_outputs(8504));
    layer2_outputs(164) <= layer1_outputs(518);
    layer2_outputs(165) <= layer1_outputs(5408);
    layer2_outputs(166) <= not(layer1_outputs(2289)) or (layer1_outputs(2428));
    layer2_outputs(167) <= (layer1_outputs(3274)) xor (layer1_outputs(5134));
    layer2_outputs(168) <= layer1_outputs(10212);
    layer2_outputs(169) <= not(layer1_outputs(5586));
    layer2_outputs(170) <= not(layer1_outputs(3525));
    layer2_outputs(171) <= not(layer1_outputs(2506)) or (layer1_outputs(7563));
    layer2_outputs(172) <= (layer1_outputs(7325)) xor (layer1_outputs(5465));
    layer2_outputs(173) <= not(layer1_outputs(9)) or (layer1_outputs(6463));
    layer2_outputs(174) <= (layer1_outputs(8265)) xor (layer1_outputs(3637));
    layer2_outputs(175) <= (layer1_outputs(40)) or (layer1_outputs(6127));
    layer2_outputs(176) <= not((layer1_outputs(2901)) xor (layer1_outputs(7270)));
    layer2_outputs(177) <= not((layer1_outputs(9958)) and (layer1_outputs(3611)));
    layer2_outputs(178) <= not((layer1_outputs(4391)) xor (layer1_outputs(1500)));
    layer2_outputs(179) <= not(layer1_outputs(1864));
    layer2_outputs(180) <= not(layer1_outputs(2738));
    layer2_outputs(181) <= layer1_outputs(4523);
    layer2_outputs(182) <= not(layer1_outputs(2994));
    layer2_outputs(183) <= not((layer1_outputs(538)) and (layer1_outputs(566)));
    layer2_outputs(184) <= (layer1_outputs(3011)) xor (layer1_outputs(8034));
    layer2_outputs(185) <= not(layer1_outputs(855));
    layer2_outputs(186) <= '1';
    layer2_outputs(187) <= not(layer1_outputs(694)) or (layer1_outputs(3226));
    layer2_outputs(188) <= not((layer1_outputs(3419)) and (layer1_outputs(9948)));
    layer2_outputs(189) <= not(layer1_outputs(8913));
    layer2_outputs(190) <= (layer1_outputs(4667)) and not (layer1_outputs(10155));
    layer2_outputs(191) <= not(layer1_outputs(5381));
    layer2_outputs(192) <= not(layer1_outputs(3727)) or (layer1_outputs(3208));
    layer2_outputs(193) <= (layer1_outputs(6890)) and not (layer1_outputs(5027));
    layer2_outputs(194) <= not((layer1_outputs(9744)) xor (layer1_outputs(2490)));
    layer2_outputs(195) <= '0';
    layer2_outputs(196) <= not(layer1_outputs(2140));
    layer2_outputs(197) <= not((layer1_outputs(2990)) and (layer1_outputs(2243)));
    layer2_outputs(198) <= layer1_outputs(9834);
    layer2_outputs(199) <= layer1_outputs(3740);
    layer2_outputs(200) <= not(layer1_outputs(980));
    layer2_outputs(201) <= not(layer1_outputs(8707));
    layer2_outputs(202) <= layer1_outputs(9722);
    layer2_outputs(203) <= not(layer1_outputs(8487));
    layer2_outputs(204) <= layer1_outputs(9733);
    layer2_outputs(205) <= not((layer1_outputs(6318)) or (layer1_outputs(1042)));
    layer2_outputs(206) <= (layer1_outputs(5191)) and (layer1_outputs(5658));
    layer2_outputs(207) <= not(layer1_outputs(7801));
    layer2_outputs(208) <= not(layer1_outputs(5737));
    layer2_outputs(209) <= (layer1_outputs(3517)) xor (layer1_outputs(8672));
    layer2_outputs(210) <= '1';
    layer2_outputs(211) <= (layer1_outputs(8211)) and (layer1_outputs(9332));
    layer2_outputs(212) <= not((layer1_outputs(6332)) and (layer1_outputs(1392)));
    layer2_outputs(213) <= not(layer1_outputs(4219));
    layer2_outputs(214) <= (layer1_outputs(3925)) or (layer1_outputs(2437));
    layer2_outputs(215) <= not(layer1_outputs(650));
    layer2_outputs(216) <= not((layer1_outputs(2882)) xor (layer1_outputs(2427)));
    layer2_outputs(217) <= (layer1_outputs(5847)) and not (layer1_outputs(5451));
    layer2_outputs(218) <= not((layer1_outputs(698)) xor (layer1_outputs(7761)));
    layer2_outputs(219) <= not(layer1_outputs(1479));
    layer2_outputs(220) <= layer1_outputs(3270);
    layer2_outputs(221) <= not(layer1_outputs(1457)) or (layer1_outputs(9088));
    layer2_outputs(222) <= not((layer1_outputs(9586)) xor (layer1_outputs(1441)));
    layer2_outputs(223) <= layer1_outputs(9809);
    layer2_outputs(224) <= not((layer1_outputs(10110)) xor (layer1_outputs(3860)));
    layer2_outputs(225) <= not((layer1_outputs(2236)) or (layer1_outputs(6896)));
    layer2_outputs(226) <= (layer1_outputs(9050)) and not (layer1_outputs(9736));
    layer2_outputs(227) <= not(layer1_outputs(5920));
    layer2_outputs(228) <= (layer1_outputs(9844)) and (layer1_outputs(7144));
    layer2_outputs(229) <= layer1_outputs(3233);
    layer2_outputs(230) <= '1';
    layer2_outputs(231) <= not((layer1_outputs(2229)) or (layer1_outputs(10228)));
    layer2_outputs(232) <= (layer1_outputs(3337)) or (layer1_outputs(9671));
    layer2_outputs(233) <= not(layer1_outputs(5500));
    layer2_outputs(234) <= not(layer1_outputs(432));
    layer2_outputs(235) <= layer1_outputs(3404);
    layer2_outputs(236) <= (layer1_outputs(1783)) or (layer1_outputs(6387));
    layer2_outputs(237) <= '0';
    layer2_outputs(238) <= (layer1_outputs(8690)) xor (layer1_outputs(4317));
    layer2_outputs(239) <= not(layer1_outputs(6158)) or (layer1_outputs(8826));
    layer2_outputs(240) <= layer1_outputs(5773);
    layer2_outputs(241) <= '0';
    layer2_outputs(242) <= not((layer1_outputs(2552)) or (layer1_outputs(3185)));
    layer2_outputs(243) <= (layer1_outputs(4299)) and (layer1_outputs(4859));
    layer2_outputs(244) <= layer1_outputs(8216);
    layer2_outputs(245) <= '0';
    layer2_outputs(246) <= layer1_outputs(6230);
    layer2_outputs(247) <= not(layer1_outputs(10040));
    layer2_outputs(248) <= not(layer1_outputs(130));
    layer2_outputs(249) <= (layer1_outputs(3608)) or (layer1_outputs(9037));
    layer2_outputs(250) <= layer1_outputs(2903);
    layer2_outputs(251) <= (layer1_outputs(1904)) xor (layer1_outputs(5073));
    layer2_outputs(252) <= (layer1_outputs(1874)) and not (layer1_outputs(250));
    layer2_outputs(253) <= not(layer1_outputs(4096));
    layer2_outputs(254) <= not(layer1_outputs(4345)) or (layer1_outputs(7734));
    layer2_outputs(255) <= not((layer1_outputs(6699)) or (layer1_outputs(3388)));
    layer2_outputs(256) <= not(layer1_outputs(3675)) or (layer1_outputs(5052));
    layer2_outputs(257) <= layer1_outputs(3497);
    layer2_outputs(258) <= not(layer1_outputs(1323)) or (layer1_outputs(732));
    layer2_outputs(259) <= (layer1_outputs(699)) or (layer1_outputs(3913));
    layer2_outputs(260) <= not((layer1_outputs(5462)) xor (layer1_outputs(9185)));
    layer2_outputs(261) <= (layer1_outputs(9191)) and not (layer1_outputs(2543));
    layer2_outputs(262) <= not(layer1_outputs(3985)) or (layer1_outputs(6420));
    layer2_outputs(263) <= layer1_outputs(4839);
    layer2_outputs(264) <= layer1_outputs(3230);
    layer2_outputs(265) <= layer1_outputs(6285);
    layer2_outputs(266) <= not((layer1_outputs(4606)) or (layer1_outputs(6790)));
    layer2_outputs(267) <= not(layer1_outputs(5993));
    layer2_outputs(268) <= layer1_outputs(6654);
    layer2_outputs(269) <= not(layer1_outputs(8782)) or (layer1_outputs(8478));
    layer2_outputs(270) <= not(layer1_outputs(9204)) or (layer1_outputs(1525));
    layer2_outputs(271) <= not(layer1_outputs(9773)) or (layer1_outputs(5502));
    layer2_outputs(272) <= not(layer1_outputs(561));
    layer2_outputs(273) <= '0';
    layer2_outputs(274) <= layer1_outputs(2269);
    layer2_outputs(275) <= not(layer1_outputs(187));
    layer2_outputs(276) <= layer1_outputs(10150);
    layer2_outputs(277) <= (layer1_outputs(394)) and not (layer1_outputs(3759));
    layer2_outputs(278) <= layer1_outputs(1294);
    layer2_outputs(279) <= layer1_outputs(1449);
    layer2_outputs(280) <= not(layer1_outputs(7934));
    layer2_outputs(281) <= layer1_outputs(2268);
    layer2_outputs(282) <= not(layer1_outputs(10079));
    layer2_outputs(283) <= not(layer1_outputs(7432));
    layer2_outputs(284) <= not((layer1_outputs(9742)) or (layer1_outputs(9825)));
    layer2_outputs(285) <= not((layer1_outputs(10025)) and (layer1_outputs(7238)));
    layer2_outputs(286) <= not(layer1_outputs(9702));
    layer2_outputs(287) <= not(layer1_outputs(5862));
    layer2_outputs(288) <= layer1_outputs(6544);
    layer2_outputs(289) <= not(layer1_outputs(3633));
    layer2_outputs(290) <= (layer1_outputs(1402)) and (layer1_outputs(998));
    layer2_outputs(291) <= layer1_outputs(2545);
    layer2_outputs(292) <= (layer1_outputs(7304)) xor (layer1_outputs(9310));
    layer2_outputs(293) <= not((layer1_outputs(1346)) and (layer1_outputs(1577)));
    layer2_outputs(294) <= layer1_outputs(4158);
    layer2_outputs(295) <= layer1_outputs(4936);
    layer2_outputs(296) <= not(layer1_outputs(10091)) or (layer1_outputs(6231));
    layer2_outputs(297) <= '1';
    layer2_outputs(298) <= not(layer1_outputs(5148));
    layer2_outputs(299) <= (layer1_outputs(6540)) and (layer1_outputs(947));
    layer2_outputs(300) <= not(layer1_outputs(7466)) or (layer1_outputs(5062));
    layer2_outputs(301) <= not(layer1_outputs(6137));
    layer2_outputs(302) <= not(layer1_outputs(9371));
    layer2_outputs(303) <= (layer1_outputs(9763)) xor (layer1_outputs(9605));
    layer2_outputs(304) <= not(layer1_outputs(2185));
    layer2_outputs(305) <= (layer1_outputs(1904)) xor (layer1_outputs(1635));
    layer2_outputs(306) <= (layer1_outputs(7996)) and not (layer1_outputs(652));
    layer2_outputs(307) <= layer1_outputs(4695);
    layer2_outputs(308) <= not((layer1_outputs(1939)) and (layer1_outputs(7579)));
    layer2_outputs(309) <= not((layer1_outputs(1295)) or (layer1_outputs(729)));
    layer2_outputs(310) <= layer1_outputs(9812);
    layer2_outputs(311) <= layer1_outputs(4067);
    layer2_outputs(312) <= layer1_outputs(6921);
    layer2_outputs(313) <= (layer1_outputs(2283)) xor (layer1_outputs(7783));
    layer2_outputs(314) <= layer1_outputs(9897);
    layer2_outputs(315) <= not(layer1_outputs(1169)) or (layer1_outputs(4284));
    layer2_outputs(316) <= not(layer1_outputs(1117)) or (layer1_outputs(7704));
    layer2_outputs(317) <= layer1_outputs(3683);
    layer2_outputs(318) <= (layer1_outputs(2749)) or (layer1_outputs(7605));
    layer2_outputs(319) <= layer1_outputs(2260);
    layer2_outputs(320) <= not((layer1_outputs(8697)) or (layer1_outputs(1544)));
    layer2_outputs(321) <= not(layer1_outputs(8948));
    layer2_outputs(322) <= '1';
    layer2_outputs(323) <= layer1_outputs(6831);
    layer2_outputs(324) <= not(layer1_outputs(683)) or (layer1_outputs(10158));
    layer2_outputs(325) <= not(layer1_outputs(7426)) or (layer1_outputs(9403));
    layer2_outputs(326) <= not(layer1_outputs(3731));
    layer2_outputs(327) <= (layer1_outputs(3951)) and (layer1_outputs(730));
    layer2_outputs(328) <= not((layer1_outputs(5735)) and (layer1_outputs(8743)));
    layer2_outputs(329) <= not(layer1_outputs(2906));
    layer2_outputs(330) <= not(layer1_outputs(9780));
    layer2_outputs(331) <= layer1_outputs(1758);
    layer2_outputs(332) <= not((layer1_outputs(6821)) and (layer1_outputs(965)));
    layer2_outputs(333) <= not((layer1_outputs(8842)) xor (layer1_outputs(1074)));
    layer2_outputs(334) <= layer1_outputs(1925);
    layer2_outputs(335) <= layer1_outputs(201);
    layer2_outputs(336) <= layer1_outputs(8628);
    layer2_outputs(337) <= not(layer1_outputs(5808)) or (layer1_outputs(7660));
    layer2_outputs(338) <= layer1_outputs(7839);
    layer2_outputs(339) <= '0';
    layer2_outputs(340) <= not(layer1_outputs(5286));
    layer2_outputs(341) <= not(layer1_outputs(7895));
    layer2_outputs(342) <= not(layer1_outputs(6488));
    layer2_outputs(343) <= not(layer1_outputs(2158));
    layer2_outputs(344) <= (layer1_outputs(7337)) or (layer1_outputs(6499));
    layer2_outputs(345) <= (layer1_outputs(3749)) or (layer1_outputs(539));
    layer2_outputs(346) <= not(layer1_outputs(6174));
    layer2_outputs(347) <= layer1_outputs(5724);
    layer2_outputs(348) <= not(layer1_outputs(1347)) or (layer1_outputs(1511));
    layer2_outputs(349) <= not((layer1_outputs(783)) and (layer1_outputs(937)));
    layer2_outputs(350) <= layer1_outputs(10007);
    layer2_outputs(351) <= not((layer1_outputs(4658)) and (layer1_outputs(8545)));
    layer2_outputs(352) <= not((layer1_outputs(3617)) or (layer1_outputs(5811)));
    layer2_outputs(353) <= not(layer1_outputs(10091)) or (layer1_outputs(6262));
    layer2_outputs(354) <= not(layer1_outputs(6572));
    layer2_outputs(355) <= not(layer1_outputs(694));
    layer2_outputs(356) <= (layer1_outputs(8328)) and (layer1_outputs(7038));
    layer2_outputs(357) <= not(layer1_outputs(6299));
    layer2_outputs(358) <= not(layer1_outputs(1814));
    layer2_outputs(359) <= layer1_outputs(3522);
    layer2_outputs(360) <= (layer1_outputs(1182)) xor (layer1_outputs(4367));
    layer2_outputs(361) <= not(layer1_outputs(8357)) or (layer1_outputs(3440));
    layer2_outputs(362) <= (layer1_outputs(3831)) or (layer1_outputs(7399));
    layer2_outputs(363) <= not(layer1_outputs(6240)) or (layer1_outputs(9806));
    layer2_outputs(364) <= layer1_outputs(4925);
    layer2_outputs(365) <= not(layer1_outputs(4125));
    layer2_outputs(366) <= layer1_outputs(2091);
    layer2_outputs(367) <= not((layer1_outputs(8993)) or (layer1_outputs(5954)));
    layer2_outputs(368) <= layer1_outputs(7722);
    layer2_outputs(369) <= not(layer1_outputs(6403));
    layer2_outputs(370) <= (layer1_outputs(3202)) and (layer1_outputs(8167));
    layer2_outputs(371) <= (layer1_outputs(2847)) and (layer1_outputs(8171));
    layer2_outputs(372) <= (layer1_outputs(5230)) and (layer1_outputs(9328));
    layer2_outputs(373) <= not(layer1_outputs(10037)) or (layer1_outputs(7114));
    layer2_outputs(374) <= not(layer1_outputs(1579));
    layer2_outputs(375) <= not(layer1_outputs(8442));
    layer2_outputs(376) <= layer1_outputs(7794);
    layer2_outputs(377) <= layer1_outputs(7941);
    layer2_outputs(378) <= layer1_outputs(7125);
    layer2_outputs(379) <= not((layer1_outputs(3103)) xor (layer1_outputs(5412)));
    layer2_outputs(380) <= (layer1_outputs(5354)) and (layer1_outputs(10031));
    layer2_outputs(381) <= not(layer1_outputs(7491)) or (layer1_outputs(9102));
    layer2_outputs(382) <= not(layer1_outputs(1197)) or (layer1_outputs(3922));
    layer2_outputs(383) <= not((layer1_outputs(1518)) and (layer1_outputs(8768)));
    layer2_outputs(384) <= not(layer1_outputs(8971));
    layer2_outputs(385) <= not((layer1_outputs(3500)) or (layer1_outputs(4280)));
    layer2_outputs(386) <= not(layer1_outputs(2650));
    layer2_outputs(387) <= (layer1_outputs(9090)) and not (layer1_outputs(5043));
    layer2_outputs(388) <= (layer1_outputs(4974)) or (layer1_outputs(1281));
    layer2_outputs(389) <= not((layer1_outputs(5015)) xor (layer1_outputs(6216)));
    layer2_outputs(390) <= not(layer1_outputs(10138));
    layer2_outputs(391) <= (layer1_outputs(3766)) or (layer1_outputs(3643));
    layer2_outputs(392) <= not(layer1_outputs(5126));
    layer2_outputs(393) <= layer1_outputs(4852);
    layer2_outputs(394) <= not((layer1_outputs(5020)) xor (layer1_outputs(9141)));
    layer2_outputs(395) <= (layer1_outputs(7725)) or (layer1_outputs(6139));
    layer2_outputs(396) <= not(layer1_outputs(8229));
    layer2_outputs(397) <= not(layer1_outputs(9209));
    layer2_outputs(398) <= not(layer1_outputs(6099));
    layer2_outputs(399) <= layer1_outputs(7443);
    layer2_outputs(400) <= not((layer1_outputs(653)) or (layer1_outputs(4554)));
    layer2_outputs(401) <= (layer1_outputs(960)) and (layer1_outputs(9666));
    layer2_outputs(402) <= layer1_outputs(4139);
    layer2_outputs(403) <= layer1_outputs(9070);
    layer2_outputs(404) <= not((layer1_outputs(420)) and (layer1_outputs(1992)));
    layer2_outputs(405) <= (layer1_outputs(7404)) and not (layer1_outputs(887));
    layer2_outputs(406) <= not(layer1_outputs(8601)) or (layer1_outputs(3326));
    layer2_outputs(407) <= not(layer1_outputs(9473));
    layer2_outputs(408) <= (layer1_outputs(5394)) and not (layer1_outputs(3292));
    layer2_outputs(409) <= layer1_outputs(2011);
    layer2_outputs(410) <= (layer1_outputs(528)) xor (layer1_outputs(10094));
    layer2_outputs(411) <= not(layer1_outputs(4178));
    layer2_outputs(412) <= (layer1_outputs(9282)) and not (layer1_outputs(7319));
    layer2_outputs(413) <= not((layer1_outputs(5444)) and (layer1_outputs(7919)));
    layer2_outputs(414) <= (layer1_outputs(3654)) and (layer1_outputs(2523));
    layer2_outputs(415) <= not(layer1_outputs(3900)) or (layer1_outputs(1975));
    layer2_outputs(416) <= not(layer1_outputs(9351)) or (layer1_outputs(6493));
    layer2_outputs(417) <= (layer1_outputs(405)) and not (layer1_outputs(7300));
    layer2_outputs(418) <= not((layer1_outputs(7777)) xor (layer1_outputs(5675)));
    layer2_outputs(419) <= '1';
    layer2_outputs(420) <= not((layer1_outputs(8352)) and (layer1_outputs(10126)));
    layer2_outputs(421) <= not(layer1_outputs(3545));
    layer2_outputs(422) <= '1';
    layer2_outputs(423) <= (layer1_outputs(3772)) and not (layer1_outputs(2939));
    layer2_outputs(424) <= not((layer1_outputs(2989)) or (layer1_outputs(5975)));
    layer2_outputs(425) <= not((layer1_outputs(6789)) xor (layer1_outputs(6417)));
    layer2_outputs(426) <= not(layer1_outputs(9136));
    layer2_outputs(427) <= not((layer1_outputs(7597)) or (layer1_outputs(1781)));
    layer2_outputs(428) <= not((layer1_outputs(10024)) xor (layer1_outputs(2635)));
    layer2_outputs(429) <= layer1_outputs(1876);
    layer2_outputs(430) <= '1';
    layer2_outputs(431) <= not(layer1_outputs(8228)) or (layer1_outputs(5526));
    layer2_outputs(432) <= not(layer1_outputs(9479));
    layer2_outputs(433) <= not(layer1_outputs(573));
    layer2_outputs(434) <= '0';
    layer2_outputs(435) <= not(layer1_outputs(5897));
    layer2_outputs(436) <= layer1_outputs(5457);
    layer2_outputs(437) <= (layer1_outputs(8472)) and not (layer1_outputs(1256));
    layer2_outputs(438) <= (layer1_outputs(9354)) and (layer1_outputs(8898));
    layer2_outputs(439) <= (layer1_outputs(4399)) or (layer1_outputs(2565));
    layer2_outputs(440) <= not(layer1_outputs(6883));
    layer2_outputs(441) <= not(layer1_outputs(586));
    layer2_outputs(442) <= not((layer1_outputs(10052)) and (layer1_outputs(6062)));
    layer2_outputs(443) <= (layer1_outputs(3458)) and (layer1_outputs(10118));
    layer2_outputs(444) <= not(layer1_outputs(1624)) or (layer1_outputs(115));
    layer2_outputs(445) <= not((layer1_outputs(523)) and (layer1_outputs(2126)));
    layer2_outputs(446) <= layer1_outputs(686);
    layer2_outputs(447) <= layer1_outputs(9398);
    layer2_outputs(448) <= '0';
    layer2_outputs(449) <= (layer1_outputs(4479)) and not (layer1_outputs(1969));
    layer2_outputs(450) <= not(layer1_outputs(5730)) or (layer1_outputs(1938));
    layer2_outputs(451) <= not((layer1_outputs(9679)) xor (layer1_outputs(4391)));
    layer2_outputs(452) <= not((layer1_outputs(6530)) and (layer1_outputs(1077)));
    layer2_outputs(453) <= not(layer1_outputs(396));
    layer2_outputs(454) <= '0';
    layer2_outputs(455) <= not(layer1_outputs(6555));
    layer2_outputs(456) <= layer1_outputs(4534);
    layer2_outputs(457) <= not((layer1_outputs(955)) xor (layer1_outputs(7661)));
    layer2_outputs(458) <= (layer1_outputs(6247)) and not (layer1_outputs(1411));
    layer2_outputs(459) <= (layer1_outputs(10067)) and not (layer1_outputs(2231));
    layer2_outputs(460) <= layer1_outputs(4154);
    layer2_outputs(461) <= layer1_outputs(8133);
    layer2_outputs(462) <= layer1_outputs(6348);
    layer2_outputs(463) <= (layer1_outputs(2221)) or (layer1_outputs(1986));
    layer2_outputs(464) <= not(layer1_outputs(6826));
    layer2_outputs(465) <= layer1_outputs(503);
    layer2_outputs(466) <= (layer1_outputs(10052)) or (layer1_outputs(1089));
    layer2_outputs(467) <= not(layer1_outputs(6989));
    layer2_outputs(468) <= not((layer1_outputs(5090)) or (layer1_outputs(10026)));
    layer2_outputs(469) <= (layer1_outputs(9644)) or (layer1_outputs(7503));
    layer2_outputs(470) <= not(layer1_outputs(5123));
    layer2_outputs(471) <= layer1_outputs(1652);
    layer2_outputs(472) <= not((layer1_outputs(1946)) or (layer1_outputs(7883)));
    layer2_outputs(473) <= not(layer1_outputs(1776)) or (layer1_outputs(7617));
    layer2_outputs(474) <= not(layer1_outputs(7252)) or (layer1_outputs(8486));
    layer2_outputs(475) <= (layer1_outputs(9001)) xor (layer1_outputs(2460));
    layer2_outputs(476) <= (layer1_outputs(3086)) and (layer1_outputs(5192));
    layer2_outputs(477) <= layer1_outputs(1740);
    layer2_outputs(478) <= not((layer1_outputs(9748)) or (layer1_outputs(9220)));
    layer2_outputs(479) <= not(layer1_outputs(6248)) or (layer1_outputs(6449));
    layer2_outputs(480) <= not((layer1_outputs(3509)) xor (layer1_outputs(8218)));
    layer2_outputs(481) <= not(layer1_outputs(2914));
    layer2_outputs(482) <= (layer1_outputs(4263)) xor (layer1_outputs(7505));
    layer2_outputs(483) <= layer1_outputs(106);
    layer2_outputs(484) <= layer1_outputs(5578);
    layer2_outputs(485) <= not(layer1_outputs(4640));
    layer2_outputs(486) <= (layer1_outputs(5810)) and (layer1_outputs(6034));
    layer2_outputs(487) <= not(layer1_outputs(9590));
    layer2_outputs(488) <= '0';
    layer2_outputs(489) <= not(layer1_outputs(7565));
    layer2_outputs(490) <= (layer1_outputs(4843)) and not (layer1_outputs(4841));
    layer2_outputs(491) <= (layer1_outputs(7822)) or (layer1_outputs(3129));
    layer2_outputs(492) <= not(layer1_outputs(6039));
    layer2_outputs(493) <= not((layer1_outputs(9931)) xor (layer1_outputs(3798)));
    layer2_outputs(494) <= '0';
    layer2_outputs(495) <= layer1_outputs(4136);
    layer2_outputs(496) <= layer1_outputs(1460);
    layer2_outputs(497) <= not(layer1_outputs(9379));
    layer2_outputs(498) <= layer1_outputs(6983);
    layer2_outputs(499) <= (layer1_outputs(7269)) and (layer1_outputs(7736));
    layer2_outputs(500) <= layer1_outputs(3419);
    layer2_outputs(501) <= not((layer1_outputs(2226)) xor (layer1_outputs(874)));
    layer2_outputs(502) <= not(layer1_outputs(1828));
    layer2_outputs(503) <= (layer1_outputs(2060)) and not (layer1_outputs(9543));
    layer2_outputs(504) <= not(layer1_outputs(4420));
    layer2_outputs(505) <= (layer1_outputs(6412)) and not (layer1_outputs(7329));
    layer2_outputs(506) <= (layer1_outputs(4213)) and not (layer1_outputs(1641));
    layer2_outputs(507) <= not(layer1_outputs(2609)) or (layer1_outputs(4302));
    layer2_outputs(508) <= (layer1_outputs(3680)) or (layer1_outputs(5772));
    layer2_outputs(509) <= not(layer1_outputs(5074)) or (layer1_outputs(6416));
    layer2_outputs(510) <= not((layer1_outputs(7024)) and (layer1_outputs(6634)));
    layer2_outputs(511) <= not(layer1_outputs(10135));
    layer2_outputs(512) <= not((layer1_outputs(6030)) xor (layer1_outputs(9879)));
    layer2_outputs(513) <= not((layer1_outputs(10110)) or (layer1_outputs(2426)));
    layer2_outputs(514) <= not(layer1_outputs(5047)) or (layer1_outputs(7219));
    layer2_outputs(515) <= layer1_outputs(10132);
    layer2_outputs(516) <= not(layer1_outputs(2689));
    layer2_outputs(517) <= not((layer1_outputs(889)) and (layer1_outputs(5946)));
    layer2_outputs(518) <= (layer1_outputs(1956)) and not (layer1_outputs(6468));
    layer2_outputs(519) <= '1';
    layer2_outputs(520) <= not((layer1_outputs(2116)) or (layer1_outputs(1920)));
    layer2_outputs(521) <= layer1_outputs(3154);
    layer2_outputs(522) <= '1';
    layer2_outputs(523) <= not(layer1_outputs(7324)) or (layer1_outputs(71));
    layer2_outputs(524) <= '1';
    layer2_outputs(525) <= layer1_outputs(4786);
    layer2_outputs(526) <= layer1_outputs(6757);
    layer2_outputs(527) <= (layer1_outputs(3986)) and not (layer1_outputs(8880));
    layer2_outputs(528) <= not(layer1_outputs(8813));
    layer2_outputs(529) <= not(layer1_outputs(4273));
    layer2_outputs(530) <= not(layer1_outputs(35));
    layer2_outputs(531) <= not(layer1_outputs(6717));
    layer2_outputs(532) <= not(layer1_outputs(1112));
    layer2_outputs(533) <= not(layer1_outputs(8208));
    layer2_outputs(534) <= layer1_outputs(6570);
    layer2_outputs(535) <= not(layer1_outputs(958));
    layer2_outputs(536) <= (layer1_outputs(2408)) and not (layer1_outputs(2980));
    layer2_outputs(537) <= (layer1_outputs(9448)) and (layer1_outputs(3612));
    layer2_outputs(538) <= (layer1_outputs(5165)) and (layer1_outputs(2500));
    layer2_outputs(539) <= not(layer1_outputs(1210));
    layer2_outputs(540) <= not(layer1_outputs(9804));
    layer2_outputs(541) <= not(layer1_outputs(3875));
    layer2_outputs(542) <= layer1_outputs(1985);
    layer2_outputs(543) <= not(layer1_outputs(7833));
    layer2_outputs(544) <= not(layer1_outputs(86)) or (layer1_outputs(4248));
    layer2_outputs(545) <= not((layer1_outputs(1266)) and (layer1_outputs(4032)));
    layer2_outputs(546) <= not(layer1_outputs(804));
    layer2_outputs(547) <= not((layer1_outputs(9038)) or (layer1_outputs(3625)));
    layer2_outputs(548) <= (layer1_outputs(813)) or (layer1_outputs(1566));
    layer2_outputs(549) <= not(layer1_outputs(9757)) or (layer1_outputs(6988));
    layer2_outputs(550) <= not(layer1_outputs(3716));
    layer2_outputs(551) <= not(layer1_outputs(4425));
    layer2_outputs(552) <= not(layer1_outputs(6202));
    layer2_outputs(553) <= not((layer1_outputs(8953)) or (layer1_outputs(1949)));
    layer2_outputs(554) <= not(layer1_outputs(6275)) or (layer1_outputs(9227));
    layer2_outputs(555) <= not(layer1_outputs(9486)) or (layer1_outputs(2531));
    layer2_outputs(556) <= (layer1_outputs(4614)) and (layer1_outputs(10215));
    layer2_outputs(557) <= '1';
    layer2_outputs(558) <= layer1_outputs(9481);
    layer2_outputs(559) <= not((layer1_outputs(5943)) and (layer1_outputs(2865)));
    layer2_outputs(560) <= layer1_outputs(1109);
    layer2_outputs(561) <= not((layer1_outputs(8018)) xor (layer1_outputs(7825)));
    layer2_outputs(562) <= (layer1_outputs(6017)) and not (layer1_outputs(10085));
    layer2_outputs(563) <= not((layer1_outputs(8964)) and (layer1_outputs(9939)));
    layer2_outputs(564) <= layer1_outputs(5786);
    layer2_outputs(565) <= (layer1_outputs(8062)) and (layer1_outputs(5574));
    layer2_outputs(566) <= not(layer1_outputs(6677));
    layer2_outputs(567) <= (layer1_outputs(3055)) and not (layer1_outputs(8073));
    layer2_outputs(568) <= not(layer1_outputs(2389));
    layer2_outputs(569) <= not(layer1_outputs(2675)) or (layer1_outputs(6906));
    layer2_outputs(570) <= not(layer1_outputs(4533));
    layer2_outputs(571) <= (layer1_outputs(10228)) xor (layer1_outputs(115));
    layer2_outputs(572) <= layer1_outputs(3345);
    layer2_outputs(573) <= '1';
    layer2_outputs(574) <= not((layer1_outputs(3294)) and (layer1_outputs(2585)));
    layer2_outputs(575) <= not((layer1_outputs(7677)) or (layer1_outputs(1679)));
    layer2_outputs(576) <= (layer1_outputs(6105)) and (layer1_outputs(2216));
    layer2_outputs(577) <= not(layer1_outputs(1549));
    layer2_outputs(578) <= layer1_outputs(8899);
    layer2_outputs(579) <= layer1_outputs(4538);
    layer2_outputs(580) <= layer1_outputs(3607);
    layer2_outputs(581) <= not(layer1_outputs(3031)) or (layer1_outputs(8780));
    layer2_outputs(582) <= (layer1_outputs(4985)) or (layer1_outputs(2497));
    layer2_outputs(583) <= not(layer1_outputs(4026)) or (layer1_outputs(2057));
    layer2_outputs(584) <= not((layer1_outputs(5101)) xor (layer1_outputs(1397)));
    layer2_outputs(585) <= layer1_outputs(2977);
    layer2_outputs(586) <= (layer1_outputs(8566)) and not (layer1_outputs(4619));
    layer2_outputs(587) <= not(layer1_outputs(8560));
    layer2_outputs(588) <= '1';
    layer2_outputs(589) <= not(layer1_outputs(4581)) or (layer1_outputs(6692));
    layer2_outputs(590) <= not(layer1_outputs(1538));
    layer2_outputs(591) <= layer1_outputs(662);
    layer2_outputs(592) <= '0';
    layer2_outputs(593) <= layer1_outputs(7776);
    layer2_outputs(594) <= not(layer1_outputs(4375));
    layer2_outputs(595) <= not((layer1_outputs(70)) or (layer1_outputs(8774)));
    layer2_outputs(596) <= not(layer1_outputs(6834));
    layer2_outputs(597) <= not(layer1_outputs(5476));
    layer2_outputs(598) <= layer1_outputs(6784);
    layer2_outputs(599) <= layer1_outputs(4189);
    layer2_outputs(600) <= not(layer1_outputs(4490)) or (layer1_outputs(854));
    layer2_outputs(601) <= (layer1_outputs(2958)) and (layer1_outputs(9592));
    layer2_outputs(602) <= not((layer1_outputs(3442)) and (layer1_outputs(4142)));
    layer2_outputs(603) <= (layer1_outputs(967)) or (layer1_outputs(5458));
    layer2_outputs(604) <= not(layer1_outputs(2007)) or (layer1_outputs(1267));
    layer2_outputs(605) <= (layer1_outputs(3547)) and not (layer1_outputs(7153));
    layer2_outputs(606) <= not(layer1_outputs(8838));
    layer2_outputs(607) <= '0';
    layer2_outputs(608) <= (layer1_outputs(2336)) and (layer1_outputs(5279));
    layer2_outputs(609) <= layer1_outputs(1251);
    layer2_outputs(610) <= not(layer1_outputs(7129));
    layer2_outputs(611) <= not(layer1_outputs(2540));
    layer2_outputs(612) <= not(layer1_outputs(8402)) or (layer1_outputs(1530));
    layer2_outputs(613) <= (layer1_outputs(6050)) and not (layer1_outputs(8496));
    layer2_outputs(614) <= not(layer1_outputs(5507));
    layer2_outputs(615) <= (layer1_outputs(2249)) and not (layer1_outputs(2015));
    layer2_outputs(616) <= '0';
    layer2_outputs(617) <= not(layer1_outputs(2669));
    layer2_outputs(618) <= (layer1_outputs(10030)) and not (layer1_outputs(178));
    layer2_outputs(619) <= not(layer1_outputs(6764));
    layer2_outputs(620) <= layer1_outputs(7601);
    layer2_outputs(621) <= (layer1_outputs(650)) xor (layer1_outputs(7528));
    layer2_outputs(622) <= (layer1_outputs(7581)) and (layer1_outputs(4130));
    layer2_outputs(623) <= layer1_outputs(4722);
    layer2_outputs(624) <= (layer1_outputs(10235)) and (layer1_outputs(10191));
    layer2_outputs(625) <= layer1_outputs(4087);
    layer2_outputs(626) <= (layer1_outputs(2839)) xor (layer1_outputs(4940));
    layer2_outputs(627) <= (layer1_outputs(5713)) and (layer1_outputs(3947));
    layer2_outputs(628) <= not((layer1_outputs(233)) and (layer1_outputs(1558)));
    layer2_outputs(629) <= (layer1_outputs(3783)) and not (layer1_outputs(4790));
    layer2_outputs(630) <= not(layer1_outputs(2891));
    layer2_outputs(631) <= (layer1_outputs(1037)) or (layer1_outputs(1797));
    layer2_outputs(632) <= not(layer1_outputs(6159));
    layer2_outputs(633) <= not(layer1_outputs(2402));
    layer2_outputs(634) <= (layer1_outputs(8772)) or (layer1_outputs(4973));
    layer2_outputs(635) <= (layer1_outputs(5525)) and not (layer1_outputs(9444));
    layer2_outputs(636) <= not((layer1_outputs(597)) or (layer1_outputs(9770)));
    layer2_outputs(637) <= not((layer1_outputs(5905)) or (layer1_outputs(500)));
    layer2_outputs(638) <= (layer1_outputs(6074)) and not (layer1_outputs(6533));
    layer2_outputs(639) <= '1';
    layer2_outputs(640) <= layer1_outputs(970);
    layer2_outputs(641) <= (layer1_outputs(2016)) and not (layer1_outputs(3156));
    layer2_outputs(642) <= layer1_outputs(9280);
    layer2_outputs(643) <= not(layer1_outputs(1772));
    layer2_outputs(644) <= (layer1_outputs(3186)) and (layer1_outputs(2972));
    layer2_outputs(645) <= (layer1_outputs(2935)) and (layer1_outputs(4862));
    layer2_outputs(646) <= not(layer1_outputs(1358));
    layer2_outputs(647) <= (layer1_outputs(1176)) xor (layer1_outputs(7248));
    layer2_outputs(648) <= not(layer1_outputs(702));
    layer2_outputs(649) <= layer1_outputs(302);
    layer2_outputs(650) <= (layer1_outputs(5940)) and (layer1_outputs(10101));
    layer2_outputs(651) <= (layer1_outputs(7837)) and (layer1_outputs(3897));
    layer2_outputs(652) <= '0';
    layer2_outputs(653) <= layer1_outputs(378);
    layer2_outputs(654) <= (layer1_outputs(10220)) xor (layer1_outputs(4129));
    layer2_outputs(655) <= '1';
    layer2_outputs(656) <= not((layer1_outputs(7878)) or (layer1_outputs(200)));
    layer2_outputs(657) <= layer1_outputs(5994);
    layer2_outputs(658) <= '0';
    layer2_outputs(659) <= not(layer1_outputs(6895));
    layer2_outputs(660) <= not(layer1_outputs(8159));
    layer2_outputs(661) <= not((layer1_outputs(1908)) and (layer1_outputs(282)));
    layer2_outputs(662) <= not((layer1_outputs(3355)) xor (layer1_outputs(6922)));
    layer2_outputs(663) <= not((layer1_outputs(2240)) or (layer1_outputs(4832)));
    layer2_outputs(664) <= layer1_outputs(5080);
    layer2_outputs(665) <= layer1_outputs(1527);
    layer2_outputs(666) <= (layer1_outputs(9736)) xor (layer1_outputs(3581));
    layer2_outputs(667) <= (layer1_outputs(2691)) xor (layer1_outputs(4474));
    layer2_outputs(668) <= not(layer1_outputs(7444));
    layer2_outputs(669) <= not((layer1_outputs(4538)) and (layer1_outputs(4706)));
    layer2_outputs(670) <= layer1_outputs(693);
    layer2_outputs(671) <= '1';
    layer2_outputs(672) <= not(layer1_outputs(5845));
    layer2_outputs(673) <= (layer1_outputs(3310)) and not (layer1_outputs(1050));
    layer2_outputs(674) <= not(layer1_outputs(6980));
    layer2_outputs(675) <= layer1_outputs(9033);
    layer2_outputs(676) <= not(layer1_outputs(1381)) or (layer1_outputs(2664));
    layer2_outputs(677) <= layer1_outputs(10218);
    layer2_outputs(678) <= not(layer1_outputs(3043)) or (layer1_outputs(9203));
    layer2_outputs(679) <= not(layer1_outputs(8182));
    layer2_outputs(680) <= (layer1_outputs(4521)) xor (layer1_outputs(5699));
    layer2_outputs(681) <= not(layer1_outputs(5370));
    layer2_outputs(682) <= (layer1_outputs(4463)) or (layer1_outputs(9577));
    layer2_outputs(683) <= layer1_outputs(1857);
    layer2_outputs(684) <= not(layer1_outputs(454));
    layer2_outputs(685) <= '0';
    layer2_outputs(686) <= not(layer1_outputs(7289)) or (layer1_outputs(386));
    layer2_outputs(687) <= (layer1_outputs(5028)) or (layer1_outputs(9518));
    layer2_outputs(688) <= not((layer1_outputs(1043)) and (layer1_outputs(441)));
    layer2_outputs(689) <= layer1_outputs(9465);
    layer2_outputs(690) <= layer1_outputs(8465);
    layer2_outputs(691) <= not(layer1_outputs(9890));
    layer2_outputs(692) <= not(layer1_outputs(6425)) or (layer1_outputs(2789));
    layer2_outputs(693) <= layer1_outputs(1343);
    layer2_outputs(694) <= (layer1_outputs(981)) or (layer1_outputs(8378));
    layer2_outputs(695) <= layer1_outputs(3709);
    layer2_outputs(696) <= not((layer1_outputs(8597)) xor (layer1_outputs(2860)));
    layer2_outputs(697) <= '0';
    layer2_outputs(698) <= layer1_outputs(6630);
    layer2_outputs(699) <= not(layer1_outputs(1216)) or (layer1_outputs(3832));
    layer2_outputs(700) <= (layer1_outputs(8021)) or (layer1_outputs(5124));
    layer2_outputs(701) <= not(layer1_outputs(6538)) or (layer1_outputs(3059));
    layer2_outputs(702) <= (layer1_outputs(6596)) and not (layer1_outputs(6343));
    layer2_outputs(703) <= layer1_outputs(963);
    layer2_outputs(704) <= (layer1_outputs(1300)) and not (layer1_outputs(8453));
    layer2_outputs(705) <= (layer1_outputs(7282)) and not (layer1_outputs(9122));
    layer2_outputs(706) <= not(layer1_outputs(5854)) or (layer1_outputs(7729));
    layer2_outputs(707) <= not(layer1_outputs(9538));
    layer2_outputs(708) <= not(layer1_outputs(5330));
    layer2_outputs(709) <= '0';
    layer2_outputs(710) <= '1';
    layer2_outputs(711) <= not(layer1_outputs(1567));
    layer2_outputs(712) <= not((layer1_outputs(7680)) xor (layer1_outputs(1537)));
    layer2_outputs(713) <= not(layer1_outputs(2514));
    layer2_outputs(714) <= not(layer1_outputs(1875));
    layer2_outputs(715) <= layer1_outputs(449);
    layer2_outputs(716) <= layer1_outputs(4145);
    layer2_outputs(717) <= '0';
    layer2_outputs(718) <= not((layer1_outputs(9764)) xor (layer1_outputs(2958)));
    layer2_outputs(719) <= layer1_outputs(567);
    layer2_outputs(720) <= layer1_outputs(7310);
    layer2_outputs(721) <= (layer1_outputs(1805)) and (layer1_outputs(9074));
    layer2_outputs(722) <= not(layer1_outputs(2461));
    layer2_outputs(723) <= (layer1_outputs(7899)) and not (layer1_outputs(4226));
    layer2_outputs(724) <= layer1_outputs(7091);
    layer2_outputs(725) <= not(layer1_outputs(222));
    layer2_outputs(726) <= layer1_outputs(8852);
    layer2_outputs(727) <= not(layer1_outputs(3887)) or (layer1_outputs(6253));
    layer2_outputs(728) <= layer1_outputs(5603);
    layer2_outputs(729) <= layer1_outputs(6229);
    layer2_outputs(730) <= layer1_outputs(3549);
    layer2_outputs(731) <= (layer1_outputs(6635)) and not (layer1_outputs(3454));
    layer2_outputs(732) <= not(layer1_outputs(8803));
    layer2_outputs(733) <= not(layer1_outputs(3429));
    layer2_outputs(734) <= '0';
    layer2_outputs(735) <= not((layer1_outputs(8490)) and (layer1_outputs(9313)));
    layer2_outputs(736) <= layer1_outputs(3818);
    layer2_outputs(737) <= not(layer1_outputs(5196)) or (layer1_outputs(5166));
    layer2_outputs(738) <= not((layer1_outputs(7811)) xor (layer1_outputs(3002)));
    layer2_outputs(739) <= layer1_outputs(6491);
    layer2_outputs(740) <= layer1_outputs(9694);
    layer2_outputs(741) <= not(layer1_outputs(4478));
    layer2_outputs(742) <= '0';
    layer2_outputs(743) <= (layer1_outputs(8566)) and (layer1_outputs(1837));
    layer2_outputs(744) <= (layer1_outputs(1956)) and (layer1_outputs(5024));
    layer2_outputs(745) <= layer1_outputs(3621);
    layer2_outputs(746) <= not((layer1_outputs(3211)) and (layer1_outputs(7851)));
    layer2_outputs(747) <= not(layer1_outputs(2952)) or (layer1_outputs(6548));
    layer2_outputs(748) <= not((layer1_outputs(4050)) and (layer1_outputs(1147)));
    layer2_outputs(749) <= not((layer1_outputs(1969)) and (layer1_outputs(10075)));
    layer2_outputs(750) <= not(layer1_outputs(9066));
    layer2_outputs(751) <= (layer1_outputs(4849)) xor (layer1_outputs(8135));
    layer2_outputs(752) <= not(layer1_outputs(6051));
    layer2_outputs(753) <= '1';
    layer2_outputs(754) <= not((layer1_outputs(6328)) or (layer1_outputs(7977)));
    layer2_outputs(755) <= (layer1_outputs(2150)) and not (layer1_outputs(2387));
    layer2_outputs(756) <= layer1_outputs(951);
    layer2_outputs(757) <= not((layer1_outputs(3889)) and (layer1_outputs(6404)));
    layer2_outputs(758) <= (layer1_outputs(5428)) and not (layer1_outputs(6046));
    layer2_outputs(759) <= '1';
    layer2_outputs(760) <= layer1_outputs(4822);
    layer2_outputs(761) <= layer1_outputs(8103);
    layer2_outputs(762) <= (layer1_outputs(6849)) and not (layer1_outputs(4655));
    layer2_outputs(763) <= (layer1_outputs(6316)) and (layer1_outputs(2776));
    layer2_outputs(764) <= layer1_outputs(1188);
    layer2_outputs(765) <= not((layer1_outputs(401)) xor (layer1_outputs(2568)));
    layer2_outputs(766) <= layer1_outputs(4183);
    layer2_outputs(767) <= not(layer1_outputs(1277));
    layer2_outputs(768) <= (layer1_outputs(3734)) or (layer1_outputs(757));
    layer2_outputs(769) <= '1';
    layer2_outputs(770) <= not((layer1_outputs(2854)) and (layer1_outputs(2613)));
    layer2_outputs(771) <= not(layer1_outputs(8231));
    layer2_outputs(772) <= not((layer1_outputs(961)) or (layer1_outputs(9928)));
    layer2_outputs(773) <= (layer1_outputs(7874)) and not (layer1_outputs(8219));
    layer2_outputs(774) <= not(layer1_outputs(9943)) or (layer1_outputs(3694));
    layer2_outputs(775) <= '1';
    layer2_outputs(776) <= layer1_outputs(8723);
    layer2_outputs(777) <= not(layer1_outputs(1690));
    layer2_outputs(778) <= layer1_outputs(3318);
    layer2_outputs(779) <= not(layer1_outputs(9588));
    layer2_outputs(780) <= layer1_outputs(6586);
    layer2_outputs(781) <= layer1_outputs(4194);
    layer2_outputs(782) <= not(layer1_outputs(1292)) or (layer1_outputs(3668));
    layer2_outputs(783) <= not(layer1_outputs(7662)) or (layer1_outputs(3629));
    layer2_outputs(784) <= '0';
    layer2_outputs(785) <= '1';
    layer2_outputs(786) <= not(layer1_outputs(5514)) or (layer1_outputs(6155));
    layer2_outputs(787) <= layer1_outputs(3191);
    layer2_outputs(788) <= not((layer1_outputs(8804)) or (layer1_outputs(8843)));
    layer2_outputs(789) <= (layer1_outputs(7962)) or (layer1_outputs(6070));
    layer2_outputs(790) <= not(layer1_outputs(4870));
    layer2_outputs(791) <= (layer1_outputs(2743)) or (layer1_outputs(2129));
    layer2_outputs(792) <= layer1_outputs(8617);
    layer2_outputs(793) <= (layer1_outputs(8164)) and not (layer1_outputs(8334));
    layer2_outputs(794) <= not(layer1_outputs(2843)) or (layer1_outputs(149));
    layer2_outputs(795) <= (layer1_outputs(8763)) and not (layer1_outputs(908));
    layer2_outputs(796) <= layer1_outputs(4655);
    layer2_outputs(797) <= (layer1_outputs(7193)) xor (layer1_outputs(9632));
    layer2_outputs(798) <= (layer1_outputs(8157)) xor (layer1_outputs(8249));
    layer2_outputs(799) <= layer1_outputs(8975);
    layer2_outputs(800) <= not(layer1_outputs(7126)) or (layer1_outputs(51));
    layer2_outputs(801) <= (layer1_outputs(6845)) or (layer1_outputs(3668));
    layer2_outputs(802) <= (layer1_outputs(5739)) or (layer1_outputs(6203));
    layer2_outputs(803) <= not(layer1_outputs(8279));
    layer2_outputs(804) <= not(layer1_outputs(8605));
    layer2_outputs(805) <= not((layer1_outputs(9160)) or (layer1_outputs(8102)));
    layer2_outputs(806) <= (layer1_outputs(2299)) xor (layer1_outputs(209));
    layer2_outputs(807) <= (layer1_outputs(4521)) and not (layer1_outputs(9256));
    layer2_outputs(808) <= layer1_outputs(7587);
    layer2_outputs(809) <= '1';
    layer2_outputs(810) <= layer1_outputs(4259);
    layer2_outputs(811) <= not((layer1_outputs(3954)) or (layer1_outputs(1045)));
    layer2_outputs(812) <= layer1_outputs(4404);
    layer2_outputs(813) <= (layer1_outputs(2453)) or (layer1_outputs(4397));
    layer2_outputs(814) <= layer1_outputs(3343);
    layer2_outputs(815) <= (layer1_outputs(5553)) and (layer1_outputs(2160));
    layer2_outputs(816) <= '0';
    layer2_outputs(817) <= not(layer1_outputs(1202));
    layer2_outputs(818) <= (layer1_outputs(7566)) and (layer1_outputs(3131));
    layer2_outputs(819) <= not(layer1_outputs(6562)) or (layer1_outputs(3018));
    layer2_outputs(820) <= '0';
    layer2_outputs(821) <= (layer1_outputs(8375)) and not (layer1_outputs(1129));
    layer2_outputs(822) <= (layer1_outputs(4712)) and (layer1_outputs(5727));
    layer2_outputs(823) <= layer1_outputs(488);
    layer2_outputs(824) <= layer1_outputs(9006);
    layer2_outputs(825) <= not((layer1_outputs(6312)) xor (layer1_outputs(7115)));
    layer2_outputs(826) <= not((layer1_outputs(4054)) xor (layer1_outputs(497)));
    layer2_outputs(827) <= (layer1_outputs(7148)) or (layer1_outputs(6010));
    layer2_outputs(828) <= layer1_outputs(5081);
    layer2_outputs(829) <= layer1_outputs(849);
    layer2_outputs(830) <= layer1_outputs(4379);
    layer2_outputs(831) <= layer1_outputs(6228);
    layer2_outputs(832) <= layer1_outputs(9218);
    layer2_outputs(833) <= not(layer1_outputs(114)) or (layer1_outputs(3742));
    layer2_outputs(834) <= not(layer1_outputs(2926));
    layer2_outputs(835) <= not(layer1_outputs(3455)) or (layer1_outputs(418));
    layer2_outputs(836) <= not(layer1_outputs(5366));
    layer2_outputs(837) <= not(layer1_outputs(6342));
    layer2_outputs(838) <= layer1_outputs(3178);
    layer2_outputs(839) <= layer1_outputs(8783);
    layer2_outputs(840) <= not((layer1_outputs(7322)) xor (layer1_outputs(3601)));
    layer2_outputs(841) <= not(layer1_outputs(9582));
    layer2_outputs(842) <= (layer1_outputs(1810)) xor (layer1_outputs(1565));
    layer2_outputs(843) <= not((layer1_outputs(1405)) and (layer1_outputs(7694)));
    layer2_outputs(844) <= '0';
    layer2_outputs(845) <= not(layer1_outputs(4863));
    layer2_outputs(846) <= '1';
    layer2_outputs(847) <= not(layer1_outputs(1536)) or (layer1_outputs(2856));
    layer2_outputs(848) <= '0';
    layer2_outputs(849) <= not(layer1_outputs(434));
    layer2_outputs(850) <= layer1_outputs(4764);
    layer2_outputs(851) <= not(layer1_outputs(6822));
    layer2_outputs(852) <= not(layer1_outputs(3149)) or (layer1_outputs(2657));
    layer2_outputs(853) <= (layer1_outputs(9640)) and not (layer1_outputs(2629));
    layer2_outputs(854) <= (layer1_outputs(4810)) or (layer1_outputs(790));
    layer2_outputs(855) <= not(layer1_outputs(9332));
    layer2_outputs(856) <= not(layer1_outputs(7746));
    layer2_outputs(857) <= not(layer1_outputs(6947));
    layer2_outputs(858) <= not(layer1_outputs(8730));
    layer2_outputs(859) <= not(layer1_outputs(4454)) or (layer1_outputs(9393));
    layer2_outputs(860) <= not(layer1_outputs(135)) or (layer1_outputs(2412));
    layer2_outputs(861) <= (layer1_outputs(8684)) and not (layer1_outputs(7450));
    layer2_outputs(862) <= (layer1_outputs(1947)) xor (layer1_outputs(4617));
    layer2_outputs(863) <= not(layer1_outputs(9025)) or (layer1_outputs(7864));
    layer2_outputs(864) <= not(layer1_outputs(7573));
    layer2_outputs(865) <= layer1_outputs(4348);
    layer2_outputs(866) <= not(layer1_outputs(3639));
    layer2_outputs(867) <= not((layer1_outputs(7311)) xor (layer1_outputs(2319)));
    layer2_outputs(868) <= not((layer1_outputs(5518)) and (layer1_outputs(9795)));
    layer2_outputs(869) <= (layer1_outputs(5055)) and not (layer1_outputs(5464));
    layer2_outputs(870) <= not(layer1_outputs(96)) or (layer1_outputs(9108));
    layer2_outputs(871) <= not(layer1_outputs(9977));
    layer2_outputs(872) <= (layer1_outputs(1595)) xor (layer1_outputs(1641));
    layer2_outputs(873) <= not(layer1_outputs(5882));
    layer2_outputs(874) <= (layer1_outputs(6267)) and not (layer1_outputs(7498));
    layer2_outputs(875) <= not(layer1_outputs(4515));
    layer2_outputs(876) <= layer1_outputs(5538);
    layer2_outputs(877) <= not(layer1_outputs(2599)) or (layer1_outputs(5480));
    layer2_outputs(878) <= not(layer1_outputs(3648));
    layer2_outputs(879) <= not((layer1_outputs(1592)) or (layer1_outputs(8913)));
    layer2_outputs(880) <= not(layer1_outputs(5753));
    layer2_outputs(881) <= not(layer1_outputs(4789)) or (layer1_outputs(213));
    layer2_outputs(882) <= layer1_outputs(1417);
    layer2_outputs(883) <= not(layer1_outputs(9390));
    layer2_outputs(884) <= (layer1_outputs(2207)) and not (layer1_outputs(2459));
    layer2_outputs(885) <= not(layer1_outputs(4122)) or (layer1_outputs(4289));
    layer2_outputs(886) <= not((layer1_outputs(2439)) and (layer1_outputs(3548)));
    layer2_outputs(887) <= not(layer1_outputs(905));
    layer2_outputs(888) <= layer1_outputs(9474);
    layer2_outputs(889) <= not(layer1_outputs(4273));
    layer2_outputs(890) <= layer1_outputs(4628);
    layer2_outputs(891) <= layer1_outputs(5515);
    layer2_outputs(892) <= not(layer1_outputs(3758));
    layer2_outputs(893) <= not((layer1_outputs(5471)) and (layer1_outputs(5938)));
    layer2_outputs(894) <= not(layer1_outputs(1076));
    layer2_outputs(895) <= layer1_outputs(1432);
    layer2_outputs(896) <= '1';
    layer2_outputs(897) <= layer1_outputs(4051);
    layer2_outputs(898) <= layer1_outputs(8728);
    layer2_outputs(899) <= not((layer1_outputs(6078)) xor (layer1_outputs(7340)));
    layer2_outputs(900) <= (layer1_outputs(1494)) xor (layer1_outputs(2072));
    layer2_outputs(901) <= layer1_outputs(5289);
    layer2_outputs(902) <= not(layer1_outputs(3840));
    layer2_outputs(903) <= not((layer1_outputs(6444)) xor (layer1_outputs(7651)));
    layer2_outputs(904) <= not(layer1_outputs(6383));
    layer2_outputs(905) <= not(layer1_outputs(9058));
    layer2_outputs(906) <= layer1_outputs(5315);
    layer2_outputs(907) <= (layer1_outputs(5472)) and (layer1_outputs(2129));
    layer2_outputs(908) <= (layer1_outputs(5765)) and (layer1_outputs(3212));
    layer2_outputs(909) <= not((layer1_outputs(1262)) or (layer1_outputs(3947)));
    layer2_outputs(910) <= not(layer1_outputs(2600));
    layer2_outputs(911) <= (layer1_outputs(8130)) and (layer1_outputs(2207));
    layer2_outputs(912) <= not((layer1_outputs(4682)) or (layer1_outputs(4291)));
    layer2_outputs(913) <= not((layer1_outputs(5022)) or (layer1_outputs(4931)));
    layer2_outputs(914) <= layer1_outputs(5568);
    layer2_outputs(915) <= not(layer1_outputs(7470));
    layer2_outputs(916) <= not(layer1_outputs(8748)) or (layer1_outputs(10114));
    layer2_outputs(917) <= (layer1_outputs(8851)) and not (layer1_outputs(9613));
    layer2_outputs(918) <= layer1_outputs(9781);
    layer2_outputs(919) <= not((layer1_outputs(3926)) or (layer1_outputs(8125)));
    layer2_outputs(920) <= not((layer1_outputs(42)) or (layer1_outputs(9484)));
    layer2_outputs(921) <= not((layer1_outputs(678)) and (layer1_outputs(8068)));
    layer2_outputs(922) <= layer1_outputs(6362);
    layer2_outputs(923) <= not((layer1_outputs(2585)) and (layer1_outputs(8133)));
    layer2_outputs(924) <= not((layer1_outputs(8160)) xor (layer1_outputs(7756)));
    layer2_outputs(925) <= '0';
    layer2_outputs(926) <= (layer1_outputs(6607)) and not (layer1_outputs(5377));
    layer2_outputs(927) <= (layer1_outputs(5685)) or (layer1_outputs(357));
    layer2_outputs(928) <= not((layer1_outputs(6976)) and (layer1_outputs(9497)));
    layer2_outputs(929) <= layer1_outputs(6794);
    layer2_outputs(930) <= not((layer1_outputs(2961)) and (layer1_outputs(7412)));
    layer2_outputs(931) <= not((layer1_outputs(9233)) and (layer1_outputs(9111)));
    layer2_outputs(932) <= not(layer1_outputs(2791));
    layer2_outputs(933) <= layer1_outputs(4232);
    layer2_outputs(934) <= not(layer1_outputs(5006)) or (layer1_outputs(2105));
    layer2_outputs(935) <= not(layer1_outputs(5708));
    layer2_outputs(936) <= layer1_outputs(4302);
    layer2_outputs(937) <= (layer1_outputs(384)) and (layer1_outputs(2048));
    layer2_outputs(938) <= (layer1_outputs(10181)) xor (layer1_outputs(4711));
    layer2_outputs(939) <= not(layer1_outputs(3909));
    layer2_outputs(940) <= not(layer1_outputs(2957));
    layer2_outputs(941) <= (layer1_outputs(4525)) or (layer1_outputs(3142));
    layer2_outputs(942) <= (layer1_outputs(1677)) and not (layer1_outputs(3205));
    layer2_outputs(943) <= not((layer1_outputs(9699)) xor (layer1_outputs(5752)));
    layer2_outputs(944) <= layer1_outputs(9758);
    layer2_outputs(945) <= not(layer1_outputs(9106));
    layer2_outputs(946) <= (layer1_outputs(7146)) and not (layer1_outputs(1898));
    layer2_outputs(947) <= (layer1_outputs(7189)) and (layer1_outputs(8991));
    layer2_outputs(948) <= not(layer1_outputs(7657)) or (layer1_outputs(3586));
    layer2_outputs(949) <= (layer1_outputs(9037)) or (layer1_outputs(1019));
    layer2_outputs(950) <= not(layer1_outputs(569));
    layer2_outputs(951) <= layer1_outputs(1536);
    layer2_outputs(952) <= not(layer1_outputs(8110)) or (layer1_outputs(1879));
    layer2_outputs(953) <= not((layer1_outputs(4195)) xor (layer1_outputs(6311)));
    layer2_outputs(954) <= (layer1_outputs(4713)) xor (layer1_outputs(5067));
    layer2_outputs(955) <= not(layer1_outputs(1783));
    layer2_outputs(956) <= not(layer1_outputs(348));
    layer2_outputs(957) <= (layer1_outputs(236)) or (layer1_outputs(738));
    layer2_outputs(958) <= not(layer1_outputs(8312));
    layer2_outputs(959) <= '1';
    layer2_outputs(960) <= not(layer1_outputs(7995));
    layer2_outputs(961) <= layer1_outputs(9441);
    layer2_outputs(962) <= not((layer1_outputs(6940)) or (layer1_outputs(5918)));
    layer2_outputs(963) <= not((layer1_outputs(867)) or (layer1_outputs(6881)));
    layer2_outputs(964) <= '0';
    layer2_outputs(965) <= (layer1_outputs(5825)) and (layer1_outputs(1408));
    layer2_outputs(966) <= '1';
    layer2_outputs(967) <= (layer1_outputs(3575)) and not (layer1_outputs(8732));
    layer2_outputs(968) <= not(layer1_outputs(8906));
    layer2_outputs(969) <= (layer1_outputs(10232)) and (layer1_outputs(4262));
    layer2_outputs(970) <= (layer1_outputs(5064)) and not (layer1_outputs(5644));
    layer2_outputs(971) <= not(layer1_outputs(7271)) or (layer1_outputs(229));
    layer2_outputs(972) <= (layer1_outputs(4559)) and not (layer1_outputs(8055));
    layer2_outputs(973) <= (layer1_outputs(1476)) and not (layer1_outputs(9472));
    layer2_outputs(974) <= not(layer1_outputs(8551)) or (layer1_outputs(1023));
    layer2_outputs(975) <= not((layer1_outputs(5401)) xor (layer1_outputs(9506)));
    layer2_outputs(976) <= '1';
    layer2_outputs(977) <= (layer1_outputs(669)) and not (layer1_outputs(2205));
    layer2_outputs(978) <= not(layer1_outputs(5396)) or (layer1_outputs(8450));
    layer2_outputs(979) <= not(layer1_outputs(664));
    layer2_outputs(980) <= layer1_outputs(2479);
    layer2_outputs(981) <= not(layer1_outputs(10217));
    layer2_outputs(982) <= (layer1_outputs(5138)) and (layer1_outputs(5401));
    layer2_outputs(983) <= layer1_outputs(6257);
    layer2_outputs(984) <= not(layer1_outputs(10048));
    layer2_outputs(985) <= '1';
    layer2_outputs(986) <= not(layer1_outputs(2288));
    layer2_outputs(987) <= not(layer1_outputs(8577)) or (layer1_outputs(7616));
    layer2_outputs(988) <= layer1_outputs(2162);
    layer2_outputs(989) <= not(layer1_outputs(7634));
    layer2_outputs(990) <= layer1_outputs(9658);
    layer2_outputs(991) <= not((layer1_outputs(4857)) or (layer1_outputs(9857)));
    layer2_outputs(992) <= not(layer1_outputs(66)) or (layer1_outputs(7203));
    layer2_outputs(993) <= not(layer1_outputs(8729));
    layer2_outputs(994) <= (layer1_outputs(1768)) and not (layer1_outputs(648));
    layer2_outputs(995) <= not(layer1_outputs(6349));
    layer2_outputs(996) <= not(layer1_outputs(2547)) or (layer1_outputs(7165));
    layer2_outputs(997) <= not(layer1_outputs(1035));
    layer2_outputs(998) <= not(layer1_outputs(7906));
    layer2_outputs(999) <= not(layer1_outputs(3520));
    layer2_outputs(1000) <= (layer1_outputs(8351)) or (layer1_outputs(5159));
    layer2_outputs(1001) <= not(layer1_outputs(6973)) or (layer1_outputs(5393));
    layer2_outputs(1002) <= layer1_outputs(1682);
    layer2_outputs(1003) <= not(layer1_outputs(3392)) or (layer1_outputs(3815));
    layer2_outputs(1004) <= (layer1_outputs(5617)) and not (layer1_outputs(6190));
    layer2_outputs(1005) <= layer1_outputs(5430);
    layer2_outputs(1006) <= not((layer1_outputs(6957)) xor (layer1_outputs(6026)));
    layer2_outputs(1007) <= (layer1_outputs(4298)) and not (layer1_outputs(3924));
    layer2_outputs(1008) <= layer1_outputs(6750);
    layer2_outputs(1009) <= layer1_outputs(4237);
    layer2_outputs(1010) <= layer1_outputs(7658);
    layer2_outputs(1011) <= not(layer1_outputs(2740));
    layer2_outputs(1012) <= not(layer1_outputs(6595)) or (layer1_outputs(2272));
    layer2_outputs(1013) <= layer1_outputs(8050);
    layer2_outputs(1014) <= '1';
    layer2_outputs(1015) <= not(layer1_outputs(8086)) or (layer1_outputs(1354));
    layer2_outputs(1016) <= not(layer1_outputs(2054)) or (layer1_outputs(7965));
    layer2_outputs(1017) <= (layer1_outputs(7650)) or (layer1_outputs(6009));
    layer2_outputs(1018) <= not((layer1_outputs(8316)) xor (layer1_outputs(134)));
    layer2_outputs(1019) <= not((layer1_outputs(9842)) and (layer1_outputs(3693)));
    layer2_outputs(1020) <= not(layer1_outputs(6077));
    layer2_outputs(1021) <= layer1_outputs(4534);
    layer2_outputs(1022) <= (layer1_outputs(6891)) or (layer1_outputs(3819));
    layer2_outputs(1023) <= layer1_outputs(3255);
    layer2_outputs(1024) <= not(layer1_outputs(878));
    layer2_outputs(1025) <= (layer1_outputs(9067)) and (layer1_outputs(1559));
    layer2_outputs(1026) <= not(layer1_outputs(6622)) or (layer1_outputs(7991));
    layer2_outputs(1027) <= '1';
    layer2_outputs(1028) <= layer1_outputs(6415);
    layer2_outputs(1029) <= not((layer1_outputs(9411)) and (layer1_outputs(8902)));
    layer2_outputs(1030) <= layer1_outputs(2752);
    layer2_outputs(1031) <= layer1_outputs(4412);
    layer2_outputs(1032) <= (layer1_outputs(1796)) and not (layer1_outputs(2071));
    layer2_outputs(1033) <= not((layer1_outputs(4305)) and (layer1_outputs(3160)));
    layer2_outputs(1034) <= (layer1_outputs(5748)) and not (layer1_outputs(9107));
    layer2_outputs(1035) <= (layer1_outputs(9827)) xor (layer1_outputs(5990));
    layer2_outputs(1036) <= layer1_outputs(6712);
    layer2_outputs(1037) <= layer1_outputs(1878);
    layer2_outputs(1038) <= (layer1_outputs(4199)) or (layer1_outputs(10106));
    layer2_outputs(1039) <= (layer1_outputs(4582)) and (layer1_outputs(1824));
    layer2_outputs(1040) <= not(layer1_outputs(9091));
    layer2_outputs(1041) <= layer1_outputs(7072);
    layer2_outputs(1042) <= not(layer1_outputs(864));
    layer2_outputs(1043) <= layer1_outputs(8985);
    layer2_outputs(1044) <= layer1_outputs(3124);
    layer2_outputs(1045) <= (layer1_outputs(8048)) and not (layer1_outputs(6660));
    layer2_outputs(1046) <= not(layer1_outputs(525)) or (layer1_outputs(4980));
    layer2_outputs(1047) <= not(layer1_outputs(5907));
    layer2_outputs(1048) <= (layer1_outputs(1885)) or (layer1_outputs(8725));
    layer2_outputs(1049) <= (layer1_outputs(3162)) and (layer1_outputs(1446));
    layer2_outputs(1050) <= layer1_outputs(8716);
    layer2_outputs(1051) <= (layer1_outputs(6447)) or (layer1_outputs(3478));
    layer2_outputs(1052) <= (layer1_outputs(3063)) and not (layer1_outputs(9601));
    layer2_outputs(1053) <= not((layer1_outputs(1250)) or (layer1_outputs(238)));
    layer2_outputs(1054) <= (layer1_outputs(6810)) and not (layer1_outputs(4936));
    layer2_outputs(1055) <= (layer1_outputs(10109)) xor (layer1_outputs(2666));
    layer2_outputs(1056) <= not(layer1_outputs(2620));
    layer2_outputs(1057) <= not((layer1_outputs(8222)) xor (layer1_outputs(6199)));
    layer2_outputs(1058) <= layer1_outputs(2796);
    layer2_outputs(1059) <= not(layer1_outputs(220));
    layer2_outputs(1060) <= not((layer1_outputs(3937)) or (layer1_outputs(8043)));
    layer2_outputs(1061) <= not(layer1_outputs(7093)) or (layer1_outputs(7341));
    layer2_outputs(1062) <= not(layer1_outputs(4424)) or (layer1_outputs(6726));
    layer2_outputs(1063) <= not((layer1_outputs(997)) or (layer1_outputs(2416)));
    layer2_outputs(1064) <= not((layer1_outputs(3689)) xor (layer1_outputs(5814)));
    layer2_outputs(1065) <= layer1_outputs(9555);
    layer2_outputs(1066) <= layer1_outputs(3372);
    layer2_outputs(1067) <= layer1_outputs(184);
    layer2_outputs(1068) <= not(layer1_outputs(2493));
    layer2_outputs(1069) <= layer1_outputs(8127);
    layer2_outputs(1070) <= '0';
    layer2_outputs(1071) <= (layer1_outputs(9618)) and (layer1_outputs(6878));
    layer2_outputs(1072) <= not(layer1_outputs(8607));
    layer2_outputs(1073) <= not(layer1_outputs(4368)) or (layer1_outputs(9028));
    layer2_outputs(1074) <= '1';
    layer2_outputs(1075) <= not(layer1_outputs(2159)) or (layer1_outputs(3351));
    layer2_outputs(1076) <= not((layer1_outputs(2353)) or (layer1_outputs(820)));
    layer2_outputs(1077) <= layer1_outputs(2933);
    layer2_outputs(1078) <= layer1_outputs(8835);
    layer2_outputs(1079) <= not(layer1_outputs(5765));
    layer2_outputs(1080) <= (layer1_outputs(613)) xor (layer1_outputs(4764));
    layer2_outputs(1081) <= not(layer1_outputs(1789)) or (layer1_outputs(2005));
    layer2_outputs(1082) <= not(layer1_outputs(5856)) or (layer1_outputs(7951));
    layer2_outputs(1083) <= layer1_outputs(1362);
    layer2_outputs(1084) <= '1';
    layer2_outputs(1085) <= layer1_outputs(501);
    layer2_outputs(1086) <= not(layer1_outputs(9026)) or (layer1_outputs(9437));
    layer2_outputs(1087) <= layer1_outputs(9772);
    layer2_outputs(1088) <= (layer1_outputs(5897)) and not (layer1_outputs(9920));
    layer2_outputs(1089) <= not(layer1_outputs(8245)) or (layer1_outputs(1295));
    layer2_outputs(1090) <= layer1_outputs(9330);
    layer2_outputs(1091) <= layer1_outputs(6194);
    layer2_outputs(1092) <= layer1_outputs(959);
    layer2_outputs(1093) <= not(layer1_outputs(3804));
    layer2_outputs(1094) <= layer1_outputs(9313);
    layer2_outputs(1095) <= not(layer1_outputs(5519));
    layer2_outputs(1096) <= not(layer1_outputs(4295));
    layer2_outputs(1097) <= not(layer1_outputs(3077));
    layer2_outputs(1098) <= '1';
    layer2_outputs(1099) <= (layer1_outputs(3565)) and (layer1_outputs(8250));
    layer2_outputs(1100) <= not(layer1_outputs(9457)) or (layer1_outputs(1707));
    layer2_outputs(1101) <= not(layer1_outputs(6189));
    layer2_outputs(1102) <= '0';
    layer2_outputs(1103) <= layer1_outputs(9412);
    layer2_outputs(1104) <= not(layer1_outputs(5469));
    layer2_outputs(1105) <= not(layer1_outputs(6771)) or (layer1_outputs(851));
    layer2_outputs(1106) <= layer1_outputs(3609);
    layer2_outputs(1107) <= (layer1_outputs(4481)) and not (layer1_outputs(6441));
    layer2_outputs(1108) <= not(layer1_outputs(7483)) or (layer1_outputs(4736));
    layer2_outputs(1109) <= (layer1_outputs(9202)) and not (layer1_outputs(4808));
    layer2_outputs(1110) <= not((layer1_outputs(8536)) or (layer1_outputs(651)));
    layer2_outputs(1111) <= not(layer1_outputs(4807));
    layer2_outputs(1112) <= not(layer1_outputs(236)) or (layer1_outputs(1382));
    layer2_outputs(1113) <= not(layer1_outputs(2266));
    layer2_outputs(1114) <= not(layer1_outputs(607)) or (layer1_outputs(7338));
    layer2_outputs(1115) <= '0';
    layer2_outputs(1116) <= not(layer1_outputs(5391));
    layer2_outputs(1117) <= layer1_outputs(6239);
    layer2_outputs(1118) <= layer1_outputs(3584);
    layer2_outputs(1119) <= (layer1_outputs(8532)) and (layer1_outputs(5847));
    layer2_outputs(1120) <= not((layer1_outputs(3078)) and (layer1_outputs(3556)));
    layer2_outputs(1121) <= not(layer1_outputs(8788));
    layer2_outputs(1122) <= not(layer1_outputs(1465));
    layer2_outputs(1123) <= not((layer1_outputs(8443)) and (layer1_outputs(553)));
    layer2_outputs(1124) <= (layer1_outputs(4917)) and not (layer1_outputs(7458));
    layer2_outputs(1125) <= not(layer1_outputs(6291));
    layer2_outputs(1126) <= (layer1_outputs(8114)) and not (layer1_outputs(6081));
    layer2_outputs(1127) <= layer1_outputs(2429);
    layer2_outputs(1128) <= not(layer1_outputs(5469));
    layer2_outputs(1129) <= not((layer1_outputs(2683)) and (layer1_outputs(9304)));
    layer2_outputs(1130) <= not(layer1_outputs(5753));
    layer2_outputs(1131) <= (layer1_outputs(6109)) and (layer1_outputs(8920));
    layer2_outputs(1132) <= not(layer1_outputs(10022));
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= not((layer1_outputs(2087)) or (layer1_outputs(1592)));
    layer2_outputs(1135) <= not(layer1_outputs(2963));
    layer2_outputs(1136) <= (layer1_outputs(2970)) or (layer1_outputs(9516));
    layer2_outputs(1137) <= not((layer1_outputs(608)) xor (layer1_outputs(5548)));
    layer2_outputs(1138) <= layer1_outputs(8582);
    layer2_outputs(1139) <= not(layer1_outputs(2689));
    layer2_outputs(1140) <= not(layer1_outputs(6524));
    layer2_outputs(1141) <= not((layer1_outputs(271)) xor (layer1_outputs(8579)));
    layer2_outputs(1142) <= layer1_outputs(9963);
    layer2_outputs(1143) <= layer1_outputs(5107);
    layer2_outputs(1144) <= '0';
    layer2_outputs(1145) <= layer1_outputs(6928);
    layer2_outputs(1146) <= '0';
    layer2_outputs(1147) <= (layer1_outputs(9012)) or (layer1_outputs(487));
    layer2_outputs(1148) <= (layer1_outputs(7096)) or (layer1_outputs(8122));
    layer2_outputs(1149) <= (layer1_outputs(7871)) xor (layer1_outputs(5969));
    layer2_outputs(1150) <= not((layer1_outputs(2645)) xor (layer1_outputs(8673)));
    layer2_outputs(1151) <= layer1_outputs(9574);
    layer2_outputs(1152) <= not(layer1_outputs(9294));
    layer2_outputs(1153) <= layer1_outputs(5154);
    layer2_outputs(1154) <= layer1_outputs(1224);
    layer2_outputs(1155) <= not(layer1_outputs(9645)) or (layer1_outputs(8324));
    layer2_outputs(1156) <= (layer1_outputs(4526)) and not (layer1_outputs(8446));
    layer2_outputs(1157) <= (layer1_outputs(5593)) xor (layer1_outputs(2411));
    layer2_outputs(1158) <= '1';
    layer2_outputs(1159) <= (layer1_outputs(6365)) and not (layer1_outputs(4714));
    layer2_outputs(1160) <= layer1_outputs(5996);
    layer2_outputs(1161) <= not(layer1_outputs(2404));
    layer2_outputs(1162) <= (layer1_outputs(4904)) and not (layer1_outputs(4851));
    layer2_outputs(1163) <= (layer1_outputs(5587)) or (layer1_outputs(7806));
    layer2_outputs(1164) <= not(layer1_outputs(17));
    layer2_outputs(1165) <= not((layer1_outputs(6628)) or (layer1_outputs(8592)));
    layer2_outputs(1166) <= layer1_outputs(787);
    layer2_outputs(1167) <= not(layer1_outputs(2684));
    layer2_outputs(1168) <= layer1_outputs(10034);
    layer2_outputs(1169) <= (layer1_outputs(8347)) and not (layer1_outputs(6212));
    layer2_outputs(1170) <= layer1_outputs(2690);
    layer2_outputs(1171) <= layer1_outputs(2049);
    layer2_outputs(1172) <= not((layer1_outputs(5357)) or (layer1_outputs(1411)));
    layer2_outputs(1173) <= (layer1_outputs(9853)) xor (layer1_outputs(4101));
    layer2_outputs(1174) <= layer1_outputs(1530);
    layer2_outputs(1175) <= layer1_outputs(2837);
    layer2_outputs(1176) <= not(layer1_outputs(6029)) or (layer1_outputs(2937));
    layer2_outputs(1177) <= layer1_outputs(4190);
    layer2_outputs(1178) <= layer1_outputs(696);
    layer2_outputs(1179) <= not((layer1_outputs(4477)) xor (layer1_outputs(5001)));
    layer2_outputs(1180) <= not(layer1_outputs(4013));
    layer2_outputs(1181) <= (layer1_outputs(5762)) or (layer1_outputs(8527));
    layer2_outputs(1182) <= not((layer1_outputs(3342)) or (layer1_outputs(6094)));
    layer2_outputs(1183) <= not(layer1_outputs(603));
    layer2_outputs(1184) <= layer1_outputs(2434);
    layer2_outputs(1185) <= layer1_outputs(4175);
    layer2_outputs(1186) <= layer1_outputs(9849);
    layer2_outputs(1187) <= not(layer1_outputs(1594));
    layer2_outputs(1188) <= '0';
    layer2_outputs(1189) <= layer1_outputs(7886);
    layer2_outputs(1190) <= not(layer1_outputs(7065));
    layer2_outputs(1191) <= not(layer1_outputs(9107));
    layer2_outputs(1192) <= not(layer1_outputs(5373));
    layer2_outputs(1193) <= layer1_outputs(7968);
    layer2_outputs(1194) <= not(layer1_outputs(896)) or (layer1_outputs(880));
    layer2_outputs(1195) <= layer1_outputs(3754);
    layer2_outputs(1196) <= (layer1_outputs(4508)) and not (layer1_outputs(1328));
    layer2_outputs(1197) <= not(layer1_outputs(4149));
    layer2_outputs(1198) <= not(layer1_outputs(5726));
    layer2_outputs(1199) <= not(layer1_outputs(5340));
    layer2_outputs(1200) <= not((layer1_outputs(5743)) and (layer1_outputs(406)));
    layer2_outputs(1201) <= layer1_outputs(10088);
    layer2_outputs(1202) <= not(layer1_outputs(6322));
    layer2_outputs(1203) <= not(layer1_outputs(9734));
    layer2_outputs(1204) <= layer1_outputs(8000);
    layer2_outputs(1205) <= layer1_outputs(3114);
    layer2_outputs(1206) <= (layer1_outputs(8616)) xor (layer1_outputs(4071));
    layer2_outputs(1207) <= (layer1_outputs(1477)) or (layer1_outputs(5410));
    layer2_outputs(1208) <= '0';
    layer2_outputs(1209) <= not(layer1_outputs(9087)) or (layer1_outputs(6068));
    layer2_outputs(1210) <= not(layer1_outputs(1420));
    layer2_outputs(1211) <= layer1_outputs(6866);
    layer2_outputs(1212) <= not((layer1_outputs(9355)) or (layer1_outputs(8608)));
    layer2_outputs(1213) <= not(layer1_outputs(10231)) or (layer1_outputs(4098));
    layer2_outputs(1214) <= not(layer1_outputs(1163));
    layer2_outputs(1215) <= not(layer1_outputs(928));
    layer2_outputs(1216) <= not(layer1_outputs(6474)) or (layer1_outputs(6200));
    layer2_outputs(1217) <= layer1_outputs(4156);
    layer2_outputs(1218) <= not(layer1_outputs(4008)) or (layer1_outputs(8760));
    layer2_outputs(1219) <= not(layer1_outputs(805)) or (layer1_outputs(6409));
    layer2_outputs(1220) <= (layer1_outputs(8257)) xor (layer1_outputs(643));
    layer2_outputs(1221) <= layer1_outputs(4356);
    layer2_outputs(1222) <= not((layer1_outputs(7419)) and (layer1_outputs(6967)));
    layer2_outputs(1223) <= not(layer1_outputs(4925));
    layer2_outputs(1224) <= not((layer1_outputs(9913)) and (layer1_outputs(6100)));
    layer2_outputs(1225) <= not(layer1_outputs(5881));
    layer2_outputs(1226) <= (layer1_outputs(8859)) or (layer1_outputs(9200));
    layer2_outputs(1227) <= not(layer1_outputs(8095)) or (layer1_outputs(7405));
    layer2_outputs(1228) <= (layer1_outputs(9756)) and not (layer1_outputs(7490));
    layer2_outputs(1229) <= (layer1_outputs(7033)) or (layer1_outputs(7066));
    layer2_outputs(1230) <= (layer1_outputs(3911)) xor (layer1_outputs(1058));
    layer2_outputs(1231) <= not((layer1_outputs(7313)) xor (layer1_outputs(2278)));
    layer2_outputs(1232) <= not(layer1_outputs(507));
    layer2_outputs(1233) <= not(layer1_outputs(2783));
    layer2_outputs(1234) <= not(layer1_outputs(5412));
    layer2_outputs(1235) <= '0';
    layer2_outputs(1236) <= not((layer1_outputs(6009)) xor (layer1_outputs(619)));
    layer2_outputs(1237) <= '1';
    layer2_outputs(1238) <= (layer1_outputs(1860)) and (layer1_outputs(5198));
    layer2_outputs(1239) <= not((layer1_outputs(4185)) and (layer1_outputs(7627)));
    layer2_outputs(1240) <= (layer1_outputs(1235)) or (layer1_outputs(1569));
    layer2_outputs(1241) <= (layer1_outputs(5870)) or (layer1_outputs(9137));
    layer2_outputs(1242) <= layer1_outputs(6162);
    layer2_outputs(1243) <= layer1_outputs(8909);
    layer2_outputs(1244) <= (layer1_outputs(6632)) xor (layer1_outputs(6931));
    layer2_outputs(1245) <= layer1_outputs(2149);
    layer2_outputs(1246) <= not(layer1_outputs(399));
    layer2_outputs(1247) <= '1';
    layer2_outputs(1248) <= (layer1_outputs(2960)) or (layer1_outputs(389));
    layer2_outputs(1249) <= (layer1_outputs(8969)) and not (layer1_outputs(5658));
    layer2_outputs(1250) <= not(layer1_outputs(3315)) or (layer1_outputs(6990));
    layer2_outputs(1251) <= layer1_outputs(1736);
    layer2_outputs(1252) <= not((layer1_outputs(6984)) xor (layer1_outputs(4196)));
    layer2_outputs(1253) <= not(layer1_outputs(477)) or (layer1_outputs(9062));
    layer2_outputs(1254) <= '0';
    layer2_outputs(1255) <= not(layer1_outputs(6814));
    layer2_outputs(1256) <= layer1_outputs(7485);
    layer2_outputs(1257) <= (layer1_outputs(4300)) and not (layer1_outputs(44));
    layer2_outputs(1258) <= (layer1_outputs(7615)) and not (layer1_outputs(1192));
    layer2_outputs(1259) <= layer1_outputs(5231);
    layer2_outputs(1260) <= (layer1_outputs(6047)) and not (layer1_outputs(10137));
    layer2_outputs(1261) <= not(layer1_outputs(8444));
    layer2_outputs(1262) <= layer1_outputs(1435);
    layer2_outputs(1263) <= not((layer1_outputs(1596)) and (layer1_outputs(3771)));
    layer2_outputs(1264) <= not((layer1_outputs(9280)) and (layer1_outputs(1915)));
    layer2_outputs(1265) <= not(layer1_outputs(3037));
    layer2_outputs(1266) <= not(layer1_outputs(9505));
    layer2_outputs(1267) <= not(layer1_outputs(5052)) or (layer1_outputs(8571));
    layer2_outputs(1268) <= not(layer1_outputs(3637)) or (layer1_outputs(2485));
    layer2_outputs(1269) <= layer1_outputs(5662);
    layer2_outputs(1270) <= not(layer1_outputs(3218));
    layer2_outputs(1271) <= '0';
    layer2_outputs(1272) <= not((layer1_outputs(2218)) xor (layer1_outputs(2470)));
    layer2_outputs(1273) <= not(layer1_outputs(7598));
    layer2_outputs(1274) <= layer1_outputs(1785);
    layer2_outputs(1275) <= layer1_outputs(663);
    layer2_outputs(1276) <= not((layer1_outputs(2665)) or (layer1_outputs(4120)));
    layer2_outputs(1277) <= not(layer1_outputs(6220));
    layer2_outputs(1278) <= layer1_outputs(9375);
    layer2_outputs(1279) <= not(layer1_outputs(7020)) or (layer1_outputs(687));
    layer2_outputs(1280) <= not(layer1_outputs(7732));
    layer2_outputs(1281) <= not(layer1_outputs(10084)) or (layer1_outputs(3526));
    layer2_outputs(1282) <= not(layer1_outputs(8287));
    layer2_outputs(1283) <= not((layer1_outputs(8658)) or (layer1_outputs(4889)));
    layer2_outputs(1284) <= (layer1_outputs(45)) and not (layer1_outputs(9717));
    layer2_outputs(1285) <= (layer1_outputs(3958)) or (layer1_outputs(7643));
    layer2_outputs(1286) <= (layer1_outputs(616)) and (layer1_outputs(4681));
    layer2_outputs(1287) <= (layer1_outputs(6646)) xor (layer1_outputs(5992));
    layer2_outputs(1288) <= not(layer1_outputs(4919)) or (layer1_outputs(1656));
    layer2_outputs(1289) <= not(layer1_outputs(1567));
    layer2_outputs(1290) <= not(layer1_outputs(6003));
    layer2_outputs(1291) <= layer1_outputs(579);
    layer2_outputs(1292) <= not((layer1_outputs(9542)) or (layer1_outputs(10120)));
    layer2_outputs(1293) <= (layer1_outputs(7142)) xor (layer1_outputs(7108));
    layer2_outputs(1294) <= (layer1_outputs(9207)) or (layer1_outputs(1282));
    layer2_outputs(1295) <= not(layer1_outputs(3451)) or (layer1_outputs(4382));
    layer2_outputs(1296) <= not(layer1_outputs(2984));
    layer2_outputs(1297) <= not((layer1_outputs(4357)) or (layer1_outputs(6162)));
    layer2_outputs(1298) <= not(layer1_outputs(6751));
    layer2_outputs(1299) <= not((layer1_outputs(3682)) or (layer1_outputs(3603)));
    layer2_outputs(1300) <= layer1_outputs(3332);
    layer2_outputs(1301) <= not((layer1_outputs(4976)) or (layer1_outputs(3083)));
    layer2_outputs(1302) <= not((layer1_outputs(1829)) xor (layer1_outputs(10087)));
    layer2_outputs(1303) <= '0';
    layer2_outputs(1304) <= (layer1_outputs(633)) and not (layer1_outputs(1285));
    layer2_outputs(1305) <= not((layer1_outputs(2999)) xor (layer1_outputs(10072)));
    layer2_outputs(1306) <= not(layer1_outputs(7144));
    layer2_outputs(1307) <= '1';
    layer2_outputs(1308) <= (layer1_outputs(1215)) and not (layer1_outputs(4343));
    layer2_outputs(1309) <= not(layer1_outputs(4271)) or (layer1_outputs(9766));
    layer2_outputs(1310) <= (layer1_outputs(9115)) and not (layer1_outputs(7462));
    layer2_outputs(1311) <= layer1_outputs(1694);
    layer2_outputs(1312) <= not(layer1_outputs(5405)) or (layer1_outputs(4003));
    layer2_outputs(1313) <= not((layer1_outputs(9872)) and (layer1_outputs(4734)));
    layer2_outputs(1314) <= (layer1_outputs(747)) and not (layer1_outputs(10097));
    layer2_outputs(1315) <= not((layer1_outputs(5839)) or (layer1_outputs(262)));
    layer2_outputs(1316) <= not((layer1_outputs(1348)) xor (layer1_outputs(4377)));
    layer2_outputs(1317) <= not((layer1_outputs(3852)) and (layer1_outputs(4803)));
    layer2_outputs(1318) <= layer1_outputs(4335);
    layer2_outputs(1319) <= (layer1_outputs(3644)) and (layer1_outputs(1450));
    layer2_outputs(1320) <= (layer1_outputs(6579)) or (layer1_outputs(3675));
    layer2_outputs(1321) <= '1';
    layer2_outputs(1322) <= not((layer1_outputs(8686)) and (layer1_outputs(9374)));
    layer2_outputs(1323) <= not((layer1_outputs(6695)) xor (layer1_outputs(3658)));
    layer2_outputs(1324) <= (layer1_outputs(9962)) and not (layer1_outputs(8161));
    layer2_outputs(1325) <= not(layer1_outputs(5670)) or (layer1_outputs(3991));
    layer2_outputs(1326) <= not(layer1_outputs(7451));
    layer2_outputs(1327) <= not((layer1_outputs(8029)) xor (layer1_outputs(3121)));
    layer2_outputs(1328) <= not(layer1_outputs(8861)) or (layer1_outputs(5614));
    layer2_outputs(1329) <= not((layer1_outputs(3609)) or (layer1_outputs(6597)));
    layer2_outputs(1330) <= layer1_outputs(2074);
    layer2_outputs(1331) <= layer1_outputs(5728);
    layer2_outputs(1332) <= layer1_outputs(9234);
    layer2_outputs(1333) <= layer1_outputs(6959);
    layer2_outputs(1334) <= not(layer1_outputs(7379));
    layer2_outputs(1335) <= not(layer1_outputs(8525));
    layer2_outputs(1336) <= not(layer1_outputs(2984));
    layer2_outputs(1337) <= not(layer1_outputs(7506));
    layer2_outputs(1338) <= (layer1_outputs(281)) xor (layer1_outputs(4622));
    layer2_outputs(1339) <= '1';
    layer2_outputs(1340) <= not(layer1_outputs(8004));
    layer2_outputs(1341) <= '0';
    layer2_outputs(1342) <= layer1_outputs(1170);
    layer2_outputs(1343) <= not(layer1_outputs(7766));
    layer2_outputs(1344) <= not(layer1_outputs(5960));
    layer2_outputs(1345) <= not((layer1_outputs(8696)) xor (layer1_outputs(7818)));
    layer2_outputs(1346) <= not(layer1_outputs(2082));
    layer2_outputs(1347) <= layer1_outputs(9841);
    layer2_outputs(1348) <= not(layer1_outputs(8348));
    layer2_outputs(1349) <= not(layer1_outputs(6258));
    layer2_outputs(1350) <= not((layer1_outputs(2487)) and (layer1_outputs(1433)));
    layer2_outputs(1351) <= not(layer1_outputs(7857));
    layer2_outputs(1352) <= (layer1_outputs(1940)) and not (layer1_outputs(3411));
    layer2_outputs(1353) <= not(layer1_outputs(4218)) or (layer1_outputs(4799));
    layer2_outputs(1354) <= layer1_outputs(9865);
    layer2_outputs(1355) <= not(layer1_outputs(9816));
    layer2_outputs(1356) <= (layer1_outputs(5856)) or (layer1_outputs(841));
    layer2_outputs(1357) <= layer1_outputs(9579);
    layer2_outputs(1358) <= not(layer1_outputs(2211));
    layer2_outputs(1359) <= not(layer1_outputs(4460)) or (layer1_outputs(3722));
    layer2_outputs(1360) <= not((layer1_outputs(5998)) or (layer1_outputs(4111)));
    layer2_outputs(1361) <= '1';
    layer2_outputs(1362) <= (layer1_outputs(1222)) and not (layer1_outputs(382));
    layer2_outputs(1363) <= not(layer1_outputs(7857)) or (layer1_outputs(4294));
    layer2_outputs(1364) <= (layer1_outputs(3336)) and not (layer1_outputs(5834));
    layer2_outputs(1365) <= layer1_outputs(4760);
    layer2_outputs(1366) <= not(layer1_outputs(5447));
    layer2_outputs(1367) <= not(layer1_outputs(4119));
    layer2_outputs(1368) <= not(layer1_outputs(7696)) or (layer1_outputs(1700));
    layer2_outputs(1369) <= not((layer1_outputs(9688)) xor (layer1_outputs(3706)));
    layer2_outputs(1370) <= not(layer1_outputs(3827));
    layer2_outputs(1371) <= layer1_outputs(4341);
    layer2_outputs(1372) <= not(layer1_outputs(3355));
    layer2_outputs(1373) <= layer1_outputs(2086);
    layer2_outputs(1374) <= layer1_outputs(4605);
    layer2_outputs(1375) <= (layer1_outputs(5019)) or (layer1_outputs(8232));
    layer2_outputs(1376) <= layer1_outputs(4449);
    layer2_outputs(1377) <= layer1_outputs(2499);
    layer2_outputs(1378) <= (layer1_outputs(9157)) xor (layer1_outputs(2189));
    layer2_outputs(1379) <= not(layer1_outputs(781)) or (layer1_outputs(8932));
    layer2_outputs(1380) <= not(layer1_outputs(9998));
    layer2_outputs(1381) <= (layer1_outputs(1136)) and not (layer1_outputs(8168));
    layer2_outputs(1382) <= not(layer1_outputs(7689));
    layer2_outputs(1383) <= not(layer1_outputs(4516)) or (layer1_outputs(88));
    layer2_outputs(1384) <= not((layer1_outputs(7750)) xor (layer1_outputs(5432)));
    layer2_outputs(1385) <= '1';
    layer2_outputs(1386) <= not(layer1_outputs(6170));
    layer2_outputs(1387) <= not(layer1_outputs(966));
    layer2_outputs(1388) <= not(layer1_outputs(77));
    layer2_outputs(1389) <= (layer1_outputs(8656)) and (layer1_outputs(3227));
    layer2_outputs(1390) <= (layer1_outputs(5890)) or (layer1_outputs(8970));
    layer2_outputs(1391) <= not((layer1_outputs(3910)) and (layer1_outputs(5732)));
    layer2_outputs(1392) <= (layer1_outputs(2513)) and not (layer1_outputs(9447));
    layer2_outputs(1393) <= not(layer1_outputs(9537));
    layer2_outputs(1394) <= not(layer1_outputs(9597));
    layer2_outputs(1395) <= (layer1_outputs(2441)) and (layer1_outputs(5499));
    layer2_outputs(1396) <= (layer1_outputs(8823)) and not (layer1_outputs(2156));
    layer2_outputs(1397) <= not(layer1_outputs(437));
    layer2_outputs(1398) <= layer1_outputs(6356);
    layer2_outputs(1399) <= not((layer1_outputs(2103)) xor (layer1_outputs(9541)));
    layer2_outputs(1400) <= not(layer1_outputs(6245));
    layer2_outputs(1401) <= (layer1_outputs(8262)) or (layer1_outputs(10083));
    layer2_outputs(1402) <= '1';
    layer2_outputs(1403) <= not((layer1_outputs(6464)) or (layer1_outputs(5402)));
    layer2_outputs(1404) <= (layer1_outputs(6576)) and (layer1_outputs(3971));
    layer2_outputs(1405) <= not(layer1_outputs(5126)) or (layer1_outputs(2761));
    layer2_outputs(1406) <= not(layer1_outputs(9124));
    layer2_outputs(1407) <= (layer1_outputs(1903)) or (layer1_outputs(9089));
    layer2_outputs(1408) <= layer1_outputs(7930);
    layer2_outputs(1409) <= layer1_outputs(5227);
    layer2_outputs(1410) <= not(layer1_outputs(6830)) or (layer1_outputs(7407));
    layer2_outputs(1411) <= not(layer1_outputs(1383));
    layer2_outputs(1412) <= layer1_outputs(6876);
    layer2_outputs(1413) <= (layer1_outputs(7875)) or (layer1_outputs(4499));
    layer2_outputs(1414) <= layer1_outputs(9583);
    layer2_outputs(1415) <= '0';
    layer2_outputs(1416) <= '1';
    layer2_outputs(1417) <= not(layer1_outputs(2009));
    layer2_outputs(1418) <= '0';
    layer2_outputs(1419) <= not(layer1_outputs(3992)) or (layer1_outputs(4466));
    layer2_outputs(1420) <= not(layer1_outputs(8873)) or (layer1_outputs(7516));
    layer2_outputs(1421) <= layer1_outputs(8844);
    layer2_outputs(1422) <= '0';
    layer2_outputs(1423) <= (layer1_outputs(3128)) xor (layer1_outputs(3175));
    layer2_outputs(1424) <= not((layer1_outputs(2422)) or (layer1_outputs(8307)));
    layer2_outputs(1425) <= not(layer1_outputs(7392)) or (layer1_outputs(5728));
    layer2_outputs(1426) <= (layer1_outputs(778)) and not (layer1_outputs(8970));
    layer2_outputs(1427) <= (layer1_outputs(9018)) and not (layer1_outputs(3439));
    layer2_outputs(1428) <= layer1_outputs(6853);
    layer2_outputs(1429) <= not((layer1_outputs(7629)) xor (layer1_outputs(9991)));
    layer2_outputs(1430) <= '0';
    layer2_outputs(1431) <= layer1_outputs(5556);
    layer2_outputs(1432) <= (layer1_outputs(2763)) or (layer1_outputs(5656));
    layer2_outputs(1433) <= not(layer1_outputs(2860));
    layer2_outputs(1434) <= (layer1_outputs(8408)) or (layer1_outputs(7997));
    layer2_outputs(1435) <= not(layer1_outputs(9190)) or (layer1_outputs(3263));
    layer2_outputs(1436) <= (layer1_outputs(2545)) or (layer1_outputs(5777));
    layer2_outputs(1437) <= layer1_outputs(6873);
    layer2_outputs(1438) <= not(layer1_outputs(5986));
    layer2_outputs(1439) <= not(layer1_outputs(398)) or (layer1_outputs(654));
    layer2_outputs(1440) <= not((layer1_outputs(7415)) xor (layer1_outputs(9417)));
    layer2_outputs(1441) <= not(layer1_outputs(8197));
    layer2_outputs(1442) <= (layer1_outputs(5295)) and not (layer1_outputs(605));
    layer2_outputs(1443) <= layer1_outputs(2108);
    layer2_outputs(1444) <= '0';
    layer2_outputs(1445) <= not(layer1_outputs(6946));
    layer2_outputs(1446) <= not(layer1_outputs(5418)) or (layer1_outputs(10090));
    layer2_outputs(1447) <= (layer1_outputs(5721)) and not (layer1_outputs(1493));
    layer2_outputs(1448) <= (layer1_outputs(5245)) and (layer1_outputs(8672));
    layer2_outputs(1449) <= layer1_outputs(6693);
    layer2_outputs(1450) <= not(layer1_outputs(1167));
    layer2_outputs(1451) <= not(layer1_outputs(5562)) or (layer1_outputs(5711));
    layer2_outputs(1452) <= (layer1_outputs(8234)) and (layer1_outputs(4361));
    layer2_outputs(1453) <= (layer1_outputs(8552)) xor (layer1_outputs(7445));
    layer2_outputs(1454) <= not(layer1_outputs(1845)) or (layer1_outputs(2166));
    layer2_outputs(1455) <= (layer1_outputs(1663)) and not (layer1_outputs(210));
    layer2_outputs(1456) <= not(layer1_outputs(3554)) or (layer1_outputs(9363));
    layer2_outputs(1457) <= not((layer1_outputs(8834)) and (layer1_outputs(7343)));
    layer2_outputs(1458) <= (layer1_outputs(164)) and (layer1_outputs(9963));
    layer2_outputs(1459) <= not(layer1_outputs(9962));
    layer2_outputs(1460) <= not((layer1_outputs(9569)) and (layer1_outputs(5553)));
    layer2_outputs(1461) <= (layer1_outputs(2277)) and (layer1_outputs(1842));
    layer2_outputs(1462) <= not(layer1_outputs(4473)) or (layer1_outputs(2879));
    layer2_outputs(1463) <= layer1_outputs(4213);
    layer2_outputs(1464) <= not(layer1_outputs(9592));
    layer2_outputs(1465) <= not(layer1_outputs(8538)) or (layer1_outputs(1047));
    layer2_outputs(1466) <= (layer1_outputs(214)) or (layer1_outputs(1979));
    layer2_outputs(1467) <= not((layer1_outputs(290)) and (layer1_outputs(4693)));
    layer2_outputs(1468) <= not(layer1_outputs(3307));
    layer2_outputs(1469) <= not(layer1_outputs(2150));
    layer2_outputs(1470) <= not((layer1_outputs(3686)) and (layer1_outputs(5534)));
    layer2_outputs(1471) <= not(layer1_outputs(1855));
    layer2_outputs(1472) <= not((layer1_outputs(7977)) xor (layer1_outputs(8146)));
    layer2_outputs(1473) <= not((layer1_outputs(9164)) or (layer1_outputs(704)));
    layer2_outputs(1474) <= not(layer1_outputs(5402)) or (layer1_outputs(6154));
    layer2_outputs(1475) <= layer1_outputs(10209);
    layer2_outputs(1476) <= (layer1_outputs(2553)) and not (layer1_outputs(1913));
    layer2_outputs(1477) <= not((layer1_outputs(4021)) and (layer1_outputs(2577)));
    layer2_outputs(1478) <= (layer1_outputs(1469)) or (layer1_outputs(4874));
    layer2_outputs(1479) <= (layer1_outputs(8524)) or (layer1_outputs(5438));
    layer2_outputs(1480) <= (layer1_outputs(4443)) and not (layer1_outputs(3141));
    layer2_outputs(1481) <= not(layer1_outputs(8570));
    layer2_outputs(1482) <= layer1_outputs(3534);
    layer2_outputs(1483) <= not(layer1_outputs(38));
    layer2_outputs(1484) <= not(layer1_outputs(8480)) or (layer1_outputs(4805));
    layer2_outputs(1485) <= (layer1_outputs(3704)) xor (layer1_outputs(575));
    layer2_outputs(1486) <= layer1_outputs(3939);
    layer2_outputs(1487) <= (layer1_outputs(3686)) xor (layer1_outputs(5996));
    layer2_outputs(1488) <= layer1_outputs(9371);
    layer2_outputs(1489) <= not(layer1_outputs(9850));
    layer2_outputs(1490) <= '0';
    layer2_outputs(1491) <= layer1_outputs(5807);
    layer2_outputs(1492) <= layer1_outputs(9061);
    layer2_outputs(1493) <= (layer1_outputs(4864)) and (layer1_outputs(3846));
    layer2_outputs(1494) <= (layer1_outputs(4941)) and not (layer1_outputs(6872));
    layer2_outputs(1495) <= layer1_outputs(9058);
    layer2_outputs(1496) <= '1';
    layer2_outputs(1497) <= (layer1_outputs(4584)) xor (layer1_outputs(5916));
    layer2_outputs(1498) <= not(layer1_outputs(1233));
    layer2_outputs(1499) <= (layer1_outputs(2477)) or (layer1_outputs(2884));
    layer2_outputs(1500) <= (layer1_outputs(6898)) and not (layer1_outputs(4806));
    layer2_outputs(1501) <= not(layer1_outputs(5015)) or (layer1_outputs(5737));
    layer2_outputs(1502) <= '0';
    layer2_outputs(1503) <= layer1_outputs(9570);
    layer2_outputs(1504) <= (layer1_outputs(9641)) and (layer1_outputs(6323));
    layer2_outputs(1505) <= '1';
    layer2_outputs(1506) <= (layer1_outputs(5163)) and not (layer1_outputs(3058));
    layer2_outputs(1507) <= (layer1_outputs(9960)) and not (layer1_outputs(8706));
    layer2_outputs(1508) <= layer1_outputs(4532);
    layer2_outputs(1509) <= not(layer1_outputs(7209));
    layer2_outputs(1510) <= (layer1_outputs(4163)) and not (layer1_outputs(3380));
    layer2_outputs(1511) <= not((layer1_outputs(8559)) or (layer1_outputs(4070)));
    layer2_outputs(1512) <= not(layer1_outputs(1646));
    layer2_outputs(1513) <= not((layer1_outputs(4621)) and (layer1_outputs(8202)));
    layer2_outputs(1514) <= not(layer1_outputs(1491));
    layer2_outputs(1515) <= not(layer1_outputs(1376));
    layer2_outputs(1516) <= layer1_outputs(2420);
    layer2_outputs(1517) <= not((layer1_outputs(1469)) or (layer1_outputs(7274)));
    layer2_outputs(1518) <= not(layer1_outputs(7816)) or (layer1_outputs(7708));
    layer2_outputs(1519) <= not(layer1_outputs(1902));
    layer2_outputs(1520) <= (layer1_outputs(1664)) and not (layer1_outputs(9674));
    layer2_outputs(1521) <= (layer1_outputs(8534)) and not (layer1_outputs(1486));
    layer2_outputs(1522) <= (layer1_outputs(3375)) or (layer1_outputs(6164));
    layer2_outputs(1523) <= (layer1_outputs(7786)) and (layer1_outputs(4819));
    layer2_outputs(1524) <= (layer1_outputs(6234)) and not (layer1_outputs(3751));
    layer2_outputs(1525) <= layer1_outputs(9760);
    layer2_outputs(1526) <= not(layer1_outputs(9201));
    layer2_outputs(1527) <= layer1_outputs(7104);
    layer2_outputs(1528) <= '0';
    layer2_outputs(1529) <= (layer1_outputs(8265)) or (layer1_outputs(6249));
    layer2_outputs(1530) <= not(layer1_outputs(6314)) or (layer1_outputs(9629));
    layer2_outputs(1531) <= not((layer1_outputs(3126)) xor (layer1_outputs(7562)));
    layer2_outputs(1532) <= not((layer1_outputs(247)) and (layer1_outputs(8720)));
    layer2_outputs(1533) <= not(layer1_outputs(9693));
    layer2_outputs(1534) <= (layer1_outputs(5964)) xor (layer1_outputs(914));
    layer2_outputs(1535) <= layer1_outputs(3696);
    layer2_outputs(1536) <= (layer1_outputs(117)) and not (layer1_outputs(4169));
    layer2_outputs(1537) <= not(layer1_outputs(360));
    layer2_outputs(1538) <= not(layer1_outputs(7219));
    layer2_outputs(1539) <= (layer1_outputs(943)) and not (layer1_outputs(9608));
    layer2_outputs(1540) <= (layer1_outputs(3632)) and not (layer1_outputs(830));
    layer2_outputs(1541) <= '0';
    layer2_outputs(1542) <= '1';
    layer2_outputs(1543) <= not(layer1_outputs(5306));
    layer2_outputs(1544) <= layer1_outputs(5170);
    layer2_outputs(1545) <= not((layer1_outputs(3395)) xor (layer1_outputs(950)));
    layer2_outputs(1546) <= not((layer1_outputs(6168)) and (layer1_outputs(2499)));
    layer2_outputs(1547) <= layer1_outputs(9178);
    layer2_outputs(1548) <= not(layer1_outputs(5010));
    layer2_outputs(1549) <= not(layer1_outputs(9049)) or (layer1_outputs(1905));
    layer2_outputs(1550) <= '0';
    layer2_outputs(1551) <= not(layer1_outputs(6936));
    layer2_outputs(1552) <= (layer1_outputs(1437)) and not (layer1_outputs(7473));
    layer2_outputs(1553) <= layer1_outputs(3546);
    layer2_outputs(1554) <= not(layer1_outputs(824));
    layer2_outputs(1555) <= '0';
    layer2_outputs(1556) <= '0';
    layer2_outputs(1557) <= not(layer1_outputs(5828));
    layer2_outputs(1558) <= layer1_outputs(9370);
    layer2_outputs(1559) <= layer1_outputs(5274);
    layer2_outputs(1560) <= (layer1_outputs(10229)) and not (layer1_outputs(6553));
    layer2_outputs(1561) <= layer1_outputs(4998);
    layer2_outputs(1562) <= not((layer1_outputs(3098)) xor (layer1_outputs(7265)));
    layer2_outputs(1563) <= (layer1_outputs(8844)) or (layer1_outputs(7226));
    layer2_outputs(1564) <= not((layer1_outputs(8190)) or (layer1_outputs(8264)));
    layer2_outputs(1565) <= (layer1_outputs(1971)) and (layer1_outputs(10029));
    layer2_outputs(1566) <= layer1_outputs(6616);
    layer2_outputs(1567) <= not((layer1_outputs(4186)) or (layer1_outputs(5764)));
    layer2_outputs(1568) <= '1';
    layer2_outputs(1569) <= not((layer1_outputs(1029)) or (layer1_outputs(7735)));
    layer2_outputs(1570) <= not(layer1_outputs(792)) or (layer1_outputs(8560));
    layer2_outputs(1571) <= layer1_outputs(4345);
    layer2_outputs(1572) <= (layer1_outputs(1080)) and not (layer1_outputs(7237));
    layer2_outputs(1573) <= not(layer1_outputs(2935));
    layer2_outputs(1574) <= (layer1_outputs(5908)) or (layer1_outputs(6468));
    layer2_outputs(1575) <= not((layer1_outputs(4752)) or (layer1_outputs(4542)));
    layer2_outputs(1576) <= not(layer1_outputs(10051)) or (layer1_outputs(1715));
    layer2_outputs(1577) <= (layer1_outputs(4723)) and (layer1_outputs(8016));
    layer2_outputs(1578) <= layer1_outputs(4039);
    layer2_outputs(1579) <= (layer1_outputs(2120)) and not (layer1_outputs(8309));
    layer2_outputs(1580) <= layer1_outputs(7812);
    layer2_outputs(1581) <= not((layer1_outputs(7044)) or (layer1_outputs(5956)));
    layer2_outputs(1582) <= not(layer1_outputs(3362));
    layer2_outputs(1583) <= layer1_outputs(9347);
    layer2_outputs(1584) <= not((layer1_outputs(2370)) xor (layer1_outputs(854)));
    layer2_outputs(1585) <= not((layer1_outputs(6182)) and (layer1_outputs(8340)));
    layer2_outputs(1586) <= not(layer1_outputs(5977)) or (layer1_outputs(8287));
    layer2_outputs(1587) <= not(layer1_outputs(3638));
    layer2_outputs(1588) <= layer1_outputs(4512);
    layer2_outputs(1589) <= (layer1_outputs(9334)) and (layer1_outputs(3620));
    layer2_outputs(1590) <= not(layer1_outputs(4284)) or (layer1_outputs(6986));
    layer2_outputs(1591) <= '1';
    layer2_outputs(1592) <= (layer1_outputs(1905)) and (layer1_outputs(9801));
    layer2_outputs(1593) <= (layer1_outputs(5341)) and not (layer1_outputs(7415));
    layer2_outputs(1594) <= (layer1_outputs(7603)) and (layer1_outputs(1899));
    layer2_outputs(1595) <= not((layer1_outputs(9845)) xor (layer1_outputs(2168)));
    layer2_outputs(1596) <= not(layer1_outputs(6855));
    layer2_outputs(1597) <= not(layer1_outputs(9413)) or (layer1_outputs(9869));
    layer2_outputs(1598) <= not((layer1_outputs(8473)) or (layer1_outputs(9798)));
    layer2_outputs(1599) <= not(layer1_outputs(554));
    layer2_outputs(1600) <= not(layer1_outputs(4356));
    layer2_outputs(1601) <= not(layer1_outputs(170)) or (layer1_outputs(2005));
    layer2_outputs(1602) <= (layer1_outputs(7711)) and not (layer1_outputs(4037));
    layer2_outputs(1603) <= not(layer1_outputs(3561)) or (layer1_outputs(7276));
    layer2_outputs(1604) <= not(layer1_outputs(8882));
    layer2_outputs(1605) <= '0';
    layer2_outputs(1606) <= '0';
    layer2_outputs(1607) <= layer1_outputs(3705);
    layer2_outputs(1608) <= not(layer1_outputs(8883));
    layer2_outputs(1609) <= not((layer1_outputs(8143)) xor (layer1_outputs(8790)));
    layer2_outputs(1610) <= not(layer1_outputs(7787));
    layer2_outputs(1611) <= (layer1_outputs(4292)) and not (layer1_outputs(3029));
    layer2_outputs(1612) <= '1';
    layer2_outputs(1613) <= not(layer1_outputs(6805));
    layer2_outputs(1614) <= not(layer1_outputs(6331));
    layer2_outputs(1615) <= layer1_outputs(1353);
    layer2_outputs(1616) <= (layer1_outputs(5452)) or (layer1_outputs(1919));
    layer2_outputs(1617) <= not(layer1_outputs(2457)) or (layer1_outputs(6640));
    layer2_outputs(1618) <= '1';
    layer2_outputs(1619) <= not((layer1_outputs(6305)) xor (layer1_outputs(174)));
    layer2_outputs(1620) <= (layer1_outputs(9706)) and (layer1_outputs(8971));
    layer2_outputs(1621) <= not(layer1_outputs(8448)) or (layer1_outputs(3127));
    layer2_outputs(1622) <= not(layer1_outputs(9137));
    layer2_outputs(1623) <= layer1_outputs(7004);
    layer2_outputs(1624) <= not(layer1_outputs(10145));
    layer2_outputs(1625) <= layer1_outputs(9114);
    layer2_outputs(1626) <= not(layer1_outputs(6431));
    layer2_outputs(1627) <= (layer1_outputs(9776)) and not (layer1_outputs(2772));
    layer2_outputs(1628) <= not(layer1_outputs(3857)) or (layer1_outputs(3012));
    layer2_outputs(1629) <= not((layer1_outputs(6290)) xor (layer1_outputs(9566)));
    layer2_outputs(1630) <= (layer1_outputs(159)) and (layer1_outputs(4690));
    layer2_outputs(1631) <= not((layer1_outputs(2309)) xor (layer1_outputs(1990)));
    layer2_outputs(1632) <= not(layer1_outputs(2786));
    layer2_outputs(1633) <= '0';
    layer2_outputs(1634) <= '0';
    layer2_outputs(1635) <= not(layer1_outputs(5253));
    layer2_outputs(1636) <= layer1_outputs(6708);
    layer2_outputs(1637) <= (layer1_outputs(9902)) and not (layer1_outputs(6899));
    layer2_outputs(1638) <= not(layer1_outputs(1760));
    layer2_outputs(1639) <= layer1_outputs(4985);
    layer2_outputs(1640) <= (layer1_outputs(9373)) or (layer1_outputs(3230));
    layer2_outputs(1641) <= layer1_outputs(6284);
    layer2_outputs(1642) <= (layer1_outputs(5924)) or (layer1_outputs(5413));
    layer2_outputs(1643) <= not((layer1_outputs(3471)) or (layer1_outputs(10093)));
    layer2_outputs(1644) <= '0';
    layer2_outputs(1645) <= (layer1_outputs(3466)) and not (layer1_outputs(1040));
    layer2_outputs(1646) <= not(layer1_outputs(4753));
    layer2_outputs(1647) <= not(layer1_outputs(6475));
    layer2_outputs(1648) <= (layer1_outputs(3774)) and not (layer1_outputs(611));
    layer2_outputs(1649) <= not(layer1_outputs(10182));
    layer2_outputs(1650) <= (layer1_outputs(9861)) or (layer1_outputs(3762));
    layer2_outputs(1651) <= '1';
    layer2_outputs(1652) <= (layer1_outputs(6498)) or (layer1_outputs(5962));
    layer2_outputs(1653) <= not((layer1_outputs(5496)) and (layer1_outputs(6121)));
    layer2_outputs(1654) <= not(layer1_outputs(9639));
    layer2_outputs(1655) <= '0';
    layer2_outputs(1656) <= not(layer1_outputs(8448));
    layer2_outputs(1657) <= layer1_outputs(6626);
    layer2_outputs(1658) <= not(layer1_outputs(167)) or (layer1_outputs(1200));
    layer2_outputs(1659) <= '0';
    layer2_outputs(1660) <= not((layer1_outputs(3082)) and (layer1_outputs(4505)));
    layer2_outputs(1661) <= not((layer1_outputs(4027)) xor (layer1_outputs(5618)));
    layer2_outputs(1662) <= (layer1_outputs(4798)) and (layer1_outputs(1095));
    layer2_outputs(1663) <= layer1_outputs(8753);
    layer2_outputs(1664) <= not(layer1_outputs(5290));
    layer2_outputs(1665) <= not((layer1_outputs(3180)) xor (layer1_outputs(7356)));
    layer2_outputs(1666) <= not(layer1_outputs(7742));
    layer2_outputs(1667) <= layer1_outputs(8749);
    layer2_outputs(1668) <= not(layer1_outputs(3946));
    layer2_outputs(1669) <= not(layer1_outputs(861)) or (layer1_outputs(916));
    layer2_outputs(1670) <= not(layer1_outputs(6564));
    layer2_outputs(1671) <= layer1_outputs(7337);
    layer2_outputs(1672) <= not((layer1_outputs(6691)) and (layer1_outputs(7355)));
    layer2_outputs(1673) <= '1';
    layer2_outputs(1674) <= layer1_outputs(6965);
    layer2_outputs(1675) <= not(layer1_outputs(6721));
    layer2_outputs(1676) <= layer1_outputs(4387);
    layer2_outputs(1677) <= layer1_outputs(8028);
    layer2_outputs(1678) <= layer1_outputs(1193);
    layer2_outputs(1679) <= not(layer1_outputs(2919));
    layer2_outputs(1680) <= not(layer1_outputs(6466)) or (layer1_outputs(1244));
    layer2_outputs(1681) <= not((layer1_outputs(9910)) or (layer1_outputs(4662)));
    layer2_outputs(1682) <= layer1_outputs(7860);
    layer2_outputs(1683) <= not(layer1_outputs(201));
    layer2_outputs(1684) <= layer1_outputs(8393);
    layer2_outputs(1685) <= not(layer1_outputs(109));
    layer2_outputs(1686) <= not((layer1_outputs(9581)) and (layer1_outputs(1007)));
    layer2_outputs(1687) <= (layer1_outputs(3810)) or (layer1_outputs(4774));
    layer2_outputs(1688) <= (layer1_outputs(7314)) and not (layer1_outputs(5880));
    layer2_outputs(1689) <= not(layer1_outputs(8424));
    layer2_outputs(1690) <= layer1_outputs(733);
    layer2_outputs(1691) <= not((layer1_outputs(4663)) xor (layer1_outputs(8345)));
    layer2_outputs(1692) <= not(layer1_outputs(2626)) or (layer1_outputs(8754));
    layer2_outputs(1693) <= (layer1_outputs(2167)) or (layer1_outputs(4483));
    layer2_outputs(1694) <= not((layer1_outputs(9551)) or (layer1_outputs(9578)));
    layer2_outputs(1695) <= not(layer1_outputs(9823)) or (layer1_outputs(5902));
    layer2_outputs(1696) <= not(layer1_outputs(6635)) or (layer1_outputs(3654));
    layer2_outputs(1697) <= '1';
    layer2_outputs(1698) <= layer1_outputs(667);
    layer2_outputs(1699) <= (layer1_outputs(3465)) and (layer1_outputs(9099));
    layer2_outputs(1700) <= not((layer1_outputs(8737)) and (layer1_outputs(3488)));
    layer2_outputs(1701) <= (layer1_outputs(2118)) xor (layer1_outputs(791));
    layer2_outputs(1702) <= not(layer1_outputs(3670)) or (layer1_outputs(8542));
    layer2_outputs(1703) <= layer1_outputs(6580);
    layer2_outputs(1704) <= not((layer1_outputs(449)) or (layer1_outputs(486)));
    layer2_outputs(1705) <= not((layer1_outputs(325)) xor (layer1_outputs(7942)));
    layer2_outputs(1706) <= '0';
    layer2_outputs(1707) <= not(layer1_outputs(4567));
    layer2_outputs(1708) <= (layer1_outputs(2190)) and not (layer1_outputs(7137));
    layer2_outputs(1709) <= layer1_outputs(9650);
    layer2_outputs(1710) <= not(layer1_outputs(9122));
    layer2_outputs(1711) <= not(layer1_outputs(740));
    layer2_outputs(1712) <= layer1_outputs(906);
    layer2_outputs(1713) <= not(layer1_outputs(381));
    layer2_outputs(1714) <= not(layer1_outputs(10150));
    layer2_outputs(1715) <= not((layer1_outputs(9459)) and (layer1_outputs(3155)));
    layer2_outputs(1716) <= not(layer1_outputs(4898)) or (layer1_outputs(3699));
    layer2_outputs(1717) <= not((layer1_outputs(1400)) and (layer1_outputs(8182)));
    layer2_outputs(1718) <= (layer1_outputs(4483)) and not (layer1_outputs(8602));
    layer2_outputs(1719) <= not(layer1_outputs(1439)) or (layer1_outputs(5736));
    layer2_outputs(1720) <= not(layer1_outputs(4732));
    layer2_outputs(1721) <= (layer1_outputs(6785)) xor (layer1_outputs(4247));
    layer2_outputs(1722) <= layer1_outputs(10144);
    layer2_outputs(1723) <= not(layer1_outputs(2871));
    layer2_outputs(1724) <= not(layer1_outputs(2243));
    layer2_outputs(1725) <= (layer1_outputs(5016)) and not (layer1_outputs(5119));
    layer2_outputs(1726) <= (layer1_outputs(8866)) and not (layer1_outputs(614));
    layer2_outputs(1727) <= '1';
    layer2_outputs(1728) <= not((layer1_outputs(5571)) and (layer1_outputs(5945)));
    layer2_outputs(1729) <= not(layer1_outputs(4671));
    layer2_outputs(1730) <= not((layer1_outputs(3740)) xor (layer1_outputs(2506)));
    layer2_outputs(1731) <= not(layer1_outputs(6259));
    layer2_outputs(1732) <= not(layer1_outputs(6289));
    layer2_outputs(1733) <= not((layer1_outputs(6664)) xor (layer1_outputs(1780)));
    layer2_outputs(1734) <= layer1_outputs(1966);
    layer2_outputs(1735) <= not(layer1_outputs(3862)) or (layer1_outputs(8105));
    layer2_outputs(1736) <= (layer1_outputs(205)) and not (layer1_outputs(3514));
    layer2_outputs(1737) <= not((layer1_outputs(82)) or (layer1_outputs(739)));
    layer2_outputs(1738) <= (layer1_outputs(9643)) xor (layer1_outputs(7283));
    layer2_outputs(1739) <= not((layer1_outputs(166)) or (layer1_outputs(7406)));
    layer2_outputs(1740) <= not((layer1_outputs(2728)) or (layer1_outputs(9217)));
    layer2_outputs(1741) <= (layer1_outputs(9677)) and not (layer1_outputs(6498));
    layer2_outputs(1742) <= not(layer1_outputs(6537));
    layer2_outputs(1743) <= not(layer1_outputs(1357)) or (layer1_outputs(4893));
    layer2_outputs(1744) <= (layer1_outputs(5859)) and not (layer1_outputs(5263));
    layer2_outputs(1745) <= not((layer1_outputs(3743)) or (layer1_outputs(7210)));
    layer2_outputs(1746) <= layer1_outputs(437);
    layer2_outputs(1747) <= layer1_outputs(2249);
    layer2_outputs(1748) <= not((layer1_outputs(5892)) xor (layer1_outputs(247)));
    layer2_outputs(1749) <= not(layer1_outputs(3530));
    layer2_outputs(1750) <= (layer1_outputs(7358)) and not (layer1_outputs(2088));
    layer2_outputs(1751) <= (layer1_outputs(1715)) and not (layer1_outputs(1279));
    layer2_outputs(1752) <= not((layer1_outputs(9352)) xor (layer1_outputs(162)));
    layer2_outputs(1753) <= '1';
    layer2_outputs(1754) <= not(layer1_outputs(2613));
    layer2_outputs(1755) <= not((layer1_outputs(8001)) xor (layer1_outputs(8948)));
    layer2_outputs(1756) <= (layer1_outputs(8697)) xor (layer1_outputs(4577));
    layer2_outputs(1757) <= not((layer1_outputs(623)) or (layer1_outputs(132)));
    layer2_outputs(1758) <= not(layer1_outputs(6151));
    layer2_outputs(1759) <= not(layer1_outputs(3197));
    layer2_outputs(1760) <= not((layer1_outputs(8796)) xor (layer1_outputs(10066)));
    layer2_outputs(1761) <= not((layer1_outputs(9877)) and (layer1_outputs(2527)));
    layer2_outputs(1762) <= (layer1_outputs(841)) or (layer1_outputs(2757));
    layer2_outputs(1763) <= not((layer1_outputs(9081)) xor (layer1_outputs(334)));
    layer2_outputs(1764) <= '0';
    layer2_outputs(1765) <= '0';
    layer2_outputs(1766) <= not(layer1_outputs(9895));
    layer2_outputs(1767) <= not(layer1_outputs(3580));
    layer2_outputs(1768) <= layer1_outputs(882);
    layer2_outputs(1769) <= layer1_outputs(7983);
    layer2_outputs(1770) <= (layer1_outputs(4768)) and not (layer1_outputs(6516));
    layer2_outputs(1771) <= not((layer1_outputs(2670)) or (layer1_outputs(4133)));
    layer2_outputs(1772) <= not(layer1_outputs(2079));
    layer2_outputs(1773) <= not(layer1_outputs(5948));
    layer2_outputs(1774) <= not((layer1_outputs(917)) and (layer1_outputs(2318)));
    layer2_outputs(1775) <= layer1_outputs(3104);
    layer2_outputs(1776) <= not(layer1_outputs(4307));
    layer2_outputs(1777) <= not(layer1_outputs(7150));
    layer2_outputs(1778) <= (layer1_outputs(3567)) or (layer1_outputs(2796));
    layer2_outputs(1779) <= not((layer1_outputs(634)) and (layer1_outputs(7730)));
    layer2_outputs(1780) <= not((layer1_outputs(60)) or (layer1_outputs(2171)));
    layer2_outputs(1781) <= not(layer1_outputs(4793)) or (layer1_outputs(1516));
    layer2_outputs(1782) <= (layer1_outputs(4522)) and not (layer1_outputs(7209));
    layer2_outputs(1783) <= (layer1_outputs(2883)) and not (layer1_outputs(4823));
    layer2_outputs(1784) <= not((layer1_outputs(5991)) xor (layer1_outputs(7533)));
    layer2_outputs(1785) <= (layer1_outputs(5585)) and not (layer1_outputs(4775));
    layer2_outputs(1786) <= layer1_outputs(755);
    layer2_outputs(1787) <= (layer1_outputs(764)) and not (layer1_outputs(5592));
    layer2_outputs(1788) <= layer1_outputs(9593);
    layer2_outputs(1789) <= (layer1_outputs(5363)) and not (layer1_outputs(6745));
    layer2_outputs(1790) <= layer1_outputs(7645);
    layer2_outputs(1791) <= layer1_outputs(3271);
    layer2_outputs(1792) <= not(layer1_outputs(8292));
    layer2_outputs(1793) <= not(layer1_outputs(4330)) or (layer1_outputs(3593));
    layer2_outputs(1794) <= not(layer1_outputs(6964));
    layer2_outputs(1795) <= '0';
    layer2_outputs(1796) <= layer1_outputs(1550);
    layer2_outputs(1797) <= (layer1_outputs(1232)) and (layer1_outputs(8586));
    layer2_outputs(1798) <= not(layer1_outputs(2426));
    layer2_outputs(1799) <= not(layer1_outputs(2445)) or (layer1_outputs(2473));
    layer2_outputs(1800) <= '1';
    layer2_outputs(1801) <= not((layer1_outputs(4975)) or (layer1_outputs(8430)));
    layer2_outputs(1802) <= not(layer1_outputs(2274));
    layer2_outputs(1803) <= layer1_outputs(6947);
    layer2_outputs(1804) <= not((layer1_outputs(3826)) xor (layer1_outputs(4772)));
    layer2_outputs(1805) <= (layer1_outputs(3921)) xor (layer1_outputs(5369));
    layer2_outputs(1806) <= (layer1_outputs(2904)) and not (layer1_outputs(405));
    layer2_outputs(1807) <= not((layer1_outputs(5510)) or (layer1_outputs(3994)));
    layer2_outputs(1808) <= not(layer1_outputs(626));
    layer2_outputs(1809) <= not(layer1_outputs(5140));
    layer2_outputs(1810) <= (layer1_outputs(8623)) and not (layer1_outputs(7912));
    layer2_outputs(1811) <= not(layer1_outputs(5116)) or (layer1_outputs(9537));
    layer2_outputs(1812) <= not(layer1_outputs(1265)) or (layer1_outputs(3888));
    layer2_outputs(1813) <= layer1_outputs(6618);
    layer2_outputs(1814) <= not((layer1_outputs(6200)) and (layer1_outputs(2029)));
    layer2_outputs(1815) <= (layer1_outputs(8784)) and (layer1_outputs(7575));
    layer2_outputs(1816) <= (layer1_outputs(5507)) or (layer1_outputs(7654));
    layer2_outputs(1817) <= not((layer1_outputs(6149)) xor (layer1_outputs(8676)));
    layer2_outputs(1818) <= layer1_outputs(8635);
    layer2_outputs(1819) <= not((layer1_outputs(1828)) or (layer1_outputs(7310)));
    layer2_outputs(1820) <= not(layer1_outputs(7456)) or (layer1_outputs(4142));
    layer2_outputs(1821) <= layer1_outputs(8358);
    layer2_outputs(1822) <= layer1_outputs(968);
    layer2_outputs(1823) <= layer1_outputs(1779);
    layer2_outputs(1824) <= not(layer1_outputs(7600));
    layer2_outputs(1825) <= layer1_outputs(604);
    layer2_outputs(1826) <= (layer1_outputs(6413)) and not (layer1_outputs(7186));
    layer2_outputs(1827) <= '0';
    layer2_outputs(1828) <= not(layer1_outputs(641));
    layer2_outputs(1829) <= layer1_outputs(6288);
    layer2_outputs(1830) <= not((layer1_outputs(10009)) or (layer1_outputs(4763)));
    layer2_outputs(1831) <= not((layer1_outputs(8542)) or (layer1_outputs(5501)));
    layer2_outputs(1832) <= (layer1_outputs(4042)) xor (layer1_outputs(7185));
    layer2_outputs(1833) <= not(layer1_outputs(8326));
    layer2_outputs(1834) <= (layer1_outputs(6829)) or (layer1_outputs(10188));
    layer2_outputs(1835) <= not(layer1_outputs(567)) or (layer1_outputs(7255));
    layer2_outputs(1836) <= (layer1_outputs(9587)) and not (layer1_outputs(1876));
    layer2_outputs(1837) <= layer1_outputs(4683);
    layer2_outputs(1838) <= (layer1_outputs(120)) and (layer1_outputs(5336));
    layer2_outputs(1839) <= (layer1_outputs(7540)) or (layer1_outputs(4771));
    layer2_outputs(1840) <= (layer1_outputs(4340)) and (layer1_outputs(7493));
    layer2_outputs(1841) <= (layer1_outputs(4645)) and not (layer1_outputs(5216));
    layer2_outputs(1842) <= '1';
    layer2_outputs(1843) <= (layer1_outputs(4477)) and (layer1_outputs(5887));
    layer2_outputs(1844) <= layer1_outputs(8092);
    layer2_outputs(1845) <= not(layer1_outputs(10043));
    layer2_outputs(1846) <= '0';
    layer2_outputs(1847) <= not((layer1_outputs(6255)) xor (layer1_outputs(4419)));
    layer2_outputs(1848) <= not(layer1_outputs(3724));
    layer2_outputs(1849) <= layer1_outputs(3568);
    layer2_outputs(1850) <= not((layer1_outputs(5481)) or (layer1_outputs(5424)));
    layer2_outputs(1851) <= (layer1_outputs(5486)) or (layer1_outputs(5615));
    layer2_outputs(1852) <= not(layer1_outputs(9131));
    layer2_outputs(1853) <= (layer1_outputs(8476)) and (layer1_outputs(6686));
    layer2_outputs(1854) <= (layer1_outputs(4826)) and (layer1_outputs(4267));
    layer2_outputs(1855) <= layer1_outputs(1978);
    layer2_outputs(1856) <= not(layer1_outputs(8399));
    layer2_outputs(1857) <= not(layer1_outputs(1666)) or (layer1_outputs(9376));
    layer2_outputs(1858) <= layer1_outputs(10184);
    layer2_outputs(1859) <= (layer1_outputs(6014)) and not (layer1_outputs(4015));
    layer2_outputs(1860) <= layer1_outputs(7206);
    layer2_outputs(1861) <= not(layer1_outputs(6857)) or (layer1_outputs(9129));
    layer2_outputs(1862) <= not((layer1_outputs(5058)) or (layer1_outputs(2845)));
    layer2_outputs(1863) <= not(layer1_outputs(3361));
    layer2_outputs(1864) <= not((layer1_outputs(6948)) and (layer1_outputs(7483)));
    layer2_outputs(1865) <= layer1_outputs(3515);
    layer2_outputs(1866) <= '0';
    layer2_outputs(1867) <= layer1_outputs(2289);
    layer2_outputs(1868) <= not(layer1_outputs(8742)) or (layer1_outputs(2168));
    layer2_outputs(1869) <= not(layer1_outputs(7870));
    layer2_outputs(1870) <= '0';
    layer2_outputs(1871) <= not(layer1_outputs(973));
    layer2_outputs(1872) <= not(layer1_outputs(3489)) or (layer1_outputs(9708));
    layer2_outputs(1873) <= layer1_outputs(4788);
    layer2_outputs(1874) <= not(layer1_outputs(8957)) or (layer1_outputs(785));
    layer2_outputs(1875) <= not(layer1_outputs(9934));
    layer2_outputs(1876) <= not((layer1_outputs(4127)) and (layer1_outputs(8659)));
    layer2_outputs(1877) <= not(layer1_outputs(3809));
    layer2_outputs(1878) <= (layer1_outputs(3948)) xor (layer1_outputs(6473));
    layer2_outputs(1879) <= (layer1_outputs(6843)) and (layer1_outputs(1870));
    layer2_outputs(1880) <= not(layer1_outputs(105));
    layer2_outputs(1881) <= not((layer1_outputs(6438)) and (layer1_outputs(1865)));
    layer2_outputs(1882) <= not(layer1_outputs(2433));
    layer2_outputs(1883) <= not(layer1_outputs(3555));
    layer2_outputs(1884) <= not(layer1_outputs(845));
    layer2_outputs(1885) <= not(layer1_outputs(1941)) or (layer1_outputs(8878));
    layer2_outputs(1886) <= not(layer1_outputs(10177)) or (layer1_outputs(5007));
    layer2_outputs(1887) <= (layer1_outputs(7955)) and not (layer1_outputs(2578));
    layer2_outputs(1888) <= (layer1_outputs(9458)) and (layer1_outputs(5350));
    layer2_outputs(1889) <= layer1_outputs(907);
    layer2_outputs(1890) <= not((layer1_outputs(1177)) xor (layer1_outputs(7208)));
    layer2_outputs(1891) <= layer1_outputs(3485);
    layer2_outputs(1892) <= not(layer1_outputs(5227));
    layer2_outputs(1893) <= not(layer1_outputs(4939));
    layer2_outputs(1894) <= not((layer1_outputs(1183)) or (layer1_outputs(8775)));
    layer2_outputs(1895) <= layer1_outputs(559);
    layer2_outputs(1896) <= layer1_outputs(7200);
    layer2_outputs(1897) <= not((layer1_outputs(4708)) or (layer1_outputs(6652)));
    layer2_outputs(1898) <= not((layer1_outputs(9855)) xor (layer1_outputs(4207)));
    layer2_outputs(1899) <= (layer1_outputs(823)) and (layer1_outputs(191));
    layer2_outputs(1900) <= layer1_outputs(7442);
    layer2_outputs(1901) <= not((layer1_outputs(1171)) and (layer1_outputs(7632)));
    layer2_outputs(1902) <= not(layer1_outputs(5226));
    layer2_outputs(1903) <= not((layer1_outputs(7031)) or (layer1_outputs(6317)));
    layer2_outputs(1904) <= layer1_outputs(2874);
    layer2_outputs(1905) <= (layer1_outputs(5755)) and not (layer1_outputs(4202));
    layer2_outputs(1906) <= layer1_outputs(6967);
    layer2_outputs(1907) <= not(layer1_outputs(774)) or (layer1_outputs(3589));
    layer2_outputs(1908) <= not(layer1_outputs(8034));
    layer2_outputs(1909) <= (layer1_outputs(8721)) or (layer1_outputs(1737));
    layer2_outputs(1910) <= (layer1_outputs(4486)) or (layer1_outputs(9803));
    layer2_outputs(1911) <= (layer1_outputs(3412)) xor (layer1_outputs(2696));
    layer2_outputs(1912) <= not((layer1_outputs(1978)) or (layer1_outputs(3055)));
    layer2_outputs(1913) <= layer1_outputs(5103);
    layer2_outputs(1914) <= not(layer1_outputs(9689)) or (layer1_outputs(2310));
    layer2_outputs(1915) <= not(layer1_outputs(4863));
    layer2_outputs(1916) <= not(layer1_outputs(3585));
    layer2_outputs(1917) <= layer1_outputs(9341);
    layer2_outputs(1918) <= layer1_outputs(4459);
    layer2_outputs(1919) <= not(layer1_outputs(6559));
    layer2_outputs(1920) <= (layer1_outputs(41)) and (layer1_outputs(8227));
    layer2_outputs(1921) <= (layer1_outputs(589)) xor (layer1_outputs(3293));
    layer2_outputs(1922) <= (layer1_outputs(1304)) and not (layer1_outputs(6928));
    layer2_outputs(1923) <= not(layer1_outputs(5638));
    layer2_outputs(1924) <= (layer1_outputs(7424)) and not (layer1_outputs(4830));
    layer2_outputs(1925) <= (layer1_outputs(1628)) and (layer1_outputs(4442));
    layer2_outputs(1926) <= not(layer1_outputs(5468)) or (layer1_outputs(1238));
    layer2_outputs(1927) <= layer1_outputs(1575);
    layer2_outputs(1928) <= (layer1_outputs(546)) and (layer1_outputs(860));
    layer2_outputs(1929) <= not(layer1_outputs(7216)) or (layer1_outputs(8664));
    layer2_outputs(1930) <= not(layer1_outputs(10206));
    layer2_outputs(1931) <= not(layer1_outputs(2353));
    layer2_outputs(1932) <= not(layer1_outputs(9844));
    layer2_outputs(1933) <= (layer1_outputs(4680)) and not (layer1_outputs(1553));
    layer2_outputs(1934) <= (layer1_outputs(5788)) or (layer1_outputs(9383));
    layer2_outputs(1935) <= (layer1_outputs(3574)) or (layer1_outputs(8920));
    layer2_outputs(1936) <= layer1_outputs(6561);
    layer2_outputs(1937) <= not((layer1_outputs(4231)) or (layer1_outputs(7332)));
    layer2_outputs(1938) <= layer1_outputs(5872);
    layer2_outputs(1939) <= layer1_outputs(6229);
    layer2_outputs(1940) <= not((layer1_outputs(2566)) or (layer1_outputs(8322)));
    layer2_outputs(1941) <= '0';
    layer2_outputs(1942) <= layer1_outputs(6462);
    layer2_outputs(1943) <= layer1_outputs(4827);
    layer2_outputs(1944) <= not(layer1_outputs(8294));
    layer2_outputs(1945) <= (layer1_outputs(8269)) and (layer1_outputs(5569));
    layer2_outputs(1946) <= '1';
    layer2_outputs(1947) <= layer1_outputs(1809);
    layer2_outputs(1948) <= (layer1_outputs(8987)) and (layer1_outputs(1447));
    layer2_outputs(1949) <= not(layer1_outputs(1708));
    layer2_outputs(1950) <= (layer1_outputs(8090)) or (layer1_outputs(3890));
    layer2_outputs(1951) <= not((layer1_outputs(3105)) and (layer1_outputs(8801)));
    layer2_outputs(1952) <= (layer1_outputs(825)) and (layer1_outputs(337));
    layer2_outputs(1953) <= not(layer1_outputs(8077)) or (layer1_outputs(4177));
    layer2_outputs(1954) <= not((layer1_outputs(9917)) or (layer1_outputs(7006)));
    layer2_outputs(1955) <= not(layer1_outputs(9360));
    layer2_outputs(1956) <= (layer1_outputs(7493)) and not (layer1_outputs(1516));
    layer2_outputs(1957) <= not(layer1_outputs(3934));
    layer2_outputs(1958) <= not((layer1_outputs(3370)) xor (layer1_outputs(4384)));
    layer2_outputs(1959) <= not(layer1_outputs(6000)) or (layer1_outputs(440));
    layer2_outputs(1960) <= (layer1_outputs(7293)) or (layer1_outputs(3521));
    layer2_outputs(1961) <= (layer1_outputs(4634)) and not (layer1_outputs(2616));
    layer2_outputs(1962) <= (layer1_outputs(2717)) and not (layer1_outputs(5944));
    layer2_outputs(1963) <= layer1_outputs(1549);
    layer2_outputs(1964) <= not(layer1_outputs(4850));
    layer2_outputs(1965) <= (layer1_outputs(1605)) and (layer1_outputs(7996));
    layer2_outputs(1966) <= not((layer1_outputs(8519)) or (layer1_outputs(9716)));
    layer2_outputs(1967) <= (layer1_outputs(468)) or (layer1_outputs(6017));
    layer2_outputs(1968) <= not(layer1_outputs(3881));
    layer2_outputs(1969) <= not(layer1_outputs(8484));
    layer2_outputs(1970) <= not((layer1_outputs(5034)) xor (layer1_outputs(529)));
    layer2_outputs(1971) <= not(layer1_outputs(4366)) or (layer1_outputs(1068));
    layer2_outputs(1972) <= (layer1_outputs(7807)) or (layer1_outputs(7180));
    layer2_outputs(1973) <= (layer1_outputs(212)) and (layer1_outputs(4210));
    layer2_outputs(1974) <= (layer1_outputs(4366)) and not (layer1_outputs(9338));
    layer2_outputs(1975) <= (layer1_outputs(10118)) xor (layer1_outputs(1125));
    layer2_outputs(1976) <= not((layer1_outputs(4524)) and (layer1_outputs(1395)));
    layer2_outputs(1977) <= not(layer1_outputs(9215)) or (layer1_outputs(8735));
    layer2_outputs(1978) <= layer1_outputs(7682);
    layer2_outputs(1979) <= (layer1_outputs(7829)) xor (layer1_outputs(8681));
    layer2_outputs(1980) <= layer1_outputs(5475);
    layer2_outputs(1981) <= (layer1_outputs(2196)) and (layer1_outputs(1401));
    layer2_outputs(1982) <= not(layer1_outputs(8954));
    layer2_outputs(1983) <= not(layer1_outputs(5861));
    layer2_outputs(1984) <= (layer1_outputs(918)) or (layer1_outputs(1075));
    layer2_outputs(1985) <= layer1_outputs(8803);
    layer2_outputs(1986) <= layer1_outputs(7752);
    layer2_outputs(1987) <= not(layer1_outputs(873));
    layer2_outputs(1988) <= not(layer1_outputs(6091));
    layer2_outputs(1989) <= '1';
    layer2_outputs(1990) <= (layer1_outputs(1528)) and not (layer1_outputs(274));
    layer2_outputs(1991) <= (layer1_outputs(3879)) and (layer1_outputs(7889));
    layer2_outputs(1992) <= '1';
    layer2_outputs(1993) <= layer1_outputs(253);
    layer2_outputs(1994) <= not((layer1_outputs(8094)) xor (layer1_outputs(4733)));
    layer2_outputs(1995) <= layer1_outputs(7720);
    layer2_outputs(1996) <= not((layer1_outputs(9408)) xor (layer1_outputs(4971)));
    layer2_outputs(1997) <= not(layer1_outputs(4362));
    layer2_outputs(1998) <= not((layer1_outputs(5867)) and (layer1_outputs(864)));
    layer2_outputs(1999) <= not(layer1_outputs(7610)) or (layer1_outputs(5081));
    layer2_outputs(2000) <= layer1_outputs(7079);
    layer2_outputs(2001) <= (layer1_outputs(434)) and not (layer1_outputs(463));
    layer2_outputs(2002) <= layer1_outputs(6092);
    layer2_outputs(2003) <= (layer1_outputs(691)) xor (layer1_outputs(517));
    layer2_outputs(2004) <= (layer1_outputs(4105)) xor (layer1_outputs(6102));
    layer2_outputs(2005) <= layer1_outputs(3919);
    layer2_outputs(2006) <= (layer1_outputs(2792)) xor (layer1_outputs(1272));
    layer2_outputs(2007) <= not((layer1_outputs(5883)) and (layer1_outputs(6927)));
    layer2_outputs(2008) <= layer1_outputs(5478);
    layer2_outputs(2009) <= not(layer1_outputs(7728)) or (layer1_outputs(7931));
    layer2_outputs(2010) <= '0';
    layer2_outputs(2011) <= (layer1_outputs(7666)) and not (layer1_outputs(2272));
    layer2_outputs(2012) <= layer1_outputs(6074);
    layer2_outputs(2013) <= layer1_outputs(2653);
    layer2_outputs(2014) <= not(layer1_outputs(9889));
    layer2_outputs(2015) <= layer1_outputs(1837);
    layer2_outputs(2016) <= layer1_outputs(1146);
    layer2_outputs(2017) <= (layer1_outputs(8392)) and (layer1_outputs(8956));
    layer2_outputs(2018) <= layer1_outputs(7548);
    layer2_outputs(2019) <= layer1_outputs(1764);
    layer2_outputs(2020) <= layer1_outputs(9070);
    layer2_outputs(2021) <= layer1_outputs(7829);
    layer2_outputs(2022) <= not(layer1_outputs(400));
    layer2_outputs(2023) <= layer1_outputs(8338);
    layer2_outputs(2024) <= layer1_outputs(5387);
    layer2_outputs(2025) <= '1';
    layer2_outputs(2026) <= not((layer1_outputs(1775)) and (layer1_outputs(1496)));
    layer2_outputs(2027) <= not(layer1_outputs(4360)) or (layer1_outputs(7346));
    layer2_outputs(2028) <= not((layer1_outputs(9222)) xor (layer1_outputs(6001)));
    layer2_outputs(2029) <= layer1_outputs(1121);
    layer2_outputs(2030) <= not((layer1_outputs(6702)) or (layer1_outputs(399)));
    layer2_outputs(2031) <= '0';
    layer2_outputs(2032) <= layer1_outputs(7189);
    layer2_outputs(2033) <= (layer1_outputs(3701)) and (layer1_outputs(4278));
    layer2_outputs(2034) <= layer1_outputs(2975);
    layer2_outputs(2035) <= (layer1_outputs(6345)) and not (layer1_outputs(6870));
    layer2_outputs(2036) <= layer1_outputs(3119);
    layer2_outputs(2037) <= not(layer1_outputs(3788));
    layer2_outputs(2038) <= layer1_outputs(9884);
    layer2_outputs(2039) <= (layer1_outputs(4276)) xor (layer1_outputs(2363));
    layer2_outputs(2040) <= not(layer1_outputs(5247));
    layer2_outputs(2041) <= not(layer1_outputs(4684));
    layer2_outputs(2042) <= (layer1_outputs(5871)) and not (layer1_outputs(1121));
    layer2_outputs(2043) <= not((layer1_outputs(3703)) xor (layer1_outputs(5809)));
    layer2_outputs(2044) <= not((layer1_outputs(8695)) and (layer1_outputs(10148)));
    layer2_outputs(2045) <= layer1_outputs(4506);
    layer2_outputs(2046) <= layer1_outputs(9987);
    layer2_outputs(2047) <= not(layer1_outputs(2791));
    layer2_outputs(2048) <= not(layer1_outputs(9600));
    layer2_outputs(2049) <= layer1_outputs(2698);
    layer2_outputs(2050) <= (layer1_outputs(5674)) and not (layer1_outputs(6591));
    layer2_outputs(2051) <= not((layer1_outputs(1812)) and (layer1_outputs(2823)));
    layer2_outputs(2052) <= not(layer1_outputs(8944)) or (layer1_outputs(1362));
    layer2_outputs(2053) <= not((layer1_outputs(6251)) or (layer1_outputs(4179)));
    layer2_outputs(2054) <= (layer1_outputs(8072)) xor (layer1_outputs(9727));
    layer2_outputs(2055) <= (layer1_outputs(9014)) and not (layer1_outputs(4238));
    layer2_outputs(2056) <= (layer1_outputs(6068)) and (layer1_outputs(3271));
    layer2_outputs(2057) <= not(layer1_outputs(2812));
    layer2_outputs(2058) <= not(layer1_outputs(2234));
    layer2_outputs(2059) <= not((layer1_outputs(1919)) or (layer1_outputs(6814)));
    layer2_outputs(2060) <= not((layer1_outputs(6812)) xor (layer1_outputs(4830)));
    layer2_outputs(2061) <= not(layer1_outputs(4964));
    layer2_outputs(2062) <= not(layer1_outputs(9047));
    layer2_outputs(2063) <= not(layer1_outputs(4346));
    layer2_outputs(2064) <= not(layer1_outputs(4472)) or (layer1_outputs(4545));
    layer2_outputs(2065) <= not(layer1_outputs(8193));
    layer2_outputs(2066) <= (layer1_outputs(171)) and not (layer1_outputs(83));
    layer2_outputs(2067) <= not(layer1_outputs(9528));
    layer2_outputs(2068) <= (layer1_outputs(4382)) and (layer1_outputs(6816));
    layer2_outputs(2069) <= layer1_outputs(6893);
    layer2_outputs(2070) <= (layer1_outputs(5688)) or (layer1_outputs(8395));
    layer2_outputs(2071) <= (layer1_outputs(3110)) and not (layer1_outputs(2466));
    layer2_outputs(2072) <= not(layer1_outputs(10125)) or (layer1_outputs(8933));
    layer2_outputs(2073) <= (layer1_outputs(5767)) and not (layer1_outputs(7915));
    layer2_outputs(2074) <= not((layer1_outputs(898)) or (layer1_outputs(4400)));
    layer2_outputs(2075) <= not(layer1_outputs(5951)) or (layer1_outputs(9066));
    layer2_outputs(2076) <= (layer1_outputs(5625)) and not (layer1_outputs(2844));
    layer2_outputs(2077) <= not((layer1_outputs(1534)) xor (layer1_outputs(6530)));
    layer2_outputs(2078) <= not((layer1_outputs(8533)) xor (layer1_outputs(2997)));
    layer2_outputs(2079) <= layer1_outputs(3483);
    layer2_outputs(2080) <= not((layer1_outputs(6484)) and (layer1_outputs(8424)));
    layer2_outputs(2081) <= not(layer1_outputs(3364));
    layer2_outputs(2082) <= layer1_outputs(9266);
    layer2_outputs(2083) <= not(layer1_outputs(5617));
    layer2_outputs(2084) <= (layer1_outputs(5063)) xor (layer1_outputs(3476));
    layer2_outputs(2085) <= (layer1_outputs(4592)) or (layer1_outputs(2039));
    layer2_outputs(2086) <= not((layer1_outputs(3057)) and (layer1_outputs(9829)));
    layer2_outputs(2087) <= not(layer1_outputs(3108));
    layer2_outputs(2088) <= layer1_outputs(8931);
    layer2_outputs(2089) <= layer1_outputs(6833);
    layer2_outputs(2090) <= not((layer1_outputs(5892)) xor (layer1_outputs(1088)));
    layer2_outputs(2091) <= not(layer1_outputs(3575));
    layer2_outputs(2092) <= not((layer1_outputs(7328)) or (layer1_outputs(2173)));
    layer2_outputs(2093) <= layer1_outputs(3430);
    layer2_outputs(2094) <= (layer1_outputs(6564)) and not (layer1_outputs(5313));
    layer2_outputs(2095) <= (layer1_outputs(5814)) and (layer1_outputs(6567));
    layer2_outputs(2096) <= layer1_outputs(4285);
    layer2_outputs(2097) <= not(layer1_outputs(2363));
    layer2_outputs(2098) <= not((layer1_outputs(6510)) and (layer1_outputs(6758)));
    layer2_outputs(2099) <= not(layer1_outputs(7959)) or (layer1_outputs(2253));
    layer2_outputs(2100) <= layer1_outputs(9683);
    layer2_outputs(2101) <= '0';
    layer2_outputs(2102) <= (layer1_outputs(3927)) and not (layer1_outputs(9060));
    layer2_outputs(2103) <= layer1_outputs(8170);
    layer2_outputs(2104) <= layer1_outputs(2723);
    layer2_outputs(2105) <= not(layer1_outputs(7087));
    layer2_outputs(2106) <= layer1_outputs(6735);
    layer2_outputs(2107) <= (layer1_outputs(8447)) xor (layer1_outputs(3733));
    layer2_outputs(2108) <= (layer1_outputs(9110)) and not (layer1_outputs(6348));
    layer2_outputs(2109) <= not(layer1_outputs(6780)) or (layer1_outputs(3737));
    layer2_outputs(2110) <= not(layer1_outputs(9703));
    layer2_outputs(2111) <= '1';
    layer2_outputs(2112) <= '1';
    layer2_outputs(2113) <= layer1_outputs(5359);
    layer2_outputs(2114) <= layer1_outputs(8769);
    layer2_outputs(2115) <= (layer1_outputs(6799)) or (layer1_outputs(9705));
    layer2_outputs(2116) <= (layer1_outputs(1663)) and not (layer1_outputs(1482));
    layer2_outputs(2117) <= not(layer1_outputs(9276));
    layer2_outputs(2118) <= (layer1_outputs(4528)) xor (layer1_outputs(4749));
    layer2_outputs(2119) <= not((layer1_outputs(9840)) and (layer1_outputs(2874)));
    layer2_outputs(2120) <= (layer1_outputs(5630)) or (layer1_outputs(6420));
    layer2_outputs(2121) <= layer1_outputs(8439);
    layer2_outputs(2122) <= (layer1_outputs(5706)) or (layer1_outputs(1665));
    layer2_outputs(2123) <= layer1_outputs(3457);
    layer2_outputs(2124) <= layer1_outputs(3531);
    layer2_outputs(2125) <= '0';
    layer2_outputs(2126) <= not((layer1_outputs(1109)) xor (layer1_outputs(7536)));
    layer2_outputs(2127) <= not(layer1_outputs(4922)) or (layer1_outputs(6681));
    layer2_outputs(2128) <= not((layer1_outputs(5791)) xor (layer1_outputs(3471)));
    layer2_outputs(2129) <= layer1_outputs(10155);
    layer2_outputs(2130) <= not(layer1_outputs(430));
    layer2_outputs(2131) <= not(layer1_outputs(7377)) or (layer1_outputs(1801));
    layer2_outputs(2132) <= (layer1_outputs(1780)) xor (layer1_outputs(4895));
    layer2_outputs(2133) <= (layer1_outputs(9933)) and not (layer1_outputs(8257));
    layer2_outputs(2134) <= not(layer1_outputs(152));
    layer2_outputs(2135) <= not((layer1_outputs(8914)) or (layer1_outputs(6234)));
    layer2_outputs(2136) <= '1';
    layer2_outputs(2137) <= layer1_outputs(2815);
    layer2_outputs(2138) <= not(layer1_outputs(8808));
    layer2_outputs(2139) <= not(layer1_outputs(2008));
    layer2_outputs(2140) <= (layer1_outputs(2186)) or (layer1_outputs(1598));
    layer2_outputs(2141) <= '1';
    layer2_outputs(2142) <= not((layer1_outputs(6438)) xor (layer1_outputs(1698)));
    layer2_outputs(2143) <= not((layer1_outputs(4099)) and (layer1_outputs(6623)));
    layer2_outputs(2144) <= layer1_outputs(1038);
    layer2_outputs(2145) <= (layer1_outputs(6064)) and not (layer1_outputs(2102));
    layer2_outputs(2146) <= not(layer1_outputs(3292));
    layer2_outputs(2147) <= not((layer1_outputs(9285)) xor (layer1_outputs(258)));
    layer2_outputs(2148) <= layer1_outputs(7914);
    layer2_outputs(2149) <= '1';
    layer2_outputs(2150) <= layer1_outputs(5984);
    layer2_outputs(2151) <= not(layer1_outputs(10234));
    layer2_outputs(2152) <= layer1_outputs(8314);
    layer2_outputs(2153) <= not((layer1_outputs(7703)) xor (layer1_outputs(2959)));
    layer2_outputs(2154) <= layer1_outputs(9811);
    layer2_outputs(2155) <= not(layer1_outputs(3223));
    layer2_outputs(2156) <= layer1_outputs(6132);
    layer2_outputs(2157) <= (layer1_outputs(4882)) and (layer1_outputs(7442));
    layer2_outputs(2158) <= not(layer1_outputs(5684)) or (layer1_outputs(5250));
    layer2_outputs(2159) <= not((layer1_outputs(9603)) xor (layer1_outputs(6134)));
    layer2_outputs(2160) <= not(layer1_outputs(3390));
    layer2_outputs(2161) <= (layer1_outputs(1984)) xor (layer1_outputs(22));
    layer2_outputs(2162) <= (layer1_outputs(5799)) and not (layer1_outputs(3507));
    layer2_outputs(2163) <= not(layer1_outputs(8410)) or (layer1_outputs(801));
    layer2_outputs(2164) <= not((layer1_outputs(5520)) and (layer1_outputs(8517)));
    layer2_outputs(2165) <= not(layer1_outputs(3590));
    layer2_outputs(2166) <= layer1_outputs(6739);
    layer2_outputs(2167) <= not(layer1_outputs(4746));
    layer2_outputs(2168) <= not(layer1_outputs(5756)) or (layer1_outputs(1067));
    layer2_outputs(2169) <= layer1_outputs(138);
    layer2_outputs(2170) <= layer1_outputs(8569);
    layer2_outputs(2171) <= not(layer1_outputs(5810)) or (layer1_outputs(4106));
    layer2_outputs(2172) <= layer1_outputs(6373);
    layer2_outputs(2173) <= '0';
    layer2_outputs(2174) <= not(layer1_outputs(2640));
    layer2_outputs(2175) <= not(layer1_outputs(1187));
    layer2_outputs(2176) <= not(layer1_outputs(6743));
    layer2_outputs(2177) <= (layer1_outputs(7763)) and (layer1_outputs(3904));
    layer2_outputs(2178) <= layer1_outputs(7663);
    layer2_outputs(2179) <= (layer1_outputs(7423)) and not (layer1_outputs(8492));
    layer2_outputs(2180) <= layer1_outputs(10099);
    layer2_outputs(2181) <= '1';
    layer2_outputs(2182) <= layer1_outputs(2124);
    layer2_outputs(2183) <= not((layer1_outputs(307)) xor (layer1_outputs(6084)));
    layer2_outputs(2184) <= not((layer1_outputs(6397)) or (layer1_outputs(5574)));
    layer2_outputs(2185) <= (layer1_outputs(1064)) and not (layer1_outputs(9640));
    layer2_outputs(2186) <= (layer1_outputs(4327)) and not (layer1_outputs(8311));
    layer2_outputs(2187) <= (layer1_outputs(7402)) and (layer1_outputs(5635));
    layer2_outputs(2188) <= not(layer1_outputs(3003));
    layer2_outputs(2189) <= not((layer1_outputs(7685)) and (layer1_outputs(4748)));
    layer2_outputs(2190) <= layer1_outputs(7472);
    layer2_outputs(2191) <= layer1_outputs(9249);
    layer2_outputs(2192) <= not((layer1_outputs(9619)) and (layer1_outputs(8728)));
    layer2_outputs(2193) <= not(layer1_outputs(8727));
    layer2_outputs(2194) <= not((layer1_outputs(5148)) and (layer1_outputs(8660)));
    layer2_outputs(2195) <= '0';
    layer2_outputs(2196) <= layer1_outputs(622);
    layer2_outputs(2197) <= not(layer1_outputs(7697));
    layer2_outputs(2198) <= layer1_outputs(8878);
    layer2_outputs(2199) <= not(layer1_outputs(174)) or (layer1_outputs(5742));
    layer2_outputs(2200) <= not(layer1_outputs(7267));
    layer2_outputs(2201) <= not((layer1_outputs(9980)) and (layer1_outputs(8345)));
    layer2_outputs(2202) <= (layer1_outputs(7739)) or (layer1_outputs(10141));
    layer2_outputs(2203) <= (layer1_outputs(3729)) and not (layer1_outputs(4077));
    layer2_outputs(2204) <= layer1_outputs(7934);
    layer2_outputs(2205) <= (layer1_outputs(1713)) or (layer1_outputs(6610));
    layer2_outputs(2206) <= (layer1_outputs(1604)) or (layer1_outputs(4506));
    layer2_outputs(2207) <= layer1_outputs(9305);
    layer2_outputs(2208) <= not(layer1_outputs(5662));
    layer2_outputs(2209) <= not((layer1_outputs(3004)) or (layer1_outputs(5821)));
    layer2_outputs(2210) <= not((layer1_outputs(3412)) or (layer1_outputs(2469)));
    layer2_outputs(2211) <= (layer1_outputs(3147)) or (layer1_outputs(8018));
    layer2_outputs(2212) <= not(layer1_outputs(7749)) or (layer1_outputs(1948));
    layer2_outputs(2213) <= (layer1_outputs(5812)) or (layer1_outputs(5860));
    layer2_outputs(2214) <= not((layer1_outputs(9672)) or (layer1_outputs(9324)));
    layer2_outputs(2215) <= not(layer1_outputs(3664));
    layer2_outputs(2216) <= (layer1_outputs(3524)) and (layer1_outputs(1714));
    layer2_outputs(2217) <= layer1_outputs(7380);
    layer2_outputs(2218) <= '1';
    layer2_outputs(2219) <= (layer1_outputs(1319)) or (layer1_outputs(3635));
    layer2_outputs(2220) <= '1';
    layer2_outputs(2221) <= layer1_outputs(8230);
    layer2_outputs(2222) <= not(layer1_outputs(2197));
    layer2_outputs(2223) <= '1';
    layer2_outputs(2224) <= (layer1_outputs(9789)) and not (layer1_outputs(8225));
    layer2_outputs(2225) <= not((layer1_outputs(4994)) and (layer1_outputs(4364)));
    layer2_outputs(2226) <= '0';
    layer2_outputs(2227) <= not((layer1_outputs(1836)) and (layer1_outputs(8828)));
    layer2_outputs(2228) <= layer1_outputs(8009);
    layer2_outputs(2229) <= not(layer1_outputs(299)) or (layer1_outputs(363));
    layer2_outputs(2230) <= not(layer1_outputs(2904)) or (layer1_outputs(9838));
    layer2_outputs(2231) <= layer1_outputs(6240);
    layer2_outputs(2232) <= not(layer1_outputs(8695));
    layer2_outputs(2233) <= layer1_outputs(7998);
    layer2_outputs(2234) <= not(layer1_outputs(7864));
    layer2_outputs(2235) <= layer1_outputs(3854);
    layer2_outputs(2236) <= not(layer1_outputs(2373));
    layer2_outputs(2237) <= '0';
    layer2_outputs(2238) <= layer1_outputs(1661);
    layer2_outputs(2239) <= (layer1_outputs(7862)) and (layer1_outputs(8647));
    layer2_outputs(2240) <= not(layer1_outputs(9696)) or (layer1_outputs(9400));
    layer2_outputs(2241) <= (layer1_outputs(7452)) or (layer1_outputs(10014));
    layer2_outputs(2242) <= not(layer1_outputs(2204));
    layer2_outputs(2243) <= layer1_outputs(7181);
    layer2_outputs(2244) <= not((layer1_outputs(1148)) and (layer1_outputs(8702)));
    layer2_outputs(2245) <= (layer1_outputs(5673)) and not (layer1_outputs(5993));
    layer2_outputs(2246) <= not(layer1_outputs(8237));
    layer2_outputs(2247) <= (layer1_outputs(5235)) and not (layer1_outputs(1218));
    layer2_outputs(2248) <= not((layer1_outputs(518)) xor (layer1_outputs(3853)));
    layer2_outputs(2249) <= layer1_outputs(8596);
    layer2_outputs(2250) <= not(layer1_outputs(5616));
    layer2_outputs(2251) <= layer1_outputs(4906);
    layer2_outputs(2252) <= not(layer1_outputs(6611)) or (layer1_outputs(800));
    layer2_outputs(2253) <= not(layer1_outputs(6581));
    layer2_outputs(2254) <= '0';
    layer2_outputs(2255) <= not(layer1_outputs(8437));
    layer2_outputs(2256) <= not((layer1_outputs(424)) or (layer1_outputs(5534)));
    layer2_outputs(2257) <= (layer1_outputs(5632)) and not (layer1_outputs(9432));
    layer2_outputs(2258) <= (layer1_outputs(7781)) and (layer1_outputs(8989));
    layer2_outputs(2259) <= (layer1_outputs(9701)) and not (layer1_outputs(5523));
    layer2_outputs(2260) <= layer1_outputs(2533);
    layer2_outputs(2261) <= not(layer1_outputs(3068));
    layer2_outputs(2262) <= not(layer1_outputs(647)) or (layer1_outputs(9765));
    layer2_outputs(2263) <= layer1_outputs(5200);
    layer2_outputs(2264) <= layer1_outputs(8666);
    layer2_outputs(2265) <= not(layer1_outputs(1367));
    layer2_outputs(2266) <= layer1_outputs(8870);
    layer2_outputs(2267) <= layer1_outputs(3989);
    layer2_outputs(2268) <= '1';
    layer2_outputs(2269) <= (layer1_outputs(7344)) and not (layer1_outputs(5646));
    layer2_outputs(2270) <= not(layer1_outputs(9338));
    layer2_outputs(2271) <= layer1_outputs(5346);
    layer2_outputs(2272) <= layer1_outputs(7272);
    layer2_outputs(2273) <= (layer1_outputs(5536)) and not (layer1_outputs(3988));
    layer2_outputs(2274) <= not(layer1_outputs(6235));
    layer2_outputs(2275) <= '1';
    layer2_outputs(2276) <= layer1_outputs(8987);
    layer2_outputs(2277) <= not((layer1_outputs(375)) or (layer1_outputs(10018)));
    layer2_outputs(2278) <= (layer1_outputs(996)) and not (layer1_outputs(4784));
    layer2_outputs(2279) <= (layer1_outputs(7190)) xor (layer1_outputs(7535));
    layer2_outputs(2280) <= (layer1_outputs(9404)) and not (layer1_outputs(7812));
    layer2_outputs(2281) <= layer1_outputs(2959);
    layer2_outputs(2282) <= not((layer1_outputs(7880)) xor (layer1_outputs(7073)));
    layer2_outputs(2283) <= (layer1_outputs(3794)) and not (layer1_outputs(9486));
    layer2_outputs(2284) <= layer1_outputs(4672);
    layer2_outputs(2285) <= not(layer1_outputs(9882));
    layer2_outputs(2286) <= layer1_outputs(746);
    layer2_outputs(2287) <= (layer1_outputs(8080)) or (layer1_outputs(2097));
    layer2_outputs(2288) <= not(layer1_outputs(6669));
    layer2_outputs(2289) <= not(layer1_outputs(8926));
    layer2_outputs(2290) <= not(layer1_outputs(2756)) or (layer1_outputs(4585));
    layer2_outputs(2291) <= not(layer1_outputs(1493));
    layer2_outputs(2292) <= '0';
    layer2_outputs(2293) <= not(layer1_outputs(3797));
    layer2_outputs(2294) <= (layer1_outputs(9194)) and not (layer1_outputs(733));
    layer2_outputs(2295) <= layer1_outputs(6570);
    layer2_outputs(2296) <= not((layer1_outputs(1103)) and (layer1_outputs(6734)));
    layer2_outputs(2297) <= layer1_outputs(7821);
    layer2_outputs(2298) <= not((layer1_outputs(7723)) and (layer1_outputs(7577)));
    layer2_outputs(2299) <= layer1_outputs(2910);
    layer2_outputs(2300) <= not(layer1_outputs(5848));
    layer2_outputs(2301) <= layer1_outputs(7243);
    layer2_outputs(2302) <= (layer1_outputs(1947)) and (layer1_outputs(2231));
    layer2_outputs(2303) <= layer1_outputs(9567);
    layer2_outputs(2304) <= not(layer1_outputs(156)) or (layer1_outputs(3951));
    layer2_outputs(2305) <= not(layer1_outputs(4677)) or (layer1_outputs(3317));
    layer2_outputs(2306) <= not((layer1_outputs(2241)) and (layer1_outputs(255)));
    layer2_outputs(2307) <= layer1_outputs(1626);
    layer2_outputs(2308) <= (layer1_outputs(2586)) and (layer1_outputs(9847));
    layer2_outputs(2309) <= not((layer1_outputs(4424)) xor (layer1_outputs(4397)));
    layer2_outputs(2310) <= (layer1_outputs(8927)) xor (layer1_outputs(8259));
    layer2_outputs(2311) <= not(layer1_outputs(1756)) or (layer1_outputs(7113));
    layer2_outputs(2312) <= not(layer1_outputs(942)) or (layer1_outputs(3435));
    layer2_outputs(2313) <= (layer1_outputs(9582)) xor (layer1_outputs(8207));
    layer2_outputs(2314) <= not((layer1_outputs(7331)) and (layer1_outputs(8961)));
    layer2_outputs(2315) <= '1';
    layer2_outputs(2316) <= not(layer1_outputs(266));
    layer2_outputs(2317) <= (layer1_outputs(2336)) xor (layer1_outputs(9469));
    layer2_outputs(2318) <= (layer1_outputs(5203)) and (layer1_outputs(9331));
    layer2_outputs(2319) <= (layer1_outputs(204)) or (layer1_outputs(4227));
    layer2_outputs(2320) <= layer1_outputs(1601);
    layer2_outputs(2321) <= (layer1_outputs(9821)) and (layer1_outputs(3423));
    layer2_outputs(2322) <= not((layer1_outputs(6388)) or (layer1_outputs(1092)));
    layer2_outputs(2323) <= not(layer1_outputs(185)) or (layer1_outputs(4576));
    layer2_outputs(2324) <= not((layer1_outputs(3876)) and (layer1_outputs(7221)));
    layer2_outputs(2325) <= layer1_outputs(5323);
    layer2_outputs(2326) <= not(layer1_outputs(4641)) or (layer1_outputs(5925));
    layer2_outputs(2327) <= (layer1_outputs(3847)) and (layer1_outputs(3210));
    layer2_outputs(2328) <= layer1_outputs(5505);
    layer2_outputs(2329) <= layer1_outputs(2404);
    layer2_outputs(2330) <= not((layer1_outputs(7992)) or (layer1_outputs(1288)));
    layer2_outputs(2331) <= (layer1_outputs(2206)) and (layer1_outputs(4911));
    layer2_outputs(2332) <= not(layer1_outputs(10013));
    layer2_outputs(2333) <= not(layer1_outputs(8535)) or (layer1_outputs(1740));
    layer2_outputs(2334) <= (layer1_outputs(8579)) or (layer1_outputs(5357));
    layer2_outputs(2335) <= not(layer1_outputs(7585));
    layer2_outputs(2336) <= layer1_outputs(5150);
    layer2_outputs(2337) <= not((layer1_outputs(9501)) or (layer1_outputs(340)));
    layer2_outputs(2338) <= (layer1_outputs(7932)) or (layer1_outputs(1728));
    layer2_outputs(2339) <= (layer1_outputs(5528)) xor (layer1_outputs(5759));
    layer2_outputs(2340) <= not((layer1_outputs(8027)) and (layer1_outputs(2632)));
    layer2_outputs(2341) <= (layer1_outputs(4540)) or (layer1_outputs(5074));
    layer2_outputs(2342) <= layer1_outputs(3572);
    layer2_outputs(2343) <= '0';
    layer2_outputs(2344) <= '1';
    layer2_outputs(2345) <= (layer1_outputs(9216)) and not (layer1_outputs(8178));
    layer2_outputs(2346) <= not(layer1_outputs(3877));
    layer2_outputs(2347) <= (layer1_outputs(4598)) and not (layer1_outputs(7395));
    layer2_outputs(2348) <= not(layer1_outputs(9755));
    layer2_outputs(2349) <= layer1_outputs(5234);
    layer2_outputs(2350) <= (layer1_outputs(8591)) and not (layer1_outputs(4041));
    layer2_outputs(2351) <= not(layer1_outputs(5863));
    layer2_outputs(2352) <= (layer1_outputs(5121)) and (layer1_outputs(6493));
    layer2_outputs(2353) <= not((layer1_outputs(6388)) xor (layer1_outputs(6416)));
    layer2_outputs(2354) <= layer1_outputs(356);
    layer2_outputs(2355) <= not(layer1_outputs(5441)) or (layer1_outputs(642));
    layer2_outputs(2356) <= not(layer1_outputs(6622));
    layer2_outputs(2357) <= layer1_outputs(7284);
    layer2_outputs(2358) <= (layer1_outputs(3144)) and not (layer1_outputs(4162));
    layer2_outputs(2359) <= (layer1_outputs(8272)) or (layer1_outputs(6671));
    layer2_outputs(2360) <= (layer1_outputs(264)) and not (layer1_outputs(4107));
    layer2_outputs(2361) <= '0';
    layer2_outputs(2362) <= not((layer1_outputs(1727)) or (layer1_outputs(4909)));
    layer2_outputs(2363) <= '1';
    layer2_outputs(2364) <= not((layer1_outputs(4597)) and (layer1_outputs(3393)));
    layer2_outputs(2365) <= '0';
    layer2_outputs(2366) <= (layer1_outputs(10233)) or (layer1_outputs(5470));
    layer2_outputs(2367) <= not((layer1_outputs(7938)) xor (layer1_outputs(5934)));
    layer2_outputs(2368) <= layer1_outputs(9690);
    layer2_outputs(2369) <= not(layer1_outputs(4407));
    layer2_outputs(2370) <= layer1_outputs(6027);
    layer2_outputs(2371) <= not(layer1_outputs(9189)) or (layer1_outputs(1488));
    layer2_outputs(2372) <= not((layer1_outputs(3976)) xor (layer1_outputs(6713)));
    layer2_outputs(2373) <= not((layer1_outputs(4002)) and (layer1_outputs(6244)));
    layer2_outputs(2374) <= layer1_outputs(9364);
    layer2_outputs(2375) <= (layer1_outputs(4974)) or (layer1_outputs(1243));
    layer2_outputs(2376) <= '0';
    layer2_outputs(2377) <= not(layer1_outputs(8221));
    layer2_outputs(2378) <= (layer1_outputs(3823)) xor (layer1_outputs(487));
    layer2_outputs(2379) <= '1';
    layer2_outputs(2380) <= (layer1_outputs(4306)) and not (layer1_outputs(9564));
    layer2_outputs(2381) <= not(layer1_outputs(1982)) or (layer1_outputs(5716));
    layer2_outputs(2382) <= (layer1_outputs(5900)) or (layer1_outputs(1053));
    layer2_outputs(2383) <= (layer1_outputs(7987)) or (layer1_outputs(996));
    layer2_outputs(2384) <= not((layer1_outputs(1650)) or (layer1_outputs(3933)));
    layer2_outputs(2385) <= (layer1_outputs(6014)) xor (layer1_outputs(7139));
    layer2_outputs(2386) <= not(layer1_outputs(4565));
    layer2_outputs(2387) <= layer1_outputs(1206);
    layer2_outputs(2388) <= not(layer1_outputs(8032)) or (layer1_outputs(9380));
    layer2_outputs(2389) <= layer1_outputs(8510);
    layer2_outputs(2390) <= (layer1_outputs(7671)) and not (layer1_outputs(3320));
    layer2_outputs(2391) <= (layer1_outputs(349)) and not (layer1_outputs(2507));
    layer2_outputs(2392) <= (layer1_outputs(2823)) or (layer1_outputs(610));
    layer2_outputs(2393) <= not(layer1_outputs(8037));
    layer2_outputs(2394) <= layer1_outputs(7564);
    layer2_outputs(2395) <= (layer1_outputs(1343)) and (layer1_outputs(4729));
    layer2_outputs(2396) <= (layer1_outputs(9902)) and not (layer1_outputs(9733));
    layer2_outputs(2397) <= layer1_outputs(6358);
    layer2_outputs(2398) <= not((layer1_outputs(230)) xor (layer1_outputs(7114)));
    layer2_outputs(2399) <= (layer1_outputs(2075)) or (layer1_outputs(9905));
    layer2_outputs(2400) <= not((layer1_outputs(6535)) xor (layer1_outputs(1517)));
    layer2_outputs(2401) <= (layer1_outputs(5868)) and (layer1_outputs(9302));
    layer2_outputs(2402) <= not(layer1_outputs(2073)) or (layer1_outputs(8604));
    layer2_outputs(2403) <= not(layer1_outputs(5119));
    layer2_outputs(2404) <= layer1_outputs(6702);
    layer2_outputs(2405) <= (layer1_outputs(4572)) and not (layer1_outputs(73));
    layer2_outputs(2406) <= '1';
    layer2_outputs(2407) <= layer1_outputs(8753);
    layer2_outputs(2408) <= not((layer1_outputs(10173)) xor (layer1_outputs(5929)));
    layer2_outputs(2409) <= not(layer1_outputs(8620)) or (layer1_outputs(7326));
    layer2_outputs(2410) <= layer1_outputs(1229);
    layer2_outputs(2411) <= not((layer1_outputs(6513)) and (layer1_outputs(4668)));
    layer2_outputs(2412) <= layer1_outputs(6805);
    layer2_outputs(2413) <= '0';
    layer2_outputs(2414) <= not(layer1_outputs(3871)) or (layer1_outputs(494));
    layer2_outputs(2415) <= not(layer1_outputs(1339));
    layer2_outputs(2416) <= (layer1_outputs(6858)) or (layer1_outputs(10175));
    layer2_outputs(2417) <= not(layer1_outputs(5429));
    layer2_outputs(2418) <= not((layer1_outputs(7429)) or (layer1_outputs(99)));
    layer2_outputs(2419) <= not((layer1_outputs(2898)) or (layer1_outputs(1340)));
    layer2_outputs(2420) <= (layer1_outputs(1857)) and not (layer1_outputs(2341));
    layer2_outputs(2421) <= not(layer1_outputs(4288));
    layer2_outputs(2422) <= layer1_outputs(7779);
    layer2_outputs(2423) <= layer1_outputs(5709);
    layer2_outputs(2424) <= not((layer1_outputs(8992)) and (layer1_outputs(8023)));
    layer2_outputs(2425) <= layer1_outputs(9504);
    layer2_outputs(2426) <= not(layer1_outputs(8526));
    layer2_outputs(2427) <= not(layer1_outputs(805));
    layer2_outputs(2428) <= layer1_outputs(9739);
    layer2_outputs(2429) <= (layer1_outputs(6816)) and (layer1_outputs(5116));
    layer2_outputs(2430) <= layer1_outputs(4769);
    layer2_outputs(2431) <= (layer1_outputs(930)) and not (layer1_outputs(5411));
    layer2_outputs(2432) <= (layer1_outputs(1226)) and not (layer1_outputs(4091));
    layer2_outputs(2433) <= not(layer1_outputs(6296)) or (layer1_outputs(3235));
    layer2_outputs(2434) <= (layer1_outputs(649)) and not (layer1_outputs(7948));
    layer2_outputs(2435) <= not((layer1_outputs(7123)) or (layer1_outputs(773)));
    layer2_outputs(2436) <= (layer1_outputs(7349)) and not (layer1_outputs(2380));
    layer2_outputs(2437) <= not((layer1_outputs(2041)) xor (layer1_outputs(5607)));
    layer2_outputs(2438) <= (layer1_outputs(4947)) and not (layer1_outputs(5072));
    layer2_outputs(2439) <= layer1_outputs(6807);
    layer2_outputs(2440) <= layer1_outputs(6077);
    layer2_outputs(2441) <= not(layer1_outputs(7070)) or (layer1_outputs(2807));
    layer2_outputs(2442) <= not((layer1_outputs(9402)) or (layer1_outputs(872)));
    layer2_outputs(2443) <= (layer1_outputs(328)) and (layer1_outputs(1412));
    layer2_outputs(2444) <= (layer1_outputs(2452)) or (layer1_outputs(6414));
    layer2_outputs(2445) <= not((layer1_outputs(9225)) or (layer1_outputs(4951)));
    layer2_outputs(2446) <= not(layer1_outputs(3489));
    layer2_outputs(2447) <= (layer1_outputs(369)) and not (layer1_outputs(10198));
    layer2_outputs(2448) <= not((layer1_outputs(5427)) xor (layer1_outputs(3120)));
    layer2_outputs(2449) <= not((layer1_outputs(3945)) and (layer1_outputs(7469)));
    layer2_outputs(2450) <= not(layer1_outputs(1166)) or (layer1_outputs(5487));
    layer2_outputs(2451) <= not(layer1_outputs(6071));
    layer2_outputs(2452) <= not((layer1_outputs(3592)) or (layer1_outputs(1261)));
    layer2_outputs(2453) <= layer1_outputs(5914);
    layer2_outputs(2454) <= not((layer1_outputs(6885)) xor (layer1_outputs(9969)));
    layer2_outputs(2455) <= (layer1_outputs(3695)) and not (layer1_outputs(2575));
    layer2_outputs(2456) <= not(layer1_outputs(1009));
    layer2_outputs(2457) <= layer1_outputs(9629);
    layer2_outputs(2458) <= not(layer1_outputs(5453)) or (layer1_outputs(1646));
    layer2_outputs(2459) <= layer1_outputs(3781);
    layer2_outputs(2460) <= layer1_outputs(7033);
    layer2_outputs(2461) <= layer1_outputs(9707);
    layer2_outputs(2462) <= layer1_outputs(2658);
    layer2_outputs(2463) <= (layer1_outputs(4638)) and not (layer1_outputs(2990));
    layer2_outputs(2464) <= not(layer1_outputs(478)) or (layer1_outputs(60));
    layer2_outputs(2465) <= layer1_outputs(158);
    layer2_outputs(2466) <= layer1_outputs(6305);
    layer2_outputs(2467) <= (layer1_outputs(2538)) and not (layer1_outputs(5058));
    layer2_outputs(2468) <= (layer1_outputs(4239)) and (layer1_outputs(6701));
    layer2_outputs(2469) <= not(layer1_outputs(5022));
    layer2_outputs(2470) <= not((layer1_outputs(3869)) and (layer1_outputs(6969)));
    layer2_outputs(2471) <= not(layer1_outputs(8853));
    layer2_outputs(2472) <= layer1_outputs(9943);
    layer2_outputs(2473) <= (layer1_outputs(365)) and not (layer1_outputs(4215));
    layer2_outputs(2474) <= (layer1_outputs(2064)) and (layer1_outputs(6662));
    layer2_outputs(2475) <= layer1_outputs(9509);
    layer2_outputs(2476) <= not(layer1_outputs(8356));
    layer2_outputs(2477) <= not((layer1_outputs(10055)) or (layer1_outputs(7780)));
    layer2_outputs(2478) <= not(layer1_outputs(2424));
    layer2_outputs(2479) <= not((layer1_outputs(1360)) and (layer1_outputs(9207)));
    layer2_outputs(2480) <= layer1_outputs(1973);
    layer2_outputs(2481) <= (layer1_outputs(5285)) xor (layer1_outputs(7567));
    layer2_outputs(2482) <= not(layer1_outputs(1674)) or (layer1_outputs(9052));
    layer2_outputs(2483) <= layer1_outputs(3900);
    layer2_outputs(2484) <= not((layer1_outputs(3618)) or (layer1_outputs(7491)));
    layer2_outputs(2485) <= not(layer1_outputs(759));
    layer2_outputs(2486) <= not((layer1_outputs(3661)) xor (layer1_outputs(5781)));
    layer2_outputs(2487) <= not(layer1_outputs(8451));
    layer2_outputs(2488) <= '1';
    layer2_outputs(2489) <= (layer1_outputs(7593)) and not (layer1_outputs(1658));
    layer2_outputs(2490) <= not((layer1_outputs(6960)) and (layer1_outputs(4312)));
    layer2_outputs(2491) <= layer1_outputs(410);
    layer2_outputs(2492) <= not(layer1_outputs(9488)) or (layer1_outputs(9094));
    layer2_outputs(2493) <= not(layer1_outputs(7112));
    layer2_outputs(2494) <= '0';
    layer2_outputs(2495) <= '1';
    layer2_outputs(2496) <= (layer1_outputs(9430)) or (layer1_outputs(342));
    layer2_outputs(2497) <= not(layer1_outputs(4233)) or (layer1_outputs(4861));
    layer2_outputs(2498) <= (layer1_outputs(5681)) or (layer1_outputs(1491));
    layer2_outputs(2499) <= layer1_outputs(3964);
    layer2_outputs(2500) <= layer1_outputs(169);
    layer2_outputs(2501) <= not(layer1_outputs(2781));
    layer2_outputs(2502) <= not(layer1_outputs(5105));
    layer2_outputs(2503) <= layer1_outputs(9399);
    layer2_outputs(2504) <= (layer1_outputs(6143)) or (layer1_outputs(6943));
    layer2_outputs(2505) <= not(layer1_outputs(9348)) or (layer1_outputs(3861));
    layer2_outputs(2506) <= (layer1_outputs(2799)) or (layer1_outputs(4921));
    layer2_outputs(2507) <= (layer1_outputs(8804)) and not (layer1_outputs(3974));
    layer2_outputs(2508) <= '0';
    layer2_outputs(2509) <= not(layer1_outputs(5684));
    layer2_outputs(2510) <= layer1_outputs(7894);
    layer2_outputs(2511) <= not(layer1_outputs(9546)) or (layer1_outputs(8367));
    layer2_outputs(2512) <= not((layer1_outputs(10112)) and (layer1_outputs(8409)));
    layer2_outputs(2513) <= not((layer1_outputs(7553)) xor (layer1_outputs(7013)));
    layer2_outputs(2514) <= (layer1_outputs(3659)) and (layer1_outputs(2421));
    layer2_outputs(2515) <= (layer1_outputs(5933)) or (layer1_outputs(5066));
    layer2_outputs(2516) <= layer1_outputs(52);
    layer2_outputs(2517) <= layer1_outputs(3628);
    layer2_outputs(2518) <= layer1_outputs(8069);
    layer2_outputs(2519) <= not(layer1_outputs(330));
    layer2_outputs(2520) <= layer1_outputs(8);
    layer2_outputs(2521) <= layer1_outputs(2349);
    layer2_outputs(2522) <= not((layer1_outputs(2018)) or (layer1_outputs(7347)));
    layer2_outputs(2523) <= not((layer1_outputs(4183)) or (layer1_outputs(962)));
    layer2_outputs(2524) <= not(layer1_outputs(7159));
    layer2_outputs(2525) <= (layer1_outputs(6638)) and not (layer1_outputs(6376));
    layer2_outputs(2526) <= (layer1_outputs(1135)) or (layer1_outputs(5397));
    layer2_outputs(2527) <= not((layer1_outputs(2416)) xor (layer1_outputs(4747)));
    layer2_outputs(2528) <= not(layer1_outputs(7973)) or (layer1_outputs(6784));
    layer2_outputs(2529) <= not(layer1_outputs(8058)) or (layer1_outputs(9721));
    layer2_outputs(2530) <= layer1_outputs(5269);
    layer2_outputs(2531) <= not((layer1_outputs(1964)) or (layer1_outputs(5665)));
    layer2_outputs(2532) <= not(layer1_outputs(1998));
    layer2_outputs(2533) <= layer1_outputs(2849);
    layer2_outputs(2534) <= layer1_outputs(10104);
    layer2_outputs(2535) <= (layer1_outputs(9401)) or (layer1_outputs(4260));
    layer2_outputs(2536) <= not(layer1_outputs(9520)) or (layer1_outputs(6459));
    layer2_outputs(2537) <= (layer1_outputs(4458)) xor (layer1_outputs(6633));
    layer2_outputs(2538) <= not(layer1_outputs(6482));
    layer2_outputs(2539) <= (layer1_outputs(3438)) or (layer1_outputs(3486));
    layer2_outputs(2540) <= (layer1_outputs(5746)) xor (layer1_outputs(2024));
    layer2_outputs(2541) <= '1';
    layer2_outputs(2542) <= not((layer1_outputs(3539)) and (layer1_outputs(7684)));
    layer2_outputs(2543) <= not(layer1_outputs(1683));
    layer2_outputs(2544) <= not(layer1_outputs(8376));
    layer2_outputs(2545) <= not(layer1_outputs(3551));
    layer2_outputs(2546) <= not((layer1_outputs(1160)) xor (layer1_outputs(4413)));
    layer2_outputs(2547) <= (layer1_outputs(6513)) and (layer1_outputs(3042));
    layer2_outputs(2548) <= not(layer1_outputs(1198)) or (layer1_outputs(3461));
    layer2_outputs(2549) <= layer1_outputs(9654);
    layer2_outputs(2550) <= (layer1_outputs(5036)) or (layer1_outputs(6001));
    layer2_outputs(2551) <= not((layer1_outputs(563)) xor (layer1_outputs(1005)));
    layer2_outputs(2552) <= not((layer1_outputs(521)) and (layer1_outputs(9856)));
    layer2_outputs(2553) <= layer1_outputs(3333);
    layer2_outputs(2554) <= not((layer1_outputs(7653)) or (layer1_outputs(6779)));
    layer2_outputs(2555) <= (layer1_outputs(3570)) and not (layer1_outputs(7869));
    layer2_outputs(2556) <= not(layer1_outputs(3484));
    layer2_outputs(2557) <= (layer1_outputs(6629)) and not (layer1_outputs(6180));
    layer2_outputs(2558) <= layer1_outputs(8434);
    layer2_outputs(2559) <= not((layer1_outputs(9999)) or (layer1_outputs(726)));
    layer2_outputs(2560) <= layer1_outputs(9073);
    layer2_outputs(2561) <= not(layer1_outputs(3323)) or (layer1_outputs(9596));
    layer2_outputs(2562) <= (layer1_outputs(1637)) and not (layer1_outputs(1540));
    layer2_outputs(2563) <= not(layer1_outputs(277));
    layer2_outputs(2564) <= layer1_outputs(253);
    layer2_outputs(2565) <= layer1_outputs(8184);
    layer2_outputs(2566) <= (layer1_outputs(1384)) or (layer1_outputs(1540));
    layer2_outputs(2567) <= (layer1_outputs(8156)) xor (layer1_outputs(5572));
    layer2_outputs(2568) <= layer1_outputs(7844);
    layer2_outputs(2569) <= not((layer1_outputs(9203)) and (layer1_outputs(4261)));
    layer2_outputs(2570) <= (layer1_outputs(2642)) and not (layer1_outputs(7284));
    layer2_outputs(2571) <= (layer1_outputs(1608)) and (layer1_outputs(989));
    layer2_outputs(2572) <= layer1_outputs(1720);
    layer2_outputs(2573) <= not((layer1_outputs(3157)) or (layer1_outputs(722)));
    layer2_outputs(2574) <= layer1_outputs(726);
    layer2_outputs(2575) <= not(layer1_outputs(7974));
    layer2_outputs(2576) <= (layer1_outputs(2965)) or (layer1_outputs(8847));
    layer2_outputs(2577) <= '0';
    layer2_outputs(2578) <= not((layer1_outputs(3111)) and (layer1_outputs(4852)));
    layer2_outputs(2579) <= (layer1_outputs(6138)) or (layer1_outputs(9800));
    layer2_outputs(2580) <= layer1_outputs(1757);
    layer2_outputs(2581) <= not((layer1_outputs(9983)) xor (layer1_outputs(3924)));
    layer2_outputs(2582) <= not((layer1_outputs(412)) xor (layer1_outputs(7370)));
    layer2_outputs(2583) <= not((layer1_outputs(3529)) xor (layer1_outputs(8862)));
    layer2_outputs(2584) <= layer1_outputs(3468);
    layer2_outputs(2585) <= layer1_outputs(10071);
    layer2_outputs(2586) <= layer1_outputs(3112);
    layer2_outputs(2587) <= (layer1_outputs(4834)) or (layer1_outputs(43));
    layer2_outputs(2588) <= not(layer1_outputs(7075));
    layer2_outputs(2589) <= (layer1_outputs(1327)) or (layer1_outputs(2354));
    layer2_outputs(2590) <= not((layer1_outputs(932)) xor (layer1_outputs(1006)));
    layer2_outputs(2591) <= (layer1_outputs(5166)) and not (layer1_outputs(510));
    layer2_outputs(2592) <= not(layer1_outputs(9720));
    layer2_outputs(2593) <= layer1_outputs(3452);
    layer2_outputs(2594) <= layer1_outputs(9468);
    layer2_outputs(2595) <= not(layer1_outputs(7624)) or (layer1_outputs(6302));
    layer2_outputs(2596) <= '0';
    layer2_outputs(2597) <= (layer1_outputs(9170)) and not (layer1_outputs(3571));
    layer2_outputs(2598) <= layer1_outputs(6136);
    layer2_outputs(2599) <= (layer1_outputs(2739)) and (layer1_outputs(10184));
    layer2_outputs(2600) <= layer1_outputs(6333);
    layer2_outputs(2601) <= (layer1_outputs(7025)) or (layer1_outputs(9013));
    layer2_outputs(2602) <= (layer1_outputs(1094)) and not (layer1_outputs(6503));
    layer2_outputs(2603) <= not(layer1_outputs(2040));
    layer2_outputs(2604) <= not(layer1_outputs(8218));
    layer2_outputs(2605) <= layer1_outputs(2246);
    layer2_outputs(2606) <= not((layer1_outputs(1950)) and (layer1_outputs(8629)));
    layer2_outputs(2607) <= not((layer1_outputs(1377)) xor (layer1_outputs(2356)));
    layer2_outputs(2608) <= '0';
    layer2_outputs(2609) <= (layer1_outputs(8150)) and not (layer1_outputs(695));
    layer2_outputs(2610) <= not(layer1_outputs(240));
    layer2_outputs(2611) <= not((layer1_outputs(1337)) xor (layer1_outputs(7635)));
    layer2_outputs(2612) <= layer1_outputs(2047);
    layer2_outputs(2613) <= not(layer1_outputs(7110)) or (layer1_outputs(5793));
    layer2_outputs(2614) <= not(layer1_outputs(3006));
    layer2_outputs(2615) <= not(layer1_outputs(420)) or (layer1_outputs(5002));
    layer2_outputs(2616) <= layer1_outputs(5808);
    layer2_outputs(2617) <= layer1_outputs(6783);
    layer2_outputs(2618) <= not(layer1_outputs(2130));
    layer2_outputs(2619) <= not((layer1_outputs(501)) or (layer1_outputs(2628)));
    layer2_outputs(2620) <= not(layer1_outputs(5858));
    layer2_outputs(2621) <= '0';
    layer2_outputs(2622) <= not(layer1_outputs(3474)) or (layer1_outputs(3098));
    layer2_outputs(2623) <= layer1_outputs(2658);
    layer2_outputs(2624) <= not(layer1_outputs(6297));
    layer2_outputs(2625) <= not(layer1_outputs(114));
    layer2_outputs(2626) <= layer1_outputs(711);
    layer2_outputs(2627) <= not(layer1_outputs(7777));
    layer2_outputs(2628) <= not(layer1_outputs(7585));
    layer2_outputs(2629) <= layer1_outputs(7330);
    layer2_outputs(2630) <= (layer1_outputs(5049)) and not (layer1_outputs(7019));
    layer2_outputs(2631) <= (layer1_outputs(8064)) or (layer1_outputs(1691));
    layer2_outputs(2632) <= not(layer1_outputs(9874)) or (layer1_outputs(5629));
    layer2_outputs(2633) <= (layer1_outputs(1329)) xor (layer1_outputs(5088));
    layer2_outputs(2634) <= not((layer1_outputs(6526)) xor (layer1_outputs(1342)));
    layer2_outputs(2635) <= layer1_outputs(9296);
    layer2_outputs(2636) <= layer1_outputs(4844);
    layer2_outputs(2637) <= '0';
    layer2_outputs(2638) <= layer1_outputs(895);
    layer2_outputs(2639) <= (layer1_outputs(784)) and not (layer1_outputs(2423));
    layer2_outputs(2640) <= not(layer1_outputs(5150));
    layer2_outputs(2641) <= not(layer1_outputs(753));
    layer2_outputs(2642) <= not(layer1_outputs(8587));
    layer2_outputs(2643) <= not(layer1_outputs(1860));
    layer2_outputs(2644) <= not(layer1_outputs(5776));
    layer2_outputs(2645) <= layer1_outputs(3036);
    layer2_outputs(2646) <= (layer1_outputs(8456)) and not (layer1_outputs(3400));
    layer2_outputs(2647) <= not(layer1_outputs(9731)) or (layer1_outputs(7030));
    layer2_outputs(2648) <= layer1_outputs(5875);
    layer2_outputs(2649) <= not(layer1_outputs(8934));
    layer2_outputs(2650) <= not((layer1_outputs(3133)) and (layer1_outputs(4202)));
    layer2_outputs(2651) <= not((layer1_outputs(1423)) xor (layer1_outputs(656)));
    layer2_outputs(2652) <= '1';
    layer2_outputs(2653) <= not(layer1_outputs(5811)) or (layer1_outputs(5530));
    layer2_outputs(2654) <= layer1_outputs(9545);
    layer2_outputs(2655) <= (layer1_outputs(2880)) and not (layer1_outputs(3140));
    layer2_outputs(2656) <= not(layer1_outputs(987)) or (layer1_outputs(2897));
    layer2_outputs(2657) <= not((layer1_outputs(1573)) xor (layer1_outputs(7272)));
    layer2_outputs(2658) <= (layer1_outputs(9499)) xor (layer1_outputs(9441));
    layer2_outputs(2659) <= layer1_outputs(3583);
    layer2_outputs(2660) <= (layer1_outputs(7611)) and not (layer1_outputs(7942));
    layer2_outputs(2661) <= layer1_outputs(2953);
    layer2_outputs(2662) <= layer1_outputs(5127);
    layer2_outputs(2663) <= (layer1_outputs(5008)) or (layer1_outputs(6768));
    layer2_outputs(2664) <= (layer1_outputs(9135)) and not (layer1_outputs(8531));
    layer2_outputs(2665) <= not(layer1_outputs(7058));
    layer2_outputs(2666) <= not(layer1_outputs(61));
    layer2_outputs(2667) <= layer1_outputs(2619);
    layer2_outputs(2668) <= layer1_outputs(1141);
    layer2_outputs(2669) <= not((layer1_outputs(2464)) or (layer1_outputs(4071)));
    layer2_outputs(2670) <= '0';
    layer2_outputs(2671) <= not((layer1_outputs(7447)) and (layer1_outputs(844)));
    layer2_outputs(2672) <= (layer1_outputs(954)) and not (layer1_outputs(1513));
    layer2_outputs(2673) <= not((layer1_outputs(404)) xor (layer1_outputs(9047)));
    layer2_outputs(2674) <= not(layer1_outputs(9141));
    layer2_outputs(2675) <= not(layer1_outputs(3421)) or (layer1_outputs(6395));
    layer2_outputs(2676) <= not((layer1_outputs(9184)) and (layer1_outputs(5483)));
    layer2_outputs(2677) <= not((layer1_outputs(3714)) and (layer1_outputs(4098)));
    layer2_outputs(2678) <= '1';
    layer2_outputs(2679) <= not((layer1_outputs(7301)) or (layer1_outputs(7257)));
    layer2_outputs(2680) <= not(layer1_outputs(2050));
    layer2_outputs(2681) <= not(layer1_outputs(9944));
    layer2_outputs(2682) <= not((layer1_outputs(5663)) or (layer1_outputs(9345)));
    layer2_outputs(2683) <= (layer1_outputs(2831)) xor (layer1_outputs(5391));
    layer2_outputs(2684) <= not(layer1_outputs(9039));
    layer2_outputs(2685) <= not(layer1_outputs(3128)) or (layer1_outputs(8862));
    layer2_outputs(2686) <= layer1_outputs(7688);
    layer2_outputs(2687) <= (layer1_outputs(986)) or (layer1_outputs(6982));
    layer2_outputs(2688) <= not(layer1_outputs(9595));
    layer2_outputs(2689) <= not((layer1_outputs(1923)) or (layer1_outputs(6741)));
    layer2_outputs(2690) <= (layer1_outputs(3776)) and (layer1_outputs(1344));
    layer2_outputs(2691) <= (layer1_outputs(614)) or (layer1_outputs(3912));
    layer2_outputs(2692) <= (layer1_outputs(8306)) xor (layer1_outputs(902));
    layer2_outputs(2693) <= '1';
    layer2_outputs(2694) <= (layer1_outputs(9852)) and not (layer1_outputs(9983));
    layer2_outputs(2695) <= not(layer1_outputs(9921));
    layer2_outputs(2696) <= not((layer1_outputs(1926)) or (layer1_outputs(1026)));
    layer2_outputs(2697) <= (layer1_outputs(1018)) and not (layer1_outputs(2821));
    layer2_outputs(2698) <= not((layer1_outputs(9043)) or (layer1_outputs(3859)));
    layer2_outputs(2699) <= not((layer1_outputs(1866)) or (layer1_outputs(347)));
    layer2_outputs(2700) <= not((layer1_outputs(1113)) or (layer1_outputs(1668)));
    layer2_outputs(2701) <= not((layer1_outputs(1387)) xor (layer1_outputs(895)));
    layer2_outputs(2702) <= (layer1_outputs(1644)) and (layer1_outputs(7273));
    layer2_outputs(2703) <= not((layer1_outputs(3000)) xor (layer1_outputs(216)));
    layer2_outputs(2704) <= (layer1_outputs(2563)) and not (layer1_outputs(6615));
    layer2_outputs(2705) <= not(layer1_outputs(4989)) or (layer1_outputs(1480));
    layer2_outputs(2706) <= not(layer1_outputs(4408)) or (layer1_outputs(5610));
    layer2_outputs(2707) <= not(layer1_outputs(9299)) or (layer1_outputs(9653));
    layer2_outputs(2708) <= not((layer1_outputs(4847)) and (layer1_outputs(949)));
    layer2_outputs(2709) <= '1';
    layer2_outputs(2710) <= not(layer1_outputs(9702));
    layer2_outputs(2711) <= not(layer1_outputs(6226));
    layer2_outputs(2712) <= not((layer1_outputs(3779)) xor (layer1_outputs(2455)));
    layer2_outputs(2713) <= '1';
    layer2_outputs(2714) <= layer1_outputs(4558);
    layer2_outputs(2715) <= (layer1_outputs(9244)) or (layer1_outputs(4875));
    layer2_outputs(2716) <= not((layer1_outputs(7805)) and (layer1_outputs(9041)));
    layer2_outputs(2717) <= not((layer1_outputs(2840)) xor (layer1_outputs(2009)));
    layer2_outputs(2718) <= not(layer1_outputs(4442));
    layer2_outputs(2719) <= not((layer1_outputs(9188)) or (layer1_outputs(5309)));
    layer2_outputs(2720) <= layer1_outputs(6460);
    layer2_outputs(2721) <= not((layer1_outputs(2982)) or (layer1_outputs(7141)));
    layer2_outputs(2722) <= not(layer1_outputs(1372));
    layer2_outputs(2723) <= layer1_outputs(6706);
    layer2_outputs(2724) <= layer1_outputs(7529);
    layer2_outputs(2725) <= (layer1_outputs(3885)) or (layer1_outputs(7432));
    layer2_outputs(2726) <= (layer1_outputs(9652)) and not (layer1_outputs(5104));
    layer2_outputs(2727) <= (layer1_outputs(2158)) or (layer1_outputs(4031));
    layer2_outputs(2728) <= layer1_outputs(931);
    layer2_outputs(2729) <= not((layer1_outputs(6552)) or (layer1_outputs(5922)));
    layer2_outputs(2730) <= (layer1_outputs(1248)) and not (layer1_outputs(5201));
    layer2_outputs(2731) <= (layer1_outputs(4858)) and not (layer1_outputs(10127));
    layer2_outputs(2732) <= not(layer1_outputs(3104));
    layer2_outputs(2733) <= (layer1_outputs(2605)) and (layer1_outputs(8937));
    layer2_outputs(2734) <= layer1_outputs(639);
    layer2_outputs(2735) <= not(layer1_outputs(572));
    layer2_outputs(2736) <= not(layer1_outputs(6931)) or (layer1_outputs(4005));
    layer2_outputs(2737) <= layer1_outputs(8932);
    layer2_outputs(2738) <= not(layer1_outputs(5515));
    layer2_outputs(2739) <= not(layer1_outputs(2444)) or (layer1_outputs(900));
    layer2_outputs(2740) <= (layer1_outputs(5449)) or (layer1_outputs(506));
    layer2_outputs(2741) <= not((layer1_outputs(3253)) or (layer1_outputs(2480)));
    layer2_outputs(2742) <= '0';
    layer2_outputs(2743) <= layer1_outputs(5179);
    layer2_outputs(2744) <= not(layer1_outputs(5872));
    layer2_outputs(2745) <= layer1_outputs(5414);
    layer2_outputs(2746) <= (layer1_outputs(3354)) and not (layer1_outputs(701));
    layer2_outputs(2747) <= not(layer1_outputs(5209));
    layer2_outputs(2748) <= layer1_outputs(8521);
    layer2_outputs(2749) <= layer1_outputs(2012);
    layer2_outputs(2750) <= not(layer1_outputs(4488)) or (layer1_outputs(6251));
    layer2_outputs(2751) <= not(layer1_outputs(2184));
    layer2_outputs(2752) <= not(layer1_outputs(4300));
    layer2_outputs(2753) <= (layer1_outputs(4635)) and not (layer1_outputs(9116));
    layer2_outputs(2754) <= (layer1_outputs(5492)) and (layer1_outputs(1450));
    layer2_outputs(2755) <= layer1_outputs(6735);
    layer2_outputs(2756) <= layer1_outputs(530);
    layer2_outputs(2757) <= not((layer1_outputs(7068)) and (layer1_outputs(4705)));
    layer2_outputs(2758) <= (layer1_outputs(3486)) or (layer1_outputs(7978));
    layer2_outputs(2759) <= layer1_outputs(222);
    layer2_outputs(2760) <= (layer1_outputs(8847)) xor (layer1_outputs(6002));
    layer2_outputs(2761) <= (layer1_outputs(4980)) or (layer1_outputs(2687));
    layer2_outputs(2762) <= not(layer1_outputs(612)) or (layer1_outputs(9776));
    layer2_outputs(2763) <= (layer1_outputs(6851)) and (layer1_outputs(257));
    layer2_outputs(2764) <= not(layer1_outputs(4471)) or (layer1_outputs(4264));
    layer2_outputs(2765) <= not(layer1_outputs(5332));
    layer2_outputs(2766) <= '0';
    layer2_outputs(2767) <= not(layer1_outputs(5959));
    layer2_outputs(2768) <= layer1_outputs(1073);
    layer2_outputs(2769) <= not((layer1_outputs(1995)) and (layer1_outputs(2765)));
    layer2_outputs(2770) <= not(layer1_outputs(7200));
    layer2_outputs(2771) <= not(layer1_outputs(7135));
    layer2_outputs(2772) <= not(layer1_outputs(137));
    layer2_outputs(2773) <= layer1_outputs(1162);
    layer2_outputs(2774) <= layer1_outputs(8606);
    layer2_outputs(2775) <= '0';
    layer2_outputs(2776) <= not((layer1_outputs(2726)) xor (layer1_outputs(8304)));
    layer2_outputs(2777) <= (layer1_outputs(2830)) or (layer1_outputs(7573));
    layer2_outputs(2778) <= (layer1_outputs(3961)) and not (layer1_outputs(7785));
    layer2_outputs(2779) <= '1';
    layer2_outputs(2780) <= layer1_outputs(4136);
    layer2_outputs(2781) <= not(layer1_outputs(6304));
    layer2_outputs(2782) <= not(layer1_outputs(4821));
    layer2_outputs(2783) <= not(layer1_outputs(7383));
    layer2_outputs(2784) <= (layer1_outputs(8134)) and not (layer1_outputs(6625));
    layer2_outputs(2785) <= not((layer1_outputs(6205)) and (layer1_outputs(8832)));
    layer2_outputs(2786) <= not((layer1_outputs(4944)) xor (layer1_outputs(8813)));
    layer2_outputs(2787) <= not(layer1_outputs(7981));
    layer2_outputs(2788) <= not((layer1_outputs(1318)) and (layer1_outputs(3685)));
    layer2_outputs(2789) <= (layer1_outputs(1117)) or (layer1_outputs(8348));
    layer2_outputs(2790) <= layer1_outputs(8889);
    layer2_outputs(2791) <= not(layer1_outputs(5439));
    layer2_outputs(2792) <= not(layer1_outputs(734));
    layer2_outputs(2793) <= not(layer1_outputs(1578)) or (layer1_outputs(1735));
    layer2_outputs(2794) <= layer1_outputs(5562);
    layer2_outputs(2795) <= layer1_outputs(8244);
    layer2_outputs(2796) <= not(layer1_outputs(6891));
    layer2_outputs(2797) <= not(layer1_outputs(8979));
    layer2_outputs(2798) <= layer1_outputs(9476);
    layer2_outputs(2799) <= (layer1_outputs(3462)) and (layer1_outputs(515));
    layer2_outputs(2800) <= (layer1_outputs(8662)) xor (layer1_outputs(3933));
    layer2_outputs(2801) <= (layer1_outputs(8979)) xor (layer1_outputs(8371));
    layer2_outputs(2802) <= not(layer1_outputs(7917));
    layer2_outputs(2803) <= not(layer1_outputs(2463));
    layer2_outputs(2804) <= (layer1_outputs(81)) xor (layer1_outputs(4882));
    layer2_outputs(2805) <= not(layer1_outputs(3578)) or (layer1_outputs(6353));
    layer2_outputs(2806) <= layer1_outputs(9766);
    layer2_outputs(2807) <= not((layer1_outputs(4095)) or (layer1_outputs(4045)));
    layer2_outputs(2808) <= (layer1_outputs(2139)) and not (layer1_outputs(2654));
    layer2_outputs(2809) <= (layer1_outputs(9628)) and not (layer1_outputs(2756));
    layer2_outputs(2810) <= '0';
    layer2_outputs(2811) <= not((layer1_outputs(9785)) or (layer1_outputs(6342)));
    layer2_outputs(2812) <= '0';
    layer2_outputs(2813) <= '1';
    layer2_outputs(2814) <= (layer1_outputs(1391)) and not (layer1_outputs(9169));
    layer2_outputs(2815) <= (layer1_outputs(72)) xor (layer1_outputs(7808));
    layer2_outputs(2816) <= not(layer1_outputs(3246));
    layer2_outputs(2817) <= not(layer1_outputs(6763)) or (layer1_outputs(7679));
    layer2_outputs(2818) <= (layer1_outputs(3415)) xor (layer1_outputs(1236));
    layer2_outputs(2819) <= (layer1_outputs(9321)) and not (layer1_outputs(2414));
    layer2_outputs(2820) <= not((layer1_outputs(1747)) or (layer1_outputs(4494)));
    layer2_outputs(2821) <= layer1_outputs(7636);
    layer2_outputs(2822) <= not(layer1_outputs(1649));
    layer2_outputs(2823) <= not(layer1_outputs(6854));
    layer2_outputs(2824) <= not(layer1_outputs(5795));
    layer2_outputs(2825) <= '0';
    layer2_outputs(2826) <= not((layer1_outputs(1233)) or (layer1_outputs(933)));
    layer2_outputs(2827) <= layer1_outputs(5067);
    layer2_outputs(2828) <= layer1_outputs(5482);
    layer2_outputs(2829) <= layer1_outputs(5442);
    layer2_outputs(2830) <= layer1_outputs(6964);
    layer2_outputs(2831) <= not(layer1_outputs(736)) or (layer1_outputs(1246));
    layer2_outputs(2832) <= '1';
    layer2_outputs(2833) <= (layer1_outputs(6827)) or (layer1_outputs(9698));
    layer2_outputs(2834) <= layer1_outputs(2955);
    layer2_outputs(2835) <= layer1_outputs(4590);
    layer2_outputs(2836) <= layer1_outputs(1429);
    layer2_outputs(2837) <= (layer1_outputs(8863)) xor (layer1_outputs(3499));
    layer2_outputs(2838) <= (layer1_outputs(9893)) and (layer1_outputs(355));
    layer2_outputs(2839) <= layer1_outputs(4583);
    layer2_outputs(2840) <= not(layer1_outputs(8815)) or (layer1_outputs(5169));
    layer2_outputs(2841) <= '0';
    layer2_outputs(2842) <= (layer1_outputs(6773)) and (layer1_outputs(5202));
    layer2_outputs(2843) <= layer1_outputs(4262);
    layer2_outputs(2844) <= not(layer1_outputs(3280)) or (layer1_outputs(6124));
    layer2_outputs(2845) <= layer1_outputs(2176);
    layer2_outputs(2846) <= (layer1_outputs(9372)) and (layer1_outputs(4131));
    layer2_outputs(2847) <= layer1_outputs(9735);
    layer2_outputs(2848) <= not(layer1_outputs(1374));
    layer2_outputs(2849) <= not(layer1_outputs(5331));
    layer2_outputs(2850) <= layer1_outputs(3267);
    layer2_outputs(2851) <= '1';
    layer2_outputs(2852) <= layer1_outputs(3923);
    layer2_outputs(2853) <= not((layer1_outputs(5039)) or (layer1_outputs(2601)));
    layer2_outputs(2854) <= (layer1_outputs(9726)) or (layer1_outputs(3391));
    layer2_outputs(2855) <= layer1_outputs(9105);
    layer2_outputs(2856) <= not(layer1_outputs(6372));
    layer2_outputs(2857) <= not((layer1_outputs(9677)) xor (layer1_outputs(5179)));
    layer2_outputs(2858) <= not((layer1_outputs(407)) xor (layer1_outputs(2516)));
    layer2_outputs(2859) <= not((layer1_outputs(7764)) or (layer1_outputs(2293)));
    layer2_outputs(2860) <= not((layer1_outputs(7265)) xor (layer1_outputs(5836)));
    layer2_outputs(2861) <= (layer1_outputs(4378)) and not (layer1_outputs(9291));
    layer2_outputs(2862) <= (layer1_outputs(4553)) and (layer1_outputs(7696));
    layer2_outputs(2863) <= '1';
    layer2_outputs(2864) <= not((layer1_outputs(8952)) or (layer1_outputs(4487)));
    layer2_outputs(2865) <= (layer1_outputs(9941)) and not (layer1_outputs(7909));
    layer2_outputs(2866) <= not(layer1_outputs(3297)) or (layer1_outputs(5642));
    layer2_outputs(2867) <= (layer1_outputs(5595)) and not (layer1_outputs(9405));
    layer2_outputs(2868) <= layer1_outputs(131);
    layer2_outputs(2869) <= (layer1_outputs(7023)) and (layer1_outputs(7596));
    layer2_outputs(2870) <= layer1_outputs(3645);
    layer2_outputs(2871) <= not((layer1_outputs(9917)) or (layer1_outputs(2359)));
    layer2_outputs(2872) <= not(layer1_outputs(9377));
    layer2_outputs(2873) <= layer1_outputs(10023);
    layer2_outputs(2874) <= (layer1_outputs(2143)) and not (layer1_outputs(2387));
    layer2_outputs(2875) <= (layer1_outputs(9293)) and not (layer1_outputs(10175));
    layer2_outputs(2876) <= not(layer1_outputs(2617));
    layer2_outputs(2877) <= (layer1_outputs(2125)) xor (layer1_outputs(1048));
    layer2_outputs(2878) <= '1';
    layer2_outputs(2879) <= (layer1_outputs(2119)) xor (layer1_outputs(596));
    layer2_outputs(2880) <= not(layer1_outputs(7220));
    layer2_outputs(2881) <= not(layer1_outputs(2273));
    layer2_outputs(2882) <= not((layer1_outputs(2176)) and (layer1_outputs(7134)));
    layer2_outputs(2883) <= (layer1_outputs(1939)) and not (layer1_outputs(6980));
    layer2_outputs(2884) <= not(layer1_outputs(2668));
    layer2_outputs(2885) <= layer1_outputs(6118);
    layer2_outputs(2886) <= not(layer1_outputs(1213)) or (layer1_outputs(110));
    layer2_outputs(2887) <= not((layer1_outputs(5970)) or (layer1_outputs(8524)));
    layer2_outputs(2888) <= (layer1_outputs(3631)) and not (layer1_outputs(1427));
    layer2_outputs(2889) <= not(layer1_outputs(1738));
    layer2_outputs(2890) <= '1';
    layer2_outputs(2891) <= not(layer1_outputs(3013));
    layer2_outputs(2892) <= not((layer1_outputs(292)) xor (layer1_outputs(6607)));
    layer2_outputs(2893) <= not((layer1_outputs(7751)) xor (layer1_outputs(1307)));
    layer2_outputs(2894) <= layer1_outputs(9394);
    layer2_outputs(2895) <= (layer1_outputs(251)) and not (layer1_outputs(2364));
    layer2_outputs(2896) <= (layer1_outputs(4457)) and not (layer1_outputs(5097));
    layer2_outputs(2897) <= (layer1_outputs(762)) xor (layer1_outputs(8762));
    layer2_outputs(2898) <= layer1_outputs(2068);
    layer2_outputs(2899) <= layer1_outputs(4065);
    layer2_outputs(2900) <= not(layer1_outputs(10068)) or (layer1_outputs(1368));
    layer2_outputs(2901) <= layer1_outputs(4560);
    layer2_outputs(2902) <= '1';
    layer2_outputs(2903) <= (layer1_outputs(200)) or (layer1_outputs(6408));
    layer2_outputs(2904) <= layer1_outputs(7561);
    layer2_outputs(2905) <= not(layer1_outputs(4530));
    layer2_outputs(2906) <= not(layer1_outputs(5135)) or (layer1_outputs(6505));
    layer2_outputs(2907) <= not(layer1_outputs(9587)) or (layer1_outputs(7974));
    layer2_outputs(2908) <= layer1_outputs(6884);
    layer2_outputs(2909) <= '1';
    layer2_outputs(2910) <= not(layer1_outputs(1961)) or (layer1_outputs(6432));
    layer2_outputs(2911) <= not(layer1_outputs(5152)) or (layer1_outputs(7105));
    layer2_outputs(2912) <= not(layer1_outputs(2929));
    layer2_outputs(2913) <= not(layer1_outputs(8838));
    layer2_outputs(2914) <= '1';
    layer2_outputs(2915) <= not(layer1_outputs(10239));
    layer2_outputs(2916) <= layer1_outputs(1079);
    layer2_outputs(2917) <= not(layer1_outputs(4953)) or (layer1_outputs(713));
    layer2_outputs(2918) <= (layer1_outputs(10095)) and not (layer1_outputs(1739));
    layer2_outputs(2919) <= '1';
    layer2_outputs(2920) <= not((layer1_outputs(7090)) xor (layer1_outputs(712)));
    layer2_outputs(2921) <= not(layer1_outputs(8158)) or (layer1_outputs(5489));
    layer2_outputs(2922) <= (layer1_outputs(1827)) xor (layer1_outputs(4049));
    layer2_outputs(2923) <= not(layer1_outputs(9039));
    layer2_outputs(2924) <= not(layer1_outputs(9653));
    layer2_outputs(2925) <= not(layer1_outputs(7973));
    layer2_outputs(2926) <= (layer1_outputs(5920)) and (layer1_outputs(4314));
    layer2_outputs(2927) <= (layer1_outputs(2648)) and (layer1_outputs(2225));
    layer2_outputs(2928) <= not(layer1_outputs(3542));
    layer2_outputs(2929) <= layer1_outputs(9260);
    layer2_outputs(2930) <= not((layer1_outputs(3614)) and (layer1_outputs(1032)));
    layer2_outputs(2931) <= '0';
    layer2_outputs(2932) <= not((layer1_outputs(1587)) xor (layer1_outputs(7551)));
    layer2_outputs(2933) <= layer1_outputs(6185);
    layer2_outputs(2934) <= not((layer1_outputs(8343)) xor (layer1_outputs(9859)));
    layer2_outputs(2935) <= (layer1_outputs(10141)) or (layer1_outputs(7475));
    layer2_outputs(2936) <= (layer1_outputs(8441)) and not (layer1_outputs(6863));
    layer2_outputs(2937) <= (layer1_outputs(6160)) and not (layer1_outputs(1483));
    layer2_outputs(2938) <= layer1_outputs(9772);
    layer2_outputs(2939) <= layer1_outputs(10084);
    layer2_outputs(2940) <= '1';
    layer2_outputs(2941) <= layer1_outputs(924);
    layer2_outputs(2942) <= (layer1_outputs(10167)) and not (layer1_outputs(2119));
    layer2_outputs(2943) <= not((layer1_outputs(2432)) or (layer1_outputs(6147)));
    layer2_outputs(2944) <= not(layer1_outputs(3523));
    layer2_outputs(2945) <= (layer1_outputs(7831)) or (layer1_outputs(7718));
    layer2_outputs(2946) <= not((layer1_outputs(2794)) or (layer1_outputs(7028)));
    layer2_outputs(2947) <= layer1_outputs(358);
    layer2_outputs(2948) <= layer1_outputs(10017);
    layer2_outputs(2949) <= layer1_outputs(5351);
    layer2_outputs(2950) <= not(layer1_outputs(9127));
    layer2_outputs(2951) <= not(layer1_outputs(4450)) or (layer1_outputs(4793));
    layer2_outputs(2952) <= '0';
    layer2_outputs(2953) <= not(layer1_outputs(1786));
    layer2_outputs(2954) <= not(layer1_outputs(5664)) or (layer1_outputs(9749));
    layer2_outputs(2955) <= (layer1_outputs(6512)) and not (layer1_outputs(2299));
    layer2_outputs(2956) <= layer1_outputs(5599);
    layer2_outputs(2957) <= not(layer1_outputs(8437));
    layer2_outputs(2958) <= not(layer1_outputs(9098));
    layer2_outputs(2959) <= '0';
    layer2_outputs(2960) <= not((layer1_outputs(435)) or (layer1_outputs(8554)));
    layer2_outputs(2961) <= (layer1_outputs(6549)) or (layer1_outputs(3926));
    layer2_outputs(2962) <= not(layer1_outputs(5174));
    layer2_outputs(2963) <= not(layer1_outputs(8912)) or (layer1_outputs(6918));
    layer2_outputs(2964) <= not(layer1_outputs(8963)) or (layer1_outputs(5436));
    layer2_outputs(2965) <= not(layer1_outputs(3849));
    layer2_outputs(2966) <= not((layer1_outputs(5834)) xor (layer1_outputs(5388)));
    layer2_outputs(2967) <= '0';
    layer2_outputs(2968) <= (layer1_outputs(7566)) and not (layer1_outputs(7508));
    layer2_outputs(2969) <= layer1_outputs(1886);
    layer2_outputs(2970) <= (layer1_outputs(9304)) and not (layer1_outputs(4138));
    layer2_outputs(2971) <= (layer1_outputs(8272)) and not (layer1_outputs(7801));
    layer2_outputs(2972) <= layer1_outputs(1535);
    layer2_outputs(2973) <= (layer1_outputs(7842)) and not (layer1_outputs(9357));
    layer2_outputs(2974) <= (layer1_outputs(10170)) and not (layer1_outputs(9420));
    layer2_outputs(2975) <= layer1_outputs(6016);
    layer2_outputs(2976) <= not(layer1_outputs(7784));
    layer2_outputs(2977) <= not(layer1_outputs(2612));
    layer2_outputs(2978) <= not(layer1_outputs(2894)) or (layer1_outputs(1859));
    layer2_outputs(2979) <= not(layer1_outputs(8640));
    layer2_outputs(2980) <= (layer1_outputs(5503)) and not (layer1_outputs(1560));
    layer2_outputs(2981) <= not((layer1_outputs(2162)) and (layer1_outputs(946)));
    layer2_outputs(2982) <= layer1_outputs(7624);
    layer2_outputs(2983) <= not((layer1_outputs(7954)) xor (layer1_outputs(2144)));
    layer2_outputs(2984) <= (layer1_outputs(10174)) and (layer1_outputs(8044));
    layer2_outputs(2985) <= layer1_outputs(9635);
    layer2_outputs(2986) <= (layer1_outputs(10065)) and (layer1_outputs(2419));
    layer2_outputs(2987) <= not((layer1_outputs(9795)) and (layer1_outputs(179)));
    layer2_outputs(2988) <= not(layer1_outputs(5769));
    layer2_outputs(2989) <= not(layer1_outputs(1831));
    layer2_outputs(2990) <= not((layer1_outputs(7496)) and (layer1_outputs(831)));
    layer2_outputs(2991) <= (layer1_outputs(5025)) xor (layer1_outputs(8599));
    layer2_outputs(2992) <= (layer1_outputs(4109)) and not (layer1_outputs(9045));
    layer2_outputs(2993) <= (layer1_outputs(4408)) and not (layer1_outputs(3648));
    layer2_outputs(2994) <= '1';
    layer2_outputs(2995) <= not(layer1_outputs(2338));
    layer2_outputs(2996) <= (layer1_outputs(7155)) and not (layer1_outputs(8865));
    layer2_outputs(2997) <= not((layer1_outputs(1196)) or (layer1_outputs(5524)));
    layer2_outputs(2998) <= not((layer1_outputs(5246)) or (layer1_outputs(4731)));
    layer2_outputs(2999) <= layer1_outputs(662);
    layer2_outputs(3000) <= not(layer1_outputs(894));
    layer2_outputs(3001) <= layer1_outputs(3892);
    layer2_outputs(3002) <= not(layer1_outputs(2094));
    layer2_outputs(3003) <= not(layer1_outputs(8691));
    layer2_outputs(3004) <= layer1_outputs(4079);
    layer2_outputs(3005) <= not(layer1_outputs(4975));
    layer2_outputs(3006) <= not(layer1_outputs(7691));
    layer2_outputs(3007) <= not(layer1_outputs(2021));
    layer2_outputs(3008) <= not(layer1_outputs(1298));
    layer2_outputs(3009) <= layer1_outputs(9624);
    layer2_outputs(3010) <= not((layer1_outputs(7154)) and (layer1_outputs(246)));
    layer2_outputs(3011) <= layer1_outputs(9308);
    layer2_outputs(3012) <= (layer1_outputs(6655)) or (layer1_outputs(6534));
    layer2_outputs(3013) <= (layer1_outputs(2285)) and not (layer1_outputs(5594));
    layer2_outputs(3014) <= not(layer1_outputs(1124));
    layer2_outputs(3015) <= not(layer1_outputs(7598));
    layer2_outputs(3016) <= not((layer1_outputs(6406)) or (layer1_outputs(2046)));
    layer2_outputs(3017) <= not(layer1_outputs(288));
    layer2_outputs(3018) <= layer1_outputs(6495);
    layer2_outputs(3019) <= not(layer1_outputs(1571)) or (layer1_outputs(2966));
    layer2_outputs(3020) <= not(layer1_outputs(7832));
    layer2_outputs(3021) <= not(layer1_outputs(5799));
    layer2_outputs(3022) <= layer1_outputs(4035);
    layer2_outputs(3023) <= not((layer1_outputs(2521)) or (layer1_outputs(7490)));
    layer2_outputs(3024) <= '0';
    layer2_outputs(3025) <= '0';
    layer2_outputs(3026) <= not(layer1_outputs(9060));
    layer2_outputs(3027) <= layer1_outputs(4465);
    layer2_outputs(3028) <= not(layer1_outputs(3066));
    layer2_outputs(3029) <= layer1_outputs(5283);
    layer2_outputs(3030) <= (layer1_outputs(1636)) xor (layer1_outputs(482));
    layer2_outputs(3031) <= (layer1_outputs(1324)) xor (layer1_outputs(9449));
    layer2_outputs(3032) <= not(layer1_outputs(7421)) or (layer1_outputs(3700));
    layer2_outputs(3033) <= not((layer1_outputs(1891)) xor (layer1_outputs(7381)));
    layer2_outputs(3034) <= not(layer1_outputs(2017));
    layer2_outputs(3035) <= not(layer1_outputs(7949));
    layer2_outputs(3036) <= (layer1_outputs(1767)) and not (layer1_outputs(7770));
    layer2_outputs(3037) <= not(layer1_outputs(531));
    layer2_outputs(3038) <= (layer1_outputs(1664)) and (layer1_outputs(7157));
    layer2_outputs(3039) <= not(layer1_outputs(2766)) or (layer1_outputs(1498));
    layer2_outputs(3040) <= not(layer1_outputs(5635)) or (layer1_outputs(8339));
    layer2_outputs(3041) <= not(layer1_outputs(4096)) or (layer1_outputs(5343));
    layer2_outputs(3042) <= not(layer1_outputs(1636));
    layer2_outputs(3043) <= not(layer1_outputs(7935));
    layer2_outputs(3044) <= not(layer1_outputs(7953)) or (layer1_outputs(1054));
    layer2_outputs(3045) <= not((layer1_outputs(2035)) and (layer1_outputs(7015)));
    layer2_outputs(3046) <= (layer1_outputs(3673)) xor (layer1_outputs(8060));
    layer2_outputs(3047) <= layer1_outputs(9018);
    layer2_outputs(3048) <= not(layer1_outputs(6381));
    layer2_outputs(3049) <= not((layer1_outputs(6649)) and (layer1_outputs(7233)));
    layer2_outputs(3050) <= '0';
    layer2_outputs(3051) <= '0';
    layer2_outputs(3052) <= not((layer1_outputs(3650)) or (layer1_outputs(7607)));
    layer2_outputs(3053) <= (layer1_outputs(6711)) and not (layer1_outputs(1766));
    layer2_outputs(3054) <= not(layer1_outputs(2604));
    layer2_outputs(3055) <= layer1_outputs(9245);
    layer2_outputs(3056) <= not(layer1_outputs(1436)) or (layer1_outputs(2170));
    layer2_outputs(3057) <= layer1_outputs(1317);
    layer2_outputs(3058) <= not(layer1_outputs(7602)) or (layer1_outputs(5605));
    layer2_outputs(3059) <= (layer1_outputs(778)) xor (layer1_outputs(245));
    layer2_outputs(3060) <= not((layer1_outputs(5488)) xor (layer1_outputs(3909)));
    layer2_outputs(3061) <= not(layer1_outputs(9714));
    layer2_outputs(3062) <= layer1_outputs(1300);
    layer2_outputs(3063) <= '1';
    layer2_outputs(3064) <= not((layer1_outputs(7550)) and (layer1_outputs(6849)));
    layer2_outputs(3065) <= not(layer1_outputs(1081)) or (layer1_outputs(5733));
    layer2_outputs(3066) <= layer1_outputs(1294);
    layer2_outputs(3067) <= layer1_outputs(4535);
    layer2_outputs(3068) <= not((layer1_outputs(5274)) xor (layer1_outputs(10135)));
    layer2_outputs(3069) <= not((layer1_outputs(8236)) xor (layer1_outputs(6367)));
    layer2_outputs(3070) <= not(layer1_outputs(7164));
    layer2_outputs(3071) <= not((layer1_outputs(5820)) or (layer1_outputs(3298)));
    layer2_outputs(3072) <= (layer1_outputs(5820)) or (layer1_outputs(796));
    layer2_outputs(3073) <= layer1_outputs(4337);
    layer2_outputs(3074) <= not((layer1_outputs(4784)) and (layer1_outputs(4126)));
    layer2_outputs(3075) <= (layer1_outputs(4829)) and not (layer1_outputs(1218));
    layer2_outputs(3076) <= not((layer1_outputs(9986)) or (layer1_outputs(6211)));
    layer2_outputs(3077) <= not(layer1_outputs(4622)) or (layer1_outputs(7411));
    layer2_outputs(3078) <= (layer1_outputs(7937)) and not (layer1_outputs(4981));
    layer2_outputs(3079) <= not((layer1_outputs(8356)) and (layer1_outputs(4897)));
    layer2_outputs(3080) <= (layer1_outputs(6122)) and not (layer1_outputs(9248));
    layer2_outputs(3081) <= not((layer1_outputs(9689)) and (layer1_outputs(828)));
    layer2_outputs(3082) <= layer1_outputs(4864);
    layer2_outputs(3083) <= '1';
    layer2_outputs(3084) <= not((layer1_outputs(3044)) or (layer1_outputs(5947)));
    layer2_outputs(3085) <= '1';
    layer2_outputs(3086) <= not(layer1_outputs(5409));
    layer2_outputs(3087) <= layer1_outputs(6537);
    layer2_outputs(3088) <= not(layer1_outputs(5252)) or (layer1_outputs(9813));
    layer2_outputs(3089) <= not((layer1_outputs(3604)) or (layer1_outputs(5070)));
    layer2_outputs(3090) <= (layer1_outputs(2)) or (layer1_outputs(5218));
    layer2_outputs(3091) <= not((layer1_outputs(54)) or (layer1_outputs(6392)));
    layer2_outputs(3092) <= not(layer1_outputs(6612)) or (layer1_outputs(6242));
    layer2_outputs(3093) <= (layer1_outputs(5889)) and not (layer1_outputs(8475));
    layer2_outputs(3094) <= not((layer1_outputs(9663)) or (layer1_outputs(1976)));
    layer2_outputs(3095) <= not((layer1_outputs(2931)) or (layer1_outputs(9319)));
    layer2_outputs(3096) <= (layer1_outputs(8747)) and not (layer1_outputs(10070));
    layer2_outputs(3097) <= (layer1_outputs(3975)) xor (layer1_outputs(9950));
    layer2_outputs(3098) <= (layer1_outputs(4724)) and not (layer1_outputs(9607));
    layer2_outputs(3099) <= not((layer1_outputs(7993)) xor (layer1_outputs(5261)));
    layer2_outputs(3100) <= not((layer1_outputs(1039)) and (layer1_outputs(1126)));
    layer2_outputs(3101) <= not(layer1_outputs(9427)) or (layer1_outputs(9784));
    layer2_outputs(3102) <= layer1_outputs(5162);
    layer2_outputs(3103) <= not(layer1_outputs(9929));
    layer2_outputs(3104) <= (layer1_outputs(4919)) and (layer1_outputs(1012));
    layer2_outputs(3105) <= (layer1_outputs(6161)) and (layer1_outputs(4189));
    layer2_outputs(3106) <= (layer1_outputs(5894)) and (layer1_outputs(6239));
    layer2_outputs(3107) <= not(layer1_outputs(8850));
    layer2_outputs(3108) <= layer1_outputs(8756);
    layer2_outputs(3109) <= layer1_outputs(2069);
    layer2_outputs(3110) <= layer1_outputs(7410);
    layer2_outputs(3111) <= not(layer1_outputs(9370)) or (layer1_outputs(2360));
    layer2_outputs(3112) <= layer1_outputs(9768);
    layer2_outputs(3113) <= layer1_outputs(7927);
    layer2_outputs(3114) <= '1';
    layer2_outputs(3115) <= not(layer1_outputs(2929));
    layer2_outputs(3116) <= layer1_outputs(2389);
    layer2_outputs(3117) <= layer1_outputs(1496);
    layer2_outputs(3118) <= not((layer1_outputs(7773)) and (layer1_outputs(37)));
    layer2_outputs(3119) <= not(layer1_outputs(6252));
    layer2_outputs(3120) <= (layer1_outputs(5981)) and (layer1_outputs(9288));
    layer2_outputs(3121) <= layer1_outputs(1928);
    layer2_outputs(3122) <= not(layer1_outputs(4418)) or (layer1_outputs(5317));
    layer2_outputs(3123) <= layer1_outputs(4104);
    layer2_outputs(3124) <= not((layer1_outputs(7029)) or (layer1_outputs(7861)));
    layer2_outputs(3125) <= not((layer1_outputs(9325)) or (layer1_outputs(793)));
    layer2_outputs(3126) <= not((layer1_outputs(8024)) xor (layer1_outputs(9045)));
    layer2_outputs(3127) <= (layer1_outputs(6920)) and not (layer1_outputs(7384));
    layer2_outputs(3128) <= '1';
    layer2_outputs(3129) <= layer1_outputs(947);
    layer2_outputs(3130) <= (layer1_outputs(6330)) and not (layer1_outputs(616));
    layer2_outputs(3131) <= layer1_outputs(6582);
    layer2_outputs(3132) <= (layer1_outputs(5988)) and (layer1_outputs(7437));
    layer2_outputs(3133) <= not(layer1_outputs(7075));
    layer2_outputs(3134) <= (layer1_outputs(3118)) xor (layer1_outputs(859));
    layer2_outputs(3135) <= (layer1_outputs(9421)) and not (layer1_outputs(6748));
    layer2_outputs(3136) <= layer1_outputs(2200);
    layer2_outputs(3137) <= not((layer1_outputs(3632)) xor (layer1_outputs(5941)));
    layer2_outputs(3138) <= not((layer1_outputs(9241)) or (layer1_outputs(8909)));
    layer2_outputs(3139) <= layer1_outputs(3634);
    layer2_outputs(3140) <= (layer1_outputs(2863)) or (layer1_outputs(4728));
    layer2_outputs(3141) <= not((layer1_outputs(3330)) or (layer1_outputs(4457)));
    layer2_outputs(3142) <= layer1_outputs(10237);
    layer2_outputs(3143) <= not((layer1_outputs(8121)) or (layer1_outputs(4644)));
    layer2_outputs(3144) <= not(layer1_outputs(9101));
    layer2_outputs(3145) <= '0';
    layer2_outputs(3146) <= not(layer1_outputs(6172));
    layer2_outputs(3147) <= not(layer1_outputs(6560));
    layer2_outputs(3148) <= layer1_outputs(2795);
    layer2_outputs(3149) <= not(layer1_outputs(4763));
    layer2_outputs(3150) <= not(layer1_outputs(9258));
    layer2_outputs(3151) <= layer1_outputs(4220);
    layer2_outputs(3152) <= layer1_outputs(9732);
    layer2_outputs(3153) <= not((layer1_outputs(6542)) and (layer1_outputs(8380)));
    layer2_outputs(3154) <= layer1_outputs(8630);
    layer2_outputs(3155) <= layer1_outputs(3676);
    layer2_outputs(3156) <= (layer1_outputs(7888)) or (layer1_outputs(9771));
    layer2_outputs(3157) <= not(layer1_outputs(679));
    layer2_outputs(3158) <= not((layer1_outputs(2078)) or (layer1_outputs(6840)));
    layer2_outputs(3159) <= '0';
    layer2_outputs(3160) <= not((layer1_outputs(208)) and (layer1_outputs(9344)));
    layer2_outputs(3161) <= (layer1_outputs(9982)) and (layer1_outputs(1968));
    layer2_outputs(3162) <= not((layer1_outputs(4132)) xor (layer1_outputs(837)));
    layer2_outputs(3163) <= '1';
    layer2_outputs(3164) <= not((layer1_outputs(2512)) and (layer1_outputs(3235)));
    layer2_outputs(3165) <= (layer1_outputs(9430)) and not (layer1_outputs(9965));
    layer2_outputs(3166) <= (layer1_outputs(1388)) and not (layer1_outputs(816));
    layer2_outputs(3167) <= (layer1_outputs(4055)) or (layer1_outputs(9476));
    layer2_outputs(3168) <= not(layer1_outputs(9410)) or (layer1_outputs(9298));
    layer2_outputs(3169) <= (layer1_outputs(7513)) xor (layer1_outputs(3993));
    layer2_outputs(3170) <= (layer1_outputs(9894)) and not (layer1_outputs(5093));
    layer2_outputs(3171) <= '0';
    layer2_outputs(3172) <= (layer1_outputs(3387)) and not (layer1_outputs(3173));
    layer2_outputs(3173) <= not(layer1_outputs(2456));
    layer2_outputs(3174) <= not(layer1_outputs(3214));
    layer2_outputs(3175) <= not((layer1_outputs(3420)) or (layer1_outputs(7640)));
    layer2_outputs(3176) <= layer1_outputs(2180);
    layer2_outputs(3177) <= not(layer1_outputs(2471));
    layer2_outputs(3178) <= not(layer1_outputs(6356));
    layer2_outputs(3179) <= layer1_outputs(393);
    layer2_outputs(3180) <= layer1_outputs(88);
    layer2_outputs(3181) <= not(layer1_outputs(3146));
    layer2_outputs(3182) <= layer1_outputs(2788);
    layer2_outputs(3183) <= not(layer1_outputs(3480));
    layer2_outputs(3184) <= layer1_outputs(8489);
    layer2_outputs(3185) <= (layer1_outputs(5185)) and not (layer1_outputs(3818));
    layer2_outputs(3186) <= not(layer1_outputs(6723));
    layer2_outputs(3187) <= not(layer1_outputs(1989)) or (layer1_outputs(1137));
    layer2_outputs(3188) <= not(layer1_outputs(1380));
    layer2_outputs(3189) <= not(layer1_outputs(9972));
    layer2_outputs(3190) <= not(layer1_outputs(9163));
    layer2_outputs(3191) <= not((layer1_outputs(7213)) and (layer1_outputs(8000)));
    layer2_outputs(3192) <= not(layer1_outputs(7168));
    layer2_outputs(3193) <= (layer1_outputs(2700)) and not (layer1_outputs(6547));
    layer2_outputs(3194) <= layer1_outputs(6150);
    layer2_outputs(3195) <= (layer1_outputs(6521)) and not (layer1_outputs(3344));
    layer2_outputs(3196) <= layer1_outputs(5896);
    layer2_outputs(3197) <= (layer1_outputs(7886)) and not (layer1_outputs(3430));
    layer2_outputs(3198) <= (layer1_outputs(6351)) or (layer1_outputs(10115));
    layer2_outputs(3199) <= not((layer1_outputs(4700)) and (layer1_outputs(1945)));
    layer2_outputs(3200) <= not(layer1_outputs(8943));
    layer2_outputs(3201) <= not(layer1_outputs(9243)) or (layer1_outputs(6868));
    layer2_outputs(3202) <= (layer1_outputs(9708)) and (layer1_outputs(10012));
    layer2_outputs(3203) <= not((layer1_outputs(1510)) or (layer1_outputs(8123)));
    layer2_outputs(3204) <= not(layer1_outputs(2329));
    layer2_outputs(3205) <= not((layer1_outputs(7450)) and (layer1_outputs(2212)));
    layer2_outputs(3206) <= '1';
    layer2_outputs(3207) <= not(layer1_outputs(1459)) or (layer1_outputs(8776));
    layer2_outputs(3208) <= layer1_outputs(682);
    layer2_outputs(3209) <= (layer1_outputs(2245)) or (layer1_outputs(3136));
    layer2_outputs(3210) <= '1';
    layer2_outputs(3211) <= not((layer1_outputs(6422)) or (layer1_outputs(6128)));
    layer2_outputs(3212) <= not(layer1_outputs(6256));
    layer2_outputs(3213) <= layer1_outputs(7660);
    layer2_outputs(3214) <= not((layer1_outputs(4814)) or (layer1_outputs(4403)));
    layer2_outputs(3215) <= layer1_outputs(8457);
    layer2_outputs(3216) <= not(layer1_outputs(4078));
    layer2_outputs(3217) <= layer1_outputs(2021);
    layer2_outputs(3218) <= not((layer1_outputs(5338)) or (layer1_outputs(10179)));
    layer2_outputs(3219) <= not((layer1_outputs(3406)) or (layer1_outputs(1856)));
    layer2_outputs(3220) <= '0';
    layer2_outputs(3221) <= not(layer1_outputs(4707));
    layer2_outputs(3222) <= '1';
    layer2_outputs(3223) <= (layer1_outputs(8897)) and not (layer1_outputs(4772));
    layer2_outputs(3224) <= '1';
    layer2_outputs(3225) <= not(layer1_outputs(5333)) or (layer1_outputs(3018));
    layer2_outputs(3226) <= (layer1_outputs(3692)) and (layer1_outputs(938));
    layer2_outputs(3227) <= layer1_outputs(2489);
    layer2_outputs(3228) <= not((layer1_outputs(2643)) and (layer1_outputs(8694)));
    layer2_outputs(3229) <= (layer1_outputs(867)) and not (layer1_outputs(7199));
    layer2_outputs(3230) <= layer1_outputs(4902);
    layer2_outputs(3231) <= layer1_outputs(5543);
    layer2_outputs(3232) <= layer1_outputs(4931);
    layer2_outputs(3233) <= (layer1_outputs(5098)) and not (layer1_outputs(3219));
    layer2_outputs(3234) <= layer1_outputs(4586);
    layer2_outputs(3235) <= not((layer1_outputs(6436)) or (layer1_outputs(8275)));
    layer2_outputs(3236) <= layer1_outputs(688);
    layer2_outputs(3237) <= not((layer1_outputs(3734)) or (layer1_outputs(4026)));
    layer2_outputs(3238) <= layer1_outputs(4986);
    layer2_outputs(3239) <= not((layer1_outputs(291)) or (layer1_outputs(6771)));
    layer2_outputs(3240) <= (layer1_outputs(3871)) and not (layer1_outputs(4344));
    layer2_outputs(3241) <= layer1_outputs(3995);
    layer2_outputs(3242) <= layer1_outputs(231);
    layer2_outputs(3243) <= '0';
    layer2_outputs(3244) <= (layer1_outputs(3488)) or (layer1_outputs(6344));
    layer2_outputs(3245) <= layer1_outputs(2937);
    layer2_outputs(3246) <= (layer1_outputs(4257)) or (layer1_outputs(6011));
    layer2_outputs(3247) <= not(layer1_outputs(8581));
    layer2_outputs(3248) <= layer1_outputs(791);
    layer2_outputs(3249) <= layer1_outputs(152);
    layer2_outputs(3250) <= not(layer1_outputs(3517));
    layer2_outputs(3251) <= not((layer1_outputs(3151)) or (layer1_outputs(4193)));
    layer2_outputs(3252) <= (layer1_outputs(6145)) and not (layer1_outputs(9526));
    layer2_outputs(3253) <= not(layer1_outputs(4117));
    layer2_outputs(3254) <= layer1_outputs(5223);
    layer2_outputs(3255) <= layer1_outputs(1962);
    layer2_outputs(3256) <= (layer1_outputs(4691)) or (layer1_outputs(9941));
    layer2_outputs(3257) <= layer1_outputs(5129);
    layer2_outputs(3258) <= (layer1_outputs(1127)) and not (layer1_outputs(2468));
    layer2_outputs(3259) <= not(layer1_outputs(4379));
    layer2_outputs(3260) <= (layer1_outputs(7414)) and not (layer1_outputs(2284));
    layer2_outputs(3261) <= not((layer1_outputs(1602)) xor (layer1_outputs(1574)));
    layer2_outputs(3262) <= not(layer1_outputs(2661)) or (layer1_outputs(6791));
    layer2_outputs(3263) <= not(layer1_outputs(4416));
    layer2_outputs(3264) <= (layer1_outputs(7168)) and not (layer1_outputs(8459));
    layer2_outputs(3265) <= not(layer1_outputs(8404)) or (layer1_outputs(7816));
    layer2_outputs(3266) <= layer1_outputs(9944);
    layer2_outputs(3267) <= (layer1_outputs(6075)) and not (layer1_outputs(7692));
    layer2_outputs(3268) <= '0';
    layer2_outputs(3269) <= (layer1_outputs(8038)) and (layer1_outputs(3352));
    layer2_outputs(3270) <= not(layer1_outputs(8651));
    layer2_outputs(3271) <= (layer1_outputs(6739)) or (layer1_outputs(2451));
    layer2_outputs(3272) <= not(layer1_outputs(3847));
    layer2_outputs(3273) <= not(layer1_outputs(4239));
    layer2_outputs(3274) <= (layer1_outputs(3618)) or (layer1_outputs(4514));
    layer2_outputs(3275) <= not(layer1_outputs(7811));
    layer2_outputs(3276) <= (layer1_outputs(8837)) and (layer1_outputs(4750));
    layer2_outputs(3277) <= not((layer1_outputs(4888)) and (layer1_outputs(325)));
    layer2_outputs(3278) <= (layer1_outputs(6754)) or (layer1_outputs(7895));
    layer2_outputs(3279) <= not((layer1_outputs(1910)) and (layer1_outputs(6764)));
    layer2_outputs(3280) <= (layer1_outputs(10077)) and (layer1_outputs(6322));
    layer2_outputs(3281) <= layer1_outputs(6613);
    layer2_outputs(3282) <= (layer1_outputs(5159)) and not (layer1_outputs(2135));
    layer2_outputs(3283) <= (layer1_outputs(9048)) or (layer1_outputs(3070));
    layer2_outputs(3284) <= not(layer1_outputs(2637));
    layer2_outputs(3285) <= layer1_outputs(8414);
    layer2_outputs(3286) <= not(layer1_outputs(9461)) or (layer1_outputs(4561));
    layer2_outputs(3287) <= (layer1_outputs(697)) and not (layer1_outputs(2818));
    layer2_outputs(3288) <= not(layer1_outputs(9290));
    layer2_outputs(3289) <= (layer1_outputs(5865)) and (layer1_outputs(7151));
    layer2_outputs(3290) <= not(layer1_outputs(8109));
    layer2_outputs(3291) <= not(layer1_outputs(9455));
    layer2_outputs(3292) <= (layer1_outputs(9995)) xor (layer1_outputs(3750));
    layer2_outputs(3293) <= (layer1_outputs(5823)) or (layer1_outputs(4933));
    layer2_outputs(3294) <= layer1_outputs(8179);
    layer2_outputs(3295) <= not((layer1_outputs(9994)) or (layer1_outputs(9192)));
    layer2_outputs(3296) <= not(layer1_outputs(9571));
    layer2_outputs(3297) <= layer1_outputs(3374);
    layer2_outputs(3298) <= layer1_outputs(3838);
    layer2_outputs(3299) <= not(layer1_outputs(322));
    layer2_outputs(3300) <= not((layer1_outputs(7162)) and (layer1_outputs(5957)));
    layer2_outputs(3301) <= '1';
    layer2_outputs(3302) <= not(layer1_outputs(2033)) or (layer1_outputs(2400));
    layer2_outputs(3303) <= not((layer1_outputs(1651)) or (layer1_outputs(1657)));
    layer2_outputs(3304) <= not(layer1_outputs(6549));
    layer2_outputs(3305) <= (layer1_outputs(7092)) and not (layer1_outputs(8291));
    layer2_outputs(3306) <= '0';
    layer2_outputs(3307) <= '0';
    layer2_outputs(3308) <= not((layer1_outputs(10193)) or (layer1_outputs(3822)));
    layer2_outputs(3309) <= layer1_outputs(2044);
    layer2_outputs(3310) <= '1';
    layer2_outputs(3311) <= not((layer1_outputs(728)) or (layer1_outputs(7082)));
    layer2_outputs(3312) <= (layer1_outputs(4005)) xor (layer1_outputs(5161));
    layer2_outputs(3313) <= not(layer1_outputs(3591)) or (layer1_outputs(8680));
    layer2_outputs(3314) <= not(layer1_outputs(549));
    layer2_outputs(3315) <= (layer1_outputs(598)) and not (layer1_outputs(3755));
    layer2_outputs(3316) <= not(layer1_outputs(9349));
    layer2_outputs(3317) <= not(layer1_outputs(922));
    layer2_outputs(3318) <= not((layer1_outputs(680)) or (layer1_outputs(4600)));
    layer2_outputs(3319) <= (layer1_outputs(5300)) and not (layer1_outputs(4438));
    layer2_outputs(3320) <= (layer1_outputs(8860)) or (layer1_outputs(5710));
    layer2_outputs(3321) <= not(layer1_outputs(9534)) or (layer1_outputs(8252));
    layer2_outputs(3322) <= '1';
    layer2_outputs(3323) <= layer1_outputs(7254);
    layer2_outputs(3324) <= layer1_outputs(5532);
    layer2_outputs(3325) <= not(layer1_outputs(401));
    layer2_outputs(3326) <= not((layer1_outputs(10235)) or (layer1_outputs(2444)));
    layer2_outputs(3327) <= not(layer1_outputs(3341));
    layer2_outputs(3328) <= (layer1_outputs(3173)) and (layer1_outputs(10076));
    layer2_outputs(3329) <= '1';
    layer2_outputs(3330) <= not((layer1_outputs(5502)) or (layer1_outputs(8352)));
    layer2_outputs(3331) <= layer1_outputs(10226);
    layer2_outputs(3332) <= layer1_outputs(4376);
    layer2_outputs(3333) <= not(layer1_outputs(8522)) or (layer1_outputs(8488));
    layer2_outputs(3334) <= layer1_outputs(1456);
    layer2_outputs(3335) <= layer1_outputs(761);
    layer2_outputs(3336) <= layer1_outputs(737);
    layer2_outputs(3337) <= not(layer1_outputs(571));
    layer2_outputs(3338) <= not((layer1_outputs(3331)) or (layer1_outputs(1589)));
    layer2_outputs(3339) <= (layer1_outputs(5000)) or (layer1_outputs(2046));
    layer2_outputs(3340) <= not(layer1_outputs(9662));
    layer2_outputs(3341) <= '1';
    layer2_outputs(3342) <= (layer1_outputs(7768)) and not (layer1_outputs(8397));
    layer2_outputs(3343) <= not((layer1_outputs(458)) xor (layer1_outputs(3602)));
    layer2_outputs(3344) <= layer1_outputs(7124);
    layer2_outputs(3345) <= not(layer1_outputs(6916));
    layer2_outputs(3346) <= not(layer1_outputs(6232));
    layer2_outputs(3347) <= (layer1_outputs(5830)) and not (layer1_outputs(4223));
    layer2_outputs(3348) <= (layer1_outputs(9389)) and (layer1_outputs(8882));
    layer2_outputs(3349) <= '0';
    layer2_outputs(3350) <= not(layer1_outputs(7430));
    layer2_outputs(3351) <= layer1_outputs(5425);
    layer2_outputs(3352) <= layer1_outputs(1106);
    layer2_outputs(3353) <= layer1_outputs(3825);
    layer2_outputs(3354) <= (layer1_outputs(2244)) and (layer1_outputs(5501));
    layer2_outputs(3355) <= (layer1_outputs(3537)) and not (layer1_outputs(8518));
    layer2_outputs(3356) <= (layer1_outputs(3810)) and not (layer1_outputs(7970));
    layer2_outputs(3357) <= layer1_outputs(10000);
    layer2_outputs(3358) <= not((layer1_outputs(9718)) and (layer1_outputs(8469)));
    layer2_outputs(3359) <= not((layer1_outputs(418)) and (layer1_outputs(7458)));
    layer2_outputs(3360) <= not(layer1_outputs(1777));
    layer2_outputs(3361) <= not((layer1_outputs(89)) or (layer1_outputs(997)));
    layer2_outputs(3362) <= not(layer1_outputs(7603)) or (layer1_outputs(6391));
    layer2_outputs(3363) <= not(layer1_outputs(579)) or (layer1_outputs(10039));
    layer2_outputs(3364) <= not(layer1_outputs(8584)) or (layer1_outputs(2457));
    layer2_outputs(3365) <= not(layer1_outputs(6905)) or (layer1_outputs(4526));
    layer2_outputs(3366) <= '0';
    layer2_outputs(3367) <= not(layer1_outputs(2867));
    layer2_outputs(3368) <= not(layer1_outputs(8116)) or (layer1_outputs(3713));
    layer2_outputs(3369) <= (layer1_outputs(6036)) and not (layer1_outputs(8075));
    layer2_outputs(3370) <= (layer1_outputs(1164)) or (layer1_outputs(823));
    layer2_outputs(3371) <= not(layer1_outputs(8693));
    layer2_outputs(3372) <= not((layer1_outputs(4296)) xor (layer1_outputs(1287)));
    layer2_outputs(3373) <= not((layer1_outputs(3989)) and (layer1_outputs(1564)));
    layer2_outputs(3374) <= not(layer1_outputs(1478));
    layer2_outputs(3375) <= (layer1_outputs(2841)) and not (layer1_outputs(9557));
    layer2_outputs(3376) <= '1';
    layer2_outputs(3377) <= not(layer1_outputs(8783));
    layer2_outputs(3378) <= layer1_outputs(10219);
    layer2_outputs(3379) <= not(layer1_outputs(7253)) or (layer1_outputs(2074));
    layer2_outputs(3380) <= layer1_outputs(3950);
    layer2_outputs(3381) <= layer1_outputs(4880);
    layer2_outputs(3382) <= '1';
    layer2_outputs(3383) <= (layer1_outputs(4624)) and not (layer1_outputs(4676));
    layer2_outputs(3384) <= not(layer1_outputs(0));
    layer2_outputs(3385) <= layer1_outputs(1229);
    layer2_outputs(3386) <= layer1_outputs(9548);
    layer2_outputs(3387) <= (layer1_outputs(1916)) and not (layer1_outputs(5468));
    layer2_outputs(3388) <= (layer1_outputs(9549)) and (layer1_outputs(4333));
    layer2_outputs(3389) <= not(layer1_outputs(3806));
    layer2_outputs(3390) <= not(layer1_outputs(3442)) or (layer1_outputs(7282));
    layer2_outputs(3391) <= '0';
    layer2_outputs(3392) <= layer1_outputs(5382);
    layer2_outputs(3393) <= (layer1_outputs(1520)) and not (layer1_outputs(4699));
    layer2_outputs(3394) <= layer1_outputs(6033);
    layer2_outputs(3395) <= not((layer1_outputs(3660)) or (layer1_outputs(3324)));
    layer2_outputs(3396) <= layer1_outputs(5483);
    layer2_outputs(3397) <= (layer1_outputs(5380)) xor (layer1_outputs(4191));
    layer2_outputs(3398) <= not(layer1_outputs(6962));
    layer2_outputs(3399) <= (layer1_outputs(2728)) and not (layer1_outputs(5264));
    layer2_outputs(3400) <= not(layer1_outputs(884));
    layer2_outputs(3401) <= (layer1_outputs(4240)) and (layer1_outputs(6139));
    layer2_outputs(3402) <= (layer1_outputs(7170)) and not (layer1_outputs(7225));
    layer2_outputs(3403) <= (layer1_outputs(7683)) and not (layer1_outputs(9333));
    layer2_outputs(3404) <= layer1_outputs(6005);
    layer2_outputs(3405) <= layer1_outputs(8041);
    layer2_outputs(3406) <= not((layer1_outputs(3427)) or (layer1_outputs(6069)));
    layer2_outputs(3407) <= layer1_outputs(412);
    layer2_outputs(3408) <= not(layer1_outputs(7865)) or (layer1_outputs(3884));
    layer2_outputs(3409) <= not(layer1_outputs(6013));
    layer2_outputs(3410) <= layer1_outputs(5290);
    layer2_outputs(3411) <= not(layer1_outputs(1562));
    layer2_outputs(3412) <= (layer1_outputs(1158)) xor (layer1_outputs(6446));
    layer2_outputs(3413) <= (layer1_outputs(8829)) and not (layer1_outputs(7640));
    layer2_outputs(3414) <= (layer1_outputs(7828)) and not (layer1_outputs(7785));
    layer2_outputs(3415) <= not(layer1_outputs(8372)) or (layer1_outputs(6321));
    layer2_outputs(3416) <= not(layer1_outputs(314));
    layer2_outputs(3417) <= (layer1_outputs(768)) and (layer1_outputs(8653));
    layer2_outputs(3418) <= not(layer1_outputs(9521));
    layer2_outputs(3419) <= not(layer1_outputs(2210));
    layer2_outputs(3420) <= not(layer1_outputs(547)) or (layer1_outputs(4181));
    layer2_outputs(3421) <= not(layer1_outputs(2320));
    layer2_outputs(3422) <= not((layer1_outputs(1679)) and (layer1_outputs(2501)));
    layer2_outputs(3423) <= (layer1_outputs(7375)) or (layer1_outputs(7220));
    layer2_outputs(3424) <= layer1_outputs(3660);
    layer2_outputs(3425) <= layer1_outputs(7513);
    layer2_outputs(3426) <= not((layer1_outputs(5636)) or (layer1_outputs(6524)));
    layer2_outputs(3427) <= (layer1_outputs(20)) and not (layer1_outputs(9306));
    layer2_outputs(3428) <= '0';
    layer2_outputs(3429) <= (layer1_outputs(4440)) xor (layer1_outputs(2274));
    layer2_outputs(3430) <= (layer1_outputs(8235)) or (layer1_outputs(3363));
    layer2_outputs(3431) <= not(layer1_outputs(9784));
    layer2_outputs(3432) <= not((layer1_outputs(4688)) xor (layer1_outputs(1953)));
    layer2_outputs(3433) <= (layer1_outputs(5603)) or (layer1_outputs(9996));
    layer2_outputs(3434) <= not(layer1_outputs(4509));
    layer2_outputs(3435) <= (layer1_outputs(5325)) and not (layer1_outputs(4665));
    layer2_outputs(3436) <= not(layer1_outputs(204)) or (layer1_outputs(3851));
    layer2_outputs(3437) <= layer1_outputs(5435);
    layer2_outputs(3438) <= (layer1_outputs(2004)) and (layer1_outputs(7911));
    layer2_outputs(3439) <= not(layer1_outputs(7030));
    layer2_outputs(3440) <= layer1_outputs(4376);
    layer2_outputs(3441) <= not((layer1_outputs(7006)) and (layer1_outputs(141)));
    layer2_outputs(3442) <= (layer1_outputs(7264)) and not (layer1_outputs(2814));
    layer2_outputs(3443) <= layer1_outputs(7595);
    layer2_outputs(3444) <= not((layer1_outputs(5721)) xor (layer1_outputs(9461)));
    layer2_outputs(3445) <= (layer1_outputs(4744)) and not (layer1_outputs(5485));
    layer2_outputs(3446) <= not(layer1_outputs(5547));
    layer2_outputs(3447) <= not(layer1_outputs(10203));
    layer2_outputs(3448) <= not((layer1_outputs(8215)) xor (layer1_outputs(3721)));
    layer2_outputs(3449) <= layer1_outputs(4952);
    layer2_outputs(3450) <= (layer1_outputs(6166)) and (layer1_outputs(2915));
    layer2_outputs(3451) <= not(layer1_outputs(8787));
    layer2_outputs(3452) <= not(layer1_outputs(5441));
    layer2_outputs(3453) <= not(layer1_outputs(3422)) or (layer1_outputs(6534));
    layer2_outputs(3454) <= not((layer1_outputs(2174)) and (layer1_outputs(278)));
    layer2_outputs(3455) <= '1';
    layer2_outputs(3456) <= not(layer1_outputs(4072));
    layer2_outputs(3457) <= not(layer1_outputs(6660)) or (layer1_outputs(7099));
    layer2_outputs(3458) <= '1';
    layer2_outputs(3459) <= (layer1_outputs(901)) and (layer1_outputs(5854));
    layer2_outputs(3460) <= layer1_outputs(2092);
    layer2_outputs(3461) <= '1';
    layer2_outputs(3462) <= not((layer1_outputs(8105)) and (layer1_outputs(4508)));
    layer2_outputs(3463) <= layer1_outputs(4507);
    layer2_outputs(3464) <= not((layer1_outputs(2172)) xor (layer1_outputs(6361)));
    layer2_outputs(3465) <= layer1_outputs(4913);
    layer2_outputs(3466) <= not(layer1_outputs(4525));
    layer2_outputs(3467) <= not(layer1_outputs(3949)) or (layer1_outputs(967));
    layer2_outputs(3468) <= not((layer1_outputs(6683)) or (layer1_outputs(3434)));
    layer2_outputs(3469) <= '0';
    layer2_outputs(3470) <= not(layer1_outputs(3927));
    layer2_outputs(3471) <= not(layer1_outputs(9984)) or (layer1_outputs(8151));
    layer2_outputs(3472) <= (layer1_outputs(4884)) and (layer1_outputs(648));
    layer2_outputs(3473) <= not(layer1_outputs(8891)) or (layer1_outputs(6096));
    layer2_outputs(3474) <= not(layer1_outputs(4438));
    layer2_outputs(3475) <= not(layer1_outputs(6243)) or (layer1_outputs(1817));
    layer2_outputs(3476) <= (layer1_outputs(2918)) or (layer1_outputs(7689));
    layer2_outputs(3477) <= layer1_outputs(5405);
    layer2_outputs(3478) <= (layer1_outputs(7296)) or (layer1_outputs(1561));
    layer2_outputs(3479) <= (layer1_outputs(7214)) and not (layer1_outputs(7612));
    layer2_outputs(3480) <= not((layer1_outputs(5829)) and (layer1_outputs(6506)));
    layer2_outputs(3481) <= not((layer1_outputs(7650)) and (layer1_outputs(8438)));
    layer2_outputs(3482) <= not(layer1_outputs(1194));
    layer2_outputs(3483) <= not((layer1_outputs(9124)) and (layer1_outputs(8365)));
    layer2_outputs(3484) <= not((layer1_outputs(8941)) xor (layer1_outputs(2663)));
    layer2_outputs(3485) <= (layer1_outputs(2867)) and not (layer1_outputs(7118));
    layer2_outputs(3486) <= (layer1_outputs(87)) and not (layer1_outputs(5377));
    layer2_outputs(3487) <= (layer1_outputs(2985)) and not (layer1_outputs(4756));
    layer2_outputs(3488) <= not((layer1_outputs(9372)) and (layer1_outputs(8704)));
    layer2_outputs(3489) <= layer1_outputs(4386);
    layer2_outputs(3490) <= (layer1_outputs(2707)) xor (layer1_outputs(537));
    layer2_outputs(3491) <= layer1_outputs(756);
    layer2_outputs(3492) <= '1';
    layer2_outputs(3493) <= layer1_outputs(6117);
    layer2_outputs(3494) <= not((layer1_outputs(7370)) and (layer1_outputs(702)));
    layer2_outputs(3495) <= (layer1_outputs(8859)) xor (layer1_outputs(9667));
    layer2_outputs(3496) <= not((layer1_outputs(2481)) and (layer1_outputs(986)));
    layer2_outputs(3497) <= (layer1_outputs(7838)) and not (layer1_outputs(4318));
    layer2_outputs(3498) <= (layer1_outputs(7488)) and not (layer1_outputs(1523));
    layer2_outputs(3499) <= not(layer1_outputs(4965)) or (layer1_outputs(6094));
    layer2_outputs(3500) <= not(layer1_outputs(6412)) or (layer1_outputs(8745));
    layer2_outputs(3501) <= (layer1_outputs(8441)) and (layer1_outputs(5757));
    layer2_outputs(3502) <= not(layer1_outputs(5952));
    layer2_outputs(3503) <= (layer1_outputs(4711)) or (layer1_outputs(3688));
    layer2_outputs(3504) <= layer1_outputs(2886);
    layer2_outputs(3505) <= (layer1_outputs(6063)) and not (layer1_outputs(2349));
    layer2_outputs(3506) <= (layer1_outputs(8173)) and not (layer1_outputs(7779));
    layer2_outputs(3507) <= not(layer1_outputs(4787)) or (layer1_outputs(8331));
    layer2_outputs(3508) <= layer1_outputs(2462);
    layer2_outputs(3509) <= '0';
    layer2_outputs(3510) <= (layer1_outputs(3915)) and (layer1_outputs(2973));
    layer2_outputs(3511) <= '0';
    layer2_outputs(3512) <= not(layer1_outputs(9636)) or (layer1_outputs(2255));
    layer2_outputs(3513) <= (layer1_outputs(1193)) and not (layer1_outputs(7647));
    layer2_outputs(3514) <= layer1_outputs(3225);
    layer2_outputs(3515) <= (layer1_outputs(6442)) or (layer1_outputs(4224));
    layer2_outputs(3516) <= layer1_outputs(3485);
    layer2_outputs(3517) <= not(layer1_outputs(10165)) or (layer1_outputs(1268));
    layer2_outputs(3518) <= '1';
    layer2_outputs(3519) <= not((layer1_outputs(5633)) and (layer1_outputs(9837)));
    layer2_outputs(3520) <= layer1_outputs(4033);
    layer2_outputs(3521) <= layer1_outputs(33);
    layer2_outputs(3522) <= not((layer1_outputs(673)) and (layer1_outputs(1637)));
    layer2_outputs(3523) <= not(layer1_outputs(8064));
    layer2_outputs(3524) <= not(layer1_outputs(8558));
    layer2_outputs(3525) <= (layer1_outputs(6271)) or (layer1_outputs(4390));
    layer2_outputs(3526) <= not(layer1_outputs(5742));
    layer2_outputs(3527) <= layer1_outputs(8432);
    layer2_outputs(3528) <= not(layer1_outputs(9808)) or (layer1_outputs(4175));
    layer2_outputs(3529) <= layer1_outputs(6159);
    layer2_outputs(3530) <= (layer1_outputs(5763)) or (layer1_outputs(408));
    layer2_outputs(3531) <= not(layer1_outputs(5999));
    layer2_outputs(3532) <= not(layer1_outputs(1554));
    layer2_outputs(3533) <= layer1_outputs(7706);
    layer2_outputs(3534) <= not((layer1_outputs(7348)) xor (layer1_outputs(2190)));
    layer2_outputs(3535) <= not((layer1_outputs(10095)) and (layer1_outputs(145)));
    layer2_outputs(3536) <= '1';
    layer2_outputs(3537) <= '1';
    layer2_outputs(3538) <= layer1_outputs(9823);
    layer2_outputs(3539) <= not(layer1_outputs(380)) or (layer1_outputs(6951));
    layer2_outputs(3540) <= not((layer1_outputs(6120)) xor (layer1_outputs(8980)));
    layer2_outputs(3541) <= not(layer1_outputs(1138));
    layer2_outputs(3542) <= (layer1_outputs(6215)) and not (layer1_outputs(6502));
    layer2_outputs(3543) <= (layer1_outputs(29)) or (layer1_outputs(8929));
    layer2_outputs(3544) <= layer1_outputs(2581);
    layer2_outputs(3545) <= not(layer1_outputs(444));
    layer2_outputs(3546) <= layer1_outputs(1692);
    layer2_outputs(3547) <= not((layer1_outputs(7086)) and (layer1_outputs(825)));
    layer2_outputs(3548) <= layer1_outputs(3188);
    layer2_outputs(3549) <= layer1_outputs(6146);
    layer2_outputs(3550) <= not((layer1_outputs(128)) xor (layer1_outputs(5463)));
    layer2_outputs(3551) <= layer1_outputs(7594);
    layer2_outputs(3552) <= layer1_outputs(8434);
    layer2_outputs(3553) <= not((layer1_outputs(3177)) xor (layer1_outputs(2220)));
    layer2_outputs(3554) <= not(layer1_outputs(3767)) or (layer1_outputs(2348));
    layer2_outputs(3555) <= (layer1_outputs(3273)) and (layer1_outputs(2923));
    layer2_outputs(3556) <= '0';
    layer2_outputs(3557) <= '1';
    layer2_outputs(3558) <= not(layer1_outputs(812)) or (layer1_outputs(5349));
    layer2_outputs(3559) <= layer1_outputs(6665);
    layer2_outputs(3560) <= not(layer1_outputs(4567)) or (layer1_outputs(4084));
    layer2_outputs(3561) <= not(layer1_outputs(3177)) or (layer1_outputs(2422));
    layer2_outputs(3562) <= (layer1_outputs(8600)) and (layer1_outputs(8700));
    layer2_outputs(3563) <= not(layer1_outputs(3072));
    layer2_outputs(3564) <= not(layer1_outputs(6127));
    layer2_outputs(3565) <= not((layer1_outputs(7106)) and (layer1_outputs(3966)));
    layer2_outputs(3566) <= (layer1_outputs(1759)) xor (layer1_outputs(4046));
    layer2_outputs(3567) <= not(layer1_outputs(3739));
    layer2_outputs(3568) <= (layer1_outputs(9954)) and (layer1_outputs(10064));
    layer2_outputs(3569) <= layer1_outputs(1906);
    layer2_outputs(3570) <= not((layer1_outputs(1134)) or (layer1_outputs(3036)));
    layer2_outputs(3571) <= (layer1_outputs(417)) and not (layer1_outputs(9956));
    layer2_outputs(3572) <= layer1_outputs(1935);
    layer2_outputs(3573) <= not(layer1_outputs(6772));
    layer2_outputs(3574) <= not((layer1_outputs(4244)) or (layer1_outputs(5637)));
    layer2_outputs(3575) <= (layer1_outputs(2833)) xor (layer1_outputs(5440));
    layer2_outputs(3576) <= layer1_outputs(9630);
    layer2_outputs(3577) <= not(layer1_outputs(5130)) or (layer1_outputs(9421));
    layer2_outputs(3578) <= layer1_outputs(600);
    layer2_outputs(3579) <= layer1_outputs(1438);
    layer2_outputs(3580) <= not(layer1_outputs(6055)) or (layer1_outputs(8960));
    layer2_outputs(3581) <= '1';
    layer2_outputs(3582) <= (layer1_outputs(6838)) or (layer1_outputs(10238));
    layer2_outputs(3583) <= not(layer1_outputs(622)) or (layer1_outputs(7247));
    layer2_outputs(3584) <= (layer1_outputs(9505)) or (layer1_outputs(4449));
    layer2_outputs(3585) <= (layer1_outputs(8659)) and not (layer1_outputs(10015));
    layer2_outputs(3586) <= not(layer1_outputs(428));
    layer2_outputs(3587) <= (layer1_outputs(7308)) and not (layer1_outputs(5815));
    layer2_outputs(3588) <= (layer1_outputs(6424)) or (layer1_outputs(7715));
    layer2_outputs(3589) <= not((layer1_outputs(8288)) or (layer1_outputs(10044)));
    layer2_outputs(3590) <= (layer1_outputs(6303)) and not (layer1_outputs(7441));
    layer2_outputs(3591) <= not(layer1_outputs(1237)) or (layer1_outputs(7992));
    layer2_outputs(3592) <= (layer1_outputs(6619)) and not (layer1_outputs(7356));
    layer2_outputs(3593) <= layer1_outputs(6306);
    layer2_outputs(3594) <= layer1_outputs(3035);
    layer2_outputs(3595) <= not(layer1_outputs(5303)) or (layer1_outputs(2576));
    layer2_outputs(3596) <= not((layer1_outputs(2061)) and (layer1_outputs(6144)));
    layer2_outputs(3597) <= not(layer1_outputs(10213)) or (layer1_outputs(6062));
    layer2_outputs(3598) <= not((layer1_outputs(4489)) or (layer1_outputs(2981)));
    layer2_outputs(3599) <= (layer1_outputs(912)) and not (layer1_outputs(8498));
    layer2_outputs(3600) <= not(layer1_outputs(53));
    layer2_outputs(3601) <= (layer1_outputs(5988)) and not (layer1_outputs(1765));
    layer2_outputs(3602) <= layer1_outputs(9812);
    layer2_outputs(3603) <= not(layer1_outputs(9978));
    layer2_outputs(3604) <= layer1_outputs(3464);
    layer2_outputs(3605) <= layer1_outputs(2339);
    layer2_outputs(3606) <= (layer1_outputs(587)) xor (layer1_outputs(1427));
    layer2_outputs(3607) <= '0';
    layer2_outputs(3608) <= (layer1_outputs(4993)) and not (layer1_outputs(6753));
    layer2_outputs(3609) <= (layer1_outputs(4343)) and not (layer1_outputs(1953));
    layer2_outputs(3610) <= not(layer1_outputs(2862));
    layer2_outputs(3611) <= (layer1_outputs(3360)) and not (layer1_outputs(1069));
    layer2_outputs(3612) <= not(layer1_outputs(1062)) or (layer1_outputs(7122));
    layer2_outputs(3613) <= (layer1_outputs(479)) and not (layer1_outputs(647));
    layer2_outputs(3614) <= not(layer1_outputs(9128));
    layer2_outputs(3615) <= (layer1_outputs(7791)) and not (layer1_outputs(868));
    layer2_outputs(3616) <= not((layer1_outputs(1260)) and (layer1_outputs(4720)));
    layer2_outputs(3617) <= layer1_outputs(9976);
    layer2_outputs(3618) <= (layer1_outputs(265)) and not (layer1_outputs(9634));
    layer2_outputs(3619) <= not((layer1_outputs(3378)) or (layer1_outputs(5906)));
    layer2_outputs(3620) <= not(layer1_outputs(4581));
    layer2_outputs(3621) <= (layer1_outputs(1238)) and not (layer1_outputs(9418));
    layer2_outputs(3622) <= (layer1_outputs(929)) and (layer1_outputs(4512));
    layer2_outputs(3623) <= not(layer1_outputs(5255));
    layer2_outputs(3624) <= not((layer1_outputs(8417)) xor (layer1_outputs(9390)));
    layer2_outputs(3625) <= (layer1_outputs(3586)) xor (layer1_outputs(5194));
    layer2_outputs(3626) <= not((layer1_outputs(8363)) and (layer1_outputs(3793)));
    layer2_outputs(3627) <= layer1_outputs(7120);
    layer2_outputs(3628) <= not(layer1_outputs(3077)) or (layer1_outputs(4143));
    layer2_outputs(3629) <= not(layer1_outputs(5138)) or (layer1_outputs(2588));
    layer2_outputs(3630) <= layer1_outputs(5272);
    layer2_outputs(3631) <= not((layer1_outputs(2467)) and (layer1_outputs(6832)));
    layer2_outputs(3632) <= not((layer1_outputs(8055)) and (layer1_outputs(6844)));
    layer2_outputs(3633) <= layer1_outputs(4528);
    layer2_outputs(3634) <= not(layer1_outputs(6994));
    layer2_outputs(3635) <= layer1_outputs(6169);
    layer2_outputs(3636) <= (layer1_outputs(5822)) and not (layer1_outputs(1575));
    layer2_outputs(3637) <= not(layer1_outputs(5172));
    layer2_outputs(3638) <= layer1_outputs(5660);
    layer2_outputs(3639) <= layer1_outputs(1483);
    layer2_outputs(3640) <= (layer1_outputs(4571)) xor (layer1_outputs(6553));
    layer2_outputs(3641) <= not(layer1_outputs(8461)) or (layer1_outputs(3775));
    layer2_outputs(3642) <= not((layer1_outputs(5120)) or (layer1_outputs(8407)));
    layer2_outputs(3643) <= not(layer1_outputs(5109)) or (layer1_outputs(2437));
    layer2_outputs(3644) <= not(layer1_outputs(4724)) or (layer1_outputs(4019));
    layer2_outputs(3645) <= (layer1_outputs(7884)) and (layer1_outputs(2517));
    layer2_outputs(3646) <= (layer1_outputs(5407)) and not (layer1_outputs(808));
    layer2_outputs(3647) <= (layer1_outputs(2202)) and not (layer1_outputs(8662));
    layer2_outputs(3648) <= not((layer1_outputs(3390)) and (layer1_outputs(2156)));
    layer2_outputs(3649) <= not(layer1_outputs(3667));
    layer2_outputs(3650) <= (layer1_outputs(8770)) or (layer1_outputs(7372));
    layer2_outputs(3651) <= layer1_outputs(627);
    layer2_outputs(3652) <= '0';
    layer2_outputs(3653) <= '1';
    layer2_outputs(3654) <= layer1_outputs(2405);
    layer2_outputs(3655) <= (layer1_outputs(2471)) or (layer1_outputs(8780));
    layer2_outputs(3656) <= not(layer1_outputs(5549));
    layer2_outputs(3657) <= not((layer1_outputs(5361)) xor (layer1_outputs(8626)));
    layer2_outputs(3658) <= (layer1_outputs(952)) and not (layer1_outputs(3653));
    layer2_outputs(3659) <= not((layer1_outputs(991)) xor (layer1_outputs(6235)));
    layer2_outputs(3660) <= (layer1_outputs(8068)) and (layer1_outputs(340));
    layer2_outputs(3661) <= (layer1_outputs(383)) xor (layer1_outputs(5919));
    layer2_outputs(3662) <= '0';
    layer2_outputs(3663) <= not(layer1_outputs(7817)) or (layer1_outputs(5372));
    layer2_outputs(3664) <= '0';
    layer2_outputs(3665) <= not((layer1_outputs(8318)) xor (layer1_outputs(6791)));
    layer2_outputs(3666) <= (layer1_outputs(6997)) and not (layer1_outputs(6230));
    layer2_outputs(3667) <= layer1_outputs(2754);
    layer2_outputs(3668) <= layer1_outputs(8036);
    layer2_outputs(3669) <= '0';
    layer2_outputs(3670) <= not(layer1_outputs(7250));
    layer2_outputs(3671) <= layer1_outputs(7716);
    layer2_outputs(3672) <= not(layer1_outputs(1507));
    layer2_outputs(3673) <= (layer1_outputs(4928)) and not (layer1_outputs(6661));
    layer2_outputs(3674) <= layer1_outputs(7790);
    layer2_outputs(3675) <= '1';
    layer2_outputs(3676) <= (layer1_outputs(6820)) xor (layer1_outputs(5403));
    layer2_outputs(3677) <= layer1_outputs(10049);
    layer2_outputs(3678) <= layer1_outputs(3920);
    layer2_outputs(3679) <= (layer1_outputs(1819)) and not (layer1_outputs(2059));
    layer2_outputs(3680) <= not(layer1_outputs(1382));
    layer2_outputs(3681) <= layer1_outputs(8706);
    layer2_outputs(3682) <= (layer1_outputs(8320)) and not (layer1_outputs(3244));
    layer2_outputs(3683) <= layer1_outputs(3482);
    layer2_outputs(3684) <= (layer1_outputs(456)) xor (layer1_outputs(9193));
    layer2_outputs(3685) <= layer1_outputs(9557);
    layer2_outputs(3686) <= (layer1_outputs(2740)) and not (layer1_outputs(840));
    layer2_outputs(3687) <= not(layer1_outputs(8749));
    layer2_outputs(3688) <= (layer1_outputs(386)) or (layer1_outputs(4715));
    layer2_outputs(3689) <= (layer1_outputs(9424)) and (layer1_outputs(8100));
    layer2_outputs(3690) <= (layer1_outputs(212)) and not (layer1_outputs(9146));
    layer2_outputs(3691) <= not(layer1_outputs(1686));
    layer2_outputs(3692) <= not(layer1_outputs(6101)) or (layer1_outputs(6842));
    layer2_outputs(3693) <= (layer1_outputs(6889)) and not (layer1_outputs(689));
    layer2_outputs(3694) <= (layer1_outputs(4358)) and not (layer1_outputs(85));
    layer2_outputs(3695) <= not(layer1_outputs(1927)) or (layer1_outputs(4558));
    layer2_outputs(3696) <= '1';
    layer2_outputs(3697) <= (layer1_outputs(1928)) xor (layer1_outputs(7915));
    layer2_outputs(3698) <= (layer1_outputs(8665)) or (layer1_outputs(2869));
    layer2_outputs(3699) <= (layer1_outputs(3497)) and (layer1_outputs(9789));
    layer2_outputs(3700) <= (layer1_outputs(6422)) xor (layer1_outputs(7158));
    layer2_outputs(3701) <= not((layer1_outputs(3599)) and (layer1_outputs(7530)));
    layer2_outputs(3702) <= layer1_outputs(7254);
    layer2_outputs(3703) <= '0';
    layer2_outputs(3704) <= (layer1_outputs(2066)) or (layer1_outputs(6134));
    layer2_outputs(3705) <= (layer1_outputs(8757)) or (layer1_outputs(4604));
    layer2_outputs(3706) <= layer1_outputs(8212);
    layer2_outputs(3707) <= not((layer1_outputs(2877)) or (layer1_outputs(5400)));
    layer2_outputs(3708) <= layer1_outputs(2737);
    layer2_outputs(3709) <= not(layer1_outputs(2062));
    layer2_outputs(3710) <= not(layer1_outputs(7919));
    layer2_outputs(3711) <= not(layer1_outputs(4603));
    layer2_outputs(3712) <= layer1_outputs(2173);
    layer2_outputs(3713) <= '1';
    layer2_outputs(3714) <= not(layer1_outputs(4210)) or (layer1_outputs(379));
    layer2_outputs(3715) <= not(layer1_outputs(7208));
    layer2_outputs(3716) <= not(layer1_outputs(10035));
    layer2_outputs(3717) <= not(layer1_outputs(1692));
    layer2_outputs(3718) <= layer1_outputs(6138);
    layer2_outputs(3719) <= not((layer1_outputs(7317)) or (layer1_outputs(8191)));
    layer2_outputs(3720) <= layer1_outputs(8986);
    layer2_outputs(3721) <= layer1_outputs(2979);
    layer2_outputs(3722) <= not(layer1_outputs(9322));
    layer2_outputs(3723) <= not(layer1_outputs(3940)) or (layer1_outputs(9167));
    layer2_outputs(3724) <= layer1_outputs(3595);
    layer2_outputs(3725) <= layer1_outputs(3373);
    layer2_outputs(3726) <= '0';
    layer2_outputs(3727) <= not((layer1_outputs(1364)) and (layer1_outputs(1467)));
    layer2_outputs(3728) <= not(layer1_outputs(1807));
    layer2_outputs(3729) <= layer1_outputs(6499);
    layer2_outputs(3730) <= layer1_outputs(7769);
    layer2_outputs(3731) <= layer1_outputs(3815);
    layer2_outputs(3732) <= layer1_outputs(9419);
    layer2_outputs(3733) <= layer1_outputs(2772);
    layer2_outputs(3734) <= not(layer1_outputs(8015)) or (layer1_outputs(3404));
    layer2_outputs(3735) <= (layer1_outputs(8494)) and not (layer1_outputs(4114));
    layer2_outputs(3736) <= layer1_outputs(7393);
    layer2_outputs(3737) <= not(layer1_outputs(4918)) or (layer1_outputs(336));
    layer2_outputs(3738) <= not(layer1_outputs(4801));
    layer2_outputs(3739) <= not((layer1_outputs(3269)) or (layer1_outputs(1546)));
    layer2_outputs(3740) <= layer1_outputs(5983);
    layer2_outputs(3741) <= '0';
    layer2_outputs(3742) <= not(layer1_outputs(6706));
    layer2_outputs(3743) <= layer1_outputs(2181);
    layer2_outputs(3744) <= not(layer1_outputs(2851));
    layer2_outputs(3745) <= layer1_outputs(7105);
    layer2_outputs(3746) <= (layer1_outputs(9996)) and (layer1_outputs(10020));
    layer2_outputs(3747) <= (layer1_outputs(9609)) and (layer1_outputs(6225));
    layer2_outputs(3748) <= not(layer1_outputs(2201));
    layer2_outputs(3749) <= '0';
    layer2_outputs(3750) <= (layer1_outputs(9462)) and (layer1_outputs(5669));
    layer2_outputs(3751) <= not(layer1_outputs(9027));
    layer2_outputs(3752) <= layer1_outputs(4982);
    layer2_outputs(3753) <= not(layer1_outputs(8717));
    layer2_outputs(3754) <= not((layer1_outputs(8362)) or (layer1_outputs(7249)));
    layer2_outputs(3755) <= layer1_outputs(992);
    layer2_outputs(3756) <= layer1_outputs(6620);
    layer2_outputs(3757) <= not((layer1_outputs(9215)) xor (layer1_outputs(4306)));
    layer2_outputs(3758) <= (layer1_outputs(9470)) xor (layer1_outputs(8453));
    layer2_outputs(3759) <= layer1_outputs(9364);
    layer2_outputs(3760) <= not(layer1_outputs(5541)) or (layer1_outputs(2525));
    layer2_outputs(3761) <= layer1_outputs(4611);
    layer2_outputs(3762) <= (layer1_outputs(9291)) and not (layer1_outputs(1820));
    layer2_outputs(3763) <= layer1_outputs(1519);
    layer2_outputs(3764) <= not(layer1_outputs(3928));
    layer2_outputs(3765) <= (layer1_outputs(5168)) and not (layer1_outputs(590));
    layer2_outputs(3766) <= not(layer1_outputs(1325));
    layer2_outputs(3767) <= layer1_outputs(9724);
    layer2_outputs(3768) <= layer1_outputs(7469);
    layer2_outputs(3769) <= not(layer1_outputs(3748));
    layer2_outputs(3770) <= (layer1_outputs(3379)) and (layer1_outputs(9283));
    layer2_outputs(3771) <= layer1_outputs(5777);
    layer2_outputs(3772) <= (layer1_outputs(3897)) and (layer1_outputs(8471));
    layer2_outputs(3773) <= not((layer1_outputs(674)) or (layer1_outputs(3193)));
    layer2_outputs(3774) <= '0';
    layer2_outputs(3775) <= (layer1_outputs(6196)) or (layer1_outputs(7957));
    layer2_outputs(3776) <= not(layer1_outputs(1748)) or (layer1_outputs(7408));
    layer2_outputs(3777) <= layer1_outputs(7525);
    layer2_outputs(3778) <= layer1_outputs(875);
    layer2_outputs(3779) <= layer1_outputs(6319);
    layer2_outputs(3780) <= not(layer1_outputs(5547));
    layer2_outputs(3781) <= not(layer1_outputs(6858)) or (layer1_outputs(5961));
    layer2_outputs(3782) <= (layer1_outputs(9465)) or (layer1_outputs(10153));
    layer2_outputs(3783) <= (layer1_outputs(5878)) or (layer1_outputs(822));
    layer2_outputs(3784) <= not((layer1_outputs(3213)) xor (layer1_outputs(9104)));
    layer2_outputs(3785) <= '0';
    layer2_outputs(3786) <= not((layer1_outputs(5621)) or (layer1_outputs(2072)));
    layer2_outputs(3787) <= not(layer1_outputs(739));
    layer2_outputs(3788) <= layer1_outputs(3850);
    layer2_outputs(3789) <= not(layer1_outputs(7232));
    layer2_outputs(3790) <= not(layer1_outputs(6355));
    layer2_outputs(3791) <= not(layer1_outputs(714));
    layer2_outputs(3792) <= not((layer1_outputs(10195)) and (layer1_outputs(4928)));
    layer2_outputs(3793) <= not(layer1_outputs(2731)) or (layer1_outputs(4778));
    layer2_outputs(3794) <= (layer1_outputs(9881)) and (layer1_outputs(7711));
    layer2_outputs(3795) <= layer1_outputs(856);
    layer2_outputs(3796) <= layer1_outputs(7867);
    layer2_outputs(3797) <= not(layer1_outputs(3684));
    layer2_outputs(3798) <= layer1_outputs(7249);
    layer2_outputs(3799) <= not(layer1_outputs(2121));
    layer2_outputs(3800) <= layer1_outputs(5140);
    layer2_outputs(3801) <= not(layer1_outputs(6181)) or (layer1_outputs(3921));
    layer2_outputs(3802) <= not(layer1_outputs(284)) or (layer1_outputs(2535));
    layer2_outputs(3803) <= (layer1_outputs(4811)) and (layer1_outputs(5710));
    layer2_outputs(3804) <= not((layer1_outputs(3150)) xor (layer1_outputs(2718)));
    layer2_outputs(3805) <= (layer1_outputs(6938)) and not (layer1_outputs(1333));
    layer2_outputs(3806) <= (layer1_outputs(9429)) and not (layer1_outputs(2947));
    layer2_outputs(3807) <= not(layer1_outputs(6287));
    layer2_outputs(3808) <= '1';
    layer2_outputs(3809) <= (layer1_outputs(6985)) and not (layer1_outputs(6057));
    layer2_outputs(3810) <= (layer1_outputs(4755)) and not (layer1_outputs(7323));
    layer2_outputs(3811) <= (layer1_outputs(4586)) xor (layer1_outputs(4871));
    layer2_outputs(3812) <= '1';
    layer2_outputs(3813) <= not(layer1_outputs(6189)) or (layer1_outputs(4651));
    layer2_outputs(3814) <= (layer1_outputs(9992)) and not (layer1_outputs(10193));
    layer2_outputs(3815) <= not(layer1_outputs(4249)) or (layer1_outputs(7465));
    layer2_outputs(3816) <= (layer1_outputs(10139)) and (layer1_outputs(6655));
    layer2_outputs(3817) <= not(layer1_outputs(500));
    layer2_outputs(3818) <= (layer1_outputs(1890)) and not (layer1_outputs(6611));
    layer2_outputs(3819) <= (layer1_outputs(10082)) xor (layer1_outputs(1059));
    layer2_outputs(3820) <= not((layer1_outputs(7870)) and (layer1_outputs(2584)));
    layer2_outputs(3821) <= (layer1_outputs(1771)) xor (layer1_outputs(6066));
    layer2_outputs(3822) <= layer1_outputs(6465);
    layer2_outputs(3823) <= not(layer1_outputs(4412));
    layer2_outputs(3824) <= not(layer1_outputs(3472)) or (layer1_outputs(6238));
    layer2_outputs(3825) <= not((layer1_outputs(148)) and (layer1_outputs(9644)));
    layer2_outputs(3826) <= layer1_outputs(1511);
    layer2_outputs(3827) <= layer1_outputs(9020);
    layer2_outputs(3828) <= '1';
    layer2_outputs(3829) <= not(layer1_outputs(8107));
    layer2_outputs(3830) <= layer1_outputs(5056);
    layer2_outputs(3831) <= '0';
    layer2_outputs(3832) <= layer1_outputs(9511);
    layer2_outputs(3833) <= not((layer1_outputs(4916)) xor (layer1_outputs(8910)));
    layer2_outputs(3834) <= not((layer1_outputs(10065)) or (layer1_outputs(2240)));
    layer2_outputs(3835) <= layer1_outputs(5236);
    layer2_outputs(3836) <= (layer1_outputs(8668)) or (layer1_outputs(9048));
    layer2_outputs(3837) <= (layer1_outputs(1541)) and (layer1_outputs(2594));
    layer2_outputs(3838) <= (layer1_outputs(495)) or (layer1_outputs(6962));
    layer2_outputs(3839) <= not(layer1_outputs(3475));
    layer2_outputs(3840) <= '1';
    layer2_outputs(3841) <= layer1_outputs(2593);
    layer2_outputs(3842) <= layer1_outputs(4223);
    layer2_outputs(3843) <= not(layer1_outputs(4884));
    layer2_outputs(3844) <= layer1_outputs(25);
    layer2_outputs(3845) <= not(layer1_outputs(4060));
    layer2_outputs(3846) <= layer1_outputs(3236);
    layer2_outputs(3847) <= layer1_outputs(8907);
    layer2_outputs(3848) <= (layer1_outputs(1143)) and not (layer1_outputs(8069));
    layer2_outputs(3849) <= layer1_outputs(55);
    layer2_outputs(3850) <= not(layer1_outputs(1849)) or (layer1_outputs(5177));
    layer2_outputs(3851) <= (layer1_outputs(9074)) and not (layer1_outputs(3975));
    layer2_outputs(3852) <= layer1_outputs(3075);
    layer2_outputs(3853) <= not(layer1_outputs(1353)) or (layer1_outputs(5704));
    layer2_outputs(3854) <= (layer1_outputs(9181)) and not (layer1_outputs(1524));
    layer2_outputs(3855) <= not((layer1_outputs(4891)) xor (layer1_outputs(8270)));
    layer2_outputs(3856) <= (layer1_outputs(6602)) and not (layer1_outputs(2630));
    layer2_outputs(3857) <= (layer1_outputs(6890)) or (layer1_outputs(7560));
    layer2_outputs(3858) <= (layer1_outputs(5167)) and (layer1_outputs(2913));
    layer2_outputs(3859) <= not(layer1_outputs(6221));
    layer2_outputs(3860) <= layer1_outputs(1150);
    layer2_outputs(3861) <= '0';
    layer2_outputs(3862) <= (layer1_outputs(4120)) and not (layer1_outputs(1937));
    layer2_outputs(3863) <= '0';
    layer2_outputs(3864) <= layer1_outputs(2417);
    layer2_outputs(3865) <= (layer1_outputs(2519)) or (layer1_outputs(5906));
    layer2_outputs(3866) <= layer1_outputs(9960);
    layer2_outputs(3867) <= not(layer1_outputs(9852)) or (layer1_outputs(9086));
    layer2_outputs(3868) <= layer1_outputs(3462);
    layer2_outputs(3869) <= (layer1_outputs(3720)) and not (layer1_outputs(3232));
    layer2_outputs(3870) <= (layer1_outputs(7951)) xor (layer1_outputs(9602));
    layer2_outputs(3871) <= layer1_outputs(6484);
    layer2_outputs(3872) <= not((layer1_outputs(9256)) and (layer1_outputs(4536)));
    layer2_outputs(3873) <= (layer1_outputs(2182)) and not (layer1_outputs(172));
    layer2_outputs(3874) <= (layer1_outputs(7443)) xor (layer1_outputs(1201));
    layer2_outputs(3875) <= not(layer1_outputs(279));
    layer2_outputs(3876) <= not(layer1_outputs(8897));
    layer2_outputs(3877) <= (layer1_outputs(6751)) and not (layer1_outputs(5580));
    layer2_outputs(3878) <= (layer1_outputs(7897)) xor (layer1_outputs(7575));
    layer2_outputs(3879) <= layer1_outputs(8264);
    layer2_outputs(3880) <= '0';
    layer2_outputs(3881) <= (layer1_outputs(5679)) or (layer1_outputs(599));
    layer2_outputs(3882) <= (layer1_outputs(8381)) and not (layer1_outputs(1339));
    layer2_outputs(3883) <= not((layer1_outputs(1442)) and (layer1_outputs(9532)));
    layer2_outputs(3884) <= not(layer1_outputs(1345));
    layer2_outputs(3885) <= not((layer1_outputs(3979)) or (layer1_outputs(2215)));
    layer2_outputs(3886) <= layer1_outputs(3095);
    layer2_outputs(3887) <= not(layer1_outputs(6040));
    layer2_outputs(3888) <= layer1_outputs(3193);
    layer2_outputs(3889) <= not(layer1_outputs(396)) or (layer1_outputs(5887));
    layer2_outputs(3890) <= layer1_outputs(3276);
    layer2_outputs(3891) <= not(layer1_outputs(3864));
    layer2_outputs(3892) <= (layer1_outputs(1317)) and not (layer1_outputs(4411));
    layer2_outputs(3893) <= layer1_outputs(9317);
    layer2_outputs(3894) <= not(layer1_outputs(1623)) or (layer1_outputs(3554));
    layer2_outputs(3895) <= (layer1_outputs(2378)) and not (layer1_outputs(1868));
    layer2_outputs(3896) <= '0';
    layer2_outputs(3897) <= not(layer1_outputs(1009)) or (layer1_outputs(9919));
    layer2_outputs(3898) <= not((layer1_outputs(242)) or (layer1_outputs(8365)));
    layer2_outputs(3899) <= not((layer1_outputs(5282)) or (layer1_outputs(1733)));
    layer2_outputs(3900) <= layer1_outputs(5287);
    layer2_outputs(3901) <= layer1_outputs(2908);
    layer2_outputs(3902) <= layer1_outputs(3019);
    layer2_outputs(3903) <= layer1_outputs(4993);
    layer2_outputs(3904) <= not(layer1_outputs(8285));
    layer2_outputs(3905) <= (layer1_outputs(1076)) or (layer1_outputs(5093));
    layer2_outputs(3906) <= (layer1_outputs(215)) and not (layer1_outputs(332));
    layer2_outputs(3907) <= not(layer1_outputs(26)) or (layer1_outputs(9002));
    layer2_outputs(3908) <= not(layer1_outputs(4848));
    layer2_outputs(3909) <= not((layer1_outputs(2194)) and (layer1_outputs(6037)));
    layer2_outputs(3910) <= not(layer1_outputs(3795));
    layer2_outputs(3911) <= not(layer1_outputs(8982)) or (layer1_outputs(10201));
    layer2_outputs(3912) <= layer1_outputs(2528);
    layer2_outputs(3913) <= (layer1_outputs(367)) or (layer1_outputs(5596));
    layer2_outputs(3914) <= not((layer1_outputs(8700)) xor (layer1_outputs(7328)));
    layer2_outputs(3915) <= not((layer1_outputs(8451)) and (layer1_outputs(6369)));
    layer2_outputs(3916) <= not(layer1_outputs(7354));
    layer2_outputs(3917) <= not((layer1_outputs(6253)) or (layer1_outputs(7055)));
    layer2_outputs(3918) <= (layer1_outputs(5051)) and (layer1_outputs(7498));
    layer2_outputs(3919) <= layer1_outputs(4773);
    layer2_outputs(3920) <= not(layer1_outputs(7278)) or (layer1_outputs(517));
    layer2_outputs(3921) <= layer1_outputs(9993);
    layer2_outputs(3922) <= not(layer1_outputs(8158));
    layer2_outputs(3923) <= layer1_outputs(6335);
    layer2_outputs(3924) <= (layer1_outputs(4806)) and (layer1_outputs(6804));
    layer2_outputs(3925) <= (layer1_outputs(5388)) xor (layer1_outputs(36));
    layer2_outputs(3926) <= layer1_outputs(7914);
    layer2_outputs(3927) <= (layer1_outputs(3642)) and not (layer1_outputs(10025));
    layer2_outputs(3928) <= not(layer1_outputs(7618));
    layer2_outputs(3929) <= layer1_outputs(3829);
    layer2_outputs(3930) <= layer1_outputs(7230);
    layer2_outputs(3931) <= layer1_outputs(8959);
    layer2_outputs(3932) <= not(layer1_outputs(4625));
    layer2_outputs(3933) <= not(layer1_outputs(8778));
    layer2_outputs(3934) <= not(layer1_outputs(7921));
    layer2_outputs(3935) <= '1';
    layer2_outputs(3936) <= layer1_outputs(8523);
    layer2_outputs(3937) <= not(layer1_outputs(10153)) or (layer1_outputs(5832));
    layer2_outputs(3938) <= layer1_outputs(169);
    layer2_outputs(3939) <= layer1_outputs(2013);
    layer2_outputs(3940) <= not(layer1_outputs(5135)) or (layer1_outputs(3526));
    layer2_outputs(3941) <= layer1_outputs(4395);
    layer2_outputs(3942) <= not((layer1_outputs(2895)) xor (layer1_outputs(10113)));
    layer2_outputs(3943) <= layer1_outputs(4163);
    layer2_outputs(3944) <= not(layer1_outputs(763)) or (layer1_outputs(10021));
    layer2_outputs(3945) <= (layer1_outputs(5741)) xor (layer1_outputs(7522));
    layer2_outputs(3946) <= '1';
    layer2_outputs(3947) <= not((layer1_outputs(1590)) or (layer1_outputs(62)));
    layer2_outputs(3948) <= (layer1_outputs(588)) and (layer1_outputs(7164));
    layer2_outputs(3949) <= '1';
    layer2_outputs(3950) <= (layer1_outputs(2386)) xor (layer1_outputs(1996));
    layer2_outputs(3951) <= not((layer1_outputs(6403)) or (layer1_outputs(5134)));
    layer2_outputs(3952) <= not(layer1_outputs(5846)) or (layer1_outputs(6754));
    layer2_outputs(3953) <= not(layer1_outputs(8493)) or (layer1_outputs(7939));
    layer2_outputs(3954) <= (layer1_outputs(6970)) and (layer1_outputs(8046));
    layer2_outputs(3955) <= layer1_outputs(7563);
    layer2_outputs(3956) <= not((layer1_outputs(7074)) and (layer1_outputs(10197)));
    layer2_outputs(3957) <= not(layer1_outputs(4681));
    layer2_outputs(3958) <= not((layer1_outputs(1527)) and (layer1_outputs(2252)));
    layer2_outputs(3959) <= (layer1_outputs(3364)) and not (layer1_outputs(5575));
    layer2_outputs(3960) <= not(layer1_outputs(5997));
    layer2_outputs(3961) <= (layer1_outputs(4006)) and not (layer1_outputs(8800));
    layer2_outputs(3962) <= layer1_outputs(2099);
    layer2_outputs(3963) <= not(layer1_outputs(9082)) or (layer1_outputs(3657));
    layer2_outputs(3964) <= (layer1_outputs(1499)) or (layer1_outputs(5204));
    layer2_outputs(3965) <= (layer1_outputs(1808)) and not (layer1_outputs(2252));
    layer2_outputs(3966) <= (layer1_outputs(7097)) or (layer1_outputs(8193));
    layer2_outputs(3967) <= (layer1_outputs(3147)) xor (layer1_outputs(1937));
    layer2_outputs(3968) <= layer1_outputs(3974);
    layer2_outputs(3969) <= not(layer1_outputs(644)) or (layer1_outputs(812));
    layer2_outputs(3970) <= not(layer1_outputs(4810)) or (layer1_outputs(7131));
    layer2_outputs(3971) <= (layer1_outputs(760)) and not (layer1_outputs(8709));
    layer2_outputs(3972) <= (layer1_outputs(8418)) and (layer1_outputs(7976));
    layer2_outputs(3973) <= not((layer1_outputs(5713)) xor (layer1_outputs(1723)));
    layer2_outputs(3974) <= not(layer1_outputs(251));
    layer2_outputs(3975) <= (layer1_outputs(6098)) and not (layer1_outputs(7695));
    layer2_outputs(3976) <= layer1_outputs(5698);
    layer2_outputs(3977) <= not((layer1_outputs(4811)) or (layer1_outputs(2032)));
    layer2_outputs(3978) <= not((layer1_outputs(2565)) and (layer1_outputs(893)));
    layer2_outputs(3979) <= (layer1_outputs(9081)) xor (layer1_outputs(8194));
    layer2_outputs(3980) <= (layer1_outputs(9233)) and not (layer1_outputs(6206));
    layer2_outputs(3981) <= not(layer1_outputs(9857)) or (layer1_outputs(8995));
    layer2_outputs(3982) <= layer1_outputs(527);
    layer2_outputs(3983) <= not((layer1_outputs(565)) or (layer1_outputs(67)));
    layer2_outputs(3984) <= not(layer1_outputs(5693)) or (layer1_outputs(3550));
    layer2_outputs(3985) <= not((layer1_outputs(1228)) or (layer1_outputs(5161)));
    layer2_outputs(3986) <= layer1_outputs(9341);
    layer2_outputs(3987) <= layer1_outputs(10016);
    layer2_outputs(3988) <= (layer1_outputs(9623)) and not (layer1_outputs(1830));
    layer2_outputs(3989) <= not(layer1_outputs(2667));
    layer2_outputs(3990) <= (layer1_outputs(10005)) xor (layer1_outputs(10059));
    layer2_outputs(3991) <= not((layer1_outputs(866)) or (layer1_outputs(3353)));
    layer2_outputs(3992) <= not((layer1_outputs(6381)) and (layer1_outputs(129)));
    layer2_outputs(3993) <= (layer1_outputs(7242)) and (layer1_outputs(1609));
    layer2_outputs(3994) <= '1';
    layer2_outputs(3995) <= not((layer1_outputs(2861)) xor (layer1_outputs(3582)));
    layer2_outputs(3996) <= layer1_outputs(4049);
    layer2_outputs(3997) <= layer1_outputs(2697);
    layer2_outputs(3998) <= not(layer1_outputs(5831)) or (layer1_outputs(3813));
    layer2_outputs(3999) <= layer1_outputs(1543);
    layer2_outputs(4000) <= not(layer1_outputs(4421));
    layer2_outputs(4001) <= not(layer1_outputs(13));
    layer2_outputs(4002) <= '1';
    layer2_outputs(4003) <= not(layer1_outputs(4197)) or (layer1_outputs(3763));
    layer2_outputs(4004) <= (layer1_outputs(7790)) and not (layer1_outputs(5682));
    layer2_outputs(4005) <= not(layer1_outputs(2900));
    layer2_outputs(4006) <= not(layer1_outputs(1060));
    layer2_outputs(4007) <= not(layer1_outputs(5185)) or (layer1_outputs(5057));
    layer2_outputs(4008) <= '0';
    layer2_outputs(4009) <= not(layer1_outputs(1805));
    layer2_outputs(4010) <= not(layer1_outputs(2460)) or (layer1_outputs(2455));
    layer2_outputs(4011) <= (layer1_outputs(9719)) and (layer1_outputs(9014));
    layer2_outputs(4012) <= layer1_outputs(5714);
    layer2_outputs(4013) <= not(layer1_outputs(1880));
    layer2_outputs(4014) <= not((layer1_outputs(3328)) and (layer1_outputs(1526)));
    layer2_outputs(4015) <= '1';
    layer2_outputs(4016) <= '0';
    layer2_outputs(4017) <= not((layer1_outputs(4652)) and (layer1_outputs(5249)));
    layer2_outputs(4018) <= layer1_outputs(9796);
    layer2_outputs(4019) <= not(layer1_outputs(6453));
    layer2_outputs(4020) <= not((layer1_outputs(6346)) or (layer1_outputs(7014)));
    layer2_outputs(4021) <= not(layer1_outputs(5474));
    layer2_outputs(4022) <= (layer1_outputs(1398)) and (layer1_outputs(2226));
    layer2_outputs(4023) <= (layer1_outputs(7903)) and not (layer1_outputs(5661));
    layer2_outputs(4024) <= not(layer1_outputs(6932));
    layer2_outputs(4025) <= not(layer1_outputs(2305)) or (layer1_outputs(8949));
    layer2_outputs(4026) <= not(layer1_outputs(3010)) or (layer1_outputs(4042));
    layer2_outputs(4027) <= layer1_outputs(8153);
    layer2_outputs(4028) <= (layer1_outputs(2084)) or (layer1_outputs(5999));
    layer2_outputs(4029) <= not(layer1_outputs(540));
    layer2_outputs(4030) <= not((layer1_outputs(4514)) and (layer1_outputs(9193)));
    layer2_outputs(4031) <= not((layer1_outputs(9627)) and (layer1_outputs(9575)));
    layer2_outputs(4032) <= not(layer1_outputs(6575)) or (layer1_outputs(7041));
    layer2_outputs(4033) <= '0';
    layer2_outputs(4034) <= layer1_outputs(361);
    layer2_outputs(4035) <= (layer1_outputs(9568)) and not (layer1_outputs(6975));
    layer2_outputs(4036) <= not((layer1_outputs(3790)) or (layer1_outputs(6840)));
    layer2_outputs(4037) <= (layer1_outputs(9325)) and not (layer1_outputs(8981));
    layer2_outputs(4038) <= not(layer1_outputs(4792));
    layer2_outputs(4039) <= not(layer1_outputs(6777));
    layer2_outputs(4040) <= layer1_outputs(1409);
    layer2_outputs(4041) <= not(layer1_outputs(6588));
    layer2_outputs(4042) <= (layer1_outputs(6457)) or (layer1_outputs(3061));
    layer2_outputs(4043) <= not(layer1_outputs(1826));
    layer2_outputs(4044) <= layer1_outputs(6333);
    layer2_outputs(4045) <= not(layer1_outputs(6700)) or (layer1_outputs(8608));
    layer2_outputs(4046) <= layer1_outputs(6191);
    layer2_outputs(4047) <= layer1_outputs(8561);
    layer2_outputs(4048) <= (layer1_outputs(8332)) and not (layer1_outputs(10056));
    layer2_outputs(4049) <= layer1_outputs(415);
    layer2_outputs(4050) <= not(layer1_outputs(9751)) or (layer1_outputs(2825));
    layer2_outputs(4051) <= (layer1_outputs(7956)) and not (layer1_outputs(6815));
    layer2_outputs(4052) <= not(layer1_outputs(3541));
    layer2_outputs(4053) <= (layer1_outputs(9796)) and (layer1_outputs(725));
    layer2_outputs(4054) <= not(layer1_outputs(9681));
    layer2_outputs(4055) <= not((layer1_outputs(2186)) or (layer1_outputs(3424)));
    layer2_outputs(4056) <= not(layer1_outputs(7474));
    layer2_outputs(4057) <= not(layer1_outputs(8817)) or (layer1_outputs(296));
    layer2_outputs(4058) <= not((layer1_outputs(2619)) or (layer1_outputs(6295)));
    layer2_outputs(4059) <= not(layer1_outputs(3198)) or (layer1_outputs(9866));
    layer2_outputs(4060) <= (layer1_outputs(1930)) and (layer1_outputs(1802));
    layer2_outputs(4061) <= not((layer1_outputs(4968)) and (layer1_outputs(1405)));
    layer2_outputs(4062) <= (layer1_outputs(2914)) or (layer1_outputs(10062));
    layer2_outputs(4063) <= (layer1_outputs(9140)) and not (layer1_outputs(5645));
    layer2_outputs(4064) <= layer1_outputs(7471);
    layer2_outputs(4065) <= layer1_outputs(7301);
    layer2_outputs(4066) <= not(layer1_outputs(10092)) or (layer1_outputs(7347));
    layer2_outputs(4067) <= not((layer1_outputs(982)) and (layer1_outputs(9450)));
    layer2_outputs(4068) <= not(layer1_outputs(8088));
    layer2_outputs(4069) <= not(layer1_outputs(7988));
    layer2_outputs(4070) <= not(layer1_outputs(884)) or (layer1_outputs(6972));
    layer2_outputs(4071) <= (layer1_outputs(315)) or (layer1_outputs(7029));
    layer2_outputs(4072) <= not((layer1_outputs(6065)) and (layer1_outputs(1002)));
    layer2_outputs(4073) <= not((layer1_outputs(245)) or (layer1_outputs(8162)));
    layer2_outputs(4074) <= (layer1_outputs(2548)) and not (layer1_outputs(5457));
    layer2_outputs(4075) <= not(layer1_outputs(5531)) or (layer1_outputs(8300));
    layer2_outputs(4076) <= layer1_outputs(6555);
    layer2_outputs(4077) <= not(layer1_outputs(3506));
    layer2_outputs(4078) <= not((layer1_outputs(9095)) xor (layer1_outputs(6047)));
    layer2_outputs(4079) <= layer1_outputs(1416);
    layer2_outputs(4080) <= not((layer1_outputs(8411)) xor (layer1_outputs(5018)));
    layer2_outputs(4081) <= not(layer1_outputs(5492)) or (layer1_outputs(9678));
    layer2_outputs(4082) <= not(layer1_outputs(5180));
    layer2_outputs(4083) <= layer1_outputs(7525);
    layer2_outputs(4084) <= not((layer1_outputs(2043)) xor (layer1_outputs(5128)));
    layer2_outputs(4085) <= not((layer1_outputs(9576)) and (layer1_outputs(2341)));
    layer2_outputs(4086) <= (layer1_outputs(4729)) and (layer1_outputs(7173));
    layer2_outputs(4087) <= not(layer1_outputs(808));
    layer2_outputs(4088) <= not((layer1_outputs(4840)) or (layer1_outputs(4903)));
    layer2_outputs(4089) <= '1';
    layer2_outputs(4090) <= layer1_outputs(557);
    layer2_outputs(4091) <= not(layer1_outputs(8284));
    layer2_outputs(4092) <= not(layer1_outputs(8557));
    layer2_outputs(4093) <= '1';
    layer2_outputs(4094) <= not(layer1_outputs(4272));
    layer2_outputs(4095) <= not((layer1_outputs(2872)) xor (layer1_outputs(6278)));
    layer2_outputs(4096) <= not(layer1_outputs(1675)) or (layer1_outputs(6694));
    layer2_outputs(4097) <= not(layer1_outputs(3386)) or (layer1_outputs(9664));
    layer2_outputs(4098) <= not((layer1_outputs(8612)) xor (layer1_outputs(2569)));
    layer2_outputs(4099) <= layer1_outputs(3893);
    layer2_outputs(4100) <= not((layer1_outputs(958)) and (layer1_outputs(6927)));
    layer2_outputs(4101) <= (layer1_outputs(7706)) xor (layer1_outputs(4960));
    layer2_outputs(4102) <= '0';
    layer2_outputs(4103) <= not((layer1_outputs(10037)) and (layer1_outputs(7110)));
    layer2_outputs(4104) <= layer1_outputs(8930);
    layer2_outputs(4105) <= (layer1_outputs(5833)) and (layer1_outputs(3394));
    layer2_outputs(4106) <= (layer1_outputs(1031)) and (layer1_outputs(5908));
    layer2_outputs(4107) <= (layer1_outputs(8740)) and not (layer1_outputs(1542));
    layer2_outputs(4108) <= not(layer1_outputs(8689)) or (layer1_outputs(8372));
    layer2_outputs(4109) <= (layer1_outputs(4969)) or (layer1_outputs(2436));
    layer2_outputs(4110) <= (layer1_outputs(809)) and (layer1_outputs(298));
    layer2_outputs(4111) <= layer1_outputs(5885);
    layer2_outputs(4112) <= (layer1_outputs(4337)) and not (layer1_outputs(2647));
    layer2_outputs(4113) <= (layer1_outputs(3852)) and not (layer1_outputs(983));
    layer2_outputs(4114) <= not((layer1_outputs(846)) or (layer1_outputs(3906)));
    layer2_outputs(4115) <= not(layer1_outputs(8834)) or (layer1_outputs(4439));
    layer2_outputs(4116) <= not((layer1_outputs(2232)) or (layer1_outputs(6871)));
    layer2_outputs(4117) <= layer1_outputs(870);
    layer2_outputs(4118) <= not((layer1_outputs(3756)) and (layer1_outputs(10107)));
    layer2_outputs(4119) <= (layer1_outputs(1934)) xor (layer1_outputs(2136));
    layer2_outputs(4120) <= (layer1_outputs(6527)) and not (layer1_outputs(410));
    layer2_outputs(4121) <= not((layer1_outputs(995)) or (layer1_outputs(1820)));
    layer2_outputs(4122) <= not(layer1_outputs(5318)) or (layer1_outputs(475));
    layer2_outputs(4123) <= not(layer1_outputs(3676));
    layer2_outputs(4124) <= layer1_outputs(3866);
    layer2_outputs(4125) <= (layer1_outputs(4007)) xor (layer1_outputs(1699));
    layer2_outputs(4126) <= layer1_outputs(7064);
    layer2_outputs(4127) <= (layer1_outputs(2505)) and (layer1_outputs(7745));
    layer2_outputs(4128) <= not(layer1_outputs(2428));
    layer2_outputs(4129) <= (layer1_outputs(6082)) and not (layer1_outputs(4243));
    layer2_outputs(4130) <= not(layer1_outputs(2450));
    layer2_outputs(4131) <= not(layer1_outputs(4717)) or (layer1_outputs(10089));
    layer2_outputs(4132) <= layer1_outputs(5523);
    layer2_outputs(4133) <= layer1_outputs(9555);
    layer2_outputs(4134) <= layer1_outputs(8191);
    layer2_outputs(4135) <= (layer1_outputs(1273)) and (layer1_outputs(2089));
    layer2_outputs(4136) <= not(layer1_outputs(8221));
    layer2_outputs(4137) <= '0';
    layer2_outputs(4138) <= layer1_outputs(7027);
    layer2_outputs(4139) <= not(layer1_outputs(2047));
    layer2_outputs(4140) <= layer1_outputs(6746);
    layer2_outputs(4141) <= not(layer1_outputs(8329)) or (layer1_outputs(1973));
    layer2_outputs(4142) <= not((layer1_outputs(9798)) xor (layer1_outputs(601)));
    layer2_outputs(4143) <= (layer1_outputs(1494)) and not (layer1_outputs(10078));
    layer2_outputs(4144) <= (layer1_outputs(7454)) xor (layer1_outputs(6854));
    layer2_outputs(4145) <= layer1_outputs(6363);
    layer2_outputs(4146) <= not(layer1_outputs(1906));
    layer2_outputs(4147) <= not((layer1_outputs(4342)) xor (layer1_outputs(6684)));
    layer2_outputs(4148) <= not((layer1_outputs(5392)) and (layer1_outputs(8576)));
    layer2_outputs(4149) <= '1';
    layer2_outputs(4150) <= (layer1_outputs(815)) and not (layer1_outputs(6338));
    layer2_outputs(4151) <= '0';
    layer2_outputs(4152) <= (layer1_outputs(5372)) and not (layer1_outputs(1293));
    layer2_outputs(4153) <= (layer1_outputs(6710)) xor (layer1_outputs(618));
    layer2_outputs(4154) <= '0';
    layer2_outputs(4155) <= (layer1_outputs(8124)) and not (layer1_outputs(1115));
    layer2_outputs(4156) <= not((layer1_outputs(7251)) and (layer1_outputs(5149)));
    layer2_outputs(4157) <= not(layer1_outputs(3153)) or (layer1_outputs(1072));
    layer2_outputs(4158) <= (layer1_outputs(1846)) and (layer1_outputs(9112));
    layer2_outputs(4159) <= layer1_outputs(508);
    layer2_outputs(4160) <= (layer1_outputs(227)) and not (layer1_outputs(3241));
    layer2_outputs(4161) <= layer1_outputs(7121);
    layer2_outputs(4162) <= (layer1_outputs(2947)) and (layer1_outputs(3225));
    layer2_outputs(4163) <= not((layer1_outputs(8426)) or (layer1_outputs(8739)));
    layer2_outputs(4164) <= not(layer1_outputs(6755));
    layer2_outputs(4165) <= layer1_outputs(3799);
    layer2_outputs(4166) <= layer1_outputs(7860);
    layer2_outputs(4167) <= layer1_outputs(990);
    layer2_outputs(4168) <= '0';
    layer2_outputs(4169) <= not((layer1_outputs(2306)) and (layer1_outputs(1169)));
    layer2_outputs(4170) <= not((layer1_outputs(8350)) or (layer1_outputs(9263)));
    layer2_outputs(4171) <= not((layer1_outputs(9846)) and (layer1_outputs(6448)));
    layer2_outputs(4172) <= (layer1_outputs(465)) xor (layer1_outputs(6821));
    layer2_outputs(4173) <= not(layer1_outputs(5088)) or (layer1_outputs(2623));
    layer2_outputs(4174) <= not((layer1_outputs(6042)) and (layer1_outputs(1167)));
    layer2_outputs(4175) <= layer1_outputs(2982);
    layer2_outputs(4176) <= layer1_outputs(3218);
    layer2_outputs(4177) <= not((layer1_outputs(9307)) xor (layer1_outputs(2235)));
    layer2_outputs(4178) <= (layer1_outputs(2141)) and not (layer1_outputs(8639));
    layer2_outputs(4179) <= not((layer1_outputs(9930)) xor (layer1_outputs(866)));
    layer2_outputs(4180) <= (layer1_outputs(6799)) and not (layer1_outputs(7823));
    layer2_outputs(4181) <= not((layer1_outputs(5592)) xor (layer1_outputs(6198)));
    layer2_outputs(4182) <= not((layer1_outputs(7487)) and (layer1_outputs(730)));
    layer2_outputs(4183) <= not(layer1_outputs(7124));
    layer2_outputs(4184) <= not(layer1_outputs(7695)) or (layer1_outputs(2807));
    layer2_outputs(4185) <= layer1_outputs(1046);
    layer2_outputs(4186) <= not(layer1_outputs(6880));
    layer2_outputs(4187) <= not(layer1_outputs(7901)) or (layer1_outputs(2079));
    layer2_outputs(4188) <= '0';
    layer2_outputs(4189) <= (layer1_outputs(6752)) and not (layer1_outputs(5425));
    layer2_outputs(4190) <= layer1_outputs(1591);
    layer2_outputs(4191) <= not(layer1_outputs(7022));
    layer2_outputs(4192) <= (layer1_outputs(9760)) and not (layer1_outputs(9145));
    layer2_outputs(4193) <= not(layer1_outputs(5231)) or (layer1_outputs(7363));
    layer2_outputs(4194) <= not((layer1_outputs(886)) and (layer1_outputs(8786)));
    layer2_outputs(4195) <= not(layer1_outputs(5641));
    layer2_outputs(4196) <= not(layer1_outputs(771)) or (layer1_outputs(9514));
    layer2_outputs(4197) <= (layer1_outputs(7629)) and (layer1_outputs(3478));
    layer2_outputs(4198) <= not(layer1_outputs(8919));
    layer2_outputs(4199) <= layer1_outputs(2534);
    layer2_outputs(4200) <= not(layer1_outputs(320));
    layer2_outputs(4201) <= not(layer1_outputs(1060));
    layer2_outputs(4202) <= not((layer1_outputs(1660)) xor (layer1_outputs(82)));
    layer2_outputs(4203) <= not(layer1_outputs(7672));
    layer2_outputs(4204) <= (layer1_outputs(8917)) and not (layer1_outputs(7729));
    layer2_outputs(4205) <= (layer1_outputs(3576)) and not (layer1_outputs(3162));
    layer2_outputs(4206) <= not((layer1_outputs(11)) xor (layer1_outputs(9914)));
    layer2_outputs(4207) <= not(layer1_outputs(4532));
    layer2_outputs(4208) <= layer1_outputs(5533);
    layer2_outputs(4209) <= not((layer1_outputs(3857)) xor (layer1_outputs(1248)));
    layer2_outputs(4210) <= not((layer1_outputs(1265)) or (layer1_outputs(4845)));
    layer2_outputs(4211) <= (layer1_outputs(9961)) and (layer1_outputs(1525));
    layer2_outputs(4212) <= not(layer1_outputs(8952));
    layer2_outputs(4213) <= not((layer1_outputs(4423)) xor (layer1_outputs(1727)));
    layer2_outputs(4214) <= '1';
    layer2_outputs(4215) <= not(layer1_outputs(8977));
    layer2_outputs(4216) <= not(layer1_outputs(3099)) or (layer1_outputs(5078));
    layer2_outputs(4217) <= not(layer1_outputs(1802));
    layer2_outputs(4218) <= not(layer1_outputs(3797));
    layer2_outputs(4219) <= not(layer1_outputs(1490)) or (layer1_outputs(3051));
    layer2_outputs(4220) <= not(layer1_outputs(5580));
    layer2_outputs(4221) <= layer1_outputs(3896);
    layer2_outputs(4222) <= not((layer1_outputs(6569)) and (layer1_outputs(8898)));
    layer2_outputs(4223) <= (layer1_outputs(3152)) or (layer1_outputs(9792));
    layer2_outputs(4224) <= (layer1_outputs(5941)) xor (layer1_outputs(6065));
    layer2_outputs(4225) <= layer1_outputs(4547);
    layer2_outputs(4226) <= not(layer1_outputs(3252));
    layer2_outputs(4227) <= not(layer1_outputs(988));
    layer2_outputs(4228) <= not(layer1_outputs(531)) or (layer1_outputs(9752));
    layer2_outputs(4229) <= layer1_outputs(2528);
    layer2_outputs(4230) <= not(layer1_outputs(3227));
    layer2_outputs(4231) <= (layer1_outputs(113)) and not (layer1_outputs(2487));
    layer2_outputs(4232) <= (layer1_outputs(3843)) xor (layer1_outputs(1425));
    layer2_outputs(4233) <= '1';
    layer2_outputs(4234) <= not(layer1_outputs(5669)) or (layer1_outputs(5146));
    layer2_outputs(4235) <= not(layer1_outputs(1609));
    layer2_outputs(4236) <= layer1_outputs(9286);
    layer2_outputs(4237) <= '0';
    layer2_outputs(4238) <= layer1_outputs(1814);
    layer2_outputs(4239) <= (layer1_outputs(2701)) and (layer1_outputs(1282));
    layer2_outputs(4240) <= layer1_outputs(5822);
    layer2_outputs(4241) <= not(layer1_outputs(1557));
    layer2_outputs(4242) <= not(layer1_outputs(4794)) or (layer1_outputs(6054));
    layer2_outputs(4243) <= not(layer1_outputs(4035));
    layer2_outputs(4244) <= (layer1_outputs(7121)) and (layer1_outputs(6465));
    layer2_outputs(4245) <= (layer1_outputs(6698)) and (layer1_outputs(7167));
    layer2_outputs(4246) <= not((layer1_outputs(6286)) xor (layer1_outputs(6577)));
    layer2_outputs(4247) <= '1';
    layer2_outputs(4248) <= '1';
    layer2_outputs(4249) <= (layer1_outputs(6286)) xor (layer1_outputs(4629));
    layer2_outputs(4250) <= not(layer1_outputs(2989));
    layer2_outputs(4251) <= (layer1_outputs(3986)) or (layer1_outputs(7019));
    layer2_outputs(4252) <= '0';
    layer2_outputs(4253) <= not(layer1_outputs(5241)) or (layer1_outputs(395));
    layer2_outputs(4254) <= (layer1_outputs(8533)) and not (layer1_outputs(5237));
    layer2_outputs(4255) <= not(layer1_outputs(7702));
    layer2_outputs(4256) <= not(layer1_outputs(4856));
    layer2_outputs(4257) <= not((layer1_outputs(3527)) and (layer1_outputs(6326)));
    layer2_outputs(4258) <= not(layer1_outputs(8928));
    layer2_outputs(4259) <= not(layer1_outputs(4560));
    layer2_outputs(4260) <= not(layer1_outputs(392)) or (layer1_outputs(10149));
    layer2_outputs(4261) <= layer1_outputs(3492);
    layer2_outputs(4262) <= '1';
    layer2_outputs(4263) <= not(layer1_outputs(2071));
    layer2_outputs(4264) <= not(layer1_outputs(3828));
    layer2_outputs(4265) <= '1';
    layer2_outputs(4266) <= layer1_outputs(8346);
    layer2_outputs(4267) <= (layer1_outputs(2171)) xor (layer1_outputs(6));
    layer2_outputs(4268) <= (layer1_outputs(8990)) xor (layer1_outputs(3807));
    layer2_outputs(4269) <= (layer1_outputs(5356)) and not (layer1_outputs(5415));
    layer2_outputs(4270) <= not(layer1_outputs(58)) or (layer1_outputs(3528));
    layer2_outputs(4271) <= not(layer1_outputs(1079));
    layer2_outputs(4272) <= layer1_outputs(9361);
    layer2_outputs(4273) <= not(layer1_outputs(8718)) or (layer1_outputs(5085));
    layer2_outputs(4274) <= layer1_outputs(4301);
    layer2_outputs(4275) <= not((layer1_outputs(3896)) or (layer1_outputs(2699)));
    layer2_outputs(4276) <= not(layer1_outputs(7371));
    layer2_outputs(4277) <= (layer1_outputs(4853)) and (layer1_outputs(8275));
    layer2_outputs(4278) <= (layer1_outputs(6490)) and not (layer1_outputs(2052));
    layer2_outputs(4279) <= layer1_outputs(4198);
    layer2_outputs(4280) <= not((layer1_outputs(8246)) or (layer1_outputs(2002)));
    layer2_outputs(4281) <= layer1_outputs(3243);
    layer2_outputs(4282) <= not(layer1_outputs(5299));
    layer2_outputs(4283) <= (layer1_outputs(4415)) and not (layer1_outputs(8091));
    layer2_outputs(4284) <= not(layer1_outputs(898)) or (layer1_outputs(9763));
    layer2_outputs(4285) <= (layer1_outputs(7280)) and not (layer1_outputs(9519));
    layer2_outputs(4286) <= not((layer1_outputs(581)) and (layer1_outputs(1964)));
    layer2_outputs(4287) <= (layer1_outputs(7496)) and (layer1_outputs(1736));
    layer2_outputs(4288) <= not(layer1_outputs(6541));
    layer2_outputs(4289) <= '1';
    layer2_outputs(4290) <= layer1_outputs(63);
    layer2_outputs(4291) <= layer1_outputs(5880);
    layer2_outputs(4292) <= not(layer1_outputs(8233));
    layer2_outputs(4293) <= (layer1_outputs(3109)) or (layer1_outputs(6577));
    layer2_outputs(4294) <= not(layer1_outputs(9680)) or (layer1_outputs(49));
    layer2_outputs(4295) <= '0';
    layer2_outputs(4296) <= (layer1_outputs(3237)) xor (layer1_outputs(2230));
    layer2_outputs(4297) <= not(layer1_outputs(8241));
    layer2_outputs(4298) <= layer1_outputs(4285);
    layer2_outputs(4299) <= (layer1_outputs(2452)) xor (layer1_outputs(9450));
    layer2_outputs(4300) <= not(layer1_outputs(3121));
    layer2_outputs(4301) <= not(layer1_outputs(1523));
    layer2_outputs(4302) <= not(layer1_outputs(697));
    layer2_outputs(4303) <= (layer1_outputs(10073)) and not (layer1_outputs(7670));
    layer2_outputs(4304) <= not(layer1_outputs(7622));
    layer2_outputs(4305) <= not(layer1_outputs(5676)) or (layer1_outputs(5156));
    layer2_outputs(4306) <= not((layer1_outputs(842)) and (layer1_outputs(8084)));
    layer2_outputs(4307) <= not(layer1_outputs(3633));
    layer2_outputs(4308) <= not(layer1_outputs(8355));
    layer2_outputs(4309) <= layer1_outputs(7705);
    layer2_outputs(4310) <= not(layer1_outputs(5293));
    layer2_outputs(4311) <= '1';
    layer2_outputs(4312) <= not(layer1_outputs(3582));
    layer2_outputs(4313) <= not(layer1_outputs(4716));
    layer2_outputs(4314) <= not(layer1_outputs(2606));
    layer2_outputs(4315) <= not((layer1_outputs(7927)) xor (layer1_outputs(9821)));
    layer2_outputs(4316) <= '0';
    layer2_outputs(4317) <= not(layer1_outputs(6696));
    layer2_outputs(4318) <= not(layer1_outputs(6405));
    layer2_outputs(4319) <= layer1_outputs(8311);
    layer2_outputs(4320) <= not((layer1_outputs(8082)) xor (layer1_outputs(5362)));
    layer2_outputs(4321) <= not((layer1_outputs(260)) and (layer1_outputs(2271)));
    layer2_outputs(4322) <= not(layer1_outputs(3194)) or (layer1_outputs(9296));
    layer2_outputs(4323) <= not(layer1_outputs(9615));
    layer2_outputs(4324) <= not(layer1_outputs(9044));
    layer2_outputs(4325) <= not(layer1_outputs(1230));
    layer2_outputs(4326) <= not(layer1_outputs(2431));
    layer2_outputs(4327) <= not(layer1_outputs(5875)) or (layer1_outputs(1605));
    layer2_outputs(4328) <= (layer1_outputs(4822)) and not (layer1_outputs(995));
    layer2_outputs(4329) <= layer1_outputs(4539);
    layer2_outputs(4330) <= (layer1_outputs(6881)) and not (layer1_outputs(9062));
    layer2_outputs(4331) <= layer1_outputs(6451);
    layer2_outputs(4332) <= (layer1_outputs(1365)) xor (layer1_outputs(5068));
    layer2_outputs(4333) <= layer1_outputs(261);
    layer2_outputs(4334) <= not((layer1_outputs(2587)) xor (layer1_outputs(1649)));
    layer2_outputs(4335) <= not(layer1_outputs(3278));
    layer2_outputs(4336) <= not((layer1_outputs(5832)) and (layer1_outputs(5601)));
    layer2_outputs(4337) <= layer1_outputs(1981);
    layer2_outputs(4338) <= layer1_outputs(2284);
    layer2_outputs(4339) <= layer1_outputs(9586);
    layer2_outputs(4340) <= not(layer1_outputs(6427));
    layer2_outputs(4341) <= (layer1_outputs(4324)) or (layer1_outputs(2968));
    layer2_outputs(4342) <= not(layer1_outputs(5394));
    layer2_outputs(4343) <= (layer1_outputs(6273)) and (layer1_outputs(7700));
    layer2_outputs(4344) <= layer1_outputs(5902);
    layer2_outputs(4345) <= (layer1_outputs(8137)) and not (layer1_outputs(9213));
    layer2_outputs(4346) <= not((layer1_outputs(3339)) and (layer1_outputs(6551)));
    layer2_outputs(4347) <= not(layer1_outputs(9535));
    layer2_outputs(4348) <= not(layer1_outputs(7554));
    layer2_outputs(4349) <= not((layer1_outputs(5199)) and (layer1_outputs(5555)));
    layer2_outputs(4350) <= not(layer1_outputs(7945)) or (layer1_outputs(4217));
    layer2_outputs(4351) <= layer1_outputs(9382);
    layer2_outputs(4352) <= not(layer1_outputs(7755));
    layer2_outputs(4353) <= not(layer1_outputs(3615)) or (layer1_outputs(459));
    layer2_outputs(4354) <= layer1_outputs(1463);
    layer2_outputs(4355) <= not(layer1_outputs(6175));
    layer2_outputs(4356) <= not(layer1_outputs(4500));
    layer2_outputs(4357) <= layer1_outputs(2320);
    layer2_outputs(4358) <= (layer1_outputs(7063)) and (layer1_outputs(5758));
    layer2_outputs(4359) <= layer1_outputs(5768);
    layer2_outputs(4360) <= not(layer1_outputs(1851));
    layer2_outputs(4361) <= not((layer1_outputs(7312)) and (layer1_outputs(4427)));
    layer2_outputs(4362) <= not(layer1_outputs(8940));
    layer2_outputs(4363) <= (layer1_outputs(3239)) and not (layer1_outputs(10116));
    layer2_outputs(4364) <= not((layer1_outputs(4079)) xor (layer1_outputs(1543)));
    layer2_outputs(4365) <= not((layer1_outputs(8152)) and (layer1_outputs(4837)));
    layer2_outputs(4366) <= not((layer1_outputs(4565)) or (layer1_outputs(9397)));
    layer2_outputs(4367) <= layer1_outputs(3698);
    layer2_outputs(4368) <= layer1_outputs(8336);
    layer2_outputs(4369) <= not((layer1_outputs(6643)) and (layer1_outputs(2366)));
    layer2_outputs(4370) <= not(layer1_outputs(1104));
    layer2_outputs(4371) <= (layer1_outputs(4242)) and not (layer1_outputs(2227));
    layer2_outputs(4372) <= (layer1_outputs(7709)) or (layer1_outputs(3343));
    layer2_outputs(4373) <= layer1_outputs(1032);
    layer2_outputs(4374) <= (layer1_outputs(6539)) or (layer1_outputs(1911));
    layer2_outputs(4375) <= layer1_outputs(8050);
    layer2_outputs(4376) <= not(layer1_outputs(5237));
    layer2_outputs(4377) <= not(layer1_outputs(3086));
    layer2_outputs(4378) <= not(layer1_outputs(4072));
    layer2_outputs(4379) <= not((layer1_outputs(750)) xor (layer1_outputs(309)));
    layer2_outputs(4380) <= layer1_outputs(2537);
    layer2_outputs(4381) <= not((layer1_outputs(5977)) or (layer1_outputs(7139)));
    layer2_outputs(4382) <= not(layer1_outputs(8537));
    layer2_outputs(4383) <= not(layer1_outputs(3894)) or (layer1_outputs(1271));
    layer2_outputs(4384) <= layer1_outputs(692);
    layer2_outputs(4385) <= layer1_outputs(7690);
    layer2_outputs(4386) <= not(layer1_outputs(7999));
    layer2_outputs(4387) <= layer1_outputs(8422);
    layer2_outputs(4388) <= (layer1_outputs(3373)) or (layer1_outputs(7083));
    layer2_outputs(4389) <= not(layer1_outputs(9483));
    layer2_outputs(4390) <= (layer1_outputs(7042)) and (layer1_outputs(2038));
    layer2_outputs(4391) <= not((layer1_outputs(8807)) or (layer1_outputs(3991)));
    layer2_outputs(4392) <= '1';
    layer2_outputs(4393) <= (layer1_outputs(9440)) or (layer1_outputs(4930));
    layer2_outputs(4394) <= not(layer1_outputs(852));
    layer2_outputs(4395) <= not(layer1_outputs(8650));
    layer2_outputs(4396) <= not(layer1_outputs(1548)) or (layer1_outputs(588));
    layer2_outputs(4397) <= layer1_outputs(4392);
    layer2_outputs(4398) <= layer1_outputs(8776);
    layer2_outputs(4399) <= (layer1_outputs(5774)) or (layer1_outputs(7136));
    layer2_outputs(4400) <= not(layer1_outputs(1421));
    layer2_outputs(4401) <= '0';
    layer2_outputs(4402) <= not(layer1_outputs(9937)) or (layer1_outputs(8506));
    layer2_outputs(4403) <= not(layer1_outputs(1734)) or (layer1_outputs(8291));
    layer2_outputs(4404) <= (layer1_outputs(5913)) xor (layer1_outputs(7844));
    layer2_outputs(4405) <= not(layer1_outputs(9814)) or (layer1_outputs(5344));
    layer2_outputs(4406) <= (layer1_outputs(7871)) and not (layer1_outputs(360));
    layer2_outputs(4407) <= not(layer1_outputs(6668));
    layer2_outputs(4408) <= layer1_outputs(5416);
    layer2_outputs(4409) <= not(layer1_outputs(4920)) or (layer1_outputs(8682));
    layer2_outputs(4410) <= not((layer1_outputs(4329)) and (layer1_outputs(78)));
    layer2_outputs(4411) <= not((layer1_outputs(195)) or (layer1_outputs(5328)));
    layer2_outputs(4412) <= '1';
    layer2_outputs(4413) <= not((layer1_outputs(8795)) xor (layer1_outputs(1428)));
    layer2_outputs(4414) <= layer1_outputs(6853);
    layer2_outputs(4415) <= (layer1_outputs(118)) or (layer1_outputs(1638));
    layer2_outputs(4416) <= (layer1_outputs(5784)) and not (layer1_outputs(8459));
    layer2_outputs(4417) <= (layer1_outputs(4986)) and (layer1_outputs(4287));
    layer2_outputs(4418) <= layer1_outputs(5686);
    layer2_outputs(4419) <= layer1_outputs(3291);
    layer2_outputs(4420) <= '1';
    layer2_outputs(4421) <= (layer1_outputs(525)) and not (layer1_outputs(4230));
    layer2_outputs(4422) <= (layer1_outputs(6624)) and not (layer1_outputs(3241));
    layer2_outputs(4423) <= (layer1_outputs(4780)) and (layer1_outputs(9129));
    layer2_outputs(4424) <= layer1_outputs(9518);
    layer2_outputs(4425) <= (layer1_outputs(5971)) or (layer1_outputs(4630));
    layer2_outputs(4426) <= (layer1_outputs(4394)) or (layer1_outputs(7455));
    layer2_outputs(4427) <= (layer1_outputs(2050)) and (layer1_outputs(8573));
    layer2_outputs(4428) <= (layer1_outputs(3559)) xor (layer1_outputs(766));
    layer2_outputs(4429) <= not(layer1_outputs(7435));
    layer2_outputs(4430) <= '1';
    layer2_outputs(4431) <= (layer1_outputs(2776)) and not (layer1_outputs(3259));
    layer2_outputs(4432) <= (layer1_outputs(5725)) or (layer1_outputs(7893));
    layer2_outputs(4433) <= not(layer1_outputs(5395));
    layer2_outputs(4434) <= (layer1_outputs(6196)) and (layer1_outputs(1896));
    layer2_outputs(4435) <= (layer1_outputs(984)) and not (layer1_outputs(17));
    layer2_outputs(4436) <= not(layer1_outputs(130));
    layer2_outputs(4437) <= (layer1_outputs(2308)) or (layer1_outputs(2491));
    layer2_outputs(4438) <= (layer1_outputs(3101)) and not (layer1_outputs(602));
    layer2_outputs(4439) <= not(layer1_outputs(4634)) or (layer1_outputs(156));
    layer2_outputs(4440) <= not((layer1_outputs(2602)) and (layer1_outputs(2806)));
    layer2_outputs(4441) <= (layer1_outputs(1972)) xor (layer1_outputs(9473));
    layer2_outputs(4442) <= (layer1_outputs(8810)) and not (layer1_outputs(7832));
    layer2_outputs(4443) <= layer1_outputs(5460);
    layer2_outputs(4444) <= layer1_outputs(1945);
    layer2_outputs(4445) <= layer1_outputs(5972);
    layer2_outputs(4446) <= layer1_outputs(6998);
    layer2_outputs(4447) <= (layer1_outputs(5661)) or (layer1_outputs(7907));
    layer2_outputs(4448) <= layer1_outputs(3033);
    layer2_outputs(4449) <= not((layer1_outputs(6609)) and (layer1_outputs(9065)));
    layer2_outputs(4450) <= (layer1_outputs(10122)) or (layer1_outputs(9033));
    layer2_outputs(4451) <= (layer1_outputs(8951)) and not (layer1_outputs(10134));
    layer2_outputs(4452) <= not((layer1_outputs(4846)) or (layer1_outputs(4253)));
    layer2_outputs(4453) <= not(layer1_outputs(4871)) or (layer1_outputs(7813));
    layer2_outputs(4454) <= not((layer1_outputs(8553)) or (layer1_outputs(4797)));
    layer2_outputs(4455) <= (layer1_outputs(9988)) and (layer1_outputs(6045));
    layer2_outputs(4456) <= layer1_outputs(224);
    layer2_outputs(4457) <= not((layer1_outputs(2198)) and (layer1_outputs(5663)));
    layer2_outputs(4458) <= not(layer1_outputs(306)) or (layer1_outputs(5045));
    layer2_outputs(4459) <= not(layer1_outputs(6901)) or (layer1_outputs(6058));
    layer2_outputs(4460) <= (layer1_outputs(8484)) xor (layer1_outputs(8884));
    layer2_outputs(4461) <= '0';
    layer2_outputs(4462) <= not(layer1_outputs(1804));
    layer2_outputs(4463) <= (layer1_outputs(1765)) and not (layer1_outputs(9246));
    layer2_outputs(4464) <= not(layer1_outputs(7831)) or (layer1_outputs(8033));
    layer2_outputs(4465) <= (layer1_outputs(2530)) xor (layer1_outputs(6335));
    layer2_outputs(4466) <= (layer1_outputs(56)) xor (layer1_outputs(2746));
    layer2_outputs(4467) <= (layer1_outputs(557)) and not (layer1_outputs(6167));
    layer2_outputs(4468) <= not((layer1_outputs(5241)) xor (layer1_outputs(1594)));
    layer2_outputs(4469) <= (layer1_outputs(9528)) xor (layer1_outputs(4856));
    layer2_outputs(4470) <= (layer1_outputs(7608)) or (layer1_outputs(122));
    layer2_outputs(4471) <= layer1_outputs(1991);
    layer2_outputs(4472) <= (layer1_outputs(7305)) and not (layer1_outputs(1165));
    layer2_outputs(4473) <= (layer1_outputs(2265)) or (layer1_outputs(8270));
    layer2_outputs(4474) <= layer1_outputs(2706);
    layer2_outputs(4475) <= not(layer1_outputs(7172));
    layer2_outputs(4476) <= not(layer1_outputs(7451)) or (layer1_outputs(1911));
    layer2_outputs(4477) <= (layer1_outputs(9690)) and not (layer1_outputs(839));
    layer2_outputs(4478) <= not(layer1_outputs(9242));
    layer2_outputs(4479) <= not(layer1_outputs(8104)) or (layer1_outputs(8716));
    layer2_outputs(4480) <= not(layer1_outputs(7802)) or (layer1_outputs(4170));
    layer2_outputs(4481) <= not((layer1_outputs(3918)) or (layer1_outputs(6782)));
    layer2_outputs(4482) <= '0';
    layer2_outputs(4483) <= not((layer1_outputs(7687)) or (layer1_outputs(507)));
    layer2_outputs(4484) <= not(layer1_outputs(45)) or (layer1_outputs(7353));
    layer2_outputs(4485) <= not(layer1_outputs(3285));
    layer2_outputs(4486) <= not(layer1_outputs(6293)) or (layer1_outputs(5348));
    layer2_outputs(4487) <= not((layer1_outputs(9175)) and (layer1_outputs(1701)));
    layer2_outputs(4488) <= layer1_outputs(223);
    layer2_outputs(4489) <= '0';
    layer2_outputs(4490) <= (layer1_outputs(2703)) and not (layer1_outputs(5878));
    layer2_outputs(4491) <= (layer1_outputs(8953)) and (layer1_outputs(3410));
    layer2_outputs(4492) <= not((layer1_outputs(91)) or (layer1_outputs(800)));
    layer2_outputs(4493) <= not(layer1_outputs(439));
    layer2_outputs(4494) <= layer1_outputs(9953);
    layer2_outputs(4495) <= (layer1_outputs(663)) xor (layer1_outputs(8231));
    layer2_outputs(4496) <= (layer1_outputs(7836)) or (layer1_outputs(9556));
    layer2_outputs(4497) <= not(layer1_outputs(2682));
    layer2_outputs(4498) <= layer1_outputs(6106);
    layer2_outputs(4499) <= not(layer1_outputs(4090));
    layer2_outputs(4500) <= not(layer1_outputs(6632)) or (layer1_outputs(9087));
    layer2_outputs(4501) <= not(layer1_outputs(8396)) or (layer1_outputs(3834));
    layer2_outputs(4502) <= not(layer1_outputs(3258));
    layer2_outputs(4503) <= not(layer1_outputs(9357));
    layer2_outputs(4504) <= layer1_outputs(1794);
    layer2_outputs(4505) <= layer1_outputs(9781);
    layer2_outputs(4506) <= (layer1_outputs(207)) or (layer1_outputs(5433));
    layer2_outputs(4507) <= (layer1_outputs(9948)) xor (layer1_outputs(1113));
    layer2_outputs(4508) <= not(layer1_outputs(18));
    layer2_outputs(4509) <= not(layer1_outputs(3996));
    layer2_outputs(4510) <= not(layer1_outputs(5247));
    layer2_outputs(4511) <= not((layer1_outputs(1512)) xor (layer1_outputs(4476)));
    layer2_outputs(4512) <= not(layer1_outputs(5104));
    layer2_outputs(4513) <= not(layer1_outputs(5472)) or (layer1_outputs(220));
    layer2_outputs(4514) <= not(layer1_outputs(2832));
    layer2_outputs(4515) <= not(layer1_outputs(669)) or (layer1_outputs(1479));
    layer2_outputs(4516) <= not(layer1_outputs(3020)) or (layer1_outputs(3119));
    layer2_outputs(4517) <= not(layer1_outputs(1293));
    layer2_outputs(4518) <= (layer1_outputs(5255)) or (layer1_outputs(7933));
    layer2_outputs(4519) <= not((layer1_outputs(451)) and (layer1_outputs(9627)));
    layer2_outputs(4520) <= not(layer1_outputs(453));
    layer2_outputs(4521) <= not(layer1_outputs(9697));
    layer2_outputs(4522) <= not(layer1_outputs(548));
    layer2_outputs(4523) <= '1';
    layer2_outputs(4524) <= not(layer1_outputs(2461));
    layer2_outputs(4525) <= not((layer1_outputs(9920)) or (layer1_outputs(8386)));
    layer2_outputs(4526) <= (layer1_outputs(8403)) and not (layer1_outputs(6974));
    layer2_outputs(4527) <= (layer1_outputs(670)) and not (layer1_outputs(5228));
    layer2_outputs(4528) <= (layer1_outputs(8969)) or (layer1_outputs(1626));
    layer2_outputs(4529) <= (layer1_outputs(7417)) and not (layer1_outputs(7306));
    layer2_outputs(4530) <= '1';
    layer2_outputs(4531) <= not(layer1_outputs(8428));
    layer2_outputs(4532) <= (layer1_outputs(10028)) and not (layer1_outputs(4274));
    layer2_outputs(4533) <= (layer1_outputs(9876)) and not (layer1_outputs(9675));
    layer2_outputs(4534) <= (layer1_outputs(8968)) xor (layer1_outputs(6876));
    layer2_outputs(4535) <= layer1_outputs(2082);
    layer2_outputs(4536) <= '1';
    layer2_outputs(4537) <= (layer1_outputs(4024)) and not (layer1_outputs(2670));
    layer2_outputs(4538) <= layer1_outputs(3169);
    layer2_outputs(4539) <= (layer1_outputs(6458)) and not (layer1_outputs(8698));
    layer2_outputs(4540) <= (layer1_outputs(3159)) or (layer1_outputs(2693));
    layer2_outputs(4541) <= layer1_outputs(7340);
    layer2_outputs(4542) <= layer1_outputs(9925);
    layer2_outputs(4543) <= not(layer1_outputs(5190)) or (layer1_outputs(4173));
    layer2_outputs(4544) <= '0';
    layer2_outputs(4545) <= layer1_outputs(9231);
    layer2_outputs(4546) <= not((layer1_outputs(2907)) or (layer1_outputs(438)));
    layer2_outputs(4547) <= not((layer1_outputs(8598)) xor (layer1_outputs(1533)));
    layer2_outputs(4548) <= '0';
    layer2_outputs(4549) <= '1';
    layer2_outputs(4550) <= layer1_outputs(3623);
    layer2_outputs(4551) <= not(layer1_outputs(9478));
    layer2_outputs(4552) <= not((layer1_outputs(4836)) or (layer1_outputs(7457)));
    layer2_outputs(4553) <= layer1_outputs(549);
    layer2_outputs(4554) <= not((layer1_outputs(1350)) or (layer1_outputs(631)));
    layer2_outputs(4555) <= '0';
    layer2_outputs(4556) <= '1';
    layer2_outputs(4557) <= layer1_outputs(7057);
    layer2_outputs(4558) <= not((layer1_outputs(3117)) or (layer1_outputs(4171)));
    layer2_outputs(4559) <= (layer1_outputs(1128)) and (layer1_outputs(3568));
    layer2_outputs(4560) <= not(layer1_outputs(7268)) or (layer1_outputs(7039));
    layer2_outputs(4561) <= not(layer1_outputs(5244));
    layer2_outputs(4562) <= layer1_outputs(1369);
    layer2_outputs(4563) <= not(layer1_outputs(3436)) or (layer1_outputs(6514));
    layer2_outputs(4564) <= layer1_outputs(158);
    layer2_outputs(4565) <= layer1_outputs(4244);
    layer2_outputs(4566) <= layer1_outputs(4792);
    layer2_outputs(4567) <= (layer1_outputs(2152)) and not (layer1_outputs(3081));
    layer2_outputs(4568) <= not((layer1_outputs(2028)) or (layer1_outputs(993)));
    layer2_outputs(4569) <= not(layer1_outputs(2023));
    layer2_outputs(4570) <= layer1_outputs(5366);
    layer2_outputs(4571) <= (layer1_outputs(7391)) and not (layer1_outputs(4579));
    layer2_outputs(4572) <= not(layer1_outputs(8487));
    layer2_outputs(4573) <= layer1_outputs(3512);
    layer2_outputs(4574) <= not(layer1_outputs(8824)) or (layer1_outputs(3823));
    layer2_outputs(4575) <= '1';
    layer2_outputs(4576) <= (layer1_outputs(8634)) or (layer1_outputs(9569));
    layer2_outputs(4577) <= (layer1_outputs(2248)) and not (layer1_outputs(5017));
    layer2_outputs(4578) <= '0';
    layer2_outputs(4579) <= layer1_outputs(3583);
    layer2_outputs(4580) <= not(layer1_outputs(9162)) or (layer1_outputs(2733));
    layer2_outputs(4581) <= not(layer1_outputs(3645)) or (layer1_outputs(9676));
    layer2_outputs(4582) <= layer1_outputs(9842);
    layer2_outputs(4583) <= not(layer1_outputs(1303));
    layer2_outputs(4584) <= not(layer1_outputs(10224));
    layer2_outputs(4585) <= (layer1_outputs(4854)) and not (layer1_outputs(8901));
    layer2_outputs(4586) <= (layer1_outputs(8313)) and not (layer1_outputs(8761));
    layer2_outputs(4587) <= (layer1_outputs(7133)) and (layer1_outputs(6236));
    layer2_outputs(4588) <= not(layer1_outputs(2049));
    layer2_outputs(4589) <= not(layer1_outputs(8779));
    layer2_outputs(4590) <= '1';
    layer2_outputs(4591) <= not((layer1_outputs(6057)) and (layer1_outputs(1746)));
    layer2_outputs(4592) <= layer1_outputs(4441);
    layer2_outputs(4593) <= not((layer1_outputs(4069)) or (layer1_outputs(7179)));
    layer2_outputs(4594) <= not((layer1_outputs(9431)) xor (layer1_outputs(7814)));
    layer2_outputs(4595) <= not(layer1_outputs(9543));
    layer2_outputs(4596) <= not(layer1_outputs(2149));
    layer2_outputs(4597) <= not(layer1_outputs(2234));
    layer2_outputs(4598) <= layer1_outputs(6352);
    layer2_outputs(4599) <= not(layer1_outputs(6429)) or (layer1_outputs(5974));
    layer2_outputs(4600) <= not((layer1_outputs(3548)) or (layer1_outputs(738)));
    layer2_outputs(4601) <= (layer1_outputs(5278)) and not (layer1_outputs(2258));
    layer2_outputs(4602) <= (layer1_outputs(3414)) or (layer1_outputs(1892));
    layer2_outputs(4603) <= (layer1_outputs(9762)) xor (layer1_outputs(5508));
    layer2_outputs(4604) <= not((layer1_outputs(8991)) or (layer1_outputs(8858)));
    layer2_outputs(4605) <= layer1_outputs(4895);
    layer2_outputs(4606) <= (layer1_outputs(6898)) and (layer1_outputs(9311));
    layer2_outputs(4607) <= layer1_outputs(4637);
    layer2_outputs(4608) <= (layer1_outputs(6554)) xor (layer1_outputs(3877));
    layer2_outputs(4609) <= (layer1_outputs(4270)) and not (layer1_outputs(7409));
    layer2_outputs(4610) <= not(layer1_outputs(5939));
    layer2_outputs(4611) <= (layer1_outputs(5187)) and not (layer1_outputs(4380));
    layer2_outputs(4612) <= (layer1_outputs(9392)) and not (layer1_outputs(5176));
    layer2_outputs(4613) <= '1';
    layer2_outputs(4614) <= '0';
    layer2_outputs(4615) <= not(layer1_outputs(533));
    layer2_outputs(4616) <= not(layer1_outputs(2731));
    layer2_outputs(4617) <= not(layer1_outputs(7639));
    layer2_outputs(4618) <= not(layer1_outputs(9271));
    layer2_outputs(4619) <= not(layer1_outputs(7463));
    layer2_outputs(4620) <= not((layer1_outputs(9544)) or (layer1_outputs(7270)));
    layer2_outputs(4621) <= not(layer1_outputs(4388)) or (layer1_outputs(558));
    layer2_outputs(4622) <= not((layer1_outputs(8681)) xor (layer1_outputs(4055)));
    layer2_outputs(4623) <= not(layer1_outputs(3391)) or (layer1_outputs(5803));
    layer2_outputs(4624) <= not((layer1_outputs(2254)) and (layer1_outputs(7561)));
    layer2_outputs(4625) <= layer1_outputs(827);
    layer2_outputs(4626) <= not((layer1_outputs(6313)) and (layer1_outputs(2948)));
    layer2_outputs(4627) <= layer1_outputs(8927);
    layer2_outputs(4628) <= not(layer1_outputs(8900)) or (layer1_outputs(8877));
    layer2_outputs(4629) <= (layer1_outputs(4247)) xor (layer1_outputs(1816));
    layer2_outputs(4630) <= (layer1_outputs(377)) xor (layer1_outputs(8512));
    layer2_outputs(4631) <= not((layer1_outputs(8557)) xor (layer1_outputs(6508)));
    layer2_outputs(4632) <= not(layer1_outputs(5199));
    layer2_outputs(4633) <= (layer1_outputs(1504)) xor (layer1_outputs(6545));
    layer2_outputs(4634) <= layer1_outputs(368);
    layer2_outputs(4635) <= not(layer1_outputs(8052)) or (layer1_outputs(6406));
    layer2_outputs(4636) <= not((layer1_outputs(2859)) or (layer1_outputs(5731)));
    layer2_outputs(4637) <= layer1_outputs(9508);
    layer2_outputs(4638) <= not(layer1_outputs(4429));
    layer2_outputs(4639) <= not(layer1_outputs(3438));
    layer2_outputs(4640) <= layer1_outputs(8);
    layer2_outputs(4641) <= (layer1_outputs(7026)) and not (layer1_outputs(5322));
    layer2_outputs(4642) <= layer1_outputs(8960);
    layer2_outputs(4643) <= not(layer1_outputs(9261));
    layer2_outputs(4644) <= not(layer1_outputs(285));
    layer2_outputs(4645) <= (layer1_outputs(6382)) or (layer1_outputs(1270));
    layer2_outputs(4646) <= layer1_outputs(6274);
    layer2_outputs(4647) <= layer1_outputs(317);
    layer2_outputs(4648) <= (layer1_outputs(9997)) and not (layer1_outputs(2098));
    layer2_outputs(4649) <= not(layer1_outputs(4761)) or (layer1_outputs(4935));
    layer2_outputs(4650) <= not(layer1_outputs(4878)) or (layer1_outputs(3286));
    layer2_outputs(4651) <= '1';
    layer2_outputs(4652) <= layer1_outputs(2086);
    layer2_outputs(4653) <= not(layer1_outputs(2943));
    layer2_outputs(4654) <= layer1_outputs(9114);
    layer2_outputs(4655) <= not(layer1_outputs(48));
    layer2_outputs(4656) <= layer1_outputs(9078);
    layer2_outputs(4657) <= (layer1_outputs(8316)) and not (layer1_outputs(3133));
    layer2_outputs(4658) <= layer1_outputs(3786);
    layer2_outputs(4659) <= (layer1_outputs(5133)) or (layer1_outputs(4467));
    layer2_outputs(4660) <= (layer1_outputs(3944)) and not (layer1_outputs(6193));
    layer2_outputs(4661) <= not((layer1_outputs(7863)) and (layer1_outputs(9054)));
    layer2_outputs(4662) <= (layer1_outputs(7060)) and not (layer1_outputs(7313));
    layer2_outputs(4663) <= not((layer1_outputs(2138)) and (layer1_outputs(8243)));
    layer2_outputs(4664) <= layer1_outputs(2846);
    layer2_outputs(4665) <= (layer1_outputs(6323)) and (layer1_outputs(4003));
    layer2_outputs(4666) <= not((layer1_outputs(2007)) and (layer1_outputs(5754)));
    layer2_outputs(4667) <= not(layer1_outputs(8200));
    layer2_outputs(4668) <= '1';
    layer2_outputs(4669) <= not((layer1_outputs(1413)) or (layer1_outputs(7263)));
    layer2_outputs(4670) <= (layer1_outputs(3677)) and (layer1_outputs(6213));
    layer2_outputs(4671) <= not((layer1_outputs(6797)) or (layer1_outputs(2747)));
    layer2_outputs(4672) <= (layer1_outputs(9899)) xor (layer1_outputs(1537));
    layer2_outputs(4673) <= not(layer1_outputs(9533));
    layer2_outputs(4674) <= not((layer1_outputs(5596)) or (layer1_outputs(1725)));
    layer2_outputs(4675) <= layer1_outputs(751);
    layer2_outputs(4676) <= not(layer1_outputs(5461));
    layer2_outputs(4677) <= (layer1_outputs(6704)) or (layer1_outputs(1227));
    layer2_outputs(4678) <= not((layer1_outputs(4126)) or (layer1_outputs(617)));
    layer2_outputs(4679) <= layer1_outputs(1287);
    layer2_outputs(4680) <= '1';
    layer2_outputs(4681) <= layer1_outputs(8889);
    layer2_outputs(4682) <= (layer1_outputs(5082)) and (layer1_outputs(7329));
    layer2_outputs(4683) <= (layer1_outputs(7195)) or (layer1_outputs(8714));
    layer2_outputs(4684) <= not(layer1_outputs(2572));
    layer2_outputs(4685) <= '1';
    layer2_outputs(4686) <= (layer1_outputs(8130)) and (layer1_outputs(6672));
    layer2_outputs(4687) <= not(layer1_outputs(654)) or (layer1_outputs(2888));
    layer2_outputs(4688) <= not(layer1_outputs(1337));
    layer2_outputs(4689) <= not(layer1_outputs(2946));
    layer2_outputs(4690) <= not((layer1_outputs(1716)) and (layer1_outputs(9221)));
    layer2_outputs(4691) <= (layer1_outputs(8635)) and not (layer1_outputs(7845));
    layer2_outputs(4692) <= (layer1_outputs(484)) and not (layer1_outputs(1234));
    layer2_outputs(4693) <= not((layer1_outputs(6149)) and (layer1_outputs(9284)));
    layer2_outputs(4694) <= not(layer1_outputs(6371)) or (layer1_outputs(9739));
    layer2_outputs(4695) <= layer1_outputs(7975);
    layer2_outputs(4696) <= layer1_outputs(1179);
    layer2_outputs(4697) <= not((layer1_outputs(1291)) and (layer1_outputs(8643)));
    layer2_outputs(4698) <= not(layer1_outputs(4147));
    layer2_outputs(4699) <= not(layer1_outputs(2486)) or (layer1_outputs(4704));
    layer2_outputs(4700) <= (layer1_outputs(2856)) and not (layer1_outputs(5271));
    layer2_outputs(4701) <= layer1_outputs(7085);
    layer2_outputs(4702) <= layer1_outputs(2142);
    layer2_outputs(4703) <= not((layer1_outputs(1180)) and (layer1_outputs(3977)));
    layer2_outputs(4704) <= (layer1_outputs(6347)) xor (layer1_outputs(5446));
    layer2_outputs(4705) <= (layer1_outputs(2698)) and not (layer1_outputs(3199));
    layer2_outputs(4706) <= layer1_outputs(3778);
    layer2_outputs(4707) <= not(layer1_outputs(5787));
    layer2_outputs(4708) <= layer1_outputs(3287);
    layer2_outputs(4709) <= layer1_outputs(7459);
    layer2_outputs(4710) <= not((layer1_outputs(1082)) xor (layer1_outputs(2099)));
    layer2_outputs(4711) <= layer1_outputs(2288);
    layer2_outputs(4712) <= '0';
    layer2_outputs(4713) <= not(layer1_outputs(3307));
    layer2_outputs(4714) <= (layer1_outputs(8517)) or (layer1_outputs(3285));
    layer2_outputs(4715) <= (layer1_outputs(8664)) and not (layer1_outputs(9826));
    layer2_outputs(4716) <= '1';
    layer2_outputs(4717) <= not(layer1_outputs(4192));
    layer2_outputs(4718) <= '1';
    layer2_outputs(4719) <= '1';
    layer2_outputs(4720) <= (layer1_outputs(6405)) and (layer1_outputs(4820));
    layer2_outputs(4721) <= (layer1_outputs(3217)) and not (layer1_outputs(4727));
    layer2_outputs(4722) <= not((layer1_outputs(4543)) or (layer1_outputs(3408)));
    layer2_outputs(4723) <= layer1_outputs(7874);
    layer2_outputs(4724) <= not(layer1_outputs(5626));
    layer2_outputs(4725) <= not(layer1_outputs(7885));
    layer2_outputs(4726) <= not((layer1_outputs(7903)) and (layer1_outputs(10001)));
    layer2_outputs(4727) <= (layer1_outputs(4385)) and not (layer1_outputs(9824));
    layer2_outputs(4728) <= not(layer1_outputs(1298)) or (layer1_outputs(8205));
    layer2_outputs(4729) <= not(layer1_outputs(3994));
    layer2_outputs(4730) <= (layer1_outputs(3844)) and not (layer1_outputs(7922));
    layer2_outputs(4731) <= not(layer1_outputs(1119));
    layer2_outputs(4732) <= layer1_outputs(7036);
    layer2_outputs(4733) <= not(layer1_outputs(7307));
    layer2_outputs(4734) <= not(layer1_outputs(1329));
    layer2_outputs(4735) <= (layer1_outputs(3843)) and (layer1_outputs(293));
    layer2_outputs(4736) <= (layer1_outputs(6648)) or (layer1_outputs(9716));
    layer2_outputs(4737) <= not((layer1_outputs(6907)) or (layer1_outputs(3057)));
    layer2_outputs(4738) <= layer1_outputs(8360);
    layer2_outputs(4739) <= not((layer1_outputs(8282)) and (layer1_outputs(9834)));
    layer2_outputs(4740) <= not((layer1_outputs(9510)) or (layer1_outputs(5870)));
    layer2_outputs(4741) <= not((layer1_outputs(5949)) and (layer1_outputs(7334)));
    layer2_outputs(4742) <= (layer1_outputs(8333)) and (layer1_outputs(75));
    layer2_outputs(4743) <= (layer1_outputs(6937)) or (layer1_outputs(2808));
    layer2_outputs(4744) <= (layer1_outputs(8196)) and (layer1_outputs(2331));
    layer2_outputs(4745) <= not(layer1_outputs(5158));
    layer2_outputs(4746) <= (layer1_outputs(1452)) and not (layer1_outputs(3836));
    layer2_outputs(4747) <= not(layer1_outputs(829));
    layer2_outputs(4748) <= not(layer1_outputs(653)) or (layer1_outputs(3257));
    layer2_outputs(4749) <= layer1_outputs(3872);
    layer2_outputs(4750) <= (layer1_outputs(7859)) and not (layer1_outputs(4728));
    layer2_outputs(4751) <= layer1_outputs(5296);
    layer2_outputs(4752) <= layer1_outputs(5564);
    layer2_outputs(4753) <= not(layer1_outputs(2582));
    layer2_outputs(4754) <= not((layer1_outputs(8051)) and (layer1_outputs(5890)));
    layer2_outputs(4755) <= layer1_outputs(8997);
    layer2_outputs(4756) <= (layer1_outputs(1744)) and not (layer1_outputs(6707));
    layer2_outputs(4757) <= layer1_outputs(2574);
    layer2_outputs(4758) <= layer1_outputs(189);
    layer2_outputs(4759) <= not(layer1_outputs(1099)) or (layer1_outputs(131));
    layer2_outputs(4760) <= (layer1_outputs(5305)) and not (layer1_outputs(4722));
    layer2_outputs(4761) <= (layer1_outputs(5557)) and (layer1_outputs(7810));
    layer2_outputs(4762) <= layer1_outputs(3786);
    layer2_outputs(4763) <= (layer1_outputs(2847)) or (layer1_outputs(5371));
    layer2_outputs(4764) <= not(layer1_outputs(7017));
    layer2_outputs(4765) <= not((layer1_outputs(6612)) and (layer1_outputs(2137)));
    layer2_outputs(4766) <= not(layer1_outputs(5998));
    layer2_outputs(4767) <= layer1_outputs(6658);
    layer2_outputs(4768) <= (layer1_outputs(6233)) and not (layer1_outputs(3481));
    layer2_outputs(4769) <= not(layer1_outputs(2702));
    layer2_outputs(4770) <= layer1_outputs(9639);
    layer2_outputs(4771) <= (layer1_outputs(5000)) and not (layer1_outputs(1681));
    layer2_outputs(4772) <= layer1_outputs(9539);
    layer2_outputs(4773) <= not(layer1_outputs(1624)) or (layer1_outputs(1654));
    layer2_outputs(4774) <= (layer1_outputs(7374)) xor (layer1_outputs(8685));
    layer2_outputs(4775) <= not(layer1_outputs(782));
    layer2_outputs(4776) <= (layer1_outputs(7477)) xor (layer1_outputs(299));
    layer2_outputs(4777) <= not(layer1_outputs(7041));
    layer2_outputs(4778) <= (layer1_outputs(8305)) and not (layer1_outputs(1387));
    layer2_outputs(4779) <= not(layer1_outputs(3851));
    layer2_outputs(4780) <= '1';
    layer2_outputs(4781) <= not(layer1_outputs(6647));
    layer2_outputs(4782) <= not(layer1_outputs(1180));
    layer2_outputs(4783) <= not((layer1_outputs(1034)) and (layer1_outputs(4450)));
    layer2_outputs(4784) <= (layer1_outputs(1517)) and (layer1_outputs(8362));
    layer2_outputs(4785) <= not(layer1_outputs(141)) or (layer1_outputs(3176));
    layer2_outputs(4786) <= (layer1_outputs(10106)) and (layer1_outputs(2147));
    layer2_outputs(4787) <= not(layer1_outputs(3995)) or (layer1_outputs(1992));
    layer2_outputs(4788) <= not(layer1_outputs(2137)) or (layer1_outputs(9491));
    layer2_outputs(4789) <= not((layer1_outputs(699)) or (layer1_outputs(9130)));
    layer2_outputs(4790) <= layer1_outputs(5028);
    layer2_outputs(4791) <= (layer1_outputs(4664)) and (layer1_outputs(532));
    layer2_outputs(4792) <= not(layer1_outputs(7258));
    layer2_outputs(4793) <= '1';
    layer2_outputs(4794) <= layer1_outputs(4255);
    layer2_outputs(4795) <= (layer1_outputs(7318)) and not (layer1_outputs(9415));
    layer2_outputs(4796) <= not(layer1_outputs(1834)) or (layer1_outputs(10214));
    layer2_outputs(4797) <= '0';
    layer2_outputs(4798) <= layer1_outputs(5797);
    layer2_outputs(4799) <= not(layer1_outputs(7820));
    layer2_outputs(4800) <= '0';
    layer2_outputs(4801) <= not(layer1_outputs(2543));
    layer2_outputs(4802) <= not(layer1_outputs(4374));
    layer2_outputs(4803) <= layer1_outputs(1254);
    layer2_outputs(4804) <= (layer1_outputs(8539)) and (layer1_outputs(255));
    layer2_outputs(4805) <= not(layer1_outputs(273));
    layer2_outputs(4806) <= layer1_outputs(3320);
    layer2_outputs(4807) <= '0';
    layer2_outputs(4808) <= not((layer1_outputs(4075)) xor (layer1_outputs(1980)));
    layer2_outputs(4809) <= not(layer1_outputs(5922));
    layer2_outputs(4810) <= not(layer1_outputs(7003));
    layer2_outputs(4811) <= (layer1_outputs(5399)) and (layer1_outputs(4932));
    layer2_outputs(4812) <= not(layer1_outputs(2482)) or (layer1_outputs(1413));
    layer2_outputs(4813) <= layer1_outputs(606);
    layer2_outputs(4814) <= not(layer1_outputs(5550));
    layer2_outputs(4815) <= layer1_outputs(5602);
    layer2_outputs(4816) <= '1';
    layer2_outputs(4817) <= not((layer1_outputs(7076)) and (layer1_outputs(1642)));
    layer2_outputs(4818) <= (layer1_outputs(4283)) and not (layer1_outputs(2380));
    layer2_outputs(4819) <= layer1_outputs(2625);
    layer2_outputs(4820) <= (layer1_outputs(3161)) and not (layer1_outputs(2577));
    layer2_outputs(4821) <= not(layer1_outputs(9439)) or (layer1_outputs(1254));
    layer2_outputs(4822) <= (layer1_outputs(4231)) or (layer1_outputs(8089));
    layer2_outputs(4823) <= layer1_outputs(7583);
    layer2_outputs(4824) <= not((layer1_outputs(4733)) and (layer1_outputs(8495)));
    layer2_outputs(4825) <= not(layer1_outputs(362));
    layer2_outputs(4826) <= layer1_outputs(8254);
    layer2_outputs(4827) <= (layer1_outputs(68)) and not (layer1_outputs(695));
    layer2_outputs(4828) <= not(layer1_outputs(3932));
    layer2_outputs(4829) <= layer1_outputs(6454);
    layer2_outputs(4830) <= not(layer1_outputs(562));
    layer2_outputs(4831) <= (layer1_outputs(1440)) and (layer1_outputs(4112));
    layer2_outputs(4832) <= not(layer1_outputs(5524));
    layer2_outputs(4833) <= '1';
    layer2_outputs(4834) <= not(layer1_outputs(4620));
    layer2_outputs(4835) <= layer1_outputs(1924);
    layer2_outputs(4836) <= (layer1_outputs(2401)) and not (layer1_outputs(5499));
    layer2_outputs(4837) <= not((layer1_outputs(5729)) and (layer1_outputs(9517)));
    layer2_outputs(4838) <= (layer1_outputs(4151)) xor (layer1_outputs(536));
    layer2_outputs(4839) <= (layer1_outputs(3249)) and (layer1_outputs(2650));
    layer2_outputs(4840) <= not((layer1_outputs(6385)) and (layer1_outputs(4751)));
    layer2_outputs(4841) <= layer1_outputs(5831);
    layer2_outputs(4842) <= not(layer1_outputs(4186)) or (layer1_outputs(1335));
    layer2_outputs(4843) <= '1';
    layer2_outputs(4844) <= (layer1_outputs(106)) and not (layer1_outputs(10218));
    layer2_outputs(4845) <= layer1_outputs(2279);
    layer2_outputs(4846) <= '1';
    layer2_outputs(4847) <= not((layer1_outputs(5252)) or (layer1_outputs(7088)));
    layer2_outputs(4848) <= not(layer1_outputs(7290));
    layer2_outputs(4849) <= '1';
    layer2_outputs(4850) <= layer1_outputs(7197);
    layer2_outputs(4851) <= not(layer1_outputs(1782));
    layer2_outputs(4852) <= not((layer1_outputs(7373)) and (layer1_outputs(5493)));
    layer2_outputs(4853) <= not((layer1_outputs(7384)) or (layer1_outputs(550)));
    layer2_outputs(4854) <= (layer1_outputs(7648)) xor (layer1_outputs(4132));
    layer2_outputs(4855) <= (layer1_outputs(8591)) and (layer1_outputs(6480));
    layer2_outputs(4856) <= not(layer1_outputs(3617)) or (layer1_outputs(5718));
    layer2_outputs(4857) <= (layer1_outputs(6389)) and (layer1_outputs(3207));
    layer2_outputs(4858) <= not(layer1_outputs(9503));
    layer2_outputs(4859) <= not((layer1_outputs(8615)) or (layer1_outputs(5287)));
    layer2_outputs(4860) <= layer1_outputs(6886);
    layer2_outputs(4861) <= layer1_outputs(7302);
    layer2_outputs(4862) <= not((layer1_outputs(4580)) or (layer1_outputs(1376)));
    layer2_outputs(4863) <= layer1_outputs(10207);
    layer2_outputs(4864) <= (layer1_outputs(5744)) xor (layer1_outputs(2521));
    layer2_outputs(4865) <= not(layer1_outputs(857));
    layer2_outputs(4866) <= not((layer1_outputs(8614)) or (layer1_outputs(3560)));
    layer2_outputs(4867) <= not((layer1_outputs(7228)) and (layer1_outputs(4737)));
    layer2_outputs(4868) <= not(layer1_outputs(7246)) or (layer1_outputs(9808));
    layer2_outputs(4869) <= layer1_outputs(3536);
    layer2_outputs(4870) <= (layer1_outputs(9730)) or (layer1_outputs(3411));
    layer2_outputs(4871) <= not(layer1_outputs(3492)) or (layer1_outputs(3498));
    layer2_outputs(4872) <= not(layer1_outputs(7840));
    layer2_outputs(4873) <= not((layer1_outputs(2608)) or (layer1_outputs(3321)));
    layer2_outputs(4874) <= not(layer1_outputs(4737));
    layer2_outputs(4875) <= layer1_outputs(9043);
    layer2_outputs(4876) <= not(layer1_outputs(2029));
    layer2_outputs(4877) <= not(layer1_outputs(8317));
    layer2_outputs(4878) <= not(layer1_outputs(5505)) or (layer1_outputs(4277));
    layer2_outputs(4879) <= (layer1_outputs(6568)) and (layer1_outputs(7721));
    layer2_outputs(4880) <= layer1_outputs(6836);
    layer2_outputs(4881) <= not(layer1_outputs(3396)) or (layer1_outputs(1881));
    layer2_outputs(4882) <= not(layer1_outputs(8269)) or (layer1_outputs(4869));
    layer2_outputs(4883) <= (layer1_outputs(2212)) and (layer1_outputs(7875));
    layer2_outputs(4884) <= '1';
    layer2_outputs(4885) <= not((layer1_outputs(5375)) xor (layer1_outputs(922)));
    layer2_outputs(4886) <= not((layer1_outputs(5984)) and (layer1_outputs(5407)));
    layer2_outputs(4887) <= not(layer1_outputs(764)) or (layer1_outputs(3835));
    layer2_outputs(4888) <= not(layer1_outputs(5494));
    layer2_outputs(4889) <= layer1_outputs(2761);
    layer2_outputs(4890) <= not(layer1_outputs(1122));
    layer2_outputs(4891) <= (layer1_outputs(3309)) and (layer1_outputs(3403));
    layer2_outputs(4892) <= not(layer1_outputs(9343));
    layer2_outputs(4893) <= layer1_outputs(875);
    layer2_outputs(4894) <= not((layer1_outputs(2753)) and (layer1_outputs(4288)));
    layer2_outputs(4895) <= not(layer1_outputs(9266));
    layer2_outputs(4896) <= '1';
    layer2_outputs(4897) <= (layer1_outputs(7644)) and not (layer1_outputs(8391));
    layer2_outputs(4898) <= (layer1_outputs(6031)) and not (layer1_outputs(5118));
    layer2_outputs(4899) <= not(layer1_outputs(782)) or (layer1_outputs(5358));
    layer2_outputs(4900) <= not((layer1_outputs(9765)) xor (layer1_outputs(6887)));
    layer2_outputs(4901) <= not(layer1_outputs(4491));
    layer2_outputs(4902) <= not(layer1_outputs(30));
    layer2_outputs(4903) <= layer1_outputs(7359);
    layer2_outputs(4904) <= '1';
    layer2_outputs(4905) <= layer1_outputs(2491);
    layer2_outputs(4906) <= (layer1_outputs(5650)) and not (layer1_outputs(5701));
    layer2_outputs(4907) <= (layer1_outputs(4103)) and not (layer1_outputs(8633));
    layer2_outputs(4908) <= not((layer1_outputs(2549)) or (layer1_outputs(9009)));
    layer2_outputs(4909) <= not((layer1_outputs(32)) or (layer1_outputs(4957)));
    layer2_outputs(4910) <= not(layer1_outputs(7464));
    layer2_outputs(4911) <= not(layer1_outputs(5769));
    layer2_outputs(4912) <= '1';
    layer2_outputs(4913) <= not(layer1_outputs(8123));
    layer2_outputs(4914) <= (layer1_outputs(155)) or (layer1_outputs(5070));
    layer2_outputs(4915) <= not(layer1_outputs(9237));
    layer2_outputs(4916) <= not((layer1_outputs(64)) and (layer1_outputs(1677)));
    layer2_outputs(4917) <= (layer1_outputs(4347)) and (layer1_outputs(672));
    layer2_outputs(4918) <= not((layer1_outputs(4564)) xor (layer1_outputs(4739)));
    layer2_outputs(4919) <= (layer1_outputs(4370)) and (layer1_outputs(4866));
    layer2_outputs(4920) <= not(layer1_outputs(1099)) or (layer1_outputs(6469));
    layer2_outputs(4921) <= not(layer1_outputs(3893));
    layer2_outputs(4922) <= (layer1_outputs(8225)) and not (layer1_outputs(1025));
    layer2_outputs(4923) <= not(layer1_outputs(2146));
    layer2_outputs(4924) <= layer1_outputs(2248);
    layer2_outputs(4925) <= not((layer1_outputs(2367)) and (layer1_outputs(2526)));
    layer2_outputs(4926) <= '0';
    layer2_outputs(4927) <= (layer1_outputs(7697)) and (layer1_outputs(9052));
    layer2_outputs(4928) <= layer1_outputs(9670);
    layer2_outputs(4929) <= not(layer1_outputs(6186));
    layer2_outputs(4930) <= layer1_outputs(2369);
    layer2_outputs(4931) <= not(layer1_outputs(6719)) or (layer1_outputs(776));
    layer2_outputs(4932) <= not(layer1_outputs(8040));
    layer2_outputs(4933) <= (layer1_outputs(8166)) xor (layer1_outputs(8930));
    layer2_outputs(4934) <= not(layer1_outputs(4326)) or (layer1_outputs(5431));
    layer2_outputs(4935) <= not((layer1_outputs(4381)) or (layer1_outputs(2919)));
    layer2_outputs(4936) <= not(layer1_outputs(7107)) or (layer1_outputs(902));
    layer2_outputs(4937) <= (layer1_outputs(8056)) or (layer1_outputs(6073));
    layer2_outputs(4938) <= not(layer1_outputs(4414));
    layer2_outputs(4939) <= (layer1_outputs(8880)) and (layer1_outputs(5796));
    layer2_outputs(4940) <= layer1_outputs(4913);
    layer2_outputs(4941) <= not(layer1_outputs(4635));
    layer2_outputs(4942) <= not((layer1_outputs(9797)) xor (layer1_outputs(2376)));
    layer2_outputs(4943) <= layer1_outputs(6565);
    layer2_outputs(4944) <= layer1_outputs(7468);
    layer2_outputs(4945) <= (layer1_outputs(9500)) and not (layer1_outputs(3551));
    layer2_outputs(4946) <= not(layer1_outputs(9888));
    layer2_outputs(4947) <= (layer1_outputs(1114)) xor (layer1_outputs(6839));
    layer2_outputs(4948) <= '1';
    layer2_outputs(4949) <= layer1_outputs(3901);
    layer2_outputs(4950) <= not(layer1_outputs(4493));
    layer2_outputs(4951) <= not(layer1_outputs(4041));
    layer2_outputs(4952) <= not((layer1_outputs(6428)) and (layer1_outputs(9386)));
    layer2_outputs(4953) <= not(layer1_outputs(9148));
    layer2_outputs(4954) <= not(layer1_outputs(2453));
    layer2_outputs(4955) <= (layer1_outputs(3487)) or (layer1_outputs(1730));
    layer2_outputs(4956) <= (layer1_outputs(6464)) and (layer1_outputs(2592));
    layer2_outputs(4957) <= not(layer1_outputs(4405));
    layer2_outputs(4958) <= not(layer1_outputs(1145));
    layer2_outputs(4959) <= not(layer1_outputs(9686)) or (layer1_outputs(1908));
    layer2_outputs(4960) <= not((layer1_outputs(8045)) or (layer1_outputs(4709)));
    layer2_outputs(4961) <= '0';
    layer2_outputs(4962) <= layer1_outputs(4016);
    layer2_outputs(4963) <= layer1_outputs(269);
    layer2_outputs(4964) <= not(layer1_outputs(4113));
    layer2_outputs(4965) <= (layer1_outputs(1370)) or (layer1_outputs(1989));
    layer2_outputs(4966) <= (layer1_outputs(1155)) and (layer1_outputs(8587));
    layer2_outputs(4967) <= not((layer1_outputs(6343)) or (layer1_outputs(9624)));
    layer2_outputs(4968) <= not(layer1_outputs(4968)) or (layer1_outputs(4225));
    layer2_outputs(4969) <= not(layer1_outputs(3289));
    layer2_outputs(4970) <= '1';
    layer2_outputs(4971) <= not((layer1_outputs(3854)) or (layer1_outputs(6987)));
    layer2_outputs(4972) <= (layer1_outputs(8101)) and (layer1_outputs(7325));
    layer2_outputs(4973) <= not(layer1_outputs(8198));
    layer2_outputs(4974) <= not(layer1_outputs(5767)) or (layer1_outputs(8404));
    layer2_outputs(4975) <= layer1_outputs(508);
    layer2_outputs(4976) <= not(layer1_outputs(219));
    layer2_outputs(4977) <= not(layer1_outputs(1205)) or (layer1_outputs(2767));
    layer2_outputs(4978) <= '0';
    layer2_outputs(4979) <= (layer1_outputs(15)) or (layer1_outputs(6334));
    layer2_outputs(4980) <= layer1_outputs(3296);
    layer2_outputs(4981) <= layer1_outputs(2474);
    layer2_outputs(4982) <= layer1_outputs(7154);
    layer2_outputs(4983) <= not(layer1_outputs(2242));
    layer2_outputs(4984) <= layer1_outputs(7120);
    layer2_outputs(4985) <= (layer1_outputs(8711)) and (layer1_outputs(2535));
    layer2_outputs(4986) <= not((layer1_outputs(3385)) or (layer1_outputs(7145)));
    layer2_outputs(4987) <= not(layer1_outputs(9229)) or (layer1_outputs(9471));
    layer2_outputs(4988) <= not(layer1_outputs(347));
    layer2_outputs(4989) <= '1';
    layer2_outputs(4990) <= not(layer1_outputs(9507));
    layer2_outputs(4991) <= layer1_outputs(2334);
    layer2_outputs(4992) <= layer1_outputs(7233);
    layer2_outputs(4993) <= layer1_outputs(2974);
    layer2_outputs(4994) <= not((layer1_outputs(4043)) and (layer1_outputs(24)));
    layer2_outputs(4995) <= '0';
    layer2_outputs(4996) <= (layer1_outputs(9126)) xor (layer1_outputs(9469));
    layer2_outputs(4997) <= not(layer1_outputs(10041)) or (layer1_outputs(7905));
    layer2_outputs(4998) <= layer1_outputs(8477);
    layer2_outputs(4999) <= layer1_outputs(6760);
    layer2_outputs(5000) <= not(layer1_outputs(6112)) or (layer1_outputs(6835));
    layer2_outputs(5001) <= not((layer1_outputs(6756)) or (layer1_outputs(6054)));
    layer2_outputs(5002) <= not((layer1_outputs(3574)) xor (layer1_outputs(824)));
    layer2_outputs(5003) <= not(layer1_outputs(4611));
    layer2_outputs(5004) <= not((layer1_outputs(1410)) and (layer1_outputs(2448)));
    layer2_outputs(5005) <= '0';
    layer2_outputs(5006) <= not((layer1_outputs(6393)) and (layer1_outputs(2729)));
    layer2_outputs(5007) <= not(layer1_outputs(81));
    layer2_outputs(5008) <= not((layer1_outputs(3117)) and (layer1_outputs(8383)));
    layer2_outputs(5009) <= not((layer1_outputs(5175)) or (layer1_outputs(5651)));
    layer2_outputs(5010) <= not(layer1_outputs(8754)) or (layer1_outputs(8885));
    layer2_outputs(5011) <= not(layer1_outputs(1051));
    layer2_outputs(5012) <= not((layer1_outputs(1731)) and (layer1_outputs(9517)));
    layer2_outputs(5013) <= not(layer1_outputs(897));
    layer2_outputs(5014) <= not(layer1_outputs(6681));
    layer2_outputs(5015) <= not(layer1_outputs(1961)) or (layer1_outputs(3963));
    layer2_outputs(5016) <= not((layer1_outputs(7512)) and (layer1_outputs(2411)));
    layer2_outputs(5017) <= '0';
    layer2_outputs(5018) <= '1';
    layer2_outputs(5019) <= (layer1_outputs(3983)) or (layer1_outputs(1227));
    layer2_outputs(5020) <= layer1_outputs(4632);
    layer2_outputs(5021) <= (layer1_outputs(5440)) and not (layer1_outputs(9211));
    layer2_outputs(5022) <= not(layer1_outputs(9665)) or (layer1_outputs(4101));
    layer2_outputs(5023) <= not(layer1_outputs(6976));
    layer2_outputs(5024) <= layer1_outputs(448);
    layer2_outputs(5025) <= not(layer1_outputs(4511)) or (layer1_outputs(344));
    layer2_outputs(5026) <= layer1_outputs(308);
    layer2_outputs(5027) <= not((layer1_outputs(3123)) and (layer1_outputs(5037)));
    layer2_outputs(5028) <= '1';
    layer2_outputs(5029) <= not(layer1_outputs(1308)) or (layer1_outputs(3563));
    layer2_outputs(5030) <= not(layer1_outputs(2672));
    layer2_outputs(5031) <= (layer1_outputs(4646)) and (layer1_outputs(7948));
    layer2_outputs(5032) <= (layer1_outputs(1297)) and not (layer1_outputs(2112));
    layer2_outputs(5033) <= (layer1_outputs(2578)) or (layer1_outputs(364));
    layer2_outputs(5034) <= not(layer1_outputs(5188));
    layer2_outputs(5035) <= (layer1_outputs(6153)) and not (layer1_outputs(941));
    layer2_outputs(5036) <= not(layer1_outputs(4332));
    layer2_outputs(5037) <= '1';
    layer2_outputs(5038) <= (layer1_outputs(10008)) and not (layer1_outputs(2279));
    layer2_outputs(5039) <= layer1_outputs(10006);
    layer2_outputs(5040) <= layer1_outputs(6226);
    layer2_outputs(5041) <= (layer1_outputs(9487)) xor (layer1_outputs(8246));
    layer2_outputs(5042) <= not((layer1_outputs(3502)) or (layer1_outputs(3743)));
    layer2_outputs(5043) <= not(layer1_outputs(9753)) or (layer1_outputs(8520));
    layer2_outputs(5044) <= not(layer1_outputs(2582));
    layer2_outputs(5045) <= not((layer1_outputs(5240)) or (layer1_outputs(319)));
    layer2_outputs(5046) <= (layer1_outputs(9922)) and not (layer1_outputs(4555));
    layer2_outputs(5047) <= not(layer1_outputs(5417)) or (layer1_outputs(6651));
    layer2_outputs(5048) <= not((layer1_outputs(8631)) and (layer1_outputs(6896)));
    layer2_outputs(5049) <= layer1_outputs(2675);
    layer2_outputs(5050) <= (layer1_outputs(8238)) and not (layer1_outputs(8308));
    layer2_outputs(5051) <= (layer1_outputs(6599)) and (layer1_outputs(2503));
    layer2_outputs(5052) <= (layer1_outputs(1157)) and not (layer1_outputs(4156));
    layer2_outputs(5053) <= (layer1_outputs(5069)) or (layer1_outputs(1743));
    layer2_outputs(5054) <= (layer1_outputs(2661)) xor (layer1_outputs(5657));
    layer2_outputs(5055) <= not(layer1_outputs(9433));
    layer2_outputs(5056) <= layer1_outputs(4519);
    layer2_outputs(5057) <= (layer1_outputs(2755)) and (layer1_outputs(6384));
    layer2_outputs(5058) <= not(layer1_outputs(636)) or (layer1_outputs(4017));
    layer2_outputs(5059) <= layer1_outputs(5602);
    layer2_outputs(5060) <= layer1_outputs(3722);
    layer2_outputs(5061) <= not(layer1_outputs(8976));
    layer2_outputs(5062) <= layer1_outputs(3138);
    layer2_outputs(5063) <= not(layer1_outputs(3850));
    layer2_outputs(5064) <= layer1_outputs(5392);
    layer2_outputs(5065) <= not(layer1_outputs(4730));
    layer2_outputs(5066) <= '1';
    layer2_outputs(5067) <= layer1_outputs(1208);
    layer2_outputs(5068) <= not(layer1_outputs(7549));
    layer2_outputs(5069) <= not((layer1_outputs(4150)) or (layer1_outputs(2192)));
    layer2_outputs(5070) <= (layer1_outputs(5815)) and (layer1_outputs(3966));
    layer2_outputs(5071) <= (layer1_outputs(9278)) and not (layer1_outputs(10105));
    layer2_outputs(5072) <= layer1_outputs(3001);
    layer2_outputs(5073) <= layer1_outputs(3642);
    layer2_outputs(5074) <= not(layer1_outputs(6491));
    layer2_outputs(5075) <= not(layer1_outputs(5439));
    layer2_outputs(5076) <= not(layer1_outputs(9594)) or (layer1_outputs(7610));
    layer2_outputs(5077) <= not(layer1_outputs(8890));
    layer2_outputs(5078) <= (layer1_outputs(9959)) and not (layer1_outputs(9656));
    layer2_outputs(5079) <= '0';
    layer2_outputs(5080) <= not((layer1_outputs(7630)) or (layer1_outputs(6496)));
    layer2_outputs(5081) <= '1';
    layer2_outputs(5082) <= '0';
    layer2_outputs(5083) <= (layer1_outputs(6377)) or (layer1_outputs(8808));
    layer2_outputs(5084) <= not((layer1_outputs(6268)) or (layer1_outputs(6430)));
    layer2_outputs(5085) <= not(layer1_outputs(2205));
    layer2_outputs(5086) <= '0';
    layer2_outputs(5087) <= layer1_outputs(1757);
    layer2_outputs(5088) <= (layer1_outputs(5297)) and not (layer1_outputs(6359));
    layer2_outputs(5089) <= not(layer1_outputs(4833)) or (layer1_outputs(9398));
    layer2_outputs(5090) <= layer1_outputs(7104);
    layer2_outputs(5091) <= (layer1_outputs(1132)) and not (layer1_outputs(8154));
    layer2_outputs(5092) <= layer1_outputs(5837);
    layer2_outputs(5093) <= not(layer1_outputs(231)) or (layer1_outputs(6313));
    layer2_outputs(5094) <= layer1_outputs(6698);
    layer2_outputs(5095) <= (layer1_outputs(3610)) and not (layer1_outputs(3197));
    layer2_outputs(5096) <= (layer1_outputs(775)) and (layer1_outputs(9530));
    layer2_outputs(5097) <= not(layer1_outputs(6665));
    layer2_outputs(5098) <= '1';
    layer2_outputs(5099) <= not(layer1_outputs(2456));
    layer2_outputs(5100) <= not(layer1_outputs(9666));
    layer2_outputs(5101) <= (layer1_outputs(2081)) and not (layer1_outputs(3366));
    layer2_outputs(5102) <= layer1_outputs(7657);
    layer2_outputs(5103) <= layer1_outputs(9970);
    layer2_outputs(5104) <= not(layer1_outputs(6043));
    layer2_outputs(5105) <= (layer1_outputs(595)) and not (layer1_outputs(9914));
    layer2_outputs(5106) <= layer1_outputs(6999);
    layer2_outputs(5107) <= (layer1_outputs(7428)) and not (layer1_outputs(9810));
    layer2_outputs(5108) <= (layer1_outputs(513)) and not (layer1_outputs(3333));
    layer2_outputs(5109) <= not(layer1_outputs(3833));
    layer2_outputs(5110) <= layer1_outputs(3827);
    layer2_outputs(5111) <= '0';
    layer2_outputs(5112) <= layer1_outputs(8746);
    layer2_outputs(5113) <= (layer1_outputs(8140)) and not (layer1_outputs(1042));
    layer2_outputs(5114) <= (layer1_outputs(1591)) and not (layer1_outputs(9396));
    layer2_outputs(5115) <= not((layer1_outputs(4984)) or (layer1_outputs(7330)));
    layer2_outputs(5116) <= (layer1_outputs(8550)) and not (layer1_outputs(8812));
    layer2_outputs(5117) <= not(layer1_outputs(5089));
    layer2_outputs(5118) <= '0';
    layer2_outputs(5119) <= not((layer1_outputs(7078)) xor (layer1_outputs(6593)));
    layer2_outputs(5120) <= (layer1_outputs(7311)) and (layer1_outputs(5540));
    layer2_outputs(5121) <= not(layer1_outputs(3848));
    layer2_outputs(5122) <= layer1_outputs(9498);
    layer2_outputs(5123) <= not(layer1_outputs(4523));
    layer2_outputs(5124) <= not(layer1_outputs(3553));
    layer2_outputs(5125) <= layer1_outputs(2621);
    layer2_outputs(5126) <= layer1_outputs(5248);
    layer2_outputs(5127) <= (layer1_outputs(47)) and not (layer1_outputs(9779));
    layer2_outputs(5128) <= not(layer1_outputs(5314));
    layer2_outputs(5129) <= not((layer1_outputs(5345)) and (layer1_outputs(9042)));
    layer2_outputs(5130) <= layer1_outputs(121);
    layer2_outputs(5131) <= not(layer1_outputs(1563));
    layer2_outputs(5132) <= (layer1_outputs(5076)) or (layer1_outputs(9257));
    layer2_outputs(5133) <= (layer1_outputs(6761)) xor (layer1_outputs(5939));
    layer2_outputs(5134) <= layer1_outputs(838);
    layer2_outputs(5135) <= (layer1_outputs(1033)) or (layer1_outputs(9361));
    layer2_outputs(5136) <= not(layer1_outputs(2132)) or (layer1_outputs(4977));
    layer2_outputs(5137) <= not(layer1_outputs(6872)) or (layer1_outputs(9288));
    layer2_outputs(5138) <= not((layer1_outputs(6327)) or (layer1_outputs(4710)));
    layer2_outputs(5139) <= (layer1_outputs(4578)) and (layer1_outputs(3308));
    layer2_outputs(5140) <= not(layer1_outputs(194));
    layer2_outputs(5141) <= not(layer1_outputs(649));
    layer2_outputs(5142) <= (layer1_outputs(3757)) and not (layer1_outputs(9464));
    layer2_outputs(5143) <= layer1_outputs(5216);
    layer2_outputs(5144) <= layer1_outputs(7918);
    layer2_outputs(5145) <= not(layer1_outputs(7259)) or (layer1_outputs(2655));
    layer2_outputs(5146) <= not(layer1_outputs(5979));
    layer2_outputs(5147) <= layer1_outputs(3622);
    layer2_outputs(5148) <= not(layer1_outputs(1852));
    layer2_outputs(5149) <= not(layer1_outputs(5542));
    layer2_outputs(5150) <= not(layer1_outputs(6767));
    layer2_outputs(5151) <= not(layer1_outputs(6215));
    layer2_outputs(5152) <= not(layer1_outputs(9349));
    layer2_outputs(5153) <= not(layer1_outputs(1473));
    layer2_outputs(5154) <= layer1_outputs(1212);
    layer2_outputs(5155) <= (layer1_outputs(1188)) and not (layer1_outputs(7497));
    layer2_outputs(5156) <= layer1_outputs(9426);
    layer2_outputs(5157) <= layer1_outputs(1283);
    layer2_outputs(5158) <= layer1_outputs(9190);
    layer2_outputs(5159) <= not((layer1_outputs(1481)) and (layer1_outputs(9044)));
    layer2_outputs(5160) <= not(layer1_outputs(1439)) or (layer1_outputs(8277));
    layer2_outputs(5161) <= not(layer1_outputs(8602));
    layer2_outputs(5162) <= not(layer1_outputs(716));
    layer2_outputs(5163) <= not((layer1_outputs(2360)) and (layer1_outputs(4359)));
    layer2_outputs(5164) <= not((layer1_outputs(8457)) or (layer1_outputs(154)));
    layer2_outputs(5165) <= not(layer1_outputs(5102));
    layer2_outputs(5166) <= layer1_outputs(3521);
    layer2_outputs(5167) <= not(layer1_outputs(3764));
    layer2_outputs(5168) <= not(layer1_outputs(7737));
    layer2_outputs(5169) <= not(layer1_outputs(3721));
    layer2_outputs(5170) <= (layer1_outputs(1800)) or (layer1_outputs(9262));
    layer2_outputs(5171) <= not(layer1_outputs(6782));
    layer2_outputs(5172) <= not(layer1_outputs(2583)) or (layer1_outputs(8071));
    layer2_outputs(5173) <= (layer1_outputs(8061)) and (layer1_outputs(3008));
    layer2_outputs(5174) <= '1';
    layer2_outputs(5175) <= not(layer1_outputs(3862));
    layer2_outputs(5176) <= layer1_outputs(8164);
    layer2_outputs(5177) <= layer1_outputs(8417);
    layer2_outputs(5178) <= not(layer1_outputs(4596)) or (layer1_outputs(7400));
    layer2_outputs(5179) <= not((layer1_outputs(9744)) and (layer1_outputs(8497)));
    layer2_outputs(5180) <= layer1_outputs(8053);
    layer2_outputs(5181) <= not(layer1_outputs(7673));
    layer2_outputs(5182) <= (layer1_outputs(7885)) and not (layer1_outputs(7668));
    layer2_outputs(5183) <= layer1_outputs(4492);
    layer2_outputs(5184) <= '1';
    layer2_outputs(5185) <= layer1_outputs(7485);
    layer2_outputs(5186) <= (layer1_outputs(5254)) and (layer1_outputs(235));
    layer2_outputs(5187) <= layer1_outputs(5195);
    layer2_outputs(5188) <= '0';
    layer2_outputs(5189) <= layer1_outputs(7302);
    layer2_outputs(5190) <= layer1_outputs(314);
    layer2_outputs(5191) <= not(layer1_outputs(5567)) or (layer1_outputs(5434));
    layer2_outputs(5192) <= not(layer1_outputs(8912)) or (layer1_outputs(4162));
    layer2_outputs(5193) <= not(layer1_outputs(3977));
    layer2_outputs(5194) <= (layer1_outputs(8714)) and not (layer1_outputs(4108));
    layer2_outputs(5195) <= layer1_outputs(272);
    layer2_outputs(5196) <= (layer1_outputs(7848)) and (layer1_outputs(913));
    layer2_outputs(5197) <= not((layer1_outputs(9807)) xor (layer1_outputs(6073)));
    layer2_outputs(5198) <= not(layer1_outputs(5311));
    layer2_outputs(5199) <= '0';
    layer2_outputs(5200) <= layer1_outputs(15);
    layer2_outputs(5201) <= '1';
    layer2_outputs(5202) <= layer1_outputs(8984);
    layer2_outputs(5203) <= layer1_outputs(1444);
    layer2_outputs(5204) <= not(layer1_outputs(3163)) or (layer1_outputs(6675));
    layer2_outputs(5205) <= layer1_outputs(5681);
    layer2_outputs(5206) <= not(layer1_outputs(1983));
    layer2_outputs(5207) <= not(layer1_outputs(6720));
    layer2_outputs(5208) <= (layer1_outputs(3116)) or (layer1_outputs(7774));
    layer2_outputs(5209) <= not(layer1_outputs(6168));
    layer2_outputs(5210) <= layer1_outputs(7031);
    layer2_outputs(5211) <= not((layer1_outputs(8699)) or (layer1_outputs(6541)));
    layer2_outputs(5212) <= not((layer1_outputs(5008)) and (layer1_outputs(9112)));
    layer2_outputs(5213) <= not((layer1_outputs(1475)) and (layer1_outputs(9281)));
    layer2_outputs(5214) <= not(layer1_outputs(4350));
    layer2_outputs(5215) <= (layer1_outputs(7765)) xor (layer1_outputs(4304));
    layer2_outputs(5216) <= (layer1_outputs(3335)) or (layer1_outputs(547));
    layer2_outputs(5217) <= not(layer1_outputs(5823)) or (layer1_outputs(10215));
    layer2_outputs(5218) <= layer1_outputs(4154);
    layer2_outputs(5219) <= not(layer1_outputs(3375));
    layer2_outputs(5220) <= (layer1_outputs(2393)) and not (layer1_outputs(4658));
    layer2_outputs(5221) <= (layer1_outputs(7978)) and (layer1_outputs(1721));
    layer2_outputs(5222) <= not(layer1_outputs(5857));
    layer2_outputs(5223) <= (layer1_outputs(5178)) or (layer1_outputs(5108));
    layer2_outputs(5224) <= not(layer1_outputs(5329));
    layer2_outputs(5225) <= not(layer1_outputs(3323));
    layer2_outputs(5226) <= layer1_outputs(5969);
    layer2_outputs(5227) <= (layer1_outputs(1745)) or (layer1_outputs(2409));
    layer2_outputs(5228) <= (layer1_outputs(1258)) xor (layer1_outputs(4966));
    layer2_outputs(5229) <= '0';
    layer2_outputs(5230) <= (layer1_outputs(4180)) or (layer1_outputs(6330));
    layer2_outputs(5231) <= layer1_outputs(542);
    layer2_outputs(5232) <= (layer1_outputs(3445)) and not (layer1_outputs(820));
    layer2_outputs(5233) <= not(layer1_outputs(2631));
    layer2_outputs(5234) <= not((layer1_outputs(2942)) and (layer1_outputs(720)));
    layer2_outputs(5235) <= (layer1_outputs(5202)) and not (layer1_outputs(9969));
    layer2_outputs(5236) <= layer1_outputs(2304);
    layer2_outputs(5237) <= not((layer1_outputs(5050)) xor (layer1_outputs(815)));
    layer2_outputs(5238) <= (layer1_outputs(8299)) and not (layer1_outputs(2191));
    layer2_outputs(5239) <= layer1_outputs(3059);
    layer2_outputs(5240) <= (layer1_outputs(2837)) or (layer1_outputs(4369));
    layer2_outputs(5241) <= layer1_outputs(6701);
    layer2_outputs(5242) <= (layer1_outputs(9493)) and not (layer1_outputs(5869));
    layer2_outputs(5243) <= not(layer1_outputs(8174));
    layer2_outputs(5244) <= layer1_outputs(1873);
    layer2_outputs(5245) <= not((layer1_outputs(4753)) or (layer1_outputs(7962)));
    layer2_outputs(5246) <= layer1_outputs(2042);
    layer2_outputs(5247) <= layer1_outputs(4874);
    layer2_outputs(5248) <= layer1_outputs(5805);
    layer2_outputs(5249) <= not((layer1_outputs(645)) or (layer1_outputs(2089)));
    layer2_outputs(5250) <= layer1_outputs(970);
    layer2_outputs(5251) <= not((layer1_outputs(2134)) or (layer1_outputs(5703)));
    layer2_outputs(5252) <= (layer1_outputs(1361)) and not (layer1_outputs(3510));
    layer2_outputs(5253) <= not((layer1_outputs(425)) or (layer1_outputs(1041)));
    layer2_outputs(5254) <= layer1_outputs(3201);
    layer2_outputs(5255) <= not((layer1_outputs(4706)) or (layer1_outputs(1252)));
    layer2_outputs(5256) <= not((layer1_outputs(1377)) xor (layer1_outputs(6201)));
    layer2_outputs(5257) <= not((layer1_outputs(5144)) or (layer1_outputs(4409)));
    layer2_outputs(5258) <= (layer1_outputs(8494)) xor (layer1_outputs(4325));
    layer2_outputs(5259) <= (layer1_outputs(4200)) and not (layer1_outputs(4842));
    layer2_outputs(5260) <= not(layer1_outputs(225));
    layer2_outputs(5261) <= layer1_outputs(2768);
    layer2_outputs(5262) <= (layer1_outputs(2094)) and not (layer1_outputs(2026));
    layer2_outputs(5263) <= not(layer1_outputs(4228));
    layer2_outputs(5264) <= not((layer1_outputs(6562)) or (layer1_outputs(9541)));
    layer2_outputs(5265) <= (layer1_outputs(506)) and not (layer1_outputs(2768));
    layer2_outputs(5266) <= (layer1_outputs(4876)) xor (layer1_outputs(3494));
    layer2_outputs(5267) <= not(layer1_outputs(5611)) or (layer1_outputs(1506));
    layer2_outputs(5268) <= not(layer1_outputs(6686)) or (layer1_outputs(965));
    layer2_outputs(5269) <= layer1_outputs(1883);
    layer2_outputs(5270) <= not(layer1_outputs(4548)) or (layer1_outputs(199));
    layer2_outputs(5271) <= layer1_outputs(9493);
    layer2_outputs(5272) <= not(layer1_outputs(8407));
    layer2_outputs(5273) <= (layer1_outputs(672)) and (layer1_outputs(3607));
    layer2_outputs(5274) <= (layer1_outputs(6266)) and (layer1_outputs(2235));
    layer2_outputs(5275) <= not(layer1_outputs(7726)) or (layer1_outputs(5466));
    layer2_outputs(5276) <= '0';
    layer2_outputs(5277) <= not((layer1_outputs(2655)) and (layer1_outputs(2344)));
    layer2_outputs(5278) <= (layer1_outputs(6961)) or (layer1_outputs(8030));
    layer2_outputs(5279) <= layer1_outputs(3260);
    layer2_outputs(5280) <= not((layer1_outputs(473)) and (layer1_outputs(8990)));
    layer2_outputs(5281) <= (layer1_outputs(122)) xor (layer1_outputs(108));
    layer2_outputs(5282) <= not((layer1_outputs(5463)) xor (layer1_outputs(4022)));
    layer2_outputs(5283) <= not(layer1_outputs(3878)) or (layer1_outputs(5702));
    layer2_outputs(5284) <= not(layer1_outputs(2608));
    layer2_outputs(5285) <= not((layer1_outputs(1987)) xor (layer1_outputs(10119)));
    layer2_outputs(5286) <= (layer1_outputs(4616)) or (layer1_outputs(1786));
    layer2_outputs(5287) <= not(layer1_outputs(3741));
    layer2_outputs(5288) <= not((layer1_outputs(5879)) and (layer1_outputs(3753)));
    layer2_outputs(5289) <= layer1_outputs(1455);
    layer2_outputs(5290) <= not(layer1_outputs(8358));
    layer2_outputs(5291) <= layer1_outputs(5059);
    layer2_outputs(5292) <= not(layer1_outputs(1150));
    layer2_outputs(5293) <= (layer1_outputs(4031)) xor (layer1_outputs(3814));
    layer2_outputs(5294) <= not(layer1_outputs(6596)) or (layer1_outputs(6315));
    layer2_outputs(5295) <= not(layer1_outputs(2651));
    layer2_outputs(5296) <= layer1_outputs(9414);
    layer2_outputs(5297) <= not((layer1_outputs(534)) and (layer1_outputs(7262)));
    layer2_outputs(5298) <= not(layer1_outputs(4685));
    layer2_outputs(5299) <= (layer1_outputs(6032)) and not (layer1_outputs(8663));
    layer2_outputs(5300) <= layer1_outputs(7051);
    layer2_outputs(5301) <= (layer1_outputs(7213)) and not (layer1_outputs(2447));
    layer2_outputs(5302) <= not(layer1_outputs(769));
    layer2_outputs(5303) <= not(layer1_outputs(1602));
    layer2_outputs(5304) <= layer1_outputs(9494);
    layer2_outputs(5305) <= not(layer1_outputs(1485));
    layer2_outputs(5306) <= (layer1_outputs(10179)) and (layer1_outputs(5613));
    layer2_outputs(5307) <= not(layer1_outputs(6503));
    layer2_outputs(5308) <= not((layer1_outputs(1142)) xor (layer1_outputs(5619)));
    layer2_outputs(5309) <= layer1_outputs(7792);
    layer2_outputs(5310) <= not((layer1_outputs(3150)) xor (layer1_outputs(927)));
    layer2_outputs(5311) <= layer1_outputs(435);
    layer2_outputs(5312) <= not(layer1_outputs(326)) or (layer1_outputs(9491));
    layer2_outputs(5313) <= not(layer1_outputs(4143));
    layer2_outputs(5314) <= (layer1_outputs(7532)) and (layer1_outputs(7288));
    layer2_outputs(5315) <= layer1_outputs(2228);
    layer2_outputs(5316) <= not(layer1_outputs(395)) or (layer1_outputs(4367));
    layer2_outputs(5317) <= (layer1_outputs(6020)) and not (layer1_outputs(8422));
    layer2_outputs(5318) <= not(layer1_outputs(9162));
    layer2_outputs(5319) <= not((layer1_outputs(9774)) and (layer1_outputs(8482)));
    layer2_outputs(5320) <= not(layer1_outputs(2251)) or (layer1_outputs(5009));
    layer2_outputs(5321) <= layer1_outputs(4614);
    layer2_outputs(5322) <= not((layer1_outputs(3253)) and (layer1_outputs(4696)));
    layer2_outputs(5323) <= layer1_outputs(6374);
    layer2_outputs(5324) <= layer1_outputs(8874);
    layer2_outputs(5325) <= not(layer1_outputs(9654));
    layer2_outputs(5326) <= not(layer1_outputs(1330)) or (layer1_outputs(6440));
    layer2_outputs(5327) <= not(layer1_outputs(3581));
    layer2_outputs(5328) <= (layer1_outputs(536)) and not (layer1_outputs(7809));
    layer2_outputs(5329) <= layer1_outputs(2066);
    layer2_outputs(5330) <= not(layer1_outputs(5398));
    layer2_outputs(5331) <= layer1_outputs(3944);
    layer2_outputs(5332) <= layer1_outputs(1349);
    layer2_outputs(5333) <= (layer1_outputs(2136)) and not (layer1_outputs(7083));
    layer2_outputs(5334) <= (layer1_outputs(9935)) or (layer1_outputs(7976));
    layer2_outputs(5335) <= (layer1_outputs(6082)) and not (layer1_outputs(4130));
    layer2_outputs(5336) <= not((layer1_outputs(637)) or (layer1_outputs(452)));
    layer2_outputs(5337) <= not(layer1_outputs(3017)) or (layer1_outputs(2864));
    layer2_outputs(5338) <= not(layer1_outputs(3712)) or (layer1_outputs(5256));
    layer2_outputs(5339) <= layer1_outputs(1601);
    layer2_outputs(5340) <= not(layer1_outputs(10088)) or (layer1_outputs(7397));
    layer2_outputs(5341) <= not(layer1_outputs(1640)) or (layer1_outputs(4110));
    layer2_outputs(5342) <= not((layer1_outputs(6915)) and (layer1_outputs(2147)));
    layer2_outputs(5343) <= layer1_outputs(8507);
    layer2_outputs(5344) <= layer1_outputs(2902);
    layer2_outputs(5345) <= (layer1_outputs(4061)) and not (layer1_outputs(5874));
    layer2_outputs(5346) <= not(layer1_outputs(3357)) or (layer1_outputs(5215));
    layer2_outputs(5347) <= (layer1_outputs(4344)) and not (layer1_outputs(4731));
    layer2_outputs(5348) <= layer1_outputs(93);
    layer2_outputs(5349) <= layer1_outputs(9676);
    layer2_outputs(5350) <= not(layer1_outputs(3945));
    layer2_outputs(5351) <= '1';
    layer2_outputs(5352) <= not((layer1_outputs(1261)) xor (layer1_outputs(3935)));
    layer2_outputs(5353) <= not((layer1_outputs(4309)) or (layer1_outputs(4089)));
    layer2_outputs(5354) <= (layer1_outputs(9843)) xor (layer1_outputs(4642));
    layer2_outputs(5355) <= '1';
    layer2_outputs(5356) <= not(layer1_outputs(3065)) or (layer1_outputs(772));
    layer2_outputs(5357) <= (layer1_outputs(9317)) and (layer1_outputs(6697));
    layer2_outputs(5358) <= not((layer1_outputs(5535)) xor (layer1_outputs(49)));
    layer2_outputs(5359) <= (layer1_outputs(3576)) xor (layer1_outputs(8724));
    layer2_outputs(5360) <= (layer1_outputs(4047)) and not (layer1_outputs(3535));
    layer2_outputs(5361) <= not(layer1_outputs(9777));
    layer2_outputs(5362) <= not(layer1_outputs(9142));
    layer2_outputs(5363) <= layer1_outputs(7455);
    layer2_outputs(5364) <= '1';
    layer2_outputs(5365) <= (layer1_outputs(9746)) or (layer1_outputs(4779));
    layer2_outputs(5366) <= not((layer1_outputs(3025)) or (layer1_outputs(7142)));
    layer2_outputs(5367) <= (layer1_outputs(832)) or (layer1_outputs(6463));
    layer2_outputs(5368) <= not((layer1_outputs(5497)) or (layer1_outputs(3382)));
    layer2_outputs(5369) <= not(layer1_outputs(3483));
    layer2_outputs(5370) <= (layer1_outputs(5195)) and (layer1_outputs(8070));
    layer2_outputs(5371) <= layer1_outputs(6213);
    layer2_outputs(5372) <= (layer1_outputs(2900)) or (layer1_outputs(7172));
    layer2_outputs(5373) <= not(layer1_outputs(7312));
    layer2_outputs(5374) <= layer1_outputs(6450);
    layer2_outputs(5375) <= layer1_outputs(6733);
    layer2_outputs(5376) <= layer1_outputs(1986);
    layer2_outputs(5377) <= '1';
    layer2_outputs(5378) <= (layer1_outputs(7165)) and not (layer1_outputs(2751));
    layer2_outputs(5379) <= '1';
    layer2_outputs(5380) <= not(layer1_outputs(3365));
    layer2_outputs(5381) <= layer1_outputs(6554);
    layer2_outputs(5382) <= not(layer1_outputs(7077)) or (layer1_outputs(35));
    layer2_outputs(5383) <= layer1_outputs(5740);
    layer2_outputs(5384) <= '0';
    layer2_outputs(5385) <= not(layer1_outputs(8213)) or (layer1_outputs(2944));
    layer2_outputs(5386) <= not(layer1_outputs(3553));
    layer2_outputs(5387) <= (layer1_outputs(8722)) or (layer1_outputs(1334));
    layer2_outputs(5388) <= layer1_outputs(107);
    layer2_outputs(5389) <= layer1_outputs(9083);
    layer2_outputs(5390) <= not(layer1_outputs(1943)) or (layer1_outputs(7527));
    layer2_outputs(5391) <= not((layer1_outputs(7767)) and (layer1_outputs(10017)));
    layer2_outputs(5392) <= (layer1_outputs(3907)) and not (layer1_outputs(4439));
    layer2_outputs(5393) <= layer1_outputs(10036);
    layer2_outputs(5394) <= (layer1_outputs(9502)) and (layer1_outputs(3541));
    layer2_outputs(5395) <= layer1_outputs(1093);
    layer2_outputs(5396) <= '0';
    layer2_outputs(5397) <= not(layer1_outputs(9659));
    layer2_outputs(5398) <= not(layer1_outputs(1361)) or (layer1_outputs(8584));
    layer2_outputs(5399) <= (layer1_outputs(10133)) and not (layer1_outputs(2850));
    layer2_outputs(5400) <= not(layer1_outputs(2431)) or (layer1_outputs(9346));
    layer2_outputs(5401) <= not(layer1_outputs(4575)) or (layer1_outputs(751));
    layer2_outputs(5402) <= not(layer1_outputs(5842)) or (layer1_outputs(8466));
    layer2_outputs(5403) <= not(layer1_outputs(1484));
    layer2_outputs(5404) <= (layer1_outputs(9435)) or (layer1_outputs(5498));
    layer2_outputs(5405) <= (layer1_outputs(879)) or (layer1_outputs(1927));
    layer2_outputs(5406) <= '1';
    layer2_outputs(5407) <= not((layer1_outputs(2793)) or (layer1_outputs(3144)));
    layer2_outputs(5408) <= (layer1_outputs(767)) or (layer1_outputs(2846));
    layer2_outputs(5409) <= not(layer1_outputs(10211));
    layer2_outputs(5410) <= '0';
    layer2_outputs(5411) <= (layer1_outputs(1296)) and (layer1_outputs(670));
    layer2_outputs(5412) <= layer1_outputs(5691);
    layer2_outputs(5413) <= '1';
    layer2_outputs(5414) <= layer1_outputs(8146);
    layer2_outputs(5415) <= layer1_outputs(822);
    layer2_outputs(5416) <= (layer1_outputs(6811)) and not (layer1_outputs(1120));
    layer2_outputs(5417) <= not(layer1_outputs(6188));
    layer2_outputs(5418) <= '0';
    layer2_outputs(5419) <= layer1_outputs(9628);
    layer2_outputs(5420) <= (layer1_outputs(2222)) and not (layer1_outputs(5704));
    layer2_outputs(5421) <= (layer1_outputs(1336)) or (layer1_outputs(9467));
    layer2_outputs(5422) <= not(layer1_outputs(7092));
    layer2_outputs(5423) <= not((layer1_outputs(3416)) xor (layer1_outputs(9927)));
    layer2_outputs(5424) <= not(layer1_outputs(2188)) or (layer1_outputs(7215));
    layer2_outputs(5425) <= not(layer1_outputs(1703));
    layer2_outputs(5426) <= not((layer1_outputs(7649)) xor (layer1_outputs(10163)));
    layer2_outputs(5427) <= layer1_outputs(5277);
    layer2_outputs(5428) <= layer1_outputs(4755);
    layer2_outputs(5429) <= layer1_outputs(3727);
    layer2_outputs(5430) <= not(layer1_outputs(2208));
    layer2_outputs(5431) <= (layer1_outputs(1707)) and (layer1_outputs(1711));
    layer2_outputs(5432) <= not(layer1_outputs(4844));
    layer2_outputs(5433) <= (layer1_outputs(2948)) and not (layer1_outputs(2885));
    layer2_outputs(5434) <= (layer1_outputs(1545)) or (layer1_outputs(5432));
    layer2_outputs(5435) <= '0';
    layer2_outputs(5436) <= not(layer1_outputs(5836));
    layer2_outputs(5437) <= not(layer1_outputs(1346));
    layer2_outputs(5438) <= '1';
    layer2_outputs(5439) <= not(layer1_outputs(8661));
    layer2_outputs(5440) <= (layer1_outputs(1126)) and not (layer1_outputs(8043));
    layer2_outputs(5441) <= layer1_outputs(613);
    layer2_outputs(5442) <= not(layer1_outputs(1151)) or (layer1_outputs(7691));
    layer2_outputs(5443) <= layer1_outputs(2964);
    layer2_outputs(5444) <= layer1_outputs(9524);
    layer2_outputs(5445) <= not((layer1_outputs(5560)) and (layer1_outputs(6467)));
    layer2_outputs(5446) <= layer1_outputs(10);
    layer2_outputs(5447) <= not(layer1_outputs(5926)) or (layer1_outputs(3725));
    layer2_outputs(5448) <= not((layer1_outputs(2097)) or (layer1_outputs(1850)));
    layer2_outputs(5449) <= layer1_outputs(8625);
    layer2_outputs(5450) <= layer1_outputs(4059);
    layer2_outputs(5451) <= (layer1_outputs(5901)) or (layer1_outputs(345));
    layer2_outputs(5452) <= layer1_outputs(7686);
    layer2_outputs(5453) <= (layer1_outputs(668)) and (layer1_outputs(2183));
    layer2_outputs(5454) <= not(layer1_outputs(2067));
    layer2_outputs(5455) <= (layer1_outputs(6370)) or (layer1_outputs(3120));
    layer2_outputs(5456) <= not(layer1_outputs(3050));
    layer2_outputs(5457) <= layer1_outputs(7997);
    layer2_outputs(5458) <= not((layer1_outputs(9196)) and (layer1_outputs(4615)));
    layer2_outputs(5459) <= not(layer1_outputs(9218)) or (layer1_outputs(3091));
    layer2_outputs(5460) <= (layer1_outputs(1206)) and not (layer1_outputs(94));
    layer2_outputs(5461) <= not(layer1_outputs(4471)) or (layer1_outputs(1056));
    layer2_outputs(5462) <= '1';
    layer2_outputs(5463) <= not(layer1_outputs(9343));
    layer2_outputs(5464) <= (layer1_outputs(3236)) and not (layer1_outputs(2782));
    layer2_outputs(5465) <= not((layer1_outputs(9723)) or (layer1_outputs(5930)));
    layer2_outputs(5466) <= not(layer1_outputs(9265)) or (layer1_outputs(8149));
    layer2_outputs(5467) <= layer1_outputs(9457);
    layer2_outputs(5468) <= (layer1_outputs(9597)) xor (layer1_outputs(5747));
    layer2_outputs(5469) <= not(layer1_outputs(8022));
    layer2_outputs(5470) <= (layer1_outputs(7843)) and not (layer1_outputs(95));
    layer2_outputs(5471) <= (layer1_outputs(1695)) and (layer1_outputs(2986));
    layer2_outputs(5472) <= not(layer1_outputs(2339));
    layer2_outputs(5473) <= (layer1_outputs(7497)) or (layer1_outputs(3212));
    layer2_outputs(5474) <= (layer1_outputs(3309)) and (layer1_outputs(9046));
    layer2_outputs(5475) <= not(layer1_outputs(9004));
    layer2_outputs(5476) <= not((layer1_outputs(171)) xor (layer1_outputs(5456)));
    layer2_outputs(5477) <= (layer1_outputs(3198)) xor (layer1_outputs(4915));
    layer2_outputs(5478) <= not(layer1_outputs(1923));
    layer2_outputs(5479) <= not((layer1_outputs(2920)) xor (layer1_outputs(9780)));
    layer2_outputs(5480) <= not((layer1_outputs(1555)) and (layer1_outputs(784)));
    layer2_outputs(5481) <= '1';
    layer2_outputs(5482) <= layer1_outputs(7332);
    layer2_outputs(5483) <= '1';
    layer2_outputs(5484) <= (layer1_outputs(9724)) and not (layer1_outputs(1818));
    layer2_outputs(5485) <= '1';
    layer2_outputs(5486) <= not((layer1_outputs(8479)) and (layer1_outputs(2522)));
    layer2_outputs(5487) <= (layer1_outputs(7368)) or (layer1_outputs(6297));
    layer2_outputs(5488) <= not((layer1_outputs(8629)) or (layer1_outputs(7949)));
    layer2_outputs(5489) <= (layer1_outputs(4112)) and (layer1_outputs(9315));
    layer2_outputs(5490) <= not(layer1_outputs(5849));
    layer2_outputs(5491) <= layer1_outputs(4825);
    layer2_outputs(5492) <= not(layer1_outputs(8220)) or (layer1_outputs(7487));
    layer2_outputs(5493) <= not(layer1_outputs(1539)) or (layer1_outputs(515));
    layer2_outputs(5494) <= '0';
    layer2_outputs(5495) <= (layer1_outputs(5634)) and not (layer1_outputs(727));
    layer2_outputs(5496) <= (layer1_outputs(550)) and not (layer1_outputs(543));
    layer2_outputs(5497) <= not((layer1_outputs(10086)) and (layer1_outputs(4232)));
    layer2_outputs(5498) <= not(layer1_outputs(4571));
    layer2_outputs(5499) <= not(layer1_outputs(5220));
    layer2_outputs(5500) <= '1';
    layer2_outputs(5501) <= not((layer1_outputs(5334)) xor (layer1_outputs(1766)));
    layer2_outputs(5502) <= (layer1_outputs(8585)) and (layer1_outputs(5197));
    layer2_outputs(5503) <= layer1_outputs(2611);
    layer2_outputs(5504) <= not(layer1_outputs(9065));
    layer2_outputs(5505) <= not(layer1_outputs(7143));
    layer2_outputs(5506) <= layer1_outputs(5408);
    layer2_outputs(5507) <= (layer1_outputs(3831)) and not (layer1_outputs(7158));
    layer2_outputs(5508) <= (layer1_outputs(9059)) or (layer1_outputs(2114));
    layer2_outputs(5509) <= layer1_outputs(1204);
    layer2_outputs(5510) <= layer1_outputs(1183);
    layer2_outputs(5511) <= (layer1_outputs(3179)) xor (layer1_outputs(8290));
    layer2_outputs(5512) <= layer1_outputs(3803);
    layer2_outputs(5513) <= (layer1_outputs(7243)) and not (layer1_outputs(1656));
    layer2_outputs(5514) <= layer1_outputs(3691);
    layer2_outputs(5515) <= (layer1_outputs(5645)) or (layer1_outputs(202));
    layer2_outputs(5516) <= (layer1_outputs(2787)) and not (layer1_outputs(4447));
    layer2_outputs(5517) <= not((layer1_outputs(4798)) and (layer1_outputs(640)));
    layer2_outputs(5518) <= not(layer1_outputs(1657)) or (layer1_outputs(4900));
    layer2_outputs(5519) <= layer1_outputs(8628);
    layer2_outputs(5520) <= not(layer1_outputs(2141));
    layer2_outputs(5521) <= (layer1_outputs(4045)) and not (layer1_outputs(1057));
    layer2_outputs(5522) <= (layer1_outputs(8389)) or (layer1_outputs(7065));
    layer2_outputs(5523) <= not(layer1_outputs(1309));
    layer2_outputs(5524) <= layer1_outputs(5626);
    layer2_outputs(5525) <= not(layer1_outputs(3690)) or (layer1_outputs(8994));
    layer2_outputs(5526) <= layer1_outputs(9134);
    layer2_outputs(5527) <= not(layer1_outputs(9178));
    layer2_outputs(5528) <= '0';
    layer2_outputs(5529) <= not((layer1_outputs(513)) xor (layer1_outputs(2630)));
    layer2_outputs(5530) <= layer1_outputs(5689);
    layer2_outputs(5531) <= (layer1_outputs(8431)) xor (layer1_outputs(8012));
    layer2_outputs(5532) <= not(layer1_outputs(6995));
    layer2_outputs(5533) <= layer1_outputs(4786);
    layer2_outputs(5534) <= (layer1_outputs(5014)) and not (layer1_outputs(4751));
    layer2_outputs(5535) <= not(layer1_outputs(9659)) or (layer1_outputs(1011));
    layer2_outputs(5536) <= layer1_outputs(182);
    layer2_outputs(5537) <= (layer1_outputs(282)) and not (layer1_outputs(1730));
    layer2_outputs(5538) <= not(layer1_outputs(7710));
    layer2_outputs(5539) <= not(layer1_outputs(6254)) or (layer1_outputs(1406));
    layer2_outputs(5540) <= (layer1_outputs(10200)) and (layer1_outputs(5249));
    layer2_outputs(5541) <= not(layer1_outputs(2748)) or (layer1_outputs(8083));
    layer2_outputs(5542) <= not(layer1_outputs(1417));
    layer2_outputs(5543) <= not(layer1_outputs(9546));
    layer2_outputs(5544) <= layer1_outputs(9013);
    layer2_outputs(5545) <= layer1_outputs(7143);
    layer2_outputs(5546) <= layer1_outputs(4671);
    layer2_outputs(5547) <= not((layer1_outputs(6380)) and (layer1_outputs(1017)));
    layer2_outputs(5548) <= not(layer1_outputs(3347));
    layer2_outputs(5549) <= not(layer1_outputs(7274));
    layer2_outputs(5550) <= '0';
    layer2_outputs(5551) <= (layer1_outputs(2263)) and not (layer1_outputs(3088));
    layer2_outputs(5552) <= layer1_outputs(1545);
    layer2_outputs(5553) <= not(layer1_outputs(6338));
    layer2_outputs(5554) <= (layer1_outputs(9322)) and (layer1_outputs(4040));
    layer2_outputs(5555) <= '0';
    layer2_outputs(5556) <= not(layer1_outputs(10));
    layer2_outputs(5557) <= not(layer1_outputs(2330));
    layer2_outputs(5558) <= layer1_outputs(5248);
    layer2_outputs(5559) <= not((layer1_outputs(3189)) xor (layer1_outputs(7586)));
    layer2_outputs(5560) <= layer1_outputs(9542);
    layer2_outputs(5561) <= '1';
    layer2_outputs(5562) <= layer1_outputs(2368);
    layer2_outputs(5563) <= layer1_outputs(5539);
    layer2_outputs(5564) <= layer1_outputs(2117);
    layer2_outputs(5565) <= not((layer1_outputs(8075)) and (layer1_outputs(4666)));
    layer2_outputs(5566) <= not(layer1_outputs(4653)) or (layer1_outputs(6522));
    layer2_outputs(5567) <= layer1_outputs(556);
    layer2_outputs(5568) <= '0';
    layer2_outputs(5569) <= layer1_outputs(7467);
    layer2_outputs(5570) <= '1';
    layer2_outputs(5571) <= layer1_outputs(7533);
    layer2_outputs(5572) <= not(layer1_outputs(390));
    layer2_outputs(5573) <= layer1_outputs(8893);
    layer2_outputs(5574) <= (layer1_outputs(5848)) and (layer1_outputs(8747));
    layer2_outputs(5575) <= (layer1_outputs(8940)) and not (layer1_outputs(8263));
    layer2_outputs(5576) <= (layer1_outputs(9272)) and not (layer1_outputs(5189));
    layer2_outputs(5577) <= not(layer1_outputs(4088)) or (layer1_outputs(2412));
    layer2_outputs(5578) <= not(layer1_outputs(3479));
    layer2_outputs(5579) <= not((layer1_outputs(3515)) or (layer1_outputs(621)));
    layer2_outputs(5580) <= (layer1_outputs(1674)) and (layer1_outputs(1669));
    layer2_outputs(5581) <= (layer1_outputs(3238)) and (layer1_outputs(6944));
    layer2_outputs(5582) <= (layer1_outputs(8600)) xor (layer1_outputs(1522));
    layer2_outputs(5583) <= layer1_outputs(7068);
    layer2_outputs(5584) <= layer1_outputs(4948);
    layer2_outputs(5585) <= layer1_outputs(6103);
    layer2_outputs(5586) <= layer1_outputs(1100);
    layer2_outputs(5587) <= not(layer1_outputs(6911));
    layer2_outputs(5588) <= layer1_outputs(7846);
    layer2_outputs(5589) <= layer1_outputs(9939);
    layer2_outputs(5590) <= '0';
    layer2_outputs(5591) <= '1';
    layer2_outputs(5592) <= not(layer1_outputs(1130));
    layer2_outputs(5593) <= not((layer1_outputs(8066)) or (layer1_outputs(3791)));
    layer2_outputs(5594) <= layer1_outputs(9359);
    layer2_outputs(5595) <= layer1_outputs(8201);
    layer2_outputs(5596) <= '0';
    layer2_outputs(5597) <= not(layer1_outputs(1851));
    layer2_outputs(5598) <= not(layer1_outputs(9922));
    layer2_outputs(5599) <= layer1_outputs(7606);
    layer2_outputs(5600) <= not(layer1_outputs(1521));
    layer2_outputs(5601) <= layer1_outputs(6421);
    layer2_outputs(5602) <= layer1_outputs(463);
    layer2_outputs(5603) <= not(layer1_outputs(10117));
    layer2_outputs(5604) <= not(layer1_outputs(3566));
    layer2_outputs(5605) <= (layer1_outputs(3615)) and (layer1_outputs(10128));
    layer2_outputs(5606) <= not(layer1_outputs(1101)) or (layer1_outputs(10187));
    layer2_outputs(5607) <= (layer1_outputs(5306)) or (layer1_outputs(3239));
    layer2_outputs(5608) <= (layer1_outputs(7558)) xor (layer1_outputs(5032));
    layer2_outputs(5609) <= (layer1_outputs(7967)) and not (layer1_outputs(7873));
    layer2_outputs(5610) <= layer1_outputs(6026);
    layer2_outputs(5611) <= (layer1_outputs(8945)) xor (layer1_outputs(3335));
    layer2_outputs(5612) <= (layer1_outputs(261)) xor (layer1_outputs(5068));
    layer2_outputs(5613) <= not(layer1_outputs(5376));
    layer2_outputs(5614) <= not((layer1_outputs(5806)) or (layer1_outputs(3795)));
    layer2_outputs(5615) <= (layer1_outputs(5194)) xor (layer1_outputs(9506));
    layer2_outputs(5616) <= layer1_outputs(3432);
    layer2_outputs(5617) <= not(layer1_outputs(6965));
    layer2_outputs(5618) <= not((layer1_outputs(5030)) or (layer1_outputs(5323)));
    layer2_outputs(5619) <= not(layer1_outputs(8388)) or (layer1_outputs(1471));
    layer2_outputs(5620) <= not((layer1_outputs(6112)) or (layer1_outputs(5966)));
    layer2_outputs(5621) <= not(layer1_outputs(2712)) or (layer1_outputs(2820));
    layer2_outputs(5622) <= (layer1_outputs(3151)) and (layer1_outputs(6119));
    layer2_outputs(5623) <= (layer1_outputs(6950)) and not (layer1_outputs(2767));
    layer2_outputs(5624) <= layer1_outputs(1433);
    layer2_outputs(5625) <= layer1_outputs(1706);
    layer2_outputs(5626) <= not(layer1_outputs(10078));
    layer2_outputs(5627) <= not(layer1_outputs(4973));
    layer2_outputs(5628) <= (layer1_outputs(3785)) and not (layer1_outputs(5182));
    layer2_outputs(5629) <= (layer1_outputs(4000)) and not (layer1_outputs(4879));
    layer2_outputs(5630) <= not((layer1_outputs(4440)) and (layer1_outputs(3042)));
    layer2_outputs(5631) <= not(layer1_outputs(181));
    layer2_outputs(5632) <= not((layer1_outputs(9684)) and (layer1_outputs(6521)));
    layer2_outputs(5633) <= (layer1_outputs(3694)) and (layer1_outputs(6285));
    layer2_outputs(5634) <= (layer1_outputs(2992)) and (layer1_outputs(7661));
    layer2_outputs(5635) <= (layer1_outputs(7793)) and (layer1_outputs(7050));
    layer2_outputs(5636) <= not((layer1_outputs(9254)) and (layer1_outputs(5744)));
    layer2_outputs(5637) <= layer1_outputs(1477);
    layer2_outputs(5638) <= layer1_outputs(5718);
    layer2_outputs(5639) <= not(layer1_outputs(1839));
    layer2_outputs(5640) <= not((layer1_outputs(6565)) or (layer1_outputs(1394)));
    layer2_outputs(5641) <= not(layer1_outputs(2647)) or (layer1_outputs(5223));
    layer2_outputs(5642) <= not(layer1_outputs(7287)) or (layer1_outputs(6834));
    layer2_outputs(5643) <= layer1_outputs(3261);
    layer2_outputs(5644) <= not(layer1_outputs(4554));
    layer2_outputs(5645) <= not(layer1_outputs(2808)) or (layer1_outputs(7453));
    layer2_outputs(5646) <= not(layer1_outputs(8973));
    layer2_outputs(5647) <= not((layer1_outputs(8949)) and (layer1_outputs(6689)));
    layer2_outputs(5648) <= not(layer1_outputs(7757)) or (layer1_outputs(1755));
    layer2_outputs(5649) <= not(layer1_outputs(7304));
    layer2_outputs(5650) <= not(layer1_outputs(10169)) or (layer1_outputs(2257));
    layer2_outputs(5651) <= not((layer1_outputs(1333)) and (layer1_outputs(2268)));
    layer2_outputs(5652) <= (layer1_outputs(2449)) xor (layer1_outputs(1724));
    layer2_outputs(5653) <= not(layer1_outputs(190)) or (layer1_outputs(3023));
    layer2_outputs(5654) <= not(layer1_outputs(5509));
    layer2_outputs(5655) <= not(layer1_outputs(43)) or (layer1_outputs(7707));
    layer2_outputs(5656) <= '0';
    layer2_outputs(5657) <= '0';
    layer2_outputs(5658) <= layer1_outputs(3332);
    layer2_outputs(5659) <= layer1_outputs(8715);
    layer2_outputs(5660) <= layer1_outputs(9725);
    layer2_outputs(5661) <= (layer1_outputs(2547)) and not (layer1_outputs(4898));
    layer2_outputs(5662) <= not(layer1_outputs(2014)) or (layer1_outputs(3941));
    layer2_outputs(5663) <= (layer1_outputs(7933)) xor (layer1_outputs(6085));
    layer2_outputs(5664) <= not(layer1_outputs(9497));
    layer2_outputs(5665) <= not(layer1_outputs(1522));
    layer2_outputs(5666) <= (layer1_outputs(5639)) and (layer1_outputs(3543));
    layer2_outputs(5667) <= layer1_outputs(5671);
    layer2_outputs(5668) <= not(layer1_outputs(6902)) or (layer1_outputs(9860));
    layer2_outputs(5669) <= (layer1_outputs(2267)) or (layer1_outputs(8738));
    layer2_outputs(5670) <= not(layer1_outputs(4732));
    layer2_outputs(5671) <= not(layer1_outputs(8418)) or (layer1_outputs(3283));
    layer2_outputs(5672) <= layer1_outputs(7724);
    layer2_outputs(5673) <= not(layer1_outputs(936));
    layer2_outputs(5674) <= (layer1_outputs(3964)) and (layer1_outputs(1529));
    layer2_outputs(5675) <= (layer1_outputs(7733)) xor (layer1_outputs(9752));
    layer2_outputs(5676) <= layer1_outputs(7828);
    layer2_outputs(5677) <= (layer1_outputs(2692)) or (layer1_outputs(5649));
    layer2_outputs(5678) <= '1';
    layer2_outputs(5679) <= layer1_outputs(1173);
    layer2_outputs(5680) <= layer1_outputs(9936);
    layer2_outputs(5681) <= layer1_outputs(5666);
    layer2_outputs(5682) <= layer1_outputs(1742);
    layer2_outputs(5683) <= not(layer1_outputs(6720)) or (layer1_outputs(2116));
    layer2_outputs(5684) <= not((layer1_outputs(3973)) xor (layer1_outputs(5262)));
    layer2_outputs(5685) <= not(layer1_outputs(5621)) or (layer1_outputs(2817));
    layer2_outputs(5686) <= layer1_outputs(5471);
    layer2_outputs(5687) <= (layer1_outputs(2695)) or (layer1_outputs(6044));
    layer2_outputs(5688) <= (layer1_outputs(9510)) xor (layer1_outputs(8935));
    layer2_outputs(5689) <= layer1_outputs(8939);
    layer2_outputs(5690) <= (layer1_outputs(7759)) and not (layer1_outputs(2311));
    layer2_outputs(5691) <= (layer1_outputs(2350)) and not (layer1_outputs(3922));
    layer2_outputs(5692) <= not(layer1_outputs(9224));
    layer2_outputs(5693) <= layer1_outputs(31);
    layer2_outputs(5694) <= (layer1_outputs(10096)) and not (layer1_outputs(4105));
    layer2_outputs(5695) <= layer1_outputs(4851);
    layer2_outputs(5696) <= layer1_outputs(257);
    layer2_outputs(5697) <= not(layer1_outputs(6961));
    layer2_outputs(5698) <= layer1_outputs(10043);
    layer2_outputs(5699) <= not((layer1_outputs(9316)) xor (layer1_outputs(2809)));
    layer2_outputs(5700) <= layer1_outputs(7416);
    layer2_outputs(5701) <= not(layer1_outputs(4818)) or (layer1_outputs(3026));
    layer2_outputs(5702) <= (layer1_outputs(239)) and not (layer1_outputs(2083));
    layer2_outputs(5703) <= (layer1_outputs(8142)) or (layer1_outputs(7841));
    layer2_outputs(5704) <= layer1_outputs(1047);
    layer2_outputs(5705) <= (layer1_outputs(1754)) and not (layer1_outputs(2239));
    layer2_outputs(5706) <= not((layer1_outputs(7952)) xor (layer1_outputs(9622)));
    layer2_outputs(5707) <= not(layer1_outputs(7753)) or (layer1_outputs(7936));
    layer2_outputs(5708) <= (layer1_outputs(7940)) and not (layer1_outputs(7156));
    layer2_outputs(5709) <= not(layer1_outputs(954));
    layer2_outputs(5710) <= not(layer1_outputs(5968));
    layer2_outputs(5711) <= (layer1_outputs(4589)) and (layer1_outputs(3982));
    layer2_outputs(5712) <= not((layer1_outputs(2169)) or (layer1_outputs(480)));
    layer2_outputs(5713) <= layer1_outputs(2568);
    layer2_outputs(5714) <= (layer1_outputs(9723)) and (layer1_outputs(1643));
    layer2_outputs(5715) <= layer1_outputs(5454);
    layer2_outputs(5716) <= layer1_outputs(9463);
    layer2_outputs(5717) <= layer1_outputs(123);
    layer2_outputs(5718) <= not(layer1_outputs(1672)) or (layer1_outputs(216));
    layer2_outputs(5719) <= layer1_outputs(8555);
    layer2_outputs(5720) <= not((layer1_outputs(9742)) xor (layer1_outputs(9886)));
    layer2_outputs(5721) <= not((layer1_outputs(2709)) and (layer1_outputs(5383)));
    layer2_outputs(5722) <= not((layer1_outputs(850)) or (layer1_outputs(6714)));
    layer2_outputs(5723) <= layer1_outputs(7551);
    layer2_outputs(5724) <= not(layer1_outputs(4139));
    layer2_outputs(5725) <= not(layer1_outputs(2719));
    layer2_outputs(5726) <= layer1_outputs(3841);
    layer2_outputs(5727) <= layer1_outputs(8545);
    layer2_outputs(5728) <= layer1_outputs(1156);
    layer2_outputs(5729) <= (layer1_outputs(6456)) and (layer1_outputs(10080));
    layer2_outputs(5730) <= '1';
    layer2_outputs(5731) <= not(layer1_outputs(7540)) or (layer1_outputs(3475));
    layer2_outputs(5732) <= not(layer1_outputs(9642));
    layer2_outputs(5733) <= not((layer1_outputs(6859)) and (layer1_outputs(6154)));
    layer2_outputs(5734) <= (layer1_outputs(1133)) xor (layer1_outputs(7589));
    layer2_outputs(5735) <= not((layer1_outputs(5859)) or (layer1_outputs(391)));
    layer2_outputs(5736) <= not(layer1_outputs(8059)) or (layer1_outputs(505));
    layer2_outputs(5737) <= not(layer1_outputs(8914));
    layer2_outputs(5738) <= not((layer1_outputs(3659)) and (layer1_outputs(3673)));
    layer2_outputs(5739) <= (layer1_outputs(4426)) and (layer1_outputs(4433));
    layer2_outputs(5740) <= (layer1_outputs(411)) xor (layer1_outputs(2466));
    layer2_outputs(5741) <= not(layer1_outputs(9401)) or (layer1_outputs(266));
    layer2_outputs(5742) <= (layer1_outputs(7479)) or (layer1_outputs(9289));
    layer2_outputs(5743) <= not(layer1_outputs(7146));
    layer2_outputs(5744) <= '0';
    layer2_outputs(5745) <= not(layer1_outputs(9940)) or (layer1_outputs(5021));
    layer2_outputs(5746) <= not((layer1_outputs(1581)) xor (layer1_outputs(7074)));
    layer2_outputs(5747) <= (layer1_outputs(8321)) or (layer1_outputs(6061));
    layer2_outputs(5748) <= layer1_outputs(4578);
    layer2_outputs(5749) <= (layer1_outputs(522)) and not (layer1_outputs(6302));
    layer2_outputs(5750) <= not(layer1_outputs(1327));
    layer2_outputs(5751) <= not(layer1_outputs(10162));
    layer2_outputs(5752) <= not((layer1_outputs(4896)) or (layer1_outputs(2490)));
    layer2_outputs(5753) <= not(layer1_outputs(3123));
    layer2_outputs(5754) <= (layer1_outputs(6888)) or (layer1_outputs(3695));
    layer2_outputs(5755) <= not((layer1_outputs(7580)) and (layer1_outputs(6979)));
    layer2_outputs(5756) <= layer1_outputs(8699);
    layer2_outputs(5757) <= '1';
    layer2_outputs(5758) <= layer1_outputs(9495);
    layer2_outputs(5759) <= not(layer1_outputs(268)) or (layer1_outputs(9558));
    layer2_outputs(5760) <= (layer1_outputs(3136)) or (layer1_outputs(1718));
    layer2_outputs(5761) <= layer1_outputs(9356);
    layer2_outputs(5762) <= layer1_outputs(9721);
    layer2_outputs(5763) <= not(layer1_outputs(10212));
    layer2_outputs(5764) <= not(layer1_outputs(1991)) or (layer1_outputs(203));
    layer2_outputs(5765) <= not(layer1_outputs(7502)) or (layer1_outputs(6386));
    layer2_outputs(5766) <= not((layer1_outputs(1332)) or (layer1_outputs(4838)));
    layer2_outputs(5767) <= (layer1_outputs(7716)) and (layer1_outputs(10222));
    layer2_outputs(5768) <= (layer1_outputs(9830)) or (layer1_outputs(8180));
    layer2_outputs(5769) <= (layer1_outputs(2733)) and not (layer1_outputs(1712));
    layer2_outputs(5770) <= not(layer1_outputs(4608));
    layer2_outputs(5771) <= layer1_outputs(8988);
    layer2_outputs(5772) <= (layer1_outputs(9533)) xor (layer1_outputs(8871));
    layer2_outputs(5773) <= layer1_outputs(265);
    layer2_outputs(5774) <= (layer1_outputs(8463)) and (layer1_outputs(4917));
    layer2_outputs(5775) <= not(layer1_outputs(4804));
    layer2_outputs(5776) <= (layer1_outputs(4301)) and not (layer1_outputs(3646));
    layer2_outputs(5777) <= (layer1_outputs(6337)) and not (layer1_outputs(1275));
    layer2_outputs(5778) <= layer1_outputs(1495);
    layer2_outputs(5779) <= (layer1_outputs(690)) xor (layer1_outputs(1718));
    layer2_outputs(5780) <= (layer1_outputs(2792)) and (layer1_outputs(5725));
    layer2_outputs(5781) <= not(layer1_outputs(1960));
    layer2_outputs(5782) <= layer1_outputs(4680);
    layer2_outputs(5783) <= not(layer1_outputs(9559)) or (layer1_outputs(10227));
    layer2_outputs(5784) <= (layer1_outputs(7714)) and not (layer1_outputs(5898));
    layer2_outputs(5785) <= not(layer1_outputs(10033));
    layer2_outputs(5786) <= not(layer1_outputs(1090)) or (layer1_outputs(6874));
    layer2_outputs(5787) <= (layer1_outputs(7080)) and not (layer1_outputs(6024));
    layer2_outputs(5788) <= not(layer1_outputs(7117));
    layer2_outputs(5789) <= layer1_outputs(5370);
    layer2_outputs(5790) <= layer1_outputs(7023);
    layer2_outputs(5791) <= (layer1_outputs(432)) and not (layer1_outputs(4597));
    layer2_outputs(5792) <= layer1_outputs(2);
    layer2_outputs(5793) <= not((layer1_outputs(2293)) and (layer1_outputs(364)));
    layer2_outputs(5794) <= not(layer1_outputs(2877)) or (layer1_outputs(8004));
    layer2_outputs(5795) <= not((layer1_outputs(2741)) or (layer1_outputs(1872)));
    layer2_outputs(5796) <= '0';
    layer2_outputs(5797) <= not(layer1_outputs(7119));
    layer2_outputs(5798) <= not(layer1_outputs(1034));
    layer2_outputs(5799) <= '1';
    layer2_outputs(5800) <= not(layer1_outputs(4157));
    layer2_outputs(5801) <= '1';
    layer2_outputs(5802) <= not(layer1_outputs(8546));
    layer2_outputs(5803) <= not(layer1_outputs(716)) or (layer1_outputs(5527));
    layer2_outputs(5804) <= not(layer1_outputs(4470));
    layer2_outputs(5805) <= not(layer1_outputs(8179));
    layer2_outputs(5806) <= (layer1_outputs(9083)) or (layer1_outputs(814));
    layer2_outputs(5807) <= layer1_outputs(4761);
    layer2_outputs(5808) <= (layer1_outputs(7519)) or (layer1_outputs(5895));
    layer2_outputs(5809) <= layer1_outputs(1940);
    layer2_outputs(5810) <= (layer1_outputs(10169)) and not (layer1_outputs(666));
    layer2_outputs(5811) <= not(layer1_outputs(6392));
    layer2_outputs(5812) <= layer1_outputs(4520);
    layer2_outputs(5813) <= layer1_outputs(3277);
    layer2_outputs(5814) <= not(layer1_outputs(3631));
    layer2_outputs(5815) <= not(layer1_outputs(5606));
    layer2_outputs(5816) <= layer1_outputs(7632);
    layer2_outputs(5817) <= not(layer1_outputs(9725));
    layer2_outputs(5818) <= (layer1_outputs(8285)) or (layer1_outputs(7567));
    layer2_outputs(5819) <= layer1_outputs(189);
    layer2_outputs(5820) <= '1';
    layer2_outputs(5821) <= not(layer1_outputs(6025));
    layer2_outputs(5822) <= '1';
    layer2_outputs(5823) <= (layer1_outputs(6280)) and not (layer1_outputs(5053));
    layer2_outputs(5824) <= not(layer1_outputs(6283)) or (layer1_outputs(5844));
    layer2_outputs(5825) <= not((layer1_outputs(7658)) xor (layer1_outputs(3340)));
    layer2_outputs(5826) <= layer1_outputs(4039);
    layer2_outputs(5827) <= not(layer1_outputs(2159));
    layer2_outputs(5828) <= (layer1_outputs(5928)) or (layer1_outputs(10134));
    layer2_outputs(5829) <= not(layer1_outputs(9871));
    layer2_outputs(5830) <= not(layer1_outputs(4308));
    layer2_outputs(5831) <= not((layer1_outputs(7796)) xor (layer1_outputs(7424)));
    layer2_outputs(5832) <= layer1_outputs(7736);
    layer2_outputs(5833) <= (layer1_outputs(641)) and (layer1_outputs(4456));
    layer2_outputs(5834) <= not((layer1_outputs(9572)) or (layer1_outputs(6425)));
    layer2_outputs(5835) <= '0';
    layer2_outputs(5836) <= '1';
    layer2_outputs(5837) <= layer1_outputs(6606);
    layer2_outputs(5838) <= not((layer1_outputs(6257)) or (layer1_outputs(3141)));
    layer2_outputs(5839) <= '0';
    layer2_outputs(5840) <= not(layer1_outputs(1488)) or (layer1_outputs(6116));
    layer2_outputs(5841) <= layer1_outputs(909);
    layer2_outputs(5842) <= layer1_outputs(8816);
    layer2_outputs(5843) <= not(layer1_outputs(6208)) or (layer1_outputs(9369));
    layer2_outputs(5844) <= layer1_outputs(2443);
    layer2_outputs(5845) <= (layer1_outputs(8857)) and (layer1_outputs(5089));
    layer2_outputs(5846) <= (layer1_outputs(6989)) and (layer1_outputs(8433));
    layer2_outputs(5847) <= (layer1_outputs(5327)) and (layer1_outputs(1846));
    layer2_outputs(5848) <= layer1_outputs(10032);
    layer2_outputs(5849) <= layer1_outputs(381);
    layer2_outputs(5850) <= layer1_outputs(2871);
    layer2_outputs(5851) <= not((layer1_outputs(9616)) and (layer1_outputs(6587)));
    layer2_outputs(5852) <= (layer1_outputs(10171)) and (layer1_outputs(2972));
    layer2_outputs(5853) <= (layer1_outputs(8109)) and (layer1_outputs(2631));
    layer2_outputs(5854) <= not(layer1_outputs(9903)) or (layer1_outputs(8020));
    layer2_outputs(5855) <= layer1_outputs(4596);
    layer2_outputs(5856) <= '0';
    layer2_outputs(5857) <= not(layer1_outputs(657));
    layer2_outputs(5858) <= (layer1_outputs(2777)) or (layer1_outputs(8496));
    layer2_outputs(5859) <= not(layer1_outputs(7246));
    layer2_outputs(5860) <= not((layer1_outputs(5163)) and (layer1_outputs(4574)));
    layer2_outputs(5861) <= layer1_outputs(92);
    layer2_outputs(5862) <= (layer1_outputs(1635)) xor (layer1_outputs(3817));
    layer2_outputs(5863) <= (layer1_outputs(7043)) and not (layer1_outputs(7171));
    layer2_outputs(5864) <= layer1_outputs(9368);
    layer2_outputs(5865) <= not(layer1_outputs(6653));
    layer2_outputs(5866) <= layer1_outputs(6097);
    layer2_outputs(5867) <= not(layer1_outputs(6984));
    layer2_outputs(5868) <= (layer1_outputs(5224)) and (layer1_outputs(632));
    layer2_outputs(5869) <= not(layer1_outputs(8872)) or (layer1_outputs(6243));
    layer2_outputs(5870) <= (layer1_outputs(4372)) and (layer1_outputs(471));
    layer2_outputs(5871) <= not(layer1_outputs(3209));
    layer2_outputs(5872) <= not((layer1_outputs(607)) xor (layer1_outputs(6294)));
    layer2_outputs(5873) <= not((layer1_outputs(4529)) and (layer1_outputs(8975)));
    layer2_outputs(5874) <= not(layer1_outputs(8995));
    layer2_outputs(5875) <= layer1_outputs(8951);
    layer2_outputs(5876) <= not((layer1_outputs(8148)) or (layer1_outputs(9038)));
    layer2_outputs(5877) <= not((layer1_outputs(1959)) and (layer1_outputs(896)));
    layer2_outputs(5878) <= not((layer1_outputs(2163)) or (layer1_outputs(1367)));
    layer2_outputs(5879) <= (layer1_outputs(4518)) and (layer1_outputs(2960));
    layer2_outputs(5880) <= not((layer1_outputs(5005)) or (layer1_outputs(4115)));
    layer2_outputs(5881) <= (layer1_outputs(5595)) or (layer1_outputs(2641));
    layer2_outputs(5882) <= not((layer1_outputs(6518)) xor (layer1_outputs(8205)));
    layer2_outputs(5883) <= not(layer1_outputs(6769));
    layer2_outputs(5884) <= (layer1_outputs(4987)) and not (layer1_outputs(1064));
    layer2_outputs(5885) <= (layer1_outputs(1915)) and not (layer1_outputs(8027));
    layer2_outputs(5886) <= not((layer1_outputs(5276)) and (layer1_outputs(5792)));
    layer2_outputs(5887) <= (layer1_outputs(1931)) or (layer1_outputs(3638));
    layer2_outputs(5888) <= not(layer1_outputs(9580));
    layer2_outputs(5889) <= '1';
    layer2_outputs(5890) <= not(layer1_outputs(8890));
    layer2_outputs(5891) <= layer1_outputs(5124);
    layer2_outputs(5892) <= not(layer1_outputs(9216)) or (layer1_outputs(5598));
    layer2_outputs(5893) <= layer1_outputs(5334);
    layer2_outputs(5894) <= layer1_outputs(470);
    layer2_outputs(5895) <= (layer1_outputs(3426)) xor (layer1_outputs(450));
    layer2_outputs(5896) <= layer1_outputs(358);
    layer2_outputs(5897) <= layer1_outputs(8053);
    layer2_outputs(5898) <= layer1_outputs(3943);
    layer2_outputs(5899) <= '1';
    layer2_outputs(5900) <= not(layer1_outputs(3401)) or (layer1_outputs(5324));
    layer2_outputs(5901) <= not(layer1_outputs(9685));
    layer2_outputs(5902) <= not(layer1_outputs(1733)) or (layer1_outputs(9354));
    layer2_outputs(5903) <= not(layer1_outputs(7898));
    layer2_outputs(5904) <= (layer1_outputs(6590)) and (layer1_outputs(9665));
    layer2_outputs(5905) <= (layer1_outputs(4281)) and not (layer1_outputs(2777));
    layer2_outputs(5906) <= not((layer1_outputs(3778)) and (layer1_outputs(8632)));
    layer2_outputs(5907) <= not(layer1_outputs(7448));
    layer2_outputs(5908) <= not((layer1_outputs(3687)) xor (layer1_outputs(6613)));
    layer2_outputs(5909) <= layer1_outputs(3955);
    layer2_outputs(5910) <= '1';
    layer2_outputs(5911) <= layer1_outputs(1441);
    layer2_outputs(5912) <= '0';
    layer2_outputs(5913) <= (layer1_outputs(6021)) xor (layer1_outputs(2827));
    layer2_outputs(5914) <= layer1_outputs(6361);
    layer2_outputs(5915) <= layer1_outputs(191);
    layer2_outputs(5916) <= not(layer1_outputs(9128));
    layer2_outputs(5917) <= not(layer1_outputs(6410));
    layer2_outputs(5918) <= (layer1_outputs(7556)) and (layer1_outputs(7054));
    layer2_outputs(5919) <= '0';
    layer2_outputs(5920) <= not(layer1_outputs(7480));
    layer2_outputs(5921) <= not(layer1_outputs(9896));
    layer2_outputs(5922) <= not(layer1_outputs(6300));
    layer2_outputs(5923) <= layer1_outputs(3258);
    layer2_outputs(5924) <= (layer1_outputs(4620)) and not (layer1_outputs(8707));
    layer2_outputs(5925) <= layer1_outputs(4280);
    layer2_outputs(5926) <= not((layer1_outputs(1898)) xor (layer1_outputs(3346)));
    layer2_outputs(5927) <= (layer1_outputs(628)) or (layer1_outputs(1016));
    layer2_outputs(5928) <= (layer1_outputs(6563)) or (layer1_outputs(1299));
    layer2_outputs(5929) <= not((layer1_outputs(5546)) xor (layer1_outputs(6207)));
    layer2_outputs(5930) <= not(layer1_outputs(8737));
    layer2_outputs(5931) <= not((layer1_outputs(4352)) or (layer1_outputs(3091)));
    layer2_outputs(5932) <= layer1_outputs(6370);
    layer2_outputs(5933) <= (layer1_outputs(451)) and (layer1_outputs(3278));
    layer2_outputs(5934) <= '0';
    layer2_outputs(5935) <= layer1_outputs(9915);
    layer2_outputs(5936) <= layer1_outputs(4741);
    layer2_outputs(5937) <= (layer1_outputs(1340)) and (layer1_outputs(7702));
    layer2_outputs(5938) <= not(layer1_outputs(5266)) or (layer1_outputs(3780));
    layer2_outputs(5939) <= not(layer1_outputs(9298)) or (layer1_outputs(6575));
    layer2_outputs(5940) <= not(layer1_outputs(2615));
    layer2_outputs(5941) <= '0';
    layer2_outputs(5942) <= '1';
    layer2_outputs(5943) <= (layer1_outputs(4552)) and not (layer1_outputs(9485));
    layer2_outputs(5944) <= layer1_outputs(1697);
    layer2_outputs(5945) <= layer1_outputs(8892);
    layer2_outputs(5946) <= not((layer1_outputs(3049)) xor (layer1_outputs(7814)));
    layer2_outputs(5947) <= not(layer1_outputs(9802)) or (layer1_outputs(2553));
    layer2_outputs(5948) <= not((layer1_outputs(5555)) and (layer1_outputs(9753)));
    layer2_outputs(5949) <= layer1_outputs(10238);
    layer2_outputs(5950) <= not(layer1_outputs(7737)) or (layer1_outputs(3305));
    layer2_outputs(5951) <= '0';
    layer2_outputs(5952) <= (layer1_outputs(10073)) and not (layer1_outputs(4901));
    layer2_outputs(5953) <= (layer1_outputs(10101)) and (layer1_outputs(2963));
    layer2_outputs(5954) <= (layer1_outputs(7440)) and not (layer1_outputs(5131));
    layer2_outputs(5955) <= not(layer1_outputs(6364)) or (layer1_outputs(5675));
    layer2_outputs(5956) <= not((layer1_outputs(5489)) or (layer1_outputs(9515)));
    layer2_outputs(5957) <= not(layer1_outputs(1066));
    layer2_outputs(5958) <= layer1_outputs(2060);
    layer2_outputs(5959) <= (layer1_outputs(8282)) xor (layer1_outputs(2084));
    layer2_outputs(5960) <= layer1_outputs(359);
    layer2_outputs(5961) <= not(layer1_outputs(5175)) or (layer1_outputs(4303));
    layer2_outputs(5962) <= not(layer1_outputs(1285)) or (layer1_outputs(2140));
    layer2_outputs(5963) <= not((layer1_outputs(10221)) and (layer1_outputs(9011)));
    layer2_outputs(5964) <= layer1_outputs(2357);
    layer2_outputs(5965) <= not(layer1_outputs(4491)) or (layer1_outputs(8214));
    layer2_outputs(5966) <= not(layer1_outputs(477));
    layer2_outputs(5967) <= not(layer1_outputs(5078));
    layer2_outputs(5968) <= (layer1_outputs(6715)) and (layer1_outputs(3326));
    layer2_outputs(5969) <= not((layer1_outputs(1699)) and (layer1_outputs(7606)));
    layer2_outputs(5970) <= (layer1_outputs(8470)) xor (layer1_outputs(9893));
    layer2_outputs(5971) <= (layer1_outputs(6705)) and not (layer1_outputs(2971));
    layer2_outputs(5972) <= layer1_outputs(6303);
    layer2_outputs(5973) <= (layer1_outputs(2802)) xor (layer1_outputs(3078));
    layer2_outputs(5974) <= layer1_outputs(7480);
    layer2_outputs(5975) <= (layer1_outputs(2045)) and (layer1_outputs(8336));
    layer2_outputs(5976) <= not((layer1_outputs(6811)) and (layer1_outputs(39)));
    layer2_outputs(5977) <= '1';
    layer2_outputs(5978) <= not((layer1_outputs(1464)) xor (layer1_outputs(8465)));
    layer2_outputs(5979) <= '1';
    layer2_outputs(5980) <= not(layer1_outputs(7550)) or (layer1_outputs(3097));
    layer2_outputs(5981) <= layer1_outputs(4881);
    layer2_outputs(5982) <= not(layer1_outputs(8836));
    layer2_outputs(5983) <= not(layer1_outputs(1380));
    layer2_outputs(5984) <= not((layer1_outputs(6232)) or (layer1_outputs(6497)));
    layer2_outputs(5985) <= not(layer1_outputs(4409)) or (layer1_outputs(5253));
    layer2_outputs(5986) <= layer1_outputs(7291);
    layer2_outputs(5987) <= layer1_outputs(1781);
    layer2_outputs(5988) <= layer1_outputs(8134);
    layer2_outputs(5989) <= layer1_outputs(5054);
    layer2_outputs(5990) <= not(layer1_outputs(4068)) or (layer1_outputs(3080));
    layer2_outputs(5991) <= not((layer1_outputs(3671)) or (layer1_outputs(9641)));
    layer2_outputs(5992) <= not((layer1_outputs(2928)) or (layer1_outputs(9915)));
    layer2_outputs(5993) <= not(layer1_outputs(492));
    layer2_outputs(5994) <= not(layer1_outputs(6802));
    layer2_outputs(5995) <= not(layer1_outputs(1454));
    layer2_outputs(5996) <= (layer1_outputs(6844)) and not (layer1_outputs(125));
    layer2_outputs(5997) <= (layer1_outputs(6752)) and not (layer1_outputs(2290));
    layer2_outputs(5998) <= '0';
    layer2_outputs(5999) <= layer1_outputs(9177);
    layer2_outputs(6000) <= not((layer1_outputs(350)) xor (layer1_outputs(2942)));
    layer2_outputs(6001) <= not(layer1_outputs(6489));
    layer2_outputs(6002) <= (layer1_outputs(7569)) xor (layer1_outputs(7760));
    layer2_outputs(6003) <= (layer1_outputs(6426)) and not (layer1_outputs(1460));
    layer2_outputs(6004) <= not(layer1_outputs(8665));
    layer2_outputs(6005) <= not((layer1_outputs(1070)) or (layer1_outputs(3490)));
    layer2_outputs(6006) <= layer1_outputs(8274);
    layer2_outputs(6007) <= not(layer1_outputs(5955)) or (layer1_outputs(7839));
    layer2_outputs(6008) <= (layer1_outputs(7163)) and (layer1_outputs(3894));
    layer2_outputs(6009) <= (layer1_outputs(5955)) and (layer1_outputs(9867));
    layer2_outputs(6010) <= not((layer1_outputs(4261)) and (layer1_outputs(4607)));
    layer2_outputs(6011) <= not(layer1_outputs(9000));
    layer2_outputs(6012) <= layer1_outputs(2579);
    layer2_outputs(6013) <= (layer1_outputs(10151)) xor (layer1_outputs(6268));
    layer2_outputs(6014) <= not((layer1_outputs(7519)) and (layer1_outputs(8021)));
    layer2_outputs(6015) <= not((layer1_outputs(8622)) or (layer1_outputs(9604)));
    layer2_outputs(6016) <= not(layer1_outputs(5972)) or (layer1_outputs(4094));
    layer2_outputs(6017) <= not(layer1_outputs(561));
    layer2_outputs(6018) <= not(layer1_outputs(8266));
    layer2_outputs(6019) <= not(layer1_outputs(8853));
    layer2_outputs(6020) <= layer1_outputs(9515);
    layer2_outputs(6021) <= (layer1_outputs(4516)) and (layer1_outputs(5100));
    layer2_outputs(6022) <= '1';
    layer2_outputs(6023) <= (layer1_outputs(8195)) xor (layer1_outputs(9699));
    layer2_outputs(6024) <= (layer1_outputs(577)) or (layer1_outputs(4184));
    layer2_outputs(6025) <= layer1_outputs(4203);
    layer2_outputs(6026) <= layer1_outputs(3587);
    layer2_outputs(6027) <= '0';
    layer2_outputs(6028) <= not(layer1_outputs(6807)) or (layer1_outputs(8562));
    layer2_outputs(6029) <= not(layer1_outputs(3245)) or (layer1_outputs(3772));
    layer2_outputs(6030) <= not((layer1_outputs(2476)) and (layer1_outputs(7058)));
    layer2_outputs(6031) <= not(layer1_outputs(2765)) or (layer1_outputs(1000));
    layer2_outputs(6032) <= not(layer1_outputs(2955)) or (layer1_outputs(7280));
    layer2_outputs(6033) <= not(layer1_outputs(5985));
    layer2_outputs(6034) <= not((layer1_outputs(9498)) xor (layer1_outputs(4776)));
    layer2_outputs(6035) <= layer1_outputs(9366);
    layer2_outputs(6036) <= not(layer1_outputs(267));
    layer2_outputs(6037) <= layer1_outputs(9152);
    layer2_outputs(6038) <= layer1_outputs(6012);
    layer2_outputs(6039) <= layer1_outputs(6354);
    layer2_outputs(6040) <= (layer1_outputs(8339)) and not (layer1_outputs(640));
    layer2_outputs(6041) <= not(layer1_outputs(6905));
    layer2_outputs(6042) <= (layer1_outputs(3754)) and not (layer1_outputs(6306));
    layer2_outputs(6043) <= '0';
    layer2_outputs(6044) <= not((layer1_outputs(5302)) or (layer1_outputs(1061)));
    layer2_outputs(6045) <= (layer1_outputs(9460)) and not (layer1_outputs(10108));
    layer2_outputs(6046) <= (layer1_outputs(2980)) xor (layer1_outputs(2351));
    layer2_outputs(6047) <= '0';
    layer2_outputs(6048) <= (layer1_outputs(2291)) and not (layer1_outputs(7355));
    layer2_outputs(6049) <= not(layer1_outputs(6809)) or (layer1_outputs(2828));
    layer2_outputs(6050) <= (layer1_outputs(9384)) or (layer1_outputs(1262));
    layer2_outputs(6051) <= not((layer1_outputs(2217)) or (layer1_outputs(2943)));
    layer2_outputs(6052) <= not(layer1_outputs(4745));
    layer2_outputs(6053) <= (layer1_outputs(2048)) xor (layer1_outputs(4828));
    layer2_outputs(6054) <= layer1_outputs(4684);
    layer2_outputs(6055) <= layer1_outputs(3108);
    layer2_outputs(6056) <= not(layer1_outputs(3803));
    layer2_outputs(6057) <= (layer1_outputs(1312)) and not (layer1_outputs(4463));
    layer2_outputs(6058) <= (layer1_outputs(5422)) and (layer1_outputs(6115));
    layer2_outputs(6059) <= layer1_outputs(4824);
    layer2_outputs(6060) <= layer1_outputs(8085);
    layer2_outputs(6061) <= (layer1_outputs(846)) and not (layer1_outputs(9700));
    layer2_outputs(6062) <= not(layer1_outputs(5346));
    layer2_outputs(6063) <= (layer1_outputs(7187)) and not (layer1_outputs(5841));
    layer2_outputs(6064) <= not(layer1_outputs(5787));
    layer2_outputs(6065) <= layer1_outputs(6886);
    layer2_outputs(6066) <= (layer1_outputs(766)) or (layer1_outputs(4135));
    layer2_outputs(6067) <= not(layer1_outputs(2020));
    layer2_outputs(6068) <= (layer1_outputs(357)) or (layer1_outputs(5316));
    layer2_outputs(6069) <= layer1_outputs(5448);
    layer2_outputs(6070) <= not(layer1_outputs(2130)) or (layer1_outputs(3208));
    layer2_outputs(6071) <= '1';
    layer2_outputs(6072) <= layer1_outputs(3433);
    layer2_outputs(6073) <= (layer1_outputs(7868)) or (layer1_outputs(9387));
    layer2_outputs(6074) <= not(layer1_outputs(1312));
    layer2_outputs(6075) <= layer1_outputs(8923);
    layer2_outputs(6076) <= (layer1_outputs(5931)) and (layer1_outputs(3980));
    layer2_outputs(6077) <= not(layer1_outputs(9161)) or (layer1_outputs(6852));
    layer2_outputs(6078) <= (layer1_outputs(946)) xor (layer1_outputs(9661));
    layer2_outputs(6079) <= layer1_outputs(9031);
    layer2_outputs(6080) <= not((layer1_outputs(116)) and (layer1_outputs(7740)));
    layer2_outputs(6081) <= not((layer1_outputs(2011)) and (layer1_outputs(8413)));
    layer2_outputs(6082) <= not(layer1_outputs(7133));
    layer2_outputs(6083) <= (layer1_outputs(7786)) or (layer1_outputs(8415));
    layer2_outputs(6084) <= not(layer1_outputs(2415)) or (layer1_outputs(9894));
    layer2_outputs(6085) <= not(layer1_outputs(7378));
    layer2_outputs(6086) <= not((layer1_outputs(8594)) or (layer1_outputs(5450)));
    layer2_outputs(6087) <= not(layer1_outputs(2720)) or (layer1_outputs(9238));
    layer2_outputs(6088) <= '0';
    layer2_outputs(6089) <= not(layer1_outputs(2281));
    layer2_outputs(6090) <= not((layer1_outputs(1877)) and (layer1_outputs(9158)));
    layer2_outputs(6091) <= (layer1_outputs(3195)) and not (layer1_outputs(5665));
    layer2_outputs(6092) <= (layer1_outputs(9358)) and not (layer1_outputs(9800));
    layer2_outputs(6093) <= not(layer1_outputs(1738));
    layer2_outputs(6094) <= not((layer1_outputs(3009)) xor (layer1_outputs(7747)));
    layer2_outputs(6095) <= (layer1_outputs(7698)) or (layer1_outputs(6910));
    layer2_outputs(6096) <= '1';
    layer2_outputs(6097) <= not(layer1_outputs(6973)) or (layer1_outputs(7687));
    layer2_outputs(6098) <= not((layer1_outputs(8344)) or (layer1_outputs(9604)));
    layer2_outputs(6099) <= layer1_outputs(3584);
    layer2_outputs(6100) <= layer1_outputs(1598);
    layer2_outputs(6101) <= not(layer1_outputs(955));
    layer2_outputs(6102) <= not(layer1_outputs(3807));
    layer2_outputs(6103) <= layer1_outputs(1070);
    layer2_outputs(6104) <= layer1_outputs(1120);
    layer2_outputs(6105) <= not(layer1_outputs(3233));
    layer2_outputs(6106) <= (layer1_outputs(5094)) and not (layer1_outputs(7439));
    layer2_outputs(6107) <= not((layer1_outputs(10096)) or (layer1_outputs(4667)));
    layer2_outputs(6108) <= not(layer1_outputs(2203));
    layer2_outputs(6109) <= layer1_outputs(6715);
    layer2_outputs(6110) <= not(layer1_outputs(8383));
    layer2_outputs(6111) <= (layer1_outputs(3089)) and not (layer1_outputs(3067));
    layer2_outputs(6112) <= not((layer1_outputs(3562)) or (layer1_outputs(7009)));
    layer2_outputs(6113) <= not(layer1_outputs(6249)) or (layer1_outputs(7981));
    layer2_outputs(6114) <= layer1_outputs(9009);
    layer2_outputs(6115) <= not(layer1_outputs(3196));
    layer2_outputs(6116) <= not((layer1_outputs(6736)) xor (layer1_outputs(6888)));
    layer2_outputs(6117) <= (layer1_outputs(10143)) and not (layer1_outputs(3625));
    layer2_outputs(6118) <= not((layer1_outputs(1036)) xor (layer1_outputs(1058)));
    layer2_outputs(6119) <= not((layer1_outputs(3732)) xor (layer1_outputs(1264)));
    layer2_outputs(6120) <= layer1_outputs(6214);
    layer2_outputs(6121) <= not(layer1_outputs(7126)) or (layer1_outputs(5987));
    layer2_outputs(6122) <= (layer1_outputs(4547)) and not (layer1_outputs(584));
    layer2_outputs(6123) <= (layer1_outputs(4677)) and not (layer1_outputs(1777));
    layer2_outputs(6124) <= not(layer1_outputs(3455));
    layer2_outputs(6125) <= '0';
    layer2_outputs(6126) <= layer1_outputs(7234);
    layer2_outputs(6127) <= layer1_outputs(4897);
    layer2_outputs(6128) <= layer1_outputs(7440);
    layer2_outputs(6129) <= not(layer1_outputs(9422));
    layer2_outputs(6130) <= (layer1_outputs(504)) and (layer1_outputs(9019));
    layer2_outputs(6131) <= layer1_outputs(7291);
    layer2_outputs(6132) <= not(layer1_outputs(9228));
    layer2_outputs(6133) <= layer1_outputs(5420);
    layer2_outputs(6134) <= not((layer1_outputs(7423)) xor (layer1_outputs(6442)));
    layer2_outputs(6135) <= not(layer1_outputs(2322)) or (layer1_outputs(4334));
    layer2_outputs(6136) <= '1';
    layer2_outputs(6137) <= (layer1_outputs(7188)) and not (layer1_outputs(9574));
    layer2_outputs(6138) <= not((layer1_outputs(2037)) xor (layer1_outputs(8260)));
    layer2_outputs(6139) <= layer1_outputs(8015);
    layer2_outputs(6140) <= (layer1_outputs(4)) or (layer1_outputs(5));
    layer2_outputs(6141) <= not(layer1_outputs(731));
    layer2_outputs(6142) <= not((layer1_outputs(9076)) and (layer1_outputs(3724)));
    layer2_outputs(6143) <= not(layer1_outputs(6354));
    layer2_outputs(6144) <= not(layer1_outputs(5813));
    layer2_outputs(6145) <= layer1_outputs(1315);
    layer2_outputs(6146) <= (layer1_outputs(8410)) xor (layer1_outputs(3259));
    layer2_outputs(6147) <= (layer1_outputs(7792)) xor (layer1_outputs(417));
    layer2_outputs(6148) <= '1';
    layer2_outputs(6149) <= not((layer1_outputs(3027)) and (layer1_outputs(2040)));
    layer2_outputs(6150) <= layer1_outputs(6069);
    layer2_outputs(6151) <= (layer1_outputs(3636)) and not (layer1_outputs(3061));
    layer2_outputs(6152) <= not((layer1_outputs(4389)) or (layer1_outputs(1885)));
    layer2_outputs(6153) <= '1';
    layer2_outputs(6154) <= layer1_outputs(603);
    layer2_outputs(6155) <= layer1_outputs(5978);
    layer2_outputs(6156) <= (layer1_outputs(8874)) and not (layer1_outputs(5060));
    layer2_outputs(6157) <= (layer1_outputs(4435)) xor (layer1_outputs(3200));
    layer2_outputs(6158) <= '1';
    layer2_outputs(6159) <= not(layer1_outputs(9815));
    layer2_outputs(6160) <= not((layer1_outputs(8833)) xor (layer1_outputs(7911)));
    layer2_outputs(6161) <= (layer1_outputs(4104)) and not (layer1_outputs(2810));
    layer2_outputs(6162) <= (layer1_outputs(2001)) xor (layer1_outputs(3245));
    layer2_outputs(6163) <= layer1_outputs(1391);
    layer2_outputs(6164) <= not(layer1_outputs(9466));
    layer2_outputs(6165) <= not(layer1_outputs(3748));
    layer2_outputs(6166) <= '0';
    layer2_outputs(6167) <= (layer1_outputs(3590)) and not (layer1_outputs(5206));
    layer2_outputs(6168) <= layer1_outputs(10038);
    layer2_outputs(6169) <= layer1_outputs(10082);
    layer2_outputs(6170) <= layer1_outputs(6271);
    layer2_outputs(6171) <= '0';
    layer2_outputs(6172) <= layer1_outputs(1751);
    layer2_outputs(6173) <= not(layer1_outputs(8024));
    layer2_outputs(6174) <= not(layer1_outputs(1190)) or (layer1_outputs(1153));
    layer2_outputs(6175) <= not(layer1_outputs(8467));
    layer2_outputs(6176) <= layer1_outputs(7647);
    layer2_outputs(6177) <= (layer1_outputs(4117)) and (layer1_outputs(625));
    layer2_outputs(6178) <= not((layer1_outputs(2282)) or (layer1_outputs(7964)));
    layer2_outputs(6179) <= not(layer1_outputs(6576));
    layer2_outputs(6180) <= '0';
    layer2_outputs(6181) <= '0';
    layer2_outputs(6182) <= not(layer1_outputs(5940)) or (layer1_outputs(4717));
    layer2_outputs(6183) <= not(layer1_outputs(818));
    layer2_outputs(6184) <= layer1_outputs(9759);
    layer2_outputs(6185) <= (layer1_outputs(2784)) or (layer1_outputs(6916));
    layer2_outputs(6186) <= (layer1_outputs(3542)) xor (layer1_outputs(4657));
    layer2_outputs(6187) <= (layer1_outputs(8544)) and not (layer1_outputs(9478));
    layer2_outputs(6188) <= layer1_outputs(2801);
    layer2_outputs(6189) <= layer1_outputs(8303);
    layer2_outputs(6190) <= not((layer1_outputs(9445)) or (layer1_outputs(10140)));
    layer2_outputs(6191) <= not(layer1_outputs(3887));
    layer2_outputs(6192) <= (layer1_outputs(3081)) and not (layer1_outputs(5446));
    layer2_outputs(6193) <= (layer1_outputs(9930)) or (layer1_outputs(3938));
    layer2_outputs(6194) <= (layer1_outputs(4206)) and not (layer1_outputs(10112));
    layer2_outputs(6195) <= '1';
    layer2_outputs(6196) <= layer1_outputs(6362);
    layer2_outputs(6197) <= layer1_outputs(909);
    layer2_outputs(6198) <= not(layer1_outputs(3344));
    layer2_outputs(6199) <= not(layer1_outputs(2318));
    layer2_outputs(6200) <= not(layer1_outputs(6205)) or (layer1_outputs(7601));
    layer2_outputs(6201) <= not(layer1_outputs(9993)) or (layer1_outputs(1116));
    layer2_outputs(6202) <= '1';
    layer2_outputs(6203) <= not(layer1_outputs(10027));
    layer2_outputs(6204) <= layer1_outputs(2858);
    layer2_outputs(6205) <= not(layer1_outputs(5016));
    layer2_outputs(6206) <= layer1_outputs(9117);
    layer2_outputs(6207) <= not(layer1_outputs(5853)) or (layer1_outputs(8016));
    layer2_outputs(6208) <= (layer1_outputs(4689)) and not (layer1_outputs(8559));
    layer2_outputs(6209) <= (layer1_outputs(5133)) and (layer1_outputs(2328));
    layer2_outputs(6210) <= layer1_outputs(6978);
    layer2_outputs(6211) <= not((layer1_outputs(6222)) and (layer1_outputs(4172)));
    layer2_outputs(6212) <= not((layer1_outputs(5646)) xor (layer1_outputs(4479)));
    layer2_outputs(6213) <= (layer1_outputs(2242)) or (layer1_outputs(3288));
    layer2_outputs(6214) <= (layer1_outputs(5409)) and (layer1_outputs(5660));
    layer2_outputs(6215) <= not(layer1_outputs(205));
    layer2_outputs(6216) <= layer1_outputs(6241);
    layer2_outputs(6217) <= not(layer1_outputs(4785)) or (layer1_outputs(5122));
    layer2_outputs(6218) <= layer1_outputs(1811);
    layer2_outputs(6219) <= layer1_outputs(8079);
    layer2_outputs(6220) <= not(layer1_outputs(4539));
    layer2_outputs(6221) <= (layer1_outputs(8957)) and not (layer1_outputs(3688));
    layer2_outputs(6222) <= (layer1_outputs(9440)) and not (layer1_outputs(8495));
    layer2_outputs(6223) <= not((layer1_outputs(5169)) or (layer1_outputs(4470)));
    layer2_outputs(6224) <= not((layer1_outputs(9057)) xor (layer1_outputs(3319)));
    layer2_outputs(6225) <= layer1_outputs(4469);
    layer2_outputs(6226) <= not(layer1_outputs(3903));
    layer2_outputs(6227) <= '1';
    layer2_outputs(6228) <= (layer1_outputs(3508)) and not (layer1_outputs(7273));
    layer2_outputs(6229) <= '1';
    layer2_outputs(6230) <= not(layer1_outputs(3183));
    layer2_outputs(6231) <= layer1_outputs(5482);
    layer2_outputs(6232) <= layer1_outputs(652);
    layer2_outputs(6233) <= not(layer1_outputs(1174));
    layer2_outputs(6234) <= (layer1_outputs(3683)) and (layer1_outputs(9202));
    layer2_outputs(6235) <= not(layer1_outputs(7653)) or (layer1_outputs(1297));
    layer2_outputs(6236) <= not(layer1_outputs(6835));
    layer2_outputs(6237) <= not(layer1_outputs(4519));
    layer2_outputs(6238) <= layer1_outputs(4485);
    layer2_outputs(6239) <= not(layer1_outputs(9907));
    layer2_outputs(6240) <= not((layer1_outputs(7778)) and (layer1_outputs(2845)));
    layer2_outputs(6241) <= not(layer1_outputs(133)) or (layer1_outputs(8896));
    layer2_outputs(6242) <= (layer1_outputs(7543)) or (layer1_outputs(198));
    layer2_outputs(6243) <= '0';
    layer2_outputs(6244) <= not(layer1_outputs(8712));
    layer2_outputs(6245) <= not(layer1_outputs(7890));
    layer2_outputs(6246) <= layer1_outputs(1089);
    layer2_outputs(6247) <= not(layer1_outputs(9323));
    layer2_outputs(6248) <= (layer1_outputs(41)) and (layer1_outputs(4501));
    layer2_outputs(6249) <= '0';
    layer2_outputs(6250) <= not((layer1_outputs(9031)) or (layer1_outputs(3274)));
    layer2_outputs(6251) <= not(layer1_outputs(9875));
    layer2_outputs(6252) <= (layer1_outputs(2195)) or (layer1_outputs(7921));
    layer2_outputs(6253) <= not(layer1_outputs(6983));
    layer2_outputs(6254) <= (layer1_outputs(8729)) and not (layer1_outputs(5423));
    layer2_outputs(6255) <= not(layer1_outputs(9649));
    layer2_outputs(6256) <= (layer1_outputs(4527)) or (layer1_outputs(8120));
    layer2_outputs(6257) <= (layer1_outputs(5760)) and not (layer1_outputs(9113));
    layer2_outputs(6258) <= not(layer1_outputs(9123)) or (layer1_outputs(9316));
    layer2_outputs(6259) <= not(layer1_outputs(9379)) or (layer1_outputs(2864));
    layer2_outputs(6260) <= not(layer1_outputs(9611));
    layer2_outputs(6261) <= (layer1_outputs(421)) or (layer1_outputs(4187));
    layer2_outputs(6262) <= (layer1_outputs(3251)) and not (layer1_outputs(1847));
    layer2_outputs(6263) <= (layer1_outputs(8764)) xor (layer1_outputs(1914));
    layer2_outputs(6264) <= layer1_outputs(5155);
    layer2_outputs(6265) <= (layer1_outputs(2816)) or (layer1_outputs(1921));
    layer2_outputs(6266) <= (layer1_outputs(7446)) or (layer1_outputs(8236));
    layer2_outputs(6267) <= '0';
    layer2_outputs(6268) <= layer1_outputs(5838);
    layer2_outputs(6269) <= '1';
    layer2_outputs(6270) <= layer1_outputs(5354);
    layer2_outputs(6271) <= layer1_outputs(4551);
    layer2_outputs(6272) <= (layer1_outputs(1647)) or (layer1_outputs(7027));
    layer2_outputs(6273) <= layer1_outputs(7261);
    layer2_outputs(6274) <= layer1_outputs(2174);
    layer2_outputs(6275) <= not(layer1_outputs(5558));
    layer2_outputs(6276) <= layer1_outputs(297);
    layer2_outputs(6277) <= (layer1_outputs(4964)) or (layer1_outputs(3327));
    layer2_outputs(6278) <= layer1_outputs(3529);
    layer2_outputs(6279) <= (layer1_outputs(8916)) and (layer1_outputs(2687));
    layer2_outputs(6280) <= (layer1_outputs(7326)) xor (layer1_outputs(2014));
    layer2_outputs(6281) <= not(layer1_outputs(6724)) or (layer1_outputs(8762));
    layer2_outputs(6282) <= (layer1_outputs(4234)) and not (layer1_outputs(4365));
    layer2_outputs(6283) <= not(layer1_outputs(7638));
    layer2_outputs(6284) <= layer1_outputs(2473);
    layer2_outputs(6285) <= '0';
    layer2_outputs(6286) <= not(layer1_outputs(2233)) or (layer1_outputs(676));
    layer2_outputs(6287) <= not(layer1_outputs(7529));
    layer2_outputs(6288) <= layer1_outputs(7888);
    layer2_outputs(6289) <= not(layer1_outputs(4978));
    layer2_outputs(6290) <= not(layer1_outputs(3039));
    layer2_outputs(6291) <= not(layer1_outputs(6398)) or (layer1_outputs(924));
    layer2_outputs(6292) <= not(layer1_outputs(3848));
    layer2_outputs(6293) <= not(layer1_outputs(5512)) or (layer1_outputs(9791));
    layer2_outputs(6294) <= (layer1_outputs(7902)) xor (layer1_outputs(6533));
    layer2_outputs(6295) <= (layer1_outputs(241)) and not (layer1_outputs(8947));
    layer2_outputs(6296) <= (layer1_outputs(6246)) and not (layer1_outputs(1394));
    layer2_outputs(6297) <= layer1_outputs(9633);
    layer2_outputs(6298) <= (layer1_outputs(3941)) or (layer1_outputs(7572));
    layer2_outputs(6299) <= (layer1_outputs(263)) and not (layer1_outputs(5));
    layer2_outputs(6300) <= not(layer1_outputs(3613));
    layer2_outputs(6301) <= (layer1_outputs(3166)) and not (layer1_outputs(5378));
    layer2_outputs(6302) <= (layer1_outputs(3076)) and (layer1_outputs(2908));
    layer2_outputs(6303) <= (layer1_outputs(5211)) xor (layer1_outputs(4089));
    layer2_outputs(6304) <= not((layer1_outputs(8595)) or (layer1_outputs(1177)));
    layer2_outputs(6305) <= not(layer1_outputs(9120));
    layer2_outputs(6306) <= (layer1_outputs(8177)) and (layer1_outputs(1930));
    layer2_outputs(6307) <= not((layer1_outputs(3556)) xor (layer1_outputs(6148)));
    layer2_outputs(6308) <= not(layer1_outputs(8689));
    layer2_outputs(6309) <= (layer1_outputs(3448)) and not (layer1_outputs(6536));
    layer2_outputs(6310) <= not(layer1_outputs(9858));
    layer2_outputs(6311) <= not((layer1_outputs(8869)) xor (layer1_outputs(5265)));
    layer2_outputs(6312) <= (layer1_outputs(5821)) and not (layer1_outputs(4245));
    layer2_outputs(6313) <= '0';
    layer2_outputs(6314) <= not(layer1_outputs(10030));
    layer2_outputs(6315) <= not((layer1_outputs(2164)) xor (layer1_outputs(7582)));
    layer2_outputs(6316) <= not(layer1_outputs(9388)) or (layer1_outputs(8041));
    layer2_outputs(6317) <= layer1_outputs(10236);
    layer2_outputs(6318) <= not(layer1_outputs(9536)) or (layer1_outputs(5304));
    layer2_outputs(6319) <= not(layer1_outputs(685)) or (layer1_outputs(9803));
    layer2_outputs(6320) <= (layer1_outputs(5899)) and (layer1_outputs(6399));
    layer2_outputs(6321) <= '0';
    layer2_outputs(6322) <= (layer1_outputs(4119)) or (layer1_outputs(4038));
    layer2_outputs(6323) <= not(layer1_outputs(4124));
    layer2_outputs(6324) <= not(layer1_outputs(8823));
    layer2_outputs(6325) <= not((layer1_outputs(4080)) and (layer1_outputs(61)));
    layer2_outputs(6326) <= not((layer1_outputs(3360)) and (layer1_outputs(3368)));
    layer2_outputs(6327) <= not(layer1_outputs(7873));
    layer2_outputs(6328) <= not((layer1_outputs(6605)) and (layer1_outputs(8456)));
    layer2_outputs(6329) <= not(layer1_outputs(4591)) or (layer1_outputs(7947));
    layer2_outputs(6330) <= (layer1_outputs(1168)) or (layer1_outputs(4914));
    layer2_outputs(6331) <= not(layer1_outputs(624));
    layer2_outputs(6332) <= layer1_outputs(1421);
    layer2_outputs(6333) <= not((layer1_outputs(9952)) or (layer1_outputs(548)));
    layer2_outputs(6334) <= (layer1_outputs(6569)) xor (layer1_outputs(1242));
    layer2_outputs(6335) <= (layer1_outputs(1239)) and not (layer1_outputs(586));
    layer2_outputs(6336) <= layer1_outputs(1729);
    layer2_outputs(6337) <= not((layer1_outputs(4636)) or (layer1_outputs(3870)));
    layer2_outputs(6338) <= '1';
    layer2_outputs(6339) <= (layer1_outputs(9149)) and (layer1_outputs(5576));
    layer2_outputs(6340) <= not(layer1_outputs(7984));
    layer2_outputs(6341) <= not(layer1_outputs(446));
    layer2_outputs(6342) <= not(layer1_outputs(8954));
    layer2_outputs(6343) <= not(layer1_outputs(9814));
    layer2_outputs(6344) <= not(layer1_outputs(2829));
    layer2_outputs(6345) <= not((layer1_outputs(3229)) or (layer1_outputs(2307)));
    layer2_outputs(6346) <= layer1_outputs(1678);
    layer2_outputs(6347) <= not(layer1_outputs(879));
    layer2_outputs(6348) <= (layer1_outputs(8806)) and (layer1_outputs(7669));
    layer2_outputs(6349) <= '1';
    layer2_outputs(6350) <= '1';
    layer2_outputs(6351) <= not(layer1_outputs(7445));
    layer2_outputs(6352) <= not((layer1_outputs(4411)) and (layer1_outputs(5697)));
    layer2_outputs(6353) <= layer1_outputs(3784);
    layer2_outputs(6354) <= layer1_outputs(1466);
    layer2_outputs(6355) <= not((layer1_outputs(9385)) or (layer1_outputs(7201)));
    layer2_outputs(6356) <= '0';
    layer2_outputs(6357) <= not(layer1_outputs(9002));
    layer2_outputs(6358) <= layer1_outputs(5403);
    layer2_outputs(6359) <= not((layer1_outputs(7841)) and (layer1_outputs(6572)));
    layer2_outputs(6360) <= (layer1_outputs(4052)) and (layer1_outputs(2612));
    layer2_outputs(6361) <= layer1_outputs(232);
    layer2_outputs(6362) <= not((layer1_outputs(2969)) and (layer1_outputs(1838)));
    layer2_outputs(6363) <= (layer1_outputs(9990)) xor (layer1_outputs(9595));
    layer2_outputs(6364) <= layer1_outputs(8761);
    layer2_outputs(6365) <= layer1_outputs(4536);
    layer2_outputs(6366) <= not(layer1_outputs(1932));
    layer2_outputs(6367) <= not((layer1_outputs(2111)) and (layer1_outputs(5664)));
    layer2_outputs(6368) <= not(layer1_outputs(2169)) or (layer1_outputs(2562));
    layer2_outputs(6369) <= layer1_outputs(765);
    layer2_outputs(6370) <= layer1_outputs(3952);
    layer2_outputs(6371) <= not(layer1_outputs(4181)) or (layer1_outputs(9738));
    layer2_outputs(6372) <= not((layer1_outputs(5014)) or (layer1_outputs(7465)));
    layer2_outputs(6373) <= not(layer1_outputs(8908));
    layer2_outputs(6374) <= layer1_outputs(9477);
    layer2_outputs(6375) <= layer1_outputs(4551);
    layer2_outputs(6376) <= (layer1_outputs(9919)) and not (layer1_outputs(4319));
    layer2_outputs(6377) <= not(layer1_outputs(5486)) or (layer1_outputs(4370));
    layer2_outputs(6378) <= not(layer1_outputs(7398)) or (layer1_outputs(3726));
    layer2_outputs(6379) <= (layer1_outputs(806)) and not (layer1_outputs(5448));
    layer2_outputs(6380) <= (layer1_outputs(923)) and not (layer1_outputs(1621));
    layer2_outputs(6381) <= not(layer1_outputs(4194));
    layer2_outputs(6382) <= not((layer1_outputs(8633)) and (layer1_outputs(4638)));
    layer2_outputs(6383) <= not((layer1_outputs(4647)) xor (layer1_outputs(1118)));
    layer2_outputs(6384) <= not(layer1_outputs(9143));
    layer2_outputs(6385) <= not(layer1_outputs(578));
    layer2_outputs(6386) <= not(layer1_outputs(8241)) or (layer1_outputs(4316));
    layer2_outputs(6387) <= '0';
    layer2_outputs(6388) <= not((layer1_outputs(2556)) xor (layer1_outputs(6455)));
    layer2_outputs(6389) <= (layer1_outputs(7751)) and not (layer1_outputs(5076));
    layer2_outputs(6390) <= not(layer1_outputs(7762));
    layer2_outputs(6391) <= not((layer1_outputs(1122)) xor (layer1_outputs(3101)));
    layer2_outputs(6392) <= (layer1_outputs(4505)) and not (layer1_outputs(9693));
    layer2_outputs(6393) <= layer1_outputs(9251);
    layer2_outputs(6394) <= layer1_outputs(63);
    layer2_outputs(6395) <= (layer1_outputs(4271)) and not (layer1_outputs(9995));
    layer2_outputs(6396) <= (layer1_outputs(6591)) xor (layer1_outputs(7631));
    layer2_outputs(6397) <= (layer1_outputs(1556)) xor (layer1_outputs(3158));
    layer2_outputs(6398) <= layer1_outputs(1830);
    layer2_outputs(6399) <= layer1_outputs(1004);
    layer2_outputs(6400) <= not((layer1_outputs(8752)) or (layer1_outputs(2257)));
    layer2_outputs(6401) <= (layer1_outputs(5546)) and not (layer1_outputs(5062));
    layer2_outputs(6402) <= (layer1_outputs(8755)) and not (layer1_outputs(4860));
    layer2_outputs(6403) <= not(layer1_outputs(6987));
    layer2_outputs(6404) <= not(layer1_outputs(5210)) or (layer1_outputs(5545));
    layer2_outputs(6405) <= (layer1_outputs(7005)) and not (layer1_outputs(4819));
    layer2_outputs(6406) <= not((layer1_outputs(3600)) or (layer1_outputs(3853)));
    layer2_outputs(6407) <= (layer1_outputs(1022)) and not (layer1_outputs(9431));
    layer2_outputs(6408) <= '0';
    layer2_outputs(6409) <= not(layer1_outputs(9878));
    layer2_outputs(6410) <= (layer1_outputs(7692)) or (layer1_outputs(8773));
    layer2_outputs(6411) <= not((layer1_outputs(3368)) and (layer1_outputs(6261)));
    layer2_outputs(6412) <= not(layer1_outputs(1001));
    layer2_outputs(6413) <= not(layer1_outputs(7599));
    layer2_outputs(6414) <= '0';
    layer2_outputs(6415) <= not((layer1_outputs(661)) or (layer1_outputs(7011)));
    layer2_outputs(6416) <= not(layer1_outputs(1071));
    layer2_outputs(6417) <= layer1_outputs(407);
    layer2_outputs(6418) <= not(layer1_outputs(732));
    layer2_outputs(6419) <= layer1_outputs(956);
    layer2_outputs(6420) <= not((layer1_outputs(2956)) and (layer1_outputs(5384)));
    layer2_outputs(6421) <= (layer1_outputs(8565)) xor (layer1_outputs(6567));
    layer2_outputs(6422) <= not(layer1_outputs(7448));
    layer2_outputs(6423) <= (layer1_outputs(4994)) and (layer1_outputs(4894));
    layer2_outputs(6424) <= not(layer1_outputs(9225)) or (layer1_outputs(8688));
    layer2_outputs(6425) <= (layer1_outputs(5606)) and (layer1_outputs(5087));
    layer2_outputs(6426) <= (layer1_outputs(5849)) and (layer1_outputs(9648));
    layer2_outputs(6427) <= layer1_outputs(9895);
    layer2_outputs(6428) <= not((layer1_outputs(5861)) or (layer1_outputs(8435)));
    layer2_outputs(6429) <= '1';
    layer2_outputs(6430) <= not(layer1_outputs(1310));
    layer2_outputs(6431) <= layer1_outputs(6707);
    layer2_outputs(6432) <= layer1_outputs(8074);
    layer2_outputs(6433) <= (layer1_outputs(6327)) or (layer1_outputs(2941));
    layer2_outputs(6434) <= (layer1_outputs(4018)) and not (layer1_outputs(4610));
    layer2_outputs(6435) <= not(layer1_outputs(1548)) or (layer1_outputs(2905));
    layer2_outputs(6436) <= (layer1_outputs(8160)) and not (layer1_outputs(921));
    layer2_outputs(6437) <= '0';
    layer2_outputs(6438) <= not((layer1_outputs(240)) and (layer1_outputs(4883)));
    layer2_outputs(6439) <= layer1_outputs(1078);
    layer2_outputs(6440) <= not(layer1_outputs(6015));
    layer2_outputs(6441) <= layer1_outputs(9171);
    layer2_outputs(6442) <= not((layer1_outputs(1907)) xor (layer1_outputs(1902)));
    layer2_outputs(6443) <= '1';
    layer2_outputs(6444) <= not((layer1_outputs(9186)) xor (layer1_outputs(4114)));
    layer2_outputs(6445) <= not(layer1_outputs(6723));
    layer2_outputs(6446) <= '0';
    layer2_outputs(6447) <= not(layer1_outputs(769));
    layer2_outputs(6448) <= not(layer1_outputs(6738));
    layer2_outputs(6449) <= (layer1_outputs(6349)) and not (layer1_outputs(3481));
    layer2_outputs(6450) <= (layer1_outputs(3960)) or (layer1_outputs(440));
    layer2_outputs(6451) <= (layer1_outputs(4054)) and not (layer1_outputs(8278));
    layer2_outputs(6452) <= not(layer1_outputs(2809));
    layer2_outputs(6453) <= not((layer1_outputs(6339)) and (layer1_outputs(8682)));
    layer2_outputs(6454) <= not((layer1_outputs(8712)) xor (layer1_outputs(5600)));
    layer2_outputs(6455) <= not((layer1_outputs(9085)) or (layer1_outputs(7518)));
    layer2_outputs(6456) <= (layer1_outputs(8078)) and not (layer1_outputs(6798));
    layer2_outputs(6457) <= not((layer1_outputs(170)) and (layer1_outputs(2362)));
    layer2_outputs(6458) <= not(layer1_outputs(4694));
    layer2_outputs(6459) <= not(layer1_outputs(1603));
    layer2_outputs(6460) <= not((layer1_outputs(8031)) or (layer1_outputs(8973)));
    layer2_outputs(6461) <= layer1_outputs(4613);
    layer2_outputs(6462) <= layer1_outputs(7694);
    layer2_outputs(6463) <= not(layer1_outputs(198)) or (layer1_outputs(7446));
    layer2_outputs(6464) <= (layer1_outputs(1861)) or (layer1_outputs(4568));
    layer2_outputs(6465) <= not((layer1_outputs(1434)) or (layer1_outputs(2446)));
    layer2_outputs(6466) <= (layer1_outputs(6292)) and not (layer1_outputs(2337));
    layer2_outputs(6467) <= not(layer1_outputs(2762)) or (layer1_outputs(6552));
    layer2_outputs(6468) <= not(layer1_outputs(9337));
    layer2_outputs(6469) <= (layer1_outputs(7127)) and not (layer1_outputs(5473));
    layer2_outputs(6470) <= not(layer1_outputs(146));
    layer2_outputs(6471) <= not(layer1_outputs(4310));
    layer2_outputs(6472) <= (layer1_outputs(10209)) and not (layer1_outputs(8980));
    layer2_outputs(6473) <= (layer1_outputs(5775)) and (layer1_outputs(9345));
    layer2_outputs(6474) <= (layer1_outputs(7869)) or (layer1_outputs(8471));
    layer2_outputs(6475) <= not(layer1_outputs(9366));
    layer2_outputs(6476) <= (layer1_outputs(2206)) and not (layer1_outputs(606));
    layer2_outputs(6477) <= not(layer1_outputs(3175)) or (layer1_outputs(7453));
    layer2_outputs(6478) <= '0';
    layer2_outputs(6479) <= (layer1_outputs(556)) or (layer1_outputs(5110));
    layer2_outputs(6480) <= not(layer1_outputs(1795));
    layer2_outputs(6481) <= (layer1_outputs(1725)) and not (layer1_outputs(9783));
    layer2_outputs(6482) <= layer1_outputs(2454);
    layer2_outputs(6483) <= not((layer1_outputs(5566)) and (layer1_outputs(6745)));
    layer2_outputs(6484) <= (layer1_outputs(6650)) and not (layer1_outputs(2058));
    layer2_outputs(6485) <= layer1_outputs(834);
    layer2_outputs(6486) <= (layer1_outputs(6604)) and (layer1_outputs(938));
    layer2_outputs(6487) <= '0';
    layer2_outputs(6488) <= not(layer1_outputs(858));
    layer2_outputs(6489) <= not(layer1_outputs(7125)) or (layer1_outputs(329));
    layer2_outputs(6490) <= not((layer1_outputs(4200)) and (layer1_outputs(1764)));
    layer2_outputs(6491) <= (layer1_outputs(4740)) xor (layer1_outputs(1863));
    layer2_outputs(6492) <= not(layer1_outputs(1210));
    layer2_outputs(6493) <= not(layer1_outputs(496)) or (layer1_outputs(10206));
    layer2_outputs(6494) <= '0';
    layer2_outputs(6495) <= (layer1_outputs(6710)) xor (layer1_outputs(5305));
    layer2_outputs(6496) <= not(layer1_outputs(6368));
    layer2_outputs(6497) <= layer1_outputs(9096);
    layer2_outputs(6498) <= (layer1_outputs(7896)) and not (layer1_outputs(8895));
    layer2_outputs(6499) <= (layer1_outputs(9711)) or (layer1_outputs(3437));
    layer2_outputs(6500) <= (layer1_outputs(5333)) and not (layer1_outputs(6281));
    layer2_outputs(6501) <= layer1_outputs(7145);
    layer2_outputs(6502) <= layer1_outputs(2327);
    layer2_outputs(6503) <= (layer1_outputs(8159)) and not (layer1_outputs(304));
    layer2_outputs(6504) <= not(layer1_outputs(2861));
    layer2_outputs(6505) <= not(layer1_outputs(4211));
    layer2_outputs(6506) <= not(layer1_outputs(426));
    layer2_outputs(6507) <= layer1_outputs(5165);
    layer2_outputs(6508) <= '0';
    layer2_outputs(6509) <= not((layer1_outputs(2475)) or (layer1_outputs(112)));
    layer2_outputs(6510) <= layer1_outputs(5801);
    layer2_outputs(6511) <= (layer1_outputs(4093)) and not (layer1_outputs(2614));
    layer2_outputs(6512) <= not(layer1_outputs(7056));
    layer2_outputs(6513) <= not((layer1_outputs(9411)) or (layer1_outputs(5042)));
    layer2_outputs(6514) <= layer1_outputs(10070);
    layer2_outputs(6515) <= not((layer1_outputs(7939)) or (layer1_outputs(6882)));
    layer2_outputs(6516) <= not((layer1_outputs(7719)) or (layer1_outputs(5964)));
    layer2_outputs(6517) <= not(layer1_outputs(940));
    layer2_outputs(6518) <= (layer1_outputs(6711)) and not (layer1_outputs(8921));
    layer2_outputs(6519) <= (layer1_outputs(103)) and not (layer1_outputs(9945));
    layer2_outputs(6520) <= not(layer1_outputs(6759));
    layer2_outputs(6521) <= not(layer1_outputs(3408));
    layer2_outputs(6522) <= (layer1_outputs(5961)) and not (layer1_outputs(3627));
    layer2_outputs(6523) <= not(layer1_outputs(1249));
    layer2_outputs(6524) <= (layer1_outputs(1551)) and not (layer1_outputs(3114));
    layer2_outputs(6525) <= not((layer1_outputs(2200)) and (layer1_outputs(8286)));
    layer2_outputs(6526) <= layer1_outputs(4804);
    layer2_outputs(6527) <= not((layer1_outputs(7656)) xor (layer1_outputs(9616)));
    layer2_outputs(6528) <= not((layer1_outputs(4629)) and (layer1_outputs(1130)));
    layer2_outputs(6529) <= '1';
    layer2_outputs(6530) <= not(layer1_outputs(9022));
    layer2_outputs(6531) <= not(layer1_outputs(933)) or (layer1_outputs(6411));
    layer2_outputs(6532) <= layer1_outputs(6829);
    layer2_outputs(6533) <= (layer1_outputs(186)) and not (layer1_outputs(313));
    layer2_outputs(6534) <= layer1_outputs(252);
    layer2_outputs(6535) <= (layer1_outputs(7321)) and not (layer1_outputs(4272));
    layer2_outputs(6536) <= not(layer1_outputs(6350));
    layer2_outputs(6537) <= not(layer1_outputs(4021));
    layer2_outputs(6538) <= (layer1_outputs(3384)) and not (layer1_outputs(4289));
    layer2_outputs(6539) <= (layer1_outputs(3458)) or (layer1_outputs(9133));
    layer2_outputs(6540) <= (layer1_outputs(681)) and (layer1_outputs(23));
    layer2_outputs(6541) <= not((layer1_outputs(2310)) and (layer1_outputs(741)));
    layer2_outputs(6542) <= layer1_outputs(975);
    layer2_outputs(6543) <= not((layer1_outputs(8929)) or (layer1_outputs(5427)));
    layer2_outputs(6544) <= not((layer1_outputs(4537)) xor (layer1_outputs(8741)));
    layer2_outputs(6545) <= not(layer1_outputs(8293)) or (layer1_outputs(4331));
    layer2_outputs(6546) <= (layer1_outputs(9554)) and not (layer1_outputs(7509));
    layer2_outputs(6547) <= '0';
    layer2_outputs(6548) <= '1';
    layer2_outputs(6549) <= not(layer1_outputs(1900));
    layer2_outputs(6550) <= (layer1_outputs(1162)) or (layer1_outputs(7342));
    layer2_outputs(6551) <= (layer1_outputs(8750)) and (layer1_outputs(10189));
    layer2_outputs(6552) <= (layer1_outputs(8563)) and (layer1_outputs(7894));
    layer2_outputs(6553) <= not((layer1_outputs(7354)) and (layer1_outputs(1798)));
    layer2_outputs(6554) <= not(layer1_outputs(4199));
    layer2_outputs(6555) <= not((layer1_outputs(835)) and (layer1_outputs(1848)));
    layer2_outputs(6556) <= not((layer1_outputs(5868)) and (layer1_outputs(6209)));
    layer2_outputs(6557) <= not((layer1_outputs(6631)) and (layer1_outputs(9388)));
    layer2_outputs(6558) <= layer1_outputs(5653);
    layer2_outputs(6559) <= not((layer1_outputs(7373)) and (layer1_outputs(4009)));
    layer2_outputs(6560) <= layer1_outputs(3680);
    layer2_outputs(6561) <= layer1_outputs(6118);
    layer2_outputs(6562) <= not(layer1_outputs(4902)) or (layer1_outputs(934));
    layer2_outputs(6563) <= not((layer1_outputs(5783)) xor (layer1_outputs(9822)));
    layer2_outputs(6564) <= not(layer1_outputs(9602));
    layer2_outputs(6565) <= '0';
    layer2_outputs(6566) <= not(layer1_outputs(7748));
    layer2_outputs(6567) <= not((layer1_outputs(10014)) or (layer1_outputs(4812)));
    layer2_outputs(6568) <= not((layer1_outputs(2264)) or (layer1_outputs(2757)));
    layer2_outputs(6569) <= (layer1_outputs(1016)) or (layer1_outputs(876));
    layer2_outputs(6570) <= not(layer1_outputs(8258)) or (layer1_outputs(7924));
    layer2_outputs(6571) <= not((layer1_outputs(3999)) xor (layer1_outputs(3640)));
    layer2_outputs(6572) <= '1';
    layer2_outputs(6573) <= layer1_outputs(8999);
    layer2_outputs(6574) <= not(layer1_outputs(1704)) or (layer1_outputs(4612));
    layer2_outputs(6575) <= '1';
    layer2_outputs(6576) <= layer1_outputs(209);
    layer2_outputs(6577) <= not((layer1_outputs(7918)) or (layer1_outputs(9015)));
    layer2_outputs(6578) <= not(layer1_outputs(7464)) or (layer1_outputs(7693));
    layer2_outputs(6579) <= (layer1_outputs(8302)) and (layer1_outputs(144));
    layer2_outputs(6580) <= (layer1_outputs(8965)) xor (layer1_outputs(2245));
    layer2_outputs(6581) <= not(layer1_outputs(23)) or (layer1_outputs(3579));
    layer2_outputs(6582) <= not(layer1_outputs(9234));
    layer2_outputs(6583) <= (layer1_outputs(1217)) and not (layer1_outputs(2880));
    layer2_outputs(6584) <= (layer1_outputs(9214)) xor (layer1_outputs(9974));
    layer2_outputs(6585) <= not(layer1_outputs(6476));
    layer2_outputs(6586) <= not(layer1_outputs(7877)) or (layer1_outputs(1044));
    layer2_outputs(6587) <= (layer1_outputs(7160)) and not (layer1_outputs(3380));
    layer2_outputs(6588) <= layer1_outputs(9782);
    layer2_outputs(6589) <= (layer1_outputs(6818)) and not (layer1_outputs(8351));
    layer2_outputs(6590) <= '0';
    layer2_outputs(6591) <= layer1_outputs(1994);
    layer2_outputs(6592) <= not(layer1_outputs(4403));
    layer2_outputs(6593) <= not(layer1_outputs(5774));
    layer2_outputs(6594) <= not(layer1_outputs(2044));
    layer2_outputs(6595) <= (layer1_outputs(1235)) and (layer1_outputs(7011));
    layer2_outputs(6596) <= layer1_outputs(6868);
    layer2_outputs(6597) <= (layer1_outputs(1313)) and (layer1_outputs(3491));
    layer2_outputs(6598) <= (layer1_outputs(5840)) xor (layer1_outputs(3562));
    layer2_outputs(6599) <= not(layer1_outputs(5147));
    layer2_outputs(6600) <= layer1_outputs(8332);
    layer2_outputs(6601) <= layer1_outputs(1414);
    layer2_outputs(6602) <= not(layer1_outputs(4348));
    layer2_outputs(6603) <= not(layer1_outputs(9239)) or (layer1_outputs(1895));
    layer2_outputs(6604) <= layer1_outputs(8572);
    layer2_outputs(6605) <= layer1_outputs(316);
    layer2_outputs(6606) <= not(layer1_outputs(2700));
    layer2_outputs(6607) <= layer1_outputs(8836);
    layer2_outputs(6608) <= '1';
    layer2_outputs(6609) <= layer1_outputs(6107);
    layer2_outputs(6610) <= not(layer1_outputs(4938)) or (layer1_outputs(7742));
    layer2_outputs(6611) <= not(layer1_outputs(2831)) or (layer1_outputs(9989));
    layer2_outputs(6612) <= not(layer1_outputs(6144));
    layer2_outputs(6613) <= '1';
    layer2_outputs(6614) <= not(layer1_outputs(5786));
    layer2_outputs(6615) <= not(layer1_outputs(4217));
    layer2_outputs(6616) <= not((layer1_outputs(2941)) and (layer1_outputs(6823)));
    layer2_outputs(6617) <= (layer1_outputs(7852)) and not (layer1_outputs(5863));
    layer2_outputs(6618) <= (layer1_outputs(3620)) or (layer1_outputs(6344));
    layer2_outputs(6619) <= (layer1_outputs(6813)) and not (layer1_outputs(4518));
    layer2_outputs(6620) <= not((layer1_outputs(563)) or (layer1_outputs(2622)));
    layer2_outputs(6621) <= not((layer1_outputs(6644)) xor (layer1_outputs(8983)));
    layer2_outputs(6622) <= not(layer1_outputs(2036)) or (layer1_outputs(9976));
    layer2_outputs(6623) <= (layer1_outputs(7517)) and not (layer1_outputs(9395));
    layer2_outputs(6624) <= not(layer1_outputs(8052)) or (layer1_outputs(8596));
    layer2_outputs(6625) <= layer1_outputs(1325);
    layer2_outputs(6626) <= not(layer1_outputs(9110));
    layer2_outputs(6627) <= (layer1_outputs(8136)) xor (layer1_outputs(5685));
    layer2_outputs(6628) <= layer1_outputs(677);
    layer2_outputs(6629) <= (layer1_outputs(0)) or (layer1_outputs(8811));
    layer2_outputs(6630) <= not(layer1_outputs(9957));
    layer2_outputs(6631) <= not(layer1_outputs(3564));
    layer2_outputs(6632) <= not((layer1_outputs(961)) or (layer1_outputs(8905)));
    layer2_outputs(6633) <= not((layer1_outputs(1632)) or (layer1_outputs(8894)));
    layer2_outputs(6634) <= not((layer1_outputs(1208)) and (layer1_outputs(821)));
    layer2_outputs(6635) <= (layer1_outputs(1942)) and not (layer1_outputs(6299));
    layer2_outputs(6636) <= not(layer1_outputs(7106)) or (layer1_outputs(6308));
    layer2_outputs(6637) <= not((layer1_outputs(762)) and (layer1_outputs(241)));
    layer2_outputs(6638) <= (layer1_outputs(5960)) and not (layer1_outputs(1185));
    layer2_outputs(6639) <= layer1_outputs(9761);
    layer2_outputs(6640) <= '1';
    layer2_outputs(6641) <= layer1_outputs(7763);
    layer2_outputs(6642) <= not(layer1_outputs(2286));
    layer2_outputs(6643) <= not(layer1_outputs(419));
    layer2_outputs(6644) <= (layer1_outputs(1224)) and not (layer1_outputs(9235));
    layer2_outputs(6645) <= layer1_outputs(7366);
    layer2_outputs(6646) <= layer1_outputs(4266);
    layer2_outputs(6647) <= not((layer1_outputs(2646)) and (layer1_outputs(700)));
    layer2_outputs(6648) <= layer1_outputs(2677);
    layer2_outputs(6649) <= (layer1_outputs(3405)) xor (layer1_outputs(3713));
    layer2_outputs(6650) <= not(layer1_outputs(8199)) or (layer1_outputs(8722));
    layer2_outputs(6651) <= layer1_outputs(3106);
    layer2_outputs(6652) <= '1';
    layer2_outputs(6653) <= layer1_outputs(2624);
    layer2_outputs(6654) <= layer1_outputs(5891);
    layer2_outputs(6655) <= (layer1_outputs(8974)) and not (layer1_outputs(9143));
    layer2_outputs(6656) <= layer1_outputs(7212);
    layer2_outputs(6657) <= (layer1_outputs(2946)) and (layer1_outputs(9661));
    layer2_outputs(6658) <= (layer1_outputs(313)) or (layer1_outputs(1611));
    layer2_outputs(6659) <= not(layer1_outputs(2098)) or (layer1_outputs(4862));
    layer2_outputs(6660) <= '0';
    layer2_outputs(6661) <= not(layer1_outputs(7898));
    layer2_outputs(6662) <= not(layer1_outputs(1385));
    layer2_outputs(6663) <= layer1_outputs(4082);
    layer2_outputs(6664) <= not((layer1_outputs(2465)) or (layer1_outputs(1842)));
    layer2_outputs(6665) <= layer1_outputs(3855);
    layer2_outputs(6666) <= (layer1_outputs(4052)) and not (layer1_outputs(2692));
    layer2_outputs(6667) <= not(layer1_outputs(2573)) or (layer1_outputs(1452));
    layer2_outputs(6668) <= (layer1_outputs(3066)) and not (layer1_outputs(1638));
    layer2_outputs(6669) <= layer1_outputs(4703);
    layer2_outputs(6670) <= (layer1_outputs(1778)) and not (layer1_outputs(8830));
    layer2_outputs(6671) <= (layer1_outputs(4048)) and (layer1_outputs(6179));
    layer2_outputs(6672) <= layer1_outputs(6941);
    layer2_outputs(6673) <= not(layer1_outputs(9032)) or (layer1_outputs(1225));
    layer2_outputs(6674) <= (layer1_outputs(9309)) and not (layer1_outputs(7166));
    layer2_outputs(6675) <= not((layer1_outputs(3513)) or (layer1_outputs(9591)));
    layer2_outputs(6676) <= '0';
    layer2_outputs(6677) <= not(layer1_outputs(806));
    layer2_outputs(6678) <= not(layer1_outputs(1447));
    layer2_outputs(6679) <= (layer1_outputs(1593)) or (layer1_outputs(7100));
    layer2_outputs(6680) <= not((layer1_outputs(4785)) and (layer1_outputs(3532)));
    layer2_outputs(6681) <= (layer1_outputs(2075)) and (layer1_outputs(1742));
    layer2_outputs(6682) <= not(layer1_outputs(5002)) or (layer1_outputs(3143));
    layer2_outputs(6683) <= not(layer1_outputs(8281));
    layer2_outputs(6684) <= (layer1_outputs(2684)) and (layer1_outputs(10205));
    layer2_outputs(6685) <= '0';
    layer2_outputs(6686) <= not((layer1_outputs(4911)) xor (layer1_outputs(5288)));
    layer2_outputs(6687) <= not((layer1_outputs(4649)) and (layer1_outputs(2340)));
    layer2_outputs(6688) <= layer1_outputs(8824);
    layer2_outputs(6689) <= (layer1_outputs(4295)) and not (layer1_outputs(7002));
    layer2_outputs(6690) <= not((layer1_outputs(8463)) and (layer1_outputs(6608)));
    layer2_outputs(6691) <= not(layer1_outputs(9275)) or (layer1_outputs(5136));
    layer2_outputs(6692) <= layer1_outputs(2746);
    layer2_outputs(6693) <= not(layer1_outputs(7089)) or (layer1_outputs(9854));
    layer2_outputs(6694) <= (layer1_outputs(6479)) and (layer1_outputs(9321));
    layer2_outputs(6695) <= layer1_outputs(535);
    layer2_outputs(6696) <= not((layer1_outputs(4047)) xor (layer1_outputs(2100)));
    layer2_outputs(6697) <= (layer1_outputs(10146)) xor (layer1_outputs(6929));
    layer2_outputs(6698) <= (layer1_outputs(5521)) or (layer1_outputs(1654));
    layer2_outputs(6699) <= layer1_outputs(1754);
    layer2_outputs(6700) <= not(layer1_outputs(767));
    layer2_outputs(6701) <= not(layer1_outputs(177));
    layer2_outputs(6702) <= (layer1_outputs(637)) xor (layer1_outputs(9712));
    layer2_outputs(6703) <= (layer1_outputs(8440)) or (layer1_outputs(7822));
    layer2_outputs(6704) <= layer1_outputs(8266);
    layer2_outputs(6705) <= layer1_outputs(5264);
    layer2_outputs(6706) <= layer1_outputs(8454);
    layer2_outputs(6707) <= layer1_outputs(4212);
    layer2_outputs(6708) <= not(layer1_outputs(4178));
    layer2_outputs(6709) <= not((layer1_outputs(8315)) or (layer1_outputs(7157)));
    layer2_outputs(6710) <= layer1_outputs(9608);
    layer2_outputs(6711) <= (layer1_outputs(978)) xor (layer1_outputs(1791));
    layer2_outputs(6712) <= (layer1_outputs(7339)) and not (layer1_outputs(10237));
    layer2_outputs(6713) <= (layer1_outputs(7641)) and (layer1_outputs(3312));
    layer2_outputs(6714) <= not(layer1_outputs(6141));
    layer2_outputs(6715) <= not((layer1_outputs(7211)) and (layer1_outputs(827)));
    layer2_outputs(6716) <= '0';
    layer2_outputs(6717) <= not(layer1_outputs(6106)) or (layer1_outputs(4066));
    layer2_outputs(6718) <= not(layer1_outputs(7056));
    layer2_outputs(6719) <= layer1_outputs(2930);
    layer2_outputs(6720) <= (layer1_outputs(1195)) or (layer1_outputs(1676));
    layer2_outputs(6721) <= layer1_outputs(6785);
    layer2_outputs(6722) <= (layer1_outputs(2301)) and not (layer1_outputs(3490));
    layer2_outputs(6723) <= (layer1_outputs(7245)) or (layer1_outputs(3969));
    layer2_outputs(6724) <= not(layer1_outputs(3161)) or (layer1_outputs(3085));
    layer2_outputs(6725) <= not(layer1_outputs(1458)) or (layer1_outputs(181));
    layer2_outputs(6726) <= not((layer1_outputs(9414)) xor (layer1_outputs(9148)));
    layer2_outputs(6727) <= not(layer1_outputs(8323));
    layer2_outputs(6728) <= layer1_outputs(737);
    layer2_outputs(6729) <= not((layer1_outputs(3557)) and (layer1_outputs(259)));
    layer2_outputs(6730) <= layer1_outputs(1893);
    layer2_outputs(6731) <= not(layer1_outputs(1189));
    layer2_outputs(6732) <= not((layer1_outputs(5273)) or (layer1_outputs(8139)));
    layer2_outputs(6733) <= (layer1_outputs(8996)) and not (layer1_outputs(2093));
    layer2_outputs(6734) <= layer1_outputs(5239);
    layer2_outputs(6735) <= not(layer1_outputs(3130));
    layer2_outputs(6736) <= '1';
    layer2_outputs(6737) <= (layer1_outputs(6724)) and (layer1_outputs(126));
    layer2_outputs(6738) <= not(layer1_outputs(6424));
    layer2_outputs(6739) <= not(layer1_outputs(4787));
    layer2_outputs(6740) <= (layer1_outputs(9773)) xor (layer1_outputs(7766));
    layer2_outputs(6741) <= not(layer1_outputs(5923)) or (layer1_outputs(2236));
    layer2_outputs(6742) <= (layer1_outputs(9981)) and not (layer1_outputs(8007));
    layer2_outputs(6743) <= not((layer1_outputs(7357)) or (layer1_outputs(8172)));
    layer2_outputs(6744) <= (layer1_outputs(100)) and not (layer1_outputs(7959));
    layer2_outputs(6745) <= (layer1_outputs(8872)) and (layer1_outputs(10170));
    layer2_outputs(6746) <= not(layer1_outputs(1456));
    layer2_outputs(6747) <= not(layer1_outputs(3032));
    layer2_outputs(6748) <= not((layer1_outputs(8074)) or (layer1_outputs(8627)));
    layer2_outputs(6749) <= not((layer1_outputs(9900)) and (layer1_outputs(413)));
    layer2_outputs(6750) <= layer1_outputs(2824);
    layer2_outputs(6751) <= layer1_outputs(5699);
    layer2_outputs(6752) <= not(layer1_outputs(1935));
    layer2_outputs(6753) <= layer1_outputs(9625);
    layer2_outputs(6754) <= not((layer1_outputs(1143)) xor (layer1_outputs(7053)));
    layer2_outputs(6755) <= not((layer1_outputs(3505)) and (layer1_outputs(9710)));
    layer2_outputs(6756) <= (layer1_outputs(4932)) and (layer1_outputs(2145));
    layer2_outputs(6757) <= layer1_outputs(7523);
    layer2_outputs(6758) <= (layer1_outputs(3538)) and not (layer1_outputs(5775));
    layer2_outputs(6759) <= not(layer1_outputs(4058)) or (layer1_outputs(203));
    layer2_outputs(6760) <= layer1_outputs(4252);
    layer2_outputs(6761) <= not((layer1_outputs(1963)) and (layer1_outputs(3540)));
    layer2_outputs(6762) <= (layer1_outputs(705)) xor (layer1_outputs(4161));
    layer2_outputs(6763) <= (layer1_outputs(376)) and (layer1_outputs(6911));
    layer2_outputs(6764) <= not(layer1_outputs(8698));
    layer2_outputs(6765) <= not((layer1_outputs(6011)) xor (layer1_outputs(1258)));
    layer2_outputs(6766) <= not((layer1_outputs(2973)) or (layer1_outputs(4850)));
    layer2_outputs(6767) <= '1';
    layer2_outputs(6768) <= '0';
    layer2_outputs(6769) <= not(layer1_outputs(3146)) or (layer1_outputs(7460));
    layer2_outputs(6770) <= not(layer1_outputs(9353));
    layer2_outputs(6771) <= layer1_outputs(3835);
    layer2_outputs(6772) <= not((layer1_outputs(9856)) and (layer1_outputs(6734)));
    layer2_outputs(6773) <= (layer1_outputs(10160)) and not (layer1_outputs(1205));
    layer2_outputs(6774) <= not(layer1_outputs(10024));
    layer2_outputs(6775) <= not(layer1_outputs(8687)) or (layer1_outputs(4001));
    layer2_outputs(6776) <= (layer1_outputs(10038)) and not (layer1_outputs(4942));
    layer2_outputs(6777) <= not(layer1_outputs(4373));
    layer2_outputs(6778) <= (layer1_outputs(5538)) xor (layer1_outputs(8138));
    layer2_outputs(6779) <= not(layer1_outputs(1257));
    layer2_outputs(6780) <= layer1_outputs(6490);
    layer2_outputs(6781) <= not(layer1_outputs(2480)) or (layer1_outputs(5570));
    layer2_outputs(6782) <= not((layer1_outputs(4735)) xor (layer1_outputs(7964)));
    layer2_outputs(6783) <= layer1_outputs(1073);
    layer2_outputs(6784) <= not((layer1_outputs(9301)) xor (layer1_outputs(7859)));
    layer2_outputs(6785) <= not(layer1_outputs(6261));
    layer2_outputs(6786) <= not(layer1_outputs(8070));
    layer2_outputs(6787) <= not((layer1_outputs(2238)) xor (layer1_outputs(8881)));
    layer2_outputs(6788) <= (layer1_outputs(3453)) and not (layer1_outputs(3048));
    layer2_outputs(6789) <= (layer1_outputs(7359)) and not (layer1_outputs(3473));
    layer2_outputs(6790) <= '1';
    layer2_outputs(6791) <= not((layer1_outputs(1084)) and (layer1_outputs(167)));
    layer2_outputs(6792) <= not(layer1_outputs(4078)) or (layer1_outputs(8502));
    layer2_outputs(6793) <= not(layer1_outputs(2602)) or (layer1_outputs(2965));
    layer2_outputs(6794) <= not((layer1_outputs(3273)) or (layer1_outputs(9404)));
    layer2_outputs(6795) <= (layer1_outputs(6875)) and not (layer1_outputs(6832));
    layer2_outputs(6796) <= layer1_outputs(339);
    layer2_outputs(6797) <= layer1_outputs(7438);
    layer2_outputs(6798) <= layer1_outputs(4474);
    layer2_outputs(6799) <= (layer1_outputs(5607)) and not (layer1_outputs(5326));
    layer2_outputs(6800) <= '1';
    layer2_outputs(6801) <= (layer1_outputs(1185)) and not (layer1_outputs(1746));
    layer2_outputs(6802) <= '0';
    layer2_outputs(6803) <= not((layer1_outputs(2180)) xor (layer1_outputs(2892)));
    layer2_outputs(6804) <= not((layer1_outputs(8798)) xor (layer1_outputs(6180)));
    layer2_outputs(6805) <= (layer1_outputs(6535)) and not (layer1_outputs(8791));
    layer2_outputs(6806) <= '1';
    layer2_outputs(6807) <= layer1_outputs(8921);
    layer2_outputs(6808) <= not(layer1_outputs(8750)) or (layer1_outputs(3182));
    layer2_outputs(6809) <= (layer1_outputs(8627)) and not (layer1_outputs(4696));
    layer2_outputs(6810) <= '1';
    layer2_outputs(6811) <= (layer1_outputs(5419)) xor (layer1_outputs(4068));
    layer2_outputs(6812) <= layer1_outputs(5573);
    layer2_outputs(6813) <= not(layer1_outputs(8821)) or (layer1_outputs(7244));
    layer2_outputs(6814) <= (layer1_outputs(8670)) or (layer1_outputs(3519));
    layer2_outputs(6815) <= layer1_outputs(7152);
    layer2_outputs(6816) <= not(layer1_outputs(230));
    layer2_outputs(6817) <= not(layer1_outputs(6639)) or (layer1_outputs(2530));
    layer2_outputs(6818) <= not(layer1_outputs(2155));
    layer2_outputs(6819) <= not((layer1_outputs(4173)) and (layer1_outputs(770)));
    layer2_outputs(6820) <= (layer1_outputs(6759)) xor (layer1_outputs(723));
    layer2_outputs(6821) <= not(layer1_outputs(3069)) or (layer1_outputs(4246));
    layer2_outputs(6822) <= (layer1_outputs(8572)) or (layer1_outputs(5460));
    layer2_outputs(6823) <= (layer1_outputs(701)) or (layer1_outputs(7929));
    layer2_outputs(6824) <= not((layer1_outputs(2712)) and (layer1_outputs(7207)));
    layer2_outputs(6825) <= (layer1_outputs(7149)) or (layer1_outputs(8564));
    layer2_outputs(6826) <= (layer1_outputs(8777)) or (layer1_outputs(2600));
    layer2_outputs(6827) <= not((layer1_outputs(7385)) or (layer1_outputs(7675)));
    layer2_outputs(6828) <= '0';
    layer2_outputs(6829) <= not((layer1_outputs(5385)) and (layer1_outputs(5973)));
    layer2_outputs(6830) <= layer1_outputs(6581);
    layer2_outputs(6831) <= not(layer1_outputs(8427)) or (layer1_outputs(9102));
    layer2_outputs(6832) <= not((layer1_outputs(8460)) xor (layer1_outputs(9171)));
    layer2_outputs(6833) <= not(layer1_outputs(3760));
    layer2_outputs(6834) <= '0';
    layer2_outputs(6835) <= not((layer1_outputs(10115)) or (layer1_outputs(6884)));
    layer2_outputs(6836) <= not((layer1_outputs(1585)) or (layer1_outputs(2294)));
    layer2_outputs(6837) <= not(layer1_outputs(6398)) or (layer1_outputs(10227));
    layer2_outputs(6838) <= not(layer1_outputs(4242));
    layer2_outputs(6839) <= (layer1_outputs(3013)) or (layer1_outputs(9767));
    layer2_outputs(6840) <= '1';
    layer2_outputs(6841) <= (layer1_outputs(3034)) and not (layer1_outputs(803));
    layer2_outputs(6842) <= '0';
    layer2_outputs(6843) <= not((layer1_outputs(6278)) xor (layer1_outputs(196)));
    layer2_outputs(6844) <= not(layer1_outputs(2509)) or (layer1_outputs(8005));
    layer2_outputs(6845) <= layer1_outputs(8935);
    layer2_outputs(6846) <= (layer1_outputs(5404)) and not (layer1_outputs(2574));
    layer2_outputs(6847) <= not(layer1_outputs(6337));
    layer2_outputs(6848) <= layer1_outputs(7681);
    layer2_outputs(6849) <= layer1_outputs(392);
    layer2_outputs(6850) <= (layer1_outputs(6173)) and (layer1_outputs(5683));
    layer2_outputs(6851) <= (layer1_outputs(3426)) and not (layer1_outputs(8669));
    layer2_outputs(6852) <= (layer1_outputs(7169)) or (layer1_outputs(802));
    layer2_outputs(6853) <= not((layer1_outputs(2560)) and (layer1_outputs(1081)));
    layer2_outputs(6854) <= not(layer1_outputs(464));
    layer2_outputs(6855) <= not(layer1_outputs(7375));
    layer2_outputs(6856) <= (layer1_outputs(2555)) and not (layer1_outputs(3689));
    layer2_outputs(6857) <= (layer1_outputs(8045)) and not (layer1_outputs(3201));
    layer2_outputs(6858) <= layer1_outputs(80);
    layer2_outputs(6859) <= not(layer1_outputs(4817));
    layer2_outputs(6860) <= not(layer1_outputs(9571));
    layer2_outputs(6861) <= not(layer1_outputs(1977));
    layer2_outputs(6862) <= not(layer1_outputs(3790));
    layer2_outputs(6863) <= not((layer1_outputs(2016)) xor (layer1_outputs(4355)));
    layer2_outputs(6864) <= not((layer1_outputs(7854)) or (layer1_outputs(1197)));
    layer2_outputs(6865) <= not(layer1_outputs(5850));
    layer2_outputs(6866) <= not(layer1_outputs(9247));
    layer2_outputs(6867) <= not((layer1_outputs(4290)) and (layer1_outputs(1190)));
    layer2_outputs(6868) <= not(layer1_outputs(9130));
    layer2_outputs(6869) <= not(layer1_outputs(1163)) or (layer1_outputs(945));
    layer2_outputs(6870) <= (layer1_outputs(9152)) or (layer1_outputs(8172));
    layer2_outputs(6871) <= not(layer1_outputs(4791));
    layer2_outputs(6872) <= not(layer1_outputs(3477)) or (layer1_outputs(3270));
    layer2_outputs(6873) <= (layer1_outputs(2127)) xor (layer1_outputs(819));
    layer2_outputs(6874) <= (layer1_outputs(7260)) and not (layer1_outputs(9277));
    layer2_outputs(6875) <= not((layer1_outputs(7579)) xor (layer1_outputs(1449)));
    layer2_outputs(6876) <= (layer1_outputs(8740)) and not (layer1_outputs(8938));
    layer2_outputs(6877) <= (layer1_outputs(1123)) and (layer1_outputs(6676));
    layer2_outputs(6878) <= (layer1_outputs(1431)) xor (layer1_outputs(429));
    layer2_outputs(6879) <= layer1_outputs(3303);
    layer2_outputs(6880) <= (layer1_outputs(7388)) or (layer1_outputs(923));
    layer2_outputs(6881) <= not(layer1_outputs(3757)) or (layer1_outputs(2325));
    layer2_outputs(6882) <= not((layer1_outputs(5556)) xor (layer1_outputs(5234)));
    layer2_outputs(6883) <= layer1_outputs(7648);
    layer2_outputs(6884) <= layer1_outputs(5098);
    layer2_outputs(6885) <= layer1_outputs(9255);
    layer2_outputs(6886) <= not(layer1_outputs(544));
    layer2_outputs(6887) <= (layer1_outputs(4417)) xor (layer1_outputs(6171));
    layer2_outputs(6888) <= layer1_outputs(9583);
    layer2_outputs(6889) <= not(layer1_outputs(2107)) or (layer1_outputs(6667));
    layer2_outputs(6890) <= layer1_outputs(5455);
    layer2_outputs(6891) <= not(layer1_outputs(3606));
    layer2_outputs(6892) <= layer1_outputs(8430);
    layer2_outputs(6893) <= (layer1_outputs(3421)) and (layer1_outputs(3328));
    layer2_outputs(6894) <= (layer1_outputs(3770)) xor (layer1_outputs(9921));
    layer2_outputs(6895) <= (layer1_outputs(3567)) and (layer1_outputs(3079));
    layer2_outputs(6896) <= layer1_outputs(8411);
    layer2_outputs(6897) <= layer1_outputs(7797);
    layer2_outputs(6898) <= (layer1_outputs(7218)) xor (layer1_outputs(5229));
    layer2_outputs(6899) <= layer1_outputs(1230);
    layer2_outputs(6900) <= not(layer1_outputs(2022));
    layer2_outputs(6901) <= not((layer1_outputs(5215)) xor (layer1_outputs(8419)));
    layer2_outputs(6902) <= not(layer1_outputs(7100));
    layer2_outputs(6903) <= not(layer1_outputs(1214));
    layer2_outputs(6904) <= (layer1_outputs(1532)) and not (layer1_outputs(5096));
    layer2_outputs(6905) <= (layer1_outputs(3527)) or (layer1_outputs(5682));
    layer2_outputs(6906) <= not((layer1_outputs(8649)) or (layer1_outputs(7559)));
    layer2_outputs(6907) <= '1';
    layer2_outputs(6908) <= (layer1_outputs(1)) or (layer1_outputs(8703));
    layer2_outputs(6909) <= not(layer1_outputs(3030));
    layer2_outputs(6910) <= not(layer1_outputs(5694));
    layer2_outputs(6911) <= not(layer1_outputs(2954)) or (layer1_outputs(4591));
    layer2_outputs(6912) <= (layer1_outputs(8755)) and (layer1_outputs(5376));
    layer2_outputs(6913) <= not(layer1_outputs(6467));
    layer2_outputs(6914) <= layer1_outputs(3187);
    layer2_outputs(6915) <= layer1_outputs(1404);
    layer2_outputs(6916) <= (layer1_outputs(2433)) and not (layer1_outputs(3605));
    layer2_outputs(6917) <= not(layer1_outputs(5415));
    layer2_outputs(6918) <= not(layer1_outputs(5191)) or (layer1_outputs(2962));
    layer2_outputs(6919) <= '0';
    layer2_outputs(6920) <= not(layer1_outputs(4086)) or (layer1_outputs(4563));
    layer2_outputs(6921) <= not(layer1_outputs(9471));
    layer2_outputs(6922) <= not(layer1_outputs(8543)) or (layer1_outputs(605));
    layer2_outputs(6923) <= (layer1_outputs(1510)) and not (layer1_outputs(6402));
    layer2_outputs(6924) <= (layer1_outputs(5390)) and (layer1_outputs(708));
    layer2_outputs(6925) <= layer1_outputs(8999);
    layer2_outputs(6926) <= (layer1_outputs(3038)) and not (layer1_outputs(5139));
    layer2_outputs(6927) <= not(layer1_outputs(2434)) or (layer1_outputs(9274));
    layer2_outputs(6928) <= (layer1_outputs(5904)) and not (layer1_outputs(1864));
    layer2_outputs(6929) <= not(layer1_outputs(8003)) or (layer1_outputs(2504));
    layer2_outputs(6930) <= not(layer1_outputs(10056)) or (layer1_outputs(3787));
    layer2_outputs(6931) <= not(layer1_outputs(1614));
    layer2_outputs(6932) <= not(layer1_outputs(476));
    layer2_outputs(6933) <= not(layer1_outputs(2677));
    layer2_outputs(6934) <= not(layer1_outputs(6141));
    layer2_outputs(6935) <= layer1_outputs(6939);
    layer2_outputs(6936) <= not((layer1_outputs(7544)) or (layer1_outputs(4029)));
    layer2_outputs(6937) <= layer1_outputs(6063);
    layer2_outputs(6938) <= not((layer1_outputs(3653)) and (layer1_outputs(1893)));
    layer2_outputs(6939) <= not(layer1_outputs(5802));
    layer2_outputs(6940) <= not(layer1_outputs(10200));
    layer2_outputs(6941) <= not(layer1_outputs(5504)) or (layer1_outputs(9286));
    layer2_outputs(6942) <= layer1_outputs(8782);
    layer2_outputs(6943) <= not((layer1_outputs(6341)) and (layer1_outputs(4122)));
    layer2_outputs(6944) <= layer1_outputs(3418);
    layer2_outputs(6945) <= (layer1_outputs(7719)) and not (layer1_outputs(9908));
    layer2_outputs(6946) <= not((layer1_outputs(5275)) or (layer1_outputs(8414)));
    layer2_outputs(6947) <= not((layer1_outputs(259)) or (layer1_outputs(4637)));
    layer2_outputs(6948) <= (layer1_outputs(1046)) and (layer1_outputs(5800));
    layer2_outputs(6949) <= (layer1_outputs(5722)) and not (layer1_outputs(9353));
    layer2_outputs(6950) <= not(layer1_outputs(2282)) or (layer1_outputs(10199));
    layer2_outputs(6951) <= layer1_outputs(9123);
    layer2_outputs(6952) <= layer1_outputs(1061);
    layer2_outputs(6953) <= not((layer1_outputs(9342)) xor (layer1_outputs(2384)));
    layer2_outputs(6954) <= layer1_outputs(1505);
    layer2_outputs(6955) <= (layer1_outputs(6473)) or (layer1_outputs(9290));
    layer2_outputs(6956) <= (layer1_outputs(6803)) or (layer1_outputs(7850));
    layer2_outputs(6957) <= not(layer1_outputs(8758));
    layer2_outputs(6958) <= (layer1_outputs(6375)) or (layer1_outputs(7224));
    layer2_outputs(6959) <= (layer1_outputs(3321)) and (layer1_outputs(6833));
    layer2_outputs(6960) <= (layer1_outputs(5363)) and not (layer1_outputs(2834));
    layer2_outputs(6961) <= not(layer1_outputs(1597));
    layer2_outputs(6962) <= (layer1_outputs(7877)) or (layer1_outputs(8478));
    layer2_outputs(6963) <= (layer1_outputs(7797)) xor (layer1_outputs(8505));
    layer2_outputs(6964) <= not((layer1_outputs(3506)) or (layer1_outputs(2916)));
    layer2_outputs(6965) <= not((layer1_outputs(7169)) xor (layer1_outputs(2508)));
    layer2_outputs(6966) <= not(layer1_outputs(2783));
    layer2_outputs(6967) <= (layer1_outputs(8583)) and not (layer1_outputs(3531));
    layer2_outputs(6968) <= not(layer1_outputs(4336));
    layer2_outputs(6969) <= (layer1_outputs(50)) and not (layer1_outputs(2529));
    layer2_outputs(6970) <= not((layer1_outputs(6458)) and (layer1_outputs(5197)));
    layer2_outputs(6971) <= (layer1_outputs(8794)) or (layer1_outputs(3598));
    layer2_outputs(6972) <= '1';
    layer2_outputs(6973) <= layer1_outputs(7682);
    layer2_outputs(6974) <= (layer1_outputs(84)) and not (layer1_outputs(5901));
    layer2_outputs(6975) <= (layer1_outputs(10016)) or (layer1_outputs(1321));
    layer2_outputs(6976) <= (layer1_outputs(2637)) or (layer1_outputs(1572));
    layer2_outputs(6977) <= (layer1_outputs(5503)) xor (layer1_outputs(5877));
    layer2_outputs(6978) <= layer1_outputs(9222);
    layer2_outputs(6979) <= (layer1_outputs(7297)) and not (layer1_outputs(7418));
    layer2_outputs(6980) <= not((layer1_outputs(2699)) or (layer1_outputs(6489)));
    layer2_outputs(6981) <= not(layer1_outputs(7638)) or (layer1_outputs(1924));
    layer2_outputs(6982) <= not(layer1_outputs(8655));
    layer2_outputs(6983) <= '0';
    layer2_outputs(6984) <= (layer1_outputs(2177)) xor (layer1_outputs(6798));
    layer2_outputs(6985) <= not(layer1_outputs(4085)) or (layer1_outputs(3383));
    layer2_outputs(6986) <= (layer1_outputs(6900)) and (layer1_outputs(8692));
    layer2_outputs(6987) <= (layer1_outputs(439)) and (layer1_outputs(8501));
    layer2_outputs(6988) <= not(layer1_outputs(6400)) or (layer1_outputs(3427));
    layer2_outputs(6989) <= not(layer1_outputs(2365));
    layer2_outputs(6990) <= not((layer1_outputs(2104)) xor (layer1_outputs(4511)));
    layer2_outputs(6991) <= layer1_outputs(7236);
    layer2_outputs(6992) <= not(layer1_outputs(5582));
    layer2_outputs(6993) <= not((layer1_outputs(7127)) and (layer1_outputs(9868)));
    layer2_outputs(6994) <= (layer1_outputs(9746)) and not (layer1_outputs(6443));
    layer2_outputs(6995) <= (layer1_outputs(6777)) and not (layer1_outputs(2270));
    layer2_outputs(6996) <= not(layer1_outputs(3167)) or (layer1_outputs(7849));
    layer2_outputs(6997) <= not(layer1_outputs(4885));
    layer2_outputs(6998) <= layer1_outputs(9862);
    layer2_outputs(6999) <= not(layer1_outputs(1815));
    layer2_outputs(7000) <= (layer1_outputs(3616)) and not (layer1_outputs(7524));
    layer2_outputs(7001) <= not((layer1_outputs(2312)) and (layer1_outputs(4008)));
    layer2_outputs(7002) <= not(layer1_outputs(6879));
    layer2_outputs(7003) <= not(layer1_outputs(9080));
    layer2_outputs(7004) <= not(layer1_outputs(5770));
    layer2_outputs(7005) <= not((layer1_outputs(8675)) xor (layer1_outputs(6035)));
    layer2_outputs(7006) <= layer1_outputs(2006);
    layer2_outputs(7007) <= not((layer1_outputs(5589)) or (layer1_outputs(5643)));
    layer2_outputs(7008) <= not(layer1_outputs(7037));
    layer2_outputs(7009) <= not(layer1_outputs(3353));
    layer2_outputs(7010) <= layer1_outputs(8526);
    layer2_outputs(7011) <= not(layer1_outputs(2843)) or (layer1_outputs(1640));
    layer2_outputs(7012) <= not((layer1_outputs(7129)) or (layer1_outputs(6925)));
    layer2_outputs(7013) <= (layer1_outputs(8666)) or (layer1_outputs(6291));
    layer2_outputs(7014) <= not((layer1_outputs(4557)) and (layer1_outputs(918)));
    layer2_outputs(7015) <= (layer1_outputs(2379)) or (layer1_outputs(3165));
    layer2_outputs(7016) <= (layer1_outputs(5622)) and not (layer1_outputs(4330));
    layer2_outputs(7017) <= not(layer1_outputs(4889));
    layer2_outputs(7018) <= layer1_outputs(592);
    layer2_outputs(7019) <= '1';
    layer2_outputs(7020) <= layer1_outputs(8886);
    layer2_outputs(7021) <= not((layer1_outputs(6941)) or (layer1_outputs(5824)));
    layer2_outputs(7022) <= (layer1_outputs(5342)) or (layer1_outputs(7506));
    layer2_outputs(7023) <= (layer1_outputs(3765)) or (layer1_outputs(3756));
    layer2_outputs(7024) <= not(layer1_outputs(8626));
    layer2_outputs(7025) <= not(layer1_outputs(6651));
    layer2_outputs(7026) <= (layer1_outputs(578)) or (layer1_outputs(8183));
    layer2_outputs(7027) <= not(layer1_outputs(10128)) or (layer1_outputs(7477));
    layer2_outputs(7028) <= not(layer1_outputs(7717));
    layer2_outputs(7029) <= not((layer1_outputs(3825)) or (layer1_outputs(3482)));
    layer2_outputs(7030) <= not(layer1_outputs(5535)) or (layer1_outputs(5271));
    layer2_outputs(7031) <= not(layer1_outputs(1404));
    layer2_outputs(7032) <= '0';
    layer2_outputs(7033) <= not(layer1_outputs(9970)) or (layer1_outputs(4373));
    layer2_outputs(7034) <= not(layer1_outputs(6093));
    layer2_outputs(7035) <= not(layer1_outputs(6120));
    layer2_outputs(7036) <= (layer1_outputs(5517)) or (layer1_outputs(5779));
    layer2_outputs(7037) <= not((layer1_outputs(3029)) and (layer1_outputs(5094)));
    layer2_outputs(7038) <= layer1_outputs(7745);
    layer2_outputs(7039) <= layer1_outputs(3387);
    layer2_outputs(7040) <= layer1_outputs(4320);
    layer2_outputs(7041) <= layer1_outputs(2483);
    layer2_outputs(7042) <= not(layer1_outputs(8972)) or (layer1_outputs(2312));
    layer2_outputs(7043) <= not(layer1_outputs(9965));
    layer2_outputs(7044) <= (layer1_outputs(7361)) and not (layer1_outputs(9778));
    layer2_outputs(7045) <= layer1_outputs(6223);
    layer2_outputs(7046) <= layer1_outputs(6461);
    layer2_outputs(7047) <= layer1_outputs(9036);
    layer2_outputs(7048) <= '1';
    layer2_outputs(7049) <= not((layer1_outputs(459)) and (layer1_outputs(7510)));
    layer2_outputs(7050) <= (layer1_outputs(5910)) xor (layer1_outputs(5358));
    layer2_outputs(7051) <= layer1_outputs(2967);
    layer2_outputs(7052) <= not(layer1_outputs(5495)) or (layer1_outputs(3374));
    layer2_outputs(7053) <= layer1_outputs(10090);
    layer2_outputs(7054) <= layer1_outputs(7192);
    layer2_outputs(7055) <= not(layer1_outputs(21)) or (layer1_outputs(2340));
    layer2_outputs(7056) <= layer1_outputs(1615);
    layer2_outputs(7057) <= not(layer1_outputs(2752)) or (layer1_outputs(6245));
    layer2_outputs(7058) <= not(layer1_outputs(4092)) or (layer1_outputs(7907));
    layer2_outputs(7059) <= '0';
    layer2_outputs(7060) <= '1';
    layer2_outputs(7061) <= layer1_outputs(8691);
    layer2_outputs(7062) <= layer1_outputs(4148);
    layer2_outputs(7063) <= (layer1_outputs(9300)) and not (layer1_outputs(9500));
    layer2_outputs(7064) <= not(layer1_outputs(8663));
    layer2_outputs(7065) <= not(layer1_outputs(856));
    layer2_outputs(7066) <= not((layer1_outputs(7830)) xor (layer1_outputs(3338)));
    layer2_outputs(7067) <= not(layer1_outputs(4827)) or (layer1_outputs(8124));
    layer2_outputs(7068) <= layer1_outputs(8187);
    layer2_outputs(7069) <= (layer1_outputs(6568)) or (layer1_outputs(8814));
    layer2_outputs(7070) <= not((layer1_outputs(9259)) and (layer1_outputs(5087)));
    layer2_outputs(7071) <= (layer1_outputs(5750)) or (layer1_outputs(6307));
    layer2_outputs(7072) <= not((layer1_outputs(3705)) and (layer1_outputs(6561)));
    layer2_outputs(7073) <= layer1_outputs(8578);
    layer2_outputs(7074) <= not((layer1_outputs(1341)) and (layer1_outputs(2438)));
    layer2_outputs(7075) <= not((layer1_outputs(5183)) or (layer1_outputs(9452)));
    layer2_outputs(7076) <= not(layer1_outputs(8462));
    layer2_outputs(7077) <= layer1_outputs(4425);
    layer2_outputs(7078) <= not(layer1_outputs(193)) or (layer1_outputs(2639));
    layer2_outputs(7079) <= not(layer1_outputs(9520)) or (layer1_outputs(6731));
    layer2_outputs(7080) <= (layer1_outputs(2679)) and not (layer1_outputs(1881));
    layer2_outputs(7081) <= not((layer1_outputs(6209)) or (layer1_outputs(4767)));
    layer2_outputs(7082) <= (layer1_outputs(7980)) or (layer1_outputs(5855));
    layer2_outputs(7083) <= not((layer1_outputs(402)) xor (layer1_outputs(9779)));
    layer2_outputs(7084) <= not(layer1_outputs(6486));
    layer2_outputs(7085) <= not(layer1_outputs(5011));
    layer2_outputs(7086) <= not(layer1_outputs(4759)) or (layer1_outputs(7963));
    layer2_outputs(7087) <= (layer1_outputs(1105)) xor (layer1_outputs(4075));
    layer2_outputs(7088) <= not(layer1_outputs(8840));
    layer2_outputs(7089) <= (layer1_outputs(8618)) and (layer1_outputs(5250));
    layer2_outputs(7090) <= not(layer1_outputs(7853));
    layer2_outputs(7091) <= '0';
    layer2_outputs(7092) <= not(layer1_outputs(5700));
    layer2_outputs(7093) <= not(layer1_outputs(5780)) or (layer1_outputs(8234));
    layer2_outputs(7094) <= not(layer1_outputs(4342));
    layer2_outputs(7095) <= layer1_outputs(6981);
    layer2_outputs(7096) <= not(layer1_outputs(227)) or (layer1_outputs(4650));
    layer2_outputs(7097) <= layer1_outputs(5091);
    layer2_outputs(7098) <= not(layer1_outputs(7799));
    layer2_outputs(7099) <= not(layer1_outputs(9984)) or (layer1_outputs(9670));
    layer2_outputs(7100) <= not((layer1_outputs(2736)) xor (layer1_outputs(6749)));
    layer2_outputs(7101) <= (layer1_outputs(425)) and not (layer1_outputs(3397));
    layer2_outputs(7102) <= not(layer1_outputs(446));
    layer2_outputs(7103) <= layer1_outputs(5429);
    layer2_outputs(7104) <= layer1_outputs(9442);
    layer2_outputs(7105) <= (layer1_outputs(5667)) and (layer1_outputs(8059));
    layer2_outputs(7106) <= '1';
    layer2_outputs(7107) <= (layer1_outputs(1106)) xor (layer1_outputs(1497));
    layer2_outputs(7108) <= (layer1_outputs(8108)) and not (layer1_outputs(5424));
    layer2_outputs(7109) <= not((layer1_outputs(9055)) or (layer1_outputs(2634)));
    layer2_outputs(7110) <= not(layer1_outputs(7958));
    layer2_outputs(7111) <= not(layer1_outputs(5891));
    layer2_outputs(7112) <= '1';
    layer2_outputs(7113) <= (layer1_outputs(10142)) or (layer1_outputs(137));
    layer2_outputs(7114) <= layer1_outputs(3443);
    layer2_outputs(7115) <= layer1_outputs(5300);
    layer2_outputs(7116) <= '0';
    layer2_outputs(7117) <= (layer1_outputs(713)) and (layer1_outputs(4014));
    layer2_outputs(7118) <= not(layer1_outputs(2373)) or (layer1_outputs(3180));
    layer2_outputs(7119) <= '0';
    layer2_outputs(7120) <= (layer1_outputs(6152)) xor (layer1_outputs(570));
    layer2_outputs(7121) <= '0';
    layer2_outputs(7122) <= (layer1_outputs(6259)) and not (layer1_outputs(5192));
    layer2_outputs(7123) <= (layer1_outputs(9647)) and not (layer1_outputs(3017));
    layer2_outputs(7124) <= (layer1_outputs(5740)) or (layer1_outputs(2832));
    layer2_outputs(7125) <= layer1_outputs(1231);
    layer2_outputs(7126) <= (layer1_outputs(765)) and not (layer1_outputs(7473));
    layer2_outputs(7127) <= (layer1_outputs(1351)) and not (layer1_outputs(7817));
    layer2_outputs(7128) <= layer1_outputs(5193);
    layer2_outputs(7129) <= (layer1_outputs(9359)) and (layer1_outputs(5198));
    layer2_outputs(7130) <= (layer1_outputs(5851)) and not (layer1_outputs(10077));
    layer2_outputs(7131) <= not(layer1_outputs(5100));
    layer2_outputs(7132) <= (layer1_outputs(8324)) and (layer1_outputs(4791));
    layer2_outputs(7133) <= not(layer1_outputs(6740));
    layer2_outputs(7134) <= not(layer1_outputs(9987));
    layer2_outputs(7135) <= not((layer1_outputs(6795)) xor (layer1_outputs(2508)));
    layer2_outputs(7136) <= not(layer1_outputs(1039)) or (layer1_outputs(7524));
    layer2_outputs(7137) <= not(layer1_outputs(3416));
    layer2_outputs(7138) <= not(layer1_outputs(6934));
    layer2_outputs(7139) <= not((layer1_outputs(8247)) or (layer1_outputs(798)));
    layer2_outputs(7140) <= not((layer1_outputs(8645)) and (layer1_outputs(6642)));
    layer2_outputs(7141) <= not(layer1_outputs(2502));
    layer2_outputs(7142) <= (layer1_outputs(112)) xor (layer1_outputs(8185));
    layer2_outputs(7143) <= layer1_outputs(8423);
    layer2_outputs(7144) <= (layer1_outputs(111)) and not (layer1_outputs(1290));
    layer2_outputs(7145) <= (layer1_outputs(5279)) or (layer1_outputs(3367));
    layer2_outputs(7146) <= (layer1_outputs(8513)) xor (layer1_outputs(9169));
    layer2_outputs(7147) <= layer1_outputs(5827);
    layer2_outputs(7148) <= (layer1_outputs(7906)) or (layer1_outputs(5146));
    layer2_outputs(7149) <= layer1_outputs(2482);
    layer2_outputs(7150) <= layer1_outputs(8167);
    layer2_outputs(7151) <= layer1_outputs(1369);
    layer2_outputs(7152) <= layer1_outputs(8502);
    layer2_outputs(7153) <= not(layer1_outputs(5141)) or (layer1_outputs(6540));
    layer2_outputs(7154) <= not((layer1_outputs(9454)) or (layer1_outputs(3503)));
    layer2_outputs(7155) <= layer1_outputs(1550);
    layer2_outputs(7156) <= layer1_outputs(9281);
    layer2_outputs(7157) <= (layer1_outputs(1803)) or (layer1_outputs(1473));
    layer2_outputs(7158) <= layer1_outputs(2916);
    layer2_outputs(7159) <= (layer1_outputs(10131)) and not (layer1_outputs(692));
    layer2_outputs(7160) <= (layer1_outputs(3299)) and (layer1_outputs(3842));
    layer2_outputs(7161) <= not(layer1_outputs(8564)) or (layer1_outputs(2775));
    layer2_outputs(7162) <= layer1_outputs(7946);
    layer2_outputs(7163) <= (layer1_outputs(8541)) or (layer1_outputs(3959));
    layer2_outputs(7164) <= not((layer1_outputs(7732)) xor (layer1_outputs(9208)));
    layer2_outputs(7165) <= (layer1_outputs(4741)) and not (layer1_outputs(8677));
    layer2_outputs(7166) <= '0';
    layer2_outputs(7167) <= not(layer1_outputs(1368)) or (layer1_outputs(975));
    layer2_outputs(7168) <= not(layer1_outputs(338)) or (layer1_outputs(6242));
    layer2_outputs(7169) <= not(layer1_outputs(2738));
    layer2_outputs(7170) <= '0';
    layer2_outputs(7171) <= not(layer1_outputs(9682)) or (layer1_outputs(498));
    layer2_outputs(7172) <= not(layer1_outputs(8521));
    layer2_outputs(7173) <= not(layer1_outputs(1068));
    layer2_outputs(7174) <= layer1_outputs(2886);
    layer2_outputs(7175) <= (layer1_outputs(195)) xor (layer1_outputs(1083));
    layer2_outputs(7176) <= not(layer1_outputs(9620)) or (layer1_outputs(431));
    layer2_outputs(7177) <= '1';
    layer2_outputs(7178) <= (layer1_outputs(1087)) or (layer1_outputs(9367));
    layer2_outputs(7179) <= layer1_outputs(770);
    layer2_outputs(7180) <= not((layer1_outputs(9580)) or (layer1_outputs(5899)));
    layer2_outputs(7181) <= not(layer1_outputs(6512));
    layer2_outputs(7182) <= not(layer1_outputs(8917));
    layer2_outputs(7183) <= not(layer1_outputs(4663));
    layer2_outputs(7184) <= not((layer1_outputs(9098)) or (layer1_outputs(9560)));
    layer2_outputs(7185) <= not(layer1_outputs(4293));
    layer2_outputs(7186) <= '1';
    layer2_outputs(7187) <= (layer1_outputs(4502)) or (layer1_outputs(4233));
    layer2_outputs(7188) <= (layer1_outputs(1653)) and not (layer1_outputs(3805));
    layer2_outputs(7189) <= layer1_outputs(5938);
    layer2_outputs(7190) <= (layer1_outputs(3010)) and (layer1_outputs(4872));
    layer2_outputs(7191) <= layer1_outputs(3792);
    layer2_outputs(7192) <= not(layer1_outputs(1666));
    layer2_outputs(7193) <= not(layer1_outputs(2361)) or (layer1_outputs(7872));
    layer2_outputs(7194) <= not(layer1_outputs(587)) or (layer1_outputs(51));
    layer2_outputs(7195) <= '0';
    layer2_outputs(7196) <= (layer1_outputs(880)) and not (layer1_outputs(3644));
    layer2_outputs(7197) <= not((layer1_outputs(6733)) xor (layer1_outputs(3901)));
    layer2_outputs(7198) <= (layer1_outputs(7015)) and not (layer1_outputs(6216));
    layer2_outputs(7199) <= not((layer1_outputs(937)) xor (layer1_outputs(1724)));
    layer2_outputs(7200) <= not(layer1_outputs(4594));
    layer2_outputs(7201) <= (layer1_outputs(4063)) and (layer1_outputs(3988));
    layer2_outputs(7202) <= (layer1_outputs(4074)) and (layer1_outputs(4341));
    layer2_outputs(7203) <= layer1_outputs(951);
    layer2_outputs(7204) <= '0';
    layer2_outputs(7205) <= (layer1_outputs(6909)) and not (layer1_outputs(9573));
    layer2_outputs(7206) <= '0';
    layer2_outputs(7207) <= layer1_outputs(1334);
    layer2_outputs(7208) <= not((layer1_outputs(7335)) and (layer1_outputs(4009)));
    layer2_outputs(7209) <= not(layer1_outputs(28)) or (layer1_outputs(10236));
    layer2_outputs(7210) <= not(layer1_outputs(2643)) or (layer1_outputs(8333));
    layer2_outputs(7211) <= (layer1_outputs(5809)) and (layer1_outputs(9880));
    layer2_outputs(7212) <= layer1_outputs(3588);
    layer2_outputs(7213) <= layer1_outputs(2978);
    layer2_outputs(7214) <= (layer1_outputs(1749)) and (layer1_outputs(6860));
    layer2_outputs(7215) <= (layer1_outputs(8289)) and not (layer1_outputs(3164));
    layer2_outputs(7216) <= (layer1_outputs(4209)) and not (layer1_outputs(1744));
    layer2_outputs(7217) <= layer1_outputs(1054);
    layer2_outputs(7218) <= not(layer1_outputs(977)) or (layer1_outputs(6423));
    layer2_outputs(7219) <= layer1_outputs(7614);
    layer2_outputs(7220) <= '1';
    layer2_outputs(7221) <= layer1_outputs(2816);
    layer2_outputs(7222) <= layer1_outputs(5322);
    layer2_outputs(7223) <= layer1_outputs(6542);
    layer2_outputs(7224) <= not(layer1_outputs(5578));
    layer2_outputs(7225) <= not(layer1_outputs(4383));
    layer2_outputs(7226) <= '0';
    layer2_outputs(7227) <= not((layer1_outputs(190)) xor (layer1_outputs(7010)));
    layer2_outputs(7228) <= layer1_outputs(9258);
    layer2_outputs(7229) <= not(layer1_outputs(6789));
    layer2_outputs(7230) <= not((layer1_outputs(7944)) and (layer1_outputs(5588)));
    layer2_outputs(7231) <= layer1_outputs(2625);
    layer2_outputs(7232) <= (layer1_outputs(2622)) and (layer1_outputs(9470));
    layer2_outputs(7233) <= '0';
    layer2_outputs(7234) <= not(layer1_outputs(3062));
    layer2_outputs(7235) <= layer1_outputs(301);
    layer2_outputs(7236) <= not((layer1_outputs(4053)) xor (layer1_outputs(5656)));
    layer2_outputs(7237) <= (layer1_outputs(356)) and not (layer1_outputs(2267));
    layer2_outputs(7238) <= not((layer1_outputs(810)) xor (layer1_outputs(4056)));
    layer2_outputs(7239) <= layer1_outputs(1629);
    layer2_outputs(7240) <= layer1_outputs(7625);
    layer2_outputs(7241) <= not(layer1_outputs(5437));
    layer2_outputs(7242) <= not((layer1_outputs(1292)) and (layer1_outputs(6893)));
    layer2_outputs(7243) <= (layer1_outputs(538)) and not (layer1_outputs(6274));
    layer2_outputs(7244) <= (layer1_outputs(1087)) and not (layer1_outputs(7908));
    layer2_outputs(7245) <= (layer1_outputs(9788)) or (layer1_outputs(7852));
    layer2_outputs(7246) <= not(layer1_outputs(657));
    layer2_outputs(7247) <= layer1_outputs(7499);
    layer2_outputs(7248) <= not(layer1_outputs(2517));
    layer2_outputs(7249) <= layer1_outputs(6265);
    layer2_outputs(7250) <= '0';
    layer2_outputs(7251) <= not(layer1_outputs(7130)) or (layer1_outputs(686));
    layer2_outputs(7252) <= (layer1_outputs(7283)) or (layer1_outputs(3504));
    layer2_outputs(7253) <= not(layer1_outputs(2627)) or (layer1_outputs(2885));
    layer2_outputs(7254) <= not(layer1_outputs(600));
    layer2_outputs(7255) <= not((layer1_outputs(3369)) xor (layer1_outputs(4236)));
    layer2_outputs(7256) <= not(layer1_outputs(6592));
    layer2_outputs(7257) <= (layer1_outputs(9269)) and (layer1_outputs(8155));
    layer2_outputs(7258) <= not(layer1_outputs(8915)) or (layer1_outputs(5504));
    layer2_outputs(7259) <= layer1_outputs(3452);
    layer2_outputs(7260) <= '1';
    layer2_outputs(7261) <= layer1_outputs(5566);
    layer2_outputs(7262) <= not(layer1_outputs(3203));
    layer2_outputs(7263) <= layer1_outputs(2745);
    layer2_outputs(7264) <= '0';
    layer2_outputs(7265) <= layer1_outputs(865);
    layer2_outputs(7266) <= layer1_outputs(3479);
    layer2_outputs(7267) <= not(layer1_outputs(2797)) or (layer1_outputs(6874));
    layer2_outputs(7268) <= (layer1_outputs(6951)) and (layer1_outputs(9489));
    layer2_outputs(7269) <= not(layer1_outputs(2706));
    layer2_outputs(7270) <= not(layer1_outputs(5321));
    layer2_outputs(7271) <= not((layer1_outputs(2952)) xor (layer1_outputs(9884)));
    layer2_outputs(7272) <= '0';
    layer2_outputs(7273) <= (layer1_outputs(877)) or (layer1_outputs(9509));
    layer2_outputs(7274) <= (layer1_outputs(6650)) and not (layer1_outputs(7993));
    layer2_outputs(7275) <= not(layer1_outputs(1831));
    layer2_outputs(7276) <= not(layer1_outputs(4110)) or (layer1_outputs(4492));
    layer2_outputs(7277) <= not(layer1_outputs(3624));
    layer2_outputs(7278) <= (layer1_outputs(1189)) or (layer1_outputs(2891));
    layer2_outputs(7279) <= not(layer1_outputs(9933));
    layer2_outputs(7280) <= '0';
    layer2_outputs(7281) <= (layer1_outputs(1997)) and (layer1_outputs(5031));
    layer2_outputs(7282) <= (layer1_outputs(4338)) xor (layer1_outputs(8679));
    layer2_outputs(7283) <= not(layer1_outputs(8734)) or (layer1_outputs(6324));
    layer2_outputs(7284) <= not((layer1_outputs(8571)) or (layer1_outputs(2558)));
    layer2_outputs(7285) <= not((layer1_outputs(8654)) and (layer1_outputs(1489)));
    layer2_outputs(7286) <= layer1_outputs(8861);
    layer2_outputs(7287) <= layer1_outputs(8169);
    layer2_outputs(7288) <= not(layer1_outputs(6822)) or (layer1_outputs(1977));
    layer2_outputs(7289) <= not((layer1_outputs(941)) and (layer1_outputs(7181)));
    layer2_outputs(7290) <= layer1_outputs(1026);
    layer2_outputs(7291) <= '1';
    layer2_outputs(7292) <= not(layer1_outputs(7936));
    layer2_outputs(7293) <= not(layer1_outputs(10121));
    layer2_outputs(7294) <= (layer1_outputs(9600)) and not (layer1_outputs(2358));
    layer2_outputs(7295) <= not(layer1_outputs(4046));
    layer2_outputs(7296) <= (layer1_outputs(3812)) or (layer1_outputs(787));
    layer2_outputs(7297) <= layer1_outputs(2451);
    layer2_outputs(7298) <= layer1_outputs(5236);
    layer2_outputs(7299) <= not(layer1_outputs(1487));
    layer2_outputs(7300) <= (layer1_outputs(1931)) and not (layer1_outputs(2993));
    layer2_outputs(7301) <= not(layer1_outputs(6925));
    layer2_outputs(7302) <= not((layer1_outputs(2465)) or (layer1_outputs(9743)));
    layer2_outputs(7303) <= '0';
    layer2_outputs(7304) <= not((layer1_outputs(6519)) or (layer1_outputs(1792)));
    layer2_outputs(7305) <= layer1_outputs(4371);
    layer2_outputs(7306) <= '1';
    layer2_outputs(7307) <= layer1_outputs(3308);
    layer2_outputs(7308) <= not(layer1_outputs(4878));
    layer2_outputs(7309) <= not(layer1_outputs(8725)) or (layer1_outputs(7565));
    layer2_outputs(7310) <= not(layer1_outputs(1220));
    layer2_outputs(7311) <= not(layer1_outputs(5615));
    layer2_outputs(7312) <= layer1_outputs(9674);
    layer2_outputs(7313) <= '0';
    layer2_outputs(7314) <= layer1_outputs(3229);
    layer2_outputs(7315) <= not(layer1_outputs(7419)) or (layer1_outputs(2588));
    layer2_outputs(7316) <= not(layer1_outputs(4718));
    layer2_outputs(7317) <= not((layer1_outputs(9239)) and (layer1_outputs(1020)));
    layer2_outputs(7318) <= layer1_outputs(7420);
    layer2_outputs(7319) <= layer1_outputs(121);
    layer2_outputs(7320) <= not((layer1_outputs(3030)) xor (layer1_outputs(7086)));
    layer2_outputs(7321) <= '0';
    layer2_outputs(7322) <= not(layer1_outputs(3753)) or (layer1_outputs(10083));
    layer2_outputs(7323) <= '1';
    layer2_outputs(7324) <= layer1_outputs(8605);
    layer2_outputs(7325) <= not(layer1_outputs(8527));
    layer2_outputs(7326) <= '1';
    layer2_outputs(7327) <= (layer1_outputs(5320)) and (layer1_outputs(7048));
    layer2_outputs(7328) <= (layer1_outputs(4077)) or (layer1_outputs(8845));
    layer2_outputs(7329) <= not(layer1_outputs(7178));
    layer2_outputs(7330) <= layer1_outputs(4381);
    layer2_outputs(7331) <= (layer1_outputs(8609)) and not (layer1_outputs(9617));
    layer2_outputs(7332) <= (layer1_outputs(4758)) and not (layer1_outputs(4057));
    layer2_outputs(7333) <= not((layer1_outputs(8307)) and (layer1_outputs(9064)));
    layer2_outputs(7334) <= not(layer1_outputs(2076));
    layer2_outputs(7335) <= (layer1_outputs(2716)) and not (layer1_outputs(7815));
    layer2_outputs(7336) <= not((layer1_outputs(9455)) and (layer1_outputs(374)));
    layer2_outputs(7337) <= '0';
    layer2_outputs(7338) <= not((layer1_outputs(3130)) xor (layer1_outputs(8981)));
    layer2_outputs(7339) <= not((layer1_outputs(9942)) or (layer1_outputs(1195)));
    layer2_outputs(7340) <= not(layer1_outputs(5548));
    layer2_outputs(7341) <= (layer1_outputs(3972)) and not (layer1_outputs(3447));
    layer2_outputs(7342) <= (layer1_outputs(7577)) and not (layer1_outputs(1794));
    layer2_outputs(7343) <= layer1_outputs(10100);
    layer2_outputs(7344) <= not(layer1_outputs(10171)) or (layer1_outputs(1618));
    layer2_outputs(7345) <= not(layer1_outputs(775));
    layer2_outputs(7346) <= not(layer1_outputs(4456));
    layer2_outputs(7347) <= not(layer1_outputs(6819)) or (layer1_outputs(5219));
    layer2_outputs(7348) <= not(layer1_outputs(6871)) or (layer1_outputs(7112));
    layer2_outputs(7349) <= not((layer1_outputs(3729)) and (layer1_outputs(8597)));
    layer2_outputs(7350) <= (layer1_outputs(306)) or (layer1_outputs(9512));
    layer2_outputs(7351) <= not((layer1_outputs(6756)) or (layer1_outputs(4803)));
    layer2_outputs(7352) <= layer1_outputs(3348);
    layer2_outputs(7353) <= (layer1_outputs(1648)) and (layer1_outputs(6846));
    layer2_outputs(7354) <= '1';
    layer2_outputs(7355) <= not(layer1_outputs(2374)) or (layer1_outputs(8865));
    layer2_outputs(7356) <= not(layer1_outputs(6427));
    layer2_outputs(7357) <= (layer1_outputs(3217)) and (layer1_outputs(2382));
    layer2_outputs(7358) <= (layer1_outputs(2730)) and not (layer1_outputs(6689));
    layer2_outputs(7359) <= (layer1_outputs(5125)) or (layer1_outputs(3808));
    layer2_outputs(7360) <= not((layer1_outputs(3735)) and (layer1_outputs(1338)));
    layer2_outputs(7361) <= not(layer1_outputs(609));
    layer2_outputs(7362) <= '0';
    layer2_outputs(7363) <= layer1_outputs(9525);
    layer2_outputs(7364) <= not((layer1_outputs(7987)) xor (layer1_outputs(87)));
    layer2_outputs(7365) <= '1';
    layer2_outputs(7366) <= (layer1_outputs(6248)) and (layer1_outputs(4828));
    layer2_outputs(7367) <= layer1_outputs(7203);
    layer2_outputs(7368) <= layer1_outputs(1203);
    layer2_outputs(7369) <= (layer1_outputs(5302)) and (layer1_outputs(4159));
    layer2_outputs(7370) <= layer1_outputs(4339);
    layer2_outputs(7371) <= not((layer1_outputs(6674)) and (layer1_outputs(6992)));
    layer2_outputs(7372) <= not(layer1_outputs(1007));
    layer2_outputs(7373) <= not(layer1_outputs(3207)) or (layer1_outputs(10104));
    layer2_outputs(7374) <= not(layer1_outputs(9790));
    layer2_outputs(7375) <= not((layer1_outputs(6256)) xor (layer1_outputs(7000)));
    layer2_outputs(7376) <= not(layer1_outputs(1772));
    layer2_outputs(7377) <= not(layer1_outputs(6346)) or (layer1_outputs(9337));
    layer2_outputs(7378) <= not(layer1_outputs(9480));
    layer2_outputs(7379) <= (layer1_outputs(5583)) and not (layer1_outputs(7752));
    layer2_outputs(7380) <= not((layer1_outputs(1984)) or (layer1_outputs(9867)));
    layer2_outputs(7381) <= not((layer1_outputs(4766)) or (layer1_outputs(4618)));
    layer2_outputs(7382) <= (layer1_outputs(5779)) and (layer1_outputs(1013));
    layer2_outputs(7383) <= (layer1_outputs(9913)) or (layer1_outputs(5599));
    layer2_outputs(7384) <= layer1_outputs(2537);
    layer2_outputs(7385) <= (layer1_outputs(4214)) or (layer1_outputs(3938));
    layer2_outputs(7386) <= not((layer1_outputs(3599)) or (layer1_outputs(5337)));
    layer2_outputs(7387) <= not(layer1_outputs(2987)) or (layer1_outputs(6027));
    layer2_outputs(7388) <= layer1_outputs(5137);
    layer2_outputs(7389) <= not(layer1_outputs(3249));
    layer2_outputs(7390) <= (layer1_outputs(1129)) or (layer1_outputs(5276));
    layer2_outputs(7391) <= not(layer1_outputs(8106));
    layer2_outputs(7392) <= not(layer1_outputs(8904)) or (layer1_outputs(912));
    layer2_outputs(7393) <= (layer1_outputs(2397)) or (layer1_outputs(10165));
    layer2_outputs(7394) <= layer1_outputs(8868);
    layer2_outputs(7395) <= layer1_outputs(4858);
    layer2_outputs(7396) <= layer1_outputs(10173);
    layer2_outputs(7397) <= not((layer1_outputs(4584)) or (layer1_outputs(9607)));
    layer2_outputs(7398) <= layer1_outputs(9777);
    layer2_outputs(7399) <= layer1_outputs(8841);
    layer2_outputs(7400) <= (layer1_outputs(4762)) and not (layer1_outputs(6819));
    layer2_outputs(7401) <= not(layer1_outputs(1840));
    layer2_outputs(7402) <= (layer1_outputs(303)) and (layer1_outputs(1138));
    layer2_outputs(7403) <= (layer1_outputs(4520)) or (layer1_outputs(2961));
    layer2_outputs(7404) <= layer1_outputs(3886);
    layer2_outputs(7405) <= (layer1_outputs(4956)) and not (layer1_outputs(4721));
    layer2_outputs(7406) <= (layer1_outputs(7234)) and not (layer1_outputs(9001));
    layer2_outputs(7407) <= not((layer1_outputs(1355)) or (layer1_outputs(780)));
    layer2_outputs(7408) <= not(layer1_outputs(2774)) or (layer1_outputs(7202));
    layer2_outputs(7409) <= layer1_outputs(7961);
    layer2_outputs(7410) <= not(layer1_outputs(1529));
    layer2_outputs(7411) <= not(layer1_outputs(4174)) or (layer1_outputs(9069));
    layer2_outputs(7412) <= (layer1_outputs(6385)) or (layer1_outputs(6732));
    layer2_outputs(7413) <= (layer1_outputs(1807)) and not (layer1_outputs(9003));
    layer2_outputs(7414) <= (layer1_outputs(9167)) or (layer1_outputs(7541));
    layer2_outputs(7415) <= layer1_outputs(301);
    layer2_outputs(7416) <= not(layer1_outputs(7782)) or (layer1_outputs(608));
    layer2_outputs(7417) <= not(layer1_outputs(3011)) or (layer1_outputs(8642));
    layer2_outputs(7418) <= not(layer1_outputs(963));
    layer2_outputs(7419) <= not(layer1_outputs(2811));
    layer2_outputs(7420) <= (layer1_outputs(1952)) and (layer1_outputs(6526));
    layer2_outputs(7421) <= not(layer1_outputs(7771));
    layer2_outputs(7422) <= not(layer1_outputs(9809)) or (layer1_outputs(3171));
    layer2_outputs(7423) <= not(layer1_outputs(5866));
    layer2_outputs(7424) <= not(layer1_outputs(2833)) or (layer1_outputs(3105));
    layer2_outputs(7425) <= not((layer1_outputs(2629)) or (layer1_outputs(7088)));
    layer2_outputs(7426) <= not((layer1_outputs(2571)) and (layer1_outputs(10210)));
    layer2_outputs(7427) <= (layer1_outputs(4972)) and not (layer1_outputs(972));
    layer2_outputs(7428) <= '0';
    layer2_outputs(7429) <= (layer1_outputs(2092)) or (layer1_outputs(7835));
    layer2_outputs(7430) <= layer1_outputs(3039);
    layer2_outputs(7431) <= not((layer1_outputs(6815)) or (layer1_outputs(3359)));
    layer2_outputs(7432) <= (layer1_outputs(1799)) and not (layer1_outputs(7633));
    layer2_outputs(7433) <= '0';
    layer2_outputs(7434) <= (layer1_outputs(351)) or (layer1_outputs(8198));
    layer2_outputs(7435) <= not(layer1_outputs(8315)) or (layer1_outputs(1277));
    layer2_outputs(7436) <= (layer1_outputs(1349)) and not (layer1_outputs(6090));
    layer2_outputs(7437) <= (layer1_outputs(4214)) and not (layer1_outputs(1223));
    layer2_outputs(7438) <= not(layer1_outputs(9818)) or (layer1_outputs(7535));
    layer2_outputs(7439) <= (layer1_outputs(229)) and (layer1_outputs(1002));
    layer2_outputs(7440) <= (layer1_outputs(3837)) and (layer1_outputs(5349));
    layer2_outputs(7441) <= not(layer1_outputs(7735)) or (layer1_outputs(4896));
    layer2_outputs(7442) <= not(layer1_outputs(10034));
    layer2_outputs(7443) <= (layer1_outputs(2892)) and (layer1_outputs(4648));
    layer2_outputs(7444) <= (layer1_outputs(7982)) and not (layer1_outputs(3984));
    layer2_outputs(7445) <= not((layer1_outputs(4316)) xor (layer1_outputs(6625)));
    layer2_outputs(7446) <= not(layer1_outputs(1932)) or (layer1_outputs(9769));
    layer2_outputs(7447) <= not((layer1_outputs(9084)) and (layer1_outputs(9051)));
    layer2_outputs(7448) <= layer1_outputs(754);
    layer2_outputs(7449) <= not(layer1_outputs(6687)) or (layer1_outputs(2819));
    layer2_outputs(7450) <= '0';
    layer2_outputs(7451) <= not(layer1_outputs(196));
    layer2_outputs(7452) <= layer1_outputs(534);
    layer2_outputs(7453) <= not(layer1_outputs(6743)) or (layer1_outputs(4842));
    layer2_outputs(7454) <= not(layer1_outputs(3998));
    layer2_outputs(7455) <= (layer1_outputs(2101)) or (layer1_outputs(7572));
    layer2_outputs(7456) <= '1';
    layer2_outputs(7457) <= not((layer1_outputs(10167)) or (layer1_outputs(5019)));
    layer2_outputs(7458) <= layer1_outputs(5511);
    layer2_outputs(7459) <= layer1_outputs(5307);
    layer2_outputs(7460) <= not(layer1_outputs(5142));
    layer2_outputs(7461) <= layer1_outputs(5189);
    layer2_outputs(7462) <= not((layer1_outputs(9916)) or (layer1_outputs(1474)));
    layer2_outputs(7463) <= not(layer1_outputs(3697));
    layer2_outputs(7464) <= layer1_outputs(664);
    layer2_outputs(7465) <= layer1_outputs(1096);
    layer2_outputs(7466) <= not((layer1_outputs(5310)) and (layer1_outputs(8405)));
    layer2_outputs(7467) <= '1';
    layer2_outputs(7468) <= layer1_outputs(9606);
    layer2_outputs(7469) <= not(layer1_outputs(7486));
    layer2_outputs(7470) <= not(layer1_outputs(4643)) or (layer1_outputs(6287));
    layer2_outputs(7471) <= not(layer1_outputs(8279));
    layer2_outputs(7472) <= (layer1_outputs(3296)) xor (layer1_outputs(9254));
    layer2_outputs(7473) <= layer1_outputs(9150);
    layer2_outputs(7474) <= not(layer1_outputs(4513));
    layer2_outputs(7475) <= (layer1_outputs(6921)) and not (layer1_outputs(6325));
    layer2_outputs(7476) <= not(layer1_outputs(6574));
    layer2_outputs(7477) <= layer1_outputs(8081);
    layer2_outputs(7478) <= not(layer1_outputs(3179));
    layer2_outputs(7479) <= not(layer1_outputs(5321)) or (layer1_outputs(502));
    layer2_outputs(7480) <= not(layer1_outputs(5221));
    layer2_outputs(7481) <= not(layer1_outputs(2663));
    layer2_outputs(7482) <= not((layer1_outputs(3928)) xor (layer1_outputs(8871)));
    layer2_outputs(7483) <= not((layer1_outputs(5442)) and (layer1_outputs(6034)));
    layer2_outputs(7484) <= not(layer1_outputs(2940));
    layer2_outputs(7485) <= (layer1_outputs(3566)) or (layer1_outputs(9769));
    layer2_outputs(7486) <= (layer1_outputs(8475)) or (layer1_outputs(9649));
    layer2_outputs(7487) <= not(layer1_outputs(4595));
    layer2_outputs(7488) <= '1';
    layer2_outputs(7489) <= not(layer1_outputs(4349));
    layer2_outputs(7490) <= not(layer1_outputs(5151));
    layer2_outputs(7491) <= (layer1_outputs(8684)) and not (layer1_outputs(4979));
    layer2_outputs(7492) <= (layer1_outputs(7420)) and not (layer1_outputs(5044));
    layer2_outputs(7493) <= (layer1_outputs(5229)) and not (layer1_outputs(6529));
    layer2_outputs(7494) <= '1';
    layer2_outputs(7495) <= layer1_outputs(6252);
    layer2_outputs(7496) <= not((layer1_outputs(4883)) xor (layer1_outputs(2026)));
    layer2_outputs(7497) <= (layer1_outputs(3504)) and not (layer1_outputs(2204));
    layer2_outputs(7498) <= not((layer1_outputs(7250)) or (layer1_outputs(4431)));
    layer2_outputs(7499) <= not(layer1_outputs(5233));
    layer2_outputs(7500) <= (layer1_outputs(5310)) xor (layer1_outputs(852));
    layer2_outputs(7501) <= not((layer1_outputs(5982)) or (layer1_outputs(6889)));
    layer2_outputs(7502) <= not(layer1_outputs(8548)) or (layer1_outputs(4051));
    layer2_outputs(7503) <= not(layer1_outputs(6272));
    layer2_outputs(7504) <= (layer1_outputs(6813)) and (layer1_outputs(7206));
    layer2_outputs(7505) <= layer1_outputs(5479);
    layer2_outputs(7506) <= '1';
    layer2_outputs(7507) <= not(layer1_outputs(7891)) or (layer1_outputs(5608));
    layer2_outputs(7508) <= not(layer1_outputs(7960));
    layer2_outputs(7509) <= layer1_outputs(8420);
    layer2_outputs(7510) <= layer1_outputs(8924);
    layer2_outputs(7511) <= not((layer1_outputs(1835)) and (layer1_outputs(2842)));
    layer2_outputs(7512) <= (layer1_outputs(1351)) and (layer1_outputs(7103));
    layer2_outputs(7513) <= not((layer1_outputs(530)) or (layer1_outputs(6728)));
    layer2_outputs(7514) <= layer1_outputs(3348);
    layer2_outputs(7515) <= layer1_outputs(8381);
    layer2_outputs(7516) <= (layer1_outputs(8686)) and not (layer1_outputs(7167));
    layer2_outputs(7517) <= (layer1_outputs(2741)) and (layer1_outputs(1782));
    layer2_outputs(7518) <= (layer1_outputs(9034)) and not (layer1_outputs(3012));
    layer2_outputs(7519) <= (layer1_outputs(1897)) and not (layer1_outputs(2836));
    layer2_outputs(7520) <= not((layer1_outputs(10164)) or (layer1_outputs(5745)));
    layer2_outputs(7521) <= not(layer1_outputs(3768));
    layer2_outputs(7522) <= not(layer1_outputs(4660));
    layer2_outputs(7523) <= (layer1_outputs(1929)) xor (layer1_outputs(8208));
    layer2_outputs(7524) <= not(layer1_outputs(3206));
    layer2_outputs(7525) <= not(layer1_outputs(6825));
    layer2_outputs(7526) <= (layer1_outputs(2992)) and (layer1_outputs(5720));
    layer2_outputs(7527) <= layer1_outputs(1204);
    layer2_outputs(7528) <= not((layer1_outputs(6639)) and (layer1_outputs(206)));
    layer2_outputs(7529) <= (layer1_outputs(7214)) and not (layer1_outputs(5613));
    layer2_outputs(7530) <= not((layer1_outputs(581)) or (layer1_outputs(249)));
    layer2_outputs(7531) <= not(layer1_outputs(5850));
    layer2_outputs(7532) <= (layer1_outputs(9819)) or (layer1_outputs(1586));
    layer2_outputs(7533) <= not(layer1_outputs(5443));
    layer2_outputs(7534) <= layer1_outputs(4076);
    layer2_outputs(7535) <= layer1_outputs(5707);
    layer2_outputs(7536) <= not(layer1_outputs(2793)) or (layer1_outputs(7800));
    layer2_outputs(7537) <= layer1_outputs(2337);
    layer2_outputs(7538) <= not(layer1_outputs(4867));
    layer2_outputs(7539) <= layer1_outputs(7807);
    layer2_outputs(7540) <= '1';
    layer2_outputs(7541) <= not(layer1_outputs(6824));
    layer2_outputs(7542) <= not(layer1_outputs(1107));
    layer2_outputs(7543) <= not(layer1_outputs(2560));
    layer2_outputs(7544) <= not((layer1_outputs(3671)) and (layer1_outputs(9159)));
    layer2_outputs(7545) <= (layer1_outputs(8751)) or (layer1_outputs(4010));
    layer2_outputs(7546) <= not(layer1_outputs(457));
    layer2_outputs(7547) <= not(layer1_outputs(3770));
    layer2_outputs(7548) <= not(layer1_outputs(4350)) or (layer1_outputs(1048));
    layer2_outputs(7549) <= not(layer1_outputs(8129));
    layer2_outputs(7550) <= (layer1_outputs(3963)) and (layer1_outputs(873));
    layer2_outputs(7551) <= not((layer1_outputs(894)) xor (layer1_outputs(5351)));
    layer2_outputs(7552) <= layer1_outputs(7084);
    layer2_outputs(7553) <= not((layer1_outputs(7590)) and (layer1_outputs(9598)));
    layer2_outputs(7554) <= not(layer1_outputs(1342));
    layer2_outputs(7555) <= (layer1_outputs(1125)) and not (layer1_outputs(4250));
    layer2_outputs(7556) <= not(layer1_outputs(8369));
    layer2_outputs(7557) <= (layer1_outputs(3987)) or (layer1_outputs(359));
    layer2_outputs(7558) <= (layer1_outputs(2913)) or (layer1_outputs(2594));
    layer2_outputs(7559) <= not((layer1_outputs(4228)) xor (layer1_outputs(1426)));
    layer2_outputs(7560) <= not(layer1_outputs(3684));
    layer2_outputs(7561) <= (layer1_outputs(1806)) or (layer1_outputs(7693));
    layer2_outputs(7562) <= layer1_outputs(8893);
    layer2_outputs(7563) <= not(layer1_outputs(5731));
    layer2_outputs(7564) <= layer1_outputs(3432);
    layer2_outputs(7565) <= not(layer1_outputs(5206)) or (layer1_outputs(1949));
    layer2_outputs(7566) <= (layer1_outputs(2552)) and not (layer1_outputs(197));
    layer2_outputs(7567) <= not(layer1_outputs(8680));
    layer2_outputs(7568) <= not(layer1_outputs(2114)) or (layer1_outputs(8840));
    layer2_outputs(7569) <= not(layer1_outputs(8289));
    layer2_outputs(7570) <= (layer1_outputs(7700)) and (layer1_outputs(7953));
    layer2_outputs(7571) <= not(layer1_outputs(7896));
    layer2_outputs(7572) <= (layer1_outputs(6087)) and not (layer1_outputs(8204));
    layer2_outputs(7573) <= not((layer1_outputs(8846)) or (layer1_outputs(6433)));
    layer2_outputs(7574) <= (layer1_outputs(5855)) xor (layer1_outputs(7466));
    layer2_outputs(7575) <= (layer1_outputs(9342)) and not (layer1_outputs(5925));
    layer2_outputs(7576) <= layer1_outputs(223);
    layer2_outputs(7577) <= layer1_outputs(876);
    layer2_outputs(7578) <= not((layer1_outputs(910)) or (layer1_outputs(8791)));
    layer2_outputs(7579) <= not(layer1_outputs(1678));
    layer2_outputs(7580) <= not((layer1_outputs(9094)) or (layer1_outputs(5222)));
    layer2_outputs(7581) <= not((layer1_outputs(4118)) xor (layer1_outputs(5594)));
    layer2_outputs(7582) <= (layer1_outputs(4004)) and not (layer1_outputs(4899));
    layer2_outputs(7583) <= (layer1_outputs(6716)) or (layer1_outputs(1124));
    layer2_outputs(7584) <= layer1_outputs(821);
    layer2_outputs(7585) <= (layer1_outputs(3749)) or (layer1_outputs(8580));
    layer2_outputs(7586) <= layer1_outputs(2873);
    layer2_outputs(7587) <= not((layer1_outputs(6193)) or (layer1_outputs(1925)));
    layer2_outputs(7588) <= layer1_outputs(9210);
    layer2_outputs(7589) <= not(layer1_outputs(3316));
    layer2_outputs(7590) <= layer1_outputs(3407);
    layer2_outputs(7591) <= layer1_outputs(1784);
    layer2_outputs(7592) <= layer1_outputs(2361);
    layer2_outputs(7593) <= layer1_outputs(2848);
    layer2_outputs(7594) <= not(layer1_outputs(6375));
    layer2_outputs(7595) <= layer1_outputs(7622);
    layer2_outputs(7596) <= layer1_outputs(7255);
    layer2_outputs(7597) <= not(layer1_outputs(952)) or (layer1_outputs(9956));
    layer2_outputs(7598) <= not(layer1_outputs(4583));
    layer2_outputs(7599) <= not((layer1_outputs(6258)) or (layer1_outputs(4943)));
    layer2_outputs(7600) <= layer1_outputs(3773);
    layer2_outputs(7601) <= not(layer1_outputs(438));
    layer2_outputs(7602) <= not(layer1_outputs(1314)) or (layer1_outputs(4165));
    layer2_outputs(7603) <= layer1_outputs(5082);
    layer2_outputs(7604) <= (layer1_outputs(1461)) and not (layer1_outputs(9898));
    layer2_outputs(7605) <= not(layer1_outputs(2209)) or (layer1_outputs(2028));
    layer2_outputs(7606) <= (layer1_outputs(3711)) and not (layer1_outputs(4393));
    layer2_outputs(7607) <= layer1_outputs(7267);
    layer2_outputs(7608) <= not((layer1_outputs(5481)) or (layer1_outputs(4955)));
    layer2_outputs(7609) <= not(layer1_outputs(8013));
    layer2_outputs(7610) <= (layer1_outputs(5261)) and not (layer1_outputs(1689));
    layer2_outputs(7611) <= (layer1_outputs(9226)) and (layer1_outputs(3027));
    layer2_outputs(7612) <= (layer1_outputs(9464)) and (layer1_outputs(9292));
    layer2_outputs(7613) <= (layer1_outputs(582)) and not (layer1_outputs(8095));
    layer2_outputs(7614) <= layer1_outputs(3474);
    layer2_outputs(7615) <= layer1_outputs(696);
    layer2_outputs(7616) <= not((layer1_outputs(4133)) or (layer1_outputs(8144)));
    layer2_outputs(7617) <= not((layer1_outputs(3537)) or (layer1_outputs(5173)));
    layer2_outputs(7618) <= not((layer1_outputs(998)) xor (layer1_outputs(4032)));
    layer2_outputs(7619) <= layer1_outputs(5011);
    layer2_outputs(7620) <= not((layer1_outputs(8271)) xor (layer1_outputs(8217)));
    layer2_outputs(7621) <= not(layer1_outputs(10211));
    layer2_outputs(7622) <= not(layer1_outputs(1179));
    layer2_outputs(7623) <= (layer1_outputs(4513)) xor (layer1_outputs(9623));
    layer2_outputs(7624) <= (layer1_outputs(5125)) or (layer1_outputs(1356));
    layer2_outputs(7625) <= layer1_outputs(2878);
    layer2_outputs(7626) <= (layer1_outputs(8895)) and not (layer1_outputs(1800));
    layer2_outputs(7627) <= not(layer1_outputs(6250)) or (layer1_outputs(5668));
    layer2_outputs(7628) <= layer1_outputs(2396);
    layer2_outputs(7629) <= layer1_outputs(4670);
    layer2_outputs(7630) <= not(layer1_outputs(3993)) or (layer1_outputs(7034));
    layer2_outputs(7631) <= not(layer1_outputs(2479));
    layer2_outputs(7632) <= (layer1_outputs(1659)) and not (layer1_outputs(5586));
    layer2_outputs(7633) <= not(layer1_outputs(660)) or (layer1_outputs(5112));
    layer2_outputs(7634) <= layer1_outputs(5298);
    layer2_outputs(7635) <= (layer1_outputs(7966)) and not (layer1_outputs(6543));
    layer2_outputs(7636) <= not(layer1_outputs(226)) or (layer1_outputs(10050));
    layer2_outputs(7637) <= not(layer1_outputs(9692));
    layer2_outputs(7638) <= not(layer1_outputs(748)) or (layer1_outputs(5343));
    layer2_outputs(7639) <= not((layer1_outputs(9397)) and (layer1_outputs(9863)));
    layer2_outputs(7640) <= not(layer1_outputs(9503)) or (layer1_outputs(953));
    layer2_outputs(7641) <= not(layer1_outputs(52)) or (layer1_outputs(957));
    layer2_outputs(7642) <= '0';
    layer2_outputs(7643) <= not(layer1_outputs(3781));
    layer2_outputs(7644) <= (layer1_outputs(5845)) and not (layer1_outputs(5270));
    layer2_outputs(7645) <= not((layer1_outputs(4331)) and (layer1_outputs(6714)));
    layer2_outputs(7646) <= (layer1_outputs(5542)) and not (layer1_outputs(6717));
    layer2_outputs(7647) <= layer1_outputs(7731);
    layer2_outputs(7648) <= not((layer1_outputs(984)) xor (layer1_outputs(3399)));
    layer2_outputs(7649) <= not(layer1_outputs(4690));
    layer2_outputs(7650) <= not(layer1_outputs(6879));
    layer2_outputs(7651) <= not(layer1_outputs(7221));
    layer2_outputs(7652) <= '1';
    layer2_outputs(7653) <= (layer1_outputs(4906)) and (layer1_outputs(1051));
    layer2_outputs(7654) <= not(layer1_outputs(1926));
    layer2_outputs(7655) <= '0';
    layer2_outputs(7656) <= layer1_outputs(3679);
    layer2_outputs(7657) <= (layer1_outputs(2369)) or (layer1_outputs(2073));
    layer2_outputs(7658) <= not((layer1_outputs(6631)) xor (layer1_outputs(5342)));
    layer2_outputs(7659) <= layer1_outputs(7076);
    layer2_outputs(7660) <= not(layer1_outputs(2262));
    layer2_outputs(7661) <= not((layer1_outputs(3925)) and (layer1_outputs(935)));
    layer2_outputs(7662) <= (layer1_outputs(8577)) and not (layer1_outputs(540));
    layer2_outputs(7663) <= not(layer1_outputs(2463));
    layer2_outputs(7664) <= layer1_outputs(4542);
    layer2_outputs(7665) <= not((layer1_outputs(4420)) or (layer1_outputs(2932)));
    layer2_outputs(7666) <= not(layer1_outputs(7433)) or (layer1_outputs(6222));
    layer2_outputs(7667) <= (layer1_outputs(5311)) and not (layer1_outputs(9075));
    layer2_outputs(7668) <= layer1_outputs(2882);
    layer2_outputs(7669) <= '0';
    layer2_outputs(7670) <= (layer1_outputs(2580)) and (layer1_outputs(6197));
    layer2_outputs(7671) <= (layer1_outputs(1610)) or (layer1_outputs(4218));
    layer2_outputs(7672) <= (layer1_outputs(9125)) and (layer1_outputs(3608));
    layer2_outputs(7673) <= not(layer1_outputs(6219));
    layer2_outputs(7674) <= not((layer1_outputs(2179)) and (layer1_outputs(1290)));
    layer2_outputs(7675) <= not(layer1_outputs(7060)) or (layer1_outputs(6379));
    layer2_outputs(7676) <= layer1_outputs(2423);
    layer2_outputs(7677) <= not((layer1_outputs(4912)) or (layer1_outputs(505)));
    layer2_outputs(7678) <= not(layer1_outputs(7047)) or (layer1_outputs(6935));
    layer2_outputs(7679) <= (layer1_outputs(9829)) and (layer1_outputs(3629));
    layer2_outputs(7680) <= (layer1_outputs(5461)) xor (layer1_outputs(3763));
    layer2_outputs(7681) <= not(layer1_outputs(6371)) or (layer1_outputs(218));
    layer2_outputs(7682) <= layer1_outputs(9184);
    layer2_outputs(7683) <= (layer1_outputs(584)) and (layer1_outputs(7813));
    layer2_outputs(7684) <= not(layer1_outputs(8787));
    layer2_outputs(7685) <= layer1_outputs(8644);
    layer2_outputs(7686) <= layer1_outputs(5644);
    layer2_outputs(7687) <= (layer1_outputs(2784)) and not (layer1_outputs(5884));
    layer2_outputs(7688) <= not(layer1_outputs(8389)) or (layer1_outputs(2550));
    layer2_outputs(7689) <= layer1_outputs(2634);
    layer2_outputs(7690) <= layer1_outputs(3626);
    layer2_outputs(7691) <= (layer1_outputs(5558)) and not (layer1_outputs(9853));
    layer2_outputs(7692) <= not(layer1_outputs(3588));
    layer2_outputs(7693) <= layer1_outputs(2703);
    layer2_outputs(7694) <= not((layer1_outputs(1662)) and (layer1_outputs(2773)));
    layer2_outputs(7695) <= (layer1_outputs(8143)) or (layer1_outputs(9368));
    layer2_outputs(7696) <= not(layer1_outputs(7082));
    layer2_outputs(7697) <= layer1_outputs(5794);
    layer2_outputs(7698) <= layer1_outputs(7294);
    layer2_outputs(7699) <= not(layer1_outputs(1755));
    layer2_outputs(7700) <= layer1_outputs(8267);
    layer2_outputs(7701) <= not(layer1_outputs(1865)) or (layer1_outputs(7495));
    layer2_outputs(7702) <= (layer1_outputs(3601)) xor (layer1_outputs(8224));
    layer2_outputs(7703) <= not(layer1_outputs(9443)) or (layer1_outputs(818));
    layer2_outputs(7704) <= not(layer1_outputs(7673)) or (layer1_outputs(6792));
    layer2_outputs(7705) <= layer1_outputs(6895);
    layer2_outputs(7706) <= not(layer1_outputs(7674));
    layer2_outputs(7707) <= (layer1_outputs(312)) or (layer1_outputs(3453));
    layer2_outputs(7708) <= (layer1_outputs(3639)) and not (layer1_outputs(8474));
    layer2_outputs(7709) <= (layer1_outputs(2895)) and not (layer1_outputs(2667));
    layer2_outputs(7710) <= not(layer1_outputs(4324)) or (layer1_outputs(5113));
    layer2_outputs(7711) <= layer1_outputs(8550);
    layer2_outputs(7712) <= not((layer1_outputs(3745)) or (layer1_outputs(7108)));
    layer2_outputs(7713) <= layer1_outputs(5638);
    layer2_outputs(7714) <= (layer1_outputs(10008)) and not (layer1_outputs(9755));
    layer2_outputs(7715) <= (layer1_outputs(9339)) xor (layer1_outputs(2492));
    layer2_outputs(7716) <= not(layer1_outputs(9166)) or (layer1_outputs(6912));
    layer2_outputs(7717) <= not(layer1_outputs(4361));
    layer2_outputs(7718) <= (layer1_outputs(4436)) xor (layer1_outputs(4153));
    layer2_outputs(7719) <= layer1_outputs(3658);
    layer2_outputs(7720) <= (layer1_outputs(8432)) and not (layer1_outputs(2505));
    layer2_outputs(7721) <= '0';
    layer2_outputs(7722) <= (layer1_outputs(7892)) xor (layer1_outputs(3745));
    layer2_outputs(7723) <= layer1_outputs(5806);
    layer2_outputs(7724) <= '0';
    layer2_outputs(7725) <= layer1_outputs(7980);
    layer2_outputs(7726) <= layer1_outputs(7197);
    layer2_outputs(7727) <= (layer1_outputs(1291)) or (layer1_outputs(4396));
    layer2_outputs(7728) <= layer1_outputs(5073);
    layer2_outputs(7729) <= not(layer1_outputs(5581));
    layer2_outputs(7730) <= not(layer1_outputs(67));
    layer2_outputs(7731) <= not((layer1_outputs(5065)) or (layer1_outputs(979)));
    layer2_outputs(7732) <= layer1_outputs(9749);
    layer2_outputs(7733) <= not(layer1_outputs(362));
    layer2_outputs(7734) <= not((layer1_outputs(6683)) or (layer1_outputs(4988)));
    layer2_outputs(7735) <= '1';
    layer2_outputs(7736) <= not(layer1_outputs(4595)) or (layer1_outputs(5624));
    layer2_outputs(7737) <= '1';
    layer2_outputs(7738) <= layer1_outputs(819);
    layer2_outputs(7739) <= layer1_outputs(2717);
    layer2_outputs(7740) <= (layer1_outputs(4956)) xor (layer1_outputs(4934));
    layer2_outputs(7741) <= layer1_outputs(9297);
    layer2_outputs(7742) <= not(layer1_outputs(8189)) or (layer1_outputs(3839));
    layer2_outputs(7743) <= not((layer1_outputs(1216)) and (layer1_outputs(7207)));
    layer2_outputs(7744) <= not(layer1_outputs(2085)) or (layer1_outputs(4088));
    layer2_outputs(7745) <= not(layer1_outputs(9720));
    layer2_outputs(7746) <= (layer1_outputs(8748)) xor (layer1_outputs(1607));
    layer2_outputs(7747) <= not(layer1_outputs(2415)) or (layer1_outputs(3148));
    layer2_outputs(7748) <= '1';
    layer2_outputs(7749) <= layer1_outputs(6667);
    layer2_outputs(7750) <= not((layer1_outputs(2893)) and (layer1_outputs(5571)));
    layer2_outputs(7751) <= not(layer1_outputs(4058));
    layer2_outputs(7752) <= not(layer1_outputs(7876));
    layer2_outputs(7753) <= not((layer1_outputs(589)) xor (layer1_outputs(7876)));
    layer2_outputs(7754) <= (layer1_outputs(665)) xor (layer1_outputs(8534));
    layer2_outputs(7755) <= layer1_outputs(496);
    layer2_outputs(7756) <= (layer1_outputs(1580)) or (layer1_outputs(3572));
    layer2_outputs(7757) <= not(layer1_outputs(7038));
    layer2_outputs(7758) <= (layer1_outputs(7985)) or (layer1_outputs(9006));
    layer2_outputs(7759) <= (layer1_outputs(4140)) and not (layer1_outputs(9833));
    layer2_outputs(7760) <= not(layer1_outputs(1003));
    layer2_outputs(7761) <= (layer1_outputs(2679)) and not (layer1_outputs(3031));
    layer2_outputs(7762) <= not((layer1_outputs(9590)) xor (layer1_outputs(3747)));
    layer2_outputs(7763) <= not((layer1_outputs(8505)) and (layer1_outputs(9235)));
    layer2_outputs(7764) <= '0';
    layer2_outputs(7765) <= not(layer1_outputs(6563));
    layer2_outputs(7766) <= (layer1_outputs(2564)) and not (layer1_outputs(9709));
    layer2_outputs(7767) <= '0';
    layer2_outputs(7768) <= layer1_outputs(1509);
    layer2_outputs(7769) <= not((layer1_outputs(6532)) and (layer1_outputs(6556)));
    layer2_outputs(7770) <= not(layer1_outputs(9197)) or (layer1_outputs(2256));
    layer2_outputs(7771) <= (layer1_outputs(10166)) and not (layer1_outputs(4550));
    layer2_outputs(7772) <= not(layer1_outputs(2722));
    layer2_outputs(7773) <= not(layer1_outputs(2991));
    layer2_outputs(7774) <= not(layer1_outputs(8355));
    layer2_outputs(7775) <= layer1_outputs(4716);
    layer2_outputs(7776) <= not(layer1_outputs(4327));
    layer2_outputs(7777) <= not((layer1_outputs(8341)) and (layer1_outputs(348)));
    layer2_outputs(7778) <= not(layer1_outputs(1251));
    layer2_outputs(7779) <= '1';
    layer2_outputs(7780) <= not((layer1_outputs(887)) and (layer1_outputs(6763)));
    layer2_outputs(7781) <= not(layer1_outputs(4507)) or (layer1_outputs(6301));
    layer2_outputs(7782) <= not(layer1_outputs(4351));
    layer2_outputs(7783) <= layer1_outputs(1817);
    layer2_outputs(7784) <= (layer1_outputs(135)) and not (layer1_outputs(9380));
    layer2_outputs(7785) <= layer1_outputs(8962);
    layer2_outputs(7786) <= not(layer1_outputs(2322)) or (layer1_outputs(2080));
    layer2_outputs(7787) <= layer1_outputs(2881);
    layer2_outputs(7788) <= not((layer1_outputs(2669)) or (layer1_outputs(388)));
    layer2_outputs(7789) <= not(layer1_outputs(9134));
    layer2_outputs(7790) <= layer1_outputs(4168);
    layer2_outputs(7791) <= not(layer1_outputs(1472));
    layer2_outputs(7792) <= layer1_outputs(8006);
    layer2_outputs(7793) <= layer1_outputs(9646);
    layer2_outputs(7794) <= not((layer1_outputs(4374)) and (layer1_outputs(7721)));
    layer2_outputs(7795) <= not(layer1_outputs(1336));
    layer2_outputs(7796) <= not((layer1_outputs(6804)) or (layer1_outputs(2536)));
    layer2_outputs(7797) <= not(layer1_outputs(9764));
    layer2_outputs(7798) <= layer1_outputs(80);
    layer2_outputs(7799) <= not(layer1_outputs(6061));
    layer2_outputs(7800) <= not(layer1_outputs(3718)) or (layer1_outputs(5041));
    layer2_outputs(7801) <= not((layer1_outputs(5454)) and (layer1_outputs(4012)));
    layer2_outputs(7802) <= layer1_outputs(7560);
    layer2_outputs(7803) <= (layer1_outputs(6377)) and not (layer1_outputs(7678));
    layer2_outputs(7804) <= not(layer1_outputs(9748)) or (layer1_outputs(1610));
    layer2_outputs(7805) <= not(layer1_outputs(6163));
    layer2_outputs(7806) <= layer1_outputs(2789);
    layer2_outputs(7807) <= (layer1_outputs(4757)) or (layer1_outputs(5212));
    layer2_outputs(7808) <= layer1_outputs(1010);
    layer2_outputs(7809) <= (layer1_outputs(59)) and not (layer1_outputs(1619));
    layer2_outputs(7810) <= (layer1_outputs(4212)) and not (layer1_outputs(3056));
    layer2_outputs(7811) <= layer1_outputs(2593);
    layer2_outputs(7812) <= not(layer1_outputs(7292)) or (layer1_outputs(9302));
    layer2_outputs(7813) <= '0';
    layer2_outputs(7814) <= (layer1_outputs(521)) and not (layer1_outputs(2329));
    layer2_outputs(7815) <= layer1_outputs(8650);
    layer2_outputs(7816) <= '0';
    layer2_outputs(7817) <= (layer1_outputs(3635)) or (layer1_outputs(36));
    layer2_outputs(7818) <= layer1_outputs(9340);
    layer2_outputs(7819) <= (layer1_outputs(5160)) or (layer1_outputs(6850));
    layer2_outputs(7820) <= not((layer1_outputs(6384)) xor (layer1_outputs(2714)));
    layer2_outputs(7821) <= not(layer1_outputs(5420)) or (layer1_outputs(1249));
    layer2_outputs(7822) <= not((layer1_outputs(6434)) xor (layer1_outputs(2424)));
    layer2_outputs(7823) <= not(layer1_outputs(6574));
    layer2_outputs(7824) <= not(layer1_outputs(2292)) or (layer1_outputs(8242));
    layer2_outputs(7825) <= '0';
    layer2_outputs(7826) <= layer1_outputs(1773);
    layer2_outputs(7827) <= (layer1_outputs(2178)) xor (layer1_outputs(8522));
    layer2_outputs(7828) <= layer1_outputs(683);
    layer2_outputs(7829) <= '1';
    layer2_outputs(7830) <= not(layer1_outputs(7418));
    layer2_outputs(7831) <= not(layer1_outputs(1160));
    layer2_outputs(7832) <= not((layer1_outputs(6837)) xor (layer1_outputs(3312)));
    layer2_outputs(7833) <= not(layer1_outputs(3882));
    layer2_outputs(7834) <= not(layer1_outputs(7478));
    layer2_outputs(7835) <= not(layer1_outputs(6244));
    layer2_outputs(7836) <= not((layer1_outputs(7017)) and (layer1_outputs(1750)));
    layer2_outputs(7837) <= layer1_outputs(4245);
    layer2_outputs(7838) <= '0';
    layer2_outputs(7839) <= not((layer1_outputs(10063)) xor (layer1_outputs(4024)));
    layer2_outputs(7840) <= (layer1_outputs(9900)) and (layer1_outputs(10127));
    layer2_outputs(7841) <= layer1_outputs(4292);
    layer2_outputs(7842) <= '1';
    layer2_outputs(7843) <= (layer1_outputs(7782)) and not (layer1_outputs(8054));
    layer2_outputs(7844) <= '1';
    layer2_outputs(7845) <= not(layer1_outputs(8132));
    layer2_outputs(7846) <= not(layer1_outputs(7183)) or (layer1_outputs(4141));
    layer2_outputs(7847) <= not(layer1_outputs(2068));
    layer2_outputs(7848) <= '1';
    layer2_outputs(7849) <= not(layer1_outputs(2739));
    layer2_outputs(7850) <= not(layer1_outputs(7103));
    layer2_outputs(7851) <= not(layer1_outputs(2523)) or (layer1_outputs(9851));
    layer2_outputs(7852) <= layer1_outputs(2678);
    layer2_outputs(7853) <= layer1_outputs(6086);
    layer2_outputs(7854) <= not(layer1_outputs(9942));
    layer2_outputs(7855) <= layer1_outputs(5826);
    layer2_outputs(7856) <= layer1_outputs(7037);
    layer2_outputs(7857) <= layer1_outputs(3961);
    layer2_outputs(7858) <= (layer1_outputs(4942)) or (layer1_outputs(5477));
    layer2_outputs(7859) <= not((layer1_outputs(2383)) xor (layer1_outputs(3978)));
    layer2_outputs(7860) <= layer1_outputs(1790);
    layer2_outputs(7861) <= layer1_outputs(2527);
    layer2_outputs(7862) <= not(layer1_outputs(8118));
    layer2_outputs(7863) <= layer1_outputs(5655);
    layer2_outputs(7864) <= not((layer1_outputs(7266)) xor (layer1_outputs(3496)));
    layer2_outputs(7865) <= not(layer1_outputs(6996));
    layer2_outputs(7866) <= not(layer1_outputs(9525));
    layer2_outputs(7867) <= not(layer1_outputs(6449));
    layer2_outputs(7868) <= not((layer1_outputs(9132)) xor (layer1_outputs(1582)));
    layer2_outputs(7869) <= not(layer1_outputs(2606)) or (layer1_outputs(7837));
    layer2_outputs(7870) <= not(layer1_outputs(5369)) or (layer1_outputs(7192));
    layer2_outputs(7871) <= not(layer1_outputs(3719));
    layer2_outputs(7872) <= (layer1_outputs(4712)) and not (layer1_outputs(6481));
    layer2_outputs(7873) <= not(layer1_outputs(2055)) or (layer1_outputs(9903));
    layer2_outputs(7874) <= '0';
    layer2_outputs(7875) <= (layer1_outputs(5361)) xor (layer1_outputs(2920));
    layer2_outputs(7876) <= (layer1_outputs(2321)) and not (layer1_outputs(7364));
    layer2_outputs(7877) <= (layer1_outputs(2720)) or (layer1_outputs(2542));
    layer2_outputs(7878) <= not(layer1_outputs(4548));
    layer2_outputs(7879) <= layer1_outputs(1570);
    layer2_outputs(7880) <= (layer1_outputs(5794)) or (layer1_outputs(4452));
    layer2_outputs(7881) <= not(layer1_outputs(6974));
    layer2_outputs(7882) <= layer1_outputs(1787);
    layer2_outputs(7883) <= not(layer1_outputs(1639));
    layer2_outputs(7884) <= not(layer1_outputs(7079));
    layer2_outputs(7885) <= (layer1_outputs(8875)) or (layer1_outputs(5952));
    layer2_outputs(7886) <= not(layer1_outputs(2148)) or (layer1_outputs(2051));
    layer2_outputs(7887) <= not(layer1_outputs(7665));
    layer2_outputs(7888) <= layer1_outputs(6642);
    layer2_outputs(7889) <= not((layer1_outputs(7413)) and (layer1_outputs(4573)));
    layer2_outputs(7890) <= not((layer1_outputs(276)) xor (layer1_outputs(1100)));
    layer2_outputs(7891) <= (layer1_outputs(423)) or (layer1_outputs(4675));
    layer2_outputs(7892) <= layer1_outputs(10225);
    layer2_outputs(7893) <= (layer1_outputs(6201)) and (layer1_outputs(6993));
    layer2_outputs(7894) <= (layer1_outputs(2844)) and not (layer1_outputs(1627));
    layer2_outputs(7895) <= layer1_outputs(9201);
    layer2_outputs(7896) <= not((layer1_outputs(8371)) xor (layer1_outputs(4545)));
    layer2_outputs(7897) <= not(layer1_outputs(2484));
    layer2_outputs(7898) <= layer1_outputs(1691);
    layer2_outputs(7899) <= not(layer1_outputs(2933));
    layer2_outputs(7900) <= not(layer1_outputs(1474));
    layer2_outputs(7901) <= not(layer1_outputs(8985));
    layer2_outputs(7902) <= layer1_outputs(9643);
    layer2_outputs(7903) <= not((layer1_outputs(3573)) and (layer1_outputs(9907)));
    layer2_outputs(7904) <= not(layer1_outputs(5374)) or (layer1_outputs(7507));
    layer2_outputs(7905) <= '1';
    layer2_outputs(7906) <= (layer1_outputs(1560)) and not (layer1_outputs(4984));
    layer2_outputs(7907) <= not(layer1_outputs(9023));
    layer2_outputs(7908) <= not(layer1_outputs(8516));
    layer2_outputs(7909) <= (layer1_outputs(422)) or (layer1_outputs(2526));
    layer2_outputs(7910) <= not(layer1_outputs(9318));
    layer2_outputs(7911) <= not(layer1_outputs(7532));
    layer2_outputs(7912) <= (layer1_outputs(7012)) and (layer1_outputs(6114));
    layer2_outputs(7913) <= layer1_outputs(7808);
    layer2_outputs(7914) <= layer1_outputs(3661);
    layer2_outputs(7915) <= layer1_outputs(7546);
    layer2_outputs(7916) <= (layer1_outputs(6788)) and not (layer1_outputs(3301));
    layer2_outputs(7917) <= (layer1_outputs(1617)) and not (layer1_outputs(1371));
    layer2_outputs(7918) <= not(layer1_outputs(2395));
    layer2_outputs(7919) <= not((layer1_outputs(5579)) or (layer1_outputs(10087)));
    layer2_outputs(7920) <= not(layer1_outputs(8679));
    layer2_outputs(7921) <= layer1_outputs(7401);
    layer2_outputs(7922) <= (layer1_outputs(4428)) and not (layer1_outputs(8137));
    layer2_outputs(7923) <= layer1_outputs(3739);
    layer2_outputs(7924) <= (layer1_outputs(5893)) and not (layer1_outputs(1611));
    layer2_outputs(7925) <= not((layer1_outputs(604)) or (layer1_outputs(2498)));
    layer2_outputs(7926) <= '1';
    layer2_outputs(7927) <= not(layer1_outputs(833));
    layer2_outputs(7928) <= (layer1_outputs(7131)) and (layer1_outputs(8349));
    layer2_outputs(7929) <= not(layer1_outputs(3237)) or (layer1_outputs(2133));
    layer2_outputs(7930) <= not(layer1_outputs(8261)) or (layer1_outputs(2418));
    layer2_outputs(7931) <= layer1_outputs(7628);
    layer2_outputs(7932) <= layer1_outputs(4579);
    layer2_outputs(7933) <= not((layer1_outputs(9180)) and (layer1_outputs(7222)));
    layer2_outputs(7934) <= (layer1_outputs(8936)) and not (layer1_outputs(6518));
    layer2_outputs(7935) <= not((layer1_outputs(1457)) and (layer1_outputs(1363)));
    layer2_outputs(7936) <= layer1_outputs(2368);
    layer2_outputs(7937) <= not((layer1_outputs(1647)) or (layer1_outputs(9261)));
    layer2_outputs(7938) <= (layer1_outputs(5921)) and (layer1_outputs(5414));
    layer2_outputs(7939) <= layer1_outputs(7771);
    layer2_outputs(7940) <= '1';
    layer2_outputs(7941) <= (layer1_outputs(2419)) and not (layer1_outputs(9153));
    layer2_outputs(7942) <= not((layer1_outputs(6496)) and (layer1_outputs(2138)));
    layer2_outputs(7943) <= not(layer1_outputs(5328)) or (layer1_outputs(6783));
    layer2_outputs(7944) <= (layer1_outputs(5776)) and not (layer1_outputs(4485));
    layer2_outputs(7945) <= (layer1_outputs(5752)) and (layer1_outputs(2036));
    layer2_outputs(7946) <= not(layer1_outputs(710)) or (layer1_outputs(5048));
    layer2_outputs(7947) <= (layer1_outputs(6856)) xor (layer1_outputs(9489));
    layer2_outputs(7948) <= layer1_outputs(8061);
    layer2_outputs(7949) <= (layer1_outputs(9378)) and not (layer1_outputs(7260));
    layer2_outputs(7950) <= not(layer1_outputs(4800));
    layer2_outputs(7951) <= not(layer1_outputs(117));
    layer2_outputs(7952) <= '0';
    layer2_outputs(7953) <= not(layer1_outputs(1583)) or (layer1_outputs(5593));
    layer2_outputs(7954) <= not((layer1_outputs(6140)) and (layer1_outputs(6520)));
    layer2_outputs(7955) <= not(layer1_outputs(6502)) or (layer1_outputs(6163));
    layer2_outputs(7956) <= layer1_outputs(4632);
    layer2_outputs(7957) <= not(layer1_outputs(7388)) or (layer1_outputs(4885));
    layer2_outputs(7958) <= layer1_outputs(5647);
    layer2_outputs(7959) <= layer1_outputs(1283);
    layer2_outputs(7960) <= not(layer1_outputs(8060));
    layer2_outputs(7961) <= layer1_outputs(3965);
    layer2_outputs(7962) <= (layer1_outputs(593)) and (layer1_outputs(6105));
    layer2_outputs(7963) <= not(layer1_outputs(3883)) or (layer1_outputs(8141));
    layer2_outputs(7964) <= layer1_outputs(4594);
    layer2_outputs(7965) <= layer1_outputs(476);
    layer2_outputs(7966) <= layer1_outputs(735);
    layer2_outputs(7967) <= not(layer1_outputs(6018));
    layer2_outputs(7968) <= not(layer1_outputs(3370));
    layer2_outputs(7969) <= layer1_outputs(5282);
    layer2_outputs(7970) <= not(layer1_outputs(2800));
    layer2_outputs(7971) <= not(layer1_outputs(1499));
    layer2_outputs(7972) <= not(layer1_outputs(7345));
    layer2_outputs(7973) <= not(layer1_outputs(1044));
    layer2_outputs(7974) <= not((layer1_outputs(572)) or (layer1_outputs(2802)));
    layer2_outputs(7975) <= not((layer1_outputs(8499)) xor (layer1_outputs(4013)));
    layer2_outputs(7976) <= layer1_outputs(7727);
    layer2_outputs(7977) <= not(layer1_outputs(8773)) or (layer1_outputs(2644));
    layer2_outputs(7978) <= (layer1_outputs(8943)) and not (layer1_outputs(7366));
    layer2_outputs(7979) <= not(layer1_outputs(1027));
    layer2_outputs(7980) <= not((layer1_outputs(4626)) or (layer1_outputs(4236)));
    layer2_outputs(7981) <= not(layer1_outputs(2627));
    layer2_outputs(7982) <= not(layer1_outputs(6592));
    layer2_outputs(7983) <= layer1_outputs(7635);
    layer2_outputs(7984) <= layer1_outputs(7336);
    layer2_outputs(7985) <= (layer1_outputs(10220)) and (layer1_outputs(6691));
    layer2_outputs(7986) <= (layer1_outputs(8726)) or (layer1_outputs(427));
    layer2_outputs(7987) <= layer1_outputs(8886);
    layer2_outputs(7988) <= not(layer1_outputs(3904));
    layer2_outputs(7989) <= not(layer1_outputs(9267));
    layer2_outputs(7990) <= not(layer1_outputs(9573));
    layer2_outputs(7991) <= not(layer1_outputs(2063));
    layer2_outputs(7992) <= not(layer1_outputs(3200));
    layer2_outputs(7993) <= not((layer1_outputs(33)) and (layer1_outputs(2676)));
    layer2_outputs(7994) <= not((layer1_outputs(1304)) or (layer1_outputs(7064)));
    layer2_outputs(7995) <= layer1_outputs(9718);
    layer2_outputs(7996) <= layer1_outputs(6902);
    layer2_outputs(7997) <= layer1_outputs(2333);
    layer2_outputs(7998) <= not(layer1_outputs(3107));
    layer2_outputs(7999) <= not(layer1_outputs(5921));
    layer2_outputs(8000) <= not(layer1_outputs(9715)) or (layer1_outputs(4587));
    layer2_outputs(8001) <= layer1_outputs(2766);
    layer2_outputs(8002) <= (layer1_outputs(6794)) or (layer1_outputs(8558));
    layer2_outputs(8003) <= (layer1_outputs(7623)) and not (layer1_outputs(8342));
    layer2_outputs(8004) <= not((layer1_outputs(5692)) and (layer1_outputs(4517)));
    layer2_outputs(8005) <= not(layer1_outputs(3371));
    layer2_outputs(8006) <= (layer1_outputs(9111)) and not (layer1_outputs(4267));
    layer2_outputs(8007) <= not(layer1_outputs(2945)) or (layer1_outputs(9034));
    layer2_outputs(8008) <= not(layer1_outputs(9729));
    layer2_outputs(8009) <= (layer1_outputs(8967)) and not (layer1_outputs(6843));
    layer2_outputs(8010) <= not(layer1_outputs(2810));
    layer2_outputs(8011) <= not(layer1_outputs(1934));
    layer2_outputs(8012) <= not(layer1_outputs(8427));
    layer2_outputs(8013) <= (layer1_outputs(10126)) xor (layer1_outputs(7865));
    layer2_outputs(8014) <= layer1_outputs(8768);
    layer2_outputs(8015) <= layer1_outputs(1308);
    layer2_outputs(8016) <= layer1_outputs(968);
    layer2_outputs(8017) <= not(layer1_outputs(636));
    layer2_outputs(8018) <= not(layer1_outputs(3160)) or (layer1_outputs(5569));
    layer2_outputs(8019) <= '0';
    layer2_outputs(8020) <= (layer1_outputs(4691)) and not (layer1_outputs(1257));
    layer2_outputs(8021) <= not(layer1_outputs(9350));
    layer2_outputs(8022) <= layer1_outputs(2556);
    layer2_outputs(8023) <= not((layer1_outputs(1576)) and (layer1_outputs(4775)));
    layer2_outputs(8024) <= not(layer1_outputs(6880));
    layer2_outputs(8025) <= (layer1_outputs(8942)) and not (layer1_outputs(4802));
    layer2_outputs(8026) <= not((layer1_outputs(2492)) or (layer1_outputs(5114)));
    layer2_outputs(8027) <= not((layer1_outputs(9403)) or (layer1_outputs(977)));
    layer2_outputs(8028) <= (layer1_outputs(1289)) and not (layer1_outputs(9565));
    layer2_outputs(8029) <= not((layer1_outputs(3143)) and (layer1_outputs(2067)));
    layer2_outputs(8030) <= '1';
    layer2_outputs(8031) <= (layer1_outputs(9806)) and (layer1_outputs(9936));
    layer2_outputs(8032) <= layer1_outputs(9229);
    layer2_outputs(8033) <= (layer1_outputs(7925)) xor (layer1_outputs(9008));
    layer2_outputs(8034) <= not(layer1_outputs(7136));
    layer2_outputs(8035) <= (layer1_outputs(4958)) and not (layer1_outputs(2405));
    layer2_outputs(8036) <= not(layer1_outputs(8610));
    layer2_outputs(8037) <= layer1_outputs(9804);
    layer2_outputs(8038) <= '1';
    layer2_outputs(8039) <= not(layer1_outputs(1706)) or (layer1_outputs(7176));
    layer2_outputs(8040) <= not((layer1_outputs(3444)) or (layer1_outputs(1422)));
    layer2_outputs(8041) <= not(layer1_outputs(6095)) or (layer1_outputs(752));
    layer2_outputs(8042) <= layer1_outputs(2595);
    layer2_outputs(8043) <= layer1_outputs(1139);
    layer2_outputs(8044) <= not(layer1_outputs(5929)) or (layer1_outputs(6227));
    layer2_outputs(8045) <= not(layer1_outputs(1655)) or (layer1_outputs(3266));
    layer2_outputs(8046) <= not(layer1_outputs(1822));
    layer2_outputs(8047) <= (layer1_outputs(5065)) xor (layer1_outputs(9832));
    layer2_outputs(8048) <= not(layer1_outputs(10148));
    layer2_outputs(8049) <= (layer1_outputs(8192)) or (layer1_outputs(128));
    layer2_outputs(8050) <= not(layer1_outputs(136)) or (layer1_outputs(8051));
    layer2_outputs(8051) <= not((layer1_outputs(974)) xor (layer1_outputs(5347)));
    layer2_outputs(8052) <= layer1_outputs(7664);
    layer2_outputs(8053) <= layer1_outputs(8025);
    layer2_outputs(8054) <= not(layer1_outputs(6233));
    layer2_outputs(8055) <= not(layer1_outputs(4930)) or (layer1_outputs(2467));
    layer2_outputs(8056) <= layer1_outputs(2314);
    layer2_outputs(8057) <= layer1_outputs(8254);
    layer2_outputs(8058) <= layer1_outputs(183);
    layer2_outputs(8059) <= layer1_outputs(5390);
    layer2_outputs(8060) <= layer1_outputs(5485);
    layer2_outputs(8061) <= not(layer1_outputs(8606)) or (layer1_outputs(2154));
    layer2_outputs(8062) <= not(layer1_outputs(810));
    layer2_outputs(8063) <= layer1_outputs(142);
    layer2_outputs(8064) <= not(layer1_outputs(9490));
    layer2_outputs(8065) <= not(layer1_outputs(5173)) or (layer1_outputs(1320));
    layer2_outputs(8066) <= not(layer1_outputs(3784));
    layer2_outputs(8067) <= (layer1_outputs(8855)) and (layer1_outputs(7591));
    layer2_outputs(8068) <= not(layer1_outputs(4742));
    layer2_outputs(8069) <= not(layer1_outputs(9195)) or (layer1_outputs(863));
    layer2_outputs(8070) <= layer1_outputs(4362);
    layer2_outputs(8071) <= not((layer1_outputs(4845)) or (layer1_outputs(4549)));
    layer2_outputs(8072) <= not(layer1_outputs(6311));
    layer2_outputs(8073) <= (layer1_outputs(5364)) and (layer1_outputs(1506));
    layer2_outputs(8074) <= layer1_outputs(8184);
    layer2_outputs(8075) <= not((layer1_outputs(9667)) or (layer1_outputs(948)));
    layer2_outputs(8076) <= not((layer1_outputs(3525)) or (layer1_outputs(9734)));
    layer2_outputs(8077) <= not((layer1_outputs(3666)) and (layer1_outputs(6556)));
    layer2_outputs(8078) <= not(layer1_outputs(107)) or (layer1_outputs(8461));
    layer2_outputs(8079) <= not(layer1_outputs(7012));
    layer2_outputs(8080) <= (layer1_outputs(6604)) or (layer1_outputs(7376));
    layer2_outputs(8081) <= (layer1_outputs(278)) and (layer1_outputs(7381));
    layer2_outputs(8082) <= layer1_outputs(1997);
    layer2_outputs(8083) <= not(layer1_outputs(7043));
    layer2_outputs(8084) <= (layer1_outputs(7394)) and (layer1_outputs(4016));
    layer2_outputs(8085) <= (layer1_outputs(2551)) or (layer1_outputs(4153));
    layer2_outputs(8086) <= not(layer1_outputs(4073));
    layer2_outputs(8087) <= (layer1_outputs(776)) and not (layer1_outputs(8256));
    layer2_outputs(8088) <= not(layer1_outputs(4603));
    layer2_outputs(8089) <= layer1_outputs(8139);
    layer2_outputs(8090) <= (layer1_outputs(6166)) and not (layer1_outputs(4427));
    layer2_outputs(8091) <= not((layer1_outputs(7726)) or (layer1_outputs(9876)));
    layer2_outputs(8092) <= not(layer1_outputs(8614));
    layer2_outputs(8093) <= not(layer1_outputs(6003));
    layer2_outputs(8094) <= (layer1_outputs(3956)) and (layer1_outputs(7621));
    layer2_outputs(8095) <= layer1_outputs(6838);
    layer2_outputs(8096) <= '1';
    layer2_outputs(8097) <= (layer1_outputs(1774)) and not (layer1_outputs(6255));
    layer2_outputs(8098) <= (layer1_outputs(184)) and not (layer1_outputs(8017));
    layer2_outputs(8099) <= (layer1_outputs(2321)) and (layer1_outputs(9336));
    layer2_outputs(8100) <= not(layer1_outputs(1156));
    layer2_outputs(8101) <= (layer1_outputs(7902)) and not (layer1_outputs(5430));
    layer2_outputs(8102) <= not((layer1_outputs(5516)) xor (layer1_outputs(10055)));
    layer2_outputs(8103) <= not(layer1_outputs(6786)) or (layer1_outputs(931));
    layer2_outputs(8104) <= (layer1_outputs(1451)) or (layer1_outputs(268));
    layer2_outputs(8105) <= '0';
    layer2_outputs(8106) <= not(layer1_outputs(5477)) or (layer1_outputs(717));
    layer2_outputs(8107) <= layer1_outputs(6039);
    layer2_outputs(8108) <= not(layer1_outputs(10160));
    layer2_outputs(8109) <= (layer1_outputs(9056)) and (layer1_outputs(5339));
    layer2_outputs(8110) <= not((layer1_outputs(5643)) xor (layer1_outputs(462)));
    layer2_outputs(8111) <= layer1_outputs(8297);
    layer2_outputs(8112) <= not((layer1_outputs(4170)) or (layer1_outputs(2420)));
    layer2_outputs(8113) <= (layer1_outputs(10161)) and not (layer1_outputs(6675));
    layer2_outputs(8114) <= not((layer1_outputs(4831)) and (layer1_outputs(8326)));
    layer2_outputs(8115) <= not((layer1_outputs(2323)) xor (layer1_outputs(6680)));
    layer2_outputs(8116) <= not((layer1_outputs(3295)) and (layer1_outputs(9140)));
    layer2_outputs(8117) <= not((layer1_outputs(7481)) or (layer1_outputs(4698)));
    layer2_outputs(8118) <= not(layer1_outputs(8296)) or (layer1_outputs(9496));
    layer2_outputs(8119) <= (layer1_outputs(9156)) or (layer1_outputs(7358));
    layer2_outputs(8120) <= not(layer1_outputs(5937));
    layer2_outputs(8121) <= not((layer1_outputs(2472)) or (layer1_outputs(1201)));
    layer2_outputs(8122) <= '0';
    layer2_outputs(8123) <= not(layer1_outputs(2484));
    layer2_outputs(8124) <= layer1_outputs(2254);
    layer2_outputs(8125) <= layer1_outputs(4754);
    layer2_outputs(8126) <= layer1_outputs(1840);
    layer2_outputs(8127) <= not(layer1_outputs(7279));
    layer2_outputs(8128) <= not(layer1_outputs(5055));
    layer2_outputs(8129) <= not(layer1_outputs(7414));
    layer2_outputs(8130) <= layer1_outputs(4219);
    layer2_outputs(8131) <= (layer1_outputs(843)) and not (layer1_outputs(5695));
    layer2_outputs(8132) <= layer1_outputs(7179);
    layer2_outputs(8133) <= layer1_outputs(7891);
    layer2_outputs(8134) <= '0';
    layer2_outputs(8135) <= not((layer1_outputs(3801)) or (layer1_outputs(6695)));
    layer2_outputs(8136) <= layer1_outputs(323);
    layer2_outputs(8137) <= (layer1_outputs(8278)) and not (layer1_outputs(5083));
    layer2_outputs(8138) <= '0';
    layer2_outputs(8139) <= not(layer1_outputs(5265));
    layer2_outputs(8140) <= (layer1_outputs(6955)) and (layer1_outputs(4704));
    layer2_outputs(8141) <= (layer1_outputs(6419)) or (layer1_outputs(1936));
    layer2_outputs(8142) <= not(layer1_outputs(4972));
    layer2_outputs(8143) <= not(layer1_outputs(8011)) or (layer1_outputs(2884));
    layer2_outputs(8144) <= not(layer1_outputs(16));
    layer2_outputs(8145) <= not(layer1_outputs(8076));
    layer2_outputs(8146) <= layer1_outputs(539);
    layer2_outputs(8147) <= (layer1_outputs(757)) and not (layer1_outputs(10204));
    layer2_outputs(8148) <= not((layer1_outputs(7515)) or (layer1_outputs(8037)));
    layer2_outputs(8149) <= layer1_outputs(1280);
    layer2_outputs(8150) <= not(layer1_outputs(8718)) or (layer1_outputs(7526));
    layer2_outputs(8151) <= (layer1_outputs(1555)) and not (layer1_outputs(10098));
    layer2_outputs(8152) <= not(layer1_outputs(1098));
    layer2_outputs(8153) <= (layer1_outputs(4961)) and (layer1_outputs(4721));
    layer2_outputs(8154) <= layer1_outputs(9199);
    layer2_outputs(8155) <= layer1_outputs(7705);
    layer2_outputs(8156) <= not((layer1_outputs(6652)) or (layer1_outputs(1870)));
    layer2_outputs(8157) <= (layer1_outputs(5981)) and not (layer1_outputs(7059));
    layer2_outputs(8158) <= layer1_outputs(7625);
    layer2_outputs(8159) <= '1';
    layer2_outputs(8160) <= not(layer1_outputs(7231));
    layer2_outputs(8161) <= (layer1_outputs(2430)) and not (layer1_outputs(8002));
    layer2_outputs(8162) <= layer1_outputs(532);
    layer2_outputs(8163) <= '0';
    layer2_outputs(8164) <= not(layer1_outputs(4318));
    layer2_outputs(8165) <= (layer1_outputs(5751)) xor (layer1_outputs(2604));
    layer2_outputs(8166) <= not(layer1_outputs(9589));
    layer2_outputs(8167) <= (layer1_outputs(9474)) or (layer1_outputs(8922));
    layer2_outputs(8168) <= not((layer1_outputs(1514)) or (layer1_outputs(2598)));
    layer2_outputs(8169) <= (layer1_outputs(9928)) or (layer1_outputs(4631));
    layer2_outputs(8170) <= not(layer1_outputs(7225));
    layer2_outputs(8171) <= (layer1_outputs(8002)) or (layer1_outputs(5220));
    layer2_outputs(8172) <= not(layer1_outputs(8866));
    layer2_outputs(8173) <= layer1_outputs(1732);
    layer2_outputs(8174) <= (layer1_outputs(6515)) and (layer1_outputs(9664));
    layer2_outputs(8175) <= not(layer1_outputs(4549));
    layer2_outputs(8176) <= (layer1_outputs(3311)) and not (layer1_outputs(6441));
    layer2_outputs(8177) <= '0';
    layer2_outputs(8178) <= not(layer1_outputs(9778)) or (layer1_outputs(2313));
    layer2_outputs(8179) <= not((layer1_outputs(9362)) or (layer1_outputs(6894)));
    layer2_outputs(8180) <= '1';
    layer2_outputs(8181) <= not((layer1_outputs(7002)) xor (layer1_outputs(4205)));
    layer2_outputs(8182) <= layer1_outputs(2896);
    layer2_outputs(8183) <= not((layer1_outputs(6913)) xor (layer1_outputs(3437)));
    layer2_outputs(8184) <= (layer1_outputs(6277)) or (layer1_outputs(5449));
    layer2_outputs(8185) <= layer1_outputs(753);
    layer2_outputs(8186) <= (layer1_outputs(3934)) and not (layer1_outputs(9550));
    layer2_outputs(8187) <= not(layer1_outputs(6557));
    layer2_outputs(8188) <= (layer1_outputs(6762)) or (layer1_outputs(564));
    layer2_outputs(8189) <= not(layer1_outputs(276));
    layer2_outputs(8190) <= not(layer1_outputs(8984));
    layer2_outputs(8191) <= layer1_outputs(8428);
    layer2_outputs(8192) <= not(layer1_outputs(6954));
    layer2_outputs(8193) <= (layer1_outputs(5029)) and (layer1_outputs(2458));
    layer2_outputs(8194) <= '1';
    layer2_outputs(8195) <= not(layer1_outputs(5668));
    layer2_outputs(8196) <= not((layer1_outputs(9610)) and (layer1_outputs(8048)));
    layer2_outputs(8197) <= (layer1_outputs(1768)) and not (layer1_outputs(7913));
    layer2_outputs(8198) <= (layer1_outputs(7305)) and (layer1_outputs(4455));
    layer2_outputs(8199) <= not((layer1_outputs(8273)) or (layer1_outputs(3070)));
    layer2_outputs(8200) <= '1';
    layer2_outputs(8201) <= (layer1_outputs(5956)) and not (layer1_outputs(651));
    layer2_outputs(8202) <= not(layer1_outputs(4121));
    layer2_outputs(8203) <= (layer1_outputs(5190)) and (layer1_outputs(3456));
    layer2_outputs(8204) <= not(layer1_outputs(1363)) or (layer1_outputs(5244));
    layer2_outputs(8205) <= (layer1_outputs(4453)) and (layer1_outputs(5528));
    layer2_outputs(8206) <= not(layer1_outputs(5893));
    layer2_outputs(8207) <= not(layer1_outputs(1954));
    layer2_outputs(8208) <= layer1_outputs(7018);
    layer2_outputs(8209) <= layer1_outputs(2198);
    layer2_outputs(8210) <= layer1_outputs(7609);
    layer2_outputs(8211) <= not(layer1_outputs(6664));
    layer2_outputs(8212) <= not(layer1_outputs(7576));
    layer2_outputs(8213) <= not(layer1_outputs(2737)) or (layer1_outputs(9700));
    layer2_outputs(8214) <= layer1_outputs(3533);
    layer2_outputs(8215) <= layer1_outputs(7539);
    layer2_outputs(8216) <= not(layer1_outputs(745));
    layer2_outputs(8217) <= not(layer1_outputs(4659));
    layer2_outputs(8218) <= (layer1_outputs(2533)) or (layer1_outputs(7362));
    layer2_outputs(8219) <= not(layer1_outputs(4515));
    layer2_outputs(8220) <= layer1_outputs(6507);
    layer2_outputs(8221) <= (layer1_outputs(8232)) and not (layer1_outputs(707));
    layer2_outputs(8222) <= not(layer1_outputs(2939));
    layer2_outputs(8223) <= (layer1_outputs(580)) and (layer1_outputs(7824));
    layer2_outputs(8224) <= not(layer1_outputs(4853));
    layer2_outputs(8225) <= '1';
    layer2_outputs(8226) <= (layer1_outputs(671)) or (layer1_outputs(187));
    layer2_outputs(8227) <= layer1_outputs(2165);
    layer2_outputs(8228) <= '0';
    layer2_outputs(8229) <= (layer1_outputs(1467)) or (layer1_outputs(1485));
    layer2_outputs(8230) <= (layer1_outputs(9453)) xor (layer1_outputs(2672));
    layer2_outputs(8231) <= (layer1_outputs(250)) and (layer1_outputs(10058));
    layer2_outputs(8232) <= not(layer1_outputs(1269)) or (layer1_outputs(8385));
    layer2_outputs(8233) <= (layer1_outputs(1587)) or (layer1_outputs(6173));
    layer2_outputs(8234) <= not(layer1_outputs(5743)) or (layer1_outputs(6340));
    layer2_outputs(8235) <= layer1_outputs(590);
    layer2_outputs(8236) <= layer1_outputs(387);
    layer2_outputs(8237) <= layer1_outputs(7147);
    layer2_outputs(8238) <= not((layer1_outputs(9446)) and (layer1_outputs(155)));
    layer2_outputs(8239) <= layer1_outputs(7472);
    layer2_outputs(8240) <= layer1_outputs(4062);
    layer2_outputs(8241) <= not(layer1_outputs(7389));
    layer2_outputs(8242) <= not(layer1_outputs(3953));
    layer2_outputs(8243) <= layer1_outputs(1787);
    layer2_outputs(8244) <= layer1_outputs(5426);
    layer2_outputs(8245) <= (layer1_outputs(9010)) and not (layer1_outputs(4208));
    layer2_outputs(8246) <= layer1_outputs(10060);
    layer2_outputs(8247) <= not(layer1_outputs(9745));
    layer2_outputs(8248) <= layer1_outputs(1052);
    layer2_outputs(8249) <= layer1_outputs(453);
    layer2_outputs(8250) <= not((layer1_outputs(5046)) and (layer1_outputs(2303)));
    layer2_outputs(8251) <= not((layer1_outputs(2607)) xor (layer1_outputs(2091)));
    layer2_outputs(8252) <= (layer1_outputs(5005)) and not (layer1_outputs(9836));
    layer2_outputs(8253) <= (layer1_outputs(104)) and (layer1_outputs(5911));
    layer2_outputs(8254) <= not((layer1_outputs(9240)) and (layer1_outputs(7756)));
    layer2_outputs(8255) <= (layer1_outputs(2676)) and (layer1_outputs(2866));
    layer2_outputs(8256) <= layer1_outputs(4395);
    layer2_outputs(8257) <= (layer1_outputs(5365)) and not (layer1_outputs(275));
    layer2_outputs(8258) <= not((layer1_outputs(1565)) and (layer1_outputs(2193)));
    layer2_outputs(8259) <= '0';
    layer2_outputs(8260) <= '1';
    layer2_outputs(8261) <= (layer1_outputs(786)) or (layer1_outputs(7152));
    layer2_outputs(8262) <= not(layer1_outputs(6963));
    layer2_outputs(8263) <= not(layer1_outputs(7215));
    layer2_outputs(8264) <= not(layer1_outputs(7584));
    layer2_outputs(8265) <= layer1_outputs(9395);
    layer2_outputs(8266) <= not(layer1_outputs(3663)) or (layer1_outputs(1199));
    layer2_outputs(8267) <= '0';
    layer2_outputs(8268) <= layer1_outputs(2956);
    layer2_outputs(8269) <= not(layer1_outputs(9187));
    layer2_outputs(8270) <= '1';
    layer2_outputs(8271) <= (layer1_outputs(4570)) and (layer1_outputs(9487));
    layer2_outputs(8272) <= not((layer1_outputs(9185)) and (layer1_outputs(9883)));
    layer2_outputs(8273) <= (layer1_outputs(2662)) or (layer1_outputs(904));
    layer2_outputs(8274) <= (layer1_outputs(2496)) and (layer1_outputs(3310));
    layer2_outputs(8275) <= layer1_outputs(6877);
    layer2_outputs(8276) <= not((layer1_outputs(3813)) and (layer1_outputs(1974)));
    layer2_outputs(8277) <= (layer1_outputs(575)) and (layer1_outputs(7527));
    layer2_outputs(8278) <= not(layer1_outputs(8863)) or (layer1_outputs(7098));
    layer2_outputs(8279) <= '0';
    layer2_outputs(8280) <= not(layer1_outputs(3997));
    layer2_outputs(8281) <= (layer1_outputs(9197)) and not (layer1_outputs(2909));
    layer2_outputs(8282) <= (layer1_outputs(5657)) and not (layer1_outputs(311));
    layer2_outputs(8283) <= (layer1_outputs(4152)) and not (layer1_outputs(1812));
    layer2_outputs(8284) <= not(layer1_outputs(3009));
    layer2_outputs(8285) <= layer1_outputs(8621);
    layer2_outputs(8286) <= layer1_outputs(1747);
    layer2_outputs(8287) <= layer1_outputs(9347);
    layer2_outputs(8288) <= not(layer1_outputs(949)) or (layer1_outputs(1844));
    layer2_outputs(8289) <= layer1_outputs(3717);
    layer2_outputs(8290) <= layer1_outputs(6744);
    layer2_outputs(8291) <= not(layer1_outputs(3215));
    layer2_outputs(8292) <= not((layer1_outputs(973)) and (layer1_outputs(9049)));
    layer2_outputs(8293) <= layer1_outputs(9389);
    layer2_outputs(8294) <= not(layer1_outputs(3967));
    layer2_outputs(8295) <= not(layer1_outputs(755));
    layer2_outputs(8296) <= not(layer1_outputs(9237));
    layer2_outputs(8297) <= not((layer1_outputs(4116)) xor (layer1_outputs(1407)));
    layer2_outputs(8298) <= not(layer1_outputs(403));
    layer2_outputs(8299) <= (layer1_outputs(6495)) and not (layer1_outputs(7835));
    layer2_outputs(8300) <= (layer1_outputs(6953)) and not (layer1_outputs(304));
    layer2_outputs(8301) <= layer1_outputs(4679);
    layer2_outputs(8302) <= not(layer1_outputs(8071));
    layer2_outputs(8303) <= not(layer1_outputs(5735));
    layer2_outputs(8304) <= not(layer1_outputs(7227));
    layer2_outputs(8305) <= not(layer1_outputs(9955));
    layer2_outputs(8306) <= not(layer1_outputs(4873));
    layer2_outputs(8307) <= not(layer1_outputs(2306));
    layer2_outputs(8308) <= layer1_outputs(7969);
    layer2_outputs(8309) <= (layer1_outputs(2616)) or (layer1_outputs(7295));
    layer2_outputs(8310) <= not(layer1_outputs(5033));
    layer2_outputs(8311) <= not(layer1_outputs(8702)) or (layer1_outputs(5171));
    layer2_outputs(8312) <= not(layer1_outputs(7731));
    layer2_outputs(8313) <= (layer1_outputs(3290)) xor (layer1_outputs(756));
    layer2_outputs(8314) <= (layer1_outputs(1981)) and not (layer1_outputs(9511));
    layer2_outputs(8315) <= not((layer1_outputs(8885)) xor (layer1_outputs(7545)));
    layer2_outputs(8316) <= not((layer1_outputs(3861)) or (layer1_outputs(7821)));
    layer2_outputs(8317) <= not(layer1_outputs(465));
    layer2_outputs(8318) <= layer1_outputs(6573);
    layer2_outputs(8319) <= '1';
    layer2_outputs(8320) <= not(layer1_outputs(2875));
    layer2_outputs(8321) <= not(layer1_outputs(7431));
    layer2_outputs(8322) <= not((layer1_outputs(3033)) and (layer1_outputs(659)));
    layer2_outputs(8323) <= not(layer1_outputs(8955)) or (layer1_outputs(9263));
    layer2_outputs(8324) <= layer1_outputs(4057);
    layer2_outputs(8325) <= not((layer1_outputs(2870)) or (layer1_outputs(9352)));
    layer2_outputs(8326) <= not(layer1_outputs(4618)) or (layer1_outputs(7923));
    layer2_outputs(8327) <= layer1_outputs(4679);
    layer2_outputs(8328) <= not((layer1_outputs(8850)) and (layer1_outputs(6124)));
    layer2_outputs(8329) <= not(layer1_outputs(3125)) or (layer1_outputs(9147));
    layer2_outputs(8330) <= layer1_outputs(9279);
    layer2_outputs(8331) <= not((layer1_outputs(1671)) xor (layer1_outputs(5186)));
    layer2_outputs(8332) <= not(layer1_outputs(2798)) or (layer1_outputs(293));
    layer2_outputs(8333) <= not(layer1_outputs(1424));
    layer2_outputs(8334) <= (layer1_outputs(419)) xor (layer1_outputs(1962));
    layer2_outputs(8335) <= (layer1_outputs(4234)) and not (layer1_outputs(2285));
    layer2_outputs(8336) <= layer1_outputs(1033);
    layer2_outputs(8337) <= (layer1_outputs(8420)) and (layer1_outputs(4015));
    layer2_outputs(8338) <= (layer1_outputs(8759)) or (layer1_outputs(5281));
    layer2_outputs(8339) <= (layer1_outputs(865)) and (layer1_outputs(2496));
    layer2_outputs(8340) <= layer1_outputs(2103);
    layer2_outputs(8341) <= (layer1_outputs(2680)) and (layer1_outputs(4177));
    layer2_outputs(8342) <= not(layer1_outputs(2497));
    layer2_outputs(8343) <= (layer1_outputs(7634)) and not (layer1_outputs(3137));
    layer2_outputs(8344) <= not((layer1_outputs(210)) xor (layer1_outputs(9003)));
    layer2_outputs(8345) <= not((layer1_outputs(3805)) and (layer1_outputs(858)));
    layer2_outputs(8346) <= not(layer1_outputs(3600));
    layer2_outputs(8347) <= '1';
    layer2_outputs(8348) <= '1';
    layer2_outputs(8349) <= (layer1_outputs(4297)) and not (layer1_outputs(37));
    layer2_outputs(8350) <= not(layer1_outputs(2680));
    layer2_outputs(8351) <= not(layer1_outputs(4465));
    layer2_outputs(8352) <= not(layer1_outputs(9496));
    layer2_outputs(8353) <= (layer1_outputs(1615)) and not (layer1_outputs(7971));
    layer2_outputs(8354) <= (layer1_outputs(10125)) and not (layer1_outputs(2840));
    layer2_outputs(8355) <= (layer1_outputs(2193)) or (layer1_outputs(2539));
    layer2_outputs(8356) <= (layer1_outputs(8764)) and (layer1_outputs(2709));
    layer2_outputs(8357) <= layer1_outputs(3987);
    layer2_outputs(8358) <= not(layer1_outputs(5174));
    layer2_outputs(8359) <= (layer1_outputs(8020)) or (layer1_outputs(6400));
    layer2_outputs(8360) <= not(layer1_outputs(4044)) or (layer1_outputs(2673));
    layer2_outputs(8361) <= not(layer1_outputs(9931)) or (layer1_outputs(3465));
    layer2_outputs(8362) <= not((layer1_outputs(4182)) xor (layer1_outputs(8831)));
    layer2_outputs(8363) <= (layer1_outputs(1871)) or (layer1_outputs(10004));
    layer2_outputs(8364) <= not(layer1_outputs(7421)) or (layer1_outputs(9180));
    layer2_outputs(8365) <= not(layer1_outputs(7229));
    layer2_outputs(8366) <= not((layer1_outputs(5756)) and (layer1_outputs(4640)));
    layer2_outputs(8367) <= layer1_outputs(1879);
    layer2_outputs(8368) <= not(layer1_outputs(9594));
    layer2_outputs(8369) <= layer1_outputs(2280);
    layer2_outputs(8370) <= (layer1_outputs(6817)) and not (layer1_outputs(10188));
    layer2_outputs(8371) <= not((layer1_outputs(2583)) and (layer1_outputs(5789)));
    layer2_outputs(8372) <= layer1_outputs(5577);
    layer2_outputs(8373) <= '1';
    layer2_outputs(8374) <= not(layer1_outputs(1175));
    layer2_outputs(8375) <= layer1_outputs(2161);
    layer2_outputs(8376) <= layer1_outputs(5785);
    layer2_outputs(8377) <= (layer1_outputs(9452)) or (layer1_outputs(4475));
    layer2_outputs(8378) <= (layer1_outputs(5153)) and (layer1_outputs(5123));
    layer2_outputs(8379) <= layer1_outputs(10145);
    layer2_outputs(8380) <= not((layer1_outputs(4726)) xor (layer1_outputs(7397)));
    layer2_outputs(8381) <= (layer1_outputs(9029)) or (layer1_outputs(1331));
    layer2_outputs(8382) <= not((layer1_outputs(9562)) xor (layer1_outputs(925)));
    layer2_outputs(8383) <= layer1_outputs(3192);
    layer2_outputs(8384) <= (layer1_outputs(7462)) or (layer1_outputs(8196));
    layer2_outputs(8385) <= layer1_outputs(5386);
    layer2_outputs(8386) <= not(layer1_outputs(7032));
    layer2_outputs(8387) <= not(layer1_outputs(8926)) or (layer1_outputs(2603));
    layer2_outputs(8388) <= (layer1_outputs(9484)) and not (layer1_outputs(6148));
    layer2_outputs(8389) <= (layer1_outputs(3499)) and (layer1_outputs(4036));
    layer2_outputs(8390) <= (layer1_outputs(1501)) xor (layer1_outputs(6174));
    layer2_outputs(8391) <= '1';
    layer2_outputs(8392) <= not(layer1_outputs(9929)) or (layer1_outputs(9055));
    layer2_outputs(8393) <= not((layer1_outputs(5771)) or (layer1_outputs(5807)));
    layer2_outputs(8394) <= not(layer1_outputs(1029));
    layer2_outputs(8395) <= (layer1_outputs(5447)) or (layer1_outputs(3723));
    layer2_outputs(8396) <= '1';
    layer2_outputs(8397) <= '0';
    layer2_outputs(8398) <= (layer1_outputs(4469)) and not (layer1_outputs(6153));
    layer2_outputs(8399) <= not(layer1_outputs(7138)) or (layer1_outputs(4625));
    layer2_outputs(8400) <= not((layer1_outputs(6165)) or (layer1_outputs(7861)));
    layer2_outputs(8401) <= not((layer1_outputs(1255)) and (layer1_outputs(3940)));
    layer2_outputs(8402) <= (layer1_outputs(7798)) and not (layer1_outputs(3534));
    layer2_outputs(8403) <= not((layer1_outputs(5576)) and (layer1_outputs(6010)));
    layer2_outputs(8404) <= '0';
    layer2_outputs(8405) <= not(layer1_outputs(8831)) or (layer1_outputs(583));
    layer2_outputs(8406) <= '0';
    layer2_outputs(8407) <= not(layer1_outputs(7009)) or (layer1_outputs(783));
    layer2_outputs(8408) <= '0';
    layer2_outputs(8409) <= not((layer1_outputs(2558)) or (layer1_outputs(3910)));
    layer2_outputs(8410) <= '0';
    layer2_outputs(8411) <= '1';
    layer2_outputs(8412) <= layer1_outputs(9146);
    layer2_outputs(8413) <= '1';
    layer2_outputs(8414) <= (layer1_outputs(837)) or (layer1_outputs(7235));
    layer2_outputs(8415) <= layer1_outputs(3441);
    layer2_outputs(8416) <= '0';
    layer2_outputs(8417) <= not(layer1_outputs(7969));
    layer2_outputs(8418) <= layer1_outputs(10196);
    layer2_outputs(8419) <= not((layer1_outputs(3178)) or (layer1_outputs(3565)));
    layer2_outputs(8420) <= (layer1_outputs(9875)) or (layer1_outputs(40));
    layer2_outputs(8421) <= (layer1_outputs(3738)) and not (layer1_outputs(5176));
    layer2_outputs(8422) <= (layer1_outputs(5314)) or (layer1_outputs(4709));
    layer2_outputs(8423) <= layer1_outputs(2366);
    layer2_outputs(8424) <= layer1_outputs(3507);
    layer2_outputs(8425) <= (layer1_outputs(6584)) and not (layer1_outputs(8786));
    layer2_outputs(8426) <= not((layer1_outputs(2981)) and (layer1_outputs(8238)));
    layer2_outputs(8427) <= not(layer1_outputs(8530));
    layer2_outputs(8428) <= not(layer1_outputs(6673)) or (layer1_outputs(4353));
    layer2_outputs(8429) <= not(layer1_outputs(127));
    layer2_outputs(8430) <= layer1_outputs(1668);
    layer2_outputs(8431) <= not(layer1_outputs(960));
    layer2_outputs(8432) <= (layer1_outputs(9374)) or (layer1_outputs(4946));
    layer2_outputs(8433) <= layer1_outputs(6052);
    layer2_outputs(8434) <= not(layer1_outputs(3377)) or (layer1_outputs(7081));
    layer2_outputs(8435) <= (layer1_outputs(10097)) and not (layer1_outputs(2881));
    layer2_outputs(8436) <= (layer1_outputs(845)) or (layer1_outputs(8364));
    layer2_outputs(8437) <= not((layer1_outputs(985)) or (layer1_outputs(9205)));
    layer2_outputs(8438) <= (layer1_outputs(2391)) or (layer1_outputs(4401));
    layer2_outputs(8439) <= not(layer1_outputs(7070));
    layer2_outputs(8440) <= (layer1_outputs(1801)) or (layer1_outputs(4282));
    layer2_outputs(8441) <= (layer1_outputs(6991)) xor (layer1_outputs(8758));
    layer2_outputs(8442) <= not((layer1_outputs(8822)) or (layer1_outputs(9032)));
    layer2_outputs(8443) <= not((layer1_outputs(1364)) or (layer1_outputs(491)));
    layer2_outputs(8444) <= not((layer1_outputs(2773)) and (layer1_outputs(724)));
    layer2_outputs(8445) <= not(layer1_outputs(1697));
    layer2_outputs(8446) <= (layer1_outputs(2859)) and not (layer1_outputs(7352));
    layer2_outputs(8447) <= layer1_outputs(5268);
    layer2_outputs(8448) <= (layer1_outputs(3905)) and (layer1_outputs(9545));
    layer2_outputs(8449) <= (layer1_outputs(2813)) or (layer1_outputs(1703));
    layer2_outputs(8450) <= not(layer1_outputs(2800));
    layer2_outputs(8451) <= not(layer1_outputs(3183)) or (layer1_outputs(3788));
    layer2_outputs(8452) <= (layer1_outputs(2406)) and not (layer1_outputs(6038));
    layer2_outputs(8453) <= (layer1_outputs(3491)) and (layer1_outputs(4953));
    layer2_outputs(8454) <= not(layer1_outputs(3916));
    layer2_outputs(8455) <= (layer1_outputs(1584)) and not (layer1_outputs(3300));
    layer2_outputs(8456) <= not(layer1_outputs(596));
    layer2_outputs(8457) <= (layer1_outputs(5654)) and not (layer1_outputs(4140));
    layer2_outputs(8458) <= not(layer1_outputs(7646)) or (layer1_outputs(10205));
    layer2_outputs(8459) <= not((layer1_outputs(9425)) xor (layer1_outputs(676)));
    layer2_outputs(8460) <= not((layer1_outputs(3252)) xor (layer1_outputs(3068)));
    layer2_outputs(8461) <= (layer1_outputs(1891)) and not (layer1_outputs(940));
    layer2_outputs(8462) <= not(layer1_outputs(4664)) or (layer1_outputs(365));
    layer2_outputs(8463) <= (layer1_outputs(3014)) and not (layer1_outputs(3738));
    layer2_outputs(8464) <= layer1_outputs(50);
    layer2_outputs(8465) <= (layer1_outputs(9759)) and not (layer1_outputs(9620));
    layer2_outputs(8466) <= not((layer1_outputs(343)) or (layer1_outputs(2247)));
    layer2_outputs(8467) <= not((layer1_outputs(2351)) and (layer1_outputs(2232)));
    layer2_outputs(8468) <= layer1_outputs(480);
    layer2_outputs(8469) <= not(layer1_outputs(2260));
    layer2_outputs(8470) <= not(layer1_outputs(8972)) or (layer1_outputs(1131));
    layer2_outputs(8471) <= layer1_outputs(7008);
    layer2_outputs(8472) <= not(layer1_outputs(5919));
    layer2_outputs(8473) <= not((layer1_outputs(9745)) or (layer1_outputs(7945)));
    layer2_outputs(8474) <= layer1_outputs(9076);
    layer2_outputs(8475) <= (layer1_outputs(9121)) and not (layer1_outputs(6636));
    layer2_outputs(8476) <= not(layer1_outputs(8310));
    layer2_outputs(8477) <= not((layer1_outputs(5509)) and (layer1_outputs(1013)));
    layer2_outputs(8478) <= not(layer1_outputs(8366));
    layer2_outputs(8479) <= layer1_outputs(4034);
    layer2_outputs(8480) <= layer1_outputs(831);
    layer2_outputs(8481) <= not(layer1_outputs(7061));
    layer2_outputs(8482) <= layer1_outputs(3789);
    layer2_outputs(8483) <= not(layer1_outputs(4383));
    layer2_outputs(8484) <= not(layer1_outputs(793));
    layer2_outputs(8485) <= (layer1_outputs(3325)) xor (layer1_outputs(4773));
    layer2_outputs(8486) <= not(layer1_outputs(9100));
    layer2_outputs(8487) <= '0';
    layer2_outputs(8488) <= layer1_outputs(8657);
    layer2_outputs(8489) <= not(layer1_outputs(3715));
    layer2_outputs(8490) <= '0';
    layer2_outputs(8491) <= (layer1_outputs(8127)) and not (layer1_outputs(3976));
    layer2_outputs(8492) <= not(layer1_outputs(1841));
    layer2_outputs(8493) <= not(layer1_outputs(9307));
    layer2_outputs(8494) <= not(layer1_outputs(8589));
    layer2_outputs(8495) <= layer1_outputs(1175);
    layer2_outputs(8496) <= not(layer1_outputs(3939));
    layer2_outputs(8497) <= layer1_outputs(1739);
    layer2_outputs(8498) <= (layer1_outputs(3293)) and not (layer1_outputs(9069));
    layer2_outputs(8499) <= (layer1_outputs(8140)) and (layer1_outputs(569));
    layer2_outputs(8500) <= not((layer1_outputs(9381)) xor (layer1_outputs(1114)));
    layer2_outputs(8501) <= (layer1_outputs(9953)) and not (layer1_outputs(5793));
    layer2_outputs(8502) <= (layer1_outputs(4834)) and not (layer1_outputs(6008));
    layer2_outputs(8503) <= not(layer1_outputs(9485));
    layer2_outputs(8504) <= layer1_outputs(5455);
    layer2_outputs(8505) <= not(layer1_outputs(4831)) or (layer1_outputs(3306));
    layer2_outputs(8506) <= '0';
    layer2_outputs(8507) <= not(layer1_outputs(2371)) or (layer1_outputs(1966));
    layer2_outputs(8508) <= not((layer1_outputs(10154)) or (layer1_outputs(8710)));
    layer2_outputs(8509) <= not(layer1_outputs(4185)) or (layer1_outputs(615));
    layer2_outputs(8510) <= (layer1_outputs(7641)) and (layer1_outputs(4623));
    layer2_outputs(8511) <= layer1_outputs(4220);
    layer2_outputs(8512) <= (layer1_outputs(2025)) xor (layer1_outputs(7198));
    layer2_outputs(8513) <= (layer1_outputs(2633)) and not (layer1_outputs(9826));
    layer2_outputs(8514) <= not(layer1_outputs(8523));
    layer2_outputs(8515) <= not(layer1_outputs(988));
    layer2_outputs(8516) <= (layer1_outputs(8619)) and (layer1_outputs(9310));
    layer2_outputs(8517) <= layer1_outputs(4064);
    layer2_outputs(8518) <= layer1_outputs(9186);
    layer2_outputs(8519) <= not(layer1_outputs(1024));
    layer2_outputs(8520) <= not(layer1_outputs(2835));
    layer2_outputs(8521) <= not((layer1_outputs(292)) or (layer1_outputs(6363)));
    layer2_outputs(8522) <= not((layer1_outputs(6459)) or (layer1_outputs(6214)));
    layer2_outputs(8523) <= not(layer1_outputs(3347)) or (layer1_outputs(2514));
    layer2_outputs(8524) <= not(layer1_outputs(4206));
    layer2_outputs(8525) <= (layer1_outputs(10042)) and not (layer1_outputs(1531));
    layer2_outputs(8526) <= (layer1_outputs(9475)) and not (layer1_outputs(2715));
    layer2_outputs(8527) <= (layer1_outputs(4988)) or (layer1_outputs(7922));
    layer2_outputs(8528) <= not((layer1_outputs(9862)) and (layer1_outputs(3891)));
    layer2_outputs(8529) <= not(layer1_outputs(321)) or (layer1_outputs(971));
    layer2_outputs(8530) <= not(layer1_outputs(6509));
    layer2_outputs(8531) <= (layer1_outputs(8338)) and (layer1_outputs(1215));
    layer2_outputs(8532) <= not(layer1_outputs(6089)) or (layer1_outputs(4886));
    layer2_outputs(8533) <= not(layer1_outputs(4392));
    layer2_outputs(8534) <= not(layer1_outputs(9959));
    layer2_outputs(8535) <= layer1_outputs(2685);
    layer2_outputs(8536) <= '1';
    layer2_outputs(8537) <= (layer1_outputs(7251)) and not (layer1_outputs(9005));
    layer2_outputs(8538) <= not(layer1_outputs(1278)) or (layer1_outputs(8578));
    layer2_outputs(8539) <= layer1_outputs(6025);
    layer2_outputs(8540) <= not(layer1_outputs(4160)) or (layer1_outputs(8660));
    layer2_outputs(8541) <= layer1_outputs(2825);
    layer2_outputs(8542) <= layer1_outputs(5584);
    layer2_outputs(8543) <= layer1_outputs(3603);
    layer2_outputs(8544) <= layer1_outputs(5077);
    layer2_outputs(8545) <= not(layer1_outputs(7893));
    layer2_outputs(8546) <= (layer1_outputs(3401)) xor (layer1_outputs(3096));
    layer2_outputs(8547) <= (layer1_outputs(7109)) and not (layer1_outputs(1055));
    layer2_outputs(8548) <= layer1_outputs(4358);
    layer2_outputs(8549) <= not((layer1_outputs(3782)) or (layer1_outputs(104)));
    layer2_outputs(8550) <= layer1_outputs(8588);
    layer2_outputs(8551) <= not(layer1_outputs(3970));
    layer2_outputs(8552) <= layer1_outputs(5086);
    layer2_outputs(8553) <= layer1_outputs(2377);
    layer2_outputs(8554) <= not(layer1_outputs(7724));
    layer2_outputs(8555) <= (layer1_outputs(4589)) and (layer1_outputs(8858));
    layer2_outputs(8556) <= not((layer1_outputs(8011)) and (layer1_outputs(8789)));
    layer2_outputs(8557) <= not(layer1_outputs(8936));
    layer2_outputs(8558) <= layer1_outputs(4268);
    layer2_outputs(8559) <= layer1_outputs(9588);
    layer2_outputs(8560) <= '1';
    layer2_outputs(8561) <= (layer1_outputs(8771)) and not (layer1_outputs(1614));
    layer2_outputs(8562) <= not(layer1_outputs(5979));
    layer2_outputs(8563) <= (layer1_outputs(2601)) and not (layer1_outputs(7552));
    layer2_outputs(8564) <= not(layer1_outputs(6507));
    layer2_outputs(8565) <= (layer1_outputs(7407)) or (layer1_outputs(6487));
    layer2_outputs(8566) <= not(layer1_outputs(7380)) or (layer1_outputs(9889));
    layer2_outputs(8567) <= '0';
    layer2_outputs(8568) <= not((layer1_outputs(5433)) xor (layer1_outputs(351)));
    layer2_outputs(8569) <= not(layer1_outputs(6982));
    layer2_outputs(8570) <= (layer1_outputs(1097)) or (layer1_outputs(6699));
    layer2_outputs(8571) <= layer1_outputs(5319);
    layer2_outputs(8572) <= (layer1_outputs(8359)) or (layer1_outputs(10129));
    layer2_outputs(8573) <= not(layer1_outputs(7117));
    layer2_outputs(8574) <= (layer1_outputs(4770)) and not (layer1_outputs(4207));
    layer2_outputs(8575) <= not(layer1_outputs(5924));
    layer2_outputs(8576) <= not((layer1_outputs(3470)) and (layer1_outputs(3776)));
    layer2_outputs(8577) <= (layer1_outputs(8708)) or (layer1_outputs(6043));
    layer2_outputs(8578) <= layer1_outputs(7929);
    layer2_outputs(8579) <= layer1_outputs(8854);
    layer2_outputs(8580) <= (layer1_outputs(6862)) and not (layer1_outputs(7904));
    layer2_outputs(8581) <= layer1_outputs(6649);
    layer2_outputs(8582) <= not(layer1_outputs(4090));
    layer2_outputs(8583) <= not(layer1_outputs(541)) or (layer1_outputs(3761));
    layer2_outputs(8584) <= layer1_outputs(8856);
    layer2_outputs(8585) <= layer1_outputs(9610);
    layer2_outputs(8586) <= not((layer1_outputs(7578)) xor (layer1_outputs(1531)));
    layer2_outputs(8587) <= not(layer1_outputs(8793)) or (layer1_outputs(9711));
    layer2_outputs(8588) <= not(layer1_outputs(677));
    layer2_outputs(8589) <= layer1_outputs(6830);
    layer2_outputs(8590) <= not(layer1_outputs(3337));
    layer2_outputs(8591) <= layer1_outputs(3880);
    layer2_outputs(8592) <= not((layer1_outputs(4444)) or (layer1_outputs(6083)));
    layer2_outputs(8593) <= not(layer1_outputs(150));
    layer2_outputs(8594) <= (layer1_outputs(7637)) xor (layer1_outputs(3796));
    layer2_outputs(8595) <= (layer1_outputs(482)) and (layer1_outputs(8209));
    layer2_outputs(8596) <= (layer1_outputs(8309)) and not (layer1_outputs(3917));
    layer2_outputs(8597) <= (layer1_outputs(4616)) or (layer1_outputs(7128));
    layer2_outputs(8598) <= (layer1_outputs(3702)) or (layer1_outputs(4251));
    layer2_outputs(8599) <= not(layer1_outputs(5108));
    layer2_outputs(8600) <= not(layer1_outputs(373)) or (layer1_outputs(2571));
    layer2_outputs(8601) <= not(layer1_outputs(8298)) or (layer1_outputs(3359));
    layer2_outputs(8602) <= (layer1_outputs(4480)) and not (layer1_outputs(5500));
    layer2_outputs(8603) <= not(layer1_outputs(2399));
    layer2_outputs(8604) <= '1';
    layer2_outputs(8605) <= layer1_outputs(9527);
    layer2_outputs(8606) <= not(layer1_outputs(4641));
    layer2_outputs(8607) <= layer1_outputs(9979);
    layer2_outputs(8608) <= not(layer1_outputs(7045));
    layer2_outputs(8609) <= not((layer1_outputs(3665)) or (layer1_outputs(8907)));
    layer2_outputs(8610) <= (layer1_outputs(9836)) or (layer1_outputs(8211));
    layer2_outputs(8611) <= not((layer1_outputs(9792)) xor (layer1_outputs(7775)));
    layer2_outputs(8612) <= not(layer1_outputs(3224));
    layer2_outputs(8613) <= '1';
    layer2_outputs(8614) <= not(layer1_outputs(5985));
    layer2_outputs(8615) <= not(layer1_outputs(5530));
    layer2_outputs(8616) <= not(layer1_outputs(928)) or (layer1_outputs(6028));
    layer2_outputs(8617) <= layer1_outputs(9824);
    layer2_outputs(8618) <= not(layer1_outputs(10177));
    layer2_outputs(8619) <= not(layer1_outputs(1687)) or (layer1_outputs(2132));
    layer2_outputs(8620) <= (layer1_outputs(3331)) and not (layer1_outputs(3744));
    layer2_outputs(8621) <= (layer1_outputs(8580)) and not (layer1_outputs(838));
    layer2_outputs(8622) <= not((layer1_outputs(533)) and (layer1_outputs(6936)));
    layer2_outputs(8623) <= not(layer1_outputs(4238));
    layer2_outputs(8624) <= not((layer1_outputs(7758)) and (layer1_outputs(8329)));
    layer2_outputs(8625) <= (layer1_outputs(7175)) and not (layer1_outputs(3826));
    layer2_outputs(8626) <= '1';
    layer2_outputs(8627) <= (layer1_outputs(8715)) and not (layer1_outputs(6328));
    layer2_outputs(8628) <= (layer1_outputs(7616)) and not (layer1_outputs(6108));
    layer2_outputs(8629) <= not(layer1_outputs(735));
    layer2_outputs(8630) <= layer1_outputs(1708);
    layer2_outputs(8631) <= not((layer1_outputs(7080)) or (layer1_outputs(3174)));
    layer2_outputs(8632) <= layer1_outputs(1475);
    layer2_outputs(8633) <= not((layer1_outputs(9817)) xor (layer1_outputs(1502)));
    layer2_outputs(8634) <= not(layer1_outputs(3076));
    layer2_outputs(8635) <= not(layer1_outputs(9575));
    layer2_outputs(8636) <= not((layer1_outputs(7633)) or (layer1_outputs(836)));
    layer2_outputs(8637) <= (layer1_outputs(585)) and (layer1_outputs(3681));
    layer2_outputs(8638) <= not((layer1_outputs(4155)) and (layer1_outputs(9951)));
    layer2_outputs(8639) <= layer1_outputs(9147);
    layer2_outputs(8640) <= (layer1_outputs(457)) and (layer1_outputs(9691));
    layer2_outputs(8641) <= not((layer1_outputs(1620)) or (layer1_outputs(3502)));
    layer2_outputs(8642) <= not((layer1_outputs(9888)) or (layer1_outputs(5046)));
    layer2_outputs(8643) <= not(layer1_outputs(9605)) or (layer1_outputs(1702));
    layer2_outputs(8644) <= (layer1_outputs(817)) and not (layer1_outputs(9075));
    layer2_outputs(8645) <= '0';
    layer2_outputs(8646) <= not(layer1_outputs(6532));
    layer2_outputs(8647) <= (layer1_outputs(10239)) or (layer1_outputs(3357));
    layer2_outputs(8648) <= not((layer1_outputs(4387)) or (layer1_outputs(8085)));
    layer2_outputs(8649) <= (layer1_outputs(6669)) and not (layer1_outputs(1057));
    layer2_outputs(8650) <= layer1_outputs(8113);
    layer2_outputs(8651) <= not(layer1_outputs(1878));
    layer2_outputs(8652) <= not(layer1_outputs(4762));
    layer2_outputs(8653) <= (layer1_outputs(1186)) and (layer1_outputs(3646));
    layer2_outputs(8654) <= (layer1_outputs(3377)) and not (layer1_outputs(70));
    layer2_outputs(8655) <= not((layer1_outputs(4752)) and (layer1_outputs(1245)));
    layer2_outputs(8656) <= (layer1_outputs(8349)) and (layer1_outputs(4879));
    layer2_outputs(8657) <= not(layer1_outputs(2805));
    layer2_outputs(8658) <= '0';
    layer2_outputs(8659) <= not(layer1_outputs(10047));
    layer2_outputs(8660) <= not((layer1_outputs(168)) xor (layer1_outputs(4599)));
    layer2_outputs(8661) <= not(layer1_outputs(6374));
    layer2_outputs(8662) <= not(layer1_outputs(8852)) or (layer1_outputs(9166));
    layer2_outputs(8663) <= not(layer1_outputs(645));
    layer2_outputs(8664) <= (layer1_outputs(860)) and not (layer1_outputs(9387));
    layer2_outputs(8665) <= layer1_outputs(4328);
    layer2_outputs(8666) <= not((layer1_outputs(7190)) xor (layer1_outputs(2219)));
    layer2_outputs(8667) <= (layer1_outputs(5618)) and not (layer1_outputs(1859));
    layer2_outputs(8668) <= (layer1_outputs(5912)) or (layer1_outputs(9925));
    layer2_outputs(8669) <= not(layer1_outputs(8421)) or (layer1_outputs(7331));
    layer2_outputs(8670) <= not(layer1_outputs(1960));
    layer2_outputs(8671) <= not(layer1_outputs(4274));
    layer2_outputs(8672) <= not((layer1_outputs(1955)) xor (layer1_outputs(2554)));
    layer2_outputs(8673) <= not(layer1_outputs(4404)) or (layer1_outputs(3170));
    layer2_outputs(8674) <= (layer1_outputs(3174)) or (layer1_outputs(8312));
    layer2_outputs(8675) <= '0';
    layer2_outputs(8676) <= not(layer1_outputs(2632)) or (layer1_outputs(8436));
    layer2_outputs(8677) <= not(layer1_outputs(2003));
    layer2_outputs(8678) <= not(layer1_outputs(4495)) or (layer1_outputs(1625));
    layer2_outputs(8679) <= not((layer1_outputs(8612)) and (layer1_outputs(1080)));
    layer2_outputs(8680) <= (layer1_outputs(577)) and not (layer1_outputs(2053));
    layer2_outputs(8681) <= (layer1_outputs(3614)) and not (layer1_outputs(4237));
    layer2_outputs(8682) <= layer1_outputs(2681);
    layer2_outputs(8683) <= not((layer1_outputs(6492)) or (layer1_outputs(7715)));
    layer2_outputs(8684) <= layer1_outputs(542);
    layer2_outputs(8685) <= not(layer1_outputs(6415)) or (layer1_outputs(1203));
    layer2_outputs(8686) <= (layer1_outputs(1882)) and not (layer1_outputs(10199));
    layer2_outputs(8687) <= not(layer1_outputs(1988));
    layer2_outputs(8688) <= '0';
    layer2_outputs(8689) <= not((layer1_outputs(9794)) xor (layer1_outputs(4436)));
    layer2_outputs(8690) <= not(layer1_outputs(5898));
    layer2_outputs(8691) <= layer1_outputs(2662);
    layer2_outputs(8692) <= layer1_outputs(2294);
    layer2_outputs(8693) <= not(layer1_outputs(143));
    layer2_outputs(8694) <= layer1_outputs(9315);
    layer2_outputs(8695) <= layer1_outputs(3569);
    layer2_outputs(8696) <= (layer1_outputs(1815)) xor (layer1_outputs(1096));
    layer2_outputs(8697) <= '1';
    layer2_outputs(8698) <= (layer1_outputs(8337)) xor (layer1_outputs(5084));
    layer2_outputs(8699) <= not(layer1_outputs(5913));
    layer2_outputs(8700) <= (layer1_outputs(2894)) and not (layer1_outputs(5604));
    layer2_outputs(8701) <= not((layer1_outputs(6996)) xor (layer1_outputs(1957)));
    layer2_outputs(8702) <= layer1_outputs(9851);
    layer2_outputs(8703) <= layer1_outputs(1478);
    layer2_outputs(8704) <= not(layer1_outputs(7297));
    layer2_outputs(8705) <= (layer1_outputs(2454)) and (layer1_outputs(9323));
    layer2_outputs(8706) <= layer1_outputs(1695);
    layer2_outputs(8707) <= not(layer1_outputs(5818));
    layer2_outputs(8708) <= (layer1_outputs(3450)) and not (layer1_outputs(8696));
    layer2_outputs(8709) <= not((layer1_outputs(5260)) or (layer1_outputs(5727)));
    layer2_outputs(8710) <= '0';
    layer2_outputs(8711) <= (layer1_outputs(2481)) and (layer1_outputs(3306));
    layer2_outputs(8712) <= not(layer1_outputs(4802)) or (layer1_outputs(5360));
    layer2_outputs(8713) <= (layer1_outputs(8529)) and not (layer1_outputs(5132));
    layer2_outputs(8714) <= not(layer1_outputs(270));
    layer2_outputs(8715) <= layer1_outputs(7147);
    layer2_outputs(8716) <= not(layer1_outputs(9785));
    layer2_outputs(8717) <= (layer1_outputs(7858)) and not (layer1_outputs(5843));
    layer2_outputs(8718) <= not((layer1_outputs(343)) or (layer1_outputs(2020)));
    layer2_outputs(8719) <= layer1_outputs(10139);
    layer2_outputs(8720) <= layer1_outputs(10053);
    layer2_outputs(8721) <= (layer1_outputs(2178)) and not (layer1_outputs(6007));
    layer2_outputs(8722) <= '1';
    layer2_outputs(8723) <= not(layer1_outputs(4074));
    layer2_outputs(8724) <= (layer1_outputs(9116)) or (layer1_outputs(6923));
    layer2_outputs(8725) <= not((layer1_outputs(8412)) or (layer1_outputs(750)));
    layer2_outputs(8726) <= not(layer1_outputs(1982));
    layer2_outputs(8727) <= layer1_outputs(3255);
    layer2_outputs(8728) <= not((layer1_outputs(4496)) or (layer1_outputs(6172)));
    layer2_outputs(8729) <= (layer1_outputs(6790)) xor (layer1_outputs(5149));
    layer2_outputs(8730) <= not((layer1_outputs(5353)) or (layer1_outputs(8322)));
    layer2_outputs(8731) <= (layer1_outputs(2673)) and not (layer1_outputs(8846));
    layer2_outputs(8732) <= (layer1_outputs(4998)) and (layer1_outputs(8391));
    layer2_outputs(8733) <= not(layer1_outputs(6357)) or (layer1_outputs(8667));
    layer2_outputs(8734) <= layer1_outputs(5103);
    layer2_outputs(8735) <= not(layer1_outputs(5060));
    layer2_outputs(8736) <= (layer1_outputs(5708)) and not (layer1_outputs(2853));
    layer2_outputs(8737) <= not((layer1_outputs(7404)) and (layer1_outputs(8856)));
    layer2_outputs(8738) <= not(layer1_outputs(5739)) or (layer1_outputs(6004));
    layer2_outputs(8739) <= not(layer1_outputs(10009));
    layer2_outputs(8740) <= not((layer1_outputs(379)) xor (layer1_outputs(5604)));
    layer2_outputs(8741) <= layer1_outputs(3984);
    layer2_outputs(8742) <= layer1_outputs(8543);
    layer2_outputs(8743) <= '1';
    layer2_outputs(8744) <= not(layer1_outputs(493));
    layer2_outputs(8745) <= not(layer1_outputs(34));
    layer2_outputs(8746) <= not(layer1_outputs(6171)) or (layer1_outputs(1356));
    layer2_outputs(8747) <= not(layer1_outputs(1722));
    layer2_outputs(8748) <= (layer1_outputs(1869)) and not (layer1_outputs(6993));
    layer2_outputs(8749) <= layer1_outputs(4363);
    layer2_outputs(8750) <= not(layer1_outputs(5335));
    layer2_outputs(8751) <= '1';
    layer2_outputs(8752) <= not(layer1_outputs(5368)) or (layer1_outputs(4268));
    layer2_outputs(8753) <= not((layer1_outputs(5995)) or (layer1_outputs(6583)));
    layer2_outputs(8754) <= (layer1_outputs(1547)) xor (layer1_outputs(9406));
    layer2_outputs(8755) <= not(layer1_outputs(4960)) or (layer1_outputs(2751));
    layer2_outputs(8756) <= not((layer1_outputs(7537)) and (layer1_outputs(5025)));
    layer2_outputs(8757) <= not(layer1_outputs(4628));
    layer2_outputs(8758) <= layer1_outputs(9071);
    layer2_outputs(8759) <= not(layer1_outputs(6954)) or (layer1_outputs(7856));
    layer2_outputs(8760) <= (layer1_outputs(3109)) or (layer1_outputs(7323));
    layer2_outputs(8761) <= (layer1_outputs(4446)) xor (layer1_outputs(4700));
    layer2_outputs(8762) <= (layer1_outputs(3284)) and (layer1_outputs(826));
    layer2_outputs(8763) <= (layer1_outputs(7549)) and not (layer1_outputs(3388));
    layer2_outputs(8764) <= layer1_outputs(4929);
    layer2_outputs(8765) <= (layer1_outputs(7188)) and (layer1_outputs(2987));
    layer2_outputs(8766) <= '1';
    layer2_outputs(8767) <= (layer1_outputs(9524)) xor (layer1_outputs(9507));
    layer2_outputs(8768) <= not((layer1_outputs(535)) xor (layer1_outputs(3317)));
    layer2_outputs(8769) <= (layer1_outputs(8911)) and (layer1_outputs(6389));
    layer2_outputs(8770) <= layer1_outputs(5537);
    layer2_outputs(8771) <= (layer1_outputs(9192)) xor (layer1_outputs(192));
    layer2_outputs(8772) <= (layer1_outputs(8500)) and not (layer1_outputs(8497));
    layer2_outputs(8773) <= not(layer1_outputs(7596));
    layer2_outputs(8774) <= layer1_outputs(5772);
    layer2_outputs(8775) <= not(layer1_outputs(8181));
    layer2_outputs(8776) <= layer1_outputs(433);
    layer2_outputs(8777) <= layer1_outputs(6146);
    layer2_outputs(8778) <= not((layer1_outputs(1823)) and (layer1_outputs(2725)));
    layer2_outputs(8779) <= layer1_outputs(5030);
    layer2_outputs(8780) <= '0';
    layer2_outputs(8781) <= not(layer1_outputs(1305));
    layer2_outputs(8782) <= '1';
    layer2_outputs(8783) <= (layer1_outputs(9271)) and not (layer1_outputs(377));
    layer2_outputs(8784) <= layer1_outputs(1194);
    layer2_outputs(8785) <= (layer1_outputs(9553)) and not (layer1_outputs(3266));
    layer2_outputs(8786) <= not(layer1_outputs(4215)) or (layer1_outputs(2356));
    layer2_outputs(8787) <= (layer1_outputs(3262)) or (layer1_outputs(5840));
    layer2_outputs(8788) <= layer1_outputs(3371);
    layer2_outputs(8789) <= not(layer1_outputs(4385)) or (layer1_outputs(2335));
    layer2_outputs(8790) <= not(layer1_outputs(8845));
    layer2_outputs(8791) <= layer1_outputs(4922);
    layer2_outputs(8792) <= '1';
    layer2_outputs(8793) <= (layer1_outputs(2398)) or (layer1_outputs(921));
    layer2_outputs(8794) <= (layer1_outputs(6742)) or (layer1_outputs(4959));
    layer2_outputs(8795) <= (layer1_outputs(5207)) or (layer1_outputs(4315));
    layer2_outputs(8796) <= not((layer1_outputs(6915)) or (layer1_outputs(5183)));
    layer2_outputs(8797) <= layer1_outputs(6861);
    layer2_outputs(8798) <= not(layer1_outputs(10047));
    layer2_outputs(8799) <= layer1_outputs(4310);
    layer2_outputs(8800) <= (layer1_outputs(4033)) and not (layer1_outputs(7484));
    layer2_outputs(8801) <= layer1_outputs(6952);
    layer2_outputs(8802) <= layer1_outputs(4568);
    layer2_outputs(8803) <= (layer1_outputs(7226)) xor (layer1_outputs(5139));
    layer2_outputs(8804) <= not(layer1_outputs(2626));
    layer2_outputs(8805) <= (layer1_outputs(7772)) and not (layer1_outputs(5911));
    layer2_outputs(8806) <= not(layer1_outputs(5214));
    layer2_outputs(8807) <= (layer1_outputs(7148)) or (layer1_outputs(6058));
    layer2_outputs(8808) <= (layer1_outputs(3)) xor (layer1_outputs(6088));
    layer2_outputs(8809) <= layer1_outputs(8661);
    layer2_outputs(8810) <= (layer1_outputs(8585)) and not (layer1_outputs(3463));
    layer2_outputs(8811) <= layer1_outputs(7531);
    layer2_outputs(8812) <= not(layer1_outputs(5896)) or (layer1_outputs(8599));
    layer2_outputs(8813) <= not((layer1_outputs(8552)) xor (layer1_outputs(1608)));
    layer2_outputs(8814) <= not(layer1_outputs(4927)) or (layer1_outputs(9005));
    layer2_outputs(8815) <= not((layer1_outputs(5095)) and (layer1_outputs(109)));
    layer2_outputs(8816) <= (layer1_outputs(1414)) xor (layer1_outputs(5256));
    layer2_outputs(8817) <= (layer1_outputs(6573)) and not (layer1_outputs(6143));
    layer2_outputs(8818) <= '1';
    layer2_outputs(8819) <= not(layer1_outputs(208)) or (layer1_outputs(8789));
    layer2_outputs(8820) <= not(layer1_outputs(6640));
    layer2_outputs(8821) <= (layer1_outputs(2524)) and not (layer1_outputs(7580));
    layer2_outputs(8822) <= not(layer1_outputs(4815));
    layer2_outputs(8823) <= not(layer1_outputs(8110));
    layer2_outputs(8824) <= layer1_outputs(2780);
    layer2_outputs(8825) <= (layer1_outputs(5494)) and not (layer1_outputs(10049));
    layer2_outputs(8826) <= not(layer1_outputs(10019));
    layer2_outputs(8827) <= '1';
    layer2_outputs(8828) <= (layer1_outputs(6578)) and not (layer1_outputs(8162));
    layer2_outputs(8829) <= layer1_outputs(2855);
    layer2_outputs(8830) <= not(layer1_outputs(1793));
    layer2_outputs(8831) <= (layer1_outputs(3874)) xor (layer1_outputs(2407));
    layer2_outputs(8832) <= (layer1_outputs(9436)) and (layer1_outputs(3297));
    layer2_outputs(8833) <= (layer1_outputs(8398)) and not (layer1_outputs(3967));
    layer2_outputs(8834) <= not(layer1_outputs(2261));
    layer2_outputs(8835) <= not(layer1_outputs(9847));
    layer2_outputs(8836) <= layer1_outputs(6932);
    layer2_outputs(8837) <= layer1_outputs(758);
    layer2_outputs(8838) <= (layer1_outputs(6437)) and (layer1_outputs(6021));
    layer2_outputs(8839) <= not(layer1_outputs(6109));
    layer2_outputs(8840) <= (layer1_outputs(1771)) and (layer1_outputs(3243));
    layer2_outputs(8841) <= layer1_outputs(188);
    layer2_outputs(8842) <= not((layer1_outputs(5479)) or (layer1_outputs(3953)));
    layer2_outputs(8843) <= not((layer1_outputs(370)) or (layer1_outputs(5294)));
    layer2_outputs(8844) <= not(layer1_outputs(9863));
    layer2_outputs(8845) <= (layer1_outputs(1585)) or (layer1_outputs(8057));
    layer2_outputs(8846) <= (layer1_outputs(8464)) xor (layer1_outputs(6182));
    layer2_outputs(8847) <= not(layer1_outputs(4184));
    layer2_outputs(8848) <= layer1_outputs(9480);
    layer2_outputs(8849) <= layer1_outputs(8727);
    layer2_outputs(8850) <= layer1_outputs(9945);
    layer2_outputs(8851) <= not((layer1_outputs(8775)) or (layer1_outputs(1658)));
    layer2_outputs(8852) <= not(layer1_outputs(6029));
    layer2_outputs(8853) <= '1';
    layer2_outputs(8854) <= not(layer1_outputs(5817));
    layer2_outputs(8855) <= not(layer1_outputs(7990)) or (layer1_outputs(1874));
    layer2_outputs(8856) <= not((layer1_outputs(4125)) or (layer1_outputs(3630)));
    layer2_outputs(8857) <= layer1_outputs(6332);
    layer2_outputs(8858) <= layer1_outputs(1617);
    layer2_outputs(8859) <= layer1_outputs(2055);
    layer2_outputs(8860) <= not((layer1_outputs(1826)) and (layer1_outputs(7508)));
    layer2_outputs(8861) <= '1';
    layer2_outputs(8862) <= not(layer1_outputs(3799)) or (layer1_outputs(74));
    layer2_outputs(8863) <= (layer1_outputs(5270)) xor (layer1_outputs(2355));
    layer2_outputs(8864) <= not((layer1_outputs(57)) or (layer1_outputs(9174)));
    layer2_outputs(8865) <= not(layer1_outputs(2488)) or (layer1_outputs(3477));
    layer2_outputs(8866) <= not((layer1_outputs(1933)) and (layer1_outputs(2876)));
    layer2_outputs(8867) <= '1';
    layer2_outputs(8868) <= not(layer1_outputs(6164));
    layer2_outputs(8869) <= not(layer1_outputs(6728));
    layer2_outputs(8870) <= not((layer1_outputs(309)) xor (layer1_outputs(13)));
    layer2_outputs(8871) <= layer1_outputs(5671);
    layer2_outputs(8872) <= not(layer1_outputs(286));
    layer2_outputs(8873) <= not((layer1_outputs(4702)) and (layer1_outputs(9830)));
    layer2_outputs(8874) <= '1';
    layer2_outputs(8875) <= (layer1_outputs(2770)) and not (layer1_outputs(8168));
    layer2_outputs(8876) <= (layer1_outputs(218)) and (layer1_outputs(2945));
    layer2_outputs(8877) <= not(layer1_outputs(7879));
    layer2_outputs(8878) <= '0';
    layer2_outputs(8879) <= layer1_outputs(8760);
    layer2_outputs(8880) <= '1';
    layer2_outputs(8881) <= layer1_outputs(3053);
    layer2_outputs(8882) <= (layer1_outputs(8185)) xor (layer1_outputs(10198));
    layer2_outputs(8883) <= layer1_outputs(1453);
    layer2_outputs(8884) <= not((layer1_outputs(1958)) and (layer1_outputs(9957)));
    layer2_outputs(8885) <= not(layer1_outputs(3393));
    layer2_outputs(8886) <= (layer1_outputs(1296)) and not (layer1_outputs(9004));
    layer2_outputs(8887) <= (layer1_outputs(4723)) xor (layer1_outputs(2928));
    layer2_outputs(8888) <= not(layer1_outputs(7626));
    layer2_outputs(8889) <= not(layer1_outputs(2077));
    layer2_outputs(8890) <= (layer1_outputs(5884)) xor (layer1_outputs(9383));
    layer2_outputs(8891) <= not((layer1_outputs(441)) xor (layer1_outputs(6387)));
    layer2_outputs(8892) <= (layer1_outputs(6423)) xor (layer1_outputs(7674));
    layer2_outputs(8893) <= not(layer1_outputs(5112)) or (layer1_outputs(1769));
    layer2_outputs(8894) <= layer1_outputs(3998);
    layer2_outputs(8895) <= (layer1_outputs(6436)) and not (layer1_outputs(6396));
    layer2_outputs(8896) <= not(layer1_outputs(8233));
    layer2_outputs(8897) <= not(layer1_outputs(2191)) or (layer1_outputs(3334));
    layer2_outputs(8898) <= '1';
    layer2_outputs(8899) <= (layer1_outputs(7036)) or (layer1_outputs(7617));
    layer2_outputs(8900) <= not(layer1_outputs(9406));
    layer2_outputs(8901) <= layer1_outputs(2015);
    layer2_outputs(8902) <= layer1_outputs(3824);
    layer2_outputs(8903) <= layer1_outputs(3902);
    layer2_outputs(8904) <= (layer1_outputs(4415)) and (layer1_outputs(9472));
    layer2_outputs(8905) <= (layer1_outputs(9138)) or (layer1_outputs(4946));
    layer2_outputs(8906) <= layer1_outputs(4027);
    layer2_outputs(8907) <= not(layer1_outputs(8213)) or (layer1_outputs(5239));
    layer2_outputs(8908) <= (layer1_outputs(3652)) and not (layer1_outputs(2401));
    layer2_outputs(8909) <= '0';
    layer2_outputs(8910) <= layer1_outputs(6407);
    layer2_outputs(8911) <= not(layer1_outputs(777));
    layer2_outputs(8912) <= not(layer1_outputs(8515));
    layer2_outputs(8913) <= not(layer1_outputs(2000)) or (layer1_outputs(7204));
    layer2_outputs(8914) <= (layer1_outputs(5511)) and not (layer1_outputs(2179));
    layer2_outputs(8915) <= not(layer1_outputs(9105));
    layer2_outputs(8916) <= not(layer1_outputs(9684));
    layer2_outputs(8917) <= layer1_outputs(8047);
    layer2_outputs(8918) <= not(layer1_outputs(7548)) or (layer1_outputs(8097));
    layer2_outputs(8919) <= layer1_outputs(5652);
    layer2_outputs(8920) <= not(layer1_outputs(7823));
    layer2_outputs(8921) <= not((layer1_outputs(6657)) and (layer1_outputs(4924)));
    layer2_outputs(8922) <= '0';
    layer2_outputs(8923) <= (layer1_outputs(2110)) and not (layer1_outputs(4796));
    layer2_outputs(8924) <= layer1_outputs(9916);
    layer2_outputs(8925) <= not(layer1_outputs(5564));
    layer2_outputs(8926) <= not((layer1_outputs(47)) and (layer1_outputs(315)));
    layer2_outputs(8927) <= not(layer1_outputs(6848)) or (layer1_outputs(3836));
    layer2_outputs(8928) <= layer1_outputs(510);
    layer2_outputs(8929) <= not(layer1_outputs(1153));
    layer2_outputs(8930) <= (layer1_outputs(6908)) xor (layer1_outputs(4668));
    layer2_outputs(8931) <= not(layer1_outputs(472)) or (layer1_outputs(7099));
    layer2_outputs(8932) <= '1';
    layer2_outputs(8933) <= layer1_outputs(3265);
    layer2_outputs(8934) <= not(layer1_outputs(1793));
    layer2_outputs(8935) <= not(layer1_outputs(1921));
    layer2_outputs(8936) <= not((layer1_outputs(1892)) or (layer1_outputs(1920)));
    layer2_outputs(8937) <= (layer1_outputs(4957)) and not (layer1_outputs(6071));
    layer2_outputs(8938) <= not(layer1_outputs(2287));
    layer2_outputs(8939) <= '1';
    layer2_outputs(8940) <= layer1_outputs(495);
    layer2_outputs(8941) <= (layer1_outputs(7712)) and not (layer1_outputs(1170));
    layer2_outputs(8942) <= not(layer1_outputs(4890));
    layer2_outputs(8943) <= not(layer1_outputs(1685)) or (layer1_outputs(3005));
    layer2_outputs(8944) <= not(layer1_outputs(6236));
    layer2_outputs(8945) <= (layer1_outputs(8072)) or (layer1_outputs(9705));
    layer2_outputs(8946) <= not(layer1_outputs(8176));
    layer2_outputs(8947) <= not(layer1_outputs(10166)) or (layer1_outputs(1107));
    layer2_outputs(8948) <= not(layer1_outputs(7223)) or (layer1_outputs(8096));
    layer2_outputs(8949) <= not((layer1_outputs(4702)) and (layer1_outputs(5367)));
    layer2_outputs(8950) <= '1';
    layer2_outputs(8951) <= layer1_outputs(5039);
    layer2_outputs(8952) <= layer1_outputs(1388);
    layer2_outputs(8953) <= not(layer1_outputs(1711));
    layer2_outputs(8954) <= (layer1_outputs(7810)) and not (layer1_outputs(1004));
    layer2_outputs(8955) <= not(layer1_outputs(2106));
    layer2_outputs(8956) <= not(layer1_outputs(4489));
    layer2_outputs(8957) <= not((layer1_outputs(2474)) or (layer1_outputs(4123)));
    layer2_outputs(8958) <= (layer1_outputs(2031)) and not (layer1_outputs(9348));
    layer2_outputs(8959) <= (layer1_outputs(3717)) xor (layer1_outputs(1214));
    layer2_outputs(8960) <= not((layer1_outputs(4642)) or (layer1_outputs(8576)));
    layer2_outputs(8961) <= (layer1_outputs(6659)) or (layer1_outputs(4461));
    layer2_outputs(8962) <= layer1_outputs(8138);
    layer2_outputs(8963) <= layer1_outputs(1518);
    layer2_outputs(8964) <= (layer1_outputs(4544)) and (layer1_outputs(3883));
    layer2_outputs(8965) <= not(layer1_outputs(4992)) or (layer1_outputs(4313));
    layer2_outputs(8966) <= not(layer1_outputs(1918));
    layer2_outputs(8967) <= not(layer1_outputs(6307));
    layer2_outputs(8968) <= (layer1_outputs(9454)) and not (layer1_outputs(6104));
    layer2_outputs(8969) <= (layer1_outputs(1430)) or (layer1_outputs(9073));
    layer2_outputs(8970) <= (layer1_outputs(9910)) xor (layer1_outputs(2758));
    layer2_outputs(8971) <= (layer1_outputs(5032)) and not (layer1_outputs(9589));
    layer2_outputs(8972) <= not((layer1_outputs(3378)) or (layer1_outputs(7232)));
    layer2_outputs(8973) <= not(layer1_outputs(2744)) or (layer1_outputs(5458));
    layer2_outputs(8974) <= not((layer1_outputs(892)) and (layer1_outputs(8830)));
    layer2_outputs(8975) <= not(layer1_outputs(8766)) or (layer1_outputs(6023));
    layer2_outputs(8976) <= not(layer1_outputs(3560)) or (layer1_outputs(6647));
    layer2_outputs(8977) <= not(layer1_outputs(9449));
    layer2_outputs(8978) <= layer1_outputs(7478);
    layer2_outputs(8979) <= not((layer1_outputs(7202)) or (layer1_outputs(166)));
    layer2_outputs(8980) <= not((layer1_outputs(545)) xor (layer1_outputs(6293)));
    layer2_outputs(8981) <= layer1_outputs(4767);
    layer2_outputs(8982) <= (layer1_outputs(5559)) or (layer1_outputs(1396));
    layer2_outputs(8983) <= not(layer1_outputs(3662));
    layer2_outputs(8984) <= (layer1_outputs(9183)) and (layer1_outputs(6382));
    layer2_outputs(8985) <= not(layer1_outputs(6318)) or (layer1_outputs(1603));
    layer2_outputs(8986) <= (layer1_outputs(9713)) and not (layer1_outputs(10051));
    layer2_outputs(8987) <= layer1_outputs(6383);
    layer2_outputs(8988) <= layer1_outputs(9646);
    layer2_outputs(8989) <= '0';
    layer2_outputs(8990) <= not(layer1_outputs(6828)) or (layer1_outputs(8007));
    layer2_outputs(8991) <= not(layer1_outputs(1751));
    layer2_outputs(8992) <= not((layer1_outputs(1314)) or (layer1_outputs(5308)));
    layer2_outputs(8993) <= not((layer1_outputs(8354)) or (layer1_outputs(3802)));
    layer2_outputs(8994) <= (layer1_outputs(464)) xor (layer1_outputs(4725));
    layer2_outputs(8995) <= layer1_outputs(6486);
    layer2_outputs(8996) <= not(layer1_outputs(8462));
    layer2_outputs(8997) <= not(layer1_outputs(7611));
    layer2_outputs(8998) <= (layer1_outputs(2515)) and not (layer1_outputs(709));
    layer2_outputs(8999) <= not((layer1_outputs(3064)) and (layer1_outputs(1171)));
    layer2_outputs(9000) <= not(layer1_outputs(9771));
    layer2_outputs(9001) <= not(layer1_outputs(3234)) or (layer1_outputs(3172));
    layer2_outputs(9002) <= layer1_outputs(6060);
    layer2_outputs(9003) <= not(layer1_outputs(684));
    layer2_outputs(9004) <= layer1_outputs(4522);
    layer2_outputs(9005) <= not(layer1_outputs(5608));
    layer2_outputs(9006) <= not(layer1_outputs(5379));
    layer2_outputs(9007) <= (layer1_outputs(3898)) and not (layer1_outputs(3154));
    layer2_outputs(9008) <= layer1_outputs(318);
    layer2_outputs(9009) <= not((layer1_outputs(324)) or (layer1_outputs(6145)));
    layer2_outputs(9010) <= (layer1_outputs(835)) and (layer1_outputs(5688));
    layer2_outputs(9011) <= (layer1_outputs(6453)) or (layer1_outputs(10007));
    layer2_outputs(9012) <= not(layer1_outputs(2645)) or (layer1_outputs(2822));
    layer2_outputs(9013) <= not((layer1_outputs(9340)) and (layer1_outputs(6919)));
    layer2_outputs(9014) <= layer1_outputs(7937);
    layer2_outputs(9015) <= (layer1_outputs(9686)) and (layer1_outputs(4796));
    layer2_outputs(9016) <= not(layer1_outputs(8240)) or (layer1_outputs(8044));
    layer2_outputs(9017) <= (layer1_outputs(2745)) and not (layer1_outputs(1468));
    layer2_outputs(9018) <= (layer1_outputs(6679)) and not (layer1_outputs(5157));
    layer2_outputs(9019) <= layer1_outputs(5573);
    layer2_outputs(9020) <= not(layer1_outputs(9219)) or (layer1_outputs(4269));
    layer2_outputs(9021) <= layer1_outputs(5616);
    layer2_outputs(9022) <= '0';
    layer2_outputs(9023) <= (layer1_outputs(3789)) and not (layer1_outputs(3917));
    layer2_outputs(9024) <= (layer1_outputs(1176)) and not (layer1_outputs(8450));
    layer2_outputs(9025) <= (layer1_outputs(4707)) and not (layer1_outputs(1253));
    layer2_outputs(9026) <= not(layer1_outputs(3929)) or (layer1_outputs(6775));
    layer2_outputs(9027) <= '1';
    layer2_outputs(9028) <= not(layer1_outputs(8563)) or (layer1_outputs(1753));
    layer2_outputs(9029) <= not(layer1_outputs(4837)) or (layer1_outputs(853));
    layer2_outputs(9030) <= (layer1_outputs(10011)) and not (layer1_outputs(3024));
    layer2_outputs(9031) <= not(layer1_outputs(8805));
    layer2_outputs(9032) <= not(layer1_outputs(22));
    layer2_outputs(9033) <= not(layer1_outputs(2707));
    layer2_outputs(9034) <= (layer1_outputs(8594)) xor (layer1_outputs(5732));
    layer2_outputs(9035) <= layer1_outputs(2826);
    layer2_outputs(9036) <= '1';
    layer2_outputs(9037) <= layer1_outputs(6195);
    layer2_outputs(9038) <= layer1_outputs(232);
    layer2_outputs(9039) <= (layer1_outputs(1917)) xor (layer1_outputs(2869));
    layer2_outputs(9040) <= not((layer1_outputs(7290)) xor (layer1_outputs(3665)));
    layer2_outputs(9041) <= not((layer1_outputs(3652)) or (layer1_outputs(8323)));
    layer2_outputs(9042) <= (layer1_outputs(3087)) xor (layer1_outputs(4674));
    layer2_outputs(9043) <= not(layer1_outputs(9878));
    layer2_outputs(9044) <= (layer1_outputs(8224)) and not (layer1_outputs(1818));
    layer2_outputs(9045) <= layer1_outputs(3456);
    layer2_outputs(9046) <= (layer1_outputs(9599)) xor (layer1_outputs(7950));
    layer2_outputs(9047) <= (layer1_outputs(2803)) or (layer1_outputs(370));
    layer2_outputs(9048) <= layer1_outputs(3662);
    layer2_outputs(9049) <= '0';
    layer2_outputs(9050) <= not(layer1_outputs(3340)) or (layer1_outputs(8544));
    layer2_outputs(9051) <= not((layer1_outputs(153)) and (layer1_outputs(484)));
    layer2_outputs(9052) <= not(layer1_outputs(4023));
    layer2_outputs(9053) <= not((layer1_outputs(9877)) or (layer1_outputs(5585)));
    layer2_outputs(9054) <= '1';
    layer2_outputs(9055) <= (layer1_outputs(829)) and not (layer1_outputs(3820));
    layer2_outputs(9056) <= not((layer1_outputs(8368)) or (layer1_outputs(814)));
    layer2_outputs(9057) <= not((layer1_outputs(4531)) or (layer1_outputs(871)));
    layer2_outputs(9058) <= (layer1_outputs(9529)) and (layer1_outputs(2797));
    layer2_outputs(9059) <= layer1_outputs(890);
    layer2_outputs(9060) <= '1';
    layer2_outputs(9061) <= not(layer1_outputs(9855));
    layer2_outputs(9062) <= not(layer1_outputs(7345)) or (layer1_outputs(7278));
    layer2_outputs(9063) <= (layer1_outputs(2901)) and not (layer1_outputs(1241));
    layer2_outputs(9064) <= not(layer1_outputs(8088)) or (layer1_outputs(2157));
    layer2_outputs(9065) <= (layer1_outputs(4011)) and not (layer1_outputs(4073));
    layer2_outputs(9066) <= (layer1_outputs(8540)) and not (layer1_outputs(9172));
    layer2_outputs(9067) <= '0';
    layer2_outputs(9068) <= layer1_outputs(4357);
    layer2_outputs(9069) <= not((layer1_outputs(872)) or (layer1_outputs(1767)));
    layer2_outputs(9070) <= layer1_outputs(7292);
    layer2_outputs(9071) <= not(layer1_outputs(124));
    layer2_outputs(9072) <= (layer1_outputs(1288)) and not (layer1_outputs(6601));
    layer2_outputs(9073) <= not((layer1_outputs(2228)) and (layer1_outputs(6131)));
    layer2_outputs(9074) <= (layer1_outputs(568)) or (layer1_outputs(1231));
    layer2_outputs(9075) <= (layer1_outputs(9544)) or (layer1_outputs(7276));
    layer2_outputs(9076) <= (layer1_outputs(2896)) and not (layer1_outputs(5791));
    layer2_outputs(9077) <= not((layer1_outputs(6865)) xor (layer1_outputs(7365)));
    layer2_outputs(9078) <= layer1_outputs(6676);
    layer2_outputs(9079) <= not((layer1_outputs(6006)) xor (layer1_outputs(7558)));
    layer2_outputs(9080) <= not(layer1_outputs(1468)) or (layer1_outputs(8767));
    layer2_outputs(9081) <= (layer1_outputs(5235)) or (layer1_outputs(8772));
    layer2_outputs(9082) <= (layer1_outputs(2238)) and not (layer1_outputs(3792));
    layer2_outputs(9083) <= not(layer1_outputs(9828));
    layer2_outputs(9084) <= not((layer1_outputs(1853)) xor (layer1_outputs(3773)));
    layer2_outputs(9085) <= not((layer1_outputs(4241)) or (layer1_outputs(2652)));
    layer2_outputs(9086) <= (layer1_outputs(4006)) or (layer1_outputs(4780));
    layer2_outputs(9087) <= layer1_outputs(9558);
    layer2_outputs(9088) <= (layer1_outputs(6217)) and (layer1_outputs(8779));
    layer2_outputs(9089) <= '0';
    layer2_outputs(9090) <= (layer1_outputs(9136)) and not (layer1_outputs(4617));
    layer2_outputs(9091) <= layer1_outputs(7819);
    layer2_outputs(9092) <= not(layer1_outputs(3869)) or (layer1_outputs(8685));
    layer2_outputs(9093) <= not((layer1_outputs(6666)) or (layer1_outputs(1688)));
    layer2_outputs(9094) <= (layer1_outputs(4053)) xor (layer1_outputs(5193));
    layer2_outputs(9095) <= not(layer1_outputs(3425));
    layer2_outputs(9096) <= (layer1_outputs(3106)) xor (layer1_outputs(2993));
    layer2_outputs(9097) <= not(layer1_outputs(8297));
    layer2_outputs(9098) <= not(layer1_outputs(5561));
    layer2_outputs(9099) <= layer1_outputs(3570);
    layer2_outputs(9100) <= (layer1_outputs(3882)) and (layer1_outputs(9663));
    layer2_outputs(9101) <= layer1_outputs(254);
    layer2_outputs(9102) <= not((layer1_outputs(3213)) or (layer1_outputs(9252)));
    layer2_outputs(9103) <= not(layer1_outputs(2056)) or (layer1_outputs(6227));
    layer2_outputs(9104) <= (layer1_outputs(2427)) and not (layer1_outputs(3498));
    layer2_outputs(9105) <= layer1_outputs(7599);
    layer2_outputs(9106) <= layer1_outputs(4918);
    layer2_outputs(9107) <= layer1_outputs(798);
    layer2_outputs(9108) <= layer1_outputs(8894);
    layer2_outputs(9109) <= (layer1_outputs(3606)) and not (layer1_outputs(1378));
    layer2_outputs(9110) <= not((layer1_outputs(1077)) xor (layer1_outputs(4305)));
    layer2_outputs(9111) <= layer1_outputs(5353);
    layer2_outputs(9112) <= (layer1_outputs(10022)) and not (layer1_outputs(2022));
    layer2_outputs(9113) <= not((layer1_outputs(3558)) or (layer1_outputs(643)));
    layer2_outputs(9114) <= (layer1_outputs(4569)) and not (layer1_outputs(2394));
    layer2_outputs(9115) <= not(layer1_outputs(9068)) or (layer1_outputs(2346));
    layer2_outputs(9116) <= not(layer1_outputs(7101));
    layer2_outputs(9117) <= not((layer1_outputs(6600)) xor (layer1_outputs(5465)));
    layer2_outputs(9118) <= layer1_outputs(620);
    layer2_outputs(9119) <= (layer1_outputs(4087)) or (layer1_outputs(6210));
    layer2_outputs(9120) <= not(layer1_outputs(7049)) or (layer1_outputs(2239));
    layer2_outputs(9121) <= (layer1_outputs(116)) or (layer1_outputs(7436));
    layer2_outputs(9122) <= not(layer1_outputs(5205));
    layer2_outputs(9123) <= layer1_outputs(9127);
    layer2_outputs(9124) <= (layer1_outputs(8102)) xor (layer1_outputs(2850));
    layer2_outputs(9125) <= not(layer1_outputs(9285));
    layer2_outputs(9126) <= not(layer1_outputs(5561)) or (layer1_outputs(1393));
    layer2_outputs(9127) <= not(layer1_outputs(4997)) or (layer1_outputs(8978));
    layer2_outputs(9128) <= layer1_outputs(4920);
    layer2_outputs(9129) <= (layer1_outputs(9079)) and not (layer1_outputs(3202));
    layer2_outputs(9130) <= not(layer1_outputs(5598));
    layer2_outputs(9131) <= (layer1_outputs(5417)) and not (layer1_outputs(3299));
    layer2_outputs(9132) <= not((layer1_outputs(355)) or (layer1_outputs(5367)));
    layer2_outputs(9133) <= not(layer1_outputs(6643)) or (layer1_outputs(1375));
    layer2_outputs(9134) <= '1';
    layer2_outputs(9135) <= layer1_outputs(3365);
    layer2_outputs(9136) <= layer1_outputs(8226);
    layer2_outputs(9137) <= layer1_outputs(1027);
    layer2_outputs(9138) <= layer1_outputs(5375);
    layer2_outputs(9139) <= layer1_outputs(2317);
    layer2_outputs(9140) <= not(layer1_outputs(6605)) or (layer1_outputs(5526));
    layer2_outputs(9141) <= layer1_outputs(2924);
    layer2_outputs(9142) <= (layer1_outputs(2653)) xor (layer1_outputs(942));
    layer2_outputs(9143) <= not(layer1_outputs(851));
    layer2_outputs(9144) <= not(layer1_outputs(138));
    layer2_outputs(9145) <= not(layer1_outputs(1731)) or (layer1_outputs(6956));
    layer2_outputs(9146) <= not(layer1_outputs(2806)) or (layer1_outputs(4892));
    layer2_outputs(9147) <= not(layer1_outputs(99));
    layer2_outputs(9148) <= layer1_outputs(354);
    layer2_outputs(9149) <= not(layer1_outputs(4501)) or (layer1_outputs(9419));
    layer2_outputs(9150) <= (layer1_outputs(4060)) and (layer1_outputs(271));
    layer2_outputs(9151) <= layer1_outputs(7489);
    layer2_outputs(9152) <= not(layer1_outputs(8361));
    layer2_outputs(9153) <= not((layer1_outputs(3782)) and (layer1_outputs(1111)));
    layer2_outputs(9154) <= layer1_outputs(7457);
    layer2_outputs(9155) <= (layer1_outputs(6225)) xor (layer1_outputs(9232));
    layer2_outputs(9156) <= not(layer1_outputs(7333)) or (layer1_outputs(9997));
    layer2_outputs(9157) <= (layer1_outputs(4703)) and (layer1_outputs(2409));
    layer2_outputs(9158) <= not((layer1_outputs(8091)) or (layer1_outputs(10032)));
    layer2_outputs(9159) <= not((layer1_outputs(6730)) and (layer1_outputs(7435)));
    layer2_outputs(9160) <= '1';
    layer2_outputs(9161) <= '1';
    layer2_outputs(9162) <= layer1_outputs(321);
    layer2_outputs(9163) <= not(layer1_outputs(1684)) or (layer1_outputs(2402));
    layer2_outputs(9164) <= not((layer1_outputs(10021)) xor (layer1_outputs(10081)));
    layer2_outputs(9165) <= layer1_outputs(7664);
    layer2_outputs(9166) <= '0';
    layer2_outputs(9167) <= not((layer1_outputs(1797)) or (layer1_outputs(9923)));
    layer2_outputs(9168) <= not((layer1_outputs(2111)) and (layer1_outputs(5778)));
    layer2_outputs(9169) <= not((layer1_outputs(9355)) xor (layer1_outputs(4286)));
    layer2_outputs(9170) <= '0';
    layer2_outputs(9171) <= not(layer1_outputs(1043));
    layer2_outputs(9172) <= (layer1_outputs(4398)) xor (layer1_outputs(9194));
    layer2_outputs(9173) <= not(layer1_outputs(6953));
    layer2_outputs(9174) <= not(layer1_outputs(7119)) or (layer1_outputs(8671));
    layer2_outputs(9175) <= (layer1_outputs(7000)) and not (layer1_outputs(2504));
    layer2_outputs(9176) <= (layer1_outputs(8603)) xor (layer1_outputs(3860));
    layer2_outputs(9177) <= (layer1_outputs(5723)) and (layer1_outputs(1806));
    layer2_outputs(9178) <= not((layer1_outputs(6780)) or (layer1_outputs(4609)));
    layer2_outputs(9179) <= not((layer1_outputs(3621)) or (layer1_outputs(1093)));
    layer2_outputs(9180) <= (layer1_outputs(3272)) or (layer1_outputs(84));
    layer2_outputs(9181) <= not((layer1_outputs(10181)) and (layer1_outputs(9)));
    layer2_outputs(9182) <= not(layer1_outputs(6386));
    layer2_outputs(9183) <= (layer1_outputs(7008)) and not (layer1_outputs(9375));
    layer2_outputs(9184) <= layer1_outputs(5620);
    layer2_outputs(9185) <= layer1_outputs(8901);
    layer2_outputs(9186) <= not(layer1_outputs(7994)) or (layer1_outputs(1778));
    layer2_outputs(9187) <= not((layer1_outputs(568)) xor (layer1_outputs(2462)));
    layer2_outputs(9188) <= layer1_outputs(1289);
    layer2_outputs(9189) <= '0';
    layer2_outputs(9190) <= not(layer1_outputs(9932));
    layer2_outputs(9191) <= not((layer1_outputs(8986)) and (layer1_outputs(877)));
    layer2_outputs(9192) <= not((layer1_outputs(7425)) or (layer1_outputs(3037)));
    layer2_outputs(9193) <= layer1_outputs(5467);
    layer2_outputs(9194) <= (layer1_outputs(7336)) or (layer1_outputs(1734));
    layer2_outputs(9195) <= '0';
    layer2_outputs(9196) <= not(layer1_outputs(400)) or (layer1_outputs(8888));
    layer2_outputs(9197) <= not((layer1_outputs(799)) xor (layer1_outputs(3793)));
    layer2_outputs(9198) <= layer1_outputs(3577);
    layer2_outputs(9199) <= not(layer1_outputs(703)) or (layer1_outputs(2343));
    layer2_outputs(9200) <= layer1_outputs(2678);
    layer2_outputs(9201) <= layer1_outputs(6097);
    layer2_outputs(9202) <= (layer1_outputs(6179)) or (layer1_outputs(3358));
    layer2_outputs(9203) <= not(layer1_outputs(7701));
    layer2_outputs(9204) <= (layer1_outputs(4360)) and not (layer1_outputs(6808));
    layer2_outputs(9205) <= '1';
    layer2_outputs(9206) <= not(layer1_outputs(3610));
    layer2_outputs(9207) <= (layer1_outputs(1999)) and not (layer1_outputs(1888));
    layer2_outputs(9208) <= layer1_outputs(9539);
    layer2_outputs(9209) <= (layer1_outputs(8821)) and not (layer1_outputs(489));
    layer2_outputs(9210) <= not(layer1_outputs(9168)) or (layer1_outputs(3226));
    layer2_outputs(9211) <= '1';
    layer2_outputs(9212) <= (layer1_outputs(7542)) xor (layer1_outputs(1894));
    layer2_outputs(9213) <= not(layer1_outputs(4909));
    layer2_outputs(9214) <= (layer1_outputs(7295)) xor (layer1_outputs(8375));
    layer2_outputs(9215) <= (layer1_outputs(7293)) and (layer1_outputs(2125));
    layer2_outputs(9216) <= not(layer1_outputs(5225));
    layer2_outputs(9217) <= not((layer1_outputs(552)) xor (layer1_outputs(8977)));
    layer2_outputs(9218) <= not(layer1_outputs(6446));
    layer2_outputs(9219) <= not(layer1_outputs(9289)) or (layer1_outputs(6431));
    layer2_outputs(9220) <= layer1_outputs(8078);
    layer2_outputs(9221) <= not(layer1_outputs(1843));
    layer2_outputs(9222) <= not(layer1_outputs(6762));
    layer2_outputs(9223) <= layer1_outputs(8625);
    layer2_outputs(9224) <= not(layer1_outputs(5031));
    layer2_outputs(9225) <= not(layer1_outputs(1407)) or (layer1_outputs(1816));
    layer2_outputs(9226) <= not(layer1_outputs(8873));
    layer2_outputs(9227) <= not(layer1_outputs(7239));
    layer2_outputs(9228) <= not(layer1_outputs(7862));
    layer2_outputs(9229) <= not(layer1_outputs(2224)) or (layer1_outputs(7434));
    layer2_outputs(9230) <= not(layer1_outputs(7746));
    layer2_outputs(9231) <= (layer1_outputs(2120)) and (layer1_outputs(1135));
    layer2_outputs(9232) <= not(layer1_outputs(4083)) or (layer1_outputs(6129));
    layer2_outputs(9233) <= not(layer1_outputs(9822));
    layer2_outputs(9234) <= not(layer1_outputs(3716));
    layer2_outputs(9235) <= not(layer1_outputs(3436)) or (layer1_outputs(2503));
    layer2_outputs(9236) <= layer1_outputs(7780);
    layer2_outputs(9237) <= not(layer1_outputs(3450));
    layer2_outputs(9238) <= not(layer1_outputs(7050)) or (layer1_outputs(4901));
    layer2_outputs(9239) <= not((layer1_outputs(338)) or (layer1_outputs(6450)));
    layer2_outputs(9240) <= not(layer1_outputs(7704)) or (layer1_outputs(9598));
    layer2_outputs(9241) <= not(layer1_outputs(3647)) or (layer1_outputs(2262));
    layer2_outputs(9242) <= layer1_outputs(469);
    layer2_outputs(9243) <= (layer1_outputs(1994)) xor (layer1_outputs(6439));
    layer2_outputs(9244) <= not(layer1_outputs(46)) or (layer1_outputs(272));
    layer2_outputs(9245) <= not(layer1_outputs(5971));
    layer2_outputs(9246) <= (layer1_outputs(9955)) and not (layer1_outputs(8344));
    layer2_outputs(9247) <= not((layer1_outputs(7409)) and (layer1_outputs(4211)));
    layer2_outputs(9248) <= '0';
    layer2_outputs(9249) <= not(layer1_outputs(932));
    layer2_outputs(9250) <= (layer1_outputs(6052)) or (layer1_outputs(3650));
    layer2_outputs(9251) <= (layer1_outputs(4480)) and not (layer1_outputs(2922));
    layer2_outputs(9252) <= layer1_outputs(7512);
    layer2_outputs(9253) <= not((layer1_outputs(2855)) or (layer1_outputs(6246)));
    layer2_outputs(9254) <= not(layer1_outputs(2839));
    layer2_outputs(9255) <= layer1_outputs(9774);
    layer2_outputs(9256) <= (layer1_outputs(91)) and (layer1_outputs(2621));
    layer2_outputs(9257) <= not((layer1_outputs(3231)) and (layer1_outputs(3303)));
    layer2_outputs(9258) <= layer1_outputs(8961);
    layer2_outputs(9259) <= layer1_outputs(760);
    layer2_outputs(9260) <= not(layer1_outputs(8964));
    layer2_outputs(9261) <= not(layer1_outputs(4394)) or (layer1_outputs(9393));
    layer2_outputs(9262) <= layer1_outputs(1788);
    layer2_outputs(9263) <= layer1_outputs(3071);
    layer2_outputs(9264) <= layer1_outputs(9548);
    layer2_outputs(9265) <= layer1_outputs(154);
    layer2_outputs(9266) <= layer1_outputs(10074);
    layer2_outputs(9267) <= not(layer1_outputs(4254));
    layer2_outputs(9268) <= '0';
    layer2_outputs(9269) <= (layer1_outputs(7761)) or (layer1_outputs(3769));
    layer2_outputs(9270) <= (layer1_outputs(1211)) and (layer1_outputs(5750));
    layer2_outputs(9271) <= not((layer1_outputs(8076)) and (layer1_outputs(1306)));
    layer2_outputs(9272) <= layer1_outputs(2425);
    layer2_outputs(9273) <= not(layer1_outputs(2435));
    layer2_outputs(9274) <= not((layer1_outputs(4570)) xor (layer1_outputs(8250)));
    layer2_outputs(9275) <= '0';
    layer2_outputs(9276) <= not(layer1_outputs(6687)) or (layer1_outputs(9966));
    layer2_outputs(9277) <= not(layer1_outputs(5597));
    layer2_outputs(9278) <= not(layer1_outputs(5888)) or (layer1_outputs(1359));
    layer2_outputs(9279) <= layer1_outputs(9968);
    layer2_outputs(9280) <= (layer1_outputs(5819)) and not (layer1_outputs(1504));
    layer2_outputs(9281) <= layer1_outputs(1320);
    layer2_outputs(9282) <= not((layer1_outputs(7393)) xor (layer1_outputs(9468)));
    layer2_outputs(9283) <= layer1_outputs(2275);
    layer2_outputs(9284) <= layer1_outputs(4688);
    layer2_outputs(9285) <= (layer1_outputs(3157)) and not (layer1_outputs(4325));
    layer2_outputs(9286) <= not(layer1_outputs(9750)) or (layer1_outputs(9521));
    layer2_outputs(9287) <= '0';
    layer2_outputs(9288) <= not(layer1_outputs(4069));
    layer2_outputs(9289) <= layer1_outputs(9947);
    layer2_outputs(9290) <= (layer1_outputs(1022)) and (layer1_outputs(2001));
    layer2_outputs(9291) <= not(layer1_outputs(2597)) or (layer1_outputs(2498));
    layer2_outputs(9292) <= layer1_outputs(5437);
    layer2_outputs(9293) <= not(layer1_outputs(1993)) or (layer1_outputs(9787));
    layer2_outputs(9294) <= layer1_outputs(346);
    layer2_outputs(9295) <= layer1_outputs(5678);
    layer2_outputs(9296) <= layer1_outputs(9567);
    layer2_outputs(9297) <= not(layer1_outputs(522));
    layer2_outputs(9298) <= layer1_outputs(1330);
    layer2_outputs(9299) <= not(layer1_outputs(8708));
    layer2_outputs(9300) <= layer1_outputs(3667);
    layer2_outputs(9301) <= not(layer1_outputs(3126)) or (layer1_outputs(8945));
    layer2_outputs(9302) <= not(layer1_outputs(6673));
    layer2_outputs(9303) <= (layer1_outputs(4407)) or (layer1_outputs(2516));
    layer2_outputs(9304) <= not(layer1_outputs(7983)) or (layer1_outputs(5242));
    layer2_outputs(9305) <= not((layer1_outputs(9756)) and (layer1_outputs(8390)));
    layer2_outputs(9306) <= not((layer1_outputs(6347)) and (layer1_outputs(2494)));
    layer2_outputs(9307) <= not(layer1_outputs(6316));
    layer2_outputs(9308) <= (layer1_outputs(1716)) and not (layer1_outputs(2464));
    layer2_outputs(9309) <= not(layer1_outputs(3841));
    layer2_outputs(9310) <= (layer1_outputs(8401)) xor (layer1_outputs(1895));
    layer2_outputs(9311) <= not(layer1_outputs(5258)) or (layer1_outputs(7063));
    layer2_outputs(9312) <= not(layer1_outputs(7883));
    layer2_outputs(9313) <= not(layer1_outputs(6558)) or (layer1_outputs(6457));
    layer2_outputs(9314) <= (layer1_outputs(7570)) or (layer1_outputs(9909));
    layer2_outputs(9315) <= (layer1_outputs(8794)) or (layer1_outputs(6997));
    layer2_outputs(9316) <= layer1_outputs(5734);
    layer2_outputs(9317) <= (layer1_outputs(4529)) and (layer1_outputs(626));
    layer2_outputs(9318) <= not(layer1_outputs(2037));
    layer2_outputs(9319) <= layer1_outputs(7162);
    layer2_outputs(9320) <= not(layer1_outputs(8713)) or (layer1_outputs(6308));
    layer2_outputs(9321) <= not(layer1_outputs(9952));
    layer2_outputs(9322) <= (layer1_outputs(4685)) xor (layer1_outputs(915));
    layer2_outputs(9323) <= (layer1_outputs(9858)) and not (layer1_outputs(9223));
    layer2_outputs(9324) <= not(layer1_outputs(5513));
    layer2_outputs(9325) <= not(layer1_outputs(6806)) or (layer1_outputs(4188));
    layer2_outputs(9326) <= not(layer1_outputs(8611));
    layer2_outputs(9327) <= layer1_outputs(9881);
    layer2_outputs(9328) <= (layer1_outputs(1454)) and not (layer1_outputs(10100));
    layer2_outputs(9329) <= (layer1_outputs(8509)) and not (layer1_outputs(416));
    layer2_outputs(9330) <= (layer1_outputs(7062)) and not (layer1_outputs(9293));
    layer2_outputs(9331) <= layer1_outputs(6284);
    layer2_outputs(9332) <= layer1_outputs(7511);
    layer2_outputs(9333) <= layer1_outputs(2458);
    layer2_outputs(9334) <= (layer1_outputs(7071)) and not (layer1_outputs(8939));
    layer2_outputs(9335) <= (layer1_outputs(8113)) or (layer1_outputs(8508));
    layer2_outputs(9336) <= '0';
    layer2_outputs(9337) <= layer1_outputs(2715);
    layer2_outputs(9338) <= not((layer1_outputs(9423)) or (layer1_outputs(7614)));
    layer2_outputs(9339) <= not(layer1_outputs(4437));
    layer2_outputs(9340) <= not(layer1_outputs(3016));
    layer2_outputs(9341) <= not(layer1_outputs(7968)) or (layer1_outputs(9210));
    layer2_outputs(9342) <= not(layer1_outputs(3007));
    layer2_outputs(9343) <= (layer1_outputs(8966)) or (layer1_outputs(1105));
    layer2_outputs(9344) <= '0';
    layer2_outputs(9345) <= (layer1_outputs(3165)) or (layer1_outputs(3704));
    layer2_outputs(9346) <= not(layer1_outputs(5833));
    layer2_outputs(9347) <= not(layer1_outputs(3830));
    layer2_outputs(9348) <= not(layer1_outputs(9363)) or (layer1_outputs(4945));
    layer2_outputs(9349) <= not((layer1_outputs(8950)) xor (layer1_outputs(3413)));
    layer2_outputs(9350) <= not((layer1_outputs(5795)) xor (layer1_outputs(9072)));
    layer2_outputs(9351) <= (layer1_outputs(4229)) or (layer1_outputs(4429));
    layer2_outputs(9352) <= not((layer1_outputs(443)) and (layer1_outputs(8586)));
    layer2_outputs(9353) <= not((layer1_outputs(5953)) xor (layer1_outputs(7552)));
    layer2_outputs(9354) <= not(layer1_outputs(679));
    layer2_outputs(9355) <= (layer1_outputs(1761)) and not (layer1_outputs(2561));
    layer2_outputs(9356) <= not((layer1_outputs(7663)) or (layer1_outputs(10002)));
    layer2_outputs(9357) <= (layer1_outputs(9530)) and not (layer1_outputs(8769));
    layer2_outputs(9358) <= (layer1_outputs(4649)) xor (layer1_outputs(6662));
    layer2_outputs(9359) <= layer1_outputs(10068);
    layer2_outputs(9360) <= not(layer1_outputs(1551)) or (layer1_outputs(7205));
    layer2_outputs(9361) <= '0';
    layer2_outputs(9362) <= not(layer1_outputs(9086));
    layer2_outputs(9363) <= not((layer1_outputs(2686)) and (layer1_outputs(2654)));
    layer2_outputs(9364) <= not(layer1_outputs(2954)) or (layer1_outputs(655));
    layer2_outputs(9365) <= not(layer1_outputs(8693));
    layer2_outputs(9366) <= not((layer1_outputs(5466)) and (layer1_outputs(761)));
    layer2_outputs(9367) <= layer1_outputs(3509);
    layer2_outputs(9368) <= layer1_outputs(5218);
    layer2_outputs(9369) <= layer1_outputs(3467);
    layer2_outputs(9370) <= layer1_outputs(7999);
    layer2_outputs(9371) <= layer1_outputs(2314);
    layer2_outputs(9372) <= layer1_outputs(7665);
    layer2_outputs(9373) <= not(layer1_outputs(6440)) or (layer1_outputs(4249));
    layer2_outputs(9374) <= '0';
    layer2_outputs(9375) <= '0';
    layer2_outputs(9376) <= not(layer1_outputs(8546));
    layer2_outputs(9377) <= not(layer1_outputs(2710)) or (layer1_outputs(1025));
    layer2_outputs(9378) <= layer1_outputs(3589);
    layer2_outputs(9379) <= not(layer1_outputs(8226));
    layer2_outputs(9380) <= (layer1_outputs(6321)) and (layer1_outputs(794));
    layer2_outputs(9381) <= not(layer1_outputs(5203)) or (layer1_outputs(5762));
    layer2_outputs(9382) <= not((layer1_outputs(5876)) and (layer1_outputs(8811)));
    layer2_outputs(9383) <= layer1_outputs(4378);
    layer2_outputs(9384) <= not((layer1_outputs(243)) and (layer1_outputs(342)));
    layer2_outputs(9385) <= not(layer1_outputs(2513));
    layer2_outputs(9386) <= not((layer1_outputs(10232)) and (layer1_outputs(3930)));
    layer2_outputs(9387) <= not(layer1_outputs(8331));
    layer2_outputs(9388) <= (layer1_outputs(9835)) and not (layer1_outputs(3594));
    layer2_outputs(9389) <= layer1_outputs(4530);
    layer2_outputs(9390) <= layer1_outputs(2617);
    layer2_outputs(9391) <= not((layer1_outputs(7390)) and (layer1_outputs(6350)));
    layer2_outputs(9392) <= (layer1_outputs(6732)) and not (layer1_outputs(5004));
    layer2_outputs(9393) <= '1';
    layer2_outputs(9394) <= not(layer1_outputs(9923)) or (layer1_outputs(3619));
    layer2_outputs(9395) <= (layer1_outputs(3627)) and not (layer1_outputs(2795));
    layer2_outputs(9396) <= layer1_outputs(5316);
    layer2_outputs(9397) <= not((layer1_outputs(4196)) xor (layer1_outputs(2641)));
    layer2_outputs(9398) <= layer1_outputs(305);
    layer2_outputs(9399) <= (layer1_outputs(2101)) and not (layer1_outputs(8364));
    layer2_outputs(9400) <= layer1_outputs(8445);
    layer2_outputs(9401) <= layer1_outputs(2371);
    layer2_outputs(9402) <= layer1_outputs(2386);
    layer2_outputs(9403) <= (layer1_outputs(183)) xor (layer1_outputs(6130));
    layer2_outputs(9404) <= not(layer1_outputs(2812));
    layer2_outputs(9405) <= layer1_outputs(8582);
    layer2_outputs(9406) <= not(layer1_outputs(6848));
    layer2_outputs(9407) <= not(layer1_outputs(9820)) or (layer1_outputs(3047));
    layer2_outputs(9408) <= layer1_outputs(5484);
    layer2_outputs(9409) <= not(layer1_outputs(2890));
    layer2_outputs(9410) <= (layer1_outputs(920)) and (layer1_outputs(8795));
    layer2_outputs(9411) <= layer1_outputs(248);
    layer2_outputs(9412) <= not(layer1_outputs(8739));
    layer2_outputs(9413) <= not(layer1_outputs(3096));
    layer2_outputs(9414) <= (layer1_outputs(2214)) and not (layer1_outputs(6919));
    layer2_outputs(9415) <= not(layer1_outputs(9279));
    layer2_outputs(9416) <= layer1_outputs(5648);
    layer2_outputs(9417) <= not((layer1_outputs(9367)) or (layer1_outputs(6202)));
    layer2_outputs(9418) <= not(layer1_outputs(2323));
    layer2_outputs(9419) <= not(layer1_outputs(4309));
    layer2_outputs(9420) <= (layer1_outputs(7391)) and (layer1_outputs(7456));
    layer2_outputs(9421) <= layer1_outputs(5948);
    layer2_outputs(9422) <= not(layer1_outputs(5943)) or (layer1_outputs(6394));
    layer2_outputs(9423) <= layer1_outputs(2546);
    layer2_outputs(9424) <= layer1_outputs(2931);
    layer2_outputs(9425) <= layer1_outputs(248);
    layer2_outputs(9426) <= layer1_outputs(1458);
    layer2_outputs(9427) <= (layer1_outputs(5275)) and not (layer1_outputs(1115));
    layer2_outputs(9428) <= not(layer1_outputs(10069)) or (layer1_outputs(780));
    layer2_outputs(9429) <= (layer1_outputs(6802)) or (layer1_outputs(7308));
    layer2_outputs(9430) <= not(layer1_outputs(5963)) or (layer1_outputs(7672));
    layer2_outputs(9431) <= layer1_outputs(6580);
    layer2_outputs(9432) <= not(layer1_outputs(7872)) or (layer1_outputs(4111));
    layer2_outputs(9433) <= layer1_outputs(3597);
    layer2_outputs(9434) <= (layer1_outputs(9843)) or (layer1_outputs(2324));
    layer2_outputs(9435) <= layer1_outputs(4643);
    layer2_outputs(9436) <= not((layer1_outputs(2211)) or (layer1_outputs(8295)));
    layer2_outputs(9437) <= not(layer1_outputs(754));
    layer2_outputs(9438) <= not(layer1_outputs(8617));
    layer2_outputs(9439) <= not(layer1_outputs(322));
    layer2_outputs(9440) <= layer1_outputs(444);
    layer2_outputs(9441) <= (layer1_outputs(516)) and (layer1_outputs(3681));
    layer2_outputs(9442) <= (layer1_outputs(6594)) or (layer1_outputs(2478));
    layer2_outputs(9443) <= (layer1_outputs(4833)) and not (layer1_outputs(10015));
    layer2_outputs(9444) <= layer1_outputs(545);
    layer2_outputs(9445) <= layer1_outputs(5170);
    layer2_outputs(9446) <= not(layer1_outputs(1629)) or (layer1_outputs(6627));
    layer2_outputs(9447) <= not(layer1_outputs(5085));
    layer2_outputs(9448) <= not(layer1_outputs(2742)) or (layer1_outputs(9954));
    layer2_outputs(9449) <= not((layer1_outputs(5368)) and (layer1_outputs(8080)));
    layer2_outputs(9450) <= layer1_outputs(2836);
    layer2_outputs(9451) <= layer1_outputs(6428);
    layer2_outputs(9452) <= not((layer1_outputs(2326)) and (layer1_outputs(2064)));
    layer2_outputs(9453) <= (layer1_outputs(9138)) or (layer1_outputs(4402));
    layer2_outputs(9454) <= not(layer1_outputs(2771));
    layer2_outputs(9455) <= not(layer1_outputs(7645));
    layer2_outputs(9456) <= (layer1_outputs(5736)) or (layer1_outputs(3946));
    layer2_outputs(9457) <= not((layer1_outputs(4059)) xor (layer1_outputs(10168)));
    layer2_outputs(9458) <= layer1_outputs(3082);
    layer2_outputs(9459) <= (layer1_outputs(10129)) and not (layer1_outputs(5950));
    layer2_outputs(9460) <= '1';
    layer2_outputs(9461) <= layer1_outputs(8777);
    layer2_outputs(9462) <= layer1_outputs(8466);
    layer2_outputs(9463) <= not(layer1_outputs(3533));
    layer2_outputs(9464) <= (layer1_outputs(7741)) and not (layer1_outputs(1933));
    layer2_outputs(9465) <= '1';
    layer2_outputs(9466) <= (layer1_outputs(790)) xor (layer1_outputs(3842));
    layer2_outputs(9467) <= not(layer1_outputs(2052));
    layer2_outputs(9468) <= (layer1_outputs(803)) or (layer1_outputs(3005));
    layer2_outputs(9469) <= not((layer1_outputs(5830)) and (layer1_outputs(333)));
    layer2_outputs(9470) <= not(layer1_outputs(2076)) or (layer1_outputs(8135));
    layer2_outputs(9471) <= '0';
    layer2_outputs(9472) <= layer1_outputs(7881);
    layer2_outputs(9473) <= not(layer1_outputs(7778)) or (layer1_outputs(7073));
    layer2_outputs(9474) <= layer1_outputs(1998);
    layer2_outputs(9475) <= not(layer1_outputs(9482));
    layer2_outputs(9476) <= layer1_outputs(9697);
    layer2_outputs(9477) <= not(layer1_outputs(5156)) or (layer1_outputs(3872));
    layer2_outputs(9478) <= not(layer1_outputs(6638));
    layer2_outputs(9479) <= (layer1_outputs(2922)) and (layer1_outputs(221));
    layer2_outputs(9480) <= not(layer1_outputs(658));
    layer2_outputs(9481) <= not(layer1_outputs(4987)) or (layer1_outputs(4396));
    layer2_outputs(9482) <= not(layer1_outputs(1619)) or (layer1_outputs(4084));
    layer2_outputs(9483) <= (layer1_outputs(2219)) and (layer1_outputs(10172));
    layer2_outputs(9484) <= (layer1_outputs(6712)) xor (layer1_outputs(197));
    layer2_outputs(9485) <= not(layer1_outputs(6900));
    layer2_outputs(9486) <= (layer1_outputs(7135)) and not (layer1_outputs(9159));
    layer2_outputs(9487) <= not(layer1_outputs(7339)) or (layer1_outputs(8286));
    layer2_outputs(9488) <= layer1_outputs(307);
    layer2_outputs(9489) <= not(layer1_outputs(9026)) or (layer1_outputs(5734));
    layer2_outputs(9490) <= not(layer1_outputs(164)) or (layer1_outputs(5387));
    layer2_outputs(9491) <= not((layer1_outputs(6857)) or (layer1_outputs(7173)));
    layer2_outputs(9492) <= not(layer1_outputs(7740)) or (layer1_outputs(2624));
    layer2_outputs(9493) <= layer1_outputs(8537);
    layer2_outputs(9494) <= (layer1_outputs(2126)) or (layer1_outputs(2157));
    layer2_outputs(9495) <= (layer1_outputs(4657)) xor (layer1_outputs(8958));
    layer2_outputs(9496) <= layer1_outputs(5105);
    layer2_outputs(9497) <= not(layer1_outputs(993));
    layer2_outputs(9498) <= not(layer1_outputs(287)) or (layer1_outputs(2726));
    layer2_outputs(9499) <= not((layer1_outputs(9027)) and (layer1_outputs(7884)));
    layer2_outputs(9500) <= not((layer1_outputs(311)) and (layer1_outputs(6765)));
    layer2_outputs(9501) <= not(layer1_outputs(9638));
    layer2_outputs(9502) <= (layer1_outputs(8251)) or (layer1_outputs(7589));
    layer2_outputs(9503) <= not(layer1_outputs(6101));
    layer2_outputs(9504) <= not(layer1_outputs(4605));
    layer2_outputs(9505) <= not(layer1_outputs(6740));
    layer2_outputs(9506) <= not((layer1_outputs(10003)) or (layer1_outputs(3410)));
    layer2_outputs(9507) <= not((layer1_outputs(5083)) and (layer1_outputs(8384)));
    layer2_outputs(9508) <= (layer1_outputs(1564)) and not (layer1_outputs(7411));
    layer2_outputs(9509) <= layer1_outputs(424);
    layer2_outputs(9510) <= layer1_outputs(10085);
    layer2_outputs(9511) <= not((layer1_outputs(3516)) and (layer1_outputs(7559)));
    layer2_outputs(9512) <= (layer1_outputs(5110)) and (layer1_outputs(9270));
    layer2_outputs(9513) <= (layer1_outputs(6359)) and not (layer1_outputs(9977));
    layer2_outputs(9514) <= not(layer1_outputs(6729));
    layer2_outputs(9515) <= not((layer1_outputs(8131)) xor (layer1_outputs(4476)));
    layer2_outputs(9516) <= (layer1_outputs(2927)) and not (layer1_outputs(3824));
    layer2_outputs(9517) <= not((layer1_outputs(371)) or (layer1_outputs(6547)));
    layer2_outputs(9518) <= not((layer1_outputs(1074)) and (layer1_outputs(10210)));
    layer2_outputs(9519) <= (layer1_outputs(8325)) and (layer1_outputs(4166));
    layer2_outputs(9520) <= not(layer1_outputs(3929)) or (layer1_outputs(8621));
    layer2_outputs(9521) <= not(layer1_outputs(48));
    layer2_outputs(9522) <= (layer1_outputs(9093)) or (layer1_outputs(2991));
    layer2_outputs(9523) <= not((layer1_outputs(6055)) and (layer1_outputs(9435)));
    layer2_outputs(9524) <= not(layer1_outputs(2927));
    layer2_outputs(9525) <= not((layer1_outputs(9975)) or (layer1_outputs(7461)));
    layer2_outputs(9526) <= layer1_outputs(7338);
    layer2_outputs(9527) <= not(layer1_outputs(2395));
    layer2_outputs(9528) <= not((layer1_outputs(526)) or (layer1_outputs(12)));
    layer2_outputs(9529) <= (layer1_outputs(9775)) and (layer1_outputs(6817));
    layer2_outputs(9530) <= layer1_outputs(1232);
    layer2_outputs(9531) <= (layer1_outputs(9635)) or (layer1_outputs(10029));
    layer2_outputs(9532) <= (layer1_outputs(4636)) xor (layer1_outputs(6892));
    layer2_outputs(9533) <= (layer1_outputs(5145)) and not (layer1_outputs(5064));
    layer2_outputs(9534) <= (layer1_outputs(6704)) xor (layer1_outputs(9330));
    layer2_outputs(9535) <= (layer1_outputs(6903)) and (layer1_outputs(7628));
    layer2_outputs(9536) <= not(layer1_outputs(9061)) or (layer1_outputs(847));
    layer2_outputs(9537) <= not((layer1_outputs(7755)) and (layer1_outputs(8370)));
    layer2_outputs(9538) <= layer1_outputs(8163);
    layer2_outputs(9539) <= not((layer1_outputs(1659)) or (layer1_outputs(4167)));
    layer2_outputs(9540) <= not(layer1_outputs(4486));
    layer2_outputs(9541) <= layer1_outputs(2788);
    layer2_outputs(9542) <= not((layer1_outputs(7571)) or (layer1_outputs(3936)));
    layer2_outputs(9543) <= layer1_outputs(3902);
    layer2_outputs(9544) <= not(layer1_outputs(8283));
    layer2_outputs(9545) <= layer1_outputs(919);
    layer2_outputs(9546) <= '1';
    layer2_outputs(9547) <= not(layer1_outputs(7346));
    layer2_outputs(9548) <= (layer1_outputs(1971)) and not (layer1_outputs(3457));
    layer2_outputs(9549) <= not(layer1_outputs(9278));
    layer2_outputs(9550) <= layer1_outputs(479);
    layer2_outputs(9551) <= not((layer1_outputs(9189)) xor (layer1_outputs(9561)));
    layer2_outputs(9552) <= (layer1_outputs(280)) and not (layer1_outputs(9947));
    layer2_outputs(9553) <= not(layer1_outputs(3880));
    layer2_outputs(9554) <= layer1_outputs(126);
    layer2_outputs(9555) <= (layer1_outputs(5722)) and not (layer1_outputs(8705));
    layer2_outputs(9556) <= not(layer1_outputs(6823)) or (layer1_outputs(4322));
    layer2_outputs(9557) <= not(layer1_outputs(2599));
    layer2_outputs(9558) <= layer1_outputs(2335);
    layer2_outputs(9559) <= not((layer1_outputs(361)) xor (layer1_outputs(7991)));
    layer2_outputs(9560) <= (layer1_outputs(1366)) and not (layer1_outputs(10093));
    layer2_outputs(9561) <= layer1_outputs(6123);
    layer2_outputs(9562) <= layer1_outputs(1198);
    layer2_outputs(9563) <= '1';
    layer2_outputs(9564) <= not(layer1_outputs(2651)) or (layer1_outputs(10057));
    layer2_outputs(9565) <= not((layer1_outputs(3728)) or (layer1_outputs(2573)));
    layer2_outputs(9566) <= not(layer1_outputs(5490));
    layer2_outputs(9567) <= layer1_outputs(10230);
    layer2_outputs(9568) <= (layer1_outputs(6885)) and (layer1_outputs(3536));
    layer2_outputs(9569) <= not((layer1_outputs(8186)) and (layer1_outputs(143)));
    layer2_outputs(9570) <= (layer1_outputs(5339)) or (layer1_outputs(9250));
    layer2_outputs(9571) <= (layer1_outputs(722)) or (layer1_outputs(8086));
    layer2_outputs(9572) <= (layer1_outputs(4650)) and not (layer1_outputs(1286));
    layer2_outputs(9573) <= not(layer1_outputs(6471));
    layer2_outputs(9574) <= layer1_outputs(718);
    layer2_outputs(9575) <= layer1_outputs(8593);
    layer2_outputs(9576) <= not((layer1_outputs(1572)) xor (layer1_outputs(3149)));
    layer2_outputs(9577) <= not((layer1_outputs(4222)) xor (layer1_outputs(3336)));
    layer2_outputs(9578) <= '1';
    layer2_outputs(9579) <= (layer1_outputs(2061)) and (layer1_outputs(7437));
    layer2_outputs(9580) <= not(layer1_outputs(4557)) or (layer1_outputs(149));
    layer2_outputs(9581) <= layer1_outputs(8849);
    layer2_outputs(9582) <= (layer1_outputs(9737)) and not (layer1_outputs(7678));
    layer2_outputs(9583) <= layer1_outputs(9924);
    layer2_outputs(9584) <= (layer1_outputs(7546)) and not (layer1_outputs(9949));
    layer2_outputs(9585) <= not((layer1_outputs(7277)) or (layer1_outputs(3918)));
    layer2_outputs(9586) <= not((layer1_outputs(2365)) or (layer1_outputs(5703)));
    layer2_outputs(9587) <= not((layer1_outputs(42)) xor (layer1_outputs(9231)));
    layer2_outputs(9588) <= layer1_outputs(5459);
    layer2_outputs(9589) <= (layer1_outputs(4970)) or (layer1_outputs(1360));
    layer2_outputs(9590) <= '1';
    layer2_outputs(9591) <= not(layer1_outputs(1645)) or (layer1_outputs(1824));
    layer2_outputs(9592) <= (layer1_outputs(6157)) and not (layer1_outputs(2418));
    layer2_outputs(9593) <= (layer1_outputs(6059)) or (layer1_outputs(7910));
    layer2_outputs(9594) <= not(layer1_outputs(7403)) or (layer1_outputs(5221));
    layer2_outputs(9595) <= '1';
    layer2_outputs(9596) <= (layer1_outputs(6587)) or (layer1_outputs(2910));
    layer2_outputs(9597) <= not((layer1_outputs(478)) xor (layer1_outputs(8756)));
    layer2_outputs(9598) <= layer1_outputs(1110);
    layer2_outputs(9599) <= not(layer1_outputs(6860));
    layer2_outputs(9600) <= layer1_outputs(551);
    layer2_outputs(9601) <= not((layer1_outputs(9794)) xor (layer1_outputs(10176)));
    layer2_outputs(9602) <= layer1_outputs(5860);
    layer2_outputs(9603) <= not((layer1_outputs(2383)) and (layer1_outputs(855)));
    layer2_outputs(9604) <= not(layer1_outputs(2298)) or (layer1_outputs(987));
    layer2_outputs(9605) <= layer1_outputs(5120);
    layer2_outputs(9606) <= (layer1_outputs(1571)) and (layer1_outputs(2666));
    layer2_outputs(9607) <= '0';
    layer2_outputs(9608) <= layer1_outputs(10137);
    layer2_outputs(9609) <= (layer1_outputs(1003)) or (layer1_outputs(5288));
    layer2_outputs(9610) <= layer1_outputs(3045);
    layer2_outputs(9611) <= not((layer1_outputs(1484)) or (layer1_outputs(6603)));
    layer2_outputs(9612) <= (layer1_outputs(9633)) or (layer1_outputs(8374));
    layer2_outputs(9613) <= layer1_outputs(8379);
    layer2_outputs(9614) <= not((layer1_outputs(4742)) or (layer1_outputs(1880)));
    layer2_outputs(9615) <= (layer1_outputs(6842)) and not (layer1_outputs(3322));
    layer2_outputs(9616) <= not((layer1_outputs(6716)) or (layer1_outputs(5013)));
    layer2_outputs(9617) <= not((layer1_outputs(9165)) xor (layer1_outputs(9417)));
    layer2_outputs(9618) <= not((layer1_outputs(3431)) xor (layer1_outputs(1476)));
    layer2_outputs(9619) <= not(layer1_outputs(202));
    layer2_outputs(9620) <= not(layer1_outputs(6930));
    layer2_outputs(9621) <= not(layer1_outputs(863));
    layer2_outputs(9622) <= (layer1_outputs(9085)) or (layer1_outputs(2710));
    layer2_outputs(9623) <= not((layer1_outputs(6192)) or (layer1_outputs(8726)));
    layer2_outputs(9624) <= not(layer1_outputs(1804));
    layer2_outputs(9625) <= (layer1_outputs(473)) xor (layer1_outputs(1260));
    layer2_outputs(9626) <= not((layer1_outputs(2724)) or (layer1_outputs(10140)));
    layer2_outputs(9627) <= (layer1_outputs(1660)) xor (layer1_outputs(8056));
    layer2_outputs(9628) <= layer1_outputs(7900);
    layer2_outputs(9629) <= layer1_outputs(9577);
    layer2_outputs(9630) <= layer1_outputs(471);
    layer2_outputs(9631) <= not(layer1_outputs(1402)) or (layer1_outputs(8731));
    layer2_outputs(9632) <= (layer1_outputs(3094)) and not (layer1_outputs(2974));
    layer2_outputs(9633) <= layer1_outputs(10142);
    layer2_outputs(9634) <= (layer1_outputs(4730)) and not (layer1_outputs(5389));
    layer2_outputs(9635) <= '1';
    layer2_outputs(9636) <= not((layer1_outputs(5320)) xor (layer1_outputs(5946)));
    layer2_outputs(9637) <= not(layer1_outputs(5291));
    layer2_outputs(9638) <= (layer1_outputs(3224)) or (layer1_outputs(2520));
    layer2_outputs(9639) <= (layer1_outputs(8520)) and (layer1_outputs(55));
    layer2_outputs(9640) <= not(layer1_outputs(7141)) or (layer1_outputs(6663));
    layer2_outputs(9641) <= (layer1_outputs(6090)) and not (layer1_outputs(7417));
    layer2_outputs(9642) <= '0';
    layer2_outputs(9643) <= (layer1_outputs(5096)) xor (layer1_outputs(7193));
    layer2_outputs(9644) <= layer1_outputs(8618);
    layer2_outputs(9645) <= not(layer1_outputs(9436));
    layer2_outputs(9646) <= not(layer1_outputs(1788));
    layer2_outputs(9647) <= (layer1_outputs(6685)) and not (layer1_outputs(5949));
    layer2_outputs(9648) <= (layer1_outputs(8962)) and not (layer1_outputs(2124));
    layer2_outputs(9649) <= layer1_outputs(10224);
    layer2_outputs(9650) <= not(layer1_outputs(7796));
    layer2_outputs(9651) <= (layer1_outputs(3023)) and not (layer1_outputs(9276));
    layer2_outputs(9652) <= not(layer1_outputs(7039)) or (layer1_outputs(2122));
    layer2_outputs(9653) <= (layer1_outputs(2735)) and not (layer1_outputs(3511));
    layer2_outputs(9654) <= (layer1_outputs(1558)) and not (layer1_outputs(9466));
    layer2_outputs(9655) <= not(layer1_outputs(3624));
    layer2_outputs(9656) <= '0';
    layer2_outputs(9657) <= not((layer1_outputs(136)) or (layer1_outputs(4369)));
    layer2_outputs(9658) <= not(layer1_outputs(1867));
    layer2_outputs(9659) <= (layer1_outputs(6280)) or (layer1_outputs(489));
    layer2_outputs(9660) <= layer1_outputs(2769);
    layer2_outputs(9661) <= not((layer1_outputs(1008)) or (layer1_outputs(4757)));
    layer2_outputs(9662) <= '0';
    layer2_outputs(9663) <= (layer1_outputs(8720)) and not (layer1_outputs(1444));
    layer2_outputs(9664) <= not(layer1_outputs(27)) or (layer1_outputs(129));
    layer2_outputs(9665) <= (layer1_outputs(8553)) and not (layer1_outputs(3484));
    layer2_outputs(9666) <= not((layer1_outputs(6955)) and (layer1_outputs(1040)));
    layer2_outputs(9667) <= not(layer1_outputs(9770)) or (layer1_outputs(3720));
    layer2_outputs(9668) <= not(layer1_outputs(1798)) or (layer1_outputs(9712));
    layer2_outputs(9669) <= not(layer1_outputs(4672));
    layer2_outputs(9670) <= '0';
    layer2_outputs(9671) <= layer1_outputs(9790);
    layer2_outputs(9672) <= not(layer1_outputs(5696));
    layer2_outputs(9673) <= not(layer1_outputs(8604));
    layer2_outputs(9674) <= not(layer1_outputs(979));
    layer2_outputs(9675) <= layer1_outputs(3957);
    layer2_outputs(9676) <= (layer1_outputs(9679)) and not (layer1_outputs(8723));
    layer2_outputs(9677) <= layer1_outputs(1985);
    layer2_outputs(9678) <= (layer1_outputs(6207)) and (layer1_outputs(1424));
    layer2_outputs(9679) <= layer1_outputs(7459);
    layer2_outputs(9680) <= not(layer1_outputs(3319));
    layer2_outputs(9681) <= not(layer1_outputs(8827));
    layer2_outputs(9682) <= (layer1_outputs(297)) and not (layer1_outputs(318));
    layer2_outputs(9683) <= (layer1_outputs(5659)) or (layer1_outputs(1743));
    layer2_outputs(9684) <= not(layer1_outputs(4062)) or (layer1_outputs(2478));
    layer2_outputs(9685) <= (layer1_outputs(1854)) xor (layer1_outputs(4197));
    layer2_outputs(9686) <= not(layer1_outputs(9358));
    layer2_outputs(9687) <= (layer1_outputs(2781)) and not (layer1_outputs(8415));
    layer2_outputs(9688) <= (layer1_outputs(4938)) and not (layer1_outputs(9386));
    layer2_outputs(9689) <= not(layer1_outputs(7500));
    layer2_outputs(9690) <= layer1_outputs(2770);
    layer2_outputs(9691) <= (layer1_outputs(5167)) and (layer1_outputs(929));
    layer2_outputs(9692) <= layer1_outputs(8107);
    layer2_outputs(9693) <= (layer1_outputs(7368)) xor (layer1_outputs(7479));
    layer2_outputs(9694) <= not(layer1_outputs(1207));
    layer2_outputs(9695) <= not((layer1_outputs(7022)) or (layer1_outputs(5825)));
    layer2_outputs(9696) <= (layer1_outputs(7588)) and (layer1_outputs(6726));
    layer2_outputs(9697) <= layer1_outputs(1266);
    layer2_outputs(9698) <= not(layer1_outputs(8770)) or (layer1_outputs(3969));
    layer2_outputs(9699) <= layer1_outputs(10060);
    layer2_outputs(9700) <= (layer1_outputs(7084)) xor (layer1_outputs(7881));
    layer2_outputs(9701) <= (layer1_outputs(7806)) and (layer1_outputs(6309));
    layer2_outputs(9702) <= not(layer1_outputs(4600)) or (layer1_outputs(8447));
    layer2_outputs(9703) <= (layer1_outputs(8042)) and (layer1_outputs(9845));
    layer2_outputs(9704) <= not(layer1_outputs(6788)) or (layer1_outputs(3577));
    layer2_outputs(9705) <= not(layer1_outputs(1776));
    layer2_outputs(9706) <= layer1_outputs(944);
    layer2_outputs(9707) <= (layer1_outputs(1269)) and (layer1_outputs(7518));
    layer2_outputs(9708) <= not((layer1_outputs(2996)) or (layer1_outputs(9549)));
    layer2_outputs(9709) <= layer1_outputs(3710);
    layer2_outputs(9710) <= (layer1_outputs(6401)) xor (layer1_outputs(9227));
    layer2_outputs(9711) <= not(layer1_outputs(8822)) or (layer1_outputs(1546));
    layer2_outputs(9712) <= layer1_outputs(4588);
    layer2_outputs(9713) <= not((layer1_outputs(3725)) or (layer1_outputs(1533)));
    layer2_outputs(9714) <= not(layer1_outputs(6677));
    layer2_outputs(9715) <= (layer1_outputs(4250)) or (layer1_outputs(4687));
    layer2_outputs(9716) <= (layer1_outputs(4562)) or (layer1_outputs(4800));
    layer2_outputs(9717) <= not(layer1_outputs(7378));
    layer2_outputs(9718) <= layer1_outputs(2002);
    layer2_outputs(9719) <= not((layer1_outputs(7335)) or (layer1_outputs(3747)));
    layer2_outputs(9720) <= layer1_outputs(1862);
    layer2_outputs(9721) <= layer1_outputs(5689);
    layer2_outputs(9722) <= not(layer1_outputs(6586));
    layer2_outputs(9723) <= not(layer1_outputs(8087));
    layer2_outputs(9724) <= not(layer1_outputs(994));
    layer2_outputs(9725) <= not(layer1_outputs(8386));
    layer2_outputs(9726) <= not(layer1_outputs(2607));
    layer2_outputs(9727) <= not((layer1_outputs(1569)) or (layer1_outputs(1832)));
    layer2_outputs(9728) <= not(layer1_outputs(2988)) or (layer1_outputs(5059));
    layer2_outputs(9729) <= not(layer1_outputs(6653));
    layer2_outputs(9730) <= not(layer1_outputs(5245));
    layer2_outputs(9731) <= (layer1_outputs(5312)) or (layer1_outputs(2053));
    layer2_outputs(9732) <= (layer1_outputs(8090)) and not (layer1_outputs(4563));
    layer2_outputs(9733) <= (layer1_outputs(5487)) and not (layer1_outputs(139));
    layer2_outputs(9734) <= (layer1_outputs(5614)) or (layer1_outputs(7334));
    layer2_outputs(9735) <= not(layer1_outputs(5883));
    layer2_outputs(9736) <= (layer1_outputs(224)) and not (layer1_outputs(5844));
    layer2_outputs(9737) <= not(layer1_outputs(5348));
    layer2_outputs(9738) <= not(layer1_outputs(7428)) or (layer1_outputs(629));
    layer2_outputs(9739) <= not(layer1_outputs(7749));
    layer2_outputs(9740) <= not(layer1_outputs(646)) or (layer1_outputs(8532));
    layer2_outputs(9741) <= not((layer1_outputs(5620)) or (layer1_outputs(9078)));
    layer2_outputs(9742) <= not(layer1_outputs(9540));
    layer2_outputs(9743) <= not(layer1_outputs(1322));
    layer2_outputs(9744) <= (layer1_outputs(5766)) and not (layer1_outputs(1017));
    layer2_outputs(9745) <= not(layer1_outputs(1521));
    layer2_outputs(9746) <= not(layer1_outputs(296));
    layer2_outputs(9747) <= not(layer1_outputs(4368)) or (layer1_outputs(6825));
    layer2_outputs(9748) <= (layer1_outputs(1631)) and (layer1_outputs(7049));
    layer2_outputs(9749) <= '0';
    layer2_outputs(9750) <= (layer1_outputs(9150)) and not (layer1_outputs(5582));
    layer2_outputs(9751) <= '1';
    layer2_outputs(9752) <= not((layer1_outputs(3886)) or (layer1_outputs(7759)));
    layer2_outputs(9753) <= not(layer1_outputs(8965));
    layer2_outputs(9754) <= not(layer1_outputs(1990)) or (layer1_outputs(2442));
    layer2_outputs(9755) <= (layer1_outputs(4347)) xor (layer1_outputs(1067));
    layer2_outputs(9756) <= '1';
    layer2_outputs(9757) <= (layer1_outputs(7855)) or (layer1_outputs(9144));
    layer2_outputs(9758) <= not(layer1_outputs(7299));
    layer2_outputs(9759) <= layer1_outputs(4286);
    layer2_outputs(9760) <= not(layer1_outputs(6019));
    layer2_outputs(9761) <= (layer1_outputs(6671)) or (layer1_outputs(2978));
    layer2_outputs(9762) <= (layer1_outputs(3139)) and (layer1_outputs(5545));
    layer2_outputs(9763) <= not(layer1_outputs(1737)) or (layer1_outputs(9536));
    layer2_outputs(9764) <= not((layer1_outputs(3891)) and (layer1_outputs(7396)));
    layer2_outputs(9765) <= layer1_outputs(9402);
    layer2_outputs(9766) <= (layer1_outputs(8089)) and not (layer1_outputs(9407));
    layer2_outputs(9767) <= not(layer1_outputs(4934));
    layer2_outputs(9768) <= '1';
    layer2_outputs(9769) <= (layer1_outputs(630)) and not (layer1_outputs(6760));
    layer2_outputs(9770) <= (layer1_outputs(7595)) and not (layer1_outputs(9696));
    layer2_outputs(9771) <= layer1_outputs(4849);
    layer2_outputs(9772) <= (layer1_outputs(4535)) xor (layer1_outputs(4809));
    layer2_outputs(9773) <= (layer1_outputs(2786)) xor (layer1_outputs(254));
    layer2_outputs(9774) <= (layer1_outputs(8005)) and not (layer1_outputs(2912));
    layer2_outputs(9775) <= layer1_outputs(3176);
    layer2_outputs(9776) <= not(layer1_outputs(4448));
    layer2_outputs(9777) <= not(layer1_outputs(1676)) or (layer1_outputs(4018));
    layer2_outputs(9778) <= '0';
    layer2_outputs(9779) <= (layer1_outputs(6178)) and (layer1_outputs(2382));
    layer2_outputs(9780) <= not(layer1_outputs(6228)) or (layer1_outputs(5677));
    layer2_outputs(9781) <= not(layer1_outputs(9106));
    layer2_outputs(9782) <= (layer1_outputs(6914)) xor (layer1_outputs(2815));
    layer2_outputs(9783) <= layer1_outputs(1338);
    layer2_outputs(9784) <= (layer1_outputs(594)) and not (layer1_outputs(337));
    layer2_outputs(9785) <= not(layer1_outputs(6407));
    layer2_outputs(9786) <= (layer1_outputs(2077)) and not (layer1_outputs(6685));
    layer2_outputs(9787) <= (layer1_outputs(3304)) and not (layer1_outputs(9719));
    layer2_outputs(9788) <= layer1_outputs(5672);
    layer2_outputs(9789) <= not(layer1_outputs(7489));
    layer2_outputs(9790) <= '0';
    layer2_outputs(9791) <= (layer1_outputs(7499)) or (layer1_outputs(436));
    layer2_outputs(9792) <= '1';
    layer2_outputs(9793) <= not(layer1_outputs(5974));
    layer2_outputs(9794) <= (layer1_outputs(7930)) and (layer1_outputs(3248));
    layer2_outputs(9795) <= not(layer1_outputs(8359));
    layer2_outputs(9796) <= not(layer1_outputs(4599)) or (layer1_outputs(8396));
    layer2_outputs(9797) <= '1';
    layer2_outputs(9798) <= (layer1_outputs(5544)) xor (layer1_outputs(1082));
    layer2_outputs(9799) <= layer1_outputs(3801);
    layer2_outputs(9800) <= not(layer1_outputs(1665));
    layer2_outputs(9801) <= layer1_outputs(7470);
    layer2_outputs(9802) <= not((layer1_outputs(1559)) and (layer1_outputs(5428)));
    layer2_outputs(9803) <= not(layer1_outputs(2917)) or (layer1_outputs(5131));
    layer2_outputs(9804) <= '0';
    layer2_outputs(9805) <= '0';
    layer2_outputs(9806) <= not((layer1_outputs(1384)) xor (layer1_outputs(2110)));
    layer2_outputs(9807) <= (layer1_outputs(7637)) or (layer1_outputs(1922));
    layer2_outputs(9808) <= not((layer1_outputs(1784)) xor (layer1_outputs(9463)));
    layer2_outputs(9809) <= layer1_outputs(1199);
    layer2_outputs(9810) <= not((layer1_outputs(2377)) and (layer1_outputs(8982)));
    layer2_outputs(9811) <= not(layer1_outputs(8950)) or (layer1_outputs(6897));
    layer2_outputs(9812) <= not((layer1_outputs(5111)) and (layer1_outputs(9572)));
    layer2_outputs(9813) <= not(layer1_outputs(796));
    layer2_outputs(9814) <= not(layer1_outputs(10081));
    layer2_outputs(9815) <= (layer1_outputs(8867)) xor (layer1_outputs(1310));
    layer2_outputs(9816) <= (layer1_outputs(5164)) and not (layer1_outputs(4393));
    layer2_outputs(9817) <= (layer1_outputs(3503)) or (layer1_outputs(9887));
    layer2_outputs(9818) <= not(layer1_outputs(7819));
    layer2_outputs(9819) <= not((layer1_outputs(1497)) xor (layer1_outputs(7904)));
    layer2_outputs(9820) <= (layer1_outputs(8607)) or (layer1_outputs(9042));
    layer2_outputs(9821) <= (layer1_outputs(5954)) and not (layer1_outputs(1890));
    layer2_outputs(9822) <= layer1_outputs(2708);
    layer2_outputs(9823) <= (layer1_outputs(2406)) or (layer1_outputs(9392));
    layer2_outputs(9824) <= (layer1_outputs(7150)) or (layer1_outputs(3276));
    layer2_outputs(9825) <= not(layer1_outputs(9839));
    layer2_outputs(9826) <= layer1_outputs(6793);
    layer2_outputs(9827) <= '1';
    layer2_outputs(9828) <= (layer1_outputs(1631)) and (layer1_outputs(7770));
    layer2_outputs(9829) <= not(layer1_outputs(406)) or (layer1_outputs(4825));
    layer2_outputs(9830) <= not(layer1_outputs(7889));
    layer2_outputs(9831) <= (layer1_outputs(7256)) and not (layer1_outputs(9408));
    layer2_outputs(9832) <= (layer1_outputs(10033)) and not (layer1_outputs(1884));
    layer2_outputs(9833) <= not(layer1_outputs(850));
    layer2_outputs(9834) <= (layer1_outputs(7367)) and (layer1_outputs(5706));
    layer2_outputs(9835) <= not((layer1_outputs(8397)) xor (layer1_outputs(3075)));
    layer2_outputs(9836) <= not(layer1_outputs(6958));
    layer2_outputs(9837) <= layer1_outputs(9882);
    layer2_outputs(9838) <= (layer1_outputs(7436)) xor (layer1_outputs(2277));
    layer2_outputs(9839) <= not(layer1_outputs(2668)) or (layer1_outputs(5857));
    layer2_outputs(9840) <= not(layer1_outputs(8444));
    layer2_outputs(9841) <= not((layer1_outputs(9981)) or (layer1_outputs(213)));
    layer2_outputs(9842) <= layer1_outputs(6022);
    layer2_outputs(9843) <= not(layer1_outputs(1430));
    layer2_outputs(9844) <= (layer1_outputs(5117)) xor (layer1_outputs(9840));
    layer2_outputs(9845) <= not((layer1_outputs(5318)) or (layer1_outputs(1306)));
    layer2_outputs(9846) <= (layer1_outputs(8924)) xor (layer1_outputs(1726));
    layer2_outputs(9847) <= not((layer1_outputs(2639)) or (layer1_outputs(9481)));
    layer2_outputs(9848) <= layer1_outputs(2063);
    layer2_outputs(9849) <= '0';
    layer2_outputs(9850) <= (layer1_outputs(5137)) and not (layer1_outputs(4323));
    layer2_outputs(9851) <= (layer1_outputs(2821)) or (layer1_outputs(7643));
    layer2_outputs(9852) <= layer1_outputs(9447);
    layer2_outputs(9853) <= not(layer1_outputs(3291));
    layer2_outputs(9854) <= not((layer1_outputs(8240)) and (layer1_outputs(7444)));
    layer2_outputs(9855) <= (layer1_outputs(868)) and (layer1_outputs(5386));
    layer2_outputs(9856) <= not(layer1_outputs(423));
    layer2_outputs(9857) <= (layer1_outputs(4735)) and not (layer1_outputs(8925));
    layer2_outputs(9858) <= (layer1_outputs(2591)) xor (layer1_outputs(4524));
    layer2_outputs(9859) <= not((layer1_outputs(468)) or (layer1_outputs(4855)));
    layer2_outputs(9860) <= (layer1_outputs(5042)) and (layer1_outputs(4037));
    layer2_outputs(9861) <= not((layer1_outputs(4877)) and (layer1_outputs(7377)));
    layer2_outputs(9862) <= layer1_outputs(2283);
    layer2_outputs(9863) <= (layer1_outputs(1741)) or (layer1_outputs(5755));
    layer2_outputs(9864) <= not(layer1_outputs(9156));
    layer2_outputs(9865) <= layer1_outputs(7257);
    layer2_outputs(9866) <= (layer1_outputs(411)) and (layer1_outputs(4020));
    layer2_outputs(9867) <= (layer1_outputs(8757)) and not (layer1_outputs(9837));
    layer2_outputs(9868) <= not(layer1_outputs(6023));
    layer2_outputs(9869) <= layer1_outputs(6506);
    layer2_outputs(9870) <= not((layer1_outputs(3712)) xor (layer1_outputs(5517)));
    layer2_outputs(9871) <= not((layer1_outputs(7195)) xor (layer1_outputs(3685)));
    layer2_outputs(9872) <= (layer1_outputs(10048)) and not (layer1_outputs(234));
    layer2_outputs(9873) <= layer1_outputs(2216);
    layer2_outputs(9874) <= (layer1_outputs(10217)) and (layer1_outputs(4839));
    layer2_outputs(9875) <= not(layer1_outputs(9115));
    layer2_outputs(9876) <= '1';
    layer2_outputs(9877) <= layer1_outputs(5410);
    layer2_outputs(9878) <= (layer1_outputs(6051)) and not (layer1_outputs(4025));
    layer2_outputs(9879) <= (layer1_outputs(2359)) and not (layer1_outputs(6492));
    layer2_outputs(9880) <= (layer1_outputs(4865)) and not (layer1_outputs(1848));
    layer2_outputs(9881) <= not((layer1_outputs(7613)) xor (layer1_outputs(3532)));
    layer2_outputs(9882) <= not(layer1_outputs(7449));
    layer2_outputs(9883) <= (layer1_outputs(10040)) or (layer1_outputs(9040));
    layer2_outputs(9884) <= '0';
    layer2_outputs(9885) <= layer1_outputs(2311);
    layer2_outputs(9886) <= '1';
    layer2_outputs(9887) <= not((layer1_outputs(9579)) or (layer1_outputs(992)));
    layer2_outputs(9888) <= not(layer1_outputs(2868));
    layer2_outputs(9889) <= layer1_outputs(1446);
    layer2_outputs(9890) <= layer1_outputs(8694);
    layer2_outputs(9891) <= layer1_outputs(1207);
    layer2_outputs(9892) <= layer1_outputs(4150);
    layer2_outputs(9893) <= (layer1_outputs(4095)) or (layer1_outputs(1490));
    layer2_outputs(9894) <= not(layer1_outputs(9551));
    layer2_outputs(9895) <= layer1_outputs(3400);
    layer2_outputs(9896) <= not(layer1_outputs(1557));
    layer2_outputs(9897) <= (layer1_outputs(5539)) and not (layer1_outputs(972));
    layer2_outputs(9898) <= not(layer1_outputs(455));
    layer2_outputs(9899) <= not(layer1_outputs(8841));
    layer2_outputs(9900) <= (layer1_outputs(1428)) or (layer1_outputs(9093));
    layer2_outputs(9901) <= not(layer1_outputs(8547)) or (layer1_outputs(4952));
    layer2_outputs(9902) <= (layer1_outputs(6847)) and (layer1_outputs(2603));
    layer2_outputs(9903) <= not(layer1_outputs(950));
    layer2_outputs(9904) <= not(layer1_outputs(3314));
    layer2_outputs(9905) <= layer1_outputs(8305);
    layer2_outputs(9906) <= not(layer1_outputs(10149));
    layer2_outputs(9907) <= not((layer1_outputs(9068)) and (layer1_outputs(9253)));
    layer2_outputs(9908) <= (layer1_outputs(3774)) and not (layer1_outputs(186));
    layer2_outputs(9909) <= not((layer1_outputs(8548)) xor (layer1_outputs(7412)));
    layer2_outputs(9910) <= layer1_outputs(7989);
    layer2_outputs(9911) <= (layer1_outputs(5411)) or (layer1_outputs(3911));
    layer2_outputs(9912) <= '1';
    layer2_outputs(9913) <= not(layer1_outputs(5587)) or (layer1_outputs(934));
    layer2_outputs(9914) <= not(layer1_outputs(4402)) or (layer1_outputs(9535));
    layer2_outputs(9915) <= layer1_outputs(6621);
    layer2_outputs(9916) <= not((layer1_outputs(7078)) and (layer1_outputs(8010)));
    layer2_outputs(9917) <= '0';
    layer2_outputs(9918) <= not(layer1_outputs(8968));
    layer2_outputs(9919) <= not(layer1_outputs(6098));
    layer2_outputs(9920) <= (layer1_outputs(5768)) and not (layer1_outputs(4349));
    layer2_outputs(9921) <= (layer1_outputs(919)) or (layer1_outputs(7604));
    layer2_outputs(9922) <= (layer1_outputs(1239)) or (layer1_outputs(75));
    layer2_outputs(9923) <= not(layer1_outputs(8046));
    layer2_outputs(9924) <= layer1_outputs(173);
    layer2_outputs(9925) <= not((layer1_outputs(1005)) xor (layer1_outputs(2887)));
    layer2_outputs(9926) <= not((layer1_outputs(4451)) or (layer1_outputs(4180)));
    layer2_outputs(9927) <= not(layer1_outputs(9394)) or (layer1_outputs(625));
    layer2_outputs(9928) <= layer1_outputs(1954);
    layer2_outputs(9929) <= not(layer1_outputs(6281));
    layer2_outputs(9930) <= not(layer1_outputs(9053));
    layer2_outputs(9931) <= not(layer1_outputs(10061)) or (layer1_outputs(9854));
    layer2_outputs(9932) <= layer1_outputs(7505);
    layer2_outputs(9933) <= not(layer1_outputs(3372));
    layer2_outputs(9934) <= layer1_outputs(7618);
    layer2_outputs(9935) <= (layer1_outputs(4025)) or (layer1_outputs(9828));
    layer2_outputs(9936) <= layer1_outputs(3231);
    layer2_outputs(9937) <= layer1_outputs(6731);
    layer2_outputs(9938) <= not((layer1_outputs(8206)) or (layer1_outputs(7855)));
    layer2_outputs(9939) <= not((layer1_outputs(2143)) or (layer1_outputs(3322)));
    layer2_outputs(9940) <= not(layer1_outputs(3110));
    layer2_outputs(9941) <= (layer1_outputs(6221)) and not (layer1_outputs(5933));
    layer2_outputs(9942) <= (layer1_outputs(8009)) xor (layer1_outputs(6081));
    layer2_outputs(9943) <= not(layer1_outputs(5700)) or (layer1_outputs(1326));
    layer2_outputs(9944) <= not(layer1_outputs(6944)) or (layer1_outputs(8535));
    layer2_outputs(9945) <= not(layer1_outputs(1398));
    layer2_outputs(9946) <= '1';
    layer2_outputs(9947) <= not(layer1_outputs(2118)) or (layer1_outputs(9816));
    layer2_outputs(9948) <= not((layer1_outputs(8701)) or (layer1_outputs(1410)));
    layer2_outputs(9949) <= not(layer1_outputs(113));
    layer2_outputs(9950) <= not(layer1_outputs(7081)) or (layer1_outputs(7882));
    layer2_outputs(9951) <= not(layer1_outputs(5597));
    layer2_outputs(9952) <= not(layer1_outputs(9023));
    layer2_outputs(9953) <= not(layer1_outputs(10001));
    layer2_outputs(9954) <= not((layer1_outputs(9084)) or (layer1_outputs(1335)));
    layer2_outputs(9955) <= layer1_outputs(8711);
    layer2_outputs(9956) <= (layer1_outputs(4029)) or (layer1_outputs(10168));
    layer2_outputs(9957) <= layer1_outputs(668);
    layer2_outputs(9958) <= layer1_outputs(7878);
    layer2_outputs(9959) <= not(layer1_outputs(2570));
    layer2_outputs(9960) <= '0';
    layer2_outputs(9961) <= '0';
    layer2_outputs(9962) <= layer1_outputs(9964);
    layer2_outputs(9963) <= '1';
    layer2_outputs(9964) <= not((layer1_outputs(353)) and (layer1_outputs(8683)));
    layer2_outputs(9965) <= not(layer1_outputs(6869));
    layer2_outputs(9966) <= not((layer1_outputs(7708)) or (layer1_outputs(288)));
    layer2_outputs(9967) <= not(layer1_outputs(6956));
    layer2_outputs(9968) <= not((layer1_outputs(2367)) or (layer1_outputs(5132)));
    layer2_outputs(9969) <= layer1_outputs(2396);
    layer2_outputs(9970) <= (layer1_outputs(6719)) and not (layer1_outputs(10164));
    layer2_outputs(9971) <= (layer1_outputs(2660)) and (layer1_outputs(10046));
    layer2_outputs(9972) <= not(layer1_outputs(6614)) or (layer1_outputs(9015));
    layer2_outputs(9973) <= layer1_outputs(2153);
    layer2_outputs(9974) <= layer1_outputs(2515);
    layer2_outputs(9975) <= not(layer1_outputs(1728)) or (layer1_outputs(3414));
    layer2_outputs(9976) <= not(layer1_outputs(6204));
    layer2_outputs(9977) <= not(layer1_outputs(8549));
    layer2_outputs(9978) <= (layer1_outputs(7005)) or (layer1_outputs(4176));
    layer2_outputs(9979) <= not(layer1_outputs(2940)) or (layer1_outputs(4967));
    layer2_outputs(9980) <= not((layer1_outputs(2054)) xor (layer1_outputs(8247)));
    layer2_outputs(9981) <= '1';
    layer2_outputs(9982) <= (layer1_outputs(2870)) or (layer1_outputs(706));
    layer2_outputs(9983) <= not((layer1_outputs(6531)) and (layer1_outputs(5021)));
    layer2_outputs(9984) <= (layer1_outputs(6806)) and (layer1_outputs(1547));
    layer2_outputs(9985) <= not(layer1_outputs(4580)) or (layer1_outputs(4750));
    layer2_outputs(9986) <= '0';
    layer2_outputs(9987) <= layer1_outputs(7686);
    layer2_outputs(9988) <= not((layer1_outputs(1508)) or (layer1_outputs(6220)));
    layer2_outputs(9989) <= not(layer1_outputs(3592));
    layer2_outputs(9990) <= not(layer1_outputs(8163));
    layer2_outputs(9991) <= layer1_outputs(7194);
    layer2_outputs(9992) <= not((layer1_outputs(5877)) xor (layer1_outputs(3898)));
    layer2_outputs(9993) <= not(layer1_outputs(5476));
    layer2_outputs(9994) <= not(layer1_outputs(9892));
    layer2_outputs(9995) <= (layer1_outputs(5782)) and (layer1_outputs(9095));
    layer2_outputs(9996) <= not(layer1_outputs(7268)) or (layer1_outputs(5050));
    layer2_outputs(9997) <= not(layer1_outputs(4926));
    layer2_outputs(9998) <= not(layer1_outputs(2705)) or (layer1_outputs(8377));
    layer2_outputs(9999) <= (layer1_outputs(8467)) xor (layer1_outputs(4552));
    layer2_outputs(10000) <= layer1_outputs(3170);
    layer2_outputs(10001) <= not(layer1_outputs(3726));
    layer2_outputs(10002) <= layer1_outputs(2925);
    layer2_outputs(10003) <= (layer1_outputs(2398)) or (layer1_outputs(9182));
    layer2_outputs(10004) <= layer1_outputs(9932);
    layer2_outputs(10005) <= '0';
    layer2_outputs(10006) <= (layer1_outputs(883)) and not (layer1_outputs(1763));
    layer2_outputs(10007) <= not(layer1_outputs(610)) or (layer1_outputs(6514));
    layer2_outputs(10008) <= not(layer1_outputs(6536)) or (layer1_outputs(4421));
    layer2_outputs(10009) <= not((layer1_outputs(5858)) and (layer1_outputs(9177)));
    layer2_outputs(10010) <= (layer1_outputs(1305)) xor (layer1_outputs(9283));
    layer2_outputs(10011) <= layer1_outputs(4899);
    layer2_outputs(10012) <= not((layer1_outputs(5117)) xor (layer1_outputs(300)));
    layer2_outputs(10013) <= (layer1_outputs(3972)) or (layer1_outputs(580));
    layer2_outputs(10014) <= (layer1_outputs(4151)) and not (layer1_outputs(6753));
    layer2_outputs(10015) <= not(layer1_outputs(7122)) or (layer1_outputs(9429));
    layer2_outputs(10016) <= not(layer1_outputs(1302));
    layer2_outputs(10017) <= not((layer1_outputs(7363)) or (layer1_outputs(8908)));
    layer2_outputs(10018) <= not(layer1_outputs(8854));
    layer2_outputs(10019) <= '0';
    layer2_outputs(10020) <= not(layer1_outputs(2638)) or (layer1_outputs(10044));
    layer2_outputs(10021) <= not(layer1_outputs(1375));
    layer2_outputs(10022) <= layer1_outputs(4537);
    layer2_outputs(10023) <= not(layer1_outputs(290));
    layer2_outputs(10024) <= not(layer1_outputs(6433)) or (layer1_outputs(6116));
    layer2_outputs(10025) <= layer1_outputs(8223);
    layer2_outputs(10026) <= (layer1_outputs(5453)) or (layer1_outputs(9344));
    layer2_outputs(10027) <= (layer1_outputs(8017)) and (layer1_outputs(1445));
    layer2_outputs(10028) <= not(layer1_outputs(1256)) or (layer1_outputs(4209));
    layer2_outputs(10029) <= (layer1_outputs(5017)) xor (layer1_outputs(5904));
    layer2_outputs(10030) <= not(layer1_outputs(665));
    layer2_outputs(10031) <= layer1_outputs(3817);
    layer2_outputs(10032) <= not(layer1_outputs(6718));
    layer2_outputs(10033) <= not(layer1_outputs(2324));
    layer2_outputs(10034) <= not(layer1_outputs(445));
    layer2_outputs(10035) <= layer1_outputs(7140);
    layer2_outputs(10036) <= (layer1_outputs(516)) xor (layer1_outputs(1303));
    layer2_outputs(10037) <= (layer1_outputs(6443)) or (layer1_outputs(6629));
    layer2_outputs(10038) <= not((layer1_outputs(4354)) and (layer1_outputs(6210)));
    layer2_outputs(10039) <= (layer1_outputs(9636)) and not (layer1_outputs(5575));
    layer2_outputs(10040) <= (layer1_outputs(1152)) xor (layer1_outputs(893));
    layer2_outputs(10041) <= (layer1_outputs(2233)) and not (layer1_outputs(3663));
    layer2_outputs(10042) <= not((layer1_outputs(4951)) xor (layer1_outputs(4116)));
    layer2_outputs(10043) <= (layer1_outputs(7592)) and not (layer1_outputs(5577));
    layer2_outputs(10044) <= (layer1_outputs(684)) xor (layer1_outputs(9783));
    layer2_outputs(10045) <= layer1_outputs(9655);
    layer2_outputs(10046) <= not((layer1_outputs(799)) and (layer1_outputs(4134)));
    layer2_outputs(10047) <= (layer1_outputs(1616)) and not (layer1_outputs(142));
    layer2_outputs(10048) <= (layer1_outputs(1038)) and not (layer1_outputs(10124));
    layer2_outputs(10049) <= not(layer1_outputs(3903));
    layer2_outputs(10050) <= layer1_outputs(6391);
    layer2_outputs(10051) <= (layer1_outputs(8647)) or (layer1_outputs(5397));
    layer2_outputs(10052) <= not(layer1_outputs(3035));
    layer2_outputs(10053) <= not((layer1_outputs(3102)) xor (layer1_outputs(4346)));
    layer2_outputs(10054) <= layer1_outputs(333);
    layer2_outputs(10055) <= not(layer1_outputs(8169));
    layer2_outputs(10056) <= '0';
    layer2_outputs(10057) <= not(layer1_outputs(8001));
    layer2_outputs(10058) <= not(layer1_outputs(2408)) or (layer1_outputs(6160));
    layer2_outputs(10059) <= not(layer1_outputs(9161));
    layer2_outputs(10060) <= '0';
    layer2_outputs(10061) <= not((layer1_outputs(1486)) xor (layer1_outputs(317)));
    layer2_outputs(10062) <= layer1_outputs(9831);
    layer2_outputs(10063) <= not(layer1_outputs(9303)) or (layer1_outputs(5591));
    layer2_outputs(10064) <= layer1_outputs(1808);
    layer2_outputs(10065) <= not(layer1_outputs(1967));
    layer2_outputs(10066) <= layer1_outputs(2096);
    layer2_outputs(10067) <= not((layer1_outputs(6589)) or (layer1_outputs(2153)));
    layer2_outputs(10068) <= not(layer1_outputs(3446));
    layer2_outputs(10069) <= layer1_outputs(7182);
    layer2_outputs(10070) <= not(layer1_outputs(2636));
    layer2_outputs(10071) <= '0';
    layer2_outputs(10072) <= not(layer1_outputs(2010)) or (layer1_outputs(6028));
    layer2_outputs(10073) <= not((layer1_outputs(6494)) and (layer1_outputs(4065)));
    layer2_outputs(10074) <= not((layer1_outputs(5729)) xor (layer1_outputs(2276)));
    layer2_outputs(10075) <= layer1_outputs(7920);
    layer2_outputs(10076) <= not(layer1_outputs(9183)) or (layer1_outputs(4670));
    layer2_outputs(10077) <= not(layer1_outputs(2154)) or (layer1_outputs(4794));
    layer2_outputs(10078) <= not((layer1_outputs(7430)) xor (layer1_outputs(9268)));
    layer2_outputs(10079) <= (layer1_outputs(8994)) and (layer1_outputs(1963));
    layer2_outputs(10080) <= layer1_outputs(9046);
    layer2_outputs(10081) <= layer1_outputs(6121);
    layer2_outputs(10082) <= not(layer1_outputs(269)) or (layer1_outputs(146));
    layer2_outputs(10083) <= not(layer1_outputs(4866));
    layer2_outputs(10084) <= (layer1_outputs(5631)) xor (layer1_outputs(4795));
    layer2_outputs(10085) <= layer1_outputs(2100);
    layer2_outputs(10086) <= not(layer1_outputs(1386));
    layer2_outputs(10087) <= '0';
    layer2_outputs(10088) <= (layer1_outputs(6329)) xor (layer1_outputs(2723));
    layer2_outputs(10089) <= (layer1_outputs(7723)) and not (layer1_outputs(2295));
    layer2_outputs(10090) <= (layer1_outputs(2759)) and not (layer1_outputs(7990));
    layer2_outputs(10091) <= (layer1_outputs(8268)) or (layer1_outputs(6364));
    layer2_outputs(10092) <= (layer1_outputs(6501)) and (layer1_outputs(4546));
    layer2_outputs(10093) <= '1';
    layer2_outputs(10094) <= (layer1_outputs(4056)) or (layer1_outputs(7655));
    layer2_outputs(10095) <= (layer1_outputs(6516)) xor (layer1_outputs(4205));
    layer2_outputs(10096) <= (layer1_outputs(3833)) and not (layer1_outputs(330));
    layer2_outputs(10097) <= (layer1_outputs(836)) and not (layer1_outputs(4694));
    layer2_outputs(10098) <= (layer1_outputs(10120)) and (layer1_outputs(7102));
    layer2_outputs(10099) <= not(layer1_outputs(2275)) or (layer1_outputs(7605));
    layer2_outputs(10100) <= (layer1_outputs(2328)) and (layer1_outputs(2475));
    layer2_outputs(10101) <= layer1_outputs(4860);
    layer2_outputs(10102) <= not(layer1_outputs(5990));
    layer2_outputs(10103) <= layer1_outputs(2265);
    layer2_outputs(10104) <= (layer1_outputs(9638)) and not (layer1_outputs(2297));
    layer2_outputs(10105) <= not(layer1_outputs(1795));
    layer2_outputs(10106) <= layer1_outputs(5026);
    layer2_outputs(10107) <= layer1_outputs(5698);
    layer2_outputs(10108) <= not(layer1_outputs(9683));
    layer2_outputs(10109) <= (layer1_outputs(2410)) or (layer1_outputs(5292));
    layer2_outputs(10110) <= (layer1_outputs(6395)) xor (layer1_outputs(3250));
    layer2_outputs(10111) <= not(layer1_outputs(3651));
    layer2_outputs(10112) <= not(layer1_outputs(9526)) or (layer1_outputs(1507));
    layer2_outputs(10113) <= (layer1_outputs(8096)) or (layer1_outputs(4959));
    layer2_outputs(10114) <= not(layer1_outputs(1841));
    layer2_outputs(10115) <= (layer1_outputs(8288)) and (layer1_outputs(4398));
    layer2_outputs(10116) <= layer1_outputs(704);
    layer2_outputs(10117) <= layer1_outputs(3856);
    layer2_outputs(10118) <= layer1_outputs(6657);
    layer2_outputs(10119) <= not((layer1_outputs(785)) xor (layer1_outputs(10111)));
    layer2_outputs(10120) <= not(layer1_outputs(10002));
    layer2_outputs(10121) <= (layer1_outputs(4504)) xor (layer1_outputs(3196));
    layer2_outputs(10122) <= (layer1_outputs(746)) or (layer1_outputs(3623));
    layer2_outputs(10123) <= not(layer1_outputs(6020)) or (layer1_outputs(6325));
    layer2_outputs(10124) <= not((layer1_outputs(9637)) xor (layer1_outputs(4743)));
    layer2_outputs(10125) <= layer1_outputs(3093);
    layer2_outputs(10126) <= not(layer1_outputs(4401));
    layer2_outputs(10127) <= (layer1_outputs(6012)) or (layer1_outputs(2170));
    layer2_outputs(10128) <= not(layer1_outputs(9657));
    layer2_outputs(10129) <= not(layer1_outputs(9650)) or (layer1_outputs(2983));
    layer2_outputs(10130) <= (layer1_outputs(7847)) and (layer1_outputs(1345));
    layer2_outputs(10131) <= (layer1_outputs(2804)) xor (layer1_outputs(3626));
    layer2_outputs(10132) <= layer1_outputs(2024);
    layer2_outputs(10133) <= not((layer1_outputs(6959)) and (layer1_outputs(2854)));
    layer2_outputs(10134) <= not((layer1_outputs(2747)) and (layer1_outputs(1014)));
    layer2_outputs(10135) <= not((layer1_outputs(3053)) and (layer1_outputs(2875)));
    layer2_outputs(10136) <= not((layer1_outputs(740)) and (layer1_outputs(4296)));
    layer2_outputs(10137) <= '0';
    layer2_outputs(10138) <= layer1_outputs(2966);
    layer2_outputs(10139) <= (layer1_outputs(9691)) or (layer1_outputs(8431));
    layer2_outputs(10140) <= not(layer1_outputs(1383)) or (layer1_outputs(6122));
    layer2_outputs(10141) <= layer1_outputs(4754);
    layer2_outputs(10142) <= not(layer1_outputs(6103));
    layer2_outputs(10143) <= (layer1_outputs(5628)) and not (layer1_outputs(8556));
    layer2_outputs(10144) <= not((layer1_outputs(5691)) and (layer1_outputs(3873)));
    layer2_outputs(10145) <= layer1_outputs(4451);
    layer2_outputs(10146) <= not(layer1_outputs(4121));
    layer2_outputs(10147) <= layer1_outputs(8569);
    layer2_outputs(10148) <= '1';
    layer2_outputs(10149) <= not((layer1_outputs(10005)) and (layer1_outputs(378)));
    layer2_outputs(10150) <= '1';
    layer2_outputs(10151) <= '1';
    layer2_outputs(10152) <= not(layer1_outputs(3878)) or (layer1_outputs(5012));
    layer2_outputs(10153) <= not((layer1_outputs(7979)) xor (layer1_outputs(8931)));
    layer2_outputs(10154) <= not((layer1_outputs(10123)) or (layer1_outputs(7531)));
    layer2_outputs(10155) <= layer1_outputs(10138);
    layer2_outputs(10156) <= layer1_outputs(3557);
    layer2_outputs(10157) <= not(layer1_outputs(1274));
    layer2_outputs(10158) <= layer1_outputs(5701);
    layer2_outputs(10159) <= not(layer1_outputs(2760));
    layer2_outputs(10160) <= (layer1_outputs(497)) and not (layer1_outputs(4654));
    layer2_outputs(10161) <= not(layer1_outputs(5640));
    layer2_outputs(10162) <= layer1_outputs(707);
    layer2_outputs(10163) <= (layer1_outputs(3318)) xor (layer1_outputs(3647));
    layer2_outputs(10164) <= layer1_outputs(562);
    layer2_outputs(10165) <= (layer1_outputs(258)) and (layer1_outputs(3210));
    layer2_outputs(10166) <= (layer1_outputs(6260)) and not (layer1_outputs(9523));
    layer2_outputs(10167) <= not(layer1_outputs(2399));
    layer2_outputs(10168) <= layer1_outputs(6151);
    layer2_outputs(10169) <= not(layer1_outputs(8195));
    layer2_outputs(10170) <= not(layer1_outputs(9025)) or (layer1_outputs(2674));
    layer2_outputs(10171) <= not(layer1_outputs(8683));
    layer2_outputs(10172) <= layer1_outputs(4371);
    layer2_outputs(10173) <= not(layer1_outputs(1789));
    layer2_outputs(10174) <= layer1_outputs(3768);
    layer2_outputs(10175) <= (layer1_outputs(10117)) xor (layer1_outputs(6088));
    layer2_outputs(10176) <= not(layer1_outputs(834));
    layer2_outputs(10177) <= not(layer1_outputs(6998)) or (layer1_outputs(2034));
    layer2_outputs(10178) <= not((layer1_outputs(5817)) or (layer1_outputs(1894)));
    layer2_outputs(10179) <= not(layer1_outputs(6178));
    layer2_outputs(10180) <= not(layer1_outputs(12)) or (layer1_outputs(7926));
    layer2_outputs(10181) <= (layer1_outputs(5319)) and (layer1_outputs(4949));
    layer2_outputs(10182) <= not((layer1_outputs(6847)) xor (layer1_outputs(3232)));
    layer2_outputs(10183) <= not(layer1_outputs(8151));
    layer2_outputs(10184) <= not((layer1_outputs(7315)) xor (layer1_outputs(7717)));
    layer2_outputs(10185) <= layer1_outputs(6877);
    layer2_outputs(10186) <= not(layer1_outputs(8319));
    layer2_outputs(10187) <= not((layer1_outputs(8092)) and (layer1_outputs(7901)));
    layer2_outputs(10188) <= layer1_outputs(3254);
    layer2_outputs(10189) <= not((layer1_outputs(9212)) or (layer1_outputs(3545)));
    layer2_outputs(10190) <= not(layer1_outputs(3651));
    layer2_outputs(10191) <= layer1_outputs(7935);
    layer2_outputs(10192) <= not(layer1_outputs(6355));
    layer2_outputs(10193) <= not((layer1_outputs(9479)) or (layer1_outputs(5426)));
    layer2_outputs(10194) <= (layer1_outputs(1157)) xor (layer1_outputs(448));
    layer2_outputs(10195) <= not((layer1_outputs(8380)) or (layer1_outputs(3088)));
    layer2_outputs(10196) <= not((layer1_outputs(3398)) or (layer1_outputs(4648)));
    layer2_outputs(10197) <= not((layer1_outputs(6254)) or (layer1_outputs(5423)));
    layer2_outputs(10198) <= (layer1_outputs(9658)) and (layer1_outputs(334));
    layer2_outputs(10199) <= layer1_outputs(6485);
    layer2_outputs(10200) <= '0';
    layer2_outputs(10201) <= (layer1_outputs(5168)) and not (layer1_outputs(1889));
    layer2_outputs(10202) <= not((layer1_outputs(1909)) and (layer1_outputs(743)));
    layer2_outputs(10203) <= not((layer1_outputs(8306)) and (layer1_outputs(7612)));
    layer2_outputs(10204) <= not(layer1_outputs(2372)) or (layer1_outputs(2534));
    layer2_outputs(10205) <= (layer1_outputs(8500)) or (layer1_outputs(8498));
    layer2_outputs(10206) <= layer1_outputs(9908);
    layer2_outputs(10207) <= layer1_outputs(2817);
    layer2_outputs(10208) <= layer1_outputs(6482);
    layer2_outputs(10209) <= (layer1_outputs(570)) xor (layer1_outputs(6379));
    layer2_outputs(10210) <= layer1_outputs(4627);
    layer2_outputs(10211) <= not(layer1_outputs(3875));
    layer2_outputs(10212) <= (layer1_outputs(3830)) or (layer1_outputs(8820));
    layer2_outputs(10213) <= (layer1_outputs(4227)) and not (layer1_outputs(2559));
    layer2_outputs(10214) <= (layer1_outputs(3182)) or (layer1_outputs(5552));
    layer2_outputs(10215) <= layer1_outputs(2391);
    layer2_outputs(10216) <= layer1_outputs(9287);
    layer2_outputs(10217) <= not(layer1_outputs(4776)) or (layer1_outputs(9619));
    layer2_outputs(10218) <= layer1_outputs(6700);
    layer2_outputs(10219) <= (layer1_outputs(9584)) and not (layer1_outputs(7046));
    layer2_outputs(10220) <= layer1_outputs(9531);
    layer2_outputs(10221) <= (layer1_outputs(7684)) and (layer1_outputs(8732));
    layer2_outputs(10222) <= not(layer1_outputs(10075));
    layer2_outputs(10223) <= '0';
    layer2_outputs(10224) <= '0';
    layer2_outputs(10225) <= not(layer1_outputs(9909)) or (layer1_outputs(8228));
    layer2_outputs(10226) <= (layer1_outputs(5001)) or (layer1_outputs(3222));
    layer2_outputs(10227) <= not((layer1_outputs(2758)) and (layer1_outputs(1883)));
    layer2_outputs(10228) <= not((layer1_outputs(1247)) or (layer1_outputs(4944)));
    layer2_outputs(10229) <= '0';
    layer2_outputs(10230) <= (layer1_outputs(4363)) and not (layer1_outputs(3552));
    layer2_outputs(10231) <= (layer1_outputs(9681)) and (layer1_outputs(7171));
    layer2_outputs(10232) <= not(layer1_outputs(3700)) or (layer1_outputs(927));
    layer2_outputs(10233) <= '1';
    layer2_outputs(10234) <= layer1_outputs(4982);
    layer2_outputs(10235) <= not(layer1_outputs(1403));
    layer2_outputs(10236) <= layer1_outputs(4921);
    layer2_outputs(10237) <= layer1_outputs(3122);
    layer2_outputs(10238) <= not(layer1_outputs(1435));
    layer2_outputs(10239) <= not(layer1_outputs(6366));
    layer3_outputs(0) <= (layer2_outputs(2299)) or (layer2_outputs(6364));
    layer3_outputs(1) <= not(layer2_outputs(8130)) or (layer2_outputs(1316));
    layer3_outputs(2) <= not(layer2_outputs(7847));
    layer3_outputs(3) <= not(layer2_outputs(5006)) or (layer2_outputs(4020));
    layer3_outputs(4) <= layer2_outputs(529);
    layer3_outputs(5) <= not(layer2_outputs(5327));
    layer3_outputs(6) <= not(layer2_outputs(7461)) or (layer2_outputs(2136));
    layer3_outputs(7) <= not(layer2_outputs(5747));
    layer3_outputs(8) <= not(layer2_outputs(2212)) or (layer2_outputs(9863));
    layer3_outputs(9) <= layer2_outputs(7090);
    layer3_outputs(10) <= not((layer2_outputs(4771)) xor (layer2_outputs(3392)));
    layer3_outputs(11) <= '0';
    layer3_outputs(12) <= not(layer2_outputs(2614));
    layer3_outputs(13) <= not(layer2_outputs(5742));
    layer3_outputs(14) <= layer2_outputs(1766);
    layer3_outputs(15) <= not(layer2_outputs(5346)) or (layer2_outputs(5242));
    layer3_outputs(16) <= not(layer2_outputs(8255));
    layer3_outputs(17) <= not(layer2_outputs(1354)) or (layer2_outputs(8369));
    layer3_outputs(18) <= not(layer2_outputs(3979));
    layer3_outputs(19) <= layer2_outputs(10050);
    layer3_outputs(20) <= '1';
    layer3_outputs(21) <= layer2_outputs(9843);
    layer3_outputs(22) <= not((layer2_outputs(3512)) or (layer2_outputs(6744)));
    layer3_outputs(23) <= not(layer2_outputs(6778));
    layer3_outputs(24) <= (layer2_outputs(476)) and (layer2_outputs(6467));
    layer3_outputs(25) <= not(layer2_outputs(5487));
    layer3_outputs(26) <= '1';
    layer3_outputs(27) <= not(layer2_outputs(5025));
    layer3_outputs(28) <= (layer2_outputs(5177)) or (layer2_outputs(4740));
    layer3_outputs(29) <= (layer2_outputs(2717)) xor (layer2_outputs(6408));
    layer3_outputs(30) <= not(layer2_outputs(3569));
    layer3_outputs(31) <= (layer2_outputs(3477)) and not (layer2_outputs(301));
    layer3_outputs(32) <= layer2_outputs(5838);
    layer3_outputs(33) <= (layer2_outputs(10170)) or (layer2_outputs(7889));
    layer3_outputs(34) <= not(layer2_outputs(6681)) or (layer2_outputs(960));
    layer3_outputs(35) <= not(layer2_outputs(8308)) or (layer2_outputs(7572));
    layer3_outputs(36) <= not(layer2_outputs(3346));
    layer3_outputs(37) <= not(layer2_outputs(5102)) or (layer2_outputs(215));
    layer3_outputs(38) <= layer2_outputs(9389);
    layer3_outputs(39) <= not((layer2_outputs(946)) and (layer2_outputs(2417)));
    layer3_outputs(40) <= not((layer2_outputs(2012)) xor (layer2_outputs(3319)));
    layer3_outputs(41) <= layer2_outputs(7044);
    layer3_outputs(42) <= not(layer2_outputs(127));
    layer3_outputs(43) <= (layer2_outputs(8385)) and not (layer2_outputs(9779));
    layer3_outputs(44) <= not(layer2_outputs(10207));
    layer3_outputs(45) <= not(layer2_outputs(8381)) or (layer2_outputs(7812));
    layer3_outputs(46) <= not(layer2_outputs(7536)) or (layer2_outputs(5032));
    layer3_outputs(47) <= layer2_outputs(1972);
    layer3_outputs(48) <= (layer2_outputs(4863)) and not (layer2_outputs(4767));
    layer3_outputs(49) <= (layer2_outputs(1965)) and (layer2_outputs(9240));
    layer3_outputs(50) <= (layer2_outputs(4166)) or (layer2_outputs(877));
    layer3_outputs(51) <= not(layer2_outputs(4312));
    layer3_outputs(52) <= layer2_outputs(1229);
    layer3_outputs(53) <= layer2_outputs(1390);
    layer3_outputs(54) <= not(layer2_outputs(754)) or (layer2_outputs(2380));
    layer3_outputs(55) <= layer2_outputs(5424);
    layer3_outputs(56) <= not(layer2_outputs(5593));
    layer3_outputs(57) <= not(layer2_outputs(4156));
    layer3_outputs(58) <= not(layer2_outputs(5993));
    layer3_outputs(59) <= layer2_outputs(8925);
    layer3_outputs(60) <= not((layer2_outputs(443)) xor (layer2_outputs(6436)));
    layer3_outputs(61) <= not(layer2_outputs(6743));
    layer3_outputs(62) <= not(layer2_outputs(3973));
    layer3_outputs(63) <= not(layer2_outputs(1407));
    layer3_outputs(64) <= not(layer2_outputs(2268));
    layer3_outputs(65) <= not(layer2_outputs(4170));
    layer3_outputs(66) <= layer2_outputs(937);
    layer3_outputs(67) <= not(layer2_outputs(4541));
    layer3_outputs(68) <= layer2_outputs(9246);
    layer3_outputs(69) <= not(layer2_outputs(3573));
    layer3_outputs(70) <= (layer2_outputs(1193)) or (layer2_outputs(8971));
    layer3_outputs(71) <= layer2_outputs(97);
    layer3_outputs(72) <= (layer2_outputs(7443)) or (layer2_outputs(2206));
    layer3_outputs(73) <= not((layer2_outputs(2112)) xor (layer2_outputs(8641)));
    layer3_outputs(74) <= layer2_outputs(3890);
    layer3_outputs(75) <= not(layer2_outputs(2368));
    layer3_outputs(76) <= not(layer2_outputs(5326)) or (layer2_outputs(4272));
    layer3_outputs(77) <= not(layer2_outputs(1615)) or (layer2_outputs(5483));
    layer3_outputs(78) <= '1';
    layer3_outputs(79) <= not(layer2_outputs(6763)) or (layer2_outputs(4404));
    layer3_outputs(80) <= not((layer2_outputs(8830)) or (layer2_outputs(1956)));
    layer3_outputs(81) <= not(layer2_outputs(8636)) or (layer2_outputs(7021));
    layer3_outputs(82) <= layer2_outputs(1168);
    layer3_outputs(83) <= not(layer2_outputs(3311)) or (layer2_outputs(3722));
    layer3_outputs(84) <= not(layer2_outputs(6836)) or (layer2_outputs(9981));
    layer3_outputs(85) <= not(layer2_outputs(6208));
    layer3_outputs(86) <= not(layer2_outputs(2015));
    layer3_outputs(87) <= (layer2_outputs(6238)) and not (layer2_outputs(9884));
    layer3_outputs(88) <= layer2_outputs(2972);
    layer3_outputs(89) <= not(layer2_outputs(9948));
    layer3_outputs(90) <= layer2_outputs(1138);
    layer3_outputs(91) <= not(layer2_outputs(5300));
    layer3_outputs(92) <= layer2_outputs(2197);
    layer3_outputs(93) <= not((layer2_outputs(4176)) xor (layer2_outputs(2762)));
    layer3_outputs(94) <= layer2_outputs(9110);
    layer3_outputs(95) <= not(layer2_outputs(4195));
    layer3_outputs(96) <= not(layer2_outputs(8727)) or (layer2_outputs(1051));
    layer3_outputs(97) <= not(layer2_outputs(1752)) or (layer2_outputs(7869));
    layer3_outputs(98) <= (layer2_outputs(7153)) xor (layer2_outputs(3585));
    layer3_outputs(99) <= '1';
    layer3_outputs(100) <= not(layer2_outputs(3246));
    layer3_outputs(101) <= (layer2_outputs(1921)) and not (layer2_outputs(4723));
    layer3_outputs(102) <= not(layer2_outputs(5415)) or (layer2_outputs(6604));
    layer3_outputs(103) <= not(layer2_outputs(8286));
    layer3_outputs(104) <= not((layer2_outputs(7565)) xor (layer2_outputs(2013)));
    layer3_outputs(105) <= layer2_outputs(1314);
    layer3_outputs(106) <= not((layer2_outputs(7620)) xor (layer2_outputs(1645)));
    layer3_outputs(107) <= not(layer2_outputs(1678)) or (layer2_outputs(598));
    layer3_outputs(108) <= not(layer2_outputs(7783)) or (layer2_outputs(5728));
    layer3_outputs(109) <= not(layer2_outputs(5158));
    layer3_outputs(110) <= (layer2_outputs(8934)) or (layer2_outputs(735));
    layer3_outputs(111) <= layer2_outputs(5911);
    layer3_outputs(112) <= not(layer2_outputs(6034));
    layer3_outputs(113) <= not(layer2_outputs(1722));
    layer3_outputs(114) <= not(layer2_outputs(6343));
    layer3_outputs(115) <= not(layer2_outputs(5867)) or (layer2_outputs(7249));
    layer3_outputs(116) <= (layer2_outputs(10072)) xor (layer2_outputs(1635));
    layer3_outputs(117) <= not((layer2_outputs(6787)) xor (layer2_outputs(5590)));
    layer3_outputs(118) <= not(layer2_outputs(8230));
    layer3_outputs(119) <= (layer2_outputs(5696)) and not (layer2_outputs(7606));
    layer3_outputs(120) <= not(layer2_outputs(10232));
    layer3_outputs(121) <= not((layer2_outputs(8629)) and (layer2_outputs(9694)));
    layer3_outputs(122) <= not(layer2_outputs(3082)) or (layer2_outputs(7346));
    layer3_outputs(123) <= layer2_outputs(6948);
    layer3_outputs(124) <= (layer2_outputs(265)) and not (layer2_outputs(7028));
    layer3_outputs(125) <= '1';
    layer3_outputs(126) <= (layer2_outputs(1976)) xor (layer2_outputs(9163));
    layer3_outputs(127) <= (layer2_outputs(6305)) or (layer2_outputs(4342));
    layer3_outputs(128) <= (layer2_outputs(10104)) or (layer2_outputs(4087));
    layer3_outputs(129) <= not(layer2_outputs(1598));
    layer3_outputs(130) <= (layer2_outputs(7983)) xor (layer2_outputs(7272));
    layer3_outputs(131) <= not((layer2_outputs(8074)) xor (layer2_outputs(1737)));
    layer3_outputs(132) <= layer2_outputs(4269);
    layer3_outputs(133) <= not(layer2_outputs(2871));
    layer3_outputs(134) <= layer2_outputs(9930);
    layer3_outputs(135) <= layer2_outputs(10096);
    layer3_outputs(136) <= not(layer2_outputs(6402));
    layer3_outputs(137) <= layer2_outputs(3452);
    layer3_outputs(138) <= (layer2_outputs(1433)) xor (layer2_outputs(1652));
    layer3_outputs(139) <= (layer2_outputs(2310)) and (layer2_outputs(9433));
    layer3_outputs(140) <= not(layer2_outputs(3080));
    layer3_outputs(141) <= not(layer2_outputs(8527));
    layer3_outputs(142) <= (layer2_outputs(9695)) xor (layer2_outputs(285));
    layer3_outputs(143) <= (layer2_outputs(837)) and not (layer2_outputs(1346));
    layer3_outputs(144) <= layer2_outputs(931);
    layer3_outputs(145) <= layer2_outputs(7275);
    layer3_outputs(146) <= not((layer2_outputs(183)) or (layer2_outputs(8331)));
    layer3_outputs(147) <= layer2_outputs(7067);
    layer3_outputs(148) <= not(layer2_outputs(3487));
    layer3_outputs(149) <= not(layer2_outputs(8651));
    layer3_outputs(150) <= not((layer2_outputs(4212)) or (layer2_outputs(2827)));
    layer3_outputs(151) <= (layer2_outputs(6382)) and (layer2_outputs(1685));
    layer3_outputs(152) <= layer2_outputs(9128);
    layer3_outputs(153) <= layer2_outputs(409);
    layer3_outputs(154) <= not(layer2_outputs(3243));
    layer3_outputs(155) <= '1';
    layer3_outputs(156) <= layer2_outputs(10176);
    layer3_outputs(157) <= not(layer2_outputs(8327));
    layer3_outputs(158) <= not((layer2_outputs(6876)) and (layer2_outputs(6254)));
    layer3_outputs(159) <= '1';
    layer3_outputs(160) <= (layer2_outputs(611)) and not (layer2_outputs(2354));
    layer3_outputs(161) <= layer2_outputs(6628);
    layer3_outputs(162) <= layer2_outputs(9776);
    layer3_outputs(163) <= not(layer2_outputs(3037));
    layer3_outputs(164) <= not(layer2_outputs(7217));
    layer3_outputs(165) <= not(layer2_outputs(1075));
    layer3_outputs(166) <= layer2_outputs(3832);
    layer3_outputs(167) <= layer2_outputs(762);
    layer3_outputs(168) <= layer2_outputs(5329);
    layer3_outputs(169) <= not((layer2_outputs(9767)) xor (layer2_outputs(8289)));
    layer3_outputs(170) <= layer2_outputs(7515);
    layer3_outputs(171) <= (layer2_outputs(5361)) and not (layer2_outputs(2660));
    layer3_outputs(172) <= layer2_outputs(4794);
    layer3_outputs(173) <= not(layer2_outputs(558));
    layer3_outputs(174) <= not((layer2_outputs(6161)) or (layer2_outputs(918)));
    layer3_outputs(175) <= (layer2_outputs(5460)) and not (layer2_outputs(5075));
    layer3_outputs(176) <= (layer2_outputs(2537)) xor (layer2_outputs(1259));
    layer3_outputs(177) <= layer2_outputs(3655);
    layer3_outputs(178) <= layer2_outputs(7989);
    layer3_outputs(179) <= layer2_outputs(4247);
    layer3_outputs(180) <= '1';
    layer3_outputs(181) <= layer2_outputs(10220);
    layer3_outputs(182) <= not(layer2_outputs(7866));
    layer3_outputs(183) <= not((layer2_outputs(6777)) xor (layer2_outputs(4457)));
    layer3_outputs(184) <= (layer2_outputs(4019)) xor (layer2_outputs(10017));
    layer3_outputs(185) <= (layer2_outputs(8522)) or (layer2_outputs(3445));
    layer3_outputs(186) <= (layer2_outputs(5091)) and not (layer2_outputs(6643));
    layer3_outputs(187) <= not(layer2_outputs(9089)) or (layer2_outputs(5191));
    layer3_outputs(188) <= (layer2_outputs(8283)) and not (layer2_outputs(2731));
    layer3_outputs(189) <= layer2_outputs(10074);
    layer3_outputs(190) <= (layer2_outputs(1715)) and (layer2_outputs(9795));
    layer3_outputs(191) <= layer2_outputs(8022);
    layer3_outputs(192) <= not(layer2_outputs(6006));
    layer3_outputs(193) <= layer2_outputs(9378);
    layer3_outputs(194) <= not((layer2_outputs(4182)) xor (layer2_outputs(2085)));
    layer3_outputs(195) <= not(layer2_outputs(3755)) or (layer2_outputs(5634));
    layer3_outputs(196) <= layer2_outputs(1730);
    layer3_outputs(197) <= layer2_outputs(8376);
    layer3_outputs(198) <= not(layer2_outputs(6470));
    layer3_outputs(199) <= (layer2_outputs(5824)) and not (layer2_outputs(3557));
    layer3_outputs(200) <= not(layer2_outputs(9361)) or (layer2_outputs(7089));
    layer3_outputs(201) <= not(layer2_outputs(3118)) or (layer2_outputs(9674));
    layer3_outputs(202) <= (layer2_outputs(4264)) and (layer2_outputs(7155));
    layer3_outputs(203) <= not(layer2_outputs(8764));
    layer3_outputs(204) <= layer2_outputs(3668);
    layer3_outputs(205) <= layer2_outputs(7589);
    layer3_outputs(206) <= not(layer2_outputs(6495)) or (layer2_outputs(10070));
    layer3_outputs(207) <= layer2_outputs(10014);
    layer3_outputs(208) <= layer2_outputs(110);
    layer3_outputs(209) <= (layer2_outputs(7669)) and not (layer2_outputs(2802));
    layer3_outputs(210) <= not((layer2_outputs(435)) or (layer2_outputs(7787)));
    layer3_outputs(211) <= not((layer2_outputs(10188)) and (layer2_outputs(3019)));
    layer3_outputs(212) <= layer2_outputs(8289);
    layer3_outputs(213) <= not(layer2_outputs(2678)) or (layer2_outputs(4325));
    layer3_outputs(214) <= not((layer2_outputs(4149)) xor (layer2_outputs(8057)));
    layer3_outputs(215) <= not(layer2_outputs(5431));
    layer3_outputs(216) <= (layer2_outputs(765)) and not (layer2_outputs(4993));
    layer3_outputs(217) <= '0';
    layer3_outputs(218) <= layer2_outputs(2932);
    layer3_outputs(219) <= (layer2_outputs(9004)) and (layer2_outputs(9911));
    layer3_outputs(220) <= layer2_outputs(5403);
    layer3_outputs(221) <= (layer2_outputs(2420)) and (layer2_outputs(1378));
    layer3_outputs(222) <= not(layer2_outputs(121));
    layer3_outputs(223) <= not((layer2_outputs(2947)) xor (layer2_outputs(8662)));
    layer3_outputs(224) <= not(layer2_outputs(9712));
    layer3_outputs(225) <= (layer2_outputs(5853)) or (layer2_outputs(9065));
    layer3_outputs(226) <= not(layer2_outputs(7077));
    layer3_outputs(227) <= not(layer2_outputs(4572));
    layer3_outputs(228) <= not(layer2_outputs(6254)) or (layer2_outputs(157));
    layer3_outputs(229) <= not(layer2_outputs(2203)) or (layer2_outputs(5814));
    layer3_outputs(230) <= '0';
    layer3_outputs(231) <= (layer2_outputs(1081)) and not (layer2_outputs(9711));
    layer3_outputs(232) <= not(layer2_outputs(7156));
    layer3_outputs(233) <= '0';
    layer3_outputs(234) <= layer2_outputs(8043);
    layer3_outputs(235) <= not(layer2_outputs(9149));
    layer3_outputs(236) <= not(layer2_outputs(7073)) or (layer2_outputs(5562));
    layer3_outputs(237) <= not((layer2_outputs(1325)) or (layer2_outputs(229)));
    layer3_outputs(238) <= not(layer2_outputs(1440));
    layer3_outputs(239) <= '1';
    layer3_outputs(240) <= (layer2_outputs(4054)) and (layer2_outputs(6319));
    layer3_outputs(241) <= layer2_outputs(9311);
    layer3_outputs(242) <= (layer2_outputs(7784)) and (layer2_outputs(1403));
    layer3_outputs(243) <= layer2_outputs(3658);
    layer3_outputs(244) <= (layer2_outputs(6848)) or (layer2_outputs(2210));
    layer3_outputs(245) <= (layer2_outputs(7457)) or (layer2_outputs(584));
    layer3_outputs(246) <= not(layer2_outputs(4642));
    layer3_outputs(247) <= not((layer2_outputs(2758)) xor (layer2_outputs(7564)));
    layer3_outputs(248) <= not((layer2_outputs(4312)) xor (layer2_outputs(6532)));
    layer3_outputs(249) <= layer2_outputs(6904);
    layer3_outputs(250) <= not(layer2_outputs(2844));
    layer3_outputs(251) <= not(layer2_outputs(3358));
    layer3_outputs(252) <= layer2_outputs(4200);
    layer3_outputs(253) <= '0';
    layer3_outputs(254) <= layer2_outputs(7036);
    layer3_outputs(255) <= (layer2_outputs(4917)) and not (layer2_outputs(4038));
    layer3_outputs(256) <= layer2_outputs(9832);
    layer3_outputs(257) <= not(layer2_outputs(7775));
    layer3_outputs(258) <= layer2_outputs(933);
    layer3_outputs(259) <= layer2_outputs(4439);
    layer3_outputs(260) <= not(layer2_outputs(110));
    layer3_outputs(261) <= not(layer2_outputs(3612));
    layer3_outputs(262) <= not((layer2_outputs(472)) or (layer2_outputs(1108)));
    layer3_outputs(263) <= not(layer2_outputs(10220));
    layer3_outputs(264) <= not(layer2_outputs(5506));
    layer3_outputs(265) <= (layer2_outputs(8906)) or (layer2_outputs(10178));
    layer3_outputs(266) <= layer2_outputs(3920);
    layer3_outputs(267) <= (layer2_outputs(6960)) xor (layer2_outputs(3363));
    layer3_outputs(268) <= layer2_outputs(1245);
    layer3_outputs(269) <= not(layer2_outputs(575)) or (layer2_outputs(3739));
    layer3_outputs(270) <= not(layer2_outputs(1456));
    layer3_outputs(271) <= (layer2_outputs(9713)) xor (layer2_outputs(2704));
    layer3_outputs(272) <= layer2_outputs(4132);
    layer3_outputs(273) <= not(layer2_outputs(4803)) or (layer2_outputs(8975));
    layer3_outputs(274) <= not(layer2_outputs(9084)) or (layer2_outputs(6306));
    layer3_outputs(275) <= not((layer2_outputs(2739)) or (layer2_outputs(2676)));
    layer3_outputs(276) <= layer2_outputs(3056);
    layer3_outputs(277) <= layer2_outputs(5338);
    layer3_outputs(278) <= layer2_outputs(1379);
    layer3_outputs(279) <= (layer2_outputs(7194)) or (layer2_outputs(9696));
    layer3_outputs(280) <= not((layer2_outputs(2939)) and (layer2_outputs(8246)));
    layer3_outputs(281) <= '1';
    layer3_outputs(282) <= (layer2_outputs(5342)) xor (layer2_outputs(1264));
    layer3_outputs(283) <= (layer2_outputs(7188)) and not (layer2_outputs(8612));
    layer3_outputs(284) <= not((layer2_outputs(7049)) xor (layer2_outputs(5381)));
    layer3_outputs(285) <= not(layer2_outputs(1835)) or (layer2_outputs(5976));
    layer3_outputs(286) <= not(layer2_outputs(5771));
    layer3_outputs(287) <= not((layer2_outputs(3656)) and (layer2_outputs(3727)));
    layer3_outputs(288) <= (layer2_outputs(2807)) and not (layer2_outputs(8082));
    layer3_outputs(289) <= not(layer2_outputs(4315));
    layer3_outputs(290) <= layer2_outputs(7494);
    layer3_outputs(291) <= (layer2_outputs(9424)) and not (layer2_outputs(6287));
    layer3_outputs(292) <= not(layer2_outputs(7105));
    layer3_outputs(293) <= layer2_outputs(2252);
    layer3_outputs(294) <= not(layer2_outputs(9528));
    layer3_outputs(295) <= layer2_outputs(1906);
    layer3_outputs(296) <= not(layer2_outputs(5721));
    layer3_outputs(297) <= not(layer2_outputs(9536));
    layer3_outputs(298) <= (layer2_outputs(9459)) xor (layer2_outputs(830));
    layer3_outputs(299) <= not(layer2_outputs(7007)) or (layer2_outputs(2949));
    layer3_outputs(300) <= (layer2_outputs(4500)) and (layer2_outputs(1924));
    layer3_outputs(301) <= not(layer2_outputs(5676));
    layer3_outputs(302) <= not(layer2_outputs(10143));
    layer3_outputs(303) <= not((layer2_outputs(9923)) xor (layer2_outputs(5306)));
    layer3_outputs(304) <= not((layer2_outputs(1753)) or (layer2_outputs(4164)));
    layer3_outputs(305) <= layer2_outputs(2691);
    layer3_outputs(306) <= layer2_outputs(2544);
    layer3_outputs(307) <= not((layer2_outputs(9412)) or (layer2_outputs(9071)));
    layer3_outputs(308) <= layer2_outputs(5366);
    layer3_outputs(309) <= (layer2_outputs(88)) and not (layer2_outputs(199));
    layer3_outputs(310) <= not((layer2_outputs(3770)) or (layer2_outputs(389)));
    layer3_outputs(311) <= not(layer2_outputs(2345));
    layer3_outputs(312) <= layer2_outputs(622);
    layer3_outputs(313) <= not((layer2_outputs(629)) or (layer2_outputs(5972)));
    layer3_outputs(314) <= not(layer2_outputs(8976));
    layer3_outputs(315) <= layer2_outputs(5574);
    layer3_outputs(316) <= (layer2_outputs(364)) and not (layer2_outputs(1208));
    layer3_outputs(317) <= (layer2_outputs(3800)) xor (layer2_outputs(5567));
    layer3_outputs(318) <= layer2_outputs(8092);
    layer3_outputs(319) <= (layer2_outputs(4446)) and not (layer2_outputs(8890));
    layer3_outputs(320) <= (layer2_outputs(3426)) and not (layer2_outputs(5));
    layer3_outputs(321) <= layer2_outputs(4066);
    layer3_outputs(322) <= layer2_outputs(3453);
    layer3_outputs(323) <= not(layer2_outputs(5660)) or (layer2_outputs(3103));
    layer3_outputs(324) <= layer2_outputs(5408);
    layer3_outputs(325) <= '0';
    layer3_outputs(326) <= not(layer2_outputs(731));
    layer3_outputs(327) <= not(layer2_outputs(2248)) or (layer2_outputs(319));
    layer3_outputs(328) <= layer2_outputs(7338);
    layer3_outputs(329) <= (layer2_outputs(3068)) and not (layer2_outputs(4224));
    layer3_outputs(330) <= layer2_outputs(1471);
    layer3_outputs(331) <= not(layer2_outputs(1062));
    layer3_outputs(332) <= not(layer2_outputs(4472));
    layer3_outputs(333) <= not(layer2_outputs(7968));
    layer3_outputs(334) <= not(layer2_outputs(8443));
    layer3_outputs(335) <= not(layer2_outputs(6678));
    layer3_outputs(336) <= (layer2_outputs(7544)) and not (layer2_outputs(6965));
    layer3_outputs(337) <= layer2_outputs(8526);
    layer3_outputs(338) <= layer2_outputs(429);
    layer3_outputs(339) <= layer2_outputs(7151);
    layer3_outputs(340) <= not(layer2_outputs(589)) or (layer2_outputs(6386));
    layer3_outputs(341) <= (layer2_outputs(3059)) or (layer2_outputs(5911));
    layer3_outputs(342) <= not((layer2_outputs(2074)) xor (layer2_outputs(9931)));
    layer3_outputs(343) <= not(layer2_outputs(4300));
    layer3_outputs(344) <= (layer2_outputs(9214)) xor (layer2_outputs(2418));
    layer3_outputs(345) <= layer2_outputs(3810);
    layer3_outputs(346) <= not((layer2_outputs(668)) or (layer2_outputs(2528)));
    layer3_outputs(347) <= not((layer2_outputs(6477)) and (layer2_outputs(8664)));
    layer3_outputs(348) <= not(layer2_outputs(5987)) or (layer2_outputs(4478));
    layer3_outputs(349) <= (layer2_outputs(6836)) and not (layer2_outputs(5153));
    layer3_outputs(350) <= not(layer2_outputs(5125));
    layer3_outputs(351) <= not(layer2_outputs(4133));
    layer3_outputs(352) <= not(layer2_outputs(3493)) or (layer2_outputs(1938));
    layer3_outputs(353) <= layer2_outputs(4569);
    layer3_outputs(354) <= not(layer2_outputs(4637));
    layer3_outputs(355) <= not(layer2_outputs(741)) or (layer2_outputs(6960));
    layer3_outputs(356) <= '1';
    layer3_outputs(357) <= not((layer2_outputs(8371)) xor (layer2_outputs(1747)));
    layer3_outputs(358) <= not((layer2_outputs(3711)) or (layer2_outputs(1483)));
    layer3_outputs(359) <= (layer2_outputs(3608)) xor (layer2_outputs(6216));
    layer3_outputs(360) <= not((layer2_outputs(3845)) or (layer2_outputs(859)));
    layer3_outputs(361) <= not((layer2_outputs(3387)) or (layer2_outputs(3276)));
    layer3_outputs(362) <= not(layer2_outputs(6205));
    layer3_outputs(363) <= (layer2_outputs(7810)) and not (layer2_outputs(6341));
    layer3_outputs(364) <= not((layer2_outputs(910)) or (layer2_outputs(4630)));
    layer3_outputs(365) <= layer2_outputs(9118);
    layer3_outputs(366) <= (layer2_outputs(7777)) and not (layer2_outputs(2079));
    layer3_outputs(367) <= layer2_outputs(311);
    layer3_outputs(368) <= layer2_outputs(5775);
    layer3_outputs(369) <= not((layer2_outputs(2134)) or (layer2_outputs(4906)));
    layer3_outputs(370) <= not(layer2_outputs(641)) or (layer2_outputs(271));
    layer3_outputs(371) <= not(layer2_outputs(2686)) or (layer2_outputs(8454));
    layer3_outputs(372) <= layer2_outputs(6933);
    layer3_outputs(373) <= not((layer2_outputs(5042)) or (layer2_outputs(6597)));
    layer3_outputs(374) <= layer2_outputs(8373);
    layer3_outputs(375) <= not(layer2_outputs(8825));
    layer3_outputs(376) <= not((layer2_outputs(10160)) or (layer2_outputs(405)));
    layer3_outputs(377) <= not((layer2_outputs(289)) xor (layer2_outputs(6174)));
    layer3_outputs(378) <= (layer2_outputs(611)) and not (layer2_outputs(7068));
    layer3_outputs(379) <= not(layer2_outputs(978));
    layer3_outputs(380) <= not(layer2_outputs(5654));
    layer3_outputs(381) <= layer2_outputs(1711);
    layer3_outputs(382) <= layer2_outputs(6760);
    layer3_outputs(383) <= not(layer2_outputs(801));
    layer3_outputs(384) <= (layer2_outputs(7427)) xor (layer2_outputs(6139));
    layer3_outputs(385) <= not(layer2_outputs(7549)) or (layer2_outputs(7093));
    layer3_outputs(386) <= not(layer2_outputs(1336));
    layer3_outputs(387) <= not((layer2_outputs(9834)) or (layer2_outputs(1978)));
    layer3_outputs(388) <= not(layer2_outputs(2176));
    layer3_outputs(389) <= (layer2_outputs(1877)) and not (layer2_outputs(1053));
    layer3_outputs(390) <= (layer2_outputs(4866)) and not (layer2_outputs(9810));
    layer3_outputs(391) <= layer2_outputs(2348);
    layer3_outputs(392) <= not((layer2_outputs(2187)) and (layer2_outputs(2599)));
    layer3_outputs(393) <= layer2_outputs(6307);
    layer3_outputs(394) <= not((layer2_outputs(4963)) xor (layer2_outputs(9994)));
    layer3_outputs(395) <= (layer2_outputs(1183)) or (layer2_outputs(6268));
    layer3_outputs(396) <= not((layer2_outputs(2002)) and (layer2_outputs(5457)));
    layer3_outputs(397) <= layer2_outputs(3602);
    layer3_outputs(398) <= layer2_outputs(2771);
    layer3_outputs(399) <= '1';
    layer3_outputs(400) <= not((layer2_outputs(3049)) or (layer2_outputs(9436)));
    layer3_outputs(401) <= (layer2_outputs(2517)) or (layer2_outputs(4186));
    layer3_outputs(402) <= (layer2_outputs(3183)) or (layer2_outputs(440));
    layer3_outputs(403) <= layer2_outputs(4368);
    layer3_outputs(404) <= layer2_outputs(789);
    layer3_outputs(405) <= layer2_outputs(2636);
    layer3_outputs(406) <= (layer2_outputs(9503)) and (layer2_outputs(6404));
    layer3_outputs(407) <= not(layer2_outputs(7935));
    layer3_outputs(408) <= not(layer2_outputs(7104));
    layer3_outputs(409) <= not(layer2_outputs(1928)) or (layer2_outputs(4677));
    layer3_outputs(410) <= (layer2_outputs(7543)) and not (layer2_outputs(7050));
    layer3_outputs(411) <= not(layer2_outputs(10121));
    layer3_outputs(412) <= not((layer2_outputs(6494)) and (layer2_outputs(9541)));
    layer3_outputs(413) <= (layer2_outputs(2243)) and not (layer2_outputs(1213));
    layer3_outputs(414) <= layer2_outputs(8293);
    layer3_outputs(415) <= not(layer2_outputs(8507));
    layer3_outputs(416) <= not((layer2_outputs(7714)) or (layer2_outputs(7754)));
    layer3_outputs(417) <= not((layer2_outputs(8565)) or (layer2_outputs(2153)));
    layer3_outputs(418) <= layer2_outputs(8374);
    layer3_outputs(419) <= not((layer2_outputs(6248)) xor (layer2_outputs(4238)));
    layer3_outputs(420) <= (layer2_outputs(5839)) and not (layer2_outputs(3992));
    layer3_outputs(421) <= '1';
    layer3_outputs(422) <= not(layer2_outputs(4769)) or (layer2_outputs(1661));
    layer3_outputs(423) <= (layer2_outputs(2764)) or (layer2_outputs(6535));
    layer3_outputs(424) <= not((layer2_outputs(4117)) xor (layer2_outputs(8415)));
    layer3_outputs(425) <= layer2_outputs(8739);
    layer3_outputs(426) <= not((layer2_outputs(6594)) xor (layer2_outputs(5701)));
    layer3_outputs(427) <= not(layer2_outputs(4316)) or (layer2_outputs(9726));
    layer3_outputs(428) <= layer2_outputs(2074);
    layer3_outputs(429) <= (layer2_outputs(5013)) xor (layer2_outputs(2222));
    layer3_outputs(430) <= not(layer2_outputs(4563));
    layer3_outputs(431) <= not((layer2_outputs(9505)) or (layer2_outputs(3362)));
    layer3_outputs(432) <= not((layer2_outputs(593)) xor (layer2_outputs(8562)));
    layer3_outputs(433) <= '0';
    layer3_outputs(434) <= (layer2_outputs(6504)) xor (layer2_outputs(3805));
    layer3_outputs(435) <= (layer2_outputs(540)) and not (layer2_outputs(6615));
    layer3_outputs(436) <= '0';
    layer3_outputs(437) <= not((layer2_outputs(982)) and (layer2_outputs(9691)));
    layer3_outputs(438) <= (layer2_outputs(1695)) and (layer2_outputs(698));
    layer3_outputs(439) <= not((layer2_outputs(2238)) xor (layer2_outputs(5317)));
    layer3_outputs(440) <= not(layer2_outputs(430)) or (layer2_outputs(9431));
    layer3_outputs(441) <= not(layer2_outputs(4444));
    layer3_outputs(442) <= layer2_outputs(4874);
    layer3_outputs(443) <= (layer2_outputs(3619)) and (layer2_outputs(5341));
    layer3_outputs(444) <= layer2_outputs(2726);
    layer3_outputs(445) <= not(layer2_outputs(1996));
    layer3_outputs(446) <= not(layer2_outputs(3675)) or (layer2_outputs(7482));
    layer3_outputs(447) <= layer2_outputs(6007);
    layer3_outputs(448) <= not(layer2_outputs(6431)) or (layer2_outputs(1977));
    layer3_outputs(449) <= layer2_outputs(863);
    layer3_outputs(450) <= (layer2_outputs(6246)) or (layer2_outputs(8112));
    layer3_outputs(451) <= (layer2_outputs(5962)) xor (layer2_outputs(2568));
    layer3_outputs(452) <= not((layer2_outputs(1169)) xor (layer2_outputs(6985)));
    layer3_outputs(453) <= not(layer2_outputs(4041)) or (layer2_outputs(2260));
    layer3_outputs(454) <= '1';
    layer3_outputs(455) <= (layer2_outputs(6190)) xor (layer2_outputs(6511));
    layer3_outputs(456) <= layer2_outputs(2856);
    layer3_outputs(457) <= (layer2_outputs(2401)) or (layer2_outputs(599));
    layer3_outputs(458) <= layer2_outputs(9225);
    layer3_outputs(459) <= (layer2_outputs(9182)) or (layer2_outputs(10123));
    layer3_outputs(460) <= not((layer2_outputs(3835)) and (layer2_outputs(8510)));
    layer3_outputs(461) <= layer2_outputs(7826);
    layer3_outputs(462) <= (layer2_outputs(5347)) and (layer2_outputs(2319));
    layer3_outputs(463) <= not(layer2_outputs(1047));
    layer3_outputs(464) <= '1';
    layer3_outputs(465) <= layer2_outputs(7726);
    layer3_outputs(466) <= not((layer2_outputs(1694)) xor (layer2_outputs(3927)));
    layer3_outputs(467) <= not(layer2_outputs(1862)) or (layer2_outputs(3878));
    layer3_outputs(468) <= layer2_outputs(1801);
    layer3_outputs(469) <= layer2_outputs(5823);
    layer3_outputs(470) <= not((layer2_outputs(8270)) or (layer2_outputs(7349)));
    layer3_outputs(471) <= not(layer2_outputs(2781));
    layer3_outputs(472) <= (layer2_outputs(249)) xor (layer2_outputs(1995));
    layer3_outputs(473) <= (layer2_outputs(3090)) xor (layer2_outputs(3558));
    layer3_outputs(474) <= not((layer2_outputs(213)) xor (layer2_outputs(9194)));
    layer3_outputs(475) <= not(layer2_outputs(2820));
    layer3_outputs(476) <= not(layer2_outputs(6759));
    layer3_outputs(477) <= not((layer2_outputs(2463)) and (layer2_outputs(7464)));
    layer3_outputs(478) <= layer2_outputs(1192);
    layer3_outputs(479) <= not(layer2_outputs(2480));
    layer3_outputs(480) <= not(layer2_outputs(4314)) or (layer2_outputs(2052));
    layer3_outputs(481) <= not(layer2_outputs(5974));
    layer3_outputs(482) <= not(layer2_outputs(2126));
    layer3_outputs(483) <= (layer2_outputs(2812)) and not (layer2_outputs(3893));
    layer3_outputs(484) <= '0';
    layer3_outputs(485) <= layer2_outputs(3788);
    layer3_outputs(486) <= (layer2_outputs(7512)) and not (layer2_outputs(2434));
    layer3_outputs(487) <= not((layer2_outputs(4036)) or (layer2_outputs(3032)));
    layer3_outputs(488) <= (layer2_outputs(8868)) and (layer2_outputs(9991));
    layer3_outputs(489) <= (layer2_outputs(4433)) xor (layer2_outputs(2611));
    layer3_outputs(490) <= layer2_outputs(314);
    layer3_outputs(491) <= (layer2_outputs(5413)) and not (layer2_outputs(7425));
    layer3_outputs(492) <= (layer2_outputs(1313)) and not (layer2_outputs(4371));
    layer3_outputs(493) <= not((layer2_outputs(1707)) or (layer2_outputs(1963)));
    layer3_outputs(494) <= '0';
    layer3_outputs(495) <= (layer2_outputs(6411)) xor (layer2_outputs(5392));
    layer3_outputs(496) <= (layer2_outputs(9164)) and not (layer2_outputs(6221));
    layer3_outputs(497) <= not(layer2_outputs(7927));
    layer3_outputs(498) <= not(layer2_outputs(3095));
    layer3_outputs(499) <= (layer2_outputs(7551)) or (layer2_outputs(735));
    layer3_outputs(500) <= not((layer2_outputs(281)) and (layer2_outputs(6990)));
    layer3_outputs(501) <= layer2_outputs(3389);
    layer3_outputs(502) <= (layer2_outputs(9141)) and not (layer2_outputs(5101));
    layer3_outputs(503) <= not((layer2_outputs(9542)) xor (layer2_outputs(2392)));
    layer3_outputs(504) <= layer2_outputs(4207);
    layer3_outputs(505) <= layer2_outputs(4486);
    layer3_outputs(506) <= (layer2_outputs(2008)) and not (layer2_outputs(3211));
    layer3_outputs(507) <= (layer2_outputs(2547)) or (layer2_outputs(7359));
    layer3_outputs(508) <= layer2_outputs(116);
    layer3_outputs(509) <= not((layer2_outputs(9862)) xor (layer2_outputs(5086)));
    layer3_outputs(510) <= not((layer2_outputs(10170)) or (layer2_outputs(2582)));
    layer3_outputs(511) <= layer2_outputs(4981);
    layer3_outputs(512) <= not(layer2_outputs(4699));
    layer3_outputs(513) <= (layer2_outputs(5693)) and not (layer2_outputs(8117));
    layer3_outputs(514) <= not(layer2_outputs(3609));
    layer3_outputs(515) <= not(layer2_outputs(3207)) or (layer2_outputs(2934));
    layer3_outputs(516) <= (layer2_outputs(8078)) and not (layer2_outputs(4199));
    layer3_outputs(517) <= layer2_outputs(2873);
    layer3_outputs(518) <= (layer2_outputs(4205)) and not (layer2_outputs(4644));
    layer3_outputs(519) <= not(layer2_outputs(2866));
    layer3_outputs(520) <= not(layer2_outputs(9068)) or (layer2_outputs(8851));
    layer3_outputs(521) <= not(layer2_outputs(8145));
    layer3_outputs(522) <= not(layer2_outputs(5132));
    layer3_outputs(523) <= '1';
    layer3_outputs(524) <= not(layer2_outputs(1980));
    layer3_outputs(525) <= layer2_outputs(878);
    layer3_outputs(526) <= not(layer2_outputs(666));
    layer3_outputs(527) <= layer2_outputs(872);
    layer3_outputs(528) <= not((layer2_outputs(5193)) xor (layer2_outputs(1279)));
    layer3_outputs(529) <= (layer2_outputs(4711)) and not (layer2_outputs(36));
    layer3_outputs(530) <= layer2_outputs(4895);
    layer3_outputs(531) <= layer2_outputs(7020);
    layer3_outputs(532) <= layer2_outputs(6773);
    layer3_outputs(533) <= not((layer2_outputs(993)) xor (layer2_outputs(9443)));
    layer3_outputs(534) <= (layer2_outputs(3935)) and not (layer2_outputs(6097));
    layer3_outputs(535) <= layer2_outputs(6466);
    layer3_outputs(536) <= not(layer2_outputs(9282));
    layer3_outputs(537) <= not(layer2_outputs(6720)) or (layer2_outputs(3394));
    layer3_outputs(538) <= not(layer2_outputs(9873)) or (layer2_outputs(8357));
    layer3_outputs(539) <= not(layer2_outputs(3184));
    layer3_outputs(540) <= (layer2_outputs(4924)) and not (layer2_outputs(1331));
    layer3_outputs(541) <= not(layer2_outputs(9883));
    layer3_outputs(542) <= not(layer2_outputs(4697)) or (layer2_outputs(2647));
    layer3_outputs(543) <= not((layer2_outputs(8226)) xor (layer2_outputs(2905)));
    layer3_outputs(544) <= layer2_outputs(8824);
    layer3_outputs(545) <= layer2_outputs(2723);
    layer3_outputs(546) <= (layer2_outputs(3367)) or (layer2_outputs(6196));
    layer3_outputs(547) <= not((layer2_outputs(8437)) and (layer2_outputs(3054)));
    layer3_outputs(548) <= not(layer2_outputs(6930));
    layer3_outputs(549) <= layer2_outputs(7220);
    layer3_outputs(550) <= (layer2_outputs(1846)) and not (layer2_outputs(9501));
    layer3_outputs(551) <= (layer2_outputs(7959)) and not (layer2_outputs(5477));
    layer3_outputs(552) <= (layer2_outputs(853)) and not (layer2_outputs(2093));
    layer3_outputs(553) <= not(layer2_outputs(9173));
    layer3_outputs(554) <= '0';
    layer3_outputs(555) <= (layer2_outputs(8984)) and not (layer2_outputs(4632));
    layer3_outputs(556) <= not(layer2_outputs(2968));
    layer3_outputs(557) <= (layer2_outputs(8819)) and (layer2_outputs(3389));
    layer3_outputs(558) <= not((layer2_outputs(8492)) or (layer2_outputs(6697)));
    layer3_outputs(559) <= not(layer2_outputs(2860)) or (layer2_outputs(2658));
    layer3_outputs(560) <= (layer2_outputs(7692)) and not (layer2_outputs(1932));
    layer3_outputs(561) <= not((layer2_outputs(7952)) or (layer2_outputs(9583)));
    layer3_outputs(562) <= (layer2_outputs(5614)) and not (layer2_outputs(9490));
    layer3_outputs(563) <= layer2_outputs(9039);
    layer3_outputs(564) <= not((layer2_outputs(1260)) or (layer2_outputs(4521)));
    layer3_outputs(565) <= not(layer2_outputs(142));
    layer3_outputs(566) <= not(layer2_outputs(4615));
    layer3_outputs(567) <= layer2_outputs(6324);
    layer3_outputs(568) <= not(layer2_outputs(1777));
    layer3_outputs(569) <= (layer2_outputs(1567)) and not (layer2_outputs(5740));
    layer3_outputs(570) <= not(layer2_outputs(8979));
    layer3_outputs(571) <= (layer2_outputs(906)) or (layer2_outputs(3279));
    layer3_outputs(572) <= not((layer2_outputs(2202)) or (layer2_outputs(160)));
    layer3_outputs(573) <= '0';
    layer3_outputs(574) <= not(layer2_outputs(6800));
    layer3_outputs(575) <= not(layer2_outputs(998)) or (layer2_outputs(3020));
    layer3_outputs(576) <= layer2_outputs(5701);
    layer3_outputs(577) <= not(layer2_outputs(2689));
    layer3_outputs(578) <= not(layer2_outputs(4136));
    layer3_outputs(579) <= not(layer2_outputs(305)) or (layer2_outputs(3332));
    layer3_outputs(580) <= not(layer2_outputs(6035));
    layer3_outputs(581) <= (layer2_outputs(7985)) or (layer2_outputs(2596));
    layer3_outputs(582) <= (layer2_outputs(9114)) and not (layer2_outputs(5208));
    layer3_outputs(583) <= (layer2_outputs(3665)) xor (layer2_outputs(5399));
    layer3_outputs(584) <= (layer2_outputs(585)) xor (layer2_outputs(1652));
    layer3_outputs(585) <= layer2_outputs(3440);
    layer3_outputs(586) <= not(layer2_outputs(9001)) or (layer2_outputs(5759));
    layer3_outputs(587) <= layer2_outputs(3914);
    layer3_outputs(588) <= not(layer2_outputs(8567));
    layer3_outputs(589) <= layer2_outputs(9463);
    layer3_outputs(590) <= layer2_outputs(8411);
    layer3_outputs(591) <= '0';
    layer3_outputs(592) <= not(layer2_outputs(5534)) or (layer2_outputs(7788));
    layer3_outputs(593) <= not((layer2_outputs(2622)) and (layer2_outputs(4420)));
    layer3_outputs(594) <= not(layer2_outputs(2605)) or (layer2_outputs(8261));
    layer3_outputs(595) <= layer2_outputs(2588);
    layer3_outputs(596) <= layer2_outputs(3181);
    layer3_outputs(597) <= layer2_outputs(8104);
    layer3_outputs(598) <= (layer2_outputs(10024)) and (layer2_outputs(9479));
    layer3_outputs(599) <= layer2_outputs(4429);
    layer3_outputs(600) <= layer2_outputs(1060);
    layer3_outputs(601) <= '1';
    layer3_outputs(602) <= layer2_outputs(2267);
    layer3_outputs(603) <= not(layer2_outputs(7992)) or (layer2_outputs(8943));
    layer3_outputs(604) <= layer2_outputs(9548);
    layer3_outputs(605) <= not((layer2_outputs(8004)) xor (layer2_outputs(9777)));
    layer3_outputs(606) <= layer2_outputs(7806);
    layer3_outputs(607) <= layer2_outputs(696);
    layer3_outputs(608) <= layer2_outputs(4933);
    layer3_outputs(609) <= (layer2_outputs(7840)) xor (layer2_outputs(2244));
    layer3_outputs(610) <= '1';
    layer3_outputs(611) <= (layer2_outputs(4013)) and (layer2_outputs(9512));
    layer3_outputs(612) <= layer2_outputs(204);
    layer3_outputs(613) <= not(layer2_outputs(7195));
    layer3_outputs(614) <= not(layer2_outputs(8935));
    layer3_outputs(615) <= layer2_outputs(5063);
    layer3_outputs(616) <= not(layer2_outputs(2322));
    layer3_outputs(617) <= layer2_outputs(10169);
    layer3_outputs(618) <= layer2_outputs(1219);
    layer3_outputs(619) <= not(layer2_outputs(3054));
    layer3_outputs(620) <= not(layer2_outputs(9835));
    layer3_outputs(621) <= layer2_outputs(5572);
    layer3_outputs(622) <= not(layer2_outputs(5256));
    layer3_outputs(623) <= not((layer2_outputs(2246)) or (layer2_outputs(4197)));
    layer3_outputs(624) <= (layer2_outputs(1484)) and not (layer2_outputs(9309));
    layer3_outputs(625) <= not(layer2_outputs(4189));
    layer3_outputs(626) <= (layer2_outputs(8999)) or (layer2_outputs(6432));
    layer3_outputs(627) <= (layer2_outputs(2859)) xor (layer2_outputs(234));
    layer3_outputs(628) <= (layer2_outputs(2308)) xor (layer2_outputs(9243));
    layer3_outputs(629) <= (layer2_outputs(8334)) xor (layer2_outputs(4715));
    layer3_outputs(630) <= (layer2_outputs(3871)) and (layer2_outputs(3261));
    layer3_outputs(631) <= layer2_outputs(5966);
    layer3_outputs(632) <= layer2_outputs(4600);
    layer3_outputs(633) <= not((layer2_outputs(7322)) or (layer2_outputs(4476)));
    layer3_outputs(634) <= not(layer2_outputs(9266));
    layer3_outputs(635) <= not(layer2_outputs(8381)) or (layer2_outputs(1638));
    layer3_outputs(636) <= not((layer2_outputs(9747)) xor (layer2_outputs(3645)));
    layer3_outputs(637) <= not(layer2_outputs(3976));
    layer3_outputs(638) <= not(layer2_outputs(8561)) or (layer2_outputs(8195));
    layer3_outputs(639) <= not(layer2_outputs(7854));
    layer3_outputs(640) <= layer2_outputs(8970);
    layer3_outputs(641) <= layer2_outputs(4222);
    layer3_outputs(642) <= not(layer2_outputs(6707));
    layer3_outputs(643) <= not(layer2_outputs(2354));
    layer3_outputs(644) <= not(layer2_outputs(3517)) or (layer2_outputs(1022));
    layer3_outputs(645) <= layer2_outputs(9275);
    layer3_outputs(646) <= not(layer2_outputs(6095));
    layer3_outputs(647) <= layer2_outputs(6947);
    layer3_outputs(648) <= not(layer2_outputs(9586));
    layer3_outputs(649) <= not(layer2_outputs(1570));
    layer3_outputs(650) <= (layer2_outputs(2233)) xor (layer2_outputs(6323));
    layer3_outputs(651) <= not(layer2_outputs(4945));
    layer3_outputs(652) <= layer2_outputs(7915);
    layer3_outputs(653) <= not(layer2_outputs(7603));
    layer3_outputs(654) <= (layer2_outputs(6256)) and not (layer2_outputs(3119));
    layer3_outputs(655) <= (layer2_outputs(4628)) and not (layer2_outputs(6448));
    layer3_outputs(656) <= (layer2_outputs(4165)) xor (layer2_outputs(4529));
    layer3_outputs(657) <= not(layer2_outputs(5181));
    layer3_outputs(658) <= (layer2_outputs(6318)) and (layer2_outputs(3189));
    layer3_outputs(659) <= not(layer2_outputs(798));
    layer3_outputs(660) <= not(layer2_outputs(6238)) or (layer2_outputs(2211));
    layer3_outputs(661) <= layer2_outputs(6512);
    layer3_outputs(662) <= not((layer2_outputs(862)) xor (layer2_outputs(8064)));
    layer3_outputs(663) <= not(layer2_outputs(5021));
    layer3_outputs(664) <= not(layer2_outputs(238));
    layer3_outputs(665) <= (layer2_outputs(6975)) and not (layer2_outputs(7386));
    layer3_outputs(666) <= layer2_outputs(6041);
    layer3_outputs(667) <= not(layer2_outputs(8052));
    layer3_outputs(668) <= not(layer2_outputs(8724));
    layer3_outputs(669) <= layer2_outputs(3250);
    layer3_outputs(670) <= layer2_outputs(3040);
    layer3_outputs(671) <= not((layer2_outputs(6465)) or (layer2_outputs(2991)));
    layer3_outputs(672) <= not(layer2_outputs(1730)) or (layer2_outputs(1611));
    layer3_outputs(673) <= (layer2_outputs(4334)) and (layer2_outputs(5213));
    layer3_outputs(674) <= layer2_outputs(7412);
    layer3_outputs(675) <= not(layer2_outputs(4524));
    layer3_outputs(676) <= (layer2_outputs(10015)) or (layer2_outputs(4932));
    layer3_outputs(677) <= not(layer2_outputs(8454));
    layer3_outputs(678) <= layer2_outputs(7283);
    layer3_outputs(679) <= layer2_outputs(1711);
    layer3_outputs(680) <= (layer2_outputs(5890)) and not (layer2_outputs(3297));
    layer3_outputs(681) <= layer2_outputs(9285);
    layer3_outputs(682) <= not(layer2_outputs(9810));
    layer3_outputs(683) <= not(layer2_outputs(7439));
    layer3_outputs(684) <= layer2_outputs(3568);
    layer3_outputs(685) <= (layer2_outputs(10093)) and (layer2_outputs(8420));
    layer3_outputs(686) <= not(layer2_outputs(9714));
    layer3_outputs(687) <= not((layer2_outputs(5528)) xor (layer2_outputs(7873)));
    layer3_outputs(688) <= not(layer2_outputs(126));
    layer3_outputs(689) <= not(layer2_outputs(5873));
    layer3_outputs(690) <= '1';
    layer3_outputs(691) <= layer2_outputs(7531);
    layer3_outputs(692) <= (layer2_outputs(6092)) or (layer2_outputs(3252));
    layer3_outputs(693) <= layer2_outputs(9731);
    layer3_outputs(694) <= (layer2_outputs(756)) xor (layer2_outputs(8929));
    layer3_outputs(695) <= not(layer2_outputs(1457)) or (layer2_outputs(4633));
    layer3_outputs(696) <= layer2_outputs(9363);
    layer3_outputs(697) <= not(layer2_outputs(8251));
    layer3_outputs(698) <= layer2_outputs(3142);
    layer3_outputs(699) <= not(layer2_outputs(5415));
    layer3_outputs(700) <= layer2_outputs(166);
    layer3_outputs(701) <= not(layer2_outputs(3498)) or (layer2_outputs(5286));
    layer3_outputs(702) <= not((layer2_outputs(9624)) and (layer2_outputs(2564)));
    layer3_outputs(703) <= not(layer2_outputs(3460));
    layer3_outputs(704) <= not((layer2_outputs(7083)) or (layer2_outputs(2627)));
    layer3_outputs(705) <= not(layer2_outputs(7635));
    layer3_outputs(706) <= '0';
    layer3_outputs(707) <= (layer2_outputs(1526)) and not (layer2_outputs(6812));
    layer3_outputs(708) <= not(layer2_outputs(1551));
    layer3_outputs(709) <= layer2_outputs(9625);
    layer3_outputs(710) <= layer2_outputs(94);
    layer3_outputs(711) <= layer2_outputs(8280);
    layer3_outputs(712) <= layer2_outputs(1277);
    layer3_outputs(713) <= not(layer2_outputs(1581)) or (layer2_outputs(9611));
    layer3_outputs(714) <= (layer2_outputs(1712)) and not (layer2_outputs(8246));
    layer3_outputs(715) <= not((layer2_outputs(5325)) and (layer2_outputs(3877)));
    layer3_outputs(716) <= not(layer2_outputs(9112));
    layer3_outputs(717) <= not(layer2_outputs(3504));
    layer3_outputs(718) <= layer2_outputs(8848);
    layer3_outputs(719) <= layer2_outputs(7341);
    layer3_outputs(720) <= '0';
    layer3_outputs(721) <= not(layer2_outputs(2257)) or (layer2_outputs(1369));
    layer3_outputs(722) <= (layer2_outputs(9083)) xor (layer2_outputs(5604));
    layer3_outputs(723) <= (layer2_outputs(3418)) and not (layer2_outputs(7455));
    layer3_outputs(724) <= '1';
    layer3_outputs(725) <= not(layer2_outputs(3493));
    layer3_outputs(726) <= layer2_outputs(5782);
    layer3_outputs(727) <= layer2_outputs(3754);
    layer3_outputs(728) <= not(layer2_outputs(6996));
    layer3_outputs(729) <= layer2_outputs(6019);
    layer3_outputs(730) <= (layer2_outputs(9434)) and not (layer2_outputs(9255));
    layer3_outputs(731) <= not(layer2_outputs(7430)) or (layer2_outputs(5956));
    layer3_outputs(732) <= not(layer2_outputs(3115)) or (layer2_outputs(4482));
    layer3_outputs(733) <= layer2_outputs(2822);
    layer3_outputs(734) <= layer2_outputs(6774);
    layer3_outputs(735) <= not((layer2_outputs(8705)) or (layer2_outputs(1123)));
    layer3_outputs(736) <= layer2_outputs(2182);
    layer3_outputs(737) <= '1';
    layer3_outputs(738) <= not(layer2_outputs(8560)) or (layer2_outputs(7160));
    layer3_outputs(739) <= not(layer2_outputs(5059));
    layer3_outputs(740) <= layer2_outputs(2983);
    layer3_outputs(741) <= layer2_outputs(5593);
    layer3_outputs(742) <= not(layer2_outputs(3688)) or (layer2_outputs(2000));
    layer3_outputs(743) <= (layer2_outputs(4237)) xor (layer2_outputs(1696));
    layer3_outputs(744) <= (layer2_outputs(5411)) and (layer2_outputs(3546));
    layer3_outputs(745) <= not(layer2_outputs(9272));
    layer3_outputs(746) <= layer2_outputs(5526);
    layer3_outputs(747) <= not((layer2_outputs(8125)) xor (layer2_outputs(5635)));
    layer3_outputs(748) <= (layer2_outputs(1312)) and not (layer2_outputs(7835));
    layer3_outputs(749) <= (layer2_outputs(4383)) and not (layer2_outputs(5759));
    layer3_outputs(750) <= '0';
    layer3_outputs(751) <= not((layer2_outputs(8769)) and (layer2_outputs(8623)));
    layer3_outputs(752) <= (layer2_outputs(371)) xor (layer2_outputs(1500));
    layer3_outputs(753) <= (layer2_outputs(44)) and not (layer2_outputs(7861));
    layer3_outputs(754) <= not(layer2_outputs(9340));
    layer3_outputs(755) <= not((layer2_outputs(6669)) or (layer2_outputs(3406)));
    layer3_outputs(756) <= not((layer2_outputs(1527)) and (layer2_outputs(8734)));
    layer3_outputs(757) <= (layer2_outputs(6330)) and (layer2_outputs(1794));
    layer3_outputs(758) <= (layer2_outputs(5019)) and not (layer2_outputs(6740));
    layer3_outputs(759) <= not(layer2_outputs(9527));
    layer3_outputs(760) <= not(layer2_outputs(8069));
    layer3_outputs(761) <= not(layer2_outputs(764));
    layer3_outputs(762) <= not(layer2_outputs(929));
    layer3_outputs(763) <= not(layer2_outputs(8235));
    layer3_outputs(764) <= not(layer2_outputs(576));
    layer3_outputs(765) <= (layer2_outputs(3462)) and not (layer2_outputs(5624));
    layer3_outputs(766) <= layer2_outputs(3094);
    layer3_outputs(767) <= (layer2_outputs(2594)) and not (layer2_outputs(9400));
    layer3_outputs(768) <= not(layer2_outputs(4236));
    layer3_outputs(769) <= not((layer2_outputs(3204)) xor (layer2_outputs(4612)));
    layer3_outputs(770) <= (layer2_outputs(5977)) and (layer2_outputs(3353));
    layer3_outputs(771) <= not((layer2_outputs(4370)) xor (layer2_outputs(782)));
    layer3_outputs(772) <= (layer2_outputs(4683)) and not (layer2_outputs(2740));
    layer3_outputs(773) <= not((layer2_outputs(623)) or (layer2_outputs(9698)));
    layer3_outputs(774) <= '1';
    layer3_outputs(775) <= (layer2_outputs(1967)) xor (layer2_outputs(9482));
    layer3_outputs(776) <= (layer2_outputs(7287)) xor (layer2_outputs(6416));
    layer3_outputs(777) <= not(layer2_outputs(4096));
    layer3_outputs(778) <= not((layer2_outputs(2665)) xor (layer2_outputs(6617)));
    layer3_outputs(779) <= (layer2_outputs(1865)) or (layer2_outputs(4410));
    layer3_outputs(780) <= not((layer2_outputs(9510)) xor (layer2_outputs(6731)));
    layer3_outputs(781) <= layer2_outputs(9242);
    layer3_outputs(782) <= (layer2_outputs(4589)) and not (layer2_outputs(9567));
    layer3_outputs(783) <= (layer2_outputs(2346)) or (layer2_outputs(8284));
    layer3_outputs(784) <= not(layer2_outputs(7879)) or (layer2_outputs(5444));
    layer3_outputs(785) <= not((layer2_outputs(2602)) xor (layer2_outputs(7680)));
    layer3_outputs(786) <= layer2_outputs(6242);
    layer3_outputs(787) <= layer2_outputs(2566);
    layer3_outputs(788) <= (layer2_outputs(8706)) and not (layer2_outputs(4802));
    layer3_outputs(789) <= layer2_outputs(8568);
    layer3_outputs(790) <= '1';
    layer3_outputs(791) <= not((layer2_outputs(8513)) or (layer2_outputs(8758)));
    layer3_outputs(792) <= (layer2_outputs(6868)) and not (layer2_outputs(10120));
    layer3_outputs(793) <= (layer2_outputs(9894)) and not (layer2_outputs(2966));
    layer3_outputs(794) <= not(layer2_outputs(93));
    layer3_outputs(795) <= not((layer2_outputs(8313)) or (layer2_outputs(4636)));
    layer3_outputs(796) <= (layer2_outputs(290)) or (layer2_outputs(5831));
    layer3_outputs(797) <= (layer2_outputs(2262)) and not (layer2_outputs(9435));
    layer3_outputs(798) <= layer2_outputs(4617);
    layer3_outputs(799) <= layer2_outputs(581);
    layer3_outputs(800) <= layer2_outputs(7857);
    layer3_outputs(801) <= not(layer2_outputs(4894));
    layer3_outputs(802) <= layer2_outputs(9555);
    layer3_outputs(803) <= (layer2_outputs(2049)) or (layer2_outputs(9749));
    layer3_outputs(804) <= (layer2_outputs(8824)) xor (layer2_outputs(3646));
    layer3_outputs(805) <= layer2_outputs(9117);
    layer3_outputs(806) <= not(layer2_outputs(1780));
    layer3_outputs(807) <= (layer2_outputs(4161)) and not (layer2_outputs(6789));
    layer3_outputs(808) <= '0';
    layer3_outputs(809) <= layer2_outputs(7078);
    layer3_outputs(810) <= not(layer2_outputs(6501));
    layer3_outputs(811) <= not(layer2_outputs(5248)) or (layer2_outputs(787));
    layer3_outputs(812) <= not(layer2_outputs(5414));
    layer3_outputs(813) <= layer2_outputs(9466);
    layer3_outputs(814) <= layer2_outputs(5146);
    layer3_outputs(815) <= not((layer2_outputs(7920)) or (layer2_outputs(6284)));
    layer3_outputs(816) <= not(layer2_outputs(3438));
    layer3_outputs(817) <= not(layer2_outputs(3031));
    layer3_outputs(818) <= '0';
    layer3_outputs(819) <= layer2_outputs(3244);
    layer3_outputs(820) <= not(layer2_outputs(6925));
    layer3_outputs(821) <= (layer2_outputs(6447)) or (layer2_outputs(4778));
    layer3_outputs(822) <= layer2_outputs(5662);
    layer3_outputs(823) <= not(layer2_outputs(2199));
    layer3_outputs(824) <= (layer2_outputs(5963)) and (layer2_outputs(33));
    layer3_outputs(825) <= layer2_outputs(455);
    layer3_outputs(826) <= (layer2_outputs(8966)) or (layer2_outputs(684));
    layer3_outputs(827) <= layer2_outputs(7958);
    layer3_outputs(828) <= layer2_outputs(9860);
    layer3_outputs(829) <= (layer2_outputs(9858)) and not (layer2_outputs(8005));
    layer3_outputs(830) <= layer2_outputs(8782);
    layer3_outputs(831) <= not(layer2_outputs(10028));
    layer3_outputs(832) <= layer2_outputs(5616);
    layer3_outputs(833) <= '1';
    layer3_outputs(834) <= (layer2_outputs(7718)) and (layer2_outputs(1829));
    layer3_outputs(835) <= '1';
    layer3_outputs(836) <= not((layer2_outputs(8016)) or (layer2_outputs(4469)));
    layer3_outputs(837) <= (layer2_outputs(1488)) and (layer2_outputs(8698));
    layer3_outputs(838) <= '0';
    layer3_outputs(839) <= (layer2_outputs(9517)) or (layer2_outputs(8893));
    layer3_outputs(840) <= layer2_outputs(2297);
    layer3_outputs(841) <= not(layer2_outputs(9227)) or (layer2_outputs(10168));
    layer3_outputs(842) <= layer2_outputs(4952);
    layer3_outputs(843) <= '0';
    layer3_outputs(844) <= not(layer2_outputs(395)) or (layer2_outputs(818));
    layer3_outputs(845) <= not(layer2_outputs(733));
    layer3_outputs(846) <= not(layer2_outputs(1314));
    layer3_outputs(847) <= '1';
    layer3_outputs(848) <= not((layer2_outputs(2377)) or (layer2_outputs(779)));
    layer3_outputs(849) <= (layer2_outputs(5915)) or (layer2_outputs(8250));
    layer3_outputs(850) <= '0';
    layer3_outputs(851) <= (layer2_outputs(6009)) and (layer2_outputs(109));
    layer3_outputs(852) <= '1';
    layer3_outputs(853) <= not((layer2_outputs(5953)) and (layer2_outputs(6487)));
    layer3_outputs(854) <= not((layer2_outputs(2237)) or (layer2_outputs(720)));
    layer3_outputs(855) <= not((layer2_outputs(8345)) xor (layer2_outputs(4892)));
    layer3_outputs(856) <= layer2_outputs(1628);
    layer3_outputs(857) <= (layer2_outputs(4778)) xor (layer2_outputs(3638));
    layer3_outputs(858) <= not(layer2_outputs(8262));
    layer3_outputs(859) <= (layer2_outputs(8091)) xor (layer2_outputs(3343));
    layer3_outputs(860) <= (layer2_outputs(8711)) and not (layer2_outputs(895));
    layer3_outputs(861) <= layer2_outputs(6573);
    layer3_outputs(862) <= (layer2_outputs(4859)) and not (layer2_outputs(6075));
    layer3_outputs(863) <= (layer2_outputs(6725)) and (layer2_outputs(851));
    layer3_outputs(864) <= layer2_outputs(6163);
    layer3_outputs(865) <= layer2_outputs(5847);
    layer3_outputs(866) <= '0';
    layer3_outputs(867) <= not((layer2_outputs(5070)) and (layer2_outputs(9042)));
    layer3_outputs(868) <= layer2_outputs(4300);
    layer3_outputs(869) <= layer2_outputs(9428);
    layer3_outputs(870) <= not(layer2_outputs(5248));
    layer3_outputs(871) <= not(layer2_outputs(8461)) or (layer2_outputs(4056));
    layer3_outputs(872) <= not(layer2_outputs(3187)) or (layer2_outputs(8652));
    layer3_outputs(873) <= layer2_outputs(9455);
    layer3_outputs(874) <= not((layer2_outputs(5828)) or (layer2_outputs(10040)));
    layer3_outputs(875) <= not(layer2_outputs(1975)) or (layer2_outputs(970));
    layer3_outputs(876) <= not(layer2_outputs(1085));
    layer3_outputs(877) <= not(layer2_outputs(9791)) or (layer2_outputs(6451));
    layer3_outputs(878) <= not(layer2_outputs(1913));
    layer3_outputs(879) <= (layer2_outputs(3668)) or (layer2_outputs(7913));
    layer3_outputs(880) <= layer2_outputs(6436);
    layer3_outputs(881) <= layer2_outputs(69);
    layer3_outputs(882) <= not(layer2_outputs(1363));
    layer3_outputs(883) <= not(layer2_outputs(6543)) or (layer2_outputs(5961));
    layer3_outputs(884) <= layer2_outputs(3773);
    layer3_outputs(885) <= '0';
    layer3_outputs(886) <= '0';
    layer3_outputs(887) <= layer2_outputs(4725);
    layer3_outputs(888) <= layer2_outputs(6769);
    layer3_outputs(889) <= not((layer2_outputs(8375)) xor (layer2_outputs(5923)));
    layer3_outputs(890) <= not(layer2_outputs(7833));
    layer3_outputs(891) <= layer2_outputs(8086);
    layer3_outputs(892) <= (layer2_outputs(6391)) and (layer2_outputs(2275));
    layer3_outputs(893) <= (layer2_outputs(2303)) or (layer2_outputs(5906));
    layer3_outputs(894) <= not(layer2_outputs(117));
    layer3_outputs(895) <= not(layer2_outputs(5610)) or (layer2_outputs(10149));
    layer3_outputs(896) <= layer2_outputs(1839);
    layer3_outputs(897) <= (layer2_outputs(9006)) and not (layer2_outputs(3136));
    layer3_outputs(898) <= not(layer2_outputs(1681));
    layer3_outputs(899) <= (layer2_outputs(2807)) xor (layer2_outputs(1222));
    layer3_outputs(900) <= (layer2_outputs(8680)) or (layer2_outputs(3906));
    layer3_outputs(901) <= layer2_outputs(3698);
    layer3_outputs(902) <= (layer2_outputs(9109)) xor (layer2_outputs(4411));
    layer3_outputs(903) <= (layer2_outputs(2463)) and (layer2_outputs(8279));
    layer3_outputs(904) <= not((layer2_outputs(8678)) or (layer2_outputs(10155)));
    layer3_outputs(905) <= layer2_outputs(3154);
    layer3_outputs(906) <= (layer2_outputs(5781)) or (layer2_outputs(2296));
    layer3_outputs(907) <= not(layer2_outputs(8203)) or (layer2_outputs(2960));
    layer3_outputs(908) <= not(layer2_outputs(9758));
    layer3_outputs(909) <= layer2_outputs(2082);
    layer3_outputs(910) <= not(layer2_outputs(9676));
    layer3_outputs(911) <= not(layer2_outputs(2454)) or (layer2_outputs(4049));
    layer3_outputs(912) <= not(layer2_outputs(5009)) or (layer2_outputs(1614));
    layer3_outputs(913) <= (layer2_outputs(6827)) and (layer2_outputs(4319));
    layer3_outputs(914) <= not(layer2_outputs(10066));
    layer3_outputs(915) <= not((layer2_outputs(2229)) xor (layer2_outputs(5695)));
    layer3_outputs(916) <= (layer2_outputs(4841)) and not (layer2_outputs(8875));
    layer3_outputs(917) <= (layer2_outputs(9844)) or (layer2_outputs(3515));
    layer3_outputs(918) <= not((layer2_outputs(7685)) and (layer2_outputs(3072)));
    layer3_outputs(919) <= layer2_outputs(6051);
    layer3_outputs(920) <= (layer2_outputs(6978)) and (layer2_outputs(5260));
    layer3_outputs(921) <= (layer2_outputs(1198)) or (layer2_outputs(1958));
    layer3_outputs(922) <= not(layer2_outputs(10031));
    layer3_outputs(923) <= not(layer2_outputs(7062)) or (layer2_outputs(7222));
    layer3_outputs(924) <= not(layer2_outputs(2539));
    layer3_outputs(925) <= not((layer2_outputs(9075)) or (layer2_outputs(395)));
    layer3_outputs(926) <= layer2_outputs(8759);
    layer3_outputs(927) <= (layer2_outputs(8777)) xor (layer2_outputs(9393));
    layer3_outputs(928) <= layer2_outputs(7281);
    layer3_outputs(929) <= layer2_outputs(9771);
    layer3_outputs(930) <= not(layer2_outputs(5434)) or (layer2_outputs(2040));
    layer3_outputs(931) <= not(layer2_outputs(2668)) or (layer2_outputs(3636));
    layer3_outputs(932) <= not((layer2_outputs(4781)) and (layer2_outputs(1963)));
    layer3_outputs(933) <= (layer2_outputs(1784)) or (layer2_outputs(7534));
    layer3_outputs(934) <= (layer2_outputs(4971)) or (layer2_outputs(8755));
    layer3_outputs(935) <= not(layer2_outputs(1009)) or (layer2_outputs(8649));
    layer3_outputs(936) <= not(layer2_outputs(4813));
    layer3_outputs(937) <= not((layer2_outputs(5833)) or (layer2_outputs(390)));
    layer3_outputs(938) <= (layer2_outputs(8713)) and not (layer2_outputs(3512));
    layer3_outputs(939) <= not(layer2_outputs(3878));
    layer3_outputs(940) <= (layer2_outputs(1014)) and not (layer2_outputs(9394));
    layer3_outputs(941) <= layer2_outputs(4884);
    layer3_outputs(942) <= (layer2_outputs(5312)) and not (layer2_outputs(7962));
    layer3_outputs(943) <= not(layer2_outputs(8144));
    layer3_outputs(944) <= layer2_outputs(2010);
    layer3_outputs(945) <= not(layer2_outputs(8046));
    layer3_outputs(946) <= layer2_outputs(4037);
    layer3_outputs(947) <= (layer2_outputs(2350)) and not (layer2_outputs(4367));
    layer3_outputs(948) <= not(layer2_outputs(10078));
    layer3_outputs(949) <= layer2_outputs(456);
    layer3_outputs(950) <= not(layer2_outputs(7270)) or (layer2_outputs(4102));
    layer3_outputs(951) <= not(layer2_outputs(570));
    layer3_outputs(952) <= layer2_outputs(690);
    layer3_outputs(953) <= not(layer2_outputs(68));
    layer3_outputs(954) <= not((layer2_outputs(8299)) and (layer2_outputs(7654)));
    layer3_outputs(955) <= (layer2_outputs(9327)) and not (layer2_outputs(6841));
    layer3_outputs(956) <= layer2_outputs(9577);
    layer3_outputs(957) <= (layer2_outputs(2586)) or (layer2_outputs(3304));
    layer3_outputs(958) <= not(layer2_outputs(1761));
    layer3_outputs(959) <= layer2_outputs(7529);
    layer3_outputs(960) <= not(layer2_outputs(979));
    layer3_outputs(961) <= not(layer2_outputs(4846)) or (layer2_outputs(4296));
    layer3_outputs(962) <= not(layer2_outputs(4561));
    layer3_outputs(963) <= layer2_outputs(1654);
    layer3_outputs(964) <= layer2_outputs(6337);
    layer3_outputs(965) <= not(layer2_outputs(5155));
    layer3_outputs(966) <= layer2_outputs(8515);
    layer3_outputs(967) <= (layer2_outputs(309)) xor (layer2_outputs(9144));
    layer3_outputs(968) <= (layer2_outputs(8607)) xor (layer2_outputs(923));
    layer3_outputs(969) <= (layer2_outputs(9230)) xor (layer2_outputs(10165));
    layer3_outputs(970) <= not(layer2_outputs(5119)) or (layer2_outputs(5936));
    layer3_outputs(971) <= (layer2_outputs(4689)) xor (layer2_outputs(1103));
    layer3_outputs(972) <= (layer2_outputs(7709)) and (layer2_outputs(9703));
    layer3_outputs(973) <= layer2_outputs(1155);
    layer3_outputs(974) <= layer2_outputs(2949);
    layer3_outputs(975) <= layer2_outputs(4030);
    layer3_outputs(976) <= not(layer2_outputs(6946));
    layer3_outputs(977) <= layer2_outputs(9058);
    layer3_outputs(978) <= layer2_outputs(8648);
    layer3_outputs(979) <= layer2_outputs(8156);
    layer3_outputs(980) <= not((layer2_outputs(6177)) and (layer2_outputs(1459)));
    layer3_outputs(981) <= not(layer2_outputs(4865));
    layer3_outputs(982) <= (layer2_outputs(1375)) and not (layer2_outputs(565));
    layer3_outputs(983) <= layer2_outputs(3791);
    layer3_outputs(984) <= not(layer2_outputs(5475));
    layer3_outputs(985) <= not(layer2_outputs(2715));
    layer3_outputs(986) <= layer2_outputs(148);
    layer3_outputs(987) <= layer2_outputs(2034);
    layer3_outputs(988) <= (layer2_outputs(9573)) or (layer2_outputs(4180));
    layer3_outputs(989) <= not((layer2_outputs(9893)) xor (layer2_outputs(7406)));
    layer3_outputs(990) <= not(layer2_outputs(4094));
    layer3_outputs(991) <= not(layer2_outputs(3705));
    layer3_outputs(992) <= layer2_outputs(3124);
    layer3_outputs(993) <= (layer2_outputs(5046)) and (layer2_outputs(5390));
    layer3_outputs(994) <= not(layer2_outputs(9942)) or (layer2_outputs(1012));
    layer3_outputs(995) <= layer2_outputs(9476);
    layer3_outputs(996) <= not(layer2_outputs(280)) or (layer2_outputs(5038));
    layer3_outputs(997) <= not(layer2_outputs(6373));
    layer3_outputs(998) <= not(layer2_outputs(8135));
    layer3_outputs(999) <= not((layer2_outputs(8622)) xor (layer2_outputs(863)));
    layer3_outputs(1000) <= not(layer2_outputs(8542));
    layer3_outputs(1001) <= (layer2_outputs(2718)) and not (layer2_outputs(3075));
    layer3_outputs(1002) <= layer2_outputs(8023);
    layer3_outputs(1003) <= layer2_outputs(6074);
    layer3_outputs(1004) <= (layer2_outputs(2362)) and not (layer2_outputs(1364));
    layer3_outputs(1005) <= layer2_outputs(9358);
    layer3_outputs(1006) <= layer2_outputs(6977);
    layer3_outputs(1007) <= (layer2_outputs(1633)) or (layer2_outputs(9327));
    layer3_outputs(1008) <= (layer2_outputs(3091)) xor (layer2_outputs(3011));
    layer3_outputs(1009) <= (layer2_outputs(2941)) xor (layer2_outputs(8083));
    layer3_outputs(1010) <= layer2_outputs(9615);
    layer3_outputs(1011) <= layer2_outputs(9289);
    layer3_outputs(1012) <= not(layer2_outputs(6889));
    layer3_outputs(1013) <= layer2_outputs(9588);
    layer3_outputs(1014) <= not(layer2_outputs(4531));
    layer3_outputs(1015) <= (layer2_outputs(4548)) and not (layer2_outputs(8864));
    layer3_outputs(1016) <= (layer2_outputs(5707)) and not (layer2_outputs(1813));
    layer3_outputs(1017) <= (layer2_outputs(6851)) and not (layer2_outputs(8994));
    layer3_outputs(1018) <= not(layer2_outputs(6569)) or (layer2_outputs(1247));
    layer3_outputs(1019) <= layer2_outputs(6530);
    layer3_outputs(1020) <= not((layer2_outputs(5907)) and (layer2_outputs(10157)));
    layer3_outputs(1021) <= not(layer2_outputs(1001)) or (layer2_outputs(8903));
    layer3_outputs(1022) <= not(layer2_outputs(3114)) or (layer2_outputs(5947));
    layer3_outputs(1023) <= (layer2_outputs(3456)) and not (layer2_outputs(821));
    layer3_outputs(1024) <= not(layer2_outputs(1920));
    layer3_outputs(1025) <= layer2_outputs(2930);
    layer3_outputs(1026) <= layer2_outputs(2506);
    layer3_outputs(1027) <= (layer2_outputs(8394)) and not (layer2_outputs(7710));
    layer3_outputs(1028) <= (layer2_outputs(5903)) and not (layer2_outputs(6376));
    layer3_outputs(1029) <= (layer2_outputs(3261)) and not (layer2_outputs(9765));
    layer3_outputs(1030) <= (layer2_outputs(3177)) or (layer2_outputs(7358));
    layer3_outputs(1031) <= '0';
    layer3_outputs(1032) <= not(layer2_outputs(6941)) or (layer2_outputs(4936));
    layer3_outputs(1033) <= not(layer2_outputs(6507));
    layer3_outputs(1034) <= not(layer2_outputs(8102)) or (layer2_outputs(3170));
    layer3_outputs(1035) <= not(layer2_outputs(3550)) or (layer2_outputs(1947));
    layer3_outputs(1036) <= not((layer2_outputs(7794)) xor (layer2_outputs(5416)));
    layer3_outputs(1037) <= not(layer2_outputs(4270)) or (layer2_outputs(768));
    layer3_outputs(1038) <= layer2_outputs(7405);
    layer3_outputs(1039) <= (layer2_outputs(6599)) xor (layer2_outputs(8962));
    layer3_outputs(1040) <= (layer2_outputs(2609)) xor (layer2_outputs(6071));
    layer3_outputs(1041) <= layer2_outputs(1939);
    layer3_outputs(1042) <= layer2_outputs(8211);
    layer3_outputs(1043) <= (layer2_outputs(5536)) and not (layer2_outputs(7944));
    layer3_outputs(1044) <= layer2_outputs(6334);
    layer3_outputs(1045) <= not(layer2_outputs(4602)) or (layer2_outputs(6397));
    layer3_outputs(1046) <= not(layer2_outputs(1777));
    layer3_outputs(1047) <= layer2_outputs(1703);
    layer3_outputs(1048) <= not((layer2_outputs(9774)) xor (layer2_outputs(6985)));
    layer3_outputs(1049) <= layer2_outputs(393);
    layer3_outputs(1050) <= not(layer2_outputs(6169));
    layer3_outputs(1051) <= not(layer2_outputs(2589));
    layer3_outputs(1052) <= layer2_outputs(6880);
    layer3_outputs(1053) <= layer2_outputs(6899);
    layer3_outputs(1054) <= layer2_outputs(7237);
    layer3_outputs(1055) <= layer2_outputs(9351);
    layer3_outputs(1056) <= (layer2_outputs(241)) and not (layer2_outputs(1640));
    layer3_outputs(1057) <= not(layer2_outputs(1349));
    layer3_outputs(1058) <= not((layer2_outputs(9886)) and (layer2_outputs(2683)));
    layer3_outputs(1059) <= (layer2_outputs(4361)) xor (layer2_outputs(8430));
    layer3_outputs(1060) <= (layer2_outputs(9379)) and not (layer2_outputs(4801));
    layer3_outputs(1061) <= not((layer2_outputs(4774)) or (layer2_outputs(9394)));
    layer3_outputs(1062) <= (layer2_outputs(5023)) or (layer2_outputs(2470));
    layer3_outputs(1063) <= not(layer2_outputs(6317)) or (layer2_outputs(651));
    layer3_outputs(1064) <= not(layer2_outputs(10239));
    layer3_outputs(1065) <= not(layer2_outputs(8808));
    layer3_outputs(1066) <= (layer2_outputs(4346)) and (layer2_outputs(1121));
    layer3_outputs(1067) <= layer2_outputs(8068);
    layer3_outputs(1068) <= layer2_outputs(2048);
    layer3_outputs(1069) <= layer2_outputs(10122);
    layer3_outputs(1070) <= layer2_outputs(8109);
    layer3_outputs(1071) <= '1';
    layer3_outputs(1072) <= layer2_outputs(7973);
    layer3_outputs(1073) <= layer2_outputs(8298);
    layer3_outputs(1074) <= not(layer2_outputs(7401));
    layer3_outputs(1075) <= not(layer2_outputs(496));
    layer3_outputs(1076) <= not(layer2_outputs(4832)) or (layer2_outputs(9437));
    layer3_outputs(1077) <= (layer2_outputs(8952)) or (layer2_outputs(4655));
    layer3_outputs(1078) <= not(layer2_outputs(1613)) or (layer2_outputs(2643));
    layer3_outputs(1079) <= layer2_outputs(2117);
    layer3_outputs(1080) <= layer2_outputs(1027);
    layer3_outputs(1081) <= not(layer2_outputs(10082));
    layer3_outputs(1082) <= layer2_outputs(6169);
    layer3_outputs(1083) <= layer2_outputs(3705);
    layer3_outputs(1084) <= not(layer2_outputs(3626));
    layer3_outputs(1085) <= not(layer2_outputs(5733)) or (layer2_outputs(8985));
    layer3_outputs(1086) <= (layer2_outputs(6188)) or (layer2_outputs(5201));
    layer3_outputs(1087) <= layer2_outputs(6162);
    layer3_outputs(1088) <= not(layer2_outputs(7391));
    layer3_outputs(1089) <= not((layer2_outputs(3861)) or (layer2_outputs(6173)));
    layer3_outputs(1090) <= not(layer2_outputs(5682)) or (layer2_outputs(9133));
    layer3_outputs(1091) <= (layer2_outputs(507)) and not (layer2_outputs(8365));
    layer3_outputs(1092) <= layer2_outputs(331);
    layer3_outputs(1093) <= not((layer2_outputs(3761)) and (layer2_outputs(3721)));
    layer3_outputs(1094) <= not(layer2_outputs(2868));
    layer3_outputs(1095) <= layer2_outputs(7771);
    layer3_outputs(1096) <= layer2_outputs(1438);
    layer3_outputs(1097) <= not((layer2_outputs(47)) and (layer2_outputs(6814)));
    layer3_outputs(1098) <= (layer2_outputs(6393)) or (layer2_outputs(1759));
    layer3_outputs(1099) <= (layer2_outputs(2675)) and not (layer2_outputs(6860));
    layer3_outputs(1100) <= not((layer2_outputs(3377)) and (layer2_outputs(1494)));
    layer3_outputs(1101) <= (layer2_outputs(4616)) and not (layer2_outputs(2292));
    layer3_outputs(1102) <= not(layer2_outputs(105)) or (layer2_outputs(159));
    layer3_outputs(1103) <= (layer2_outputs(3224)) and not (layer2_outputs(612));
    layer3_outputs(1104) <= (layer2_outputs(4571)) or (layer2_outputs(6481));
    layer3_outputs(1105) <= (layer2_outputs(2900)) and (layer2_outputs(3215));
    layer3_outputs(1106) <= (layer2_outputs(7458)) or (layer2_outputs(3466));
    layer3_outputs(1107) <= layer2_outputs(2849);
    layer3_outputs(1108) <= not(layer2_outputs(9651));
    layer3_outputs(1109) <= not((layer2_outputs(7003)) and (layer2_outputs(5770)));
    layer3_outputs(1110) <= (layer2_outputs(8620)) or (layer2_outputs(871));
    layer3_outputs(1111) <= (layer2_outputs(3568)) xor (layer2_outputs(6077));
    layer3_outputs(1112) <= layer2_outputs(2962);
    layer3_outputs(1113) <= not((layer2_outputs(7182)) and (layer2_outputs(515)));
    layer3_outputs(1114) <= not((layer2_outputs(5516)) or (layer2_outputs(3440)));
    layer3_outputs(1115) <= layer2_outputs(5335);
    layer3_outputs(1116) <= layer2_outputs(4335);
    layer3_outputs(1117) <= (layer2_outputs(8743)) xor (layer2_outputs(6593));
    layer3_outputs(1118) <= '1';
    layer3_outputs(1119) <= not(layer2_outputs(3941));
    layer3_outputs(1120) <= (layer2_outputs(6597)) or (layer2_outputs(6299));
    layer3_outputs(1121) <= not(layer2_outputs(9449));
    layer3_outputs(1122) <= not(layer2_outputs(1294));
    layer3_outputs(1123) <= not(layer2_outputs(4263));
    layer3_outputs(1124) <= (layer2_outputs(8155)) and not (layer2_outputs(6714));
    layer3_outputs(1125) <= layer2_outputs(8317);
    layer3_outputs(1126) <= layer2_outputs(7209);
    layer3_outputs(1127) <= not(layer2_outputs(2207));
    layer3_outputs(1128) <= layer2_outputs(8754);
    layer3_outputs(1129) <= not(layer2_outputs(9568));
    layer3_outputs(1130) <= layer2_outputs(6782);
    layer3_outputs(1131) <= layer2_outputs(2);
    layer3_outputs(1132) <= layer2_outputs(4910);
    layer3_outputs(1133) <= not(layer2_outputs(2688));
    layer3_outputs(1134) <= layer2_outputs(8856);
    layer3_outputs(1135) <= layer2_outputs(1681);
    layer3_outputs(1136) <= (layer2_outputs(2950)) and not (layer2_outputs(606));
    layer3_outputs(1137) <= not(layer2_outputs(5129));
    layer3_outputs(1138) <= layer2_outputs(4696);
    layer3_outputs(1139) <= not(layer2_outputs(4643));
    layer3_outputs(1140) <= not(layer2_outputs(10020)) or (layer2_outputs(871));
    layer3_outputs(1141) <= (layer2_outputs(683)) xor (layer2_outputs(4066));
    layer3_outputs(1142) <= not(layer2_outputs(1290));
    layer3_outputs(1143) <= not(layer2_outputs(6356));
    layer3_outputs(1144) <= (layer2_outputs(6194)) and not (layer2_outputs(6882));
    layer3_outputs(1145) <= (layer2_outputs(5057)) xor (layer2_outputs(7075));
    layer3_outputs(1146) <= not((layer2_outputs(7587)) or (layer2_outputs(5975)));
    layer3_outputs(1147) <= layer2_outputs(7981);
    layer3_outputs(1148) <= not(layer2_outputs(1243)) or (layer2_outputs(1990));
    layer3_outputs(1149) <= (layer2_outputs(5680)) xor (layer2_outputs(1725));
    layer3_outputs(1150) <= not(layer2_outputs(1677)) or (layer2_outputs(3467));
    layer3_outputs(1151) <= not(layer2_outputs(504));
    layer3_outputs(1152) <= not(layer2_outputs(349)) or (layer2_outputs(954));
    layer3_outputs(1153) <= layer2_outputs(9297);
    layer3_outputs(1154) <= not(layer2_outputs(7133));
    layer3_outputs(1155) <= not(layer2_outputs(9456)) or (layer2_outputs(4670));
    layer3_outputs(1156) <= (layer2_outputs(4765)) or (layer2_outputs(5645));
    layer3_outputs(1157) <= not(layer2_outputs(3135)) or (layer2_outputs(9862));
    layer3_outputs(1158) <= (layer2_outputs(10183)) xor (layer2_outputs(1657));
    layer3_outputs(1159) <= not(layer2_outputs(1651)) or (layer2_outputs(4170));
    layer3_outputs(1160) <= not(layer2_outputs(9923));
    layer3_outputs(1161) <= layer2_outputs(8043);
    layer3_outputs(1162) <= (layer2_outputs(506)) or (layer2_outputs(1757));
    layer3_outputs(1163) <= (layer2_outputs(8674)) and not (layer2_outputs(10026));
    layer3_outputs(1164) <= layer2_outputs(4759);
    layer3_outputs(1165) <= (layer2_outputs(173)) and not (layer2_outputs(7908));
    layer3_outputs(1166) <= not(layer2_outputs(3227));
    layer3_outputs(1167) <= (layer2_outputs(5874)) xor (layer2_outputs(258));
    layer3_outputs(1168) <= not((layer2_outputs(688)) and (layer2_outputs(9153)));
    layer3_outputs(1169) <= (layer2_outputs(7587)) and (layer2_outputs(9856));
    layer3_outputs(1170) <= (layer2_outputs(3234)) and not (layer2_outputs(5700));
    layer3_outputs(1171) <= not(layer2_outputs(4691)) or (layer2_outputs(1699));
    layer3_outputs(1172) <= not(layer2_outputs(9579)) or (layer2_outputs(6564));
    layer3_outputs(1173) <= not(layer2_outputs(9092));
    layer3_outputs(1174) <= layer2_outputs(4567);
    layer3_outputs(1175) <= (layer2_outputs(8968)) xor (layer2_outputs(2834));
    layer3_outputs(1176) <= (layer2_outputs(593)) and (layer2_outputs(3317));
    layer3_outputs(1177) <= not(layer2_outputs(5957)) or (layer2_outputs(10094));
    layer3_outputs(1178) <= (layer2_outputs(6651)) and not (layer2_outputs(1216));
    layer3_outputs(1179) <= not((layer2_outputs(2336)) xor (layer2_outputs(9204)));
    layer3_outputs(1180) <= layer2_outputs(4724);
    layer3_outputs(1181) <= layer2_outputs(8456);
    layer3_outputs(1182) <= (layer2_outputs(3606)) and not (layer2_outputs(2992));
    layer3_outputs(1183) <= not(layer2_outputs(1054));
    layer3_outputs(1184) <= '0';
    layer3_outputs(1185) <= (layer2_outputs(6797)) xor (layer2_outputs(8701));
    layer3_outputs(1186) <= not(layer2_outputs(358));
    layer3_outputs(1187) <= layer2_outputs(4570);
    layer3_outputs(1188) <= not(layer2_outputs(3942));
    layer3_outputs(1189) <= layer2_outputs(9283);
    layer3_outputs(1190) <= not(layer2_outputs(4046));
    layer3_outputs(1191) <= layer2_outputs(2129);
    layer3_outputs(1192) <= '1';
    layer3_outputs(1193) <= not(layer2_outputs(8339));
    layer3_outputs(1194) <= layer2_outputs(3051);
    layer3_outputs(1195) <= not(layer2_outputs(3355)) or (layer2_outputs(4800));
    layer3_outputs(1196) <= (layer2_outputs(6991)) xor (layer2_outputs(5420));
    layer3_outputs(1197) <= not(layer2_outputs(6113)) or (layer2_outputs(2098));
    layer3_outputs(1198) <= not((layer2_outputs(9376)) and (layer2_outputs(5578)));
    layer3_outputs(1199) <= layer2_outputs(254);
    layer3_outputs(1200) <= not(layer2_outputs(10100)) or (layer2_outputs(9624));
    layer3_outputs(1201) <= not(layer2_outputs(6951)) or (layer2_outputs(7672));
    layer3_outputs(1202) <= not(layer2_outputs(7616)) or (layer2_outputs(7724));
    layer3_outputs(1203) <= (layer2_outputs(8011)) and not (layer2_outputs(3800));
    layer3_outputs(1204) <= not(layer2_outputs(4631));
    layer3_outputs(1205) <= (layer2_outputs(2640)) and not (layer2_outputs(5659));
    layer3_outputs(1206) <= not(layer2_outputs(7699)) or (layer2_outputs(9841));
    layer3_outputs(1207) <= not((layer2_outputs(590)) xor (layer2_outputs(260)));
    layer3_outputs(1208) <= not(layer2_outputs(7374));
    layer3_outputs(1209) <= (layer2_outputs(8242)) or (layer2_outputs(1055));
    layer3_outputs(1210) <= layer2_outputs(4004);
    layer3_outputs(1211) <= not(layer2_outputs(7510)) or (layer2_outputs(1593));
    layer3_outputs(1212) <= (layer2_outputs(327)) and not (layer2_outputs(9706));
    layer3_outputs(1213) <= layer2_outputs(2939);
    layer3_outputs(1214) <= layer2_outputs(732);
    layer3_outputs(1215) <= (layer2_outputs(1033)) xor (layer2_outputs(3763));
    layer3_outputs(1216) <= (layer2_outputs(8468)) xor (layer2_outputs(3666));
    layer3_outputs(1217) <= not(layer2_outputs(8262));
    layer3_outputs(1218) <= not(layer2_outputs(2586));
    layer3_outputs(1219) <= not(layer2_outputs(2180)) or (layer2_outputs(1463));
    layer3_outputs(1220) <= not(layer2_outputs(76));
    layer3_outputs(1221) <= layer2_outputs(8514);
    layer3_outputs(1222) <= layer2_outputs(6042);
    layer3_outputs(1223) <= (layer2_outputs(6739)) and (layer2_outputs(3881));
    layer3_outputs(1224) <= not(layer2_outputs(7027));
    layer3_outputs(1225) <= not(layer2_outputs(8464)) or (layer2_outputs(2655));
    layer3_outputs(1226) <= not(layer2_outputs(834));
    layer3_outputs(1227) <= layer2_outputs(6911);
    layer3_outputs(1228) <= not(layer2_outputs(7062));
    layer3_outputs(1229) <= (layer2_outputs(2412)) and not (layer2_outputs(6413));
    layer3_outputs(1230) <= (layer2_outputs(3191)) and (layer2_outputs(2359));
    layer3_outputs(1231) <= not((layer2_outputs(4749)) or (layer2_outputs(9595)));
    layer3_outputs(1232) <= layer2_outputs(9848);
    layer3_outputs(1233) <= not((layer2_outputs(9882)) and (layer2_outputs(9258)));
    layer3_outputs(1234) <= layer2_outputs(10173);
    layer3_outputs(1235) <= not(layer2_outputs(6995)) or (layer2_outputs(5494));
    layer3_outputs(1236) <= not(layer2_outputs(1684));
    layer3_outputs(1237) <= (layer2_outputs(333)) and (layer2_outputs(3543));
    layer3_outputs(1238) <= layer2_outputs(1185);
    layer3_outputs(1239) <= layer2_outputs(5916);
    layer3_outputs(1240) <= (layer2_outputs(4856)) and (layer2_outputs(4591));
    layer3_outputs(1241) <= layer2_outputs(1425);
    layer3_outputs(1242) <= not(layer2_outputs(9860));
    layer3_outputs(1243) <= layer2_outputs(8670);
    layer3_outputs(1244) <= not(layer2_outputs(4840));
    layer3_outputs(1245) <= (layer2_outputs(6359)) and not (layer2_outputs(9368));
    layer3_outputs(1246) <= (layer2_outputs(317)) and not (layer2_outputs(1744));
    layer3_outputs(1247) <= not((layer2_outputs(7086)) and (layer2_outputs(10179)));
    layer3_outputs(1248) <= not(layer2_outputs(8073)) or (layer2_outputs(8897));
    layer3_outputs(1249) <= not((layer2_outputs(3039)) or (layer2_outputs(9797)));
    layer3_outputs(1250) <= not(layer2_outputs(8820));
    layer3_outputs(1251) <= (layer2_outputs(2357)) and not (layer2_outputs(2993));
    layer3_outputs(1252) <= not(layer2_outputs(4244)) or (layer2_outputs(4943));
    layer3_outputs(1253) <= layer2_outputs(5225);
    layer3_outputs(1254) <= (layer2_outputs(374)) or (layer2_outputs(306));
    layer3_outputs(1255) <= (layer2_outputs(1232)) or (layer2_outputs(7252));
    layer3_outputs(1256) <= not(layer2_outputs(7664));
    layer3_outputs(1257) <= layer2_outputs(7913);
    layer3_outputs(1258) <= not(layer2_outputs(294));
    layer3_outputs(1259) <= layer2_outputs(9247);
    layer3_outputs(1260) <= (layer2_outputs(7842)) xor (layer2_outputs(5195));
    layer3_outputs(1261) <= not(layer2_outputs(8973));
    layer3_outputs(1262) <= not(layer2_outputs(7097));
    layer3_outputs(1263) <= layer2_outputs(1300);
    layer3_outputs(1264) <= layer2_outputs(6127);
    layer3_outputs(1265) <= not(layer2_outputs(1796)) or (layer2_outputs(7629));
    layer3_outputs(1266) <= not(layer2_outputs(2381)) or (layer2_outputs(2733));
    layer3_outputs(1267) <= not(layer2_outputs(4038));
    layer3_outputs(1268) <= (layer2_outputs(8439)) and not (layer2_outputs(3579));
    layer3_outputs(1269) <= not(layer2_outputs(604)) or (layer2_outputs(3843));
    layer3_outputs(1270) <= (layer2_outputs(6373)) and (layer2_outputs(8241));
    layer3_outputs(1271) <= not(layer2_outputs(711)) or (layer2_outputs(3360));
    layer3_outputs(1272) <= (layer2_outputs(4231)) and not (layer2_outputs(7011));
    layer3_outputs(1273) <= (layer2_outputs(2027)) and (layer2_outputs(4537));
    layer3_outputs(1274) <= layer2_outputs(4202);
    layer3_outputs(1275) <= layer2_outputs(913);
    layer3_outputs(1276) <= layer2_outputs(4375);
    layer3_outputs(1277) <= layer2_outputs(6264);
    layer3_outputs(1278) <= not(layer2_outputs(9574));
    layer3_outputs(1279) <= (layer2_outputs(8214)) or (layer2_outputs(9438));
    layer3_outputs(1280) <= not((layer2_outputs(6002)) xor (layer2_outputs(693)));
    layer3_outputs(1281) <= layer2_outputs(5456);
    layer3_outputs(1282) <= (layer2_outputs(9669)) or (layer2_outputs(625));
    layer3_outputs(1283) <= not(layer2_outputs(1072));
    layer3_outputs(1284) <= not(layer2_outputs(1105));
    layer3_outputs(1285) <= layer2_outputs(2007);
    layer3_outputs(1286) <= (layer2_outputs(9178)) or (layer2_outputs(6082));
    layer3_outputs(1287) <= (layer2_outputs(3789)) and not (layer2_outputs(10152));
    layer3_outputs(1288) <= (layer2_outputs(5121)) and (layer2_outputs(6667));
    layer3_outputs(1289) <= '0';
    layer3_outputs(1290) <= not(layer2_outputs(7428)) or (layer2_outputs(1950));
    layer3_outputs(1291) <= (layer2_outputs(5711)) and not (layer2_outputs(6631));
    layer3_outputs(1292) <= layer2_outputs(8910);
    layer3_outputs(1293) <= not(layer2_outputs(4016));
    layer3_outputs(1294) <= (layer2_outputs(9814)) xor (layer2_outputs(2083));
    layer3_outputs(1295) <= layer2_outputs(4557);
    layer3_outputs(1296) <= layer2_outputs(3802);
    layer3_outputs(1297) <= not(layer2_outputs(375));
    layer3_outputs(1298) <= not(layer2_outputs(8218));
    layer3_outputs(1299) <= not((layer2_outputs(3404)) and (layer2_outputs(8798)));
    layer3_outputs(1300) <= layer2_outputs(4079);
    layer3_outputs(1301) <= not(layer2_outputs(9816));
    layer3_outputs(1302) <= layer2_outputs(8340);
    layer3_outputs(1303) <= (layer2_outputs(4618)) xor (layer2_outputs(971));
    layer3_outputs(1304) <= not((layer2_outputs(9468)) or (layer2_outputs(6240)));
    layer3_outputs(1305) <= (layer2_outputs(6463)) or (layer2_outputs(7409));
    layer3_outputs(1306) <= (layer2_outputs(1084)) and not (layer2_outputs(2895));
    layer3_outputs(1307) <= not(layer2_outputs(6019));
    layer3_outputs(1308) <= not((layer2_outputs(4050)) or (layer2_outputs(1799)));
    layer3_outputs(1309) <= layer2_outputs(2045);
    layer3_outputs(1310) <= not(layer2_outputs(4905));
    layer3_outputs(1311) <= (layer2_outputs(4344)) xor (layer2_outputs(9628));
    layer3_outputs(1312) <= not(layer2_outputs(9288)) or (layer2_outputs(6655));
    layer3_outputs(1313) <= not(layer2_outputs(6639));
    layer3_outputs(1314) <= (layer2_outputs(7630)) and not (layer2_outputs(9650));
    layer3_outputs(1315) <= (layer2_outputs(3993)) and (layer2_outputs(2108));
    layer3_outputs(1316) <= not(layer2_outputs(317));
    layer3_outputs(1317) <= (layer2_outputs(2841)) and not (layer2_outputs(8712));
    layer3_outputs(1318) <= layer2_outputs(5224);
    layer3_outputs(1319) <= (layer2_outputs(4522)) and (layer2_outputs(10084));
    layer3_outputs(1320) <= not(layer2_outputs(7426));
    layer3_outputs(1321) <= not((layer2_outputs(5311)) xor (layer2_outputs(10013)));
    layer3_outputs(1322) <= layer2_outputs(8114);
    layer3_outputs(1323) <= (layer2_outputs(2149)) and (layer2_outputs(6702));
    layer3_outputs(1324) <= not((layer2_outputs(7219)) and (layer2_outputs(9381)));
    layer3_outputs(1325) <= (layer2_outputs(4413)) and (layer2_outputs(4249));
    layer3_outputs(1326) <= not(layer2_outputs(5582));
    layer3_outputs(1327) <= '1';
    layer3_outputs(1328) <= not(layer2_outputs(713)) or (layer2_outputs(7040));
    layer3_outputs(1329) <= not((layer2_outputs(10058)) and (layer2_outputs(4281)));
    layer3_outputs(1330) <= not(layer2_outputs(7390));
    layer3_outputs(1331) <= not(layer2_outputs(5060));
    layer3_outputs(1332) <= not(layer2_outputs(7199));
    layer3_outputs(1333) <= not(layer2_outputs(217));
    layer3_outputs(1334) <= '1';
    layer3_outputs(1335) <= not(layer2_outputs(10000));
    layer3_outputs(1336) <= (layer2_outputs(7633)) or (layer2_outputs(3554));
    layer3_outputs(1337) <= not(layer2_outputs(9180));
    layer3_outputs(1338) <= layer2_outputs(2150);
    layer3_outputs(1339) <= not((layer2_outputs(7818)) or (layer2_outputs(8223)));
    layer3_outputs(1340) <= (layer2_outputs(1835)) and not (layer2_outputs(6684));
    layer3_outputs(1341) <= layer2_outputs(7613);
    layer3_outputs(1342) <= layer2_outputs(1464);
    layer3_outputs(1343) <= not((layer2_outputs(6780)) xor (layer2_outputs(8318)));
    layer3_outputs(1344) <= (layer2_outputs(4711)) or (layer2_outputs(2177));
    layer3_outputs(1345) <= layer2_outputs(10113);
    layer3_outputs(1346) <= (layer2_outputs(1688)) and (layer2_outputs(6946));
    layer3_outputs(1347) <= not((layer2_outputs(2286)) xor (layer2_outputs(3535)));
    layer3_outputs(1348) <= not(layer2_outputs(2455));
    layer3_outputs(1349) <= not(layer2_outputs(9739));
    layer3_outputs(1350) <= not(layer2_outputs(10135));
    layer3_outputs(1351) <= not((layer2_outputs(8265)) xor (layer2_outputs(9779)));
    layer3_outputs(1352) <= not(layer2_outputs(1071));
    layer3_outputs(1353) <= (layer2_outputs(5725)) and not (layer2_outputs(3163));
    layer3_outputs(1354) <= not(layer2_outputs(9807));
    layer3_outputs(1355) <= layer2_outputs(4869);
    layer3_outputs(1356) <= not((layer2_outputs(4131)) or (layer2_outputs(9778)));
    layer3_outputs(1357) <= layer2_outputs(9904);
    layer3_outputs(1358) <= not(layer2_outputs(9607)) or (layer2_outputs(537));
    layer3_outputs(1359) <= (layer2_outputs(9273)) and (layer2_outputs(8969));
    layer3_outputs(1360) <= (layer2_outputs(5897)) and not (layer2_outputs(4314));
    layer3_outputs(1361) <= (layer2_outputs(6546)) and not (layer2_outputs(9160));
    layer3_outputs(1362) <= not(layer2_outputs(2120)) or (layer2_outputs(3672));
    layer3_outputs(1363) <= (layer2_outputs(2596)) and (layer2_outputs(6063));
    layer3_outputs(1364) <= not(layer2_outputs(5758));
    layer3_outputs(1365) <= not(layer2_outputs(5323));
    layer3_outputs(1366) <= (layer2_outputs(7139)) xor (layer2_outputs(5241));
    layer3_outputs(1367) <= not(layer2_outputs(1618));
    layer3_outputs(1368) <= layer2_outputs(3834);
    layer3_outputs(1369) <= not(layer2_outputs(5731));
    layer3_outputs(1370) <= (layer2_outputs(2783)) or (layer2_outputs(4426));
    layer3_outputs(1371) <= not(layer2_outputs(6630));
    layer3_outputs(1372) <= layer2_outputs(3640);
    layer3_outputs(1373) <= not((layer2_outputs(6715)) xor (layer2_outputs(9569)));
    layer3_outputs(1374) <= layer2_outputs(1940);
    layer3_outputs(1375) <= not(layer2_outputs(2542)) or (layer2_outputs(2620));
    layer3_outputs(1376) <= not(layer2_outputs(6921));
    layer3_outputs(1377) <= layer2_outputs(400);
    layer3_outputs(1378) <= (layer2_outputs(9601)) and (layer2_outputs(8312));
    layer3_outputs(1379) <= not(layer2_outputs(452)) or (layer2_outputs(7106));
    layer3_outputs(1380) <= not((layer2_outputs(4111)) or (layer2_outputs(7770)));
    layer3_outputs(1381) <= layer2_outputs(2402);
    layer3_outputs(1382) <= '0';
    layer3_outputs(1383) <= not((layer2_outputs(3051)) and (layer2_outputs(2072)));
    layer3_outputs(1384) <= (layer2_outputs(834)) and not (layer2_outputs(5706));
    layer3_outputs(1385) <= not(layer2_outputs(6527)) or (layer2_outputs(1709));
    layer3_outputs(1386) <= not(layer2_outputs(6631));
    layer3_outputs(1387) <= layer2_outputs(1521);
    layer3_outputs(1388) <= layer2_outputs(2623);
    layer3_outputs(1389) <= (layer2_outputs(9598)) and not (layer2_outputs(855));
    layer3_outputs(1390) <= (layer2_outputs(7708)) and not (layer2_outputs(1903));
    layer3_outputs(1391) <= layer2_outputs(3549);
    layer3_outputs(1392) <= layer2_outputs(3764);
    layer3_outputs(1393) <= not(layer2_outputs(867));
    layer3_outputs(1394) <= layer2_outputs(3293);
    layer3_outputs(1395) <= not(layer2_outputs(9374));
    layer3_outputs(1396) <= (layer2_outputs(4607)) and (layer2_outputs(7353));
    layer3_outputs(1397) <= not(layer2_outputs(5845));
    layer3_outputs(1398) <= not(layer2_outputs(1894));
    layer3_outputs(1399) <= layer2_outputs(5128);
    layer3_outputs(1400) <= (layer2_outputs(1531)) and not (layer2_outputs(10229));
    layer3_outputs(1401) <= layer2_outputs(9461);
    layer3_outputs(1402) <= not(layer2_outputs(8336));
    layer3_outputs(1403) <= not(layer2_outputs(9818)) or (layer2_outputs(7052));
    layer3_outputs(1404) <= (layer2_outputs(5875)) xor (layer2_outputs(3865));
    layer3_outputs(1405) <= not((layer2_outputs(3249)) and (layer2_outputs(8723)));
    layer3_outputs(1406) <= not((layer2_outputs(7459)) and (layer2_outputs(7368)));
    layer3_outputs(1407) <= not(layer2_outputs(8343));
    layer3_outputs(1408) <= (layer2_outputs(5369)) and (layer2_outputs(2895));
    layer3_outputs(1409) <= not((layer2_outputs(4135)) xor (layer2_outputs(124)));
    layer3_outputs(1410) <= not((layer2_outputs(8675)) or (layer2_outputs(152)));
    layer3_outputs(1411) <= (layer2_outputs(7671)) xor (layer2_outputs(4384));
    layer3_outputs(1412) <= not(layer2_outputs(8856));
    layer3_outputs(1413) <= not(layer2_outputs(4706));
    layer3_outputs(1414) <= (layer2_outputs(6509)) and not (layer2_outputs(956));
    layer3_outputs(1415) <= not(layer2_outputs(7697));
    layer3_outputs(1416) <= (layer2_outputs(3305)) and not (layer2_outputs(6703));
    layer3_outputs(1417) <= layer2_outputs(9238);
    layer3_outputs(1418) <= layer2_outputs(6165);
    layer3_outputs(1419) <= layer2_outputs(1240);
    layer3_outputs(1420) <= not(layer2_outputs(1790));
    layer3_outputs(1421) <= not(layer2_outputs(6830));
    layer3_outputs(1422) <= not(layer2_outputs(4448)) or (layer2_outputs(7935));
    layer3_outputs(1423) <= (layer2_outputs(3925)) and (layer2_outputs(9335));
    layer3_outputs(1424) <= not(layer2_outputs(4861));
    layer3_outputs(1425) <= not((layer2_outputs(9097)) and (layer2_outputs(9715)));
    layer3_outputs(1426) <= layer2_outputs(3258);
    layer3_outputs(1427) <= layer2_outputs(131);
    layer3_outputs(1428) <= layer2_outputs(9276);
    layer3_outputs(1429) <= (layer2_outputs(669)) xor (layer2_outputs(5316));
    layer3_outputs(1430) <= not(layer2_outputs(814));
    layer3_outputs(1431) <= not(layer2_outputs(5909));
    layer3_outputs(1432) <= not(layer2_outputs(7585));
    layer3_outputs(1433) <= '1';
    layer3_outputs(1434) <= not((layer2_outputs(2629)) xor (layer2_outputs(3359)));
    layer3_outputs(1435) <= not(layer2_outputs(6766));
    layer3_outputs(1436) <= not((layer2_outputs(7345)) xor (layer2_outputs(709)));
    layer3_outputs(1437) <= '0';
    layer3_outputs(1438) <= (layer2_outputs(5913)) or (layer2_outputs(4954));
    layer3_outputs(1439) <= not(layer2_outputs(9295)) or (layer2_outputs(4642));
    layer3_outputs(1440) <= (layer2_outputs(5867)) and not (layer2_outputs(7282));
    layer3_outputs(1441) <= layer2_outputs(1571);
    layer3_outputs(1442) <= (layer2_outputs(981)) and (layer2_outputs(7984));
    layer3_outputs(1443) <= not(layer2_outputs(4397));
    layer3_outputs(1444) <= layer2_outputs(1758);
    layer3_outputs(1445) <= not(layer2_outputs(328));
    layer3_outputs(1446) <= layer2_outputs(9712);
    layer3_outputs(1447) <= not(layer2_outputs(4734));
    layer3_outputs(1448) <= not(layer2_outputs(1107));
    layer3_outputs(1449) <= layer2_outputs(5313);
    layer3_outputs(1450) <= layer2_outputs(3177);
    layer3_outputs(1451) <= layer2_outputs(7908);
    layer3_outputs(1452) <= not(layer2_outputs(7976));
    layer3_outputs(1453) <= not(layer2_outputs(3764));
    layer3_outputs(1454) <= not(layer2_outputs(6191));
    layer3_outputs(1455) <= layer2_outputs(1454);
    layer3_outputs(1456) <= not((layer2_outputs(9485)) or (layer2_outputs(1146)));
    layer3_outputs(1457) <= (layer2_outputs(549)) and not (layer2_outputs(2213));
    layer3_outputs(1458) <= not(layer2_outputs(421));
    layer3_outputs(1459) <= not(layer2_outputs(2208));
    layer3_outputs(1460) <= layer2_outputs(4509);
    layer3_outputs(1461) <= not(layer2_outputs(711));
    layer3_outputs(1462) <= not(layer2_outputs(7528));
    layer3_outputs(1463) <= layer2_outputs(9882);
    layer3_outputs(1464) <= '1';
    layer3_outputs(1465) <= not(layer2_outputs(3860));
    layer3_outputs(1466) <= '0';
    layer3_outputs(1467) <= not(layer2_outputs(8523));
    layer3_outputs(1468) <= layer2_outputs(4268);
    layer3_outputs(1469) <= not(layer2_outputs(9)) or (layer2_outputs(4518));
    layer3_outputs(1470) <= layer2_outputs(2264);
    layer3_outputs(1471) <= not(layer2_outputs(1002));
    layer3_outputs(1472) <= (layer2_outputs(6963)) and not (layer2_outputs(3823));
    layer3_outputs(1473) <= '0';
    layer3_outputs(1474) <= layer2_outputs(6812);
    layer3_outputs(1475) <= not((layer2_outputs(3313)) or (layer2_outputs(6586)));
    layer3_outputs(1476) <= not(layer2_outputs(2826)) or (layer2_outputs(5547));
    layer3_outputs(1477) <= layer2_outputs(2415);
    layer3_outputs(1478) <= not(layer2_outputs(9086)) or (layer2_outputs(1489));
    layer3_outputs(1479) <= not(layer2_outputs(9801));
    layer3_outputs(1480) <= (layer2_outputs(7427)) or (layer2_outputs(8243));
    layer3_outputs(1481) <= layer2_outputs(1976);
    layer3_outputs(1482) <= not(layer2_outputs(3145));
    layer3_outputs(1483) <= not(layer2_outputs(1100)) or (layer2_outputs(1523));
    layer3_outputs(1484) <= not(layer2_outputs(8707)) or (layer2_outputs(7112));
    layer3_outputs(1485) <= not((layer2_outputs(1129)) or (layer2_outputs(8655)));
    layer3_outputs(1486) <= (layer2_outputs(3933)) or (layer2_outputs(9891));
    layer3_outputs(1487) <= layer2_outputs(9128);
    layer3_outputs(1488) <= (layer2_outputs(6181)) and not (layer2_outputs(5534));
    layer3_outputs(1489) <= not((layer2_outputs(10070)) or (layer2_outputs(5739)));
    layer3_outputs(1490) <= (layer2_outputs(4764)) xor (layer2_outputs(8099));
    layer3_outputs(1491) <= not(layer2_outputs(4948)) or (layer2_outputs(1754));
    layer3_outputs(1492) <= (layer2_outputs(9354)) and not (layer2_outputs(9864));
    layer3_outputs(1493) <= (layer2_outputs(625)) xor (layer2_outputs(3904));
    layer3_outputs(1494) <= (layer2_outputs(9622)) xor (layer2_outputs(9656));
    layer3_outputs(1495) <= (layer2_outputs(4350)) and (layer2_outputs(496));
    layer3_outputs(1496) <= (layer2_outputs(9658)) xor (layer2_outputs(6295));
    layer3_outputs(1497) <= layer2_outputs(6733);
    layer3_outputs(1498) <= layer2_outputs(7832);
    layer3_outputs(1499) <= (layer2_outputs(578)) and not (layer2_outputs(4876));
    layer3_outputs(1500) <= not(layer2_outputs(1139));
    layer3_outputs(1501) <= not(layer2_outputs(8497));
    layer3_outputs(1502) <= (layer2_outputs(850)) and not (layer2_outputs(6356));
    layer3_outputs(1503) <= '0';
    layer3_outputs(1504) <= not(layer2_outputs(7167)) or (layer2_outputs(3453));
    layer3_outputs(1505) <= '0';
    layer3_outputs(1506) <= not(layer2_outputs(450)) or (layer2_outputs(9708));
    layer3_outputs(1507) <= not(layer2_outputs(6026));
    layer3_outputs(1508) <= layer2_outputs(254);
    layer3_outputs(1509) <= (layer2_outputs(499)) xor (layer2_outputs(6087));
    layer3_outputs(1510) <= not(layer2_outputs(4545));
    layer3_outputs(1511) <= layer2_outputs(9564);
    layer3_outputs(1512) <= layer2_outputs(2356);
    layer3_outputs(1513) <= layer2_outputs(5430);
    layer3_outputs(1514) <= not((layer2_outputs(5061)) and (layer2_outputs(9264)));
    layer3_outputs(1515) <= not((layer2_outputs(653)) xor (layer2_outputs(2261)));
    layer3_outputs(1516) <= (layer2_outputs(535)) or (layer2_outputs(2274));
    layer3_outputs(1517) <= not(layer2_outputs(8103)) or (layer2_outputs(3639));
    layer3_outputs(1518) <= not(layer2_outputs(5595));
    layer3_outputs(1519) <= layer2_outputs(7826);
    layer3_outputs(1520) <= not(layer2_outputs(6121));
    layer3_outputs(1521) <= layer2_outputs(7885);
    layer3_outputs(1522) <= not((layer2_outputs(9111)) xor (layer2_outputs(1964)));
    layer3_outputs(1523) <= layer2_outputs(1704);
    layer3_outputs(1524) <= layer2_outputs(1306);
    layer3_outputs(1525) <= not(layer2_outputs(8565)) or (layer2_outputs(2887));
    layer3_outputs(1526) <= not((layer2_outputs(6571)) and (layer2_outputs(740)));
    layer3_outputs(1527) <= not((layer2_outputs(5750)) xor (layer2_outputs(5832)));
    layer3_outputs(1528) <= not(layer2_outputs(3406));
    layer3_outputs(1529) <= (layer2_outputs(9601)) xor (layer2_outputs(6107));
    layer3_outputs(1530) <= not(layer2_outputs(2351));
    layer3_outputs(1531) <= not(layer2_outputs(4983));
    layer3_outputs(1532) <= layer2_outputs(6994);
    layer3_outputs(1533) <= (layer2_outputs(5952)) or (layer2_outputs(4572));
    layer3_outputs(1534) <= (layer2_outputs(1697)) or (layer2_outputs(1043));
    layer3_outputs(1535) <= not(layer2_outputs(364));
    layer3_outputs(1536) <= not(layer2_outputs(6875));
    layer3_outputs(1537) <= layer2_outputs(708);
    layer3_outputs(1538) <= not(layer2_outputs(2501));
    layer3_outputs(1539) <= not((layer2_outputs(4712)) or (layer2_outputs(9664)));
    layer3_outputs(1540) <= not((layer2_outputs(6130)) and (layer2_outputs(1073)));
    layer3_outputs(1541) <= layer2_outputs(5130);
    layer3_outputs(1542) <= not(layer2_outputs(3100));
    layer3_outputs(1543) <= layer2_outputs(2393);
    layer3_outputs(1544) <= not(layer2_outputs(1685));
    layer3_outputs(1545) <= not(layer2_outputs(7230));
    layer3_outputs(1546) <= layer2_outputs(2096);
    layer3_outputs(1547) <= not(layer2_outputs(5046));
    layer3_outputs(1548) <= not(layer2_outputs(542)) or (layer2_outputs(6498));
    layer3_outputs(1549) <= not(layer2_outputs(1747)) or (layer2_outputs(7276));
    layer3_outputs(1550) <= not((layer2_outputs(1050)) or (layer2_outputs(1204)));
    layer3_outputs(1551) <= not(layer2_outputs(5103));
    layer3_outputs(1552) <= layer2_outputs(161);
    layer3_outputs(1553) <= layer2_outputs(3636);
    layer3_outputs(1554) <= (layer2_outputs(10055)) and (layer2_outputs(4291));
    layer3_outputs(1555) <= (layer2_outputs(6177)) xor (layer2_outputs(6770));
    layer3_outputs(1556) <= (layer2_outputs(2866)) and (layer2_outputs(1642));
    layer3_outputs(1557) <= layer2_outputs(9782);
    layer3_outputs(1558) <= layer2_outputs(7744);
    layer3_outputs(1559) <= layer2_outputs(3970);
    layer3_outputs(1560) <= not(layer2_outputs(3605));
    layer3_outputs(1561) <= (layer2_outputs(6431)) and not (layer2_outputs(6500));
    layer3_outputs(1562) <= not((layer2_outputs(7187)) xor (layer2_outputs(10000)));
    layer3_outputs(1563) <= not(layer2_outputs(7252));
    layer3_outputs(1564) <= '0';
    layer3_outputs(1565) <= '1';
    layer3_outputs(1566) <= not(layer2_outputs(8365));
    layer3_outputs(1567) <= not((layer2_outputs(1770)) and (layer2_outputs(8252)));
    layer3_outputs(1568) <= not(layer2_outputs(3426));
    layer3_outputs(1569) <= not(layer2_outputs(3138));
    layer3_outputs(1570) <= (layer2_outputs(5864)) xor (layer2_outputs(2251));
    layer3_outputs(1571) <= not(layer2_outputs(819));
    layer3_outputs(1572) <= layer2_outputs(120);
    layer3_outputs(1573) <= '1';
    layer3_outputs(1574) <= (layer2_outputs(2325)) xor (layer2_outputs(7519));
    layer3_outputs(1575) <= (layer2_outputs(7796)) or (layer2_outputs(4589));
    layer3_outputs(1576) <= not((layer2_outputs(5350)) or (layer2_outputs(508)));
    layer3_outputs(1577) <= (layer2_outputs(1382)) and not (layer2_outputs(3999));
    layer3_outputs(1578) <= not(layer2_outputs(6306));
    layer3_outputs(1579) <= (layer2_outputs(6566)) or (layer2_outputs(3491));
    layer3_outputs(1580) <= layer2_outputs(3062);
    layer3_outputs(1581) <= not(layer2_outputs(3300));
    layer3_outputs(1582) <= (layer2_outputs(4710)) xor (layer2_outputs(7686));
    layer3_outputs(1583) <= not((layer2_outputs(5456)) xor (layer2_outputs(4726)));
    layer3_outputs(1584) <= (layer2_outputs(3034)) and not (layer2_outputs(8324));
    layer3_outputs(1585) <= layer2_outputs(7921);
    layer3_outputs(1586) <= not((layer2_outputs(5375)) xor (layer2_outputs(10102)));
    layer3_outputs(1587) <= not(layer2_outputs(7890));
    layer3_outputs(1588) <= (layer2_outputs(8528)) xor (layer2_outputs(3320));
    layer3_outputs(1589) <= layer2_outputs(3968);
    layer3_outputs(1590) <= not(layer2_outputs(6056));
    layer3_outputs(1591) <= not((layer2_outputs(631)) xor (layer2_outputs(175)));
    layer3_outputs(1592) <= not((layer2_outputs(5058)) or (layer2_outputs(6788)));
    layer3_outputs(1593) <= (layer2_outputs(6742)) or (layer2_outputs(10167));
    layer3_outputs(1594) <= not((layer2_outputs(8311)) xor (layer2_outputs(9364)));
    layer3_outputs(1595) <= (layer2_outputs(8985)) and not (layer2_outputs(1019));
    layer3_outputs(1596) <= not(layer2_outputs(2755)) or (layer2_outputs(3604));
    layer3_outputs(1597) <= not((layer2_outputs(1175)) or (layer2_outputs(9415)));
    layer3_outputs(1598) <= not(layer2_outputs(3516));
    layer3_outputs(1599) <= layer2_outputs(2890);
    layer3_outputs(1600) <= (layer2_outputs(7134)) and not (layer2_outputs(2151));
    layer3_outputs(1601) <= not((layer2_outputs(96)) xor (layer2_outputs(9621)));
    layer3_outputs(1602) <= not(layer2_outputs(812));
    layer3_outputs(1603) <= (layer2_outputs(3723)) or (layer2_outputs(5174));
    layer3_outputs(1604) <= layer2_outputs(6164);
    layer3_outputs(1605) <= layer2_outputs(2555);
    layer3_outputs(1606) <= layer2_outputs(3861);
    layer3_outputs(1607) <= (layer2_outputs(6390)) xor (layer2_outputs(58));
    layer3_outputs(1608) <= '1';
    layer3_outputs(1609) <= layer2_outputs(213);
    layer3_outputs(1610) <= (layer2_outputs(1971)) and not (layer2_outputs(6101));
    layer3_outputs(1611) <= layer2_outputs(4288);
    layer3_outputs(1612) <= (layer2_outputs(5002)) and not (layer2_outputs(7887));
    layer3_outputs(1613) <= not(layer2_outputs(8775));
    layer3_outputs(1614) <= layer2_outputs(2727);
    layer3_outputs(1615) <= not((layer2_outputs(2388)) and (layer2_outputs(2091)));
    layer3_outputs(1616) <= (layer2_outputs(7626)) and not (layer2_outputs(6336));
    layer3_outputs(1617) <= not(layer2_outputs(596));
    layer3_outputs(1618) <= (layer2_outputs(8101)) or (layer2_outputs(10137));
    layer3_outputs(1619) <= not(layer2_outputs(5523)) or (layer2_outputs(3748));
    layer3_outputs(1620) <= not(layer2_outputs(7125)) or (layer2_outputs(2457));
    layer3_outputs(1621) <= not(layer2_outputs(7729));
    layer3_outputs(1622) <= layer2_outputs(7838);
    layer3_outputs(1623) <= not(layer2_outputs(2316));
    layer3_outputs(1624) <= layer2_outputs(967);
    layer3_outputs(1625) <= not(layer2_outputs(8669)) or (layer2_outputs(6058));
    layer3_outputs(1626) <= not(layer2_outputs(3484));
    layer3_outputs(1627) <= layer2_outputs(1744);
    layer3_outputs(1628) <= layer2_outputs(9815);
    layer3_outputs(1629) <= layer2_outputs(7060);
    layer3_outputs(1630) <= not((layer2_outputs(2155)) xor (layer2_outputs(4701)));
    layer3_outputs(1631) <= not((layer2_outputs(3854)) or (layer2_outputs(7371)));
    layer3_outputs(1632) <= (layer2_outputs(8948)) and not (layer2_outputs(8428));
    layer3_outputs(1633) <= layer2_outputs(4779);
    layer3_outputs(1634) <= layer2_outputs(1647);
    layer3_outputs(1635) <= not(layer2_outputs(757));
    layer3_outputs(1636) <= layer2_outputs(1922);
    layer3_outputs(1637) <= not((layer2_outputs(8396)) or (layer2_outputs(9537)));
    layer3_outputs(1638) <= layer2_outputs(9064);
    layer3_outputs(1639) <= '1';
    layer3_outputs(1640) <= (layer2_outputs(3316)) and not (layer2_outputs(9926));
    layer3_outputs(1641) <= (layer2_outputs(4808)) and not (layer2_outputs(9884));
    layer3_outputs(1642) <= not(layer2_outputs(5602)) or (layer2_outputs(5215));
    layer3_outputs(1643) <= not((layer2_outputs(7221)) or (layer2_outputs(7793)));
    layer3_outputs(1644) <= not((layer2_outputs(5955)) xor (layer2_outputs(8089)));
    layer3_outputs(1645) <= not(layer2_outputs(4467));
    layer3_outputs(1646) <= (layer2_outputs(5544)) or (layer2_outputs(9013));
    layer3_outputs(1647) <= not((layer2_outputs(4109)) and (layer2_outputs(4594)));
    layer3_outputs(1648) <= not(layer2_outputs(5054));
    layer3_outputs(1649) <= (layer2_outputs(3212)) and (layer2_outputs(7740));
    layer3_outputs(1650) <= not(layer2_outputs(3929)) or (layer2_outputs(2288));
    layer3_outputs(1651) <= not(layer2_outputs(8656));
    layer3_outputs(1652) <= layer2_outputs(10195);
    layer3_outputs(1653) <= (layer2_outputs(966)) xor (layer2_outputs(2808));
    layer3_outputs(1654) <= not(layer2_outputs(925));
    layer3_outputs(1655) <= layer2_outputs(5908);
    layer3_outputs(1656) <= (layer2_outputs(3018)) xor (layer2_outputs(8064));
    layer3_outputs(1657) <= (layer2_outputs(3138)) and not (layer2_outputs(7245));
    layer3_outputs(1658) <= not((layer2_outputs(2027)) or (layer2_outputs(714)));
    layer3_outputs(1659) <= not(layer2_outputs(5296));
    layer3_outputs(1660) <= not(layer2_outputs(8167));
    layer3_outputs(1661) <= not(layer2_outputs(5853));
    layer3_outputs(1662) <= not(layer2_outputs(573)) or (layer2_outputs(10034));
    layer3_outputs(1663) <= layer2_outputs(4125);
    layer3_outputs(1664) <= not(layer2_outputs(9748));
    layer3_outputs(1665) <= layer2_outputs(1912);
    layer3_outputs(1666) <= layer2_outputs(1984);
    layer3_outputs(1667) <= not(layer2_outputs(2334));
    layer3_outputs(1668) <= not((layer2_outputs(3996)) or (layer2_outputs(5492)));
    layer3_outputs(1669) <= (layer2_outputs(10053)) xor (layer2_outputs(2447));
    layer3_outputs(1670) <= not(layer2_outputs(2489)) or (layer2_outputs(2848));
    layer3_outputs(1671) <= not(layer2_outputs(1833));
    layer3_outputs(1672) <= not(layer2_outputs(1740));
    layer3_outputs(1673) <= not((layer2_outputs(6944)) xor (layer2_outputs(4242)));
    layer3_outputs(1674) <= not(layer2_outputs(9609));
    layer3_outputs(1675) <= not((layer2_outputs(2901)) or (layer2_outputs(1144)));
    layer3_outputs(1676) <= (layer2_outputs(3337)) or (layer2_outputs(5109));
    layer3_outputs(1677) <= (layer2_outputs(8935)) and (layer2_outputs(3659));
    layer3_outputs(1678) <= layer2_outputs(7421);
    layer3_outputs(1679) <= not(layer2_outputs(5170));
    layer3_outputs(1680) <= not(layer2_outputs(2923));
    layer3_outputs(1681) <= layer2_outputs(8114);
    layer3_outputs(1682) <= layer2_outputs(77);
    layer3_outputs(1683) <= not((layer2_outputs(3171)) or (layer2_outputs(559)));
    layer3_outputs(1684) <= (layer2_outputs(8182)) and (layer2_outputs(4751));
    layer3_outputs(1685) <= layer2_outputs(2703);
    layer3_outputs(1686) <= (layer2_outputs(4303)) xor (layer2_outputs(2153));
    layer3_outputs(1687) <= not(layer2_outputs(8670));
    layer3_outputs(1688) <= (layer2_outputs(8879)) and not (layer2_outputs(5524));
    layer3_outputs(1689) <= not(layer2_outputs(2456)) or (layer2_outputs(8757));
    layer3_outputs(1690) <= not(layer2_outputs(6166));
    layer3_outputs(1691) <= layer2_outputs(8324);
    layer3_outputs(1692) <= not(layer2_outputs(3423)) or (layer2_outputs(4692));
    layer3_outputs(1693) <= not((layer2_outputs(8625)) or (layer2_outputs(6067)));
    layer3_outputs(1694) <= (layer2_outputs(2809)) and not (layer2_outputs(7081));
    layer3_outputs(1695) <= not(layer2_outputs(9633));
    layer3_outputs(1696) <= layer2_outputs(6234);
    layer3_outputs(1697) <= (layer2_outputs(9004)) and not (layer2_outputs(166));
    layer3_outputs(1698) <= layer2_outputs(8537);
    layer3_outputs(1699) <= layer2_outputs(953);
    layer3_outputs(1700) <= layer2_outputs(7537);
    layer3_outputs(1701) <= not(layer2_outputs(9012));
    layer3_outputs(1702) <= not(layer2_outputs(5793));
    layer3_outputs(1703) <= '0';
    layer3_outputs(1704) <= layer2_outputs(429);
    layer3_outputs(1705) <= not(layer2_outputs(6645)) or (layer2_outputs(6369));
    layer3_outputs(1706) <= (layer2_outputs(1036)) or (layer2_outputs(4517));
    layer3_outputs(1707) <= not((layer2_outputs(6279)) and (layer2_outputs(3905)));
    layer3_outputs(1708) <= not(layer2_outputs(7560));
    layer3_outputs(1709) <= not((layer2_outputs(1320)) or (layer2_outputs(5287)));
    layer3_outputs(1710) <= layer2_outputs(2033);
    layer3_outputs(1711) <= '1';
    layer3_outputs(1712) <= not(layer2_outputs(8563));
    layer3_outputs(1713) <= not(layer2_outputs(2800));
    layer3_outputs(1714) <= not(layer2_outputs(5704));
    layer3_outputs(1715) <= '1';
    layer3_outputs(1716) <= (layer2_outputs(5326)) and not (layer2_outputs(8029));
    layer3_outputs(1717) <= (layer2_outputs(8984)) or (layer2_outputs(7215));
    layer3_outputs(1718) <= (layer2_outputs(7576)) and not (layer2_outputs(6919));
    layer3_outputs(1719) <= layer2_outputs(5224);
    layer3_outputs(1720) <= (layer2_outputs(5242)) xor (layer2_outputs(6111));
    layer3_outputs(1721) <= not(layer2_outputs(2706));
    layer3_outputs(1722) <= not(layer2_outputs(396));
    layer3_outputs(1723) <= not(layer2_outputs(6143));
    layer3_outputs(1724) <= not(layer2_outputs(8681));
    layer3_outputs(1725) <= layer2_outputs(3043);
    layer3_outputs(1726) <= not((layer2_outputs(6225)) xor (layer2_outputs(9930)));
    layer3_outputs(1727) <= layer2_outputs(8795);
    layer3_outputs(1728) <= layer2_outputs(2665);
    layer3_outputs(1729) <= layer2_outputs(3567);
    layer3_outputs(1730) <= layer2_outputs(6955);
    layer3_outputs(1731) <= layer2_outputs(9370);
    layer3_outputs(1732) <= not((layer2_outputs(3116)) and (layer2_outputs(1638)));
    layer3_outputs(1733) <= '1';
    layer3_outputs(1734) <= layer2_outputs(8433);
    layer3_outputs(1735) <= not(layer2_outputs(1097)) or (layer2_outputs(899));
    layer3_outputs(1736) <= layer2_outputs(3532);
    layer3_outputs(1737) <= layer2_outputs(8862);
    layer3_outputs(1738) <= (layer2_outputs(1147)) and (layer2_outputs(6067));
    layer3_outputs(1739) <= not(layer2_outputs(8393)) or (layer2_outputs(4248));
    layer3_outputs(1740) <= (layer2_outputs(1607)) xor (layer2_outputs(6202));
    layer3_outputs(1741) <= not((layer2_outputs(1536)) xor (layer2_outputs(2625)));
    layer3_outputs(1742) <= layer2_outputs(6704);
    layer3_outputs(1743) <= layer2_outputs(1442);
    layer3_outputs(1744) <= not(layer2_outputs(4565));
    layer3_outputs(1745) <= layer2_outputs(3726);
    layer3_outputs(1746) <= (layer2_outputs(5476)) xor (layer2_outputs(8600));
    layer3_outputs(1747) <= not((layer2_outputs(4414)) or (layer2_outputs(6108)));
    layer3_outputs(1748) <= (layer2_outputs(7661)) and (layer2_outputs(5014));
    layer3_outputs(1749) <= '0';
    layer3_outputs(1750) <= layer2_outputs(1684);
    layer3_outputs(1751) <= layer2_outputs(1899);
    layer3_outputs(1752) <= layer2_outputs(6210);
    layer3_outputs(1753) <= (layer2_outputs(2390)) and (layer2_outputs(3967));
    layer3_outputs(1754) <= (layer2_outputs(1146)) or (layer2_outputs(7511));
    layer3_outputs(1755) <= (layer2_outputs(9260)) xor (layer2_outputs(7524));
    layer3_outputs(1756) <= not((layer2_outputs(2535)) and (layer2_outputs(3460)));
    layer3_outputs(1757) <= not(layer2_outputs(3599));
    layer3_outputs(1758) <= not(layer2_outputs(8465));
    layer3_outputs(1759) <= not(layer2_outputs(4475));
    layer3_outputs(1760) <= not((layer2_outputs(1699)) xor (layer2_outputs(2710)));
    layer3_outputs(1761) <= not(layer2_outputs(8975)) or (layer2_outputs(1128));
    layer3_outputs(1762) <= '1';
    layer3_outputs(1763) <= not(layer2_outputs(9680));
    layer3_outputs(1764) <= (layer2_outputs(2522)) and not (layer2_outputs(6298));
    layer3_outputs(1765) <= (layer2_outputs(3482)) and not (layer2_outputs(9730));
    layer3_outputs(1766) <= not(layer2_outputs(6286)) or (layer2_outputs(9345));
    layer3_outputs(1767) <= not(layer2_outputs(6909));
    layer3_outputs(1768) <= not(layer2_outputs(7956));
    layer3_outputs(1769) <= not((layer2_outputs(6529)) xor (layer2_outputs(9208)));
    layer3_outputs(1770) <= not(layer2_outputs(74));
    layer3_outputs(1771) <= not(layer2_outputs(5940));
    layer3_outputs(1772) <= (layer2_outputs(10132)) xor (layer2_outputs(577));
    layer3_outputs(1773) <= not(layer2_outputs(6310));
    layer3_outputs(1774) <= not(layer2_outputs(6923)) or (layer2_outputs(337));
    layer3_outputs(1775) <= not(layer2_outputs(3633));
    layer3_outputs(1776) <= layer2_outputs(3402);
    layer3_outputs(1777) <= not(layer2_outputs(5416));
    layer3_outputs(1778) <= not(layer2_outputs(2753)) or (layer2_outputs(9220));
    layer3_outputs(1779) <= layer2_outputs(4706);
    layer3_outputs(1780) <= not(layer2_outputs(5409));
    layer3_outputs(1781) <= not(layer2_outputs(5439));
    layer3_outputs(1782) <= not(layer2_outputs(2600)) or (layer2_outputs(6262));
    layer3_outputs(1783) <= (layer2_outputs(7848)) xor (layer2_outputs(139));
    layer3_outputs(1784) <= layer2_outputs(5063);
    layer3_outputs(1785) <= not(layer2_outputs(8110));
    layer3_outputs(1786) <= (layer2_outputs(9150)) and not (layer2_outputs(1428));
    layer3_outputs(1787) <= (layer2_outputs(4332)) xor (layer2_outputs(7659));
    layer3_outputs(1788) <= not(layer2_outputs(2089)) or (layer2_outputs(8450));
    layer3_outputs(1789) <= (layer2_outputs(543)) and (layer2_outputs(5899));
    layer3_outputs(1790) <= not(layer2_outputs(5731)) or (layer2_outputs(8258));
    layer3_outputs(1791) <= layer2_outputs(5264);
    layer3_outputs(1792) <= not(layer2_outputs(3793));
    layer3_outputs(1793) <= layer2_outputs(7322);
    layer3_outputs(1794) <= (layer2_outputs(3466)) and (layer2_outputs(1850));
    layer3_outputs(1795) <= not(layer2_outputs(7163));
    layer3_outputs(1796) <= (layer2_outputs(8149)) and not (layer2_outputs(4662));
    layer3_outputs(1797) <= layer2_outputs(3230);
    layer3_outputs(1798) <= not((layer2_outputs(5407)) or (layer2_outputs(2309)));
    layer3_outputs(1799) <= layer2_outputs(6560);
    layer3_outputs(1800) <= not((layer2_outputs(5659)) xor (layer2_outputs(9357)));
    layer3_outputs(1801) <= layer2_outputs(9855);
    layer3_outputs(1802) <= not(layer2_outputs(582));
    layer3_outputs(1803) <= not(layer2_outputs(9491));
    layer3_outputs(1804) <= (layer2_outputs(5971)) and (layer2_outputs(3959));
    layer3_outputs(1805) <= (layer2_outputs(9356)) and (layer2_outputs(5093));
    layer3_outputs(1806) <= (layer2_outputs(4776)) and not (layer2_outputs(7899));
    layer3_outputs(1807) <= not((layer2_outputs(2170)) xor (layer2_outputs(4192)));
    layer3_outputs(1808) <= not((layer2_outputs(6397)) or (layer2_outputs(5688)));
    layer3_outputs(1809) <= layer2_outputs(5348);
    layer3_outputs(1810) <= not(layer2_outputs(7643));
    layer3_outputs(1811) <= layer2_outputs(5981);
    layer3_outputs(1812) <= not((layer2_outputs(5263)) and (layer2_outputs(8138)));
    layer3_outputs(1813) <= layer2_outputs(6105);
    layer3_outputs(1814) <= (layer2_outputs(8966)) or (layer2_outputs(3274));
    layer3_outputs(1815) <= '0';
    layer3_outputs(1816) <= layer2_outputs(8344);
    layer3_outputs(1817) <= '0';
    layer3_outputs(1818) <= not(layer2_outputs(5000));
    layer3_outputs(1819) <= not((layer2_outputs(4357)) or (layer2_outputs(486)));
    layer3_outputs(1820) <= not(layer2_outputs(3767));
    layer3_outputs(1821) <= (layer2_outputs(4376)) xor (layer2_outputs(7115));
    layer3_outputs(1822) <= layer2_outputs(9661);
    layer3_outputs(1823) <= not(layer2_outputs(6600));
    layer3_outputs(1824) <= not(layer2_outputs(8168)) or (layer2_outputs(5406));
    layer3_outputs(1825) <= layer2_outputs(5773);
    layer3_outputs(1826) <= '0';
    layer3_outputs(1827) <= layer2_outputs(5943);
    layer3_outputs(1828) <= not(layer2_outputs(5945)) or (layer2_outputs(1518));
    layer3_outputs(1829) <= (layer2_outputs(4073)) xor (layer2_outputs(4851));
    layer3_outputs(1830) <= not((layer2_outputs(6461)) xor (layer2_outputs(2693)));
    layer3_outputs(1831) <= not(layer2_outputs(5237)) or (layer2_outputs(4676));
    layer3_outputs(1832) <= not(layer2_outputs(6244));
    layer3_outputs(1833) <= layer2_outputs(10049);
    layer3_outputs(1834) <= not(layer2_outputs(6761));
    layer3_outputs(1835) <= not(layer2_outputs(6365)) or (layer2_outputs(7231));
    layer3_outputs(1836) <= not((layer2_outputs(5489)) xor (layer2_outputs(8813)));
    layer3_outputs(1837) <= layer2_outputs(7604);
    layer3_outputs(1838) <= layer2_outputs(4922);
    layer3_outputs(1839) <= not(layer2_outputs(8920));
    layer3_outputs(1840) <= layer2_outputs(7293);
    layer3_outputs(1841) <= (layer2_outputs(5760)) xor (layer2_outputs(5381));
    layer3_outputs(1842) <= (layer2_outputs(397)) and not (layer2_outputs(5691));
    layer3_outputs(1843) <= (layer2_outputs(4151)) and not (layer2_outputs(7748));
    layer3_outputs(1844) <= not(layer2_outputs(1031));
    layer3_outputs(1845) <= layer2_outputs(482);
    layer3_outputs(1846) <= layer2_outputs(6548);
    layer3_outputs(1847) <= not(layer2_outputs(4491));
    layer3_outputs(1848) <= not((layer2_outputs(7666)) xor (layer2_outputs(7300)));
    layer3_outputs(1849) <= not(layer2_outputs(1875));
    layer3_outputs(1850) <= not(layer2_outputs(6707));
    layer3_outputs(1851) <= not((layer2_outputs(9345)) or (layer2_outputs(2591)));
    layer3_outputs(1852) <= (layer2_outputs(9005)) xor (layer2_outputs(1649));
    layer3_outputs(1853) <= not((layer2_outputs(3203)) and (layer2_outputs(9110)));
    layer3_outputs(1854) <= (layer2_outputs(9067)) or (layer2_outputs(8626));
    layer3_outputs(1855) <= not((layer2_outputs(1279)) or (layer2_outputs(6477)));
    layer3_outputs(1856) <= not(layer2_outputs(9545));
    layer3_outputs(1857) <= layer2_outputs(4946);
    layer3_outputs(1858) <= (layer2_outputs(5851)) and not (layer2_outputs(8529));
    layer3_outputs(1859) <= (layer2_outputs(3978)) or (layer2_outputs(6223));
    layer3_outputs(1860) <= (layer2_outputs(9799)) and not (layer2_outputs(5355));
    layer3_outputs(1861) <= layer2_outputs(8602);
    layer3_outputs(1862) <= layer2_outputs(5313);
    layer3_outputs(1863) <= not(layer2_outputs(10054));
    layer3_outputs(1864) <= (layer2_outputs(8550)) and not (layer2_outputs(5831));
    layer3_outputs(1865) <= not((layer2_outputs(5114)) and (layer2_outputs(453)));
    layer3_outputs(1866) <= (layer2_outputs(379)) xor (layer2_outputs(4002));
    layer3_outputs(1867) <= not(layer2_outputs(7204));
    layer3_outputs(1868) <= not((layer2_outputs(5940)) xor (layer2_outputs(827)));
    layer3_outputs(1869) <= not(layer2_outputs(6752)) or (layer2_outputs(3099));
    layer3_outputs(1870) <= layer2_outputs(3456);
    layer3_outputs(1871) <= not(layer2_outputs(8109)) or (layer2_outputs(4539));
    layer3_outputs(1872) <= (layer2_outputs(4504)) and not (layer2_outputs(1013));
    layer3_outputs(1873) <= layer2_outputs(194);
    layer3_outputs(1874) <= layer2_outputs(6225);
    layer3_outputs(1875) <= layer2_outputs(1043);
    layer3_outputs(1876) <= not((layer2_outputs(9603)) and (layer2_outputs(4265)));
    layer3_outputs(1877) <= (layer2_outputs(111)) and not (layer2_outputs(5582));
    layer3_outputs(1878) <= '1';
    layer3_outputs(1879) <= not(layer2_outputs(3562)) or (layer2_outputs(6654));
    layer3_outputs(1880) <= (layer2_outputs(5811)) and (layer2_outputs(2324));
    layer3_outputs(1881) <= (layer2_outputs(6761)) xor (layer2_outputs(2509));
    layer3_outputs(1882) <= (layer2_outputs(8942)) and (layer2_outputs(2171));
    layer3_outputs(1883) <= not((layer2_outputs(6976)) and (layer2_outputs(35)));
    layer3_outputs(1884) <= '1';
    layer3_outputs(1885) <= '1';
    layer3_outputs(1886) <= layer2_outputs(3421);
    layer3_outputs(1887) <= layer2_outputs(2525);
    layer3_outputs(1888) <= not(layer2_outputs(2842)) or (layer2_outputs(9076));
    layer3_outputs(1889) <= not((layer2_outputs(922)) and (layer2_outputs(5283)));
    layer3_outputs(1890) <= not(layer2_outputs(7306));
    layer3_outputs(1891) <= not(layer2_outputs(10043));
    layer3_outputs(1892) <= layer2_outputs(7542);
    layer3_outputs(1893) <= not(layer2_outputs(9030)) or (layer2_outputs(7878));
    layer3_outputs(1894) <= (layer2_outputs(478)) and not (layer2_outputs(1173));
    layer3_outputs(1895) <= layer2_outputs(3101);
    layer3_outputs(1896) <= (layer2_outputs(173)) and not (layer2_outputs(9000));
    layer3_outputs(1897) <= (layer2_outputs(164)) xor (layer2_outputs(8389));
    layer3_outputs(1898) <= (layer2_outputs(8891)) and not (layer2_outputs(7828));
    layer3_outputs(1899) <= '1';
    layer3_outputs(1900) <= not((layer2_outputs(9736)) and (layer2_outputs(2485)));
    layer3_outputs(1901) <= not(layer2_outputs(2654));
    layer3_outputs(1902) <= not(layer2_outputs(29));
    layer3_outputs(1903) <= (layer2_outputs(277)) and not (layer2_outputs(6897));
    layer3_outputs(1904) <= not(layer2_outputs(4277));
    layer3_outputs(1905) <= '0';
    layer3_outputs(1906) <= not((layer2_outputs(9382)) and (layer2_outputs(1751)));
    layer3_outputs(1907) <= (layer2_outputs(8816)) and not (layer2_outputs(5802));
    layer3_outputs(1908) <= not(layer2_outputs(1537)) or (layer2_outputs(4740));
    layer3_outputs(1909) <= (layer2_outputs(9155)) and (layer2_outputs(2696));
    layer3_outputs(1910) <= not(layer2_outputs(6186));
    layer3_outputs(1911) <= layer2_outputs(601);
    layer3_outputs(1912) <= not(layer2_outputs(8257));
    layer3_outputs(1913) <= '1';
    layer3_outputs(1914) <= not((layer2_outputs(660)) xor (layer2_outputs(6509)));
    layer3_outputs(1915) <= not(layer2_outputs(3481));
    layer3_outputs(1916) <= not(layer2_outputs(9966)) or (layer2_outputs(916));
    layer3_outputs(1917) <= (layer2_outputs(2644)) xor (layer2_outputs(4253));
    layer3_outputs(1918) <= (layer2_outputs(8461)) and not (layer2_outputs(375));
    layer3_outputs(1919) <= (layer2_outputs(9045)) xor (layer2_outputs(8007));
    layer3_outputs(1920) <= not(layer2_outputs(9666));
    layer3_outputs(1921) <= not((layer2_outputs(6771)) xor (layer2_outputs(7721)));
    layer3_outputs(1922) <= not((layer2_outputs(10171)) xor (layer2_outputs(9320)));
    layer3_outputs(1923) <= (layer2_outputs(8607)) or (layer2_outputs(1546));
    layer3_outputs(1924) <= (layer2_outputs(7107)) and not (layer2_outputs(6504));
    layer3_outputs(1925) <= not(layer2_outputs(5071));
    layer3_outputs(1926) <= layer2_outputs(566);
    layer3_outputs(1927) <= layer2_outputs(9859);
    layer3_outputs(1928) <= (layer2_outputs(7786)) and not (layer2_outputs(338));
    layer3_outputs(1929) <= not(layer2_outputs(2065));
    layer3_outputs(1930) <= '0';
    layer3_outputs(1931) <= (layer2_outputs(4318)) and not (layer2_outputs(649));
    layer3_outputs(1932) <= (layer2_outputs(8865)) and not (layer2_outputs(9932));
    layer3_outputs(1933) <= '1';
    layer3_outputs(1934) <= not((layer2_outputs(2929)) or (layer2_outputs(4959)));
    layer3_outputs(1935) <= layer2_outputs(9916);
    layer3_outputs(1936) <= not(layer2_outputs(8005));
    layer3_outputs(1937) <= not(layer2_outputs(3690));
    layer3_outputs(1938) <= not(layer2_outputs(8865));
    layer3_outputs(1939) <= not(layer2_outputs(7961)) or (layer2_outputs(10077));
    layer3_outputs(1940) <= layer2_outputs(9974);
    layer3_outputs(1941) <= not(layer2_outputs(10115));
    layer3_outputs(1942) <= (layer2_outputs(5669)) and (layer2_outputs(4010));
    layer3_outputs(1943) <= not((layer2_outputs(6842)) and (layer2_outputs(5555)));
    layer3_outputs(1944) <= not((layer2_outputs(6104)) xor (layer2_outputs(7477)));
    layer3_outputs(1945) <= (layer2_outputs(995)) or (layer2_outputs(8749));
    layer3_outputs(1946) <= not(layer2_outputs(8568));
    layer3_outputs(1947) <= layer2_outputs(33);
    layer3_outputs(1948) <= not(layer2_outputs(6152)) or (layer2_outputs(8833));
    layer3_outputs(1949) <= (layer2_outputs(7822)) xor (layer2_outputs(7184));
    layer3_outputs(1950) <= (layer2_outputs(6850)) and not (layer2_outputs(35));
    layer3_outputs(1951) <= not(layer2_outputs(8432));
    layer3_outputs(1952) <= layer2_outputs(9916);
    layer3_outputs(1953) <= layer2_outputs(5297);
    layer3_outputs(1954) <= not(layer2_outputs(4999));
    layer3_outputs(1955) <= (layer2_outputs(2371)) or (layer2_outputs(7267));
    layer3_outputs(1956) <= not(layer2_outputs(10172));
    layer3_outputs(1957) <= not(layer2_outputs(6457));
    layer3_outputs(1958) <= layer2_outputs(7602);
    layer3_outputs(1959) <= not((layer2_outputs(7359)) and (layer2_outputs(95)));
    layer3_outputs(1960) <= not(layer2_outputs(9482)) or (layer2_outputs(211));
    layer3_outputs(1961) <= layer2_outputs(397);
    layer3_outputs(1962) <= '1';
    layer3_outputs(1963) <= layer2_outputs(1500);
    layer3_outputs(1964) <= not(layer2_outputs(5212));
    layer3_outputs(1965) <= not(layer2_outputs(767));
    layer3_outputs(1966) <= not(layer2_outputs(10002)) or (layer2_outputs(5690));
    layer3_outputs(1967) <= layer2_outputs(3237);
    layer3_outputs(1968) <= not(layer2_outputs(5192)) or (layer2_outputs(4216));
    layer3_outputs(1969) <= '0';
    layer3_outputs(1970) <= not(layer2_outputs(8390));
    layer3_outputs(1971) <= not(layer2_outputs(9824));
    layer3_outputs(1972) <= (layer2_outputs(7776)) and not (layer2_outputs(518));
    layer3_outputs(1973) <= (layer2_outputs(3299)) or (layer2_outputs(652));
    layer3_outputs(1974) <= '1';
    layer3_outputs(1975) <= layer2_outputs(4442);
    layer3_outputs(1976) <= (layer2_outputs(2722)) and not (layer2_outputs(5527));
    layer3_outputs(1977) <= layer2_outputs(7369);
    layer3_outputs(1978) <= not((layer2_outputs(9473)) xor (layer2_outputs(966)));
    layer3_outputs(1979) <= layer2_outputs(2068);
    layer3_outputs(1980) <= layer2_outputs(5078);
    layer3_outputs(1981) <= not((layer2_outputs(9200)) and (layer2_outputs(2065)));
    layer3_outputs(1982) <= (layer2_outputs(9366)) xor (layer2_outputs(1568));
    layer3_outputs(1983) <= (layer2_outputs(9542)) or (layer2_outputs(9938));
    layer3_outputs(1984) <= not((layer2_outputs(3700)) and (layer2_outputs(6798)));
    layer3_outputs(1985) <= not((layer2_outputs(6531)) xor (layer2_outputs(1424)));
    layer3_outputs(1986) <= layer2_outputs(41);
    layer3_outputs(1987) <= (layer2_outputs(656)) or (layer2_outputs(6517));
    layer3_outputs(1988) <= layer2_outputs(5187);
    layer3_outputs(1989) <= layer2_outputs(5760);
    layer3_outputs(1990) <= (layer2_outputs(4207)) xor (layer2_outputs(9485));
    layer3_outputs(1991) <= layer2_outputs(7731);
    layer3_outputs(1992) <= '0';
    layer3_outputs(1993) <= not(layer2_outputs(10021));
    layer3_outputs(1994) <= not(layer2_outputs(8548));
    layer3_outputs(1995) <= not(layer2_outputs(2759));
    layer3_outputs(1996) <= not(layer2_outputs(5768));
    layer3_outputs(1997) <= layer2_outputs(280);
    layer3_outputs(1998) <= not(layer2_outputs(6804));
    layer3_outputs(1999) <= not(layer2_outputs(550));
    layer3_outputs(2000) <= not((layer2_outputs(5892)) or (layer2_outputs(3225)));
    layer3_outputs(2001) <= not(layer2_outputs(56));
    layer3_outputs(2002) <= not(layer2_outputs(7854));
    layer3_outputs(2003) <= (layer2_outputs(5814)) or (layer2_outputs(5265));
    layer3_outputs(2004) <= '1';
    layer3_outputs(2005) <= not(layer2_outputs(3759));
    layer3_outputs(2006) <= not((layer2_outputs(6313)) and (layer2_outputs(387)));
    layer3_outputs(2007) <= not(layer2_outputs(828)) or (layer2_outputs(6214));
    layer3_outputs(2008) <= (layer2_outputs(2379)) and not (layer2_outputs(7626));
    layer3_outputs(2009) <= (layer2_outputs(9433)) and not (layer2_outputs(7294));
    layer3_outputs(2010) <= (layer2_outputs(7319)) or (layer2_outputs(6000));
    layer3_outputs(2011) <= not(layer2_outputs(3230)) or (layer2_outputs(2793));
    layer3_outputs(2012) <= not(layer2_outputs(2493));
    layer3_outputs(2013) <= not(layer2_outputs(8726));
    layer3_outputs(2014) <= layer2_outputs(1311);
    layer3_outputs(2015) <= not(layer2_outputs(8496));
    layer3_outputs(2016) <= not((layer2_outputs(4849)) xor (layer2_outputs(4460)));
    layer3_outputs(2017) <= not(layer2_outputs(7185));
    layer3_outputs(2018) <= layer2_outputs(810);
    layer3_outputs(2019) <= (layer2_outputs(1199)) and not (layer2_outputs(7882));
    layer3_outputs(2020) <= (layer2_outputs(5960)) and (layer2_outputs(1126));
    layer3_outputs(2021) <= not(layer2_outputs(6578));
    layer3_outputs(2022) <= not(layer2_outputs(7765)) or (layer2_outputs(7354));
    layer3_outputs(2023) <= not(layer2_outputs(1572));
    layer3_outputs(2024) <= '1';
    layer3_outputs(2025) <= not((layer2_outputs(2851)) xor (layer2_outputs(2583)));
    layer3_outputs(2026) <= '1';
    layer3_outputs(2027) <= (layer2_outputs(3928)) and not (layer2_outputs(4165));
    layer3_outputs(2028) <= layer2_outputs(8645);
    layer3_outputs(2029) <= not((layer2_outputs(8479)) and (layer2_outputs(4626)));
    layer3_outputs(2030) <= not(layer2_outputs(6172));
    layer3_outputs(2031) <= not(layer2_outputs(4177));
    layer3_outputs(2032) <= not((layer2_outputs(9108)) and (layer2_outputs(1024)));
    layer3_outputs(2033) <= not((layer2_outputs(6670)) or (layer2_outputs(6506)));
    layer3_outputs(2034) <= (layer2_outputs(1625)) and not (layer2_outputs(3149));
    layer3_outputs(2035) <= not(layer2_outputs(8708));
    layer3_outputs(2036) <= (layer2_outputs(2823)) and not (layer2_outputs(5386));
    layer3_outputs(2037) <= (layer2_outputs(2484)) or (layer2_outputs(3340));
    layer3_outputs(2038) <= layer2_outputs(5250);
    layer3_outputs(2039) <= layer2_outputs(9016);
    layer3_outputs(2040) <= not((layer2_outputs(8802)) or (layer2_outputs(4664)));
    layer3_outputs(2041) <= (layer2_outputs(1848)) or (layer2_outputs(7070));
    layer3_outputs(2042) <= (layer2_outputs(9115)) or (layer2_outputs(7717));
    layer3_outputs(2043) <= (layer2_outputs(2766)) and (layer2_outputs(6245));
    layer3_outputs(2044) <= layer2_outputs(9974);
    layer3_outputs(2045) <= layer2_outputs(5360);
    layer3_outputs(2046) <= layer2_outputs(7671);
    layer3_outputs(2047) <= not(layer2_outputs(1296));
    layer3_outputs(2048) <= (layer2_outputs(7258)) and not (layer2_outputs(1057));
    layer3_outputs(2049) <= (layer2_outputs(7058)) and not (layer2_outputs(6700));
    layer3_outputs(2050) <= not(layer2_outputs(2409));
    layer3_outputs(2051) <= layer2_outputs(8221);
    layer3_outputs(2052) <= layer2_outputs(719);
    layer3_outputs(2053) <= not(layer2_outputs(3566));
    layer3_outputs(2054) <= not((layer2_outputs(4592)) or (layer2_outputs(5401)));
    layer3_outputs(2055) <= layer2_outputs(7664);
    layer3_outputs(2056) <= (layer2_outputs(5282)) xor (layer2_outputs(9500));
    layer3_outputs(2057) <= not((layer2_outputs(6522)) and (layer2_outputs(312)));
    layer3_outputs(2058) <= (layer2_outputs(8347)) xor (layer2_outputs(2963));
    layer3_outputs(2059) <= (layer2_outputs(788)) or (layer2_outputs(9597));
    layer3_outputs(2060) <= (layer2_outputs(9451)) xor (layer2_outputs(7705));
    layer3_outputs(2061) <= not(layer2_outputs(2276)) or (layer2_outputs(4279));
    layer3_outputs(2062) <= layer2_outputs(7749);
    layer3_outputs(2063) <= not(layer2_outputs(2714));
    layer3_outputs(2064) <= not(layer2_outputs(9134)) or (layer2_outputs(6440));
    layer3_outputs(2065) <= not((layer2_outputs(5565)) and (layer2_outputs(3603)));
    layer3_outputs(2066) <= (layer2_outputs(3525)) and not (layer2_outputs(1005));
    layer3_outputs(2067) <= (layer2_outputs(3788)) and not (layer2_outputs(3321));
    layer3_outputs(2068) <= (layer2_outputs(8983)) xor (layer2_outputs(9095));
    layer3_outputs(2069) <= not((layer2_outputs(3955)) and (layer2_outputs(3478)));
    layer3_outputs(2070) <= '1';
    layer3_outputs(2071) <= not(layer2_outputs(2374));
    layer3_outputs(2072) <= (layer2_outputs(2123)) xor (layer2_outputs(4813));
    layer3_outputs(2073) <= not(layer2_outputs(8476));
    layer3_outputs(2074) <= (layer2_outputs(9819)) and (layer2_outputs(3753));
    layer3_outputs(2075) <= not((layer2_outputs(233)) xor (layer2_outputs(5888)));
    layer3_outputs(2076) <= (layer2_outputs(4752)) xor (layer2_outputs(339));
    layer3_outputs(2077) <= not(layer2_outputs(366)) or (layer2_outputs(9332));
    layer3_outputs(2078) <= not((layer2_outputs(3734)) and (layer2_outputs(8241)));
    layer3_outputs(2079) <= layer2_outputs(5529);
    layer3_outputs(2080) <= not((layer2_outputs(1788)) and (layer2_outputs(7498)));
    layer3_outputs(2081) <= (layer2_outputs(3550)) xor (layer2_outputs(8048));
    layer3_outputs(2082) <= (layer2_outputs(5695)) xor (layer2_outputs(1708));
    layer3_outputs(2083) <= layer2_outputs(3717);
    layer3_outputs(2084) <= layer2_outputs(8488);
    layer3_outputs(2085) <= not(layer2_outputs(253));
    layer3_outputs(2086) <= layer2_outputs(1151);
    layer3_outputs(2087) <= layer2_outputs(5154);
    layer3_outputs(2088) <= not((layer2_outputs(5722)) or (layer2_outputs(6277)));
    layer3_outputs(2089) <= not(layer2_outputs(6718)) or (layer2_outputs(8465));
    layer3_outputs(2090) <= not(layer2_outputs(8510));
    layer3_outputs(2091) <= not(layer2_outputs(4360));
    layer3_outputs(2092) <= '1';
    layer3_outputs(2093) <= not(layer2_outputs(5720)) or (layer2_outputs(10029));
    layer3_outputs(2094) <= not(layer2_outputs(9553));
    layer3_outputs(2095) <= layer2_outputs(7517);
    layer3_outputs(2096) <= layer2_outputs(7009);
    layer3_outputs(2097) <= not(layer2_outputs(9007));
    layer3_outputs(2098) <= (layer2_outputs(4153)) and not (layer2_outputs(9793));
    layer3_outputs(2099) <= (layer2_outputs(5845)) and (layer2_outputs(833));
    layer3_outputs(2100) <= not(layer2_outputs(2254)) or (layer2_outputs(1093));
    layer3_outputs(2101) <= (layer2_outputs(9498)) and not (layer2_outputs(1653));
    layer3_outputs(2102) <= (layer2_outputs(8612)) xor (layer2_outputs(5708));
    layer3_outputs(2103) <= not((layer2_outputs(1977)) xor (layer2_outputs(9029)));
    layer3_outputs(2104) <= layer2_outputs(3362);
    layer3_outputs(2105) <= layer2_outputs(1729);
    layer3_outputs(2106) <= not((layer2_outputs(7289)) or (layer2_outputs(9404)));
    layer3_outputs(2107) <= not((layer2_outputs(6665)) and (layer2_outputs(5449)));
    layer3_outputs(2108) <= not(layer2_outputs(9457));
    layer3_outputs(2109) <= not(layer2_outputs(4351)) or (layer2_outputs(9928));
    layer3_outputs(2110) <= not((layer2_outputs(7713)) or (layer2_outputs(5466)));
    layer3_outputs(2111) <= not(layer2_outputs(3582));
    layer3_outputs(2112) <= (layer2_outputs(2914)) and not (layer2_outputs(1086));
    layer3_outputs(2113) <= layer2_outputs(6086);
    layer3_outputs(2114) <= not(layer2_outputs(459)) or (layer2_outputs(6352));
    layer3_outputs(2115) <= '1';
    layer3_outputs(2116) <= layer2_outputs(10142);
    layer3_outputs(2117) <= not(layer2_outputs(9934));
    layer3_outputs(2118) <= not(layer2_outputs(4503)) or (layer2_outputs(3410));
    layer3_outputs(2119) <= layer2_outputs(4424);
    layer3_outputs(2120) <= layer2_outputs(1600);
    layer3_outputs(2121) <= '0';
    layer3_outputs(2122) <= layer2_outputs(6050);
    layer3_outputs(2123) <= not(layer2_outputs(1545));
    layer3_outputs(2124) <= not(layer2_outputs(2362)) or (layer2_outputs(3765));
    layer3_outputs(2125) <= (layer2_outputs(1817)) and not (layer2_outputs(10012));
    layer3_outputs(2126) <= layer2_outputs(8449);
    layer3_outputs(2127) <= not((layer2_outputs(566)) and (layer2_outputs(4492)));
    layer3_outputs(2128) <= not((layer2_outputs(7757)) xor (layer2_outputs(3634)));
    layer3_outputs(2129) <= layer2_outputs(8763);
    layer3_outputs(2130) <= (layer2_outputs(4499)) and (layer2_outputs(8144));
    layer3_outputs(2131) <= (layer2_outputs(7383)) and (layer2_outputs(4356));
    layer3_outputs(2132) <= not((layer2_outputs(3844)) and (layer2_outputs(1077)));
    layer3_outputs(2133) <= not((layer2_outputs(6476)) and (layer2_outputs(5769)));
    layer3_outputs(2134) <= not(layer2_outputs(7318));
    layer3_outputs(2135) <= layer2_outputs(408);
    layer3_outputs(2136) <= not(layer2_outputs(4311)) or (layer2_outputs(1124));
    layer3_outputs(2137) <= layer2_outputs(5794);
    layer3_outputs(2138) <= not(layer2_outputs(4348));
    layer3_outputs(2139) <= layer2_outputs(5526);
    layer3_outputs(2140) <= not((layer2_outputs(865)) and (layer2_outputs(1501)));
    layer3_outputs(2141) <= not((layer2_outputs(4438)) or (layer2_outputs(6310)));
    layer3_outputs(2142) <= not(layer2_outputs(461));
    layer3_outputs(2143) <= layer2_outputs(5357);
    layer3_outputs(2144) <= not((layer2_outputs(1059)) and (layer2_outputs(2034)));
    layer3_outputs(2145) <= (layer2_outputs(1504)) or (layer2_outputs(5585));
    layer3_outputs(2146) <= not(layer2_outputs(789)) or (layer2_outputs(8869));
    layer3_outputs(2147) <= (layer2_outputs(509)) and not (layer2_outputs(290));
    layer3_outputs(2148) <= (layer2_outputs(5982)) and not (layer2_outputs(336));
    layer3_outputs(2149) <= layer2_outputs(8679);
    layer3_outputs(2150) <= not(layer2_outputs(7396));
    layer3_outputs(2151) <= layer2_outputs(2460);
    layer3_outputs(2152) <= (layer2_outputs(1610)) xor (layer2_outputs(4235));
    layer3_outputs(2153) <= layer2_outputs(9847);
    layer3_outputs(2154) <= not(layer2_outputs(2148));
    layer3_outputs(2155) <= not(layer2_outputs(3507)) or (layer2_outputs(7493));
    layer3_outputs(2156) <= '0';
    layer3_outputs(2157) <= (layer2_outputs(242)) and not (layer2_outputs(6396));
    layer3_outputs(2158) <= not((layer2_outputs(3557)) and (layer2_outputs(6096)));
    layer3_outputs(2159) <= '1';
    layer3_outputs(2160) <= (layer2_outputs(810)) or (layer2_outputs(10221));
    layer3_outputs(2161) <= not(layer2_outputs(9270));
    layer3_outputs(2162) <= layer2_outputs(9596);
    layer3_outputs(2163) <= not(layer2_outputs(8267)) or (layer2_outputs(6733));
    layer3_outputs(2164) <= not(layer2_outputs(2236));
    layer3_outputs(2165) <= not(layer2_outputs(354));
    layer3_outputs(2166) <= (layer2_outputs(390)) and not (layer2_outputs(10045));
    layer3_outputs(2167) <= layer2_outputs(9719);
    layer3_outputs(2168) <= (layer2_outputs(636)) xor (layer2_outputs(3047));
    layer3_outputs(2169) <= (layer2_outputs(2334)) and not (layer2_outputs(3006));
    layer3_outputs(2170) <= layer2_outputs(1048);
    layer3_outputs(2171) <= not(layer2_outputs(1255));
    layer3_outputs(2172) <= not(layer2_outputs(8376));
    layer3_outputs(2173) <= not(layer2_outputs(1214));
    layer3_outputs(2174) <= not(layer2_outputs(5478));
    layer3_outputs(2175) <= (layer2_outputs(5412)) and not (layer2_outputs(6276));
    layer3_outputs(2176) <= '1';
    layer3_outputs(2177) <= layer2_outputs(299);
    layer3_outputs(2178) <= layer2_outputs(2883);
    layer3_outputs(2179) <= (layer2_outputs(4034)) and not (layer2_outputs(1048));
    layer3_outputs(2180) <= layer2_outputs(1516);
    layer3_outputs(2181) <= (layer2_outputs(2846)) and not (layer2_outputs(4167));
    layer3_outputs(2182) <= (layer2_outputs(9352)) or (layer2_outputs(3447));
    layer3_outputs(2183) <= not((layer2_outputs(932)) and (layer2_outputs(6847)));
    layer3_outputs(2184) <= not((layer2_outputs(7381)) and (layer2_outputs(5452)));
    layer3_outputs(2185) <= not(layer2_outputs(5957));
    layer3_outputs(2186) <= layer2_outputs(3414);
    layer3_outputs(2187) <= layer2_outputs(4806);
    layer3_outputs(2188) <= layer2_outputs(8604);
    layer3_outputs(2189) <= (layer2_outputs(5365)) xor (layer2_outputs(5519));
    layer3_outputs(2190) <= layer2_outputs(1958);
    layer3_outputs(2191) <= (layer2_outputs(6593)) or (layer2_outputs(2280));
    layer3_outputs(2192) <= '0';
    layer3_outputs(2193) <= not((layer2_outputs(6933)) xor (layer2_outputs(705)));
    layer3_outputs(2194) <= (layer2_outputs(1458)) and not (layer2_outputs(9550));
    layer3_outputs(2195) <= not(layer2_outputs(4275)) or (layer2_outputs(552));
    layer3_outputs(2196) <= not(layer2_outputs(253));
    layer3_outputs(2197) <= layer2_outputs(8653);
    layer3_outputs(2198) <= '1';
    layer3_outputs(2199) <= not((layer2_outputs(3719)) xor (layer2_outputs(5186)));
    layer3_outputs(2200) <= not((layer2_outputs(2770)) xor (layer2_outputs(4093)));
    layer3_outputs(2201) <= (layer2_outputs(2174)) and not (layer2_outputs(400));
    layer3_outputs(2202) <= not((layer2_outputs(2687)) or (layer2_outputs(3646)));
    layer3_outputs(2203) <= not(layer2_outputs(4665));
    layer3_outputs(2204) <= not((layer2_outputs(4464)) or (layer2_outputs(3982)));
    layer3_outputs(2205) <= (layer2_outputs(6370)) and not (layer2_outputs(6012));
    layer3_outputs(2206) <= not(layer2_outputs(7002));
    layer3_outputs(2207) <= layer2_outputs(24);
    layer3_outputs(2208) <= not(layer2_outputs(6326));
    layer3_outputs(2209) <= not(layer2_outputs(2850));
    layer3_outputs(2210) <= not(layer2_outputs(8847)) or (layer2_outputs(8896));
    layer3_outputs(2211) <= not(layer2_outputs(4189));
    layer3_outputs(2212) <= not(layer2_outputs(9926));
    layer3_outputs(2213) <= layer2_outputs(1938);
    layer3_outputs(2214) <= not(layer2_outputs(9008));
    layer3_outputs(2215) <= not(layer2_outputs(5037));
    layer3_outputs(2216) <= (layer2_outputs(958)) and not (layer2_outputs(308));
    layer3_outputs(2217) <= not(layer2_outputs(9286));
    layer3_outputs(2218) <= layer2_outputs(2394);
    layer3_outputs(2219) <= layer2_outputs(851);
    layer3_outputs(2220) <= layer2_outputs(3381);
    layer3_outputs(2221) <= not(layer2_outputs(327));
    layer3_outputs(2222) <= (layer2_outputs(10226)) xor (layer2_outputs(2896));
    layer3_outputs(2223) <= (layer2_outputs(10087)) and (layer2_outputs(900));
    layer3_outputs(2224) <= (layer2_outputs(2696)) xor (layer2_outputs(393));
    layer3_outputs(2225) <= not((layer2_outputs(1983)) or (layer2_outputs(9401)));
    layer3_outputs(2226) <= (layer2_outputs(6685)) or (layer2_outputs(7743));
    layer3_outputs(2227) <= (layer2_outputs(9510)) and (layer2_outputs(1069));
    layer3_outputs(2228) <= not((layer2_outputs(3113)) and (layer2_outputs(5841)));
    layer3_outputs(2229) <= layer2_outputs(8473);
    layer3_outputs(2230) <= not(layer2_outputs(5067));
    layer3_outputs(2231) <= not(layer2_outputs(9043));
    layer3_outputs(2232) <= not(layer2_outputs(2160));
    layer3_outputs(2233) <= not(layer2_outputs(8640));
    layer3_outputs(2234) <= '0';
    layer3_outputs(2235) <= layer2_outputs(2491);
    layer3_outputs(2236) <= (layer2_outputs(9802)) and (layer2_outputs(5558));
    layer3_outputs(2237) <= not(layer2_outputs(3232));
    layer3_outputs(2238) <= not(layer2_outputs(9929)) or (layer2_outputs(250));
    layer3_outputs(2239) <= (layer2_outputs(6412)) or (layer2_outputs(7481));
    layer3_outputs(2240) <= (layer2_outputs(6604)) and not (layer2_outputs(9375));
    layer3_outputs(2241) <= not(layer2_outputs(1662));
    layer3_outputs(2242) <= (layer2_outputs(1868)) and not (layer2_outputs(1016));
    layer3_outputs(2243) <= layer2_outputs(8863);
    layer3_outputs(2244) <= layer2_outputs(5630);
    layer3_outputs(2245) <= (layer2_outputs(5449)) or (layer2_outputs(4935));
    layer3_outputs(2246) <= not(layer2_outputs(6255)) or (layer2_outputs(5581));
    layer3_outputs(2247) <= not((layer2_outputs(4796)) and (layer2_outputs(3352)));
    layer3_outputs(2248) <= (layer2_outputs(7794)) or (layer2_outputs(3079));
    layer3_outputs(2249) <= (layer2_outputs(6844)) xor (layer2_outputs(5077));
    layer3_outputs(2250) <= layer2_outputs(9216);
    layer3_outputs(2251) <= layer2_outputs(4653);
    layer3_outputs(2252) <= not((layer2_outputs(7605)) and (layer2_outputs(1942)));
    layer3_outputs(2253) <= not((layer2_outputs(5908)) xor (layer2_outputs(6209)));
    layer3_outputs(2254) <= (layer2_outputs(1824)) and not (layer2_outputs(2233));
    layer3_outputs(2255) <= not((layer2_outputs(8897)) or (layer2_outputs(1553)));
    layer3_outputs(2256) <= layer2_outputs(10224);
    layer3_outputs(2257) <= not(layer2_outputs(5426));
    layer3_outputs(2258) <= not((layer2_outputs(10086)) and (layer2_outputs(8464)));
    layer3_outputs(2259) <= not((layer2_outputs(7295)) xor (layer2_outputs(1481)));
    layer3_outputs(2260) <= layer2_outputs(6807);
    layer3_outputs(2261) <= not(layer2_outputs(5175));
    layer3_outputs(2262) <= not(layer2_outputs(6897));
    layer3_outputs(2263) <= not(layer2_outputs(7739));
    layer3_outputs(2264) <= not((layer2_outputs(3813)) and (layer2_outputs(9846)));
    layer3_outputs(2265) <= not(layer2_outputs(6797));
    layer3_outputs(2266) <= layer2_outputs(7231);
    layer3_outputs(2267) <= not((layer2_outputs(9625)) and (layer2_outputs(4682)));
    layer3_outputs(2268) <= (layer2_outputs(1785)) or (layer2_outputs(3748));
    layer3_outputs(2269) <= not(layer2_outputs(8316)) or (layer2_outputs(9908));
    layer3_outputs(2270) <= not(layer2_outputs(484));
    layer3_outputs(2271) <= not(layer2_outputs(1326));
    layer3_outputs(2272) <= layer2_outputs(6938);
    layer3_outputs(2273) <= not(layer2_outputs(1944)) or (layer2_outputs(6267));
    layer3_outputs(2274) <= not((layer2_outputs(6375)) and (layer2_outputs(2773)));
    layer3_outputs(2275) <= layer2_outputs(685);
    layer3_outputs(2276) <= layer2_outputs(7713);
    layer3_outputs(2277) <= not((layer2_outputs(8051)) and (layer2_outputs(5783)));
    layer3_outputs(2278) <= not(layer2_outputs(5188));
    layer3_outputs(2279) <= layer2_outputs(3806);
    layer3_outputs(2280) <= layer2_outputs(8688);
    layer3_outputs(2281) <= not(layer2_outputs(6500));
    layer3_outputs(2282) <= layer2_outputs(4749);
    layer3_outputs(2283) <= (layer2_outputs(5905)) and (layer2_outputs(7066));
    layer3_outputs(2284) <= '0';
    layer3_outputs(2285) <= layer2_outputs(4843);
    layer3_outputs(2286) <= not(layer2_outputs(6832));
    layer3_outputs(2287) <= not((layer2_outputs(898)) or (layer2_outputs(5226)));
    layer3_outputs(2288) <= '1';
    layer3_outputs(2289) <= layer2_outputs(4152);
    layer3_outputs(2290) <= (layer2_outputs(3064)) xor (layer2_outputs(5141));
    layer3_outputs(2291) <= not(layer2_outputs(1187));
    layer3_outputs(2292) <= (layer2_outputs(8486)) and (layer2_outputs(4147));
    layer3_outputs(2293) <= (layer2_outputs(7471)) or (layer2_outputs(3108));
    layer3_outputs(2294) <= not(layer2_outputs(9689));
    layer3_outputs(2295) <= not(layer2_outputs(3073)) or (layer2_outputs(7564));
    layer3_outputs(2296) <= (layer2_outputs(6484)) and (layer2_outputs(4937));
    layer3_outputs(2297) <= not((layer2_outputs(3025)) xor (layer2_outputs(4208)));
    layer3_outputs(2298) <= (layer2_outputs(9227)) xor (layer2_outputs(2857));
    layer3_outputs(2299) <= not(layer2_outputs(10106));
    layer3_outputs(2300) <= (layer2_outputs(417)) and (layer2_outputs(8370));
    layer3_outputs(2301) <= (layer2_outputs(8041)) or (layer2_outputs(202));
    layer3_outputs(2302) <= not(layer2_outputs(9713)) or (layer2_outputs(7795));
    layer3_outputs(2303) <= not(layer2_outputs(3644));
    layer3_outputs(2304) <= layer2_outputs(4377);
    layer3_outputs(2305) <= not(layer2_outputs(6605)) or (layer2_outputs(8162));
    layer3_outputs(2306) <= not((layer2_outputs(4447)) and (layer2_outputs(3042)));
    layer3_outputs(2307) <= (layer2_outputs(7685)) and not (layer2_outputs(6483));
    layer3_outputs(2308) <= layer2_outputs(9722);
    layer3_outputs(2309) <= not(layer2_outputs(1266)) or (layer2_outputs(3438));
    layer3_outputs(2310) <= not(layer2_outputs(7674));
    layer3_outputs(2311) <= layer2_outputs(3930);
    layer3_outputs(2312) <= (layer2_outputs(2881)) xor (layer2_outputs(4490));
    layer3_outputs(2313) <= not(layer2_outputs(7895));
    layer3_outputs(2314) <= layer2_outputs(8368);
    layer3_outputs(2315) <= not((layer2_outputs(9493)) or (layer2_outputs(5785)));
    layer3_outputs(2316) <= not(layer2_outputs(646));
    layer3_outputs(2317) <= not(layer2_outputs(2858)) or (layer2_outputs(1686));
    layer3_outputs(2318) <= layer2_outputs(4077);
    layer3_outputs(2319) <= layer2_outputs(1933);
    layer3_outputs(2320) <= not(layer2_outputs(2757)) or (layer2_outputs(6133));
    layer3_outputs(2321) <= not(layer2_outputs(1061));
    layer3_outputs(2322) <= not((layer2_outputs(10237)) or (layer2_outputs(2558)));
    layer3_outputs(2323) <= layer2_outputs(5530);
    layer3_outputs(2324) <= not(layer2_outputs(8973)) or (layer2_outputs(7088));
    layer3_outputs(2325) <= layer2_outputs(5210);
    layer3_outputs(2326) <= layer2_outputs(1469);
    layer3_outputs(2327) <= layer2_outputs(2882);
    layer3_outputs(2328) <= (layer2_outputs(3131)) and not (layer2_outputs(1542));
    layer3_outputs(2329) <= layer2_outputs(2872);
    layer3_outputs(2330) <= not((layer2_outputs(9902)) or (layer2_outputs(8498)));
    layer3_outputs(2331) <= not(layer2_outputs(3005));
    layer3_outputs(2332) <= not((layer2_outputs(9072)) or (layer2_outputs(3207)));
    layer3_outputs(2333) <= layer2_outputs(2574);
    layer3_outputs(2334) <= '0';
    layer3_outputs(2335) <= (layer2_outputs(1579)) and not (layer2_outputs(4742));
    layer3_outputs(2336) <= not(layer2_outputs(9403)) or (layer2_outputs(6559));
    layer3_outputs(2337) <= not((layer2_outputs(7114)) and (layer2_outputs(7201)));
    layer3_outputs(2338) <= layer2_outputs(2797);
    layer3_outputs(2339) <= not(layer2_outputs(1879));
    layer3_outputs(2340) <= not((layer2_outputs(1891)) and (layer2_outputs(751)));
    layer3_outputs(2341) <= (layer2_outputs(89)) or (layer2_outputs(10119));
    layer3_outputs(2342) <= layer2_outputs(7011);
    layer3_outputs(2343) <= layer2_outputs(781);
    layer3_outputs(2344) <= layer2_outputs(1126);
    layer3_outputs(2345) <= layer2_outputs(4453);
    layer3_outputs(2346) <= layer2_outputs(4437);
    layer3_outputs(2347) <= '1';
    layer3_outputs(2348) <= (layer2_outputs(9469)) and (layer2_outputs(980));
    layer3_outputs(2349) <= layer2_outputs(7514);
    layer3_outputs(2350) <= layer2_outputs(4276);
    layer3_outputs(2351) <= layer2_outputs(9692);
    layer3_outputs(2352) <= not(layer2_outputs(2804));
    layer3_outputs(2353) <= (layer2_outputs(9539)) or (layer2_outputs(9230));
    layer3_outputs(2354) <= (layer2_outputs(9465)) and (layer2_outputs(9872));
    layer3_outputs(2355) <= not(layer2_outputs(7238)) or (layer2_outputs(5211));
    layer3_outputs(2356) <= layer2_outputs(3044);
    layer3_outputs(2357) <= (layer2_outputs(6809)) xor (layer2_outputs(4081));
    layer3_outputs(2358) <= not((layer2_outputs(1877)) and (layer2_outputs(4666)));
    layer3_outputs(2359) <= not((layer2_outputs(759)) xor (layer2_outputs(119)));
    layer3_outputs(2360) <= layer2_outputs(6239);
    layer3_outputs(2361) <= not(layer2_outputs(8765));
    layer3_outputs(2362) <= not(layer2_outputs(6496));
    layer3_outputs(2363) <= not(layer2_outputs(8928));
    layer3_outputs(2364) <= not((layer2_outputs(7032)) xor (layer2_outputs(1299)));
    layer3_outputs(2365) <= not((layer2_outputs(6232)) or (layer2_outputs(4148)));
    layer3_outputs(2366) <= (layer2_outputs(4114)) and (layer2_outputs(7637));
    layer3_outputs(2367) <= not(layer2_outputs(3716));
    layer3_outputs(2368) <= not(layer2_outputs(5203)) or (layer2_outputs(5));
    layer3_outputs(2369) <= layer2_outputs(8596);
    layer3_outputs(2370) <= (layer2_outputs(4341)) xor (layer2_outputs(2870));
    layer3_outputs(2371) <= (layer2_outputs(2397)) and (layer2_outputs(7191));
    layer3_outputs(2372) <= not(layer2_outputs(5052));
    layer3_outputs(2373) <= layer2_outputs(8611);
    layer3_outputs(2374) <= layer2_outputs(8172);
    layer3_outputs(2375) <= '0';
    layer3_outputs(2376) <= not((layer2_outputs(4625)) or (layer2_outputs(2916)));
    layer3_outputs(2377) <= not(layer2_outputs(3851)) or (layer2_outputs(9907));
    layer3_outputs(2378) <= layer2_outputs(4857);
    layer3_outputs(2379) <= layer2_outputs(8779);
    layer3_outputs(2380) <= not((layer2_outputs(9012)) xor (layer2_outputs(5815)));
    layer3_outputs(2381) <= (layer2_outputs(8839)) or (layer2_outputs(5293));
    layer3_outputs(2382) <= not(layer2_outputs(8623)) or (layer2_outputs(8598));
    layer3_outputs(2383) <= not((layer2_outputs(6125)) or (layer2_outputs(1497)));
    layer3_outputs(2384) <= layer2_outputs(7810);
    layer3_outputs(2385) <= not((layer2_outputs(979)) or (layer2_outputs(1029)));
    layer3_outputs(2386) <= not(layer2_outputs(2245));
    layer3_outputs(2387) <= not(layer2_outputs(565));
    layer3_outputs(2388) <= (layer2_outputs(9197)) or (layer2_outputs(4343));
    layer3_outputs(2389) <= not(layer2_outputs(6426));
    layer3_outputs(2390) <= (layer2_outputs(6388)) and not (layer2_outputs(6206));
    layer3_outputs(2391) <= layer2_outputs(2888);
    layer3_outputs(2392) <= not(layer2_outputs(7877)) or (layer2_outputs(8790));
    layer3_outputs(2393) <= layer2_outputs(7410);
    layer3_outputs(2394) <= not((layer2_outputs(7103)) xor (layer2_outputs(9795)));
    layer3_outputs(2395) <= layer2_outputs(8743);
    layer3_outputs(2396) <= not(layer2_outputs(5245));
    layer3_outputs(2397) <= layer2_outputs(2884);
    layer3_outputs(2398) <= not((layer2_outputs(137)) or (layer2_outputs(82)));
    layer3_outputs(2399) <= not(layer2_outputs(5193));
    layer3_outputs(2400) <= not(layer2_outputs(9417));
    layer3_outputs(2401) <= layer2_outputs(878);
    layer3_outputs(2402) <= not(layer2_outputs(4094));
    layer3_outputs(2403) <= (layer2_outputs(3579)) and not (layer2_outputs(8782));
    layer3_outputs(2404) <= layer2_outputs(2668);
    layer3_outputs(2405) <= not((layer2_outputs(9962)) and (layer2_outputs(4114)));
    layer3_outputs(2406) <= not((layer2_outputs(6970)) xor (layer2_outputs(4250)));
    layer3_outputs(2407) <= not((layer2_outputs(4874)) or (layer2_outputs(2935)));
    layer3_outputs(2408) <= not(layer2_outputs(1515));
    layer3_outputs(2409) <= (layer2_outputs(4939)) and (layer2_outputs(519));
    layer3_outputs(2410) <= '1';
    layer3_outputs(2411) <= (layer2_outputs(2047)) or (layer2_outputs(9147));
    layer3_outputs(2412) <= (layer2_outputs(4872)) and (layer2_outputs(9423));
    layer3_outputs(2413) <= (layer2_outputs(1846)) or (layer2_outputs(6021));
    layer3_outputs(2414) <= not(layer2_outputs(6592));
    layer3_outputs(2415) <= not(layer2_outputs(2081)) or (layer2_outputs(4273));
    layer3_outputs(2416) <= not(layer2_outputs(7134));
    layer3_outputs(2417) <= not(layer2_outputs(6033));
    layer3_outputs(2418) <= not(layer2_outputs(5226));
    layer3_outputs(2419) <= not(layer2_outputs(7467));
    layer3_outputs(2420) <= (layer2_outputs(232)) or (layer2_outputs(8457));
    layer3_outputs(2421) <= (layer2_outputs(7979)) and not (layer2_outputs(5484));
    layer3_outputs(2422) <= not((layer2_outputs(6535)) or (layer2_outputs(1376)));
    layer3_outputs(2423) <= (layer2_outputs(3508)) and not (layer2_outputs(6375));
    layer3_outputs(2424) <= layer2_outputs(3099);
    layer3_outputs(2425) <= not(layer2_outputs(4563)) or (layer2_outputs(8158));
    layer3_outputs(2426) <= layer2_outputs(2769);
    layer3_outputs(2427) <= layer2_outputs(6239);
    layer3_outputs(2428) <= (layer2_outputs(2769)) and not (layer2_outputs(1063));
    layer3_outputs(2429) <= (layer2_outputs(5073)) and not (layer2_outputs(4288));
    layer3_outputs(2430) <= not((layer2_outputs(974)) xor (layer2_outputs(2183)));
    layer3_outputs(2431) <= not(layer2_outputs(3459));
    layer3_outputs(2432) <= (layer2_outputs(6572)) or (layer2_outputs(2331));
    layer3_outputs(2433) <= not((layer2_outputs(3384)) or (layer2_outputs(8946)));
    layer3_outputs(2434) <= not((layer2_outputs(8823)) or (layer2_outputs(1436)));
    layer3_outputs(2435) <= not(layer2_outputs(619));
    layer3_outputs(2436) <= layer2_outputs(2232);
    layer3_outputs(2437) <= layer2_outputs(7077);
    layer3_outputs(2438) <= not((layer2_outputs(3649)) xor (layer2_outputs(6623)));
    layer3_outputs(2439) <= not(layer2_outputs(613));
    layer3_outputs(2440) <= layer2_outputs(2587);
    layer3_outputs(2441) <= not(layer2_outputs(2523));
    layer3_outputs(2442) <= (layer2_outputs(4887)) or (layer2_outputs(5894));
    layer3_outputs(2443) <= layer2_outputs(8596);
    layer3_outputs(2444) <= '0';
    layer3_outputs(2445) <= (layer2_outputs(5349)) or (layer2_outputs(9323));
    layer3_outputs(2446) <= not((layer2_outputs(6966)) or (layer2_outputs(8906)));
    layer3_outputs(2447) <= not(layer2_outputs(891));
    layer3_outputs(2448) <= not(layer2_outputs(1087));
    layer3_outputs(2449) <= not(layer2_outputs(7548));
    layer3_outputs(2450) <= layer2_outputs(7343);
    layer3_outputs(2451) <= not(layer2_outputs(3320));
    layer3_outputs(2452) <= (layer2_outputs(8401)) and not (layer2_outputs(1450));
    layer3_outputs(2453) <= (layer2_outputs(8696)) and not (layer2_outputs(2777));
    layer3_outputs(2454) <= (layer2_outputs(1865)) xor (layer2_outputs(3164));
    layer3_outputs(2455) <= (layer2_outputs(6554)) xor (layer2_outputs(5537));
    layer3_outputs(2456) <= (layer2_outputs(6962)) and not (layer2_outputs(3120));
    layer3_outputs(2457) <= (layer2_outputs(9041)) xor (layer2_outputs(4977));
    layer3_outputs(2458) <= layer2_outputs(5117);
    layer3_outputs(2459) <= (layer2_outputs(7451)) or (layer2_outputs(8177));
    layer3_outputs(2460) <= not(layer2_outputs(6512));
    layer3_outputs(2461) <= not(layer2_outputs(3200));
    layer3_outputs(2462) <= not(layer2_outputs(1080));
    layer3_outputs(2463) <= (layer2_outputs(3778)) xor (layer2_outputs(6267));
    layer3_outputs(2464) <= layer2_outputs(10162);
    layer3_outputs(2465) <= not((layer2_outputs(7980)) and (layer2_outputs(10)));
    layer3_outputs(2466) <= layer2_outputs(7356);
    layer3_outputs(2467) <= (layer2_outputs(2984)) xor (layer2_outputs(9159));
    layer3_outputs(2468) <= layer2_outputs(8482);
    layer3_outputs(2469) <= (layer2_outputs(6255)) and (layer2_outputs(8835));
    layer3_outputs(2470) <= (layer2_outputs(10076)) xor (layer2_outputs(5096));
    layer3_outputs(2471) <= '0';
    layer3_outputs(2472) <= layer2_outputs(5732);
    layer3_outputs(2473) <= (layer2_outputs(4860)) xor (layer2_outputs(8425));
    layer3_outputs(2474) <= not(layer2_outputs(2523));
    layer3_outputs(2475) <= not((layer2_outputs(1599)) or (layer2_outputs(2484)));
    layer3_outputs(2476) <= not(layer2_outputs(2500));
    layer3_outputs(2477) <= (layer2_outputs(10159)) and not (layer2_outputs(4585));
    layer3_outputs(2478) <= layer2_outputs(10140);
    layer3_outputs(2479) <= '0';
    layer3_outputs(2480) <= not(layer2_outputs(5522));
    layer3_outputs(2481) <= not(layer2_outputs(4546)) or (layer2_outputs(10072));
    layer3_outputs(2482) <= not(layer2_outputs(7290));
    layer3_outputs(2483) <= '0';
    layer3_outputs(2484) <= (layer2_outputs(1704)) or (layer2_outputs(8530));
    layer3_outputs(2485) <= not(layer2_outputs(2448));
    layer3_outputs(2486) <= not((layer2_outputs(736)) xor (layer2_outputs(4118)));
    layer3_outputs(2487) <= '0';
    layer3_outputs(2488) <= layer2_outputs(3106);
    layer3_outputs(2489) <= layer2_outputs(326);
    layer3_outputs(2490) <= layer2_outputs(5268);
    layer3_outputs(2491) <= not(layer2_outputs(1750));
    layer3_outputs(2492) <= not(layer2_outputs(7224));
    layer3_outputs(2493) <= not(layer2_outputs(2441)) or (layer2_outputs(3874));
    layer3_outputs(2494) <= not(layer2_outputs(8555));
    layer3_outputs(2495) <= layer2_outputs(9888);
    layer3_outputs(2496) <= not(layer2_outputs(1395));
    layer3_outputs(2497) <= (layer2_outputs(5791)) xor (layer2_outputs(3594));
    layer3_outputs(2498) <= not(layer2_outputs(8582)) or (layer2_outputs(6618));
    layer3_outputs(2499) <= layer2_outputs(3980);
    layer3_outputs(2500) <= (layer2_outputs(8441)) and not (layer2_outputs(9799));
    layer3_outputs(2501) <= layer2_outputs(3367);
    layer3_outputs(2502) <= '0';
    layer3_outputs(2503) <= not(layer2_outputs(4519)) or (layer2_outputs(8642));
    layer3_outputs(2504) <= not((layer2_outputs(6040)) and (layer2_outputs(752)));
    layer3_outputs(2505) <= layer2_outputs(261);
    layer3_outputs(2506) <= not(layer2_outputs(9874));
    layer3_outputs(2507) <= layer2_outputs(4552);
    layer3_outputs(2508) <= not(layer2_outputs(9782));
    layer3_outputs(2509) <= '1';
    layer3_outputs(2510) <= not((layer2_outputs(2422)) xor (layer2_outputs(8046)));
    layer3_outputs(2511) <= (layer2_outputs(6313)) xor (layer2_outputs(3454));
    layer3_outputs(2512) <= layer2_outputs(9444);
    layer3_outputs(2513) <= layer2_outputs(6687);
    layer3_outputs(2514) <= not(layer2_outputs(7923));
    layer3_outputs(2515) <= (layer2_outputs(5126)) or (layer2_outputs(1270));
    layer3_outputs(2516) <= not(layer2_outputs(4437));
    layer3_outputs(2517) <= not((layer2_outputs(3222)) and (layer2_outputs(2399)));
    layer3_outputs(2518) <= not(layer2_outputs(6398));
    layer3_outputs(2519) <= layer2_outputs(5085);
    layer3_outputs(2520) <= '1';
    layer3_outputs(2521) <= not((layer2_outputs(5448)) or (layer2_outputs(6337)));
    layer3_outputs(2522) <= not((layer2_outputs(4173)) xor (layer2_outputs(8779)));
    layer3_outputs(2523) <= not(layer2_outputs(1268));
    layer3_outputs(2524) <= (layer2_outputs(7628)) xor (layer2_outputs(9893));
    layer3_outputs(2525) <= not(layer2_outputs(3357));
    layer3_outputs(2526) <= not(layer2_outputs(7539));
    layer3_outputs(2527) <= not(layer2_outputs(5812)) or (layer2_outputs(3781));
    layer3_outputs(2528) <= not(layer2_outputs(70));
    layer3_outputs(2529) <= not(layer2_outputs(3621)) or (layer2_outputs(2053));
    layer3_outputs(2530) <= not(layer2_outputs(2294));
    layer3_outputs(2531) <= (layer2_outputs(6964)) and not (layer2_outputs(7617));
    layer3_outputs(2532) <= not(layer2_outputs(8379));
    layer3_outputs(2533) <= not((layer2_outputs(4078)) and (layer2_outputs(7131)));
    layer3_outputs(2534) <= '0';
    layer3_outputs(2535) <= (layer2_outputs(8447)) and not (layer2_outputs(6468));
    layer3_outputs(2536) <= (layer2_outputs(2613)) xor (layer2_outputs(1760));
    layer3_outputs(2537) <= layer2_outputs(1789);
    layer3_outputs(2538) <= layer2_outputs(2299);
    layer3_outputs(2539) <= not(layer2_outputs(8826));
    layer3_outputs(2540) <= (layer2_outputs(2565)) and not (layer2_outputs(926));
    layer3_outputs(2541) <= not(layer2_outputs(6378)) or (layer2_outputs(4783));
    layer3_outputs(2542) <= layer2_outputs(8919);
    layer3_outputs(2543) <= (layer2_outputs(3428)) xor (layer2_outputs(4985));
    layer3_outputs(2544) <= layer2_outputs(3183);
    layer3_outputs(2545) <= not(layer2_outputs(1264)) or (layer2_outputs(2774));
    layer3_outputs(2546) <= not(layer2_outputs(6102));
    layer3_outputs(2547) <= not(layer2_outputs(5048)) or (layer2_outputs(5391));
    layer3_outputs(2548) <= (layer2_outputs(9131)) xor (layer2_outputs(5160));
    layer3_outputs(2549) <= not((layer2_outputs(2279)) xor (layer2_outputs(3614)));
    layer3_outputs(2550) <= not(layer2_outputs(2727)) or (layer2_outputs(196));
    layer3_outputs(2551) <= (layer2_outputs(7599)) xor (layer2_outputs(562));
    layer3_outputs(2552) <= (layer2_outputs(6281)) or (layer2_outputs(5365));
    layer3_outputs(2553) <= not(layer2_outputs(3334)) or (layer2_outputs(5514));
    layer3_outputs(2554) <= layer2_outputs(7954);
    layer3_outputs(2555) <= layer2_outputs(3834);
    layer3_outputs(2556) <= (layer2_outputs(4015)) xor (layer2_outputs(7650));
    layer3_outputs(2557) <= (layer2_outputs(9761)) and not (layer2_outputs(1798));
    layer3_outputs(2558) <= not(layer2_outputs(843));
    layer3_outputs(2559) <= (layer2_outputs(2681)) xor (layer2_outputs(7196));
    layer3_outputs(2560) <= layer2_outputs(5565);
    layer3_outputs(2561) <= not(layer2_outputs(5060));
    layer3_outputs(2562) <= layer2_outputs(1935);
    layer3_outputs(2563) <= not((layer2_outputs(149)) and (layer2_outputs(8969)));
    layer3_outputs(2564) <= (layer2_outputs(7221)) and not (layer2_outputs(2295));
    layer3_outputs(2565) <= '1';
    layer3_outputs(2566) <= not(layer2_outputs(7887));
    layer3_outputs(2567) <= (layer2_outputs(8676)) and not (layer2_outputs(9885));
    layer3_outputs(2568) <= not(layer2_outputs(8601));
    layer3_outputs(2569) <= (layer2_outputs(47)) and not (layer2_outputs(2643));
    layer3_outputs(2570) <= not((layer2_outputs(9302)) xor (layer2_outputs(2768)));
    layer3_outputs(2571) <= (layer2_outputs(2570)) and (layer2_outputs(10109));
    layer3_outputs(2572) <= not(layer2_outputs(2853));
    layer3_outputs(2573) <= layer2_outputs(6413);
    layer3_outputs(2574) <= not(layer2_outputs(5161));
    layer3_outputs(2575) <= not(layer2_outputs(6024));
    layer3_outputs(2576) <= (layer2_outputs(3434)) and not (layer2_outputs(792));
    layer3_outputs(2577) <= (layer2_outputs(7949)) or (layer2_outputs(999));
    layer3_outputs(2578) <= not(layer2_outputs(3575)) or (layer2_outputs(155));
    layer3_outputs(2579) <= not(layer2_outputs(6902));
    layer3_outputs(2580) <= not(layer2_outputs(5812));
    layer3_outputs(2581) <= layer2_outputs(3873);
    layer3_outputs(2582) <= not(layer2_outputs(8564));
    layer3_outputs(2583) <= (layer2_outputs(4349)) or (layer2_outputs(8871));
    layer3_outputs(2584) <= layer2_outputs(4760);
    layer3_outputs(2585) <= layer2_outputs(8696);
    layer3_outputs(2586) <= layer2_outputs(1559);
    layer3_outputs(2587) <= (layer2_outputs(7933)) and not (layer2_outputs(3879));
    layer3_outputs(2588) <= not((layer2_outputs(5791)) or (layer2_outputs(3611)));
    layer3_outputs(2589) <= not((layer2_outputs(9463)) or (layer2_outputs(999)));
    layer3_outputs(2590) <= not(layer2_outputs(1329));
    layer3_outputs(2591) <= '1';
    layer3_outputs(2592) <= (layer2_outputs(1412)) and not (layer2_outputs(7164));
    layer3_outputs(2593) <= not(layer2_outputs(2142)) or (layer2_outputs(5587));
    layer3_outputs(2594) <= (layer2_outputs(8802)) and (layer2_outputs(1523));
    layer3_outputs(2595) <= not((layer2_outputs(1432)) or (layer2_outputs(8951)));
    layer3_outputs(2596) <= (layer2_outputs(7308)) or (layer2_outputs(9716));
    layer3_outputs(2597) <= not(layer2_outputs(8541)) or (layer2_outputs(4285));
    layer3_outputs(2598) <= not((layer2_outputs(1772)) xor (layer2_outputs(1761)));
    layer3_outputs(2599) <= layer2_outputs(7604);
    layer3_outputs(2600) <= layer2_outputs(7193);
    layer3_outputs(2601) <= not((layer2_outputs(1716)) xor (layer2_outputs(4154)));
    layer3_outputs(2602) <= layer2_outputs(7052);
    layer3_outputs(2603) <= not((layer2_outputs(6168)) or (layer2_outputs(5404)));
    layer3_outputs(2604) <= layer2_outputs(10045);
    layer3_outputs(2605) <= layer2_outputs(6553);
    layer3_outputs(2606) <= (layer2_outputs(763)) and (layer2_outputs(6455));
    layer3_outputs(2607) <= not((layer2_outputs(7610)) and (layer2_outputs(6697)));
    layer3_outputs(2608) <= not((layer2_outputs(1312)) or (layer2_outputs(5433)));
    layer3_outputs(2609) <= (layer2_outputs(10095)) and not (layer2_outputs(8316));
    layer3_outputs(2610) <= (layer2_outputs(1078)) and not (layer2_outputs(1209));
    layer3_outputs(2611) <= layer2_outputs(1682);
    layer3_outputs(2612) <= layer2_outputs(5566);
    layer3_outputs(2613) <= layer2_outputs(6662);
    layer3_outputs(2614) <= '0';
    layer3_outputs(2615) <= (layer2_outputs(4534)) and not (layer2_outputs(6138));
    layer3_outputs(2616) <= not(layer2_outputs(5741));
    layer3_outputs(2617) <= layer2_outputs(2253);
    layer3_outputs(2618) <= not(layer2_outputs(8702));
    layer3_outputs(2619) <= (layer2_outputs(513)) and not (layer2_outputs(6657));
    layer3_outputs(2620) <= layer2_outputs(153);
    layer3_outputs(2621) <= (layer2_outputs(3209)) and not (layer2_outputs(214));
    layer3_outputs(2622) <= not(layer2_outputs(3112));
    layer3_outputs(2623) <= layer2_outputs(9223);
    layer3_outputs(2624) <= not(layer2_outputs(1525));
    layer3_outputs(2625) <= not(layer2_outputs(4479));
    layer3_outputs(2626) <= '1';
    layer3_outputs(2627) <= (layer2_outputs(2630)) and not (layer2_outputs(6590));
    layer3_outputs(2628) <= not(layer2_outputs(5589)) or (layer2_outputs(349));
    layer3_outputs(2629) <= (layer2_outputs(9965)) and not (layer2_outputs(2855));
    layer3_outputs(2630) <= not(layer2_outputs(3302));
    layer3_outputs(2631) <= (layer2_outputs(1631)) and (layer2_outputs(8160));
    layer3_outputs(2632) <= (layer2_outputs(9589)) xor (layer2_outputs(2304));
    layer3_outputs(2633) <= (layer2_outputs(5916)) and not (layer2_outputs(1135));
    layer3_outputs(2634) <= not(layer2_outputs(2968));
    layer3_outputs(2635) <= not(layer2_outputs(4015)) or (layer2_outputs(1078));
    layer3_outputs(2636) <= not(layer2_outputs(7518));
    layer3_outputs(2637) <= layer2_outputs(776);
    layer3_outputs(2638) <= layer2_outputs(10231);
    layer3_outputs(2639) <= not(layer2_outputs(5138));
    layer3_outputs(2640) <= not((layer2_outputs(4059)) xor (layer2_outputs(9983)));
    layer3_outputs(2641) <= not((layer2_outputs(4838)) or (layer2_outputs(5178)));
    layer3_outputs(2642) <= '1';
    layer3_outputs(2643) <= layer2_outputs(7399);
    layer3_outputs(2644) <= not(layer2_outputs(7625));
    layer3_outputs(2645) <= (layer2_outputs(7462)) and not (layer2_outputs(8827));
    layer3_outputs(2646) <= layer2_outputs(5595);
    layer3_outputs(2647) <= (layer2_outputs(8586)) xor (layer2_outputs(6603));
    layer3_outputs(2648) <= not(layer2_outputs(5767)) or (layer2_outputs(7941));
    layer3_outputs(2649) <= (layer2_outputs(7433)) and not (layer2_outputs(5341));
    layer3_outputs(2650) <= (layer2_outputs(1929)) xor (layer2_outputs(2206));
    layer3_outputs(2651) <= not(layer2_outputs(7922));
    layer3_outputs(2652) <= (layer2_outputs(10014)) or (layer2_outputs(1573));
    layer3_outputs(2653) <= (layer2_outputs(5775)) and (layer2_outputs(3600));
    layer3_outputs(2654) <= not(layer2_outputs(8021));
    layer3_outputs(2655) <= not(layer2_outputs(7669));
    layer3_outputs(2656) <= not(layer2_outputs(5993));
    layer3_outputs(2657) <= (layer2_outputs(4669)) and not (layer2_outputs(8214));
    layer3_outputs(2658) <= layer2_outputs(9001);
    layer3_outputs(2659) <= (layer2_outputs(4368)) xor (layer2_outputs(4358));
    layer3_outputs(2660) <= not((layer2_outputs(7871)) or (layer2_outputs(3881)));
    layer3_outputs(2661) <= not(layer2_outputs(10234));
    layer3_outputs(2662) <= not((layer2_outputs(9248)) or (layer2_outputs(9552)));
    layer3_outputs(2663) <= layer2_outputs(9447);
    layer3_outputs(2664) <= not((layer2_outputs(158)) and (layer2_outputs(268)));
    layer3_outputs(2665) <= (layer2_outputs(5316)) and not (layer2_outputs(6198));
    layer3_outputs(2666) <= layer2_outputs(2960);
    layer3_outputs(2667) <= not((layer2_outputs(5427)) or (layer2_outputs(2449)));
    layer3_outputs(2668) <= not(layer2_outputs(6979));
    layer3_outputs(2669) <= (layer2_outputs(3430)) or (layer2_outputs(6403));
    layer3_outputs(2670) <= not(layer2_outputs(6954));
    layer3_outputs(2671) <= layer2_outputs(7621);
    layer3_outputs(2672) <= layer2_outputs(9367);
    layer3_outputs(2673) <= layer2_outputs(6673);
    layer3_outputs(2674) <= layer2_outputs(4296);
    layer3_outputs(2675) <= not(layer2_outputs(2995)) or (layer2_outputs(2802));
    layer3_outputs(2676) <= (layer2_outputs(3357)) and not (layer2_outputs(9509));
    layer3_outputs(2677) <= not(layer2_outputs(5358));
    layer3_outputs(2678) <= layer2_outputs(1150);
    layer3_outputs(2679) <= not((layer2_outputs(92)) or (layer2_outputs(9090)));
    layer3_outputs(2680) <= not(layer2_outputs(7));
    layer3_outputs(2681) <= layer2_outputs(7580);
    layer3_outputs(2682) <= not(layer2_outputs(8708));
    layer3_outputs(2683) <= not((layer2_outputs(1200)) xor (layer2_outputs(6726)));
    layer3_outputs(2684) <= layer2_outputs(1265);
    layer3_outputs(2685) <= layer2_outputs(942);
    layer3_outputs(2686) <= not((layer2_outputs(6774)) xor (layer2_outputs(8763)));
    layer3_outputs(2687) <= not((layer2_outputs(2931)) and (layer2_outputs(9602)));
    layer3_outputs(2688) <= not((layer2_outputs(2268)) and (layer2_outputs(9616)));
    layer3_outputs(2689) <= '1';
    layer3_outputs(2690) <= not(layer2_outputs(5830));
    layer3_outputs(2691) <= (layer2_outputs(8377)) and not (layer2_outputs(394));
    layer3_outputs(2692) <= not(layer2_outputs(9693));
    layer3_outputs(2693) <= (layer2_outputs(10200)) and not (layer2_outputs(2330));
    layer3_outputs(2694) <= (layer2_outputs(8950)) and (layer2_outputs(3196));
    layer3_outputs(2695) <= not(layer2_outputs(6956));
    layer3_outputs(2696) <= not(layer2_outputs(9550));
    layer3_outputs(2697) <= not(layer2_outputs(6068));
    layer3_outputs(2698) <= layer2_outputs(4764);
    layer3_outputs(2699) <= layer2_outputs(489);
    layer3_outputs(2700) <= not(layer2_outputs(3840));
    layer3_outputs(2701) <= not(layer2_outputs(856));
    layer3_outputs(2702) <= (layer2_outputs(807)) or (layer2_outputs(6384));
    layer3_outputs(2703) <= (layer2_outputs(8181)) and (layer2_outputs(423));
    layer3_outputs(2704) <= not((layer2_outputs(2127)) xor (layer2_outputs(3884)));
    layer3_outputs(2705) <= (layer2_outputs(8056)) or (layer2_outputs(1201));
    layer3_outputs(2706) <= not(layer2_outputs(77));
    layer3_outputs(2707) <= not(layer2_outputs(6765));
    layer3_outputs(2708) <= (layer2_outputs(7745)) and (layer2_outputs(5909));
    layer3_outputs(2709) <= layer2_outputs(2571);
    layer3_outputs(2710) <= layer2_outputs(1365);
    layer3_outputs(2711) <= not(layer2_outputs(2397));
    layer3_outputs(2712) <= layer2_outputs(1363);
    layer3_outputs(2713) <= layer2_outputs(2977);
    layer3_outputs(2714) <= not(layer2_outputs(8809));
    layer3_outputs(2715) <= layer2_outputs(6635);
    layer3_outputs(2716) <= not(layer2_outputs(6976)) or (layer2_outputs(8353));
    layer3_outputs(2717) <= (layer2_outputs(6185)) xor (layer2_outputs(7133));
    layer3_outputs(2718) <= not((layer2_outputs(6896)) or (layer2_outputs(4753)));
    layer3_outputs(2719) <= not(layer2_outputs(3645));
    layer3_outputs(2720) <= (layer2_outputs(4089)) and not (layer2_outputs(7729));
    layer3_outputs(2721) <= not(layer2_outputs(6662));
    layer3_outputs(2722) <= layer2_outputs(6163);
    layer3_outputs(2723) <= '0';
    layer3_outputs(2724) <= not((layer2_outputs(8659)) and (layer2_outputs(1630)));
    layer3_outputs(2725) <= not((layer2_outputs(6010)) and (layer2_outputs(6480)));
    layer3_outputs(2726) <= layer2_outputs(7298);
    layer3_outputs(2727) <= (layer2_outputs(1534)) and (layer2_outputs(7884));
    layer3_outputs(2728) <= layer2_outputs(10089);
    layer3_outputs(2729) <= (layer2_outputs(9811)) and not (layer2_outputs(4145));
    layer3_outputs(2730) <= layer2_outputs(6852);
    layer3_outputs(2731) <= not(layer2_outputs(4651));
    layer3_outputs(2732) <= layer2_outputs(8719);
    layer3_outputs(2733) <= not((layer2_outputs(8783)) or (layer2_outputs(9551)));
    layer3_outputs(2734) <= not((layer2_outputs(6643)) xor (layer2_outputs(5030)));
    layer3_outputs(2735) <= (layer2_outputs(5136)) or (layer2_outputs(1074));
    layer3_outputs(2736) <= not(layer2_outputs(6433));
    layer3_outputs(2737) <= (layer2_outputs(6381)) and not (layer2_outputs(4618));
    layer3_outputs(2738) <= layer2_outputs(3277);
    layer3_outputs(2739) <= '0';
    layer3_outputs(2740) <= layer2_outputs(10202);
    layer3_outputs(2741) <= '1';
    layer3_outputs(2742) <= not(layer2_outputs(6837));
    layer3_outputs(2743) <= (layer2_outputs(7621)) or (layer2_outputs(6524));
    layer3_outputs(2744) <= not((layer2_outputs(8071)) xor (layer2_outputs(7722)));
    layer3_outputs(2745) <= not(layer2_outputs(9842));
    layer3_outputs(2746) <= (layer2_outputs(6735)) xor (layer2_outputs(4127));
    layer3_outputs(2747) <= (layer2_outputs(2867)) or (layer2_outputs(1070));
    layer3_outputs(2748) <= (layer2_outputs(4404)) xor (layer2_outputs(2832));
    layer3_outputs(2749) <= (layer2_outputs(4842)) or (layer2_outputs(726));
    layer3_outputs(2750) <= not(layer2_outputs(4580));
    layer3_outputs(2751) <= not(layer2_outputs(5601));
    layer3_outputs(2752) <= not(layer2_outputs(4331)) or (layer2_outputs(2609));
    layer3_outputs(2753) <= not(layer2_outputs(554));
    layer3_outputs(2754) <= not(layer2_outputs(6839)) or (layer2_outputs(7485));
    layer3_outputs(2755) <= (layer2_outputs(7307)) xor (layer2_outputs(4173));
    layer3_outputs(2756) <= not(layer2_outputs(9171));
    layer3_outputs(2757) <= (layer2_outputs(865)) and not (layer2_outputs(4228));
    layer3_outputs(2758) <= not(layer2_outputs(1382));
    layer3_outputs(2759) <= not((layer2_outputs(3477)) or (layer2_outputs(8638)));
    layer3_outputs(2760) <= not(layer2_outputs(6824));
    layer3_outputs(2761) <= (layer2_outputs(9846)) xor (layer2_outputs(7868));
    layer3_outputs(2762) <= (layer2_outputs(984)) or (layer2_outputs(3691));
    layer3_outputs(2763) <= (layer2_outputs(2192)) and (layer2_outputs(2917));
    layer3_outputs(2764) <= (layer2_outputs(370)) and not (layer2_outputs(6624));
    layer3_outputs(2765) <= layer2_outputs(738);
    layer3_outputs(2766) <= not((layer2_outputs(3443)) xor (layer2_outputs(6899)));
    layer3_outputs(2767) <= '1';
    layer3_outputs(2768) <= not(layer2_outputs(1478));
    layer3_outputs(2769) <= not(layer2_outputs(2479));
    layer3_outputs(2770) <= not(layer2_outputs(343)) or (layer2_outputs(4139));
    layer3_outputs(2771) <= '0';
    layer3_outputs(2772) <= (layer2_outputs(3712)) or (layer2_outputs(1639));
    layer3_outputs(2773) <= not(layer2_outputs(8256));
    layer3_outputs(2774) <= (layer2_outputs(4591)) xor (layer2_outputs(304));
    layer3_outputs(2775) <= layer2_outputs(3949);
    layer3_outputs(2776) <= layer2_outputs(7651);
    layer3_outputs(2777) <= not(layer2_outputs(4099));
    layer3_outputs(2778) <= not(layer2_outputs(5594));
    layer3_outputs(2779) <= not(layer2_outputs(9717));
    layer3_outputs(2780) <= not(layer2_outputs(1494));
    layer3_outputs(2781) <= not(layer2_outputs(8551));
    layer3_outputs(2782) <= layer2_outputs(8284);
    layer3_outputs(2783) <= not((layer2_outputs(6569)) and (layer2_outputs(3291)));
    layer3_outputs(2784) <= layer2_outputs(2906);
    layer3_outputs(2785) <= not(layer2_outputs(4538));
    layer3_outputs(2786) <= layer2_outputs(6815);
    layer3_outputs(2787) <= (layer2_outputs(8094)) and not (layer2_outputs(2161));
    layer3_outputs(2788) <= not(layer2_outputs(8788));
    layer3_outputs(2789) <= not((layer2_outputs(2953)) xor (layer2_outputs(2997)));
    layer3_outputs(2790) <= '1';
    layer3_outputs(2791) <= '1';
    layer3_outputs(2792) <= (layer2_outputs(243)) xor (layer2_outputs(8516));
    layer3_outputs(2793) <= not(layer2_outputs(2562));
    layer3_outputs(2794) <= (layer2_outputs(1941)) and not (layer2_outputs(4334));
    layer3_outputs(2795) <= (layer2_outputs(3680)) and not (layer2_outputs(2893));
    layer3_outputs(2796) <= (layer2_outputs(3558)) and not (layer2_outputs(3745));
    layer3_outputs(2797) <= not(layer2_outputs(3035));
    layer3_outputs(2798) <= not(layer2_outputs(7682));
    layer3_outputs(2799) <= not(layer2_outputs(2102));
    layer3_outputs(2800) <= (layer2_outputs(3576)) and not (layer2_outputs(2073));
    layer3_outputs(2801) <= (layer2_outputs(3312)) xor (layer2_outputs(4370));
    layer3_outputs(2802) <= '1';
    layer3_outputs(2803) <= not(layer2_outputs(9803));
    layer3_outputs(2804) <= layer2_outputs(2892);
    layer3_outputs(2805) <= not((layer2_outputs(9821)) and (layer2_outputs(2647)));
    layer3_outputs(2806) <= layer2_outputs(7028);
    layer3_outputs(2807) <= not((layer2_outputs(4031)) or (layer2_outputs(9943)));
    layer3_outputs(2808) <= (layer2_outputs(1633)) xor (layer2_outputs(2794));
    layer3_outputs(2809) <= (layer2_outputs(22)) or (layer2_outputs(7063));
    layer3_outputs(2810) <= (layer2_outputs(4702)) and (layer2_outputs(8874));
    layer3_outputs(2811) <= layer2_outputs(9868);
    layer3_outputs(2812) <= layer2_outputs(2774);
    layer3_outputs(2813) <= '0';
    layer3_outputs(2814) <= (layer2_outputs(5363)) and not (layer2_outputs(585));
    layer3_outputs(2815) <= '1';
    layer3_outputs(2816) <= not(layer2_outputs(7328));
    layer3_outputs(2817) <= not((layer2_outputs(7356)) xor (layer2_outputs(1818)));
    layer3_outputs(2818) <= not(layer2_outputs(9738));
    layer3_outputs(2819) <= not(layer2_outputs(9937));
    layer3_outputs(2820) <= not(layer2_outputs(4584));
    layer3_outputs(2821) <= not(layer2_outputs(1667));
    layer3_outputs(2822) <= (layer2_outputs(9771)) and not (layer2_outputs(3657));
    layer3_outputs(2823) <= (layer2_outputs(7001)) and not (layer2_outputs(790));
    layer3_outputs(2824) <= (layer2_outputs(8818)) and (layer2_outputs(2152));
    layer3_outputs(2825) <= (layer2_outputs(4258)) and not (layer2_outputs(9353));
    layer3_outputs(2826) <= not(layer2_outputs(7856));
    layer3_outputs(2827) <= not(layer2_outputs(6230));
    layer3_outputs(2828) <= not(layer2_outputs(2690));
    layer3_outputs(2829) <= (layer2_outputs(8616)) and (layer2_outputs(480));
    layer3_outputs(2830) <= not(layer2_outputs(268));
    layer3_outputs(2831) <= (layer2_outputs(4791)) and (layer2_outputs(7937));
    layer3_outputs(2832) <= (layer2_outputs(1317)) or (layer2_outputs(1509));
    layer3_outputs(2833) <= layer2_outputs(1968);
    layer3_outputs(2834) <= not((layer2_outputs(8933)) or (layer2_outputs(2418)));
    layer3_outputs(2835) <= not(layer2_outputs(3160));
    layer3_outputs(2836) <= (layer2_outputs(9048)) and not (layer2_outputs(5108));
    layer3_outputs(2837) <= not((layer2_outputs(2796)) and (layer2_outputs(6170)));
    layer3_outputs(2838) <= not(layer2_outputs(3587));
    layer3_outputs(2839) <= layer2_outputs(9321);
    layer3_outputs(2840) <= layer2_outputs(9845);
    layer3_outputs(2841) <= layer2_outputs(9975);
    layer3_outputs(2842) <= not(layer2_outputs(4716)) or (layer2_outputs(4781));
    layer3_outputs(2843) <= not(layer2_outputs(7611));
    layer3_outputs(2844) <= not((layer2_outputs(6437)) xor (layer2_outputs(6231)));
    layer3_outputs(2845) <= layer2_outputs(7951);
    layer3_outputs(2846) <= not(layer2_outputs(7113)) or (layer2_outputs(5197));
    layer3_outputs(2847) <= layer2_outputs(3217);
    layer3_outputs(2848) <= not(layer2_outputs(5807));
    layer3_outputs(2849) <= not((layer2_outputs(9707)) xor (layer2_outputs(6764)));
    layer3_outputs(2850) <= not(layer2_outputs(7129));
    layer3_outputs(2851) <= (layer2_outputs(1335)) or (layer2_outputs(7483));
    layer3_outputs(2852) <= layer2_outputs(9648);
    layer3_outputs(2853) <= layer2_outputs(2836);
    layer3_outputs(2854) <= (layer2_outputs(3794)) or (layer2_outputs(8503));
    layer3_outputs(2855) <= not(layer2_outputs(8164));
    layer3_outputs(2856) <= layer2_outputs(777);
    layer3_outputs(2857) <= (layer2_outputs(3643)) xor (layer2_outputs(2928));
    layer3_outputs(2858) <= (layer2_outputs(7135)) and not (layer2_outputs(8491));
    layer3_outputs(2859) <= layer2_outputs(2593);
    layer3_outputs(2860) <= layer2_outputs(3604);
    layer3_outputs(2861) <= '0';
    layer3_outputs(2862) <= (layer2_outputs(4248)) and not (layer2_outputs(9583));
    layer3_outputs(2863) <= not((layer2_outputs(8088)) or (layer2_outputs(4295)));
    layer3_outputs(2864) <= layer2_outputs(1518);
    layer3_outputs(2865) <= (layer2_outputs(6815)) and not (layer2_outputs(8172));
    layer3_outputs(2866) <= not((layer2_outputs(2122)) xor (layer2_outputs(8178)));
    layer3_outputs(2867) <= layer2_outputs(74);
    layer3_outputs(2868) <= not((layer2_outputs(2599)) and (layer2_outputs(8610)));
    layer3_outputs(2869) <= not((layer2_outputs(1527)) xor (layer2_outputs(802)));
    layer3_outputs(2870) <= not(layer2_outputs(1899));
    layer3_outputs(2871) <= layer2_outputs(9242);
    layer3_outputs(2872) <= '0';
    layer3_outputs(2873) <= (layer2_outputs(1052)) and not (layer2_outputs(1616));
    layer3_outputs(2874) <= not(layer2_outputs(6997));
    layer3_outputs(2875) <= (layer2_outputs(4384)) or (layer2_outputs(10113));
    layer3_outputs(2876) <= not(layer2_outputs(9586));
    layer3_outputs(2877) <= '1';
    layer3_outputs(2878) <= layer2_outputs(6222);
    layer3_outputs(2879) <= layer2_outputs(2683);
    layer3_outputs(2880) <= not(layer2_outputs(2545));
    layer3_outputs(2881) <= not(layer2_outputs(5490));
    layer3_outputs(2882) <= not(layer2_outputs(6787));
    layer3_outputs(2883) <= (layer2_outputs(7918)) and not (layer2_outputs(5862));
    layer3_outputs(2884) <= not(layer2_outputs(8229));
    layer3_outputs(2885) <= layer2_outputs(4067);
    layer3_outputs(2886) <= not(layer2_outputs(6980));
    layer3_outputs(2887) <= not(layer2_outputs(2800));
    layer3_outputs(2888) <= layer2_outputs(1800);
    layer3_outputs(2889) <= (layer2_outputs(2133)) xor (layer2_outputs(6602));
    layer3_outputs(2890) <= (layer2_outputs(5926)) and not (layer2_outputs(7809));
    layer3_outputs(2891) <= not((layer2_outputs(2270)) and (layer2_outputs(9367)));
    layer3_outputs(2892) <= not(layer2_outputs(31)) or (layer2_outputs(7176));
    layer3_outputs(2893) <= '1';
    layer3_outputs(2894) <= layer2_outputs(345);
    layer3_outputs(2895) <= not(layer2_outputs(550)) or (layer2_outputs(8375));
    layer3_outputs(2896) <= layer2_outputs(7452);
    layer3_outputs(2897) <= (layer2_outputs(2038)) or (layer2_outputs(6439));
    layer3_outputs(2898) <= not(layer2_outputs(6817));
    layer3_outputs(2899) <= layer2_outputs(3433);
    layer3_outputs(2900) <= layer2_outputs(9987);
    layer3_outputs(2901) <= not(layer2_outputs(2453));
    layer3_outputs(2902) <= not(layer2_outputs(1618));
    layer3_outputs(2903) <= not(layer2_outputs(3017)) or (layer2_outputs(1499));
    layer3_outputs(2904) <= not(layer2_outputs(5809));
    layer3_outputs(2905) <= not(layer2_outputs(8128));
    layer3_outputs(2906) <= not(layer2_outputs(7436));
    layer3_outputs(2907) <= not(layer2_outputs(10085));
    layer3_outputs(2908) <= not(layer2_outputs(10235)) or (layer2_outputs(5139));
    layer3_outputs(2909) <= layer2_outputs(2571);
    layer3_outputs(2910) <= layer2_outputs(3731);
    layer3_outputs(2911) <= (layer2_outputs(969)) or (layer2_outputs(6083));
    layer3_outputs(2912) <= not(layer2_outputs(9494));
    layer3_outputs(2913) <= (layer2_outputs(7257)) and not (layer2_outputs(303));
    layer3_outputs(2914) <= not(layer2_outputs(4661)) or (layer2_outputs(5652));
    layer3_outputs(2915) <= (layer2_outputs(7086)) and not (layer2_outputs(1966));
    layer3_outputs(2916) <= not((layer2_outputs(2531)) or (layer2_outputs(4984)));
    layer3_outputs(2917) <= layer2_outputs(7742);
    layer3_outputs(2918) <= layer2_outputs(5337);
    layer3_outputs(2919) <= layer2_outputs(2589);
    layer3_outputs(2920) <= not((layer2_outputs(1205)) and (layer2_outputs(2070)));
    layer3_outputs(2921) <= not(layer2_outputs(198)) or (layer2_outputs(5585));
    layer3_outputs(2922) <= not(layer2_outputs(3955));
    layer3_outputs(2923) <= (layer2_outputs(2032)) and not (layer2_outputs(7724));
    layer3_outputs(2924) <= not(layer2_outputs(9521));
    layer3_outputs(2925) <= (layer2_outputs(239)) and not (layer2_outputs(561));
    layer3_outputs(2926) <= layer2_outputs(7159);
    layer3_outputs(2927) <= layer2_outputs(7782);
    layer3_outputs(2928) <= layer2_outputs(2588);
    layer3_outputs(2929) <= not(layer2_outputs(3905));
    layer3_outputs(2930) <= layer2_outputs(4159);
    layer3_outputs(2931) <= (layer2_outputs(7835)) xor (layer2_outputs(10233));
    layer3_outputs(2932) <= '1';
    layer3_outputs(2933) <= not(layer2_outputs(4255));
    layer3_outputs(2934) <= not((layer2_outputs(6803)) and (layer2_outputs(3822)));
    layer3_outputs(2935) <= not(layer2_outputs(2353));
    layer3_outputs(2936) <= not(layer2_outputs(8635));
    layer3_outputs(2937) <= layer2_outputs(9519);
    layer3_outputs(2938) <= not(layer2_outputs(6335));
    layer3_outputs(2939) <= not((layer2_outputs(6880)) xor (layer2_outputs(10002)));
    layer3_outputs(2940) <= layer2_outputs(9852);
    layer3_outputs(2941) <= layer2_outputs(10212);
    layer3_outputs(2942) <= not(layer2_outputs(2264));
    layer3_outputs(2943) <= (layer2_outputs(2471)) or (layer2_outputs(8494));
    layer3_outputs(2944) <= layer2_outputs(6688);
    layer3_outputs(2945) <= not(layer2_outputs(380)) or (layer2_outputs(5692));
    layer3_outputs(2946) <= not(layer2_outputs(1887));
    layer3_outputs(2947) <= (layer2_outputs(3105)) and not (layer2_outputs(621));
    layer3_outputs(2948) <= '1';
    layer3_outputs(2949) <= not(layer2_outputs(626));
    layer3_outputs(2950) <= '0';
    layer3_outputs(2951) <= layer2_outputs(743);
    layer3_outputs(2952) <= (layer2_outputs(7309)) and not (layer2_outputs(5535));
    layer3_outputs(2953) <= not((layer2_outputs(1068)) and (layer2_outputs(3254)));
    layer3_outputs(2954) <= layer2_outputs(1355);
    layer3_outputs(2955) <= (layer2_outputs(135)) xor (layer2_outputs(7704));
    layer3_outputs(2956) <= not((layer2_outputs(7569)) xor (layer2_outputs(9342)));
    layer3_outputs(2957) <= layer2_outputs(3574);
    layer3_outputs(2958) <= (layer2_outputs(4401)) xor (layer2_outputs(5377));
    layer3_outputs(2959) <= '0';
    layer3_outputs(2960) <= not(layer2_outputs(9983));
    layer3_outputs(2961) <= (layer2_outputs(7256)) and (layer2_outputs(542));
    layer3_outputs(2962) <= not((layer2_outputs(4694)) and (layer2_outputs(2131)));
    layer3_outputs(2963) <= layer2_outputs(5747);
    layer3_outputs(2964) <= not((layer2_outputs(9065)) and (layer2_outputs(1690)));
    layer3_outputs(2965) <= layer2_outputs(48);
    layer3_outputs(2966) <= not(layer2_outputs(1674)) or (layer2_outputs(4080));
    layer3_outputs(2967) <= (layer2_outputs(198)) and not (layer2_outputs(6070));
    layer3_outputs(2968) <= layer2_outputs(4809);
    layer3_outputs(2969) <= (layer2_outputs(548)) and not (layer2_outputs(7282));
    layer3_outputs(2970) <= layer2_outputs(7559);
    layer3_outputs(2971) <= not(layer2_outputs(10158));
    layer3_outputs(2972) <= (layer2_outputs(1848)) or (layer2_outputs(2025));
    layer3_outputs(2973) <= (layer2_outputs(2298)) xor (layer2_outputs(4631));
    layer3_outputs(2974) <= layer2_outputs(9371);
    layer3_outputs(2975) <= layer2_outputs(5208);
    layer3_outputs(2976) <= (layer2_outputs(2637)) and not (layer2_outputs(2218));
    layer3_outputs(2977) <= not(layer2_outputs(9526));
    layer3_outputs(2978) <= not(layer2_outputs(2944));
    layer3_outputs(2979) <= not((layer2_outputs(2203)) and (layer2_outputs(4931)));
    layer3_outputs(2980) <= not(layer2_outputs(10174)) or (layer2_outputs(6304));
    layer3_outputs(2981) <= (layer2_outputs(6070)) and not (layer2_outputs(10084));
    layer3_outputs(2982) <= (layer2_outputs(2689)) and (layer2_outputs(10236));
    layer3_outputs(2983) <= not((layer2_outputs(6521)) and (layer2_outputs(8807)));
    layer3_outputs(2984) <= '0';
    layer3_outputs(2985) <= not(layer2_outputs(3103));
    layer3_outputs(2986) <= layer2_outputs(2097);
    layer3_outputs(2987) <= layer2_outputs(5785);
    layer3_outputs(2988) <= not((layer2_outputs(1094)) or (layer2_outputs(5896)));
    layer3_outputs(2989) <= not((layer2_outputs(4042)) or (layer2_outputs(8675)));
    layer3_outputs(2990) <= layer2_outputs(4681);
    layer3_outputs(2991) <= not(layer2_outputs(8088));
    layer3_outputs(2992) <= not(layer2_outputs(9725)) or (layer2_outputs(2461));
    layer3_outputs(2993) <= not((layer2_outputs(2291)) xor (layer2_outputs(3098)));
    layer3_outputs(2994) <= (layer2_outputs(3076)) and not (layer2_outputs(5023));
    layer3_outputs(2995) <= layer2_outputs(6081);
    layer3_outputs(2996) <= not((layer2_outputs(9425)) and (layer2_outputs(3264)));
    layer3_outputs(2997) <= layer2_outputs(1535);
    layer3_outputs(2998) <= not(layer2_outputs(7397));
    layer3_outputs(2999) <= not(layer2_outputs(8306));
    layer3_outputs(3000) <= '1';
    layer3_outputs(3001) <= not(layer2_outputs(2045));
    layer3_outputs(3002) <= (layer2_outputs(3985)) and not (layer2_outputs(7998));
    layer3_outputs(3003) <= '1';
    layer3_outputs(3004) <= not(layer2_outputs(1837));
    layer3_outputs(3005) <= (layer2_outputs(7333)) or (layer2_outputs(2178));
    layer3_outputs(3006) <= not(layer2_outputs(2891));
    layer3_outputs(3007) <= not(layer2_outputs(5297));
    layer3_outputs(3008) <= not((layer2_outputs(7829)) and (layer2_outputs(8154)));
    layer3_outputs(3009) <= layer2_outputs(4147);
    layer3_outputs(3010) <= not(layer2_outputs(4502));
    layer3_outputs(3011) <= not(layer2_outputs(1221)) or (layer2_outputs(6913));
    layer3_outputs(3012) <= layer2_outputs(2249);
    layer3_outputs(3013) <= not(layer2_outputs(1799)) or (layer2_outputs(9397));
    layer3_outputs(3014) <= not((layer2_outputs(8882)) or (layer2_outputs(5540)));
    layer3_outputs(3015) <= not(layer2_outputs(450)) or (layer2_outputs(9418));
    layer3_outputs(3016) <= not(layer2_outputs(7575));
    layer3_outputs(3017) <= not(layer2_outputs(3197));
    layer3_outputs(3018) <= layer2_outputs(883);
    layer3_outputs(3019) <= not(layer2_outputs(4689));
    layer3_outputs(3020) <= not(layer2_outputs(9448));
    layer3_outputs(3021) <= not(layer2_outputs(1178));
    layer3_outputs(3022) <= layer2_outputs(6150);
    layer3_outputs(3023) <= not(layer2_outputs(8766));
    layer3_outputs(3024) <= not((layer2_outputs(8588)) or (layer2_outputs(6123)));
    layer3_outputs(3025) <= not((layer2_outputs(5019)) and (layer2_outputs(9609)));
    layer3_outputs(3026) <= '1';
    layer3_outputs(3027) <= (layer2_outputs(8405)) xor (layer2_outputs(7655));
    layer3_outputs(3028) <= not((layer2_outputs(2877)) xor (layer2_outputs(27)));
    layer3_outputs(3029) <= (layer2_outputs(9753)) and (layer2_outputs(8002));
    layer3_outputs(3030) <= not(layer2_outputs(8216));
    layer3_outputs(3031) <= layer2_outputs(1888);
    layer3_outputs(3032) <= (layer2_outputs(6144)) and (layer2_outputs(2447));
    layer3_outputs(3033) <= not((layer2_outputs(3160)) and (layer2_outputs(4653)));
    layer3_outputs(3034) <= not(layer2_outputs(1531)) or (layer2_outputs(4060));
    layer3_outputs(3035) <= layer2_outputs(1582);
    layer3_outputs(3036) <= layer2_outputs(2927);
    layer3_outputs(3037) <= (layer2_outputs(1203)) and not (layer2_outputs(6317));
    layer3_outputs(3038) <= (layer2_outputs(9504)) and not (layer2_outputs(9702));
    layer3_outputs(3039) <= not(layer2_outputs(10101));
    layer3_outputs(3040) <= (layer2_outputs(9414)) and not (layer2_outputs(1232));
    layer3_outputs(3041) <= not(layer2_outputs(4555)) or (layer2_outputs(2679));
    layer3_outputs(3042) <= layer2_outputs(5085);
    layer3_outputs(3043) <= (layer2_outputs(4606)) and not (layer2_outputs(620));
    layer3_outputs(3044) <= layer2_outputs(5805);
    layer3_outputs(3045) <= (layer2_outputs(7)) and not (layer2_outputs(9630));
    layer3_outputs(3046) <= (layer2_outputs(9962)) and (layer2_outputs(7593));
    layer3_outputs(3047) <= layer2_outputs(7503);
    layer3_outputs(3048) <= (layer2_outputs(471)) and not (layer2_outputs(2138));
    layer3_outputs(3049) <= not(layer2_outputs(357));
    layer3_outputs(3050) <= not(layer2_outputs(522));
    layer3_outputs(3051) <= (layer2_outputs(5863)) and not (layer2_outputs(2191));
    layer3_outputs(3052) <= (layer2_outputs(6653)) xor (layer2_outputs(6282));
    layer3_outputs(3053) <= layer2_outputs(5209);
    layer3_outputs(3054) <= layer2_outputs(1979);
    layer3_outputs(3055) <= not((layer2_outputs(7441)) xor (layer2_outputs(7189)));
    layer3_outputs(3056) <= layer2_outputs(8020);
    layer3_outputs(3057) <= not((layer2_outputs(9963)) and (layer2_outputs(9789)));
    layer3_outputs(3058) <= layer2_outputs(3025);
    layer3_outputs(3059) <= (layer2_outputs(2762)) and not (layer2_outputs(790));
    layer3_outputs(3060) <= not((layer2_outputs(8751)) xor (layer2_outputs(3043)));
    layer3_outputs(3061) <= (layer2_outputs(2849)) and not (layer2_outputs(8974));
    layer3_outputs(3062) <= not(layer2_outputs(770)) or (layer2_outputs(1753));
    layer3_outputs(3063) <= not(layer2_outputs(7778));
    layer3_outputs(3064) <= not(layer2_outputs(4649));
    layer3_outputs(3065) <= not(layer2_outputs(6538));
    layer3_outputs(3066) <= (layer2_outputs(8593)) or (layer2_outputs(10217));
    layer3_outputs(3067) <= layer2_outputs(9843);
    layer3_outputs(3068) <= layer2_outputs(8427);
    layer3_outputs(3069) <= not(layer2_outputs(6730));
    layer3_outputs(3070) <= not((layer2_outputs(1460)) or (layer2_outputs(9802)));
    layer3_outputs(3071) <= not(layer2_outputs(1002));
    layer3_outputs(3072) <= (layer2_outputs(7797)) or (layer2_outputs(3190));
    layer3_outputs(3073) <= (layer2_outputs(2664)) and not (layer2_outputs(6));
    layer3_outputs(3074) <= layer2_outputs(9290);
    layer3_outputs(3075) <= (layer2_outputs(7928)) or (layer2_outputs(7492));
    layer3_outputs(3076) <= layer2_outputs(814);
    layer3_outputs(3077) <= not((layer2_outputs(3772)) and (layer2_outputs(6814)));
    layer3_outputs(3078) <= (layer2_outputs(44)) xor (layer2_outputs(10216));
    layer3_outputs(3079) <= not(layer2_outputs(344));
    layer3_outputs(3080) <= not(layer2_outputs(9002));
    layer3_outputs(3081) <= not(layer2_outputs(9989));
    layer3_outputs(3082) <= '0';
    layer3_outputs(3083) <= '0';
    layer3_outputs(3084) <= (layer2_outputs(3749)) and not (layer2_outputs(1876));
    layer3_outputs(3085) <= not(layer2_outputs(4488)) or (layer2_outputs(4601));
    layer3_outputs(3086) <= (layer2_outputs(7997)) or (layer2_outputs(3094));
    layer3_outputs(3087) <= (layer2_outputs(8318)) and (layer2_outputs(9439));
    layer3_outputs(3088) <= not(layer2_outputs(7124));
    layer3_outputs(3089) <= layer2_outputs(9003);
    layer3_outputs(3090) <= layer2_outputs(8957);
    layer3_outputs(3091) <= not(layer2_outputs(3586));
    layer3_outputs(3092) <= not(layer2_outputs(1785));
    layer3_outputs(3093) <= layer2_outputs(5564);
    layer3_outputs(3094) <= not(layer2_outputs(9009));
    layer3_outputs(3095) <= not((layer2_outputs(9599)) xor (layer2_outputs(9823)));
    layer3_outputs(3096) <= not(layer2_outputs(3199));
    layer3_outputs(3097) <= not(layer2_outputs(410)) or (layer2_outputs(4357));
    layer3_outputs(3098) <= layer2_outputs(1646);
    layer3_outputs(3099) <= not(layer2_outputs(9337));
    layer3_outputs(3100) <= layer2_outputs(9496);
    layer3_outputs(3101) <= not((layer2_outputs(6930)) or (layer2_outputs(1083)));
    layer3_outputs(3102) <= layer2_outputs(381);
    layer3_outputs(3103) <= (layer2_outputs(6237)) xor (layer2_outputs(3513));
    layer3_outputs(3104) <= (layer2_outputs(4061)) xor (layer2_outputs(8483));
    layer3_outputs(3105) <= not(layer2_outputs(6272)) or (layer2_outputs(2336));
    layer3_outputs(3106) <= not((layer2_outputs(2221)) or (layer2_outputs(2302)));
    layer3_outputs(3107) <= not(layer2_outputs(9096));
    layer3_outputs(3108) <= '0';
    layer3_outputs(3109) <= layer2_outputs(3187);
    layer3_outputs(3110) <= layer2_outputs(5792);
    layer3_outputs(3111) <= (layer2_outputs(1944)) and (layer2_outputs(4321));
    layer3_outputs(3112) <= layer2_outputs(4574);
    layer3_outputs(3113) <= not(layer2_outputs(2130));
    layer3_outputs(3114) <= (layer2_outputs(4382)) and not (layer2_outputs(9813));
    layer3_outputs(3115) <= (layer2_outputs(8425)) xor (layer2_outputs(3937));
    layer3_outputs(3116) <= not(layer2_outputs(279));
    layer3_outputs(3117) <= layer2_outputs(4987);
    layer3_outputs(3118) <= not(layer2_outputs(3517));
    layer3_outputs(3119) <= layer2_outputs(6333);
    layer3_outputs(3120) <= layer2_outputs(8015);
    layer3_outputs(3121) <= not(layer2_outputs(4825)) or (layer2_outputs(6200));
    layer3_outputs(3122) <= not(layer2_outputs(3093)) or (layer2_outputs(855));
    layer3_outputs(3123) <= not(layer2_outputs(615));
    layer3_outputs(3124) <= layer2_outputs(1098);
    layer3_outputs(3125) <= not(layer2_outputs(2235));
    layer3_outputs(3126) <= layer2_outputs(2650);
    layer3_outputs(3127) <= not((layer2_outputs(10194)) and (layer2_outputs(8846)));
    layer3_outputs(3128) <= layer2_outputs(2830);
    layer3_outputs(3129) <= layer2_outputs(6550);
    layer3_outputs(3130) <= not(layer2_outputs(5343));
    layer3_outputs(3131) <= '0';
    layer3_outputs(3132) <= not(layer2_outputs(5710));
    layer3_outputs(3133) <= not(layer2_outputs(7673));
    layer3_outputs(3134) <= (layer2_outputs(117)) or (layer2_outputs(1787));
    layer3_outputs(3135) <= not(layer2_outputs(1596)) or (layer2_outputs(7108));
    layer3_outputs(3136) <= not(layer2_outputs(10117));
    layer3_outputs(3137) <= (layer2_outputs(7695)) and (layer2_outputs(5192));
    layer3_outputs(3138) <= not((layer2_outputs(3441)) xor (layer2_outputs(8672)));
    layer3_outputs(3139) <= not((layer2_outputs(8062)) or (layer2_outputs(8408)));
    layer3_outputs(3140) <= not(layer2_outputs(7480));
    layer3_outputs(3141) <= (layer2_outputs(9499)) and not (layer2_outputs(1557));
    layer3_outputs(3142) <= not(layer2_outputs(7082)) or (layer2_outputs(7450));
    layer3_outputs(3143) <= not(layer2_outputs(1545));
    layer3_outputs(3144) <= not((layer2_outputs(635)) or (layer2_outputs(5629)));
    layer3_outputs(3145) <= not((layer2_outputs(260)) or (layer2_outputs(2409)));
    layer3_outputs(3146) <= (layer2_outputs(2580)) and (layer2_outputs(5997));
    layer3_outputs(3147) <= not(layer2_outputs(8710)) or (layer2_outputs(1082));
    layer3_outputs(3148) <= not(layer2_outputs(7973));
    layer3_outputs(3149) <= layer2_outputs(9631);
    layer3_outputs(3150) <= (layer2_outputs(2138)) and (layer2_outputs(26));
    layer3_outputs(3151) <= (layer2_outputs(9175)) xor (layer2_outputs(3576));
    layer3_outputs(3152) <= not(layer2_outputs(9059)) or (layer2_outputs(8091));
    layer3_outputs(3153) <= layer2_outputs(5333);
    layer3_outputs(3154) <= (layer2_outputs(1931)) xor (layer2_outputs(4399));
    layer3_outputs(3155) <= layer2_outputs(4256);
    layer3_outputs(3156) <= (layer2_outputs(9727)) and not (layer2_outputs(1605));
    layer3_outputs(3157) <= not((layer2_outputs(4137)) xor (layer2_outputs(4588)));
    layer3_outputs(3158) <= layer2_outputs(4729);
    layer3_outputs(3159) <= (layer2_outputs(4536)) xor (layer2_outputs(5574));
    layer3_outputs(3160) <= layer2_outputs(6248);
    layer3_outputs(3161) <= layer2_outputs(5614);
    layer3_outputs(3162) <= layer2_outputs(9038);
    layer3_outputs(3163) <= not(layer2_outputs(2511));
    layer3_outputs(3164) <= not((layer2_outputs(7478)) and (layer2_outputs(3198)));
    layer3_outputs(3165) <= (layer2_outputs(2851)) xor (layer2_outputs(6093));
    layer3_outputs(3166) <= (layer2_outputs(975)) and not (layer2_outputs(4488));
    layer3_outputs(3167) <= not(layer2_outputs(6495)) or (layer2_outputs(6282));
    layer3_outputs(3168) <= not(layer2_outputs(8431));
    layer3_outputs(3169) <= not((layer2_outputs(3425)) xor (layer2_outputs(2505)));
    layer3_outputs(3170) <= not(layer2_outputs(6805));
    layer3_outputs(3171) <= (layer2_outputs(4479)) or (layer2_outputs(65));
    layer3_outputs(3172) <= (layer2_outputs(1506)) and (layer2_outputs(8646));
    layer3_outputs(3173) <= '0';
    layer3_outputs(3174) <= not(layer2_outputs(1167));
    layer3_outputs(3175) <= not(layer2_outputs(3601));
    layer3_outputs(3176) <= '0';
    layer3_outputs(3177) <= not((layer2_outputs(4827)) and (layer2_outputs(249)));
    layer3_outputs(3178) <= not(layer2_outputs(5195));
    layer3_outputs(3179) <= (layer2_outputs(3768)) and not (layer2_outputs(1249));
    layer3_outputs(3180) <= not(layer2_outputs(8960));
    layer3_outputs(3181) <= (layer2_outputs(1780)) and (layer2_outputs(9474));
    layer3_outputs(3182) <= layer2_outputs(5073);
    layer3_outputs(3183) <= layer2_outputs(7243);
    layer3_outputs(3184) <= not(layer2_outputs(9388));
    layer3_outputs(3185) <= layer2_outputs(8472);
    layer3_outputs(3186) <= '0';
    layer3_outputs(3187) <= layer2_outputs(8135);
    layer3_outputs(3188) <= (layer2_outputs(7161)) and (layer2_outputs(9700));
    layer3_outputs(3189) <= (layer2_outputs(8430)) and not (layer2_outputs(7925));
    layer3_outputs(3190) <= (layer2_outputs(3638)) xor (layer2_outputs(3449));
    layer3_outputs(3191) <= not(layer2_outputs(4209)) or (layer2_outputs(6251));
    layer3_outputs(3192) <= not((layer2_outputs(2786)) xor (layer2_outputs(5272)));
    layer3_outputs(3193) <= not((layer2_outputs(8606)) and (layer2_outputs(5113)));
    layer3_outputs(3194) <= layer2_outputs(2335);
    layer3_outputs(3195) <= (layer2_outputs(4720)) xor (layer2_outputs(545));
    layer3_outputs(3196) <= not(layer2_outputs(3010));
    layer3_outputs(3197) <= layer2_outputs(6160);
    layer3_outputs(3198) <= (layer2_outputs(1167)) xor (layer2_outputs(8391));
    layer3_outputs(3199) <= layer2_outputs(3092);
    layer3_outputs(3200) <= not((layer2_outputs(9193)) xor (layer2_outputs(8382)));
    layer3_outputs(3201) <= not(layer2_outputs(3839));
    layer3_outputs(3202) <= layer2_outputs(3903);
    layer3_outputs(3203) <= layer2_outputs(673);
    layer3_outputs(3204) <= not(layer2_outputs(1855));
    layer3_outputs(3205) <= not(layer2_outputs(7468));
    layer3_outputs(3206) <= layer2_outputs(3463);
    layer3_outputs(3207) <= layer2_outputs(3179);
    layer3_outputs(3208) <= (layer2_outputs(3168)) or (layer2_outputs(7919));
    layer3_outputs(3209) <= layer2_outputs(3315);
    layer3_outputs(3210) <= not((layer2_outputs(2248)) xor (layer2_outputs(3293)));
    layer3_outputs(3211) <= (layer2_outputs(8344)) or (layer2_outputs(9899));
    layer3_outputs(3212) <= layer2_outputs(6173);
    layer3_outputs(3213) <= not(layer2_outputs(6078));
    layer3_outputs(3214) <= not(layer2_outputs(8572)) or (layer2_outputs(2555));
    layer3_outputs(3215) <= layer2_outputs(4053);
    layer3_outputs(3216) <= (layer2_outputs(1851)) and not (layer2_outputs(5708));
    layer3_outputs(3217) <= layer2_outputs(7094);
    layer3_outputs(3218) <= not(layer2_outputs(9141)) or (layer2_outputs(5144));
    layer3_outputs(3219) <= (layer2_outputs(1814)) xor (layer2_outputs(1584));
    layer3_outputs(3220) <= '0';
    layer3_outputs(3221) <= not((layer2_outputs(10033)) and (layer2_outputs(5891)));
    layer3_outputs(3222) <= layer2_outputs(9722);
    layer3_outputs(3223) <= not((layer2_outputs(7130)) and (layer2_outputs(186)));
    layer3_outputs(3224) <= not(layer2_outputs(9222)) or (layer2_outputs(8986));
    layer3_outputs(3225) <= (layer2_outputs(3961)) or (layer2_outputs(7116));
    layer3_outputs(3226) <= not((layer2_outputs(7620)) xor (layer2_outputs(6520)));
    layer3_outputs(3227) <= not(layer2_outputs(9622));
    layer3_outputs(3228) <= layer2_outputs(2058);
    layer3_outputs(3229) <= (layer2_outputs(3736)) and not (layer2_outputs(223));
    layer3_outputs(3230) <= (layer2_outputs(832)) xor (layer2_outputs(6489));
    layer3_outputs(3231) <= layer2_outputs(2667);
    layer3_outputs(3232) <= layer2_outputs(2451);
    layer3_outputs(3233) <= (layer2_outputs(1748)) and not (layer2_outputs(2902));
    layer3_outputs(3234) <= not(layer2_outputs(8392));
    layer3_outputs(3235) <= not(layer2_outputs(6197));
    layer3_outputs(3236) <= not(layer2_outputs(6480));
    layer3_outputs(3237) <= not(layer2_outputs(7046));
    layer3_outputs(3238) <= not(layer2_outputs(1292));
    layer3_outputs(3239) <= layer2_outputs(2171);
    layer3_outputs(3240) <= not((layer2_outputs(8632)) xor (layer2_outputs(8538)));
    layer3_outputs(3241) <= not((layer2_outputs(9988)) xor (layer2_outputs(8186)));
    layer3_outputs(3242) <= not(layer2_outputs(5294)) or (layer2_outputs(1260));
    layer3_outputs(3243) <= not(layer2_outputs(347));
    layer3_outputs(3244) <= '0';
    layer3_outputs(3245) <= not(layer2_outputs(6470));
    layer3_outputs(3246) <= not((layer2_outputs(3010)) and (layer2_outputs(6871)));
    layer3_outputs(3247) <= not((layer2_outputs(10188)) or (layer2_outputs(5115)));
    layer3_outputs(3248) <= layer2_outputs(8737);
    layer3_outputs(3249) <= not(layer2_outputs(2093));
    layer3_outputs(3250) <= layer2_outputs(4337);
    layer3_outputs(3251) <= not(layer2_outputs(7022));
    layer3_outputs(3252) <= (layer2_outputs(4430)) xor (layer2_outputs(1233));
    layer3_outputs(3253) <= not(layer2_outputs(7169));
    layer3_outputs(3254) <= not(layer2_outputs(373));
    layer3_outputs(3255) <= not((layer2_outputs(1406)) and (layer2_outputs(6695)));
    layer3_outputs(3256) <= layer2_outputs(9035);
    layer3_outputs(3257) <= (layer2_outputs(8800)) and not (layer2_outputs(3162));
    layer3_outputs(3258) <= not(layer2_outputs(1587)) or (layer2_outputs(8682));
    layer3_outputs(3259) <= not(layer2_outputs(8693));
    layer3_outputs(3260) <= not(layer2_outputs(8927));
    layer3_outputs(3261) <= not(layer2_outputs(5261));
    layer3_outputs(3262) <= layer2_outputs(746);
    layer3_outputs(3263) <= not(layer2_outputs(7898));
    layer3_outputs(3264) <= not(layer2_outputs(4101)) or (layer2_outputs(8941));
    layer3_outputs(3265) <= not((layer2_outputs(4980)) and (layer2_outputs(3218)));
    layer3_outputs(3266) <= layer2_outputs(3849);
    layer3_outputs(3267) <= (layer2_outputs(6586)) xor (layer2_outputs(3180));
    layer3_outputs(3268) <= layer2_outputs(2964);
    layer3_outputs(3269) <= not(layer2_outputs(1910));
    layer3_outputs(3270) <= not(layer2_outputs(9585));
    layer3_outputs(3271) <= layer2_outputs(3149);
    layer3_outputs(3272) <= '1';
    layer3_outputs(3273) <= (layer2_outputs(610)) and (layer2_outputs(3441));
    layer3_outputs(3274) <= (layer2_outputs(5051)) and not (layer2_outputs(7617));
    layer3_outputs(3275) <= not(layer2_outputs(6791)) or (layer2_outputs(3498));
    layer3_outputs(3276) <= layer2_outputs(715);
    layer3_outputs(3277) <= '1';
    layer3_outputs(3278) <= '1';
    layer3_outputs(3279) <= not(layer2_outputs(2527));
    layer3_outputs(3280) <= not(layer2_outputs(2304));
    layer3_outputs(3281) <= (layer2_outputs(6533)) and not (layer2_outputs(5427));
    layer3_outputs(3282) <= (layer2_outputs(3464)) or (layer2_outputs(6915));
    layer3_outputs(3283) <= not(layer2_outputs(10134));
    layer3_outputs(3284) <= not(layer2_outputs(4930));
    layer3_outputs(3285) <= (layer2_outputs(2044)) and not (layer2_outputs(9120));
    layer3_outputs(3286) <= not(layer2_outputs(7521));
    layer3_outputs(3287) <= not(layer2_outputs(5288));
    layer3_outputs(3288) <= (layer2_outputs(3486)) and not (layer2_outputs(8679));
    layer3_outputs(3289) <= not((layer2_outputs(659)) xor (layer2_outputs(10160)));
    layer3_outputs(3290) <= not(layer2_outputs(6162)) or (layer2_outputs(9450));
    layer3_outputs(3291) <= not(layer2_outputs(10191));
    layer3_outputs(3292) <= layer2_outputs(1662);
    layer3_outputs(3293) <= layer2_outputs(9924);
    layer3_outputs(3294) <= not((layer2_outputs(7310)) xor (layer2_outputs(5653)));
    layer3_outputs(3295) <= (layer2_outputs(7392)) and (layer2_outputs(5576));
    layer3_outputs(3296) <= layer2_outputs(1276);
    layer3_outputs(3297) <= not(layer2_outputs(1257));
    layer3_outputs(3298) <= layer2_outputs(5573);
    layer3_outputs(3299) <= layer2_outputs(2386);
    layer3_outputs(3300) <= (layer2_outputs(8127)) or (layer2_outputs(5168));
    layer3_outputs(3301) <= layer2_outputs(7404);
    layer3_outputs(3302) <= layer2_outputs(3799);
    layer3_outputs(3303) <= layer2_outputs(8559);
    layer3_outputs(3304) <= not(layer2_outputs(2154));
    layer3_outputs(3305) <= layer2_outputs(6283);
    layer3_outputs(3306) <= layer2_outputs(2592);
    layer3_outputs(3307) <= not((layer2_outputs(120)) or (layer2_outputs(4163)));
    layer3_outputs(3308) <= not(layer2_outputs(699)) or (layer2_outputs(3635));
    layer3_outputs(3309) <= not(layer2_outputs(4795));
    layer3_outputs(3310) <= not(layer2_outputs(4899)) or (layer2_outputs(210));
    layer3_outputs(3311) <= not(layer2_outputs(7988));
    layer3_outputs(3312) <= (layer2_outputs(8184)) xor (layer2_outputs(9629));
    layer3_outputs(3313) <= (layer2_outputs(6191)) xor (layer2_outputs(10211));
    layer3_outputs(3314) <= (layer2_outputs(2524)) and not (layer2_outputs(1015));
    layer3_outputs(3315) <= not(layer2_outputs(7014));
    layer3_outputs(3316) <= (layer2_outputs(6948)) and (layer2_outputs(1444));
    layer3_outputs(3317) <= not(layer2_outputs(758));
    layer3_outputs(3318) <= layer2_outputs(1065);
    layer3_outputs(3319) <= not((layer2_outputs(1136)) xor (layer2_outputs(2480)));
    layer3_outputs(3320) <= '1';
    layer3_outputs(3321) <= not((layer2_outputs(1827)) or (layer2_outputs(6014)));
    layer3_outputs(3322) <= layer2_outputs(362);
    layer3_outputs(3323) <= not(layer2_outputs(1844)) or (layer2_outputs(10103));
    layer3_outputs(3324) <= not(layer2_outputs(8060));
    layer3_outputs(3325) <= layer2_outputs(7160);
    layer3_outputs(3326) <= not(layer2_outputs(5511));
    layer3_outputs(3327) <= not(layer2_outputs(5187));
    layer3_outputs(3328) <= layer2_outputs(8397);
    layer3_outputs(3329) <= not(layer2_outputs(3870)) or (layer2_outputs(1661));
    layer3_outputs(3330) <= not(layer2_outputs(10076)) or (layer2_outputs(5507));
    layer3_outputs(3331) <= '1';
    layer3_outputs(3332) <= (layer2_outputs(5171)) and not (layer2_outputs(3387));
    layer3_outputs(3333) <= '1';
    layer3_outputs(3334) <= layer2_outputs(94);
    layer3_outputs(3335) <= not(layer2_outputs(5039));
    layer3_outputs(3336) <= not((layer2_outputs(7909)) and (layer2_outputs(8752)));
    layer3_outputs(3337) <= layer2_outputs(5923);
    layer3_outputs(3338) <= not((layer2_outputs(6552)) or (layer2_outputs(1560)));
    layer3_outputs(3339) <= not((layer2_outputs(534)) and (layer2_outputs(8958)));
    layer3_outputs(3340) <= not(layer2_outputs(7870));
    layer3_outputs(3341) <= (layer2_outputs(6233)) and not (layer2_outputs(9835));
    layer3_outputs(3342) <= not(layer2_outputs(1589));
    layer3_outputs(3343) <= (layer2_outputs(6894)) and (layer2_outputs(968));
    layer3_outputs(3344) <= not(layer2_outputs(4222));
    layer3_outputs(3345) <= not(layer2_outputs(2173));
    layer3_outputs(3346) <= not((layer2_outputs(2079)) xor (layer2_outputs(782)));
    layer3_outputs(3347) <= not(layer2_outputs(2977));
    layer3_outputs(3348) <= layer2_outputs(2365);
    layer3_outputs(3349) <= not((layer2_outputs(83)) and (layer2_outputs(1361)));
    layer3_outputs(3350) <= not((layer2_outputs(2746)) or (layer2_outputs(7894)));
    layer3_outputs(3351) <= not((layer2_outputs(6335)) and (layer2_outputs(2128)));
    layer3_outputs(3352) <= (layer2_outputs(5651)) and (layer2_outputs(1733));
    layer3_outputs(3353) <= (layer2_outputs(5337)) xor (layer2_outputs(7007));
    layer3_outputs(3354) <= not((layer2_outputs(1687)) xor (layer2_outputs(7508)));
    layer3_outputs(3355) <= (layer2_outputs(1400)) and not (layer2_outputs(10023));
    layer3_outputs(3356) <= layer2_outputs(9750);
    layer3_outputs(3357) <= not(layer2_outputs(7567));
    layer3_outputs(3358) <= not((layer2_outputs(3037)) or (layer2_outputs(9840)));
    layer3_outputs(3359) <= not(layer2_outputs(6536));
    layer3_outputs(3360) <= not(layer2_outputs(6689));
    layer3_outputs(3361) <= layer2_outputs(2601);
    layer3_outputs(3362) <= (layer2_outputs(8129)) or (layer2_outputs(2061));
    layer3_outputs(3363) <= not((layer2_outputs(3112)) or (layer2_outputs(5947)));
    layer3_outputs(3364) <= not(layer2_outputs(3900));
    layer3_outputs(3365) <= not(layer2_outputs(2855));
    layer3_outputs(3366) <= layer2_outputs(5493);
    layer3_outputs(3367) <= (layer2_outputs(1355)) or (layer2_outputs(8741));
    layer3_outputs(3368) <= not(layer2_outputs(10156));
    layer3_outputs(3369) <= not(layer2_outputs(2058));
    layer3_outputs(3370) <= (layer2_outputs(1631)) or (layer2_outputs(9928));
    layer3_outputs(3371) <= layer2_outputs(8075);
    layer3_outputs(3372) <= not(layer2_outputs(1311));
    layer3_outputs(3373) <= not((layer2_outputs(1220)) or (layer2_outputs(5340)));
    layer3_outputs(3374) <= (layer2_outputs(2289)) xor (layer2_outputs(8390));
    layer3_outputs(3375) <= not(layer2_outputs(9009));
    layer3_outputs(3376) <= layer2_outputs(5577);
    layer3_outputs(3377) <= '0';
    layer3_outputs(3378) <= layer2_outputs(6468);
    layer3_outputs(3379) <= not(layer2_outputs(9989));
    layer3_outputs(3380) <= not((layer2_outputs(765)) or (layer2_outputs(6915)));
    layer3_outputs(3381) <= (layer2_outputs(8667)) and not (layer2_outputs(4760));
    layer3_outputs(3382) <= layer2_outputs(6740);
    layer3_outputs(3383) <= not(layer2_outputs(6683));
    layer3_outputs(3384) <= not(layer2_outputs(3004)) or (layer2_outputs(9729));
    layer3_outputs(3385) <= '1';
    layer3_outputs(3386) <= layer2_outputs(1621);
    layer3_outputs(3387) <= (layer2_outputs(8664)) and (layer2_outputs(3378));
    layer3_outputs(3388) <= not(layer2_outputs(6762));
    layer3_outputs(3389) <= (layer2_outputs(4974)) and (layer2_outputs(4098));
    layer3_outputs(3390) <= (layer2_outputs(7403)) and (layer2_outputs(2054));
    layer3_outputs(3391) <= (layer2_outputs(3434)) or (layer2_outputs(2725));
    layer3_outputs(3392) <= not((layer2_outputs(10089)) or (layer2_outputs(5998)));
    layer3_outputs(3393) <= not(layer2_outputs(7753)) or (layer2_outputs(7020));
    layer3_outputs(3394) <= '0';
    layer3_outputs(3395) <= not(layer2_outputs(9055));
    layer3_outputs(3396) <= (layer2_outputs(7827)) and not (layer2_outputs(729));
    layer3_outputs(3397) <= layer2_outputs(9965);
    layer3_outputs(3398) <= layer2_outputs(6383);
    layer3_outputs(3399) <= (layer2_outputs(7813)) and (layer2_outputs(6243));
    layer3_outputs(3400) <= layer2_outputs(3309);
    layer3_outputs(3401) <= not(layer2_outputs(1131));
    layer3_outputs(3402) <= layer2_outputs(3864);
    layer3_outputs(3403) <= not((layer2_outputs(4423)) or (layer2_outputs(594)));
    layer3_outputs(3404) <= (layer2_outputs(8351)) and not (layer2_outputs(7298));
    layer3_outputs(3405) <= not(layer2_outputs(7387));
    layer3_outputs(3406) <= layer2_outputs(212);
    layer3_outputs(3407) <= not(layer2_outputs(9410)) or (layer2_outputs(1074));
    layer3_outputs(3408) <= layer2_outputs(5605);
    layer3_outputs(3409) <= layer2_outputs(7382);
    layer3_outputs(3410) <= layer2_outputs(5189);
    layer3_outputs(3411) <= (layer2_outputs(3939)) or (layer2_outputs(8753));
    layer3_outputs(3412) <= layer2_outputs(5205);
    layer3_outputs(3413) <= not(layer2_outputs(724));
    layer3_outputs(3414) <= layer2_outputs(3672);
    layer3_outputs(3415) <= (layer2_outputs(3997)) xor (layer2_outputs(580));
    layer3_outputs(3416) <= layer2_outputs(3610);
    layer3_outputs(3417) <= layer2_outputs(9221);
    layer3_outputs(3418) <= not((layer2_outputs(8932)) and (layer2_outputs(4684)));
    layer3_outputs(3419) <= (layer2_outputs(9872)) xor (layer2_outputs(6505));
    layer3_outputs(3420) <= not(layer2_outputs(4848));
    layer3_outputs(3421) <= not((layer2_outputs(46)) or (layer2_outputs(2042)));
    layer3_outputs(3422) <= not((layer2_outputs(5688)) and (layer2_outputs(300)));
    layer3_outputs(3423) <= not(layer2_outputs(754));
    layer3_outputs(3424) <= (layer2_outputs(3058)) or (layer2_outputs(956));
    layer3_outputs(3425) <= (layer2_outputs(7880)) and not (layer2_outputs(8599));
    layer3_outputs(3426) <= not(layer2_outputs(8491)) or (layer2_outputs(671));
    layer3_outputs(3427) <= (layer2_outputs(6904)) and not (layer2_outputs(1740));
    layer3_outputs(3428) <= (layer2_outputs(266)) and not (layer2_outputs(8934));
    layer3_outputs(3429) <= not(layer2_outputs(9249));
    layer3_outputs(3430) <= layer2_outputs(3598);
    layer3_outputs(3431) <= layer2_outputs(7330);
    layer3_outputs(3432) <= not((layer2_outputs(4559)) xor (layer2_outputs(712)));
    layer3_outputs(3433) <= layer2_outputs(6794);
    layer3_outputs(3434) <= layer2_outputs(2386);
    layer3_outputs(3435) <= layer2_outputs(6314);
    layer3_outputs(3436) <= layer2_outputs(9427);
    layer3_outputs(3437) <= (layer2_outputs(7084)) and (layer2_outputs(2902));
    layer3_outputs(3438) <= layer2_outputs(4639);
    layer3_outputs(3439) <= not(layer2_outputs(8769));
    layer3_outputs(3440) <= (layer2_outputs(4720)) and not (layer2_outputs(5129));
    layer3_outputs(3441) <= not(layer2_outputs(3030));
    layer3_outputs(3442) <= (layer2_outputs(5214)) or (layer2_outputs(8548));
    layer3_outputs(3443) <= not(layer2_outputs(1117));
    layer3_outputs(3444) <= not(layer2_outputs(7391));
    layer3_outputs(3445) <= '1';
    layer3_outputs(3446) <= not(layer2_outputs(3090));
    layer3_outputs(3447) <= not(layer2_outputs(1948));
    layer3_outputs(3448) <= not((layer2_outputs(2446)) or (layer2_outputs(9875)));
    layer3_outputs(3449) <= (layer2_outputs(2657)) and (layer2_outputs(4135));
    layer3_outputs(3450) <= '0';
    layer3_outputs(3451) <= layer2_outputs(5556);
    layer3_outputs(3452) <= layer2_outputs(1679);
    layer3_outputs(3453) <= (layer2_outputs(7999)) and (layer2_outputs(8209));
    layer3_outputs(3454) <= '0';
    layer3_outputs(3455) <= (layer2_outputs(8512)) and (layer2_outputs(9617));
    layer3_outputs(3456) <= not(layer2_outputs(6572)) or (layer2_outputs(2186));
    layer3_outputs(3457) <= not(layer2_outputs(7733));
    layer3_outputs(3458) <= (layer2_outputs(8936)) or (layer2_outputs(67));
    layer3_outputs(3459) <= layer2_outputs(1486);
    layer3_outputs(3460) <= layer2_outputs(2838);
    layer3_outputs(3461) <= not(layer2_outputs(4063));
    layer3_outputs(3462) <= (layer2_outputs(6320)) and (layer2_outputs(6016));
    layer3_outputs(3463) <= not(layer2_outputs(3424)) or (layer2_outputs(5913));
    layer3_outputs(3464) <= not(layer2_outputs(6916)) or (layer2_outputs(3380));
    layer3_outputs(3465) <= not((layer2_outputs(2307)) xor (layer2_outputs(4440)));
    layer3_outputs(3466) <= not((layer2_outputs(5479)) or (layer2_outputs(3654)));
    layer3_outputs(3467) <= not((layer2_outputs(9949)) or (layer2_outputs(1617)));
    layer3_outputs(3468) <= '0';
    layer3_outputs(3469) <= not(layer2_outputs(9503));
    layer3_outputs(3470) <= not(layer2_outputs(2840));
    layer3_outputs(3471) <= (layer2_outputs(4733)) and (layer2_outputs(676));
    layer3_outputs(3472) <= not(layer2_outputs(7667));
    layer3_outputs(3473) <= not(layer2_outputs(1271)) or (layer2_outputs(350));
    layer3_outputs(3474) <= not((layer2_outputs(1449)) and (layer2_outputs(2467)));
    layer3_outputs(3475) <= not(layer2_outputs(985)) or (layer2_outputs(7400));
    layer3_outputs(3476) <= not(layer2_outputs(2113));
    layer3_outputs(3477) <= not(layer2_outputs(511)) or (layer2_outputs(3188));
    layer3_outputs(3478) <= not(layer2_outputs(5532)) or (layer2_outputs(9642));
    layer3_outputs(3479) <= not(layer2_outputs(4448)) or (layer2_outputs(5099));
    layer3_outputs(3480) <= not(layer2_outputs(2326)) or (layer2_outputs(2020));
    layer3_outputs(3481) <= (layer2_outputs(4227)) and not (layer2_outputs(4078));
    layer3_outputs(3482) <= (layer2_outputs(6276)) xor (layer2_outputs(6876));
    layer3_outputs(3483) <= (layer2_outputs(6521)) and (layer2_outputs(9190));
    layer3_outputs(3484) <= layer2_outputs(6371);
    layer3_outputs(3485) <= layer2_outputs(3225);
    layer3_outputs(3486) <= layer2_outputs(5552);
    layer3_outputs(3487) <= not((layer2_outputs(2379)) xor (layer2_outputs(9455)));
    layer3_outputs(3488) <= not(layer2_outputs(2666)) or (layer2_outputs(10130));
    layer3_outputs(3489) <= layer2_outputs(7805);
    layer3_outputs(3490) <= layer2_outputs(561);
    layer3_outputs(3491) <= (layer2_outputs(7444)) or (layer2_outputs(6863));
    layer3_outputs(3492) <= not(layer2_outputs(8097)) or (layer2_outputs(785));
    layer3_outputs(3493) <= not(layer2_outputs(5808)) or (layer2_outputs(4680));
    layer3_outputs(3494) <= '0';
    layer3_outputs(3495) <= (layer2_outputs(3199)) or (layer2_outputs(1052));
    layer3_outputs(3496) <= (layer2_outputs(2446)) xor (layer2_outputs(6760));
    layer3_outputs(3497) <= (layer2_outputs(9187)) and (layer2_outputs(4484));
    layer3_outputs(3498) <= not(layer2_outputs(3259));
    layer3_outputs(3499) <= layer2_outputs(9735);
    layer3_outputs(3500) <= layer2_outputs(9334);
    layer3_outputs(3501) <= layer2_outputs(5288);
    layer3_outputs(3502) <= (layer2_outputs(2885)) and (layer2_outputs(5014));
    layer3_outputs(3503) <= (layer2_outputs(7995)) and not (layer2_outputs(358));
    layer3_outputs(3504) <= (layer2_outputs(3310)) xor (layer2_outputs(10172));
    layer3_outputs(3505) <= not((layer2_outputs(1118)) and (layer2_outputs(2193)));
    layer3_outputs(3506) <= layer2_outputs(7064);
    layer3_outputs(3507) <= layer2_outputs(1755);
    layer3_outputs(3508) <= layer2_outputs(6869);
    layer3_outputs(3509) <= not((layer2_outputs(8506)) or (layer2_outputs(4183)));
    layer3_outputs(3510) <= not(layer2_outputs(8954));
    layer3_outputs(3511) <= (layer2_outputs(9313)) xor (layer2_outputs(8730));
    layer3_outputs(3512) <= not((layer2_outputs(5714)) and (layer2_outputs(6878)));
    layer3_outputs(3513) <= not(layer2_outputs(7321));
    layer3_outputs(3514) <= (layer2_outputs(3766)) or (layer2_outputs(1924));
    layer3_outputs(3515) <= layer2_outputs(640);
    layer3_outputs(3516) <= not(layer2_outputs(3423));
    layer3_outputs(3517) <= (layer2_outputs(6051)) xor (layer2_outputs(8644));
    layer3_outputs(3518) <= layer2_outputs(5984);
    layer3_outputs(3519) <= not(layer2_outputs(3952));
    layer3_outputs(3520) <= layer2_outputs(9855);
    layer3_outputs(3521) <= (layer2_outputs(1781)) and not (layer2_outputs(292));
    layer3_outputs(3522) <= layer2_outputs(1803);
    layer3_outputs(3523) <= not(layer2_outputs(8767));
    layer3_outputs(3524) <= (layer2_outputs(6841)) and not (layer2_outputs(9831));
    layer3_outputs(3525) <= (layer2_outputs(1417)) and (layer2_outputs(5011));
    layer3_outputs(3526) <= not(layer2_outputs(7373));
    layer3_outputs(3527) <= (layer2_outputs(10180)) or (layer2_outputs(930));
    layer3_outputs(3528) <= (layer2_outputs(4796)) and not (layer2_outputs(2876));
    layer3_outputs(3529) <= not((layer2_outputs(8367)) and (layer2_outputs(7270)));
    layer3_outputs(3530) <= not(layer2_outputs(4067));
    layer3_outputs(3531) <= not(layer2_outputs(4645));
    layer3_outputs(3532) <= not((layer2_outputs(5559)) xor (layer2_outputs(2705)));
    layer3_outputs(3533) <= '1';
    layer3_outputs(3534) <= not(layer2_outputs(8161));
    layer3_outputs(3535) <= not(layer2_outputs(6868));
    layer3_outputs(3536) <= (layer2_outputs(8647)) and not (layer2_outputs(9565));
    layer3_outputs(3537) <= (layer2_outputs(705)) and (layer2_outputs(6274));
    layer3_outputs(3538) <= not((layer2_outputs(8498)) and (layer2_outputs(9384)));
    layer3_outputs(3539) <= (layer2_outputs(2981)) and not (layer2_outputs(4470));
    layer3_outputs(3540) <= not(layer2_outputs(2214)) or (layer2_outputs(7965));
    layer3_outputs(3541) <= layer2_outputs(9317);
    layer3_outputs(3542) <= not(layer2_outputs(10202));
    layer3_outputs(3543) <= not(layer2_outputs(2714));
    layer3_outputs(3544) <= (layer2_outputs(4668)) and (layer2_outputs(3096));
    layer3_outputs(3545) <= (layer2_outputs(3316)) and (layer2_outputs(2567));
    layer3_outputs(3546) <= '0';
    layer3_outputs(3547) <= layer2_outputs(9265);
    layer3_outputs(3548) <= not(layer2_outputs(7408)) or (layer2_outputs(3497));
    layer3_outputs(3549) <= not(layer2_outputs(948));
    layer3_outputs(3550) <= (layer2_outputs(9018)) xor (layer2_outputs(2158));
    layer3_outputs(3551) <= not(layer2_outputs(3370));
    layer3_outputs(3552) <= not(layer2_outputs(2404));
    layer3_outputs(3553) <= layer2_outputs(1371);
    layer3_outputs(3554) <= not(layer2_outputs(893));
    layer3_outputs(3555) <= not((layer2_outputs(1054)) and (layer2_outputs(223)));
    layer3_outputs(3556) <= layer2_outputs(2756);
    layer3_outputs(3557) <= (layer2_outputs(6801)) and not (layer2_outputs(5041));
    layer3_outputs(3558) <= '0';
    layer3_outputs(3559) <= not(layer2_outputs(3787));
    layer3_outputs(3560) <= not((layer2_outputs(1120)) xor (layer2_outputs(4410)));
    layer3_outputs(3561) <= layer2_outputs(5598);
    layer3_outputs(3562) <= not((layer2_outputs(5568)) or (layer2_outputs(4741)));
    layer3_outputs(3563) <= not(layer2_outputs(6355));
    layer3_outputs(3564) <= (layer2_outputs(10124)) xor (layer2_outputs(8724));
    layer3_outputs(3565) <= (layer2_outputs(7789)) and not (layer2_outputs(8881));
    layer3_outputs(3566) <= not(layer2_outputs(801));
    layer3_outputs(3567) <= layer2_outputs(670);
    layer3_outputs(3568) <= (layer2_outputs(9078)) and (layer2_outputs(4975));
    layer3_outputs(3569) <= not((layer2_outputs(527)) or (layer2_outputs(4282)));
    layer3_outputs(3570) <= not(layer2_outputs(4817)) or (layer2_outputs(5716));
    layer3_outputs(3571) <= not((layer2_outputs(7688)) xor (layer2_outputs(451)));
    layer3_outputs(3572) <= layer2_outputs(5801);
    layer3_outputs(3573) <= not(layer2_outputs(2124));
    layer3_outputs(3574) <= not((layer2_outputs(4851)) and (layer2_outputs(5948)));
    layer3_outputs(3575) <= '1';
    layer3_outputs(3576) <= layer2_outputs(6807);
    layer3_outputs(3577) <= not((layer2_outputs(3495)) xor (layer2_outputs(4709)));
    layer3_outputs(3578) <= layer2_outputs(8967);
    layer3_outputs(3579) <= (layer2_outputs(8130)) and not (layer2_outputs(7932));
    layer3_outputs(3580) <= (layer2_outputs(1732)) and not (layer2_outputs(6576));
    layer3_outputs(3581) <= not(layer2_outputs(6625));
    layer3_outputs(3582) <= (layer2_outputs(3613)) and not (layer2_outputs(1712));
    layer3_outputs(3583) <= not(layer2_outputs(4923));
    layer3_outputs(3584) <= not(layer2_outputs(1446));
    layer3_outputs(3585) <= not((layer2_outputs(7181)) and (layer2_outputs(3102)));
    layer3_outputs(3586) <= not((layer2_outputs(6458)) xor (layer2_outputs(4451)));
    layer3_outputs(3587) <= not(layer2_outputs(572));
    layer3_outputs(3588) <= layer2_outputs(6154);
    layer3_outputs(3589) <= not(layer2_outputs(5727));
    layer3_outputs(3590) <= not(layer2_outputs(1413)) or (layer2_outputs(9932));
    layer3_outputs(3591) <= not(layer2_outputs(9460));
    layer3_outputs(3592) <= (layer2_outputs(8415)) and not (layer2_outputs(830));
    layer3_outputs(3593) <= not(layer2_outputs(7544));
    layer3_outputs(3594) <= (layer2_outputs(7326)) or (layer2_outputs(9051));
    layer3_outputs(3595) <= layer2_outputs(5777);
    layer3_outputs(3596) <= (layer2_outputs(1686)) and (layer2_outputs(374));
    layer3_outputs(3597) <= (layer2_outputs(5569)) xor (layer2_outputs(8702));
    layer3_outputs(3598) <= layer2_outputs(9080);
    layer3_outputs(3599) <= layer2_outputs(9243);
    layer3_outputs(3600) <= not(layer2_outputs(9662)) or (layer2_outputs(37));
    layer3_outputs(3601) <= layer2_outputs(8036);
    layer3_outputs(3602) <= (layer2_outputs(6898)) or (layer2_outputs(8997));
    layer3_outputs(3603) <= layer2_outputs(3572);
    layer3_outputs(3604) <= layer2_outputs(4541);
    layer3_outputs(3605) <= layer2_outputs(6258);
    layer3_outputs(3606) <= (layer2_outputs(7822)) and (layer2_outputs(7165));
    layer3_outputs(3607) <= not((layer2_outputs(4104)) and (layer2_outputs(1308)));
    layer3_outputs(3608) <= layer2_outputs(2700);
    layer3_outputs(3609) <= layer2_outputs(4620);
    layer3_outputs(3610) <= not(layer2_outputs(7834));
    layer3_outputs(3611) <= (layer2_outputs(10087)) or (layer2_outputs(6026));
    layer3_outputs(3612) <= not(layer2_outputs(3587));
    layer3_outputs(3613) <= not(layer2_outputs(1098)) or (layer2_outputs(7027));
    layer3_outputs(3614) <= not(layer2_outputs(8201));
    layer3_outputs(3615) <= layer2_outputs(6449);
    layer3_outputs(3616) <= not((layer2_outputs(7720)) xor (layer2_outputs(4389)));
    layer3_outputs(3617) <= not(layer2_outputs(3918));
    layer3_outputs(3618) <= (layer2_outputs(2578)) or (layer2_outputs(8652));
    layer3_outputs(3619) <= layer2_outputs(4882);
    layer3_outputs(3620) <= not((layer2_outputs(969)) xor (layer2_outputs(6819)));
    layer3_outputs(3621) <= (layer2_outputs(1212)) and not (layer2_outputs(2219));
    layer3_outputs(3622) <= not(layer2_outputs(7439));
    layer3_outputs(3623) <= (layer2_outputs(6076)) and not (layer2_outputs(613));
    layer3_outputs(3624) <= not(layer2_outputs(5677)) or (layer2_outputs(1510));
    layer3_outputs(3625) <= not(layer2_outputs(3862)) or (layer2_outputs(9013));
    layer3_outputs(3626) <= not(layer2_outputs(7519));
    layer3_outputs(3627) <= not(layer2_outputs(917)) or (layer2_outputs(5259));
    layer3_outputs(3628) <= layer2_outputs(4520);
    layer3_outputs(3629) <= layer2_outputs(1571);
    layer3_outputs(3630) <= (layer2_outputs(2918)) and not (layer2_outputs(5113));
    layer3_outputs(3631) <= '1';
    layer3_outputs(3632) <= not(layer2_outputs(2989));
    layer3_outputs(3633) <= layer2_outputs(3455);
    layer3_outputs(3634) <= not(layer2_outputs(1011)) or (layer2_outputs(7087));
    layer3_outputs(3635) <= not(layer2_outputs(9820));
    layer3_outputs(3636) <= not((layer2_outputs(1525)) or (layer2_outputs(65)));
    layer3_outputs(3637) <= (layer2_outputs(6783)) and (layer2_outputs(6158));
    layer3_outputs(3638) <= not(layer2_outputs(8093));
    layer3_outputs(3639) <= (layer2_outputs(7711)) and not (layer2_outputs(927));
    layer3_outputs(3640) <= not((layer2_outputs(1435)) or (layer2_outputs(5137)));
    layer3_outputs(3641) <= not(layer2_outputs(3740));
    layer3_outputs(3642) <= layer2_outputs(208);
    layer3_outputs(3643) <= layer2_outputs(6809);
    layer3_outputs(3644) <= not(layer2_outputs(10080));
    layer3_outputs(3645) <= not(layer2_outputs(9186));
    layer3_outputs(3646) <= layer2_outputs(3063);
    layer3_outputs(3647) <= not((layer2_outputs(3855)) and (layer2_outputs(5423)));
    layer3_outputs(3648) <= layer2_outputs(86);
    layer3_outputs(3649) <= not(layer2_outputs(6723));
    layer3_outputs(3650) <= '1';
    layer3_outputs(3651) <= (layer2_outputs(5244)) xor (layer2_outputs(1567));
    layer3_outputs(3652) <= not(layer2_outputs(767)) or (layer2_outputs(3747));
    layer3_outputs(3653) <= not((layer2_outputs(7451)) and (layer2_outputs(6770)));
    layer3_outputs(3654) <= '0';
    layer3_outputs(3655) <= (layer2_outputs(9446)) and not (layer2_outputs(1502));
    layer3_outputs(3656) <= not(layer2_outputs(2767));
    layer3_outputs(3657) <= layer2_outputs(3107);
    layer3_outputs(3658) <= not(layer2_outputs(6186));
    layer3_outputs(3659) <= not(layer2_outputs(6000)) or (layer2_outputs(8949));
    layer3_outputs(3660) <= not(layer2_outputs(6542));
    layer3_outputs(3661) <= '1';
    layer3_outputs(3662) <= layer2_outputs(7525);
    layer3_outputs(3663) <= not(layer2_outputs(2602));
    layer3_outputs(3664) <= (layer2_outputs(1109)) and not (layer2_outputs(9343));
    layer3_outputs(3665) <= not((layer2_outputs(2497)) and (layer2_outputs(6759)));
    layer3_outputs(3666) <= (layer2_outputs(470)) and not (layer2_outputs(7262));
    layer3_outputs(3667) <= (layer2_outputs(1677)) and not (layer2_outputs(1934));
    layer3_outputs(3668) <= layer2_outputs(6855);
    layer3_outputs(3669) <= (layer2_outputs(7597)) and not (layer2_outputs(1925));
    layer3_outputs(3670) <= (layer2_outputs(8259)) or (layer2_outputs(9657));
    layer3_outputs(3671) <= (layer2_outputs(8471)) and (layer2_outputs(3278));
    layer3_outputs(3672) <= layer2_outputs(7248);
    layer3_outputs(3673) <= layer2_outputs(9396);
    layer3_outputs(3674) <= (layer2_outputs(9410)) xor (layer2_outputs(7832));
    layer3_outputs(3675) <= layer2_outputs(8817);
    layer3_outputs(3676) <= not(layer2_outputs(1828)) or (layer2_outputs(4023));
    layer3_outputs(3677) <= '1';
    layer3_outputs(3678) <= not((layer2_outputs(4511)) xor (layer2_outputs(8870)));
    layer3_outputs(3679) <= '1';
    layer3_outputs(3680) <= not(layer2_outputs(5655));
    layer3_outputs(3681) <= not(layer2_outputs(2744));
    layer3_outputs(3682) <= not(layer2_outputs(5411));
    layer3_outputs(3683) <= layer2_outputs(8150);
    layer3_outputs(3684) <= layer2_outputs(4562);
    layer3_outputs(3685) <= not(layer2_outputs(210)) or (layer2_outputs(3958));
    layer3_outputs(3686) <= (layer2_outputs(2432)) and not (layer2_outputs(7446));
    layer3_outputs(3687) <= (layer2_outputs(7489)) and not (layer2_outputs(2191));
    layer3_outputs(3688) <= (layer2_outputs(6412)) or (layer2_outputs(8467));
    layer3_outputs(3689) <= (layer2_outputs(1179)) or (layer2_outputs(5545));
    layer3_outputs(3690) <= layer2_outputs(1124);
    layer3_outputs(3691) <= not(layer2_outputs(4757)) or (layer2_outputs(9953));
    layer3_outputs(3692) <= (layer2_outputs(952)) or (layer2_outputs(6088));
    layer3_outputs(3693) <= (layer2_outputs(6145)) and not (layer2_outputs(2790));
    layer3_outputs(3694) <= (layer2_outputs(5606)) or (layer2_outputs(3560));
    layer3_outputs(3695) <= '1';
    layer3_outputs(3696) <= (layer2_outputs(9544)) and (layer2_outputs(3783));
    layer3_outputs(3697) <= not(layer2_outputs(1734));
    layer3_outputs(3698) <= (layer2_outputs(7402)) and not (layer2_outputs(1957));
    layer3_outputs(3699) <= not(layer2_outputs(4330)) or (layer2_outputs(8205));
    layer3_outputs(3700) <= '1';
    layer3_outputs(3701) <= (layer2_outputs(7487)) and not (layer2_outputs(7014));
    layer3_outputs(3702) <= '1';
    layer3_outputs(3703) <= (layer2_outputs(5194)) or (layer2_outputs(9741));
    layer3_outputs(3704) <= (layer2_outputs(8244)) and not (layer2_outputs(922));
    layer3_outputs(3705) <= (layer2_outputs(5077)) and not (layer2_outputs(5455));
    layer3_outputs(3706) <= not(layer2_outputs(5340)) or (layer2_outputs(7290));
    layer3_outputs(3707) <= not((layer2_outputs(9129)) xor (layer2_outputs(5252)));
    layer3_outputs(3708) <= (layer2_outputs(6435)) and not (layer2_outputs(1280));
    layer3_outputs(3709) <= (layer2_outputs(2549)) xor (layer2_outputs(4948));
    layer3_outputs(3710) <= (layer2_outputs(2749)) xor (layer2_outputs(2899));
    layer3_outputs(3711) <= not(layer2_outputs(531));
    layer3_outputs(3712) <= (layer2_outputs(9535)) or (layer2_outputs(5098));
    layer3_outputs(3713) <= not(layer2_outputs(6909));
    layer3_outputs(3714) <= not(layer2_outputs(7019)) or (layer2_outputs(9729));
    layer3_outputs(3715) <= not(layer2_outputs(1152));
    layer3_outputs(3716) <= not(layer2_outputs(4693));
    layer3_outputs(3717) <= layer2_outputs(4083);
    layer3_outputs(3718) <= not(layer2_outputs(8442));
    layer3_outputs(3719) <= layer2_outputs(1871);
    layer3_outputs(3720) <= not(layer2_outputs(6609)) or (layer2_outputs(6638));
    layer3_outputs(3721) <= not((layer2_outputs(8990)) xor (layer2_outputs(8367)));
    layer3_outputs(3722) <= layer2_outputs(2648);
    layer3_outputs(3723) <= not((layer2_outputs(7911)) xor (layer2_outputs(8431)));
    layer3_outputs(3724) <= not((layer2_outputs(888)) xor (layer2_outputs(288)));
    layer3_outputs(3725) <= not(layer2_outputs(8904));
    layer3_outputs(3726) <= (layer2_outputs(315)) and not (layer2_outputs(1792));
    layer3_outputs(3727) <= not(layer2_outputs(494));
    layer3_outputs(3728) <= not(layer2_outputs(9347));
    layer3_outputs(3729) <= (layer2_outputs(6571)) xor (layer2_outputs(4748));
    layer3_outputs(3730) <= (layer2_outputs(8058)) or (layer2_outputs(4587));
    layer3_outputs(3731) <= (layer2_outputs(5194)) and not (layer2_outputs(7802));
    layer3_outputs(3732) <= not(layer2_outputs(9405));
    layer3_outputs(3733) <= layer2_outputs(8757);
    layer3_outputs(3734) <= layer2_outputs(5636);
    layer3_outputs(3735) <= (layer2_outputs(5575)) and not (layer2_outputs(3640));
    layer3_outputs(3736) <= layer2_outputs(4652);
    layer3_outputs(3737) <= (layer2_outputs(1775)) xor (layer2_outputs(4829));
    layer3_outputs(3738) <= not((layer2_outputs(2051)) xor (layer2_outputs(3648)));
    layer3_outputs(3739) <= not(layer2_outputs(6538));
    layer3_outputs(3740) <= (layer2_outputs(4498)) and not (layer2_outputs(9671));
    layer3_outputs(3741) <= not(layer2_outputs(402)) or (layer2_outputs(6627));
    layer3_outputs(3742) <= '0';
    layer3_outputs(3743) <= not(layer2_outputs(2179));
    layer3_outputs(3744) <= (layer2_outputs(1511)) and not (layer2_outputs(9677));
    layer3_outputs(3745) <= not((layer2_outputs(3924)) xor (layer2_outputs(8600)));
    layer3_outputs(3746) <= layer2_outputs(7785);
    layer3_outputs(3747) <= layer2_outputs(6545);
    layer3_outputs(3748) <= layer2_outputs(5000);
    layer3_outputs(3749) <= not(layer2_outputs(1137));
    layer3_outputs(3750) <= not(layer2_outputs(9226));
    layer3_outputs(3751) <= (layer2_outputs(3238)) and not (layer2_outputs(9176));
    layer3_outputs(3752) <= (layer2_outputs(4106)) and not (layer2_outputs(900));
    layer3_outputs(3753) <= not(layer2_outputs(6600));
    layer3_outputs(3754) <= not(layer2_outputs(6873));
    layer3_outputs(3755) <= not(layer2_outputs(3188));
    layer3_outputs(3756) <= (layer2_outputs(7694)) xor (layer2_outputs(376));
    layer3_outputs(3757) <= not(layer2_outputs(4938));
    layer3_outputs(3758) <= not(layer2_outputs(3704)) or (layer2_outputs(6874));
    layer3_outputs(3759) <= (layer2_outputs(4609)) and not (layer2_outputs(1644));
    layer3_outputs(3760) <= not(layer2_outputs(125)) or (layer2_outputs(4344));
    layer3_outputs(3761) <= layer2_outputs(960);
    layer3_outputs(3762) <= layer2_outputs(218);
    layer3_outputs(3763) <= layer2_outputs(5207);
    layer3_outputs(3764) <= (layer2_outputs(1632)) and not (layer2_outputs(8597));
    layer3_outputs(3765) <= not(layer2_outputs(7197));
    layer3_outputs(3766) <= not(layer2_outputs(7755)) or (layer2_outputs(619));
    layer3_outputs(3767) <= layer2_outputs(7179);
    layer3_outputs(3768) <= not((layer2_outputs(8412)) and (layer2_outputs(1297)));
    layer3_outputs(3769) <= not(layer2_outputs(9812)) or (layer2_outputs(1959));
    layer3_outputs(3770) <= layer2_outputs(8203);
    layer3_outputs(3771) <= (layer2_outputs(5436)) and not (layer2_outputs(3202));
    layer3_outputs(3772) <= not(layer2_outputs(9080));
    layer3_outputs(3773) <= layer2_outputs(9191);
    layer3_outputs(3774) <= (layer2_outputs(3971)) and (layer2_outputs(3514));
    layer3_outputs(3775) <= (layer2_outputs(915)) and not (layer2_outputs(5749));
    layer3_outputs(3776) <= not(layer2_outputs(10099));
    layer3_outputs(3777) <= layer2_outputs(936);
    layer3_outputs(3778) <= layer2_outputs(1283);
    layer3_outputs(3779) <= not(layer2_outputs(3693));
    layer3_outputs(3780) <= (layer2_outputs(3825)) and not (layer2_outputs(7937));
    layer3_outputs(3781) <= not(layer2_outputs(8992));
    layer3_outputs(3782) <= '0';
    layer3_outputs(3783) <= (layer2_outputs(1957)) or (layer2_outputs(4857));
    layer3_outputs(3784) <= not((layer2_outputs(3733)) or (layer2_outputs(4546)));
    layer3_outputs(3785) <= (layer2_outputs(1111)) or (layer2_outputs(2708));
    layer3_outputs(3786) <= (layer2_outputs(8404)) and not (layer2_outputs(887));
    layer3_outputs(3787) <= layer2_outputs(1203);
    layer3_outputs(3788) <= layer2_outputs(10162);
    layer3_outputs(3789) <= layer2_outputs(4052);
    layer3_outputs(3790) <= not((layer2_outputs(3782)) or (layer2_outputs(9089)));
    layer3_outputs(3791) <= (layer2_outputs(6629)) and (layer2_outputs(3048));
    layer3_outputs(3792) <= layer2_outputs(2038);
    layer3_outputs(3793) <= not(layer2_outputs(1211));
    layer3_outputs(3794) <= (layer2_outputs(9474)) or (layer2_outputs(3589));
    layer3_outputs(3795) <= layer2_outputs(5677);
    layer3_outputs(3796) <= not(layer2_outputs(7385)) or (layer2_outputs(6349));
    layer3_outputs(3797) <= '1';
    layer3_outputs(3798) <= not(layer2_outputs(1504)) or (layer2_outputs(9341));
    layer3_outputs(3799) <= not((layer2_outputs(2438)) or (layer2_outputs(2163)));
    layer3_outputs(3800) <= not((layer2_outputs(875)) xor (layer2_outputs(2401)));
    layer3_outputs(3801) <= (layer2_outputs(6820)) xor (layer2_outputs(9146));
    layer3_outputs(3802) <= not(layer2_outputs(9966)) or (layer2_outputs(8085));
    layer3_outputs(3803) <= not((layer2_outputs(3049)) xor (layer2_outputs(10161)));
    layer3_outputs(3804) <= layer2_outputs(9566);
    layer3_outputs(3805) <= layer2_outputs(7558);
    layer3_outputs(3806) <= not(layer2_outputs(3360));
    layer3_outputs(3807) <= not(layer2_outputs(3615));
    layer3_outputs(3808) <= layer2_outputs(5257);
    layer3_outputs(3809) <= layer2_outputs(5262);
    layer3_outputs(3810) <= not((layer2_outputs(9155)) or (layer2_outputs(955)));
    layer3_outputs(3811) <= (layer2_outputs(4726)) xor (layer2_outputs(7137));
    layer3_outputs(3812) <= layer2_outputs(2980);
    layer3_outputs(3813) <= not(layer2_outputs(9470));
    layer3_outputs(3814) <= not((layer2_outputs(2295)) xor (layer2_outputs(5563)));
    layer3_outputs(3815) <= not(layer2_outputs(5324));
    layer3_outputs(3816) <= not(layer2_outputs(5389));
    layer3_outputs(3817) <= not(layer2_outputs(5204)) or (layer2_outputs(7860));
    layer3_outputs(3818) <= not((layer2_outputs(4843)) xor (layer2_outputs(8863)));
    layer3_outputs(3819) <= (layer2_outputs(6657)) xor (layer2_outputs(5551));
    layer3_outputs(3820) <= not(layer2_outputs(8105));
    layer3_outputs(3821) <= (layer2_outputs(9895)) or (layer2_outputs(9943));
    layer3_outputs(3822) <= (layer2_outputs(7574)) and not (layer2_outputs(1020));
    layer3_outputs(3823) <= not(layer2_outputs(6211));
    layer3_outputs(3824) <= not(layer2_outputs(8131));
    layer3_outputs(3825) <= (layer2_outputs(9102)) or (layer2_outputs(8010));
    layer3_outputs(3826) <= layer2_outputs(1557);
    layer3_outputs(3827) <= not((layer2_outputs(1422)) xor (layer2_outputs(7972)));
    layer3_outputs(3828) <= not((layer2_outputs(8776)) and (layer2_outputs(50)));
    layer3_outputs(3829) <= layer2_outputs(3549);
    layer3_outputs(3830) <= layer2_outputs(1648);
    layer3_outputs(3831) <= (layer2_outputs(6611)) and (layer2_outputs(6316));
    layer3_outputs(3832) <= '1';
    layer3_outputs(3833) <= (layer2_outputs(4186)) and not (layer2_outputs(614));
    layer3_outputs(3834) <= not(layer2_outputs(451));
    layer3_outputs(3835) <= layer2_outputs(3319);
    layer3_outputs(3836) <= not(layer2_outputs(1763));
    layer3_outputs(3837) <= layer2_outputs(10052);
    layer3_outputs(3838) <= '0';
    layer3_outputs(3839) <= (layer2_outputs(7752)) and not (layer2_outputs(7049));
    layer3_outputs(3840) <= (layer2_outputs(4770)) or (layer2_outputs(6260));
    layer3_outputs(3841) <= not(layer2_outputs(1532));
    layer3_outputs(3842) <= not((layer2_outputs(2105)) or (layer2_outputs(3714)));
    layer3_outputs(3843) <= not(layer2_outputs(3015));
    layer3_outputs(3844) <= not((layer2_outputs(5131)) and (layer2_outputs(3898)));
    layer3_outputs(3845) <= not(layer2_outputs(4793)) or (layer2_outputs(4510));
    layer3_outputs(3846) <= (layer2_outputs(750)) and not (layer2_outputs(4877));
    layer3_outputs(3847) <= layer2_outputs(3879);
    layer3_outputs(3848) <= layer2_outputs(5091);
    layer3_outputs(3849) <= not(layer2_outputs(457));
    layer3_outputs(3850) <= layer2_outputs(5520);
    layer3_outputs(3851) <= layer2_outputs(5973);
    layer3_outputs(3852) <= (layer2_outputs(10167)) and not (layer2_outputs(7660));
    layer3_outputs(3853) <= (layer2_outputs(4904)) and not (layer2_outputs(3616));
    layer3_outputs(3854) <= not((layer2_outputs(5398)) and (layer2_outputs(6908)));
    layer3_outputs(3855) <= (layer2_outputs(9647)) and not (layer2_outputs(5675));
    layer3_outputs(3856) <= not((layer2_outputs(8544)) xor (layer2_outputs(9887)));
    layer3_outputs(3857) <= layer2_outputs(5118);
    layer3_outputs(3858) <= not(layer2_outputs(1514)) or (layer2_outputs(9562));
    layer3_outputs(3859) <= layer2_outputs(6568);
    layer3_outputs(3860) <= layer2_outputs(2973);
    layer3_outputs(3861) <= layer2_outputs(2590);
    layer3_outputs(3862) <= not(layer2_outputs(3016));
    layer3_outputs(3863) <= layer2_outputs(4292);
    layer3_outputs(3864) <= not(layer2_outputs(795));
    layer3_outputs(3865) <= layer2_outputs(7344);
    layer3_outputs(3866) <= not(layer2_outputs(1778)) or (layer2_outputs(6425));
    layer3_outputs(3867) <= (layer2_outputs(10197)) and (layer2_outputs(7798));
    layer3_outputs(3868) <= not(layer2_outputs(2520));
    layer3_outputs(3869) <= (layer2_outputs(1926)) or (layer2_outputs(791));
    layer3_outputs(3870) <= (layer2_outputs(4039)) and not (layer2_outputs(6588));
    layer3_outputs(3871) <= layer2_outputs(6734);
    layer3_outputs(3872) <= (layer2_outputs(383)) and not (layer2_outputs(4245));
    layer3_outputs(3873) <= layer2_outputs(5432);
    layer3_outputs(3874) <= not(layer2_outputs(7917)) or (layer2_outputs(3847));
    layer3_outputs(3875) <= '1';
    layer3_outputs(3876) <= not((layer2_outputs(7916)) and (layer2_outputs(6428)));
    layer3_outputs(3877) <= not(layer2_outputs(3352));
    layer3_outputs(3878) <= layer2_outputs(2464);
    layer3_outputs(3879) <= not(layer2_outputs(1894));
    layer3_outputs(3880) <= '0';
    layer3_outputs(3881) <= (layer2_outputs(3147)) and (layer2_outputs(1820));
    layer3_outputs(3882) <= (layer2_outputs(8589)) or (layer2_outputs(4647));
    layer3_outputs(3883) <= layer2_outputs(6025);
    layer3_outputs(3884) <= layer2_outputs(2222);
    layer3_outputs(3885) <= not(layer2_outputs(2475));
    layer3_outputs(3886) <= layer2_outputs(5758);
    layer3_outputs(3887) <= layer2_outputs(5104);
    layer3_outputs(3888) <= not(layer2_outputs(9405));
    layer3_outputs(3889) <= not(layer2_outputs(340)) or (layer2_outputs(9346));
    layer3_outputs(3890) <= not(layer2_outputs(1643));
    layer3_outputs(3891) <= (layer2_outputs(3627)) and not (layer2_outputs(8133));
    layer3_outputs(3892) <= not(layer2_outputs(9352));
    layer3_outputs(3893) <= layer2_outputs(1396);
    layer3_outputs(3894) <= '1';
    layer3_outputs(3895) <= (layer2_outputs(7540)) or (layer2_outputs(3815));
    layer3_outputs(3896) <= (layer2_outputs(1779)) xor (layer2_outputs(5109));
    layer3_outputs(3897) <= not((layer2_outputs(2235)) and (layer2_outputs(7946)));
    layer3_outputs(3898) <= not(layer2_outputs(4699)) or (layer2_outputs(9285));
    layer3_outputs(3899) <= layer2_outputs(9400);
    layer3_outputs(3900) <= not(layer2_outputs(7547));
    layer3_outputs(3901) <= not(layer2_outputs(8264)) or (layer2_outputs(6497));
    layer3_outputs(3902) <= not(layer2_outputs(4721)) or (layer2_outputs(5597));
    layer3_outputs(3903) <= layer2_outputs(3184);
    layer3_outputs(3904) <= (layer2_outputs(8764)) xor (layer2_outputs(4673));
    layer3_outputs(3905) <= not(layer2_outputs(9851));
    layer3_outputs(3906) <= not(layer2_outputs(7899));
    layer3_outputs(3907) <= not(layer2_outputs(7727)) or (layer2_outputs(22));
    layer3_outputs(3908) <= not(layer2_outputs(7682));
    layer3_outputs(3909) <= (layer2_outputs(7957)) and not (layer2_outputs(2493));
    layer3_outputs(3910) <= not((layer2_outputs(9087)) xor (layer2_outputs(4022)));
    layer3_outputs(3911) <= not(layer2_outputs(3777));
    layer3_outputs(3912) <= not(layer2_outputs(8793));
    layer3_outputs(3913) <= layer2_outputs(5440);
    layer3_outputs(3914) <= not(layer2_outputs(2573)) or (layer2_outputs(7319));
    layer3_outputs(3915) <= layer2_outputs(2111);
    layer3_outputs(3916) <= not(layer2_outputs(2934)) or (layer2_outputs(1421));
    layer3_outputs(3917) <= (layer2_outputs(9152)) and not (layer2_outputs(1360));
    layer3_outputs(3918) <= (layer2_outputs(9788)) and (layer2_outputs(9737));
    layer3_outputs(3919) <= not((layer2_outputs(3931)) xor (layer2_outputs(7867)));
    layer3_outputs(3920) <= not(layer2_outputs(7324));
    layer3_outputs(3921) <= not((layer2_outputs(3442)) or (layer2_outputs(9017)));
    layer3_outputs(3922) <= layer2_outputs(5938);
    layer3_outputs(3923) <= layer2_outputs(914);
    layer3_outputs(3924) <= (layer2_outputs(1115)) and not (layer2_outputs(2503));
    layer3_outputs(3925) <= layer2_outputs(3586);
    layer3_outputs(3926) <= layer2_outputs(9047);
    layer3_outputs(3927) <= layer2_outputs(4960);
    layer3_outputs(3928) <= layer2_outputs(5315);
    layer3_outputs(3929) <= not(layer2_outputs(2831)) or (layer2_outputs(7013));
    layer3_outputs(3930) <= (layer2_outputs(8691)) and not (layer2_outputs(6610));
    layer3_outputs(3931) <= not((layer2_outputs(7018)) or (layer2_outputs(8128)));
    layer3_outputs(3932) <= layer2_outputs(3564);
    layer3_outputs(3933) <= not(layer2_outputs(4422));
    layer3_outputs(3934) <= layer2_outputs(2160);
    layer3_outputs(3935) <= not((layer2_outputs(1902)) xor (layer2_outputs(10048)));
    layer3_outputs(3936) <= not(layer2_outputs(5141));
    layer3_outputs(3937) <= not((layer2_outputs(9125)) xor (layer2_outputs(7858)));
    layer3_outputs(3938) <= not(layer2_outputs(8661));
    layer3_outputs(3939) <= not(layer2_outputs(5166));
    layer3_outputs(3940) <= not((layer2_outputs(8893)) or (layer2_outputs(7446)));
    layer3_outputs(3941) <= '1';
    layer3_outputs(3942) <= not((layer2_outputs(2865)) xor (layer2_outputs(4275)));
    layer3_outputs(3943) <= layer2_outputs(6301);
    layer3_outputs(3944) <= not((layer2_outputs(5079)) xor (layer2_outputs(1863)));
    layer3_outputs(3945) <= not(layer2_outputs(6081));
    layer3_outputs(3946) <= layer2_outputs(9423);
    layer3_outputs(3947) <= '0';
    layer3_outputs(3948) <= not(layer2_outputs(4)) or (layer2_outputs(5649));
    layer3_outputs(3949) <= not((layer2_outputs(9302)) or (layer2_outputs(608)));
    layer3_outputs(3950) <= not((layer2_outputs(9365)) xor (layer2_outputs(3617)));
    layer3_outputs(3951) <= not(layer2_outputs(832));
    layer3_outputs(3952) <= (layer2_outputs(84)) and not (layer2_outputs(1763));
    layer3_outputs(3953) <= not(layer2_outputs(1493)) or (layer2_outputs(3153));
    layer3_outputs(3954) <= not(layer2_outputs(1323));
    layer3_outputs(3955) <= layer2_outputs(9967);
    layer3_outputs(3956) <= layer2_outputs(5164);
    layer3_outputs(3957) <= (layer2_outputs(5767)) or (layer2_outputs(7292));
    layer3_outputs(3958) <= not(layer2_outputs(4146));
    layer3_outputs(3959) <= layer2_outputs(895);
    layer3_outputs(3960) <= layer2_outputs(1959);
    layer3_outputs(3961) <= not(layer2_outputs(6813));
    layer3_outputs(3962) <= layer2_outputs(7120);
    layer3_outputs(3963) <= not(layer2_outputs(4571));
    layer3_outputs(3964) <= not((layer2_outputs(1399)) or (layer2_outputs(1576)));
    layer3_outputs(3965) <= not(layer2_outputs(1669)) or (layer2_outputs(1590));
    layer3_outputs(3966) <= '0';
    layer3_outputs(3967) <= (layer2_outputs(2146)) and not (layer2_outputs(4457));
    layer3_outputs(3968) <= layer2_outputs(1915);
    layer3_outputs(3969) <= '1';
    layer3_outputs(3970) <= not((layer2_outputs(8609)) xor (layer2_outputs(602)));
    layer3_outputs(3971) <= (layer2_outputs(1692)) and (layer2_outputs(415));
    layer3_outputs(3972) <= not(layer2_outputs(8945)) or (layer2_outputs(2259));
    layer3_outputs(3973) <= layer2_outputs(1570);
    layer3_outputs(3974) <= not(layer2_outputs(7516));
    layer3_outputs(3975) <= not(layer2_outputs(7538));
    layer3_outputs(3976) <= not(layer2_outputs(2179)) or (layer2_outputs(425));
    layer3_outputs(3977) <= not(layer2_outputs(2520));
    layer3_outputs(3978) <= not(layer2_outputs(7948)) or (layer2_outputs(5210));
    layer3_outputs(3979) <= (layer2_outputs(1773)) xor (layer2_outputs(1900));
    layer3_outputs(3980) <= layer2_outputs(8789);
    layer3_outputs(3981) <= (layer2_outputs(7800)) xor (layer2_outputs(6301));
    layer3_outputs(3982) <= not(layer2_outputs(7261));
    layer3_outputs(3983) <= not(layer2_outputs(7431)) or (layer2_outputs(2810));
    layer3_outputs(3984) <= '0';
    layer3_outputs(3985) <= not((layer2_outputs(4361)) and (layer2_outputs(477)));
    layer3_outputs(3986) <= not(layer2_outputs(5567));
    layer3_outputs(3987) <= (layer2_outputs(3021)) or (layer2_outputs(6636));
    layer3_outputs(3988) <= layer2_outputs(669);
    layer3_outputs(3989) <= not(layer2_outputs(5481));
    layer3_outputs(3990) <= layer2_outputs(4514);
    layer3_outputs(3991) <= (layer2_outputs(665)) and not (layer2_outputs(5059));
    layer3_outputs(3992) <= not(layer2_outputs(4119)) or (layer2_outputs(3941));
    layer3_outputs(3993) <= layer2_outputs(3737);
    layer3_outputs(3994) <= layer2_outputs(424);
    layer3_outputs(3995) <= (layer2_outputs(2129)) xor (layer2_outputs(7783));
    layer3_outputs(3996) <= not(layer2_outputs(6299));
    layer3_outputs(3997) <= not(layer2_outputs(7080));
    layer3_outputs(3998) <= (layer2_outputs(6467)) and not (layer2_outputs(8621));
    layer3_outputs(3999) <= layer2_outputs(2507);
    layer3_outputs(4000) <= layer2_outputs(1387);
    layer3_outputs(4001) <= not((layer2_outputs(9682)) xor (layer2_outputs(3085)));
    layer3_outputs(4002) <= not(layer2_outputs(2141)) or (layer2_outputs(9114));
    layer3_outputs(4003) <= not(layer2_outputs(7030));
    layer3_outputs(4004) <= (layer2_outputs(2628)) xor (layer2_outputs(7963));
    layer3_outputs(4005) <= layer2_outputs(1826);
    layer3_outputs(4006) <= not(layer2_outputs(3246));
    layer3_outputs(4007) <= (layer2_outputs(8330)) xor (layer2_outputs(341));
    layer3_outputs(4008) <= layer2_outputs(6053);
    layer3_outputs(4009) <= (layer2_outputs(6374)) and not (layer2_outputs(5328));
    layer3_outputs(4010) <= (layer2_outputs(4732)) and not (layer2_outputs(3348));
    layer3_outputs(4011) <= layer2_outputs(5648);
    layer3_outputs(4012) <= not(layer2_outputs(2125)) or (layer2_outputs(3782));
    layer3_outputs(4013) <= not(layer2_outputs(3841));
    layer3_outputs(4014) <= not((layer2_outputs(3678)) and (layer2_outputs(4045)));
    layer3_outputs(4015) <= (layer2_outputs(1498)) xor (layer2_outputs(4553));
    layer3_outputs(4016) <= layer2_outputs(6124);
    layer3_outputs(4017) <= not(layer2_outputs(1735));
    layer3_outputs(4018) <= (layer2_outputs(5027)) xor (layer2_outputs(3439));
    layer3_outputs(4019) <= layer2_outputs(692);
    layer3_outputs(4020) <= (layer2_outputs(3045)) and not (layer2_outputs(6139));
    layer3_outputs(4021) <= not(layer2_outputs(5854)) or (layer2_outputs(2039));
    layer3_outputs(4022) <= not(layer2_outputs(9409)) or (layer2_outputs(3083));
    layer3_outputs(4023) <= '1';
    layer3_outputs(4024) <= not(layer2_outputs(5872));
    layer3_outputs(4025) <= not(layer2_outputs(9431));
    layer3_outputs(4026) <= not(layer2_outputs(203)) or (layer2_outputs(2959));
    layer3_outputs(4027) <= not(layer2_outputs(8273));
    layer3_outputs(4028) <= layer2_outputs(8677);
    layer3_outputs(4029) <= not(layer2_outputs(9811));
    layer3_outputs(4030) <= layer2_outputs(1600);
    layer3_outputs(4031) <= not((layer2_outputs(7031)) or (layer2_outputs(8628)));
    layer3_outputs(4032) <= layer2_outputs(911);
    layer3_outputs(4033) <= not(layer2_outputs(1191)) or (layer2_outputs(446));
    layer3_outputs(4034) <= not((layer2_outputs(5894)) or (layer2_outputs(4021)));
    layer3_outputs(4035) <= not((layer2_outputs(3971)) and (layer2_outputs(1348)));
    layer3_outputs(4036) <= (layer2_outputs(1776)) xor (layer2_outputs(7164));
    layer3_outputs(4037) <= not(layer2_outputs(1916));
    layer3_outputs(4038) <= layer2_outputs(7335);
    layer3_outputs(4039) <= not(layer2_outputs(3908));
    layer3_outputs(4040) <= not((layer2_outputs(6902)) and (layer2_outputs(1574)));
    layer3_outputs(4041) <= not(layer2_outputs(9291));
    layer3_outputs(4042) <= not(layer2_outputs(1830));
    layer3_outputs(4043) <= layer2_outputs(6045);
    layer3_outputs(4044) <= not(layer2_outputs(9244));
    layer3_outputs(4045) <= not((layer2_outputs(3781)) and (layer2_outputs(2903)));
    layer3_outputs(4046) <= layer2_outputs(7407);
    layer3_outputs(4047) <= layer2_outputs(886);
    layer3_outputs(4048) <= not(layer2_outputs(143));
    layer3_outputs(4049) <= not(layer2_outputs(7422));
    layer3_outputs(4050) <= layer2_outputs(9124);
    layer3_outputs(4051) <= not(layer2_outputs(487));
    layer3_outputs(4052) <= layer2_outputs(8369);
    layer3_outputs(4053) <= (layer2_outputs(8684)) xor (layer2_outputs(4280));
    layer3_outputs(4054) <= (layer2_outputs(8469)) and (layer2_outputs(1081));
    layer3_outputs(4055) <= not(layer2_outputs(6015));
    layer3_outputs(4056) <= (layer2_outputs(8096)) xor (layer2_outputs(8118));
    layer3_outputs(4057) <= not(layer2_outputs(5859)) or (layer2_outputs(7978));
    layer3_outputs(4058) <= layer2_outputs(9068);
    layer3_outputs(4059) <= not((layer2_outputs(3754)) xor (layer2_outputs(6208)));
    layer3_outputs(4060) <= not((layer2_outputs(9011)) or (layer2_outputs(5840)));
    layer3_outputs(4061) <= (layer2_outputs(9008)) and not (layer2_outputs(9904));
    layer3_outputs(4062) <= layer2_outputs(9805);
    layer3_outputs(4063) <= (layer2_outputs(5869)) and not (layer2_outputs(2277));
    layer3_outputs(4064) <= not(layer2_outputs(6987)) or (layer2_outputs(9271));
    layer3_outputs(4065) <= layer2_outputs(728);
    layer3_outputs(4066) <= (layer2_outputs(2616)) xor (layer2_outputs(9605));
    layer3_outputs(4067) <= not(layer2_outputs(6520));
    layer3_outputs(4068) <= not((layer2_outputs(576)) or (layer2_outputs(6829)));
    layer3_outputs(4069) <= not((layer2_outputs(2656)) or (layer2_outputs(8238)));
    layer3_outputs(4070) <= not((layer2_outputs(3671)) and (layer2_outputs(1542)));
    layer3_outputs(4071) <= (layer2_outputs(495)) and not (layer2_outputs(6686));
    layer3_outputs(4072) <= not(layer2_outputs(427)) or (layer2_outputs(3804));
    layer3_outputs(4073) <= (layer2_outputs(7804)) and not (layer2_outputs(3014));
    layer3_outputs(4074) <= layer2_outputs(10169);
    layer3_outputs(4075) <= not(layer2_outputs(3390));
    layer3_outputs(4076) <= not((layer2_outputs(9775)) xor (layer2_outputs(2290)));
    layer3_outputs(4077) <= (layer2_outputs(6961)) and (layer2_outputs(2837));
    layer3_outputs(4078) <= (layer2_outputs(9945)) xor (layer2_outputs(5571));
    layer3_outputs(4079) <= (layer2_outputs(1365)) and not (layer2_outputs(4927));
    layer3_outputs(4080) <= layer2_outputs(1508);
    layer3_outputs(4081) <= not((layer2_outputs(2403)) and (layer2_outputs(1731)));
    layer3_outputs(4082) <= (layer2_outputs(4454)) and not (layer2_outputs(7216));
    layer3_outputs(4083) <= layer2_outputs(9868);
    layer3_outputs(4084) <= layer2_outputs(4363);
    layer3_outputs(4085) <= not(layer2_outputs(6018)) or (layer2_outputs(9710));
    layer3_outputs(4086) <= not((layer2_outputs(4058)) or (layer2_outputs(8132)));
    layer3_outputs(4087) <= not(layer2_outputs(853));
    layer3_outputs(4088) <= not(layer2_outputs(4178));
    layer3_outputs(4089) <= not(layer2_outputs(6609));
    layer3_outputs(4090) <= not((layer2_outputs(2478)) or (layer2_outputs(9753)));
    layer3_outputs(4091) <= not((layer2_outputs(2543)) xor (layer2_outputs(10058)));
    layer3_outputs(4092) <= (layer2_outputs(1961)) and not (layer2_outputs(6273));
    layer3_outputs(4093) <= (layer2_outputs(8314)) and not (layer2_outputs(567));
    layer3_outputs(4094) <= not(layer2_outputs(5766)) or (layer2_outputs(6219));
    layer3_outputs(4095) <= not(layer2_outputs(7338));
    layer3_outputs(4096) <= not(layer2_outputs(1735));
    layer3_outputs(4097) <= (layer2_outputs(8038)) and (layer2_outputs(9646));
    layer3_outputs(4098) <= not(layer2_outputs(7239));
    layer3_outputs(4099) <= not(layer2_outputs(2711));
    layer3_outputs(4100) <= layer2_outputs(8100);
    layer3_outputs(4101) <= layer2_outputs(2431);
    layer3_outputs(4102) <= not(layer2_outputs(4261));
    layer3_outputs(4103) <= layer2_outputs(3157);
    layer3_outputs(4104) <= layer2_outputs(433);
    layer3_outputs(4105) <= layer2_outputs(5230);
    layer3_outputs(4106) <= not((layer2_outputs(3836)) or (layer2_outputs(9977)));
    layer3_outputs(4107) <= (layer2_outputs(6894)) xor (layer2_outputs(1831));
    layer3_outputs(4108) <= not(layer2_outputs(5498));
    layer3_outputs(4109) <= '1';
    layer3_outputs(4110) <= not(layer2_outputs(4116));
    layer3_outputs(4111) <= (layer2_outputs(4806)) or (layer2_outputs(8590));
    layer3_outputs(4112) <= not(layer2_outputs(5353));
    layer3_outputs(4113) <= (layer2_outputs(653)) and (layer2_outputs(9025));
    layer3_outputs(4114) <= layer2_outputs(2818);
    layer3_outputs(4115) <= '1';
    layer3_outputs(4116) <= layer2_outputs(7705);
    layer3_outputs(4117) <= not(layer2_outputs(4836));
    layer3_outputs(4118) <= layer2_outputs(2831);
    layer3_outputs(4119) <= not((layer2_outputs(8752)) or (layer2_outputs(9440)));
    layer3_outputs(4120) <= layer2_outputs(1676);
    layer3_outputs(4121) <= not((layer2_outputs(4980)) and (layer2_outputs(7509)));
    layer3_outputs(4122) <= layer2_outputs(6278);
    layer3_outputs(4123) <= not(layer2_outputs(9399));
    layer3_outputs(4124) <= (layer2_outputs(4885)) and (layer2_outputs(4697));
    layer3_outputs(4125) <= not(layer2_outputs(1707));
    layer3_outputs(4126) <= layer2_outputs(8402);
    layer3_outputs(4127) <= layer2_outputs(9996);
    layer3_outputs(4128) <= not(layer2_outputs(8249));
    layer3_outputs(4129) <= '0';
    layer3_outputs(4130) <= not(layer2_outputs(6351));
    layer3_outputs(4131) <= not((layer2_outputs(4995)) or (layer2_outputs(1295)));
    layer3_outputs(4132) <= not(layer2_outputs(6140));
    layer3_outputs(4133) <= layer2_outputs(9982);
    layer3_outputs(4134) <= not(layer2_outputs(8978));
    layer3_outputs(4135) <= layer2_outputs(3429);
    layer3_outputs(4136) <= (layer2_outputs(7468)) and not (layer2_outputs(6859));
    layer3_outputs(4137) <= (layer2_outputs(5846)) and not (layer2_outputs(4474));
    layer3_outputs(4138) <= not((layer2_outputs(7917)) and (layer2_outputs(2791)));
    layer3_outputs(4139) <= not(layer2_outputs(3686));
    layer3_outputs(4140) <= layer2_outputs(857);
    layer3_outputs(4141) <= layer2_outputs(1539);
    layer3_outputs(4142) <= layer2_outputs(3637);
    layer3_outputs(4143) <= not(layer2_outputs(1360));
    layer3_outputs(4144) <= (layer2_outputs(9007)) and (layer2_outputs(718));
    layer3_outputs(4145) <= not(layer2_outputs(5501));
    layer3_outputs(4146) <= not(layer2_outputs(4433));
    layer3_outputs(4147) <= '1';
    layer3_outputs(4148) <= layer2_outputs(9566);
    layer3_outputs(4149) <= layer2_outputs(1007);
    layer3_outputs(4150) <= '1';
    layer3_outputs(4151) <= (layer2_outputs(6303)) and not (layer2_outputs(5285));
    layer3_outputs(4152) <= (layer2_outputs(7678)) and (layer2_outputs(221));
    layer3_outputs(4153) <= (layer2_outputs(6925)) xor (layer2_outputs(8051));
    layer3_outputs(4154) <= not(layer2_outputs(9658));
    layer3_outputs(4155) <= layer2_outputs(5835);
    layer3_outputs(4156) <= '1';
    layer3_outputs(4157) <= (layer2_outputs(9744)) xor (layer2_outputs(1875));
    layer3_outputs(4158) <= (layer2_outputs(8419)) and (layer2_outputs(2385));
    layer3_outputs(4159) <= (layer2_outputs(4756)) xor (layer2_outputs(49));
    layer3_outputs(4160) <= not(layer2_outputs(2419)) or (layer2_outputs(3805));
    layer3_outputs(4161) <= not(layer2_outputs(8546));
    layer3_outputs(4162) <= layer2_outputs(5716);
    layer3_outputs(4163) <= not(layer2_outputs(7615)) or (layer2_outputs(3972));
    layer3_outputs(4164) <= (layer2_outputs(6170)) and (layer2_outputs(9621));
    layer3_outputs(4165) <= not(layer2_outputs(7584)) or (layer2_outputs(6446));
    layer3_outputs(4166) <= (layer2_outputs(9600)) xor (layer2_outputs(9752));
    layer3_outputs(4167) <= not((layer2_outputs(5169)) xor (layer2_outputs(4064)));
    layer3_outputs(4168) <= layer2_outputs(5038);
    layer3_outputs(4169) <= not(layer2_outputs(2731));
    layer3_outputs(4170) <= (layer2_outputs(4755)) and not (layer2_outputs(8632));
    layer3_outputs(4171) <= (layer2_outputs(5196)) and not (layer2_outputs(6528));
    layer3_outputs(4172) <= (layer2_outputs(4554)) or (layer2_outputs(4515));
    layer3_outputs(4173) <= layer2_outputs(252);
    layer3_outputs(4174) <= not(layer2_outputs(226));
    layer3_outputs(4175) <= layer2_outputs(3769);
    layer3_outputs(4176) <= (layer2_outputs(6878)) or (layer2_outputs(1116));
    layer3_outputs(4177) <= '0';
    layer3_outputs(4178) <= not(layer2_outputs(5249));
    layer3_outputs(4179) <= (layer2_outputs(1332)) and (layer2_outputs(1592));
    layer3_outputs(4180) <= layer2_outputs(5369);
    layer3_outputs(4181) <= layer2_outputs(5922);
    layer3_outputs(4182) <= not((layer2_outputs(85)) or (layer2_outputs(2445)));
    layer3_outputs(4183) <= not(layer2_outputs(8756));
    layer3_outputs(4184) <= layer2_outputs(3932);
    layer3_outputs(4185) <= not((layer2_outputs(10154)) xor (layer2_outputs(2991)));
    layer3_outputs(4186) <= layer2_outputs(7849);
    layer3_outputs(4187) <= layer2_outputs(4615);
    layer3_outputs(4188) <= not(layer2_outputs(6165)) or (layer2_outputs(9807));
    layer3_outputs(4189) <= '1';
    layer3_outputs(4190) <= not(layer2_outputs(913)) or (layer2_outputs(3165));
    layer3_outputs(4191) <= not(layer2_outputs(5277)) or (layer2_outputs(6484));
    layer3_outputs(4192) <= (layer2_outputs(4921)) and not (layer2_outputs(3591));
    layer3_outputs(4193) <= not(layer2_outputs(5852));
    layer3_outputs(4194) <= layer2_outputs(6534);
    layer3_outputs(4195) <= (layer2_outputs(8555)) and not (layer2_outputs(435));
    layer3_outputs(4196) <= (layer2_outputs(5591)) xor (layer2_outputs(7876));
    layer3_outputs(4197) <= layer2_outputs(3109);
    layer3_outputs(4198) <= (layer2_outputs(5030)) xor (layer2_outputs(5703));
    layer3_outputs(4199) <= not(layer2_outputs(4638));
    layer3_outputs(4200) <= (layer2_outputs(7577)) and not (layer2_outputs(5876));
    layer3_outputs(4201) <= layer2_outputs(7087);
    layer3_outputs(4202) <= layer2_outputs(5280);
    layer3_outputs(4203) <= (layer2_outputs(6574)) and (layer2_outputs(4217));
    layer3_outputs(4204) <= not(layer2_outputs(1398));
    layer3_outputs(4205) <= (layer2_outputs(1287)) or (layer2_outputs(9143));
    layer3_outputs(4206) <= not((layer2_outputs(5181)) and (layer2_outputs(9220)));
    layer3_outputs(4207) <= not((layer2_outputs(9342)) or (layer2_outputs(1683)));
    layer3_outputs(4208) <= layer2_outputs(2861);
    layer3_outputs(4209) <= not(layer2_outputs(1207)) or (layer2_outputs(2965));
    layer3_outputs(4210) <= (layer2_outputs(7244)) or (layer2_outputs(5732));
    layer3_outputs(4211) <= (layer2_outputs(10073)) or (layer2_outputs(518));
    layer3_outputs(4212) <= '1';
    layer3_outputs(4213) <= layer2_outputs(8055);
    layer3_outputs(4214) <= (layer2_outputs(5920)) xor (layer2_outputs(914));
    layer3_outputs(4215) <= layer2_outputs(9859);
    layer3_outputs(4216) <= not((layer2_outputs(1197)) xor (layer2_outputs(240)));
    layer3_outputs(4217) <= not((layer2_outputs(9518)) xor (layer2_outputs(4976)));
    layer3_outputs(4218) <= not(layer2_outputs(2208));
    layer3_outputs(4219) <= not(layer2_outputs(1003)) or (layer2_outputs(8290));
    layer3_outputs(4220) <= not(layer2_outputs(3687));
    layer3_outputs(4221) <= (layer2_outputs(4675)) or (layer2_outputs(9850));
    layer3_outputs(4222) <= (layer2_outputs(3020)) and not (layer2_outputs(9338));
    layer3_outputs(4223) <= layer2_outputs(9021);
    layer3_outputs(4224) <= layer2_outputs(1887);
    layer3_outputs(4225) <= (layer2_outputs(2969)) xor (layer2_outputs(1659));
    layer3_outputs(4226) <= layer2_outputs(8755);
    layer3_outputs(4227) <= not(layer2_outputs(8190)) or (layer2_outputs(7735));
    layer3_outputs(4228) <= layer2_outputs(1858);
    layer3_outputs(4229) <= (layer2_outputs(4902)) and (layer2_outputs(749));
    layer3_outputs(4230) <= layer2_outputs(6496);
    layer3_outputs(4231) <= (layer2_outputs(694)) or (layer2_outputs(8160));
    layer3_outputs(4232) <= not(layer2_outputs(6548)) or (layer2_outputs(1038));
    layer3_outputs(4233) <= layer2_outputs(5544);
    layer3_outputs(4234) <= layer2_outputs(8480);
    layer3_outputs(4235) <= layer2_outputs(4438);
    layer3_outputs(4236) <= layer2_outputs(5417);
    layer3_outputs(4237) <= layer2_outputs(2089);
    layer3_outputs(4238) <= layer2_outputs(5057);
    layer3_outputs(4239) <= not((layer2_outputs(5185)) xor (layer2_outputs(9032)));
    layer3_outputs(4240) <= not(layer2_outputs(5269));
    layer3_outputs(4241) <= not(layer2_outputs(3245));
    layer3_outputs(4242) <= '1';
    layer3_outputs(4243) <= '0';
    layer3_outputs(4244) <= (layer2_outputs(8089)) or (layer2_outputs(1614));
    layer3_outputs(4245) <= layer2_outputs(8911);
    layer3_outputs(4246) <= not((layer2_outputs(4547)) xor (layer2_outputs(944)));
    layer3_outputs(4247) <= layer2_outputs(6465);
    layer3_outputs(4248) <= layer2_outputs(1056);
    layer3_outputs(4249) <= (layer2_outputs(1257)) and not (layer2_outputs(1869));
    layer3_outputs(4250) <= not(layer2_outputs(6410));
    layer3_outputs(4251) <= not(layer2_outputs(9956)) or (layer2_outputs(3970));
    layer3_outputs(4252) <= not(layer2_outputs(5627));
    layer3_outputs(4253) <= not(layer2_outputs(8176));
    layer3_outputs(4254) <= (layer2_outputs(4719)) or (layer2_outputs(9430));
    layer3_outputs(4255) <= layer2_outputs(2481);
    layer3_outputs(4256) <= not((layer2_outputs(9322)) and (layer2_outputs(5696)));
    layer3_outputs(4257) <= (layer2_outputs(544)) xor (layer2_outputs(8850));
    layer3_outputs(4258) <= layer2_outputs(9457);
    layer3_outputs(4259) <= not(layer2_outputs(477));
    layer3_outputs(4260) <= '0';
    layer3_outputs(4261) <= (layer2_outputs(732)) and not (layer2_outputs(8460));
    layer3_outputs(4262) <= layer2_outputs(5078);
    layer3_outputs(4263) <= not(layer2_outputs(4155));
    layer3_outputs(4264) <= layer2_outputs(905);
    layer3_outputs(4265) <= not(layer2_outputs(8954));
    layer3_outputs(4266) <= not(layer2_outputs(8737)) or (layer2_outputs(8885));
    layer3_outputs(4267) <= not(layer2_outputs(6159)) or (layer2_outputs(5503));
    layer3_outputs(4268) <= not(layer2_outputs(6746));
    layer3_outputs(4269) <= not((layer2_outputs(2290)) and (layer2_outputs(961)));
    layer3_outputs(4270) <= (layer2_outputs(9380)) and (layer2_outputs(9865));
    layer3_outputs(4271) <= layer2_outputs(9594);
    layer3_outputs(4272) <= layer2_outputs(415);
    layer3_outputs(4273) <= not(layer2_outputs(4574));
    layer3_outputs(4274) <= layer2_outputs(3060);
    layer3_outputs(4275) <= not(layer2_outputs(4799));
    layer3_outputs(4276) <= layer2_outputs(4136);
    layer3_outputs(4277) <= not(layer2_outputs(2279));
    layer3_outputs(4278) <= not(layer2_outputs(1128)) or (layer2_outputs(6514));
    layer3_outputs(4279) <= (layer2_outputs(5680)) or (layer2_outputs(1645));
    layer3_outputs(4280) <= not((layer2_outputs(9296)) xor (layer2_outputs(3542)));
    layer3_outputs(4281) <= not(layer2_outputs(4268));
    layer3_outputs(4282) <= not((layer2_outputs(2566)) and (layer2_outputs(6127)));
    layer3_outputs(4283) <= (layer2_outputs(3821)) and not (layer2_outputs(4125));
    layer3_outputs(4284) <= layer2_outputs(2154);
    layer3_outputs(4285) <= not((layer2_outputs(2985)) xor (layer2_outputs(9851)));
    layer3_outputs(4286) <= (layer2_outputs(659)) xor (layer2_outputs(1637));
    layer3_outputs(4287) <= '1';
    layer3_outputs(4288) <= not((layer2_outputs(5849)) or (layer2_outputs(8539)));
    layer3_outputs(4289) <= layer2_outputs(583);
    layer3_outputs(4290) <= (layer2_outputs(9608)) and not (layer2_outputs(4301));
    layer3_outputs(4291) <= (layer2_outputs(310)) and (layer2_outputs(1696));
    layer3_outputs(4292) <= not(layer2_outputs(4059));
    layer3_outputs(4293) <= not((layer2_outputs(9870)) xor (layer2_outputs(8072)));
    layer3_outputs(4294) <= not(layer2_outputs(1467)) or (layer2_outputs(8781));
    layer3_outputs(4295) <= not(layer2_outputs(7627)) or (layer2_outputs(3464));
    layer3_outputs(4296) <= not(layer2_outputs(3806)) or (layer2_outputs(7137));
    layer3_outputs(4297) <= not(layer2_outputs(1285)) or (layer2_outputs(3909));
    layer3_outputs(4298) <= not((layer2_outputs(2028)) xor (layer2_outputs(8891)));
    layer3_outputs(4299) <= layer2_outputs(750);
    layer3_outputs(4300) <= layer2_outputs(5227);
    layer3_outputs(4301) <= layer2_outputs(9237);
    layer3_outputs(4302) <= not(layer2_outputs(2887)) or (layer2_outputs(119));
    layer3_outputs(4303) <= layer2_outputs(6857);
    layer3_outputs(4304) <= (layer2_outputs(4917)) and not (layer2_outputs(4211));
    layer3_outputs(4305) <= not(layer2_outputs(3281));
    layer3_outputs(4306) <= layer2_outputs(5543);
    layer3_outputs(4307) <= not(layer2_outputs(3858));
    layer3_outputs(4308) <= layer2_outputs(3032);
    layer3_outputs(4309) <= (layer2_outputs(516)) xor (layer2_outputs(6993));
    layer3_outputs(4310) <= layer2_outputs(4570);
    layer3_outputs(4311) <= (layer2_outputs(4407)) and not (layer2_outputs(9419));
    layer3_outputs(4312) <= not(layer2_outputs(4961)) or (layer2_outputs(9014));
    layer3_outputs(4313) <= layer2_outputs(5668);
    layer3_outputs(4314) <= layer2_outputs(6464);
    layer3_outputs(4315) <= layer2_outputs(3932);
    layer3_outputs(4316) <= (layer2_outputs(5888)) and not (layer2_outputs(1115));
    layer3_outputs(4317) <= not(layer2_outputs(7910)) or (layer2_outputs(1841));
    layer3_outputs(4318) <= layer2_outputs(9554);
    layer3_outputs(4319) <= (layer2_outputs(7214)) xor (layer2_outputs(10136));
    layer3_outputs(4320) <= not(layer2_outputs(5503));
    layer3_outputs(4321) <= (layer2_outputs(3564)) and not (layer2_outputs(1273));
    layer3_outputs(4322) <= '0';
    layer3_outputs(4323) <= layer2_outputs(594);
    layer3_outputs(4324) <= not(layer2_outputs(6503));
    layer3_outputs(4325) <= not((layer2_outputs(7441)) and (layer2_outputs(8669)));
    layer3_outputs(4326) <= (layer2_outputs(4623)) and not (layer2_outputs(7457));
    layer3_outputs(4327) <= not(layer2_outputs(4468));
    layer3_outputs(4328) <= not((layer2_outputs(4839)) xor (layer2_outputs(8013)));
    layer3_outputs(4329) <= not(layer2_outputs(3273));
    layer3_outputs(4330) <= layer2_outputs(5003);
    layer3_outputs(4331) <= layer2_outputs(4559);
    layer3_outputs(4332) <= layer2_outputs(1974);
    layer3_outputs(4333) <= '1';
    layer3_outputs(4334) <= (layer2_outputs(9181)) xor (layer2_outputs(6105));
    layer3_outputs(4335) <= not(layer2_outputs(1358));
    layer3_outputs(4336) <= not(layer2_outputs(5183)) or (layer2_outputs(1218));
    layer3_outputs(4337) <= '0';
    layer3_outputs(4338) <= not((layer2_outputs(7738)) xor (layer2_outputs(9168)));
    layer3_outputs(4339) <= layer2_outputs(6987);
    layer3_outputs(4340) <= not(layer2_outputs(7343));
    layer3_outputs(4341) <= not((layer2_outputs(9582)) xor (layer2_outputs(7912)));
    layer3_outputs(4342) <= not(layer2_outputs(192)) or (layer2_outputs(4040));
    layer3_outputs(4343) <= (layer2_outputs(2404)) and (layer2_outputs(1461));
    layer3_outputs(4344) <= layer2_outputs(9540);
    layer3_outputs(4345) <= (layer2_outputs(6939)) or (layer2_outputs(1569));
    layer3_outputs(4346) <= layer2_outputs(4000);
    layer3_outputs(4347) <= (layer2_outputs(3442)) and not (layer2_outputs(650));
    layer3_outputs(4348) <= not(layer2_outputs(9171));
    layer3_outputs(4349) <= (layer2_outputs(5523)) and (layer2_outputs(7824));
    layer3_outputs(4350) <= not(layer2_outputs(1644));
    layer3_outputs(4351) <= layer2_outputs(4383);
    layer3_outputs(4352) <= (layer2_outputs(6295)) and not (layer2_outputs(844));
    layer3_outputs(4353) <= (layer2_outputs(486)) and (layer2_outputs(8914));
    layer3_outputs(4354) <= not(layer2_outputs(4520));
    layer3_outputs(4355) <= layer2_outputs(9495);
    layer3_outputs(4356) <= not(layer2_outputs(947)) or (layer2_outputs(6854));
    layer3_outputs(4357) <= not(layer2_outputs(2913));
    layer3_outputs(4358) <= layer2_outputs(113);
    layer3_outputs(4359) <= not(layer2_outputs(7413));
    layer3_outputs(4360) <= not(layer2_outputs(9777));
    layer3_outputs(4361) <= layer2_outputs(6358);
    layer3_outputs(4362) <= not((layer2_outputs(5071)) and (layer2_outputs(8851)));
    layer3_outputs(4363) <= layer2_outputs(877);
    layer3_outputs(4364) <= not(layer2_outputs(456));
    layer3_outputs(4365) <= layer2_outputs(5428);
    layer3_outputs(4366) <= not(layer2_outputs(2672)) or (layer2_outputs(8647));
    layer3_outputs(4367) <= layer2_outputs(7101);
    layer3_outputs(4368) <= not(layer2_outputs(10184));
    layer3_outputs(4369) <= layer2_outputs(1552);
    layer3_outputs(4370) <= (layer2_outputs(7485)) xor (layer2_outputs(5572));
    layer3_outputs(4371) <= not(layer2_outputs(6710));
    layer3_outputs(4372) <= not(layer2_outputs(7503));
    layer3_outputs(4373) <= layer2_outputs(3600);
    layer3_outputs(4374) <= (layer2_outputs(5879)) or (layer2_outputs(5122));
    layer3_outputs(4375) <= (layer2_outputs(1705)) and not (layer2_outputs(4121));
    layer3_outputs(4376) <= (layer2_outputs(4868)) and not (layer2_outputs(3213));
    layer3_outputs(4377) <= layer2_outputs(3075);
    layer3_outputs(4378) <= not(layer2_outputs(6226));
    layer3_outputs(4379) <= not((layer2_outputs(8391)) xor (layer2_outputs(8250)));
    layer3_outputs(4380) <= not(layer2_outputs(2545)) or (layer2_outputs(9023));
    layer3_outputs(4381) <= not(layer2_outputs(4978)) or (layer2_outputs(786));
    layer3_outputs(4382) <= (layer2_outputs(3869)) and not (layer2_outputs(4021));
    layer3_outputs(4383) <= layer2_outputs(9443);
    layer3_outputs(4384) <= layer2_outputs(9840);
    layer3_outputs(4385) <= '1';
    layer3_outputs(4386) <= (layer2_outputs(6567)) or (layer2_outputs(1086));
    layer3_outputs(4387) <= not((layer2_outputs(2395)) and (layer2_outputs(665)));
    layer3_outputs(4388) <= layer2_outputs(9964);
    layer3_outputs(4389) <= (layer2_outputs(176)) and not (layer2_outputs(3328));
    layer3_outputs(4390) <= not(layer2_outputs(9627));
    layer3_outputs(4391) <= layer2_outputs(4815);
    layer3_outputs(4392) <= layer2_outputs(9575);
    layer3_outputs(4393) <= layer2_outputs(2162);
    layer3_outputs(4394) <= layer2_outputs(7329);
    layer3_outputs(4395) <= not(layer2_outputs(10108));
    layer3_outputs(4396) <= not((layer2_outputs(9303)) and (layer2_outputs(8413)));
    layer3_outputs(4397) <= not((layer2_outputs(4949)) or (layer2_outputs(3975)));
    layer3_outputs(4398) <= not(layer2_outputs(7476));
    layer3_outputs(4399) <= (layer2_outputs(5463)) and not (layer2_outputs(9825));
    layer3_outputs(4400) <= (layer2_outputs(9191)) and not (layer2_outputs(4829));
    layer3_outputs(4401) <= not(layer2_outputs(3272));
    layer3_outputs(4402) <= not(layer2_outputs(4525));
    layer3_outputs(4403) <= not(layer2_outputs(1322));
    layer3_outputs(4404) <= (layer2_outputs(4408)) or (layer2_outputs(5576));
    layer3_outputs(4405) <= (layer2_outputs(7535)) or (layer2_outputs(9513));
    layer3_outputs(4406) <= not((layer2_outputs(1488)) or (layer2_outputs(8566)));
    layer3_outputs(4407) <= (layer2_outputs(10205)) and not (layer2_outputs(2349));
    layer3_outputs(4408) <= layer2_outputs(9140);
    layer3_outputs(4409) <= not(layer2_outputs(9614)) or (layer2_outputs(3279));
    layer3_outputs(4410) <= layer2_outputs(5838);
    layer3_outputs(4411) <= layer2_outputs(115);
    layer3_outputs(4412) <= not(layer2_outputs(9557));
    layer3_outputs(4413) <= (layer2_outputs(2576)) and not (layer2_outputs(6581));
    layer3_outputs(4414) <= (layer2_outputs(9056)) and not (layer2_outputs(582));
    layer3_outputs(4415) <= not(layer2_outputs(3842));
    layer3_outputs(4416) <= layer2_outputs(8829);
    layer3_outputs(4417) <= layer2_outputs(5654);
    layer3_outputs(4418) <= (layer2_outputs(9702)) and not (layer2_outputs(5636));
    layer3_outputs(4419) <= (layer2_outputs(3965)) and not (layer2_outputs(860));
    layer3_outputs(4420) <= (layer2_outputs(9546)) and not (layer2_outputs(3022));
    layer3_outputs(4421) <= (layer2_outputs(3614)) and not (layer2_outputs(1823));
    layer3_outputs(4422) <= not((layer2_outputs(2443)) or (layer2_outputs(8183)));
    layer3_outputs(4423) <= (layer2_outputs(4830)) and (layer2_outputs(4458));
    layer3_outputs(4424) <= (layer2_outputs(4583)) or (layer2_outputs(9637));
    layer3_outputs(4425) <= '1';
    layer3_outputs(4426) <= (layer2_outputs(8327)) or (layer2_outputs(4950));
    layer3_outputs(4427) <= layer2_outputs(3684);
    layer3_outputs(4428) <= not(layer2_outputs(1743));
    layer3_outputs(4429) <= not(layer2_outputs(2123));
    layer3_outputs(4430) <= not(layer2_outputs(1390));
    layer3_outputs(4431) <= (layer2_outputs(9524)) and not (layer2_outputs(1741));
    layer3_outputs(4432) <= not(layer2_outputs(1663));
    layer3_outputs(4433) <= layer2_outputs(7799);
    layer3_outputs(4434) <= not((layer2_outputs(2216)) xor (layer2_outputs(1085)));
    layer3_outputs(4435) <= not(layer2_outputs(2374));
    layer3_outputs(4436) <= not(layer2_outputs(8996));
    layer3_outputs(4437) <= layer2_outputs(4019);
    layer3_outputs(4438) <= not((layer2_outputs(2737)) xor (layer2_outputs(9160)));
    layer3_outputs(4439) <= not(layer2_outputs(4388));
    layer3_outputs(4440) <= not(layer2_outputs(8553));
    layer3_outputs(4441) <= not((layer2_outputs(103)) or (layer2_outputs(8858)));
    layer3_outputs(4442) <= (layer2_outputs(178)) xor (layer2_outputs(8035));
    layer3_outputs(4443) <= layer2_outputs(823);
    layer3_outputs(4444) <= not(layer2_outputs(8219));
    layer3_outputs(4445) <= not((layer2_outputs(291)) and (layer2_outputs(8227)));
    layer3_outputs(4446) <= not(layer2_outputs(8860));
    layer3_outputs(4447) <= layer2_outputs(4086);
    layer3_outputs(4448) <= (layer2_outputs(412)) or (layer2_outputs(6358));
    layer3_outputs(4449) <= not(layer2_outputs(2339));
    layer3_outputs(4450) <= (layer2_outputs(4890)) and not (layer2_outputs(9292));
    layer3_outputs(4451) <= '1';
    layer3_outputs(4452) <= (layer2_outputs(8614)) or (layer2_outputs(3571));
    layer3_outputs(4453) <= (layer2_outputs(5882)) xor (layer2_outputs(748));
    layer3_outputs(4454) <= layer2_outputs(7082);
    layer3_outputs(4455) <= not((layer2_outputs(3768)) and (layer2_outputs(3865)));
    layer3_outputs(4456) <= not((layer2_outputs(2938)) and (layer2_outputs(6126)));
    layer3_outputs(4457) <= (layer2_outputs(8121)) and not (layer2_outputs(9053));
    layer3_outputs(4458) <= layer2_outputs(9870);
    layer3_outputs(4459) <= not(layer2_outputs(10232));
    layer3_outputs(4460) <= not((layer2_outputs(7675)) xor (layer2_outputs(3735)));
    layer3_outputs(4461) <= not((layer2_outputs(1282)) or (layer2_outputs(6004)));
    layer3_outputs(4462) <= not(layer2_outputs(3300)) or (layer2_outputs(1341));
    layer3_outputs(4463) <= layer2_outputs(7530);
    layer3_outputs(4464) <= (layer2_outputs(5657)) and (layer2_outputs(4535));
    layer3_outputs(4465) <= not((layer2_outputs(9535)) xor (layer2_outputs(3713)));
    layer3_outputs(4466) <= layer2_outputs(5247);
    layer3_outputs(4467) <= layer2_outputs(4761);
    layer3_outputs(4468) <= not(layer2_outputs(9606));
    layer3_outputs(4469) <= not(layer2_outputs(4473)) or (layer2_outputs(2723));
    layer3_outputs(4470) <= not(layer2_outputs(6414));
    layer3_outputs(4471) <= (layer2_outputs(4873)) xor (layer2_outputs(5094));
    layer3_outputs(4472) <= not(layer2_outputs(7263));
    layer3_outputs(4473) <= not(layer2_outputs(126));
    layer3_outputs(4474) <= layer2_outputs(3695);
    layer3_outputs(4475) <= (layer2_outputs(9848)) and not (layer2_outputs(4748));
    layer3_outputs(4476) <= layer2_outputs(2291);
    layer3_outputs(4477) <= not(layer2_outputs(8165)) or (layer2_outputs(5976));
    layer3_outputs(4478) <= (layer2_outputs(4835)) and not (layer2_outputs(8659));
    layer3_outputs(4479) <= not(layer2_outputs(7026)) or (layer2_outputs(5140));
    layer3_outputs(4480) <= '1';
    layer3_outputs(4481) <= layer2_outputs(1252);
    layer3_outputs(4482) <= (layer2_outputs(6182)) and not (layer2_outputs(438));
    layer3_outputs(4483) <= not((layer2_outputs(9885)) xor (layer2_outputs(2595)));
    layer3_outputs(4484) <= layer2_outputs(9446);
    layer3_outputs(4485) <= (layer2_outputs(9251)) and (layer2_outputs(1242));
    layer3_outputs(4486) <= not(layer2_outputs(9897));
    layer3_outputs(4487) <= not(layer2_outputs(3944));
    layer3_outputs(4488) <= layer2_outputs(1498);
    layer3_outputs(4489) <= not(layer2_outputs(3875));
    layer3_outputs(4490) <= layer2_outputs(5546);
    layer3_outputs(4491) <= not(layer2_outputs(4505));
    layer3_outputs(4492) <= not(layer2_outputs(570));
    layer3_outputs(4493) <= not((layer2_outputs(8453)) xor (layer2_outputs(5409)));
    layer3_outputs(4494) <= not(layer2_outputs(6244));
    layer3_outputs(4495) <= not((layer2_outputs(6781)) xor (layer2_outputs(2099)));
    layer3_outputs(4496) <= not(layer2_outputs(6390)) or (layer2_outputs(7561));
    layer3_outputs(4497) <= not(layer2_outputs(5318));
    layer3_outputs(4498) <= not(layer2_outputs(4395));
    layer3_outputs(4499) <= layer2_outputs(9290);
    layer3_outputs(4500) <= not(layer2_outputs(10138));
    layer3_outputs(4501) <= layer2_outputs(3275);
    layer3_outputs(4502) <= not((layer2_outputs(8309)) xor (layer2_outputs(8307)));
    layer3_outputs(4503) <= not(layer2_outputs(5040)) or (layer2_outputs(8718));
    layer3_outputs(4504) <= not(layer2_outputs(8868));
    layer3_outputs(4505) <= (layer2_outputs(2611)) and not (layer2_outputs(3966));
    layer3_outputs(4506) <= not((layer2_outputs(6885)) and (layer2_outputs(1215)));
    layer3_outputs(4507) <= layer2_outputs(4085);
    layer3_outputs(4508) <= not((layer2_outputs(6588)) xor (layer2_outputs(8999)));
    layer3_outputs(4509) <= (layer2_outputs(8120)) and (layer2_outputs(574));
    layer3_outputs(4510) <= not(layer2_outputs(107));
    layer3_outputs(4511) <= not((layer2_outputs(8066)) and (layer2_outputs(957)));
    layer3_outputs(4512) <= '1';
    layer3_outputs(4513) <= (layer2_outputs(10088)) and not (layer2_outputs(584));
    layer3_outputs(4514) <= not(layer2_outputs(8335)) or (layer2_outputs(9355));
    layer3_outputs(4515) <= (layer2_outputs(5225)) xor (layer2_outputs(1728));
    layer3_outputs(4516) <= not(layer2_outputs(1672)) or (layer2_outputs(9368));
    layer3_outputs(4517) <= (layer2_outputs(3654)) and not (layer2_outputs(2867));
    layer3_outputs(4518) <= not(layer2_outputs(156));
    layer3_outputs(4519) <= not(layer2_outputs(8519));
    layer3_outputs(4520) <= '1';
    layer3_outputs(4521) <= (layer2_outputs(9826)) and not (layer2_outputs(3530));
    layer3_outputs(4522) <= layer2_outputs(3718);
    layer3_outputs(4523) <= not((layer2_outputs(4493)) xor (layer2_outputs(10044)));
    layer3_outputs(4524) <= not(layer2_outputs(6250));
    layer3_outputs(4525) <= not((layer2_outputs(846)) or (layer2_outputs(7636)));
    layer3_outputs(4526) <= layer2_outputs(3015);
    layer3_outputs(4527) <= (layer2_outputs(10201)) and (layer2_outputs(4283));
    layer3_outputs(4528) <= not(layer2_outputs(8263));
    layer3_outputs(4529) <= (layer2_outputs(9294)) xor (layer2_outputs(4134));
    layer3_outputs(4530) <= layer2_outputs(7609);
    layer3_outputs(4531) <= layer2_outputs(3073);
    layer3_outputs(4532) <= not(layer2_outputs(7321));
    layer3_outputs(4533) <= (layer2_outputs(1175)) and (layer2_outputs(7442));
    layer3_outputs(4534) <= not(layer2_outputs(1611));
    layer3_outputs(4535) <= not(layer2_outputs(6227)) or (layer2_outputs(5770));
    layer3_outputs(4536) <= not(layer2_outputs(2467));
    layer3_outputs(4537) <= (layer2_outputs(5550)) and not (layer2_outputs(2514));
    layer3_outputs(4538) <= not(layer2_outputs(2989));
    layer3_outputs(4539) <= not(layer2_outputs(9709));
    layer3_outputs(4540) <= layer2_outputs(10131);
    layer3_outputs(4541) <= layer2_outputs(9218);
    layer3_outputs(4542) <= not(layer2_outputs(7238));
    layer3_outputs(4543) <= not(layer2_outputs(3065));
    layer3_outputs(4544) <= layer2_outputs(323);
    layer3_outputs(4545) <= not(layer2_outputs(3350));
    layer3_outputs(4546) <= not(layer2_outputs(2069)) or (layer2_outputs(4966));
    layer3_outputs(4547) <= layer2_outputs(2204);
    layer3_outputs(4548) <= not(layer2_outputs(2529));
    layer3_outputs(4549) <= (layer2_outputs(8070)) and not (layer2_outputs(1218));
    layer3_outputs(4550) <= layer2_outputs(4241);
    layer3_outputs(4551) <= layer2_outputs(7085);
    layer3_outputs(4552) <= not(layer2_outputs(3378));
    layer3_outputs(4553) <= (layer2_outputs(9181)) and not (layer2_outputs(3139));
    layer3_outputs(4554) <= layer2_outputs(1316);
    layer3_outputs(4555) <= layer2_outputs(9082);
    layer3_outputs(4556) <= (layer2_outputs(5470)) or (layer2_outputs(5988));
    layer3_outputs(4557) <= not(layer2_outputs(1493));
    layer3_outputs(4558) <= not((layer2_outputs(8358)) xor (layer2_outputs(1041)));
    layer3_outputs(4559) <= not(layer2_outputs(4728));
    layer3_outputs(4560) <= not(layer2_outputs(4542));
    layer3_outputs(4561) <= not(layer2_outputs(3712)) or (layer2_outputs(5382));
    layer3_outputs(4562) <= layer2_outputs(1647);
    layer3_outputs(4563) <= layer2_outputs(4723);
    layer3_outputs(4564) <= layer2_outputs(5605);
    layer3_outputs(4565) <= not(layer2_outputs(1247)) or (layer2_outputs(994));
    layer3_outputs(4566) <= not((layer2_outputs(3247)) and (layer2_outputs(7689)));
    layer3_outputs(4567) <= not(layer2_outputs(1246)) or (layer2_outputs(7820));
    layer3_outputs(4568) <= not(layer2_outputs(3794));
    layer3_outputs(4569) <= not(layer2_outputs(4708));
    layer3_outputs(4570) <= not(layer2_outputs(43));
    layer3_outputs(4571) <= (layer2_outputs(7012)) xor (layer2_outputs(5264));
    layer3_outputs(4572) <= not(layer2_outputs(2502));
    layer3_outputs(4573) <= (layer2_outputs(601)) and not (layer2_outputs(5827));
    layer3_outputs(4574) <= not((layer2_outputs(8791)) and (layer2_outputs(4266)));
    layer3_outputs(4575) <= not((layer2_outputs(7602)) or (layer2_outputs(1528)));
    layer3_outputs(4576) <= (layer2_outputs(9643)) and not (layer2_outputs(7958));
    layer3_outputs(4577) <= layer2_outputs(9157);
    layer3_outputs(4578) <= (layer2_outputs(8699)) and not (layer2_outputs(8487));
    layer3_outputs(4579) <= not(layer2_outputs(2276));
    layer3_outputs(4580) <= not(layer2_outputs(3539)) or (layer2_outputs(9521));
    layer3_outputs(4581) <= not(layer2_outputs(9876)) or (layer2_outputs(4075));
    layer3_outputs(4582) <= not(layer2_outputs(6973)) or (layer2_outputs(4391));
    layer3_outputs(4583) <= (layer2_outputs(8258)) xor (layer2_outputs(9104));
    layer3_outputs(4584) <= layer2_outputs(8936);
    layer3_outputs(4585) <= layer2_outputs(7375);
    layer3_outputs(4586) <= not(layer2_outputs(8079));
    layer3_outputs(4587) <= (layer2_outputs(607)) or (layer2_outputs(7575));
    layer3_outputs(4588) <= (layer2_outputs(6679)) and not (layer2_outputs(9416));
    layer3_outputs(4589) <= not((layer2_outputs(3796)) and (layer2_outputs(1430)));
    layer3_outputs(4590) <= layer2_outputs(5344);
    layer3_outputs(4591) <= layer2_outputs(2739);
    layer3_outputs(4592) <= not(layer2_outputs(4187));
    layer3_outputs(4593) <= (layer2_outputs(7775)) xor (layer2_outputs(9560));
    layer3_outputs(4594) <= not(layer2_outputs(372));
    layer3_outputs(4595) <= not((layer2_outputs(78)) xor (layer2_outputs(1601)));
    layer3_outputs(4596) <= layer2_outputs(7198);
    layer3_outputs(4597) <= (layer2_outputs(137)) or (layer2_outputs(5664));
    layer3_outputs(4598) <= not(layer2_outputs(5477));
    layer3_outputs(4599) <= not((layer2_outputs(1628)) xor (layer2_outputs(3749)));
    layer3_outputs(4600) <= not(layer2_outputs(1130)) or (layer2_outputs(1090));
    layer3_outputs(4601) <= (layer2_outputs(1890)) or (layer2_outputs(221));
    layer3_outputs(4602) <= not(layer2_outputs(6632));
    layer3_outputs(4603) <= (layer2_outputs(1927)) or (layer2_outputs(3302));
    layer3_outputs(4604) <= not(layer2_outputs(6038));
    layer3_outputs(4605) <= not(layer2_outputs(6199)) or (layer2_outputs(5566));
    layer3_outputs(4606) <= layer2_outputs(7038);
    layer3_outputs(4607) <= layer2_outputs(1954);
    layer3_outputs(4608) <= not(layer2_outputs(8747));
    layer3_outputs(4609) <= not(layer2_outputs(646));
    layer3_outputs(4610) <= (layer2_outputs(8052)) or (layer2_outputs(2043));
    layer3_outputs(4611) <= not((layer2_outputs(3868)) xor (layer2_outputs(2532)));
    layer3_outputs(4612) <= not(layer2_outputs(3415));
    layer3_outputs(4613) <= layer2_outputs(3342);
    layer3_outputs(4614) <= (layer2_outputs(9311)) xor (layer2_outputs(72));
    layer3_outputs(4615) <= layer2_outputs(6515);
    layer3_outputs(4616) <= not(layer2_outputs(8303));
    layer3_outputs(4617) <= not(layer2_outputs(3872));
    layer3_outputs(4618) <= (layer2_outputs(9755)) and (layer2_outputs(8364));
    layer3_outputs(4619) <= (layer2_outputs(5442)) xor (layer2_outputs(4533));
    layer3_outputs(4620) <= not(layer2_outputs(9035));
    layer3_outputs(4621) <= layer2_outputs(1213);
    layer3_outputs(4622) <= not(layer2_outputs(6042)) or (layer2_outputs(1792));
    layer3_outputs(4623) <= not((layer2_outputs(5678)) xor (layer2_outputs(8671)));
    layer3_outputs(4624) <= (layer2_outputs(8296)) xor (layer2_outputs(406));
    layer3_outputs(4625) <= not(layer2_outputs(5827));
    layer3_outputs(4626) <= layer2_outputs(2004);
    layer3_outputs(4627) <= not((layer2_outputs(8142)) and (layer2_outputs(123)));
    layer3_outputs(4628) <= layer2_outputs(165);
    layer3_outputs(4629) <= not((layer2_outputs(7232)) and (layer2_outputs(8204)));
    layer3_outputs(4630) <= not(layer2_outputs(7193));
    layer3_outputs(4631) <= '0';
    layer3_outputs(4632) <= '0';
    layer3_outputs(4633) <= layer2_outputs(7520);
    layer3_outputs(4634) <= layer2_outputs(8277);
    layer3_outputs(4635) <= not((layer2_outputs(430)) xor (layer2_outputs(8663)));
    layer3_outputs(4636) <= layer2_outputs(4943);
    layer3_outputs(4637) <= not((layer2_outputs(168)) and (layer2_outputs(1186)));
    layer3_outputs(4638) <= (layer2_outputs(7283)) and (layer2_outputs(1816));
    layer3_outputs(4639) <= (layer2_outputs(401)) and not (layer2_outputs(2260));
    layer3_outputs(4640) <= (layer2_outputs(7773)) or (layer2_outputs(8579));
    layer3_outputs(4641) <= layer2_outputs(4240);
    layer3_outputs(4642) <= '1';
    layer3_outputs(4643) <= not(layer2_outputs(4975)) or (layer2_outputs(9971));
    layer3_outputs(4644) <= not(layer2_outputs(7888));
    layer3_outputs(4645) <= not(layer2_outputs(6231));
    layer3_outputs(4646) <= not(layer2_outputs(1714)) or (layer2_outputs(4061));
    layer3_outputs(4647) <= not(layer2_outputs(8185));
    layer3_outputs(4648) <= not(layer2_outputs(8359));
    layer3_outputs(4649) <= (layer2_outputs(5685)) and (layer2_outputs(8553));
    layer3_outputs(4650) <= not(layer2_outputs(4782));
    layer3_outputs(4651) <= (layer2_outputs(8025)) and (layer2_outputs(1492));
    layer3_outputs(4652) <= layer2_outputs(8424);
    layer3_outputs(4653) <= not(layer2_outputs(2419)) or (layer2_outputs(3936));
    layer3_outputs(4654) <= not((layer2_outputs(2398)) or (layer2_outputs(1880)));
    layer3_outputs(4655) <= (layer2_outputs(1212)) and (layer2_outputs(8922));
    layer3_outputs(4656) <= not(layer2_outputs(6955));
    layer3_outputs(4657) <= not(layer2_outputs(10136));
    layer3_outputs(4658) <= not((layer2_outputs(1802)) xor (layer2_outputs(3152)));
    layer3_outputs(4659) <= (layer2_outputs(3938)) and not (layer2_outputs(125));
    layer3_outputs(4660) <= layer2_outputs(8726);
    layer3_outputs(4661) <= (layer2_outputs(273)) and not (layer2_outputs(6444));
    layer3_outputs(4662) <= layer2_outputs(5665);
    layer3_outputs(4663) <= not(layer2_outputs(5051));
    layer3_outputs(4664) <= layer2_outputs(7531);
    layer3_outputs(4665) <= (layer2_outputs(3057)) and (layer2_outputs(2569));
    layer3_outputs(4666) <= (layer2_outputs(7915)) or (layer2_outputs(133));
    layer3_outputs(4667) <= not(layer2_outputs(5679));
    layer3_outputs(4668) <= not(layer2_outputs(8333)) or (layer2_outputs(4219));
    layer3_outputs(4669) <= (layer2_outputs(8218)) and not (layer2_outputs(2261));
    layer3_outputs(4670) <= layer2_outputs(8967);
    layer3_outputs(4671) <= not(layer2_outputs(9056));
    layer3_outputs(4672) <= not(layer2_outputs(4768));
    layer3_outputs(4673) <= not(layer2_outputs(2925));
    layer3_outputs(4674) <= not(layer2_outputs(5631));
    layer3_outputs(4675) <= not(layer2_outputs(7158));
    layer3_outputs(4676) <= not(layer2_outputs(487)) or (layer2_outputs(9978));
    layer3_outputs(4677) <= '1';
    layer3_outputs(4678) <= not(layer2_outputs(4029));
    layer3_outputs(4679) <= layer2_outputs(8388);
    layer3_outputs(4680) <= (layer2_outputs(3437)) and not (layer2_outputs(1252));
    layer3_outputs(4681) <= not(layer2_outputs(538));
    layer3_outputs(4682) <= layer2_outputs(6974);
    layer3_outputs(4683) <= layer2_outputs(4380);
    layer3_outputs(4684) <= not(layer2_outputs(9679));
    layer3_outputs(4685) <= (layer2_outputs(9479)) and not (layer2_outputs(6220));
    layer3_outputs(4686) <= not(layer2_outputs(9081));
    layer3_outputs(4687) <= layer2_outputs(4501);
    layer3_outputs(4688) <= (layer2_outputs(7706)) and (layer2_outputs(4583));
    layer3_outputs(4689) <= not(layer2_outputs(702));
    layer3_outputs(4690) <= layer2_outputs(4270);
    layer3_outputs(4691) <= not((layer2_outputs(7374)) or (layer2_outputs(7982)));
    layer3_outputs(4692) <= layer2_outputs(5295);
    layer3_outputs(4693) <= not((layer2_outputs(4691)) or (layer2_outputs(4039)));
    layer3_outputs(4694) <= layer2_outputs(9078);
    layer3_outputs(4695) <= layer2_outputs(8357);
    layer3_outputs(4696) <= '0';
    layer3_outputs(4697) <= (layer2_outputs(3910)) xor (layer2_outputs(4920));
    layer3_outputs(4698) <= not(layer2_outputs(10159));
    layer3_outputs(4699) <= (layer2_outputs(2060)) and not (layer2_outputs(8544));
    layer3_outputs(4700) <= not((layer2_outputs(9993)) xor (layer2_outputs(6982)));
    layer3_outputs(4701) <= not(layer2_outputs(5699)) or (layer2_outputs(1733));
    layer3_outputs(4702) <= not((layer2_outputs(6808)) xor (layer2_outputs(2708)));
    layer3_outputs(4703) <= (layer2_outputs(7488)) and (layer2_outputs(7927));
    layer3_outputs(4704) <= layer2_outputs(5611);
    layer3_outputs(4705) <= layer2_outputs(4727);
    layer3_outputs(4706) <= (layer2_outputs(624)) and not (layer2_outputs(8879));
    layer3_outputs(4707) <= not(layer2_outputs(2827));
    layer3_outputs(4708) <= not((layer2_outputs(1839)) and (layer2_outputs(1683)));
    layer3_outputs(4709) <= not(layer2_outputs(5043));
    layer3_outputs(4710) <= (layer2_outputs(9533)) or (layer2_outputs(2465));
    layer3_outputs(4711) <= not(layer2_outputs(7471));
    layer3_outputs(4712) <= not(layer2_outputs(4245));
    layer3_outputs(4713) <= (layer2_outputs(3009)) and not (layer2_outputs(4168));
    layer3_outputs(4714) <= not(layer2_outputs(475)) or (layer2_outputs(8074));
    layer3_outputs(4715) <= layer2_outputs(2330);
    layer3_outputs(4716) <= not(layer2_outputs(6011));
    layer3_outputs(4717) <= layer2_outputs(9516);
    layer3_outputs(4718) <= '0';
    layer3_outputs(4719) <= layer2_outputs(6291);
    layer3_outputs(4720) <= (layer2_outputs(9997)) xor (layer2_outputs(6990));
    layer3_outputs(4721) <= layer2_outputs(3695);
    layer3_outputs(4722) <= not(layer2_outputs(5021));
    layer3_outputs(4723) <= not((layer2_outputs(2433)) and (layer2_outputs(1955)));
    layer3_outputs(4724) <= not((layer2_outputs(4483)) or (layer2_outputs(3257)));
    layer3_outputs(4725) <= not(layer2_outputs(3634));
    layer3_outputs(4726) <= not((layer2_outputs(214)) and (layer2_outputs(6362)));
    layer3_outputs(4727) <= not(layer2_outputs(9417)) or (layer2_outputs(9170));
    layer3_outputs(4728) <= not((layer2_outputs(7127)) or (layer2_outputs(2551)));
    layer3_outputs(4729) <= layer2_outputs(1253);
    layer3_outputs(4730) <= not(layer2_outputs(2522));
    layer3_outputs(4731) <= layer2_outputs(2090);
    layer3_outputs(4732) <= not((layer2_outputs(6529)) and (layer2_outputs(7191)));
    layer3_outputs(4733) <= not((layer2_outputs(7851)) or (layer2_outputs(1025)));
    layer3_outputs(4734) <= not(layer2_outputs(5378));
    layer3_outputs(4735) <= layer2_outputs(882);
    layer3_outputs(4736) <= not((layer2_outputs(2904)) xor (layer2_outputs(2389)));
    layer3_outputs(4737) <= (layer2_outputs(8176)) xor (layer2_outputs(108));
    layer3_outputs(4738) <= not((layer2_outputs(1261)) and (layer2_outputs(4447)));
    layer3_outputs(4739) <= (layer2_outputs(779)) and not (layer2_outputs(5425));
    layer3_outputs(4740) <= not(layer2_outputs(6059));
    layer3_outputs(4741) <= layer2_outputs(102);
    layer3_outputs(4742) <= not(layer2_outputs(6472)) or (layer2_outputs(4319));
    layer3_outputs(4743) <= not((layer2_outputs(7470)) and (layer2_outputs(609)));
    layer3_outputs(4744) <= not((layer2_outputs(5140)) xor (layer2_outputs(3419)));
    layer3_outputs(4745) <= (layer2_outputs(1561)) or (layer2_outputs(5334));
    layer3_outputs(4746) <= (layer2_outputs(2662)) xor (layer2_outputs(541));
    layer3_outputs(4747) <= (layer2_outputs(2249)) and not (layer2_outputs(1120));
    layer3_outputs(4748) <= not(layer2_outputs(1896)) or (layer2_outputs(4051));
    layer3_outputs(4749) <= layer2_outputs(3929);
    layer3_outputs(4750) <= not(layer2_outputs(1238));
    layer3_outputs(4751) <= '0';
    layer3_outputs(4752) <= layer2_outputs(4535);
    layer3_outputs(4753) <= (layer2_outputs(5255)) xor (layer2_outputs(5963));
    layer3_outputs(4754) <= not(layer2_outputs(2269)) or (layer2_outputs(7350));
    layer3_outputs(4755) <= '1';
    layer3_outputs(4756) <= layer2_outputs(3266);
    layer3_outputs(4757) <= not(layer2_outputs(7056));
    layer3_outputs(4758) <= (layer2_outputs(6544)) and not (layer2_outputs(6028));
    layer3_outputs(4759) <= (layer2_outputs(8959)) and not (layer2_outputs(8192));
    layer3_outputs(4760) <= (layer2_outputs(4087)) and not (layer2_outputs(7571));
    layer3_outputs(4761) <= layer2_outputs(6223);
    layer3_outputs(4762) <= (layer2_outputs(5794)) or (layer2_outputs(7961));
    layer3_outputs(4763) <= layer2_outputs(7047);
    layer3_outputs(4764) <= (layer2_outputs(1850)) and (layer2_outputs(1690));
    layer3_outputs(4765) <= not(layer2_outputs(8700));
    layer3_outputs(4766) <= not(layer2_outputs(128)) or (layer2_outputs(6758));
    layer3_outputs(4767) <= not((layer2_outputs(9224)) and (layer2_outputs(4736)));
    layer3_outputs(4768) <= not(layer2_outputs(890));
    layer3_outputs(4769) <= not(layer2_outputs(304));
    layer3_outputs(4770) <= not(layer2_outputs(10218));
    layer3_outputs(4771) <= layer2_outputs(7690);
    layer3_outputs(4772) <= not(layer2_outputs(7092));
    layer3_outputs(4773) <= layer2_outputs(6226);
    layer3_outputs(4774) <= (layer2_outputs(9383)) xor (layer2_outputs(9132));
    layer3_outputs(4775) <= not(layer2_outputs(8570)) or (layer2_outputs(5408));
    layer3_outputs(4776) <= layer2_outputs(5737);
    layer3_outputs(4777) <= not((layer2_outputs(9073)) and (layer2_outputs(4788)));
    layer3_outputs(4778) <= not(layer2_outputs(1125));
    layer3_outputs(4779) <= layer2_outputs(7502);
    layer3_outputs(4780) <= (layer2_outputs(6873)) xor (layer2_outputs(8923));
    layer3_outputs(4781) <= (layer2_outputs(6314)) and (layer2_outputs(6690));
    layer3_outputs(4782) <= layer2_outputs(8295);
    layer3_outputs(4783) <= not(layer2_outputs(7697));
    layer3_outputs(4784) <= not(layer2_outputs(6968));
    layer3_outputs(4785) <= layer2_outputs(3755);
    layer3_outputs(4786) <= not((layer2_outputs(9331)) xor (layer2_outputs(9652)));
    layer3_outputs(4787) <= not(layer2_outputs(7444)) or (layer2_outputs(6474));
    layer3_outputs(4788) <= (layer2_outputs(3102)) and not (layer2_outputs(876));
    layer3_outputs(4789) <= layer2_outputs(5674);
    layer3_outputs(4790) <= not(layer2_outputs(2098));
    layer3_outputs(4791) <= not(layer2_outputs(7173)) or (layer2_outputs(513));
    layer3_outputs(4792) <= layer2_outputs(4934);
    layer3_outputs(4793) <= layer2_outputs(1489);
    layer3_outputs(4794) <= not((layer2_outputs(1970)) xor (layer2_outputs(8549)));
    layer3_outputs(4795) <= (layer2_outputs(3508)) and not (layer2_outputs(1843));
    layer3_outputs(4796) <= not(layer2_outputs(8588)) or (layer2_outputs(3826));
    layer3_outputs(4797) <= (layer2_outputs(4100)) and not (layer2_outputs(6968));
    layer3_outputs(4798) <= not((layer2_outputs(6219)) xor (layer2_outputs(9049)));
    layer3_outputs(4799) <= (layer2_outputs(10147)) and (layer2_outputs(6450));
    layer3_outputs(4800) <= not(layer2_outputs(3823));
    layer3_outputs(4801) <= (layer2_outputs(4436)) and not (layer2_outputs(6634));
    layer3_outputs(4802) <= not((layer2_outputs(5497)) or (layer2_outputs(9339)));
    layer3_outputs(4803) <= not(layer2_outputs(10180));
    layer3_outputs(4804) <= (layer2_outputs(278)) and (layer2_outputs(437));
    layer3_outputs(4805) <= (layer2_outputs(10057)) xor (layer2_outputs(2392));
    layer3_outputs(4806) <= layer2_outputs(455);
    layer3_outputs(4807) <= layer2_outputs(8363);
    layer3_outputs(4808) <= not(layer2_outputs(1804));
    layer3_outputs(4809) <= layer2_outputs(799);
    layer3_outputs(4810) <= (layer2_outputs(5512)) and (layer2_outputs(6271));
    layer3_outputs(4811) <= not((layer2_outputs(8306)) and (layer2_outputs(9931)));
    layer3_outputs(4812) <= layer2_outputs(9249);
    layer3_outputs(4813) <= layer2_outputs(4443);
    layer3_outputs(4814) <= not((layer2_outputs(6341)) or (layer2_outputs(5514)));
    layer3_outputs(4815) <= not(layer2_outputs(563));
    layer3_outputs(4816) <= not(layer2_outputs(9471));
    layer3_outputs(4817) <= (layer2_outputs(4735)) and not (layer2_outputs(6071));
    layer3_outputs(4818) <= not(layer2_outputs(7019)) or (layer2_outputs(4933));
    layer3_outputs(4819) <= not((layer2_outputs(338)) xor (layer2_outputs(8591)));
    layer3_outputs(4820) <= layer2_outputs(5478);
    layer3_outputs(4821) <= layer2_outputs(7981);
    layer3_outputs(4822) <= not((layer2_outputs(6183)) xor (layer2_outputs(4221)));
    layer3_outputs(4823) <= '1';
    layer3_outputs(4824) <= not((layer2_outputs(4640)) xor (layer2_outputs(6490)));
    layer3_outputs(4825) <= layer2_outputs(9512);
    layer3_outputs(4826) <= not(layer2_outputs(2772)) or (layer2_outputs(5946));
    layer3_outputs(4827) <= (layer2_outputs(3509)) xor (layer2_outputs(9529));
    layer3_outputs(4828) <= (layer2_outputs(3242)) and (layer2_outputs(7278));
    layer3_outputs(4829) <= layer2_outputs(4202);
    layer3_outputs(4830) <= (layer2_outputs(5648)) and not (layer2_outputs(598));
    layer3_outputs(4831) <= (layer2_outputs(5338)) xor (layer2_outputs(5524));
    layer3_outputs(4832) <= not(layer2_outputs(4227));
    layer3_outputs(4833) <= layer2_outputs(9086);
    layer3_outputs(4834) <= (layer2_outputs(6560)) and not (layer2_outputs(7394));
    layer3_outputs(4835) <= not(layer2_outputs(3500));
    layer3_outputs(4836) <= (layer2_outputs(9879)) and not (layer2_outputs(4968));
    layer3_outputs(4837) <= layer2_outputs(2898);
    layer3_outputs(4838) <= not(layer2_outputs(989));
    layer3_outputs(4839) <= (layer2_outputs(840)) and not (layer2_outputs(5206));
    layer3_outputs(4840) <= not(layer2_outputs(3944));
    layer3_outputs(4841) <= layer2_outputs(2948);
    layer3_outputs(4842) <= (layer2_outputs(5346)) and not (layer2_outputs(4414));
    layer3_outputs(4843) <= (layer2_outputs(6428)) or (layer2_outputs(1836));
    layer3_outputs(4844) <= not(layer2_outputs(2194));
    layer3_outputs(4845) <= not((layer2_outputs(4203)) or (layer2_outputs(1108)));
    layer3_outputs(4846) <= layer2_outputs(7527);
    layer3_outputs(4847) <= not((layer2_outputs(902)) and (layer2_outputs(6585)));
    layer3_outputs(4848) <= layer2_outputs(9279);
    layer3_outputs(4849) <= layer2_outputs(5865);
    layer3_outputs(4850) <= (layer2_outputs(4984)) or (layer2_outputs(8081));
    layer3_outputs(4851) <= (layer2_outputs(9365)) xor (layer2_outputs(9130));
    layer3_outputs(4852) <= not(layer2_outputs(3193)) or (layer2_outputs(3876));
    layer3_outputs(4853) <= (layer2_outputs(7100)) xor (layer2_outputs(9649));
    layer3_outputs(4854) <= not(layer2_outputs(8156));
    layer3_outputs(4855) <= not(layer2_outputs(1333));
    layer3_outputs(4856) <= not((layer2_outputs(5951)) and (layer2_outputs(7146)));
    layer3_outputs(4857) <= layer2_outputs(581);
    layer3_outputs(4858) <= layer2_outputs(5672);
    layer3_outputs(4859) <= '1';
    layer3_outputs(4860) <= layer2_outputs(7599);
    layer3_outputs(4861) <= (layer2_outputs(8497)) or (layer2_outputs(7683));
    layer3_outputs(4862) <= not(layer2_outputs(6533));
    layer3_outputs(4863) <= not(layer2_outputs(7986)) or (layer2_outputs(1466));
    layer3_outputs(4864) <= not(layer2_outputs(6389)) or (layer2_outputs(5591));
    layer3_outputs(4865) <= not(layer2_outputs(4597));
    layer3_outputs(4866) <= (layer2_outputs(5986)) and (layer2_outputs(3575));
    layer3_outputs(4867) <= layer2_outputs(507);
    layer3_outputs(4868) <= layer2_outputs(9589);
    layer3_outputs(4869) <= (layer2_outputs(8323)) and not (layer2_outputs(2064));
    layer3_outputs(4870) <= not(layer2_outputs(2922));
    layer3_outputs(4871) <= (layer2_outputs(2430)) or (layer2_outputs(8716));
    layer3_outputs(4872) <= (layer2_outputs(4807)) or (layer2_outputs(8741));
    layer3_outputs(4873) <= '0';
    layer3_outputs(4874) <= not(layer2_outputs(1447));
    layer3_outputs(4875) <= (layer2_outputs(1882)) xor (layer2_outputs(5700));
    layer3_outputs(4876) <= not((layer2_outputs(6910)) xor (layer2_outputs(7128)));
    layer3_outputs(4877) <= not(layer2_outputs(1594));
    layer3_outputs(4878) <= not(layer2_outputs(7214));
    layer3_outputs(4879) <= not(layer2_outputs(7653)) or (layer2_outputs(2474));
    layer3_outputs(4880) <= layer2_outputs(6482);
    layer3_outputs(4881) <= not(layer2_outputs(8520)) or (layer2_outputs(4252));
    layer3_outputs(4882) <= layer2_outputs(9935);
    layer3_outputs(4883) <= not((layer2_outputs(9333)) or (layer2_outputs(4396)));
    layer3_outputs(4884) <= not(layer2_outputs(7836));
    layer3_outputs(4885) <= (layer2_outputs(4842)) xor (layer2_outputs(4001));
    layer3_outputs(4886) <= layer2_outputs(3484);
    layer3_outputs(4887) <= layer2_outputs(3178);
    layer3_outputs(4888) <= not(layer2_outputs(2513));
    layer3_outputs(4889) <= not(layer2_outputs(9533)) or (layer2_outputs(1860));
    layer3_outputs(4890) <= layer2_outputs(1810);
    layer3_outputs(4891) <= not((layer2_outputs(4634)) xor (layer2_outputs(2124)));
    layer3_outputs(4892) <= not(layer2_outputs(5608));
    layer3_outputs(4893) <= (layer2_outputs(2687)) and not (layer2_outputs(4958));
    layer3_outputs(4894) <= not(layer2_outputs(5084)) or (layer2_outputs(4743));
    layer3_outputs(4895) <= not(layer2_outputs(8866));
    layer3_outputs(4896) <= layer2_outputs(6322);
    layer3_outputs(4897) <= not(layer2_outputs(2426));
    layer3_outputs(4898) <= not((layer2_outputs(3775)) xor (layer2_outputs(7645)));
    layer3_outputs(4899) <= not(layer2_outputs(2437));
    layer3_outputs(4900) <= not(layer2_outputs(3647)) or (layer2_outputs(4105));
    layer3_outputs(4901) <= not((layer2_outputs(2921)) or (layer2_outputs(6739)));
    layer3_outputs(4902) <= layer2_outputs(10177);
    layer3_outputs(4903) <= (layer2_outputs(9462)) and not (layer2_outputs(4408));
    layer3_outputs(4904) <= not((layer2_outputs(1011)) xor (layer2_outputs(391)));
    layer3_outputs(4905) <= not(layer2_outputs(8328)) or (layer2_outputs(2764));
    layer3_outputs(4906) <= (layer2_outputs(473)) and (layer2_outputs(6505));
    layer3_outputs(4907) <= not((layer2_outputs(7781)) or (layer2_outputs(1838)));
    layer3_outputs(4908) <= (layer2_outputs(1864)) xor (layer2_outputs(4385));
    layer3_outputs(4909) <= not(layer2_outputs(1250)) or (layer2_outputs(9105));
    layer3_outputs(4910) <= layer2_outputs(7085);
    layer3_outputs(4911) <= (layer2_outputs(3676)) and not (layer2_outputs(7132));
    layer3_outputs(4912) <= layer2_outputs(9413);
    layer3_outputs(4913) <= not(layer2_outputs(7846)) or (layer2_outputs(9464));
    layer3_outputs(4914) <= not((layer2_outputs(3706)) and (layer2_outputs(7576)));
    layer3_outputs(4915) <= not(layer2_outputs(421));
    layer3_outputs(4916) <= layer2_outputs(1423);
    layer3_outputs(4917) <= layer2_outputs(5372);
    layer3_outputs(4918) <= (layer2_outputs(4780)) and not (layer2_outputs(9283));
    layer3_outputs(4919) <= (layer2_outputs(667)) and not (layer2_outputs(2875));
    layer3_outputs(4920) <= (layer2_outputs(2716)) xor (layer2_outputs(6886));
    layer3_outputs(4921) <= not((layer2_outputs(8504)) xor (layer2_outputs(1427)));
    layer3_outputs(4922) <= layer2_outputs(3919);
    layer3_outputs(4923) <= not((layer2_outputs(6232)) and (layer2_outputs(6486)));
    layer3_outputs(4924) <= not(layer2_outputs(7248));
    layer3_outputs(4925) <= (layer2_outputs(4480)) and not (layer2_outputs(8438));
    layer3_outputs(4926) <= not(layer2_outputs(546)) or (layer2_outputs(8903));
    layer3_outputs(4927) <= (layer2_outputs(3871)) or (layer2_outputs(3644));
    layer3_outputs(4928) <= not(layer2_outputs(10047));
    layer3_outputs(4929) <= not((layer2_outputs(7432)) or (layer2_outputs(1526)));
    layer3_outputs(4930) <= layer2_outputs(203);
    layer3_outputs(4931) <= not(layer2_outputs(1884)) or (layer2_outputs(10007));
    layer3_outputs(4932) <= '1';
    layer3_outputs(4933) <= not((layer2_outputs(3142)) and (layer2_outputs(5926)));
    layer3_outputs(4934) <= not(layer2_outputs(9085));
    layer3_outputs(4935) <= not((layer2_outputs(5615)) or (layer2_outputs(1603)));
    layer3_outputs(4936) <= not(layer2_outputs(2511));
    layer3_outputs(4937) <= layer2_outputs(4815);
    layer3_outputs(4938) <= layer2_outputs(7158);
    layer3_outputs(4939) <= (layer2_outputs(8476)) or (layer2_outputs(9563));
    layer3_outputs(4940) <= (layer2_outputs(8928)) or (layer2_outputs(5066));
    layer3_outputs(4941) <= '0';
    layer3_outputs(4942) <= (layer2_outputs(51)) xor (layer2_outputs(2242));
    layer3_outputs(4943) <= layer2_outputs(7467);
    layer3_outputs(4944) <= not(layer2_outputs(2100));
    layer3_outputs(4945) <= layer2_outputs(4814);
    layer3_outputs(4946) <= (layer2_outputs(4508)) and (layer2_outputs(8294));
    layer3_outputs(4947) <= not(layer2_outputs(7008));
    layer3_outputs(4948) <= not(layer2_outputs(3588));
    layer3_outputs(4949) <= not(layer2_outputs(514)) or (layer2_outputs(9939));
    layer3_outputs(4950) <= not((layer2_outputs(6905)) and (layer2_outputs(3959)));
    layer3_outputs(4951) <= (layer2_outputs(6077)) and (layer2_outputs(9605));
    layer3_outputs(4952) <= not(layer2_outputs(3762));
    layer3_outputs(4953) <= (layer2_outputs(1709)) and not (layer2_outputs(7149));
    layer3_outputs(4954) <= not((layer2_outputs(1111)) and (layer2_outputs(1693)));
    layer3_outputs(4955) <= layer2_outputs(2735);
    layer3_outputs(4956) <= (layer2_outputs(8615)) and not (layer2_outputs(9120));
    layer3_outputs(4957) <= not((layer2_outputs(1346)) xor (layer2_outputs(5202)));
    layer3_outputs(4958) <= not((layer2_outputs(8474)) or (layer2_outputs(3792)));
    layer3_outputs(4959) <= layer2_outputs(700);
    layer3_outputs(4960) <= not(layer2_outputs(6338)) or (layer2_outputs(7883));
    layer3_outputs(4961) <= not((layer2_outputs(7357)) and (layer2_outputs(9785)));
    layer3_outputs(4962) <= layer2_outputs(774);
    layer3_outputs(4963) <= not(layer2_outputs(1464));
    layer3_outputs(4964) <= not(layer2_outputs(9668)) or (layer2_outputs(1370));
    layer3_outputs(4965) <= not((layer2_outputs(5811)) or (layer2_outputs(9506)));
    layer3_outputs(4966) <= not((layer2_outputs(4523)) xor (layer2_outputs(4084)));
    layer3_outputs(4967) <= (layer2_outputs(10011)) or (layer2_outputs(8665));
    layer3_outputs(4968) <= not((layer2_outputs(8617)) xor (layer2_outputs(9747)));
    layer3_outputs(4969) <= (layer2_outputs(6816)) or (layer2_outputs(9226));
    layer3_outputs(4970) <= not((layer2_outputs(457)) or (layer2_outputs(760)));
    layer3_outputs(4971) <= (layer2_outputs(768)) xor (layer2_outputs(1507));
    layer3_outputs(4972) <= not((layer2_outputs(3574)) xor (layer2_outputs(7474)));
    layer3_outputs(4973) <= not(layer2_outputs(1340));
    layer3_outputs(4974) <= not(layer2_outputs(7971));
    layer3_outputs(4975) <= (layer2_outputs(952)) xor (layer2_outputs(6151));
    layer3_outputs(4976) <= (layer2_outputs(4914)) and not (layer2_outputs(3991));
    layer3_outputs(4977) <= (layer2_outputs(1135)) and (layer2_outputs(1162));
    layer3_outputs(4978) <= not((layer2_outputs(3065)) and (layer2_outputs(6038)));
    layer3_outputs(4979) <= not(layer2_outputs(7787));
    layer3_outputs(4980) <= (layer2_outputs(7568)) xor (layer2_outputs(6622));
    layer3_outputs(4981) <= layer2_outputs(4826);
    layer3_outputs(4982) <= not(layer2_outputs(5002));
    layer3_outputs(4983) <= not(layer2_outputs(904)) or (layer2_outputs(8750));
    layer3_outputs(4984) <= layer2_outputs(1980);
    layer3_outputs(4985) <= not(layer2_outputs(2519));
    layer3_outputs(4986) <= (layer2_outputs(8838)) and not (layer2_outputs(2024));
    layer3_outputs(4987) <= layer2_outputs(8799);
    layer3_outputs(4988) <= (layer2_outputs(6242)) or (layer2_outputs(1221));
    layer3_outputs(4989) <= not((layer2_outputs(10028)) xor (layer2_outputs(1797)));
    layer3_outputs(4990) <= layer2_outputs(9867);
    layer3_outputs(4991) <= (layer2_outputs(1480)) or (layer2_outputs(8678));
    layer3_outputs(4992) <= layer2_outputs(8173);
    layer3_outputs(4993) <= (layer2_outputs(89)) or (layer2_outputs(1064));
    layer3_outputs(4994) <= not((layer2_outputs(2850)) or (layer2_outputs(5332)));
    layer3_outputs(4995) <= (layer2_outputs(2709)) and (layer2_outputs(6716));
    layer3_outputs(4996) <= layer2_outputs(466);
    layer3_outputs(4997) <= layer2_outputs(983);
    layer3_outputs(4998) <= not(layer2_outputs(3502));
    layer3_outputs(4999) <= not(layer2_outputs(4326)) or (layer2_outputs(10008));
    layer3_outputs(5000) <= layer2_outputs(6489);
    layer3_outputs(5001) <= not(layer2_outputs(712));
    layer3_outputs(5002) <= not((layer2_outputs(5956)) and (layer2_outputs(8421)));
    layer3_outputs(5003) <= (layer2_outputs(1049)) or (layer2_outputs(808));
    layer3_outputs(5004) <= layer2_outputs(4883);
    layer3_outputs(5005) <= not((layer2_outputs(2280)) or (layer2_outputs(2297)));
    layer3_outputs(5006) <= not((layer2_outputs(7579)) or (layer2_outputs(8785)));
    layer3_outputs(5007) <= not(layer2_outputs(9427));
    layer3_outputs(5008) <= (layer2_outputs(4682)) and not (layer2_outputs(2984));
    layer3_outputs(5009) <= '0';
    layer3_outputs(5010) <= not(layer2_outputs(4317));
    layer3_outputs(5011) <= not(layer2_outputs(4409));
    layer3_outputs(5012) <= not(layer2_outputs(6519));
    layer3_outputs(5013) <= (layer2_outputs(7855)) and (layer2_outputs(83));
    layer3_outputs(5014) <= (layer2_outputs(4646)) or (layer2_outputs(3975));
    layer3_outputs(5015) <= layer2_outputs(1694);
    layer3_outputs(5016) <= not(layer2_outputs(1021));
    layer3_outputs(5017) <= not((layer2_outputs(193)) or (layer2_outputs(8699)));
    layer3_outputs(5018) <= not((layer2_outputs(352)) and (layer2_outputs(9487)));
    layer3_outputs(5019) <= (layer2_outputs(2504)) and not (layer2_outputs(2974));
    layer3_outputs(5020) <= not(layer2_outputs(7227));
    layer3_outputs(5021) <= not(layer2_outputs(7746)) or (layer2_outputs(7931));
    layer3_outputs(5022) <= not(layer2_outputs(3915));
    layer3_outputs(5023) <= (layer2_outputs(4958)) xor (layer2_outputs(7092));
    layer3_outputs(5024) <= not(layer2_outputs(7797));
    layer3_outputs(5025) <= not(layer2_outputs(46));
    layer3_outputs(5026) <= (layer2_outputs(3849)) and (layer2_outputs(6536));
    layer3_outputs(5027) <= not(layer2_outputs(3111));
    layer3_outputs(5028) <= layer2_outputs(1322);
    layer3_outputs(5029) <= not(layer2_outputs(746));
    layer3_outputs(5030) <= layer2_outputs(8734);
    layer3_outputs(5031) <= not(layer2_outputs(8995));
    layer3_outputs(5032) <= not(layer2_outputs(5417));
    layer3_outputs(5033) <= not(layer2_outputs(9651));
    layer3_outputs(5034) <= not(layer2_outputs(7111));
    layer3_outputs(5035) <= not((layer2_outputs(8354)) xor (layer2_outputs(5997)));
    layer3_outputs(5036) <= not(layer2_outputs(1337));
    layer3_outputs(5037) <= not(layer2_outputs(4634));
    layer3_outputs(5038) <= (layer2_outputs(8495)) xor (layer2_outputs(5143));
    layer3_outputs(5039) <= layer2_outputs(8558);
    layer3_outputs(5040) <= layer2_outputs(3201);
    layer3_outputs(5041) <= (layer2_outputs(3842)) and not (layer2_outputs(2999));
    layer3_outputs(5042) <= layer2_outputs(695);
    layer3_outputs(5043) <= not(layer2_outputs(3856));
    layer3_outputs(5044) <= '1';
    layer3_outputs(5045) <= not(layer2_outputs(37)) or (layer2_outputs(2633));
    layer3_outputs(5046) <= not(layer2_outputs(3385));
    layer3_outputs(5047) <= not(layer2_outputs(3704));
    layer3_outputs(5048) <= layer2_outputs(3335);
    layer3_outputs(5049) <= (layer2_outputs(10077)) and not (layer2_outputs(6614));
    layer3_outputs(5050) <= not(layer2_outputs(4043));
    layer3_outputs(5051) <= (layer2_outputs(9350)) and (layer2_outputs(4616));
    layer3_outputs(5052) <= '1';
    layer3_outputs(5053) <= layer2_outputs(3765);
    layer3_outputs(5054) <= not(layer2_outputs(6866));
    layer3_outputs(5055) <= layer2_outputs(1339);
    layer3_outputs(5056) <= layer2_outputs(718);
    layer3_outputs(5057) <= (layer2_outputs(6595)) and (layer2_outputs(1458));
    layer3_outputs(5058) <= not(layer2_outputs(9245));
    layer3_outputs(5059) <= not((layer2_outputs(3041)) and (layer2_outputs(10207)));
    layer3_outputs(5060) <= not((layer2_outputs(7821)) or (layer2_outputs(6675)));
    layer3_outputs(5061) <= not(layer2_outputs(3531)) or (layer2_outputs(7662));
    layer3_outputs(5062) <= not((layer2_outputs(8810)) xor (layer2_outputs(1768)));
    layer3_outputs(5063) <= (layer2_outputs(6646)) or (layer2_outputs(5723));
    layer3_outputs(5064) <= layer2_outputs(5587);
    layer3_outputs(5065) <= not(layer2_outputs(9267));
    layer3_outputs(5066) <= (layer2_outputs(2707)) or (layer2_outputs(8488));
    layer3_outputs(5067) <= not((layer2_outputs(4739)) or (layer2_outputs(5156)));
    layer3_outputs(5068) <= layer2_outputs(2631);
    layer3_outputs(5069) <= (layer2_outputs(1432)) and not (layer2_outputs(5452));
    layer3_outputs(5070) <= (layer2_outputs(7025)) and not (layer2_outputs(2424));
    layer3_outputs(5071) <= not(layer2_outputs(3267));
    layer3_outputs(5072) <= layer2_outputs(6832);
    layer3_outputs(5073) <= (layer2_outputs(1059)) and not (layer2_outputs(9617));
    layer3_outputs(5074) <= not(layer2_outputs(1819));
    layer3_outputs(5075) <= not(layer2_outputs(7613));
    layer3_outputs(5076) <= not(layer2_outputs(6585));
    layer3_outputs(5077) <= not((layer2_outputs(3152)) and (layer2_outputs(2862)));
    layer3_outputs(5078) <= layer2_outputs(7076);
    layer3_outputs(5079) <= (layer2_outputs(2472)) or (layer2_outputs(4987));
    layer3_outputs(5080) <= layer2_outputs(9360);
    layer3_outputs(5081) <= not(layer2_outputs(6736)) or (layer2_outputs(9020));
    layer3_outputs(5082) <= (layer2_outputs(586)) xor (layer2_outputs(2931));
    layer3_outputs(5083) <= not(layer2_outputs(4459)) or (layer2_outputs(8513));
    layer3_outputs(5084) <= layer2_outputs(4191);
    layer3_outputs(5085) <= (layer2_outputs(7886)) xor (layer2_outputs(4893));
    layer3_outputs(5086) <= not(layer2_outputs(5076));
    layer3_outputs(5087) <= (layer2_outputs(2605)) and not (layer2_outputs(1986));
    layer3_outputs(5088) <= not(layer2_outputs(1910));
    layer3_outputs(5089) <= layer2_outputs(20);
    layer3_outputs(5090) <= not(layer2_outputs(3515)) or (layer2_outputs(7313));
    layer3_outputs(5091) <= layer2_outputs(9097);
    layer3_outputs(5092) <= layer2_outputs(1190);
    layer3_outputs(5093) <= not(layer2_outputs(651));
    layer3_outputs(5094) <= not(layer2_outputs(9875));
    layer3_outputs(5095) <= layer2_outputs(1164);
    layer3_outputs(5096) <= (layer2_outputs(5102)) and not (layer2_outputs(852));
    layer3_outputs(5097) <= not(layer2_outputs(2342));
    layer3_outputs(5098) <= not(layer2_outputs(6498)) or (layer2_outputs(6123));
    layer3_outputs(5099) <= not((layer2_outputs(6110)) and (layer2_outputs(7998)));
    layer3_outputs(5100) <= layer2_outputs(9678);
    layer3_outputs(5101) <= not((layer2_outputs(4831)) xor (layer2_outputs(5511)));
    layer3_outputs(5102) <= (layer2_outputs(10209)) or (layer2_outputs(7417));
    layer3_outputs(5103) <= (layer2_outputs(9092)) and (layer2_outputs(9185));
    layer3_outputs(5104) <= not(layer2_outputs(6641));
    layer3_outputs(5105) <= layer2_outputs(5331);
    layer3_outputs(5106) <= not(layer2_outputs(8239));
    layer3_outputs(5107) <= not(layer2_outputs(7991));
    layer3_outputs(5108) <= not(layer2_outputs(3714));
    layer3_outputs(5109) <= (layer2_outputs(8575)) xor (layer2_outputs(7065));
    layer3_outputs(5110) <= (layer2_outputs(5132)) and (layer2_outputs(4358));
    layer3_outputs(5111) <= not(layer2_outputs(5154)) or (layer2_outputs(2592));
    layer3_outputs(5112) <= not((layer2_outputs(2691)) or (layer2_outputs(7760)));
    layer3_outputs(5113) <= layer2_outputs(4692);
    layer3_outputs(5114) <= layer2_outputs(8535);
    layer3_outputs(5115) <= not(layer2_outputs(8210)) or (layer2_outputs(3520));
    layer3_outputs(5116) <= '0';
    layer3_outputs(5117) <= not(layer2_outputs(4400));
    layer3_outputs(5118) <= layer2_outputs(3858);
    layer3_outputs(5119) <= (layer2_outputs(6943)) and not (layer2_outputs(8896));
    layer3_outputs(5120) <= not((layer2_outputs(7161)) or (layer2_outputs(2642)));
    layer3_outputs(5121) <= layer2_outputs(2347);
    layer3_outputs(5122) <= not(layer2_outputs(8310)) or (layer2_outputs(4101));
    layer3_outputs(5123) <= not(layer2_outputs(9397));
    layer3_outputs(5124) <= not((layer2_outputs(736)) xor (layer2_outputs(2465)));
    layer3_outputs(5125) <= (layer2_outputs(9074)) and not (layer2_outputs(5216));
    layer3_outputs(5126) <= not(layer2_outputs(2382)) or (layer2_outputs(5637));
    layer3_outputs(5127) <= not(layer2_outputs(6260));
    layer3_outputs(5128) <= not((layer2_outputs(6885)) or (layer2_outputs(436)));
    layer3_outputs(5129) <= layer2_outputs(286);
    layer3_outputs(5130) <= not(layer2_outputs(893));
    layer3_outputs(5131) <= not((layer2_outputs(1811)) and (layer2_outputs(1985)));
    layer3_outputs(5132) <= not(layer2_outputs(7560)) or (layer2_outputs(8001));
    layer3_outputs(5133) <= layer2_outputs(2826);
    layer3_outputs(5134) <= layer2_outputs(8886);
    layer3_outputs(5135) <= not(layer2_outputs(4503)) or (layer2_outputs(5686));
    layer3_outputs(5136) <= not(layer2_outputs(825));
    layer3_outputs(5137) <= not((layer2_outputs(5495)) and (layer2_outputs(721)));
    layer3_outputs(5138) <= layer2_outputs(687);
    layer3_outputs(5139) <= layer2_outputs(4485);
    layer3_outputs(5140) <= not(layer2_outputs(3052));
    layer3_outputs(5141) <= (layer2_outputs(172)) or (layer2_outputs(182));
    layer3_outputs(5142) <= not(layer2_outputs(3799));
    layer3_outputs(5143) <= not((layer2_outputs(1658)) or (layer2_outputs(4687)));
    layer3_outputs(5144) <= not(layer2_outputs(2204));
    layer3_outputs(5145) <= not((layer2_outputs(8320)) or (layer2_outputs(707)));
    layer3_outputs(5146) <= not(layer2_outputs(6327));
    layer3_outputs(5147) <= (layer2_outputs(8065)) and not (layer2_outputs(1168));
    layer3_outputs(5148) <= not(layer2_outputs(6331)) or (layer2_outputs(7655));
    layer3_outputs(5149) <= layer2_outputs(4171);
    layer3_outputs(5150) <= not(layer2_outputs(2378));
    layer3_outputs(5151) <= not(layer2_outputs(4576));
    layer3_outputs(5152) <= not(layer2_outputs(2763));
    layer3_outputs(5153) <= (layer2_outputs(2087)) and (layer2_outputs(3827));
    layer3_outputs(5154) <= (layer2_outputs(2721)) xor (layer2_outputs(4628));
    layer3_outputs(5155) <= not((layer2_outputs(3166)) and (layer2_outputs(1235)));
    layer3_outputs(5156) <= not((layer2_outputs(2738)) and (layer2_outputs(5424)));
    layer3_outputs(5157) <= not((layer2_outputs(3221)) and (layer2_outputs(4656)));
    layer3_outputs(5158) <= not(layer2_outputs(3465)) or (layer2_outputs(1946));
    layer3_outputs(5159) <= layer2_outputs(3655);
    layer3_outputs(5160) <= layer2_outputs(3846);
    layer3_outputs(5161) <= layer2_outputs(4104);
    layer3_outputs(5162) <= layer2_outputs(1178);
    layer3_outputs(5163) <= layer2_outputs(5765);
    layer3_outputs(5164) <= layer2_outputs(7562);
    layer3_outputs(5165) <= not(layer2_outputs(8211)) or (layer2_outputs(3890));
    layer3_outputs(5166) <= not((layer2_outputs(9558)) and (layer2_outputs(3850)));
    layer3_outputs(5167) <= '0';
    layer3_outputs(5168) <= layer2_outputs(9252);
    layer3_outputs(5169) <= not(layer2_outputs(4828)) or (layer2_outputs(10186));
    layer3_outputs(5170) <= (layer2_outputs(1981)) xor (layer2_outputs(5937));
    layer3_outputs(5171) <= (layer2_outputs(209)) and not (layer2_outputs(1793));
    layer3_outputs(5172) <= not((layer2_outputs(3127)) and (layer2_outputs(9062)));
    layer3_outputs(5173) <= not(layer2_outputs(2375));
    layer3_outputs(5174) <= (layer2_outputs(609)) and not (layer2_outputs(7433));
    layer3_outputs(5175) <= '1';
    layer3_outputs(5176) <= not(layer2_outputs(9679));
    layer3_outputs(5177) <= not((layer2_outputs(8739)) or (layer2_outputs(7045)));
    layer3_outputs(5178) <= not(layer2_outputs(9448));
    layer3_outputs(5179) <= not(layer2_outputs(8710)) or (layer2_outputs(950));
    layer3_outputs(5180) <= layer2_outputs(796);
    layer3_outputs(5181) <= not(layer2_outputs(7901));
    layer3_outputs(5182) <= (layer2_outputs(3595)) and not (layer2_outputs(6189));
    layer3_outputs(5183) <= '0';
    layer3_outputs(5184) <= layer2_outputs(8268);
    layer3_outputs(5185) <= layer2_outputs(3308);
    layer3_outputs(5186) <= not(layer2_outputs(2915));
    layer3_outputs(5187) <= not((layer2_outputs(2008)) xor (layer2_outputs(1462)));
    layer3_outputs(5188) <= not((layer2_outputs(1742)) and (layer2_outputs(8821)));
    layer3_outputs(5189) <= not((layer2_outputs(6143)) and (layer2_outputs(9325)));
    layer3_outputs(5190) <= not(layer2_outputs(2766)) or (layer2_outputs(985));
    layer3_outputs(5191) <= not(layer2_outputs(9892)) or (layer2_outputs(2512));
    layer3_outputs(5192) <= '0';
    layer3_outputs(5193) <= not(layer2_outputs(3175));
    layer3_outputs(5194) <= not(layer2_outputs(9749)) or (layer2_outputs(549));
    layer3_outputs(5195) <= not(layer2_outputs(3444));
    layer3_outputs(5196) <= not(layer2_outputs(9412));
    layer3_outputs(5197) <= (layer2_outputs(5250)) and not (layer2_outputs(279));
    layer3_outputs(5198) <= layer2_outputs(1149);
    layer3_outputs(5199) <= (layer2_outputs(5180)) and not (layer2_outputs(7642));
    layer3_outputs(5200) <= (layer2_outputs(954)) and not (layer2_outputs(8770));
    layer3_outputs(5201) <= layer2_outputs(2630);
    layer3_outputs(5202) <= layer2_outputs(7053);
    layer3_outputs(5203) <= not((layer2_outputs(4586)) xor (layer2_outputs(10198)));
    layer3_outputs(5204) <= layer2_outputs(2610);
    layer3_outputs(5205) <= layer2_outputs(6844);
    layer3_outputs(5206) <= not(layer2_outputs(4512)) or (layer2_outputs(6644));
    layer3_outputs(5207) <= not(layer2_outputs(2654));
    layer3_outputs(5208) <= not((layer2_outputs(8038)) and (layer2_outputs(4091)));
    layer3_outputs(5209) <= (layer2_outputs(10052)) and not (layer2_outputs(5292));
    layer3_outputs(5210) <= layer2_outputs(6279);
    layer3_outputs(5211) <= not(layer2_outputs(9299)) or (layer2_outputs(3829));
    layer3_outputs(5212) <= layer2_outputs(1970);
    layer3_outputs(5213) <= not(layer2_outputs(8136));
    layer3_outputs(5214) <= not((layer2_outputs(2619)) or (layer2_outputs(7445)));
    layer3_outputs(5215) <= layer2_outputs(5620);
    layer3_outputs(5216) <= layer2_outputs(3743);
    layer3_outputs(5217) <= not(layer2_outputs(3396));
    layer3_outputs(5218) <= layer2_outputs(1842);
    layer3_outputs(5219) <= not(layer2_outputs(9300));
    layer3_outputs(5220) <= layer2_outputs(7034);
    layer3_outputs(5221) <= not(layer2_outputs(45));
    layer3_outputs(5222) <= (layer2_outputs(8008)) and not (layer2_outputs(1060));
    layer3_outputs(5223) <= not(layer2_outputs(5306)) or (layer2_outputs(5672));
    layer3_outputs(5224) <= not(layer2_outputs(6950)) or (layer2_outputs(3078));
    layer3_outputs(5225) <= not(layer2_outputs(2272));
    layer3_outputs(5226) <= layer2_outputs(8110);
    layer3_outputs(5227) <= '1';
    layer3_outputs(5228) <= not(layer2_outputs(81));
    layer3_outputs(5229) <= (layer2_outputs(9757)) or (layer2_outputs(7443));
    layer3_outputs(5230) <= (layer2_outputs(1288)) and (layer2_outputs(7140));
    layer3_outputs(5231) <= (layer2_outputs(6713)) and not (layer2_outputs(8617));
    layer3_outputs(5232) <= (layer2_outputs(2063)) xor (layer2_outputs(10044));
    layer3_outputs(5233) <= layer2_outputs(4309);
    layer3_outputs(5234) <= not((layer2_outputs(4983)) or (layer2_outputs(1427)));
    layer3_outputs(5235) <= not(layer2_outputs(8104)) or (layer2_outputs(1702));
    layer3_outputs(5236) <= layer2_outputs(9206);
    layer3_outputs(5237) <= not((layer2_outputs(9666)) xor (layer2_outputs(7583)));
    layer3_outputs(5238) <= '1';
    layer3_outputs(5239) <= layer2_outputs(6693);
    layer3_outputs(5240) <= not(layer2_outputs(7384)) or (layer2_outputs(7308));
    layer3_outputs(5241) <= layer2_outputs(3412);
    layer3_outputs(5242) <= (layer2_outputs(9386)) and not (layer2_outputs(1566));
    layer3_outputs(5243) <= not((layer2_outputs(2055)) xor (layer2_outputs(7219)));
    layer3_outputs(5244) <= layer2_outputs(6270);
    layer3_outputs(5245) <= not((layer2_outputs(4513)) and (layer2_outputs(1869)));
    layer3_outputs(5246) <= not(layer2_outputs(8811)) or (layer2_outputs(3731));
    layer3_outputs(5247) <= layer2_outputs(3624);
    layer3_outputs(5248) <= not(layer2_outputs(4443)) or (layer2_outputs(4818));
    layer3_outputs(5249) <= layer2_outputs(3061);
    layer3_outputs(5250) <= not(layer2_outputs(8774));
    layer3_outputs(5251) <= not(layer2_outputs(1632));
    layer3_outputs(5252) <= not(layer2_outputs(7563)) or (layer2_outputs(1902));
    layer3_outputs(5253) <= not(layer2_outputs(6046));
    layer3_outputs(5254) <= '1';
    layer3_outputs(5255) <= (layer2_outputs(8661)) and not (layer2_outputs(1408));
    layer3_outputs(5256) <= layer2_outputs(3000);
    layer3_outputs(5257) <= not(layer2_outputs(7203));
    layer3_outputs(5258) <= (layer2_outputs(5473)) or (layer2_outputs(10222));
    layer3_outputs(5259) <= not((layer2_outputs(5723)) xor (layer2_outputs(5402)));
    layer3_outputs(5260) <= layer2_outputs(4444);
    layer3_outputs(5261) <= '1';
    layer3_outputs(5262) <= not((layer2_outputs(8134)) and (layer2_outputs(925)));
    layer3_outputs(5263) <= not(layer2_outputs(6073));
    layer3_outputs(5264) <= layer2_outputs(3569);
    layer3_outputs(5265) <= (layer2_outputs(1764)) and (layer2_outputs(10078));
    layer3_outputs(5266) <= not((layer2_outputs(5505)) xor (layer2_outputs(3715)));
    layer3_outputs(5267) <= (layer2_outputs(7799)) xor (layer2_outputs(6354));
    layer3_outputs(5268) <= (layer2_outputs(2475)) xor (layer2_outputs(2956));
    layer3_outputs(5269) <= not((layer2_outputs(5257)) xor (layer2_outputs(7408)));
    layer3_outputs(5270) <= (layer2_outputs(671)) xor (layer2_outputs(2854));
    layer3_outputs(5271) <= not((layer2_outputs(8991)) or (layer2_outputs(9274)));
    layer3_outputs(5272) <= layer2_outputs(4201);
    layer3_outputs(5273) <= not(layer2_outputs(3728)) or (layer2_outputs(4373));
    layer3_outputs(5274) <= '1';
    layer3_outputs(5275) <= (layer2_outputs(484)) and not (layer2_outputs(5322));
    layer3_outputs(5276) <= layer2_outputs(910);
    layer3_outputs(5277) <= not(layer2_outputs(7663));
    layer3_outputs(5278) <= not(layer2_outputs(1170)) or (layer2_outputs(885));
    layer3_outputs(5279) <= layer2_outputs(4888);
    layer3_outputs(5280) <= not(layer2_outputs(9796)) or (layer2_outputs(6764));
    layer3_outputs(5281) <= not(layer2_outputs(5606));
    layer3_outputs(5282) <= not(layer2_outputs(1179));
    layer3_outputs(5283) <= layer2_outputs(2172);
    layer3_outputs(5284) <= not(layer2_outputs(1377));
    layer3_outputs(5285) <= not((layer2_outputs(6921)) and (layer2_outputs(8291)));
    layer3_outputs(5286) <= not(layer2_outputs(2870)) or (layer2_outputs(8164));
    layer3_outputs(5287) <= (layer2_outputs(6476)) or (layer2_outputs(4805));
    layer3_outputs(5288) <= not((layer2_outputs(3544)) and (layer2_outputs(5516)));
    layer3_outputs(5289) <= layer2_outputs(9372);
    layer3_outputs(5290) <= not(layer2_outputs(1626));
    layer3_outputs(5291) <= layer2_outputs(7667);
    layer3_outputs(5292) <= '1';
    layer3_outputs(5293) <= (layer2_outputs(9634)) and not (layer2_outputs(4934));
    layer3_outputs(5294) <= not(layer2_outputs(171));
    layer3_outputs(5295) <= layer2_outputs(9228);
    layer3_outputs(5296) <= not((layer2_outputs(1941)) or (layer2_outputs(4547)));
    layer3_outputs(5297) <= layer2_outputs(8504);
    layer3_outputs(5298) <= (layer2_outputs(6830)) xor (layer2_outputs(3891));
    layer3_outputs(5299) <= not(layer2_outputs(16)) or (layer2_outputs(9121));
    layer3_outputs(5300) <= not(layer2_outputs(804)) or (layer2_outputs(3977));
    layer3_outputs(5301) <= layer2_outputs(704);
    layer3_outputs(5302) <= (layer2_outputs(9192)) or (layer2_outputs(591));
    layer3_outputs(5303) <= layer2_outputs(3000);
    layer3_outputs(5304) <= not((layer2_outputs(1841)) and (layer2_outputs(6660)));
    layer3_outputs(5305) <= (layer2_outputs(2192)) and not (layer2_outputs(8469));
    layer3_outputs(5306) <= layer2_outputs(2530);
    layer3_outputs(5307) <= not(layer2_outputs(9136));
    layer3_outputs(5308) <= not((layer2_outputs(2046)) and (layer2_outputs(10176)));
    layer3_outputs(5309) <= (layer2_outputs(5012)) xor (layer2_outputs(6788));
    layer3_outputs(5310) <= not(layer2_outputs(2697)) or (layer2_outputs(6448));
    layer3_outputs(5311) <= not(layer2_outputs(8275));
    layer3_outputs(5312) <= not((layer2_outputs(2615)) and (layer2_outputs(5339)));
    layer3_outputs(5313) <= not(layer2_outputs(3556));
    layer3_outputs(5314) <= not(layer2_outputs(9130));
    layer3_outputs(5315) <= layer2_outputs(4323);
    layer3_outputs(5316) <= not(layer2_outputs(2930));
    layer3_outputs(5317) <= not((layer2_outputs(9969)) or (layer2_outputs(5235)));
    layer3_outputs(5318) <= not((layer2_outputs(9432)) xor (layer2_outputs(8578)));
    layer3_outputs(5319) <= not(layer2_outputs(8092));
    layer3_outputs(5320) <= not(layer2_outputs(128)) or (layer2_outputs(5919));
    layer3_outputs(5321) <= not(layer2_outputs(9295));
    layer3_outputs(5322) <= (layer2_outputs(8361)) and (layer2_outputs(4938));
    layer3_outputs(5323) <= not((layer2_outputs(7540)) xor (layer2_outputs(2384)));
    layer3_outputs(5324) <= (layer2_outputs(302)) and not (layer2_outputs(5096));
    layer3_outputs(5325) <= not(layer2_outputs(2805));
    layer3_outputs(5326) <= layer2_outputs(8107);
    layer3_outputs(5327) <= layer2_outputs(8079);
    layer3_outputs(5328) <= not((layer2_outputs(690)) xor (layer2_outputs(5780)));
    layer3_outputs(5329) <= (layer2_outputs(6194)) or (layer2_outputs(2699));
    layer3_outputs(5330) <= not(layer2_outputs(8264));
    layer3_outputs(5331) <= not(layer2_outputs(3028));
    layer3_outputs(5332) <= not(layer2_outputs(1477)) or (layer2_outputs(9677));
    layer3_outputs(5333) <= (layer2_outputs(6549)) xor (layer2_outputs(7896));
    layer3_outputs(5334) <= not(layer2_outputs(7185));
    layer3_outputs(5335) <= not((layer2_outputs(5473)) or (layer2_outputs(7659)));
    layer3_outputs(5336) <= layer2_outputs(7869);
    layer3_outputs(5337) <= not(layer2_outputs(6839));
    layer3_outputs(5338) <= not(layer2_outputs(3750)) or (layer2_outputs(2684));
    layer3_outputs(5339) <= layer2_outputs(7561);
    layer3_outputs(5340) <= not((layer2_outputs(4160)) and (layer2_outputs(1992)));
    layer3_outputs(5341) <= (layer2_outputs(5155)) xor (layer2_outputs(1448));
    layer3_outputs(5342) <= not((layer2_outputs(8571)) and (layer2_outputs(6401)));
    layer3_outputs(5343) <= not((layer2_outputs(1397)) xor (layer2_outputs(2918)));
    layer3_outputs(5344) <= '1';
    layer3_outputs(5345) <= not(layer2_outputs(2407));
    layer3_outputs(5346) <= not(layer2_outputs(6005));
    layer3_outputs(5347) <= (layer2_outputs(3492)) and (layer2_outputs(2305));
    layer3_outputs(5348) <= not((layer2_outputs(7016)) xor (layer2_outputs(2857)));
    layer3_outputs(5349) <= (layer2_outputs(5240)) and not (layer2_outputs(1058));
    layer3_outputs(5350) <= (layer2_outputs(2912)) or (layer2_outputs(8687));
    layer3_outputs(5351) <= layer2_outputs(5175);
    layer3_outputs(5352) <= not(layer2_outputs(7225));
    layer3_outputs(5353) <= (layer2_outputs(9911)) and not (layer2_outputs(3009));
    layer3_outputs(5354) <= layer2_outputs(6870);
    layer3_outputs(5355) <= (layer2_outputs(9087)) or (layer2_outputs(5093));
    layer3_outputs(5356) <= not((layer2_outputs(1543)) or (layer2_outputs(7267)));
    layer3_outputs(5357) <= layer2_outputs(3086);
    layer3_outputs(5358) <= '1';
    layer3_outputs(5359) <= layer2_outputs(4246);
    layer3_outputs(5360) <= not(layer2_outputs(2946)) or (layer2_outputs(292));
    layer3_outputs(5361) <= not(layer2_outputs(6617)) or (layer2_outputs(3059));
    layer3_outputs(5362) <= not(layer2_outputs(2852));
    layer3_outputs(5363) <= layer2_outputs(1127);
    layer3_outputs(5364) <= not(layer2_outputs(7760));
    layer3_outputs(5365) <= layer2_outputs(8500);
    layer3_outputs(5366) <= not(layer2_outputs(108));
    layer3_outputs(5367) <= layer2_outputs(4996);
    layer3_outputs(5368) <= '1';
    layer3_outputs(5369) <= not(layer2_outputs(1878));
    layer3_outputs(5370) <= not(layer2_outputs(5481)) or (layer2_outputs(3337));
    layer3_outputs(5371) <= not(layer2_outputs(4736)) or (layer2_outputs(6487));
    layer3_outputs(5372) <= (layer2_outputs(3577)) xor (layer2_outputs(6082));
    layer3_outputs(5373) <= (layer2_outputs(3730)) or (layer2_outputs(7843));
    layer3_outputs(5374) <= not(layer2_outputs(282));
    layer3_outputs(5375) <= not((layer2_outputs(1228)) or (layer2_outputs(6427)));
    layer3_outputs(5376) <= (layer2_outputs(7320)) xor (layer2_outputs(7241));
    layer3_outputs(5377) <= not(layer2_outputs(4063));
    layer3_outputs(5378) <= not((layer2_outputs(1743)) xor (layer2_outputs(5711)));
    layer3_outputs(5379) <= not((layer2_outputs(7816)) or (layer2_outputs(163)));
    layer3_outputs(5380) <= layer2_outputs(861);
    layer3_outputs(5381) <= not(layer2_outputs(2017));
    layer3_outputs(5382) <= (layer2_outputs(5507)) or (layer2_outputs(6795));
    layer3_outputs(5383) <= not(layer2_outputs(4713));
    layer3_outputs(5384) <= '1';
    layer3_outputs(5385) <= not((layer2_outputs(3688)) and (layer2_outputs(5875)));
    layer3_outputs(5386) <= not(layer2_outputs(6666));
    layer3_outputs(5387) <= '1';
    layer3_outputs(5388) <= not(layer2_outputs(7340));
    layer3_outputs(5389) <= layer2_outputs(3613);
    layer3_outputs(5390) <= not(layer2_outputs(9831));
    layer3_outputs(5391) <= layer2_outputs(4956);
    layer3_outputs(5392) <= not(layer2_outputs(1786));
    layer3_outputs(5393) <= '0';
    layer3_outputs(5394) <= (layer2_outputs(3946)) or (layer2_outputs(4440));
    layer3_outputs(5395) <= not(layer2_outputs(5292));
    layer3_outputs(5396) <= layer2_outputs(3390);
    layer3_outputs(5397) <= layer2_outputs(4927);
    layer3_outputs(5398) <= not(layer2_outputs(6420));
    layer3_outputs(5399) <= (layer2_outputs(1538)) and (layer2_outputs(1358));
    layer3_outputs(5400) <= (layer2_outputs(6580)) xor (layer2_outputs(4169));
    layer3_outputs(5401) <= not((layer2_outputs(5944)) xor (layer2_outputs(9984)));
    layer3_outputs(5402) <= layer2_outputs(6321);
    layer3_outputs(5403) <= layer2_outputs(9623);
    layer3_outputs(5404) <= not((layer2_outputs(7741)) xor (layer2_outputs(4593)));
    layer3_outputs(5405) <= layer2_outputs(9213);
    layer3_outputs(5406) <= not(layer2_outputs(1738)) or (layer2_outputs(3432));
    layer3_outputs(5407) <= not(layer2_outputs(6566));
    layer3_outputs(5408) <= layer2_outputs(1806);
    layer3_outputs(5409) <= layer2_outputs(4427);
    layer3_outputs(5410) <= (layer2_outputs(50)) or (layer2_outputs(1883));
    layer3_outputs(5411) <= not(layer2_outputs(868));
    layer3_outputs(5412) <= not(layer2_outputs(7929));
    layer3_outputs(5413) <= not((layer2_outputs(3866)) or (layer2_outputs(4880)));
    layer3_outputs(5414) <= not(layer2_outputs(627));
    layer3_outputs(5415) <= layer2_outputs(8222);
    layer3_outputs(5416) <= not(layer2_outputs(3650));
    layer3_outputs(5417) <= layer2_outputs(5454);
    layer3_outputs(5418) <= not(layer2_outputs(244));
    layer3_outputs(5419) <= (layer2_outputs(9002)) xor (layer2_outputs(4995));
    layer3_outputs(5420) <= layer2_outputs(3547);
    layer3_outputs(5421) <= not(layer2_outputs(5370));
    layer3_outputs(5422) <= not(layer2_outputs(8017));
    layer3_outputs(5423) <= not(layer2_outputs(4158));
    layer3_outputs(5424) <= layer2_outputs(9026);
    layer3_outputs(5425) <= not(layer2_outputs(8368)) or (layer2_outputs(8329));
    layer3_outputs(5426) <= (layer2_outputs(8587)) and not (layer2_outputs(9458));
    layer3_outputs(5427) <= (layer2_outputs(7694)) and not (layer2_outputs(3974));
    layer3_outputs(5428) <= (layer2_outputs(8315)) and (layer2_outputs(5784));
    layer3_outputs(5429) <= not((layer2_outputs(1186)) or (layer2_outputs(4171)));
    layer3_outputs(5430) <= layer2_outputs(2813);
    layer3_outputs(5431) <= '1';
    layer3_outputs(5432) <= not(layer2_outputs(1603));
    layer3_outputs(5433) <= layer2_outputs(8167);
    layer3_outputs(5434) <= (layer2_outputs(4141)) or (layer2_outputs(3189));
    layer3_outputs(5435) <= '0';
    layer3_outputs(5436) <= (layer2_outputs(4204)) and (layer2_outputs(8194));
    layer3_outputs(5437) <= '0';
    layer3_outputs(5438) <= layer2_outputs(6130);
    layer3_outputs(5439) <= not(layer2_outputs(9395)) or (layer2_outputs(9237));
    layer3_outputs(5440) <= layer2_outputs(4387);
    layer3_outputs(5441) <= not(layer2_outputs(2771));
    layer3_outputs(5442) <= not(layer2_outputs(7681));
    layer3_outputs(5443) <= (layer2_outputs(2509)) and not (layer2_outputs(443));
    layer3_outputs(5444) <= (layer2_outputs(7183)) and not (layer2_outputs(1244));
    layer3_outputs(5445) <= not((layer2_outputs(3538)) xor (layer2_outputs(569)));
    layer3_outputs(5446) <= (layer2_outputs(9339)) xor (layer2_outputs(383));
    layer3_outputs(5447) <= (layer2_outputs(2073)) and not (layer2_outputs(5086));
    layer3_outputs(5448) <= layer2_outputs(9620);
    layer3_outputs(5449) <= (layer2_outputs(5294)) and not (layer2_outputs(9675));
    layer3_outputs(5450) <= (layer2_outputs(4506)) xor (layer2_outputs(179));
    layer3_outputs(5451) <= not((layer2_outputs(2997)) or (layer2_outputs(4530)));
    layer3_outputs(5452) <= (layer2_outputs(2961)) and not (layer2_outputs(7473));
    layer3_outputs(5453) <= layer2_outputs(403);
    layer3_outputs(5454) <= not(layer2_outputs(5312));
    layer3_outputs(5455) <= (layer2_outputs(6060)) or (layer2_outputs(392));
    layer3_outputs(5456) <= not(layer2_outputs(9183)) or (layer2_outputs(2685));
    layer3_outputs(5457) <= not(layer2_outputs(6218));
    layer3_outputs(5458) <= layer2_outputs(9122);
    layer3_outputs(5459) <= (layer2_outputs(1455)) xor (layer2_outputs(9927));
    layer3_outputs(5460) <= (layer2_outputs(4932)) and (layer2_outputs(9288));
    layer3_outputs(5461) <= layer2_outputs(6435);
    layer3_outputs(5462) <= (layer2_outputs(6259)) and not (layer2_outputs(1774));
    layer3_outputs(5463) <= (layer2_outputs(1439)) and not (layer2_outputs(6230));
    layer3_outputs(5464) <= not(layer2_outputs(9703)) or (layer2_outputs(9373));
    layer3_outputs(5465) <= layer2_outputs(7549);
    layer3_outputs(5466) <= (layer2_outputs(9199)) xor (layer2_outputs(862));
    layer3_outputs(5467) <= not(layer2_outputs(691));
    layer3_outputs(5468) <= layer2_outputs(4537);
    layer3_outputs(5469) <= '1';
    layer3_outputs(5470) <= not((layer2_outputs(7634)) xor (layer2_outputs(6727)));
    layer3_outputs(5471) <= not(layer2_outputs(4190));
    layer3_outputs(5472) <= not(layer2_outputs(6918));
    layer3_outputs(5473) <= (layer2_outputs(4727)) xor (layer2_outputs(9060));
    layer3_outputs(5474) <= layer2_outputs(7656);
    layer3_outputs(5475) <= layer2_outputs(2417);
    layer3_outputs(5476) <= not(layer2_outputs(9475));
    layer3_outputs(5477) <= not((layer2_outputs(2550)) or (layer2_outputs(3824)));
    layer3_outputs(5478) <= (layer2_outputs(10004)) xor (layer2_outputs(6423));
    layer3_outputs(5479) <= not((layer2_outputs(5437)) xor (layer2_outputs(5560)));
    layer3_outputs(5480) <= (layer2_outputs(8878)) and not (layer2_outputs(1454));
    layer3_outputs(5481) <= not(layer2_outputs(10154)) or (layer2_outputs(934));
    layer3_outputs(5482) <= not(layer2_outputs(7898));
    layer3_outputs(5483) <= not((layer2_outputs(6923)) xor (layer2_outputs(1795)));
    layer3_outputs(5484) <= layer2_outputs(4184);
    layer3_outputs(5485) <= not(layer2_outputs(5156));
    layer3_outputs(5486) <= (layer2_outputs(647)) xor (layer2_outputs(2139));
    layer3_outputs(5487) <= (layer2_outputs(6778)) and not (layer2_outputs(4302));
    layer3_outputs(5488) <= layer2_outputs(8448);
    layer3_outputs(5489) <= not(layer2_outputs(2526)) or (layer2_outputs(7533));
    layer3_outputs(5490) <= not(layer2_outputs(8857)) or (layer2_outputs(3595));
    layer3_outputs(5491) <= (layer2_outputs(1746)) and not (layer2_outputs(6790));
    layer3_outputs(5492) <= layer2_outputs(1391);
    layer3_outputs(5493) <= (layer2_outputs(2730)) and (layer2_outputs(3053));
    layer3_outputs(5494) <= layer2_outputs(4474);
    layer3_outputs(5495) <= not(layer2_outputs(7914));
    layer3_outputs(5496) <= layer2_outputs(7102);
    layer3_outputs(5497) <= layer2_outputs(792);
    layer3_outputs(5498) <= (layer2_outputs(3760)) xor (layer2_outputs(9418));
    layer3_outputs(5499) <= not(layer2_outputs(7888));
    layer3_outputs(5500) <= (layer2_outputs(6978)) and (layer2_outputs(6818));
    layer3_outputs(5501) <= (layer2_outputs(6901)) and not (layer2_outputs(6821));
    layer3_outputs(5502) <= not(layer2_outputs(7068)) or (layer2_outputs(6041));
    layer3_outputs(5503) <= not(layer2_outputs(1253));
    layer3_outputs(5504) <= not((layer2_outputs(2626)) and (layer2_outputs(5289)));
    layer3_outputs(5505) <= not((layer2_outputs(5159)) and (layer2_outputs(495)));
    layer3_outputs(5506) <= not((layer2_outputs(8711)) xor (layer2_outputs(3674)));
    layer3_outputs(5507) <= (layer2_outputs(7104)) and not (layer2_outputs(2669));
    layer3_outputs(5508) <= (layer2_outputs(5882)) xor (layer2_outputs(7790));
    layer3_outputs(5509) <= not((layer2_outputs(872)) or (layer2_outputs(2815)));
    layer3_outputs(5510) <= (layer2_outputs(2486)) and not (layer2_outputs(4006));
    layer3_outputs(5511) <= (layer2_outputs(3007)) and not (layer2_outputs(6419));
    layer3_outputs(5512) <= (layer2_outputs(9029)) and not (layer2_outputs(9580));
    layer3_outputs(5513) <= not(layer2_outputs(2064));
    layer3_outputs(5514) <= not(layer2_outputs(1767));
    layer3_outputs(5515) <= not(layer2_outputs(7398));
    layer3_outputs(5516) <= not(layer2_outputs(8087));
    layer3_outputs(5517) <= not((layer2_outputs(2413)) and (layer2_outputs(5127)));
    layer3_outputs(5518) <= (layer2_outputs(9584)) and not (layer2_outputs(7494));
    layer3_outputs(5519) <= (layer2_outputs(5234)) xor (layer2_outputs(1164));
    layer3_outputs(5520) <= (layer2_outputs(5068)) or (layer2_outputs(489));
    layer3_outputs(5521) <= not(layer2_outputs(3966)) or (layer2_outputs(823));
    layer3_outputs(5522) <= (layer2_outputs(5362)) and (layer2_outputs(3882));
    layer3_outputs(5523) <= (layer2_outputs(4560)) xor (layer2_outputs(9863));
    layer3_outputs(5524) <= (layer2_outputs(6227)) and not (layer2_outputs(4481));
    layer3_outputs(5525) <= layer2_outputs(1853);
    layer3_outputs(5526) <= not(layer2_outputs(8946));
    layer3_outputs(5527) <= (layer2_outputs(6015)) and not (layer2_outputs(6432));
    layer3_outputs(5528) <= layer2_outputs(10054);
    layer3_outputs(5529) <= layer2_outputs(8456);
    layer3_outputs(5530) <= not(layer2_outputs(3463));
    layer3_outputs(5531) <= not(layer2_outputs(8356));
    layer3_outputs(5532) <= not(layer2_outputs(2889));
    layer3_outputs(5533) <= not(layer2_outputs(8657));
    layer3_outputs(5534) <= layer2_outputs(6829);
    layer3_outputs(5535) <= '1';
    layer3_outputs(5536) <= not(layer2_outputs(206)) or (layer2_outputs(8978));
    layer3_outputs(5537) <= layer2_outputs(6439);
    layer3_outputs(5538) <= not((layer2_outputs(7833)) or (layer2_outputs(3237)));
    layer3_outputs(5539) <= layer2_outputs(6992);
    layer3_outputs(5540) <= not(layer2_outputs(9156));
    layer3_outputs(5541) <= not(layer2_outputs(7750)) or (layer2_outputs(7592));
    layer3_outputs(5542) <= layer2_outputs(1700);
    layer3_outputs(5543) <= (layer2_outputs(10139)) and not (layer2_outputs(9785));
    layer3_outputs(5544) <= not(layer2_outputs(3882));
    layer3_outputs(5545) <= not((layer2_outputs(2814)) and (layer2_outputs(7144)));
    layer3_outputs(5546) <= not(layer2_outputs(3596));
    layer3_outputs(5547) <= layer2_outputs(5039);
    layer3_outputs(5548) <= not(layer2_outputs(8689));
    layer3_outputs(5549) <= not(layer2_outputs(4657)) or (layer2_outputs(674));
    layer3_outputs(5550) <= not(layer2_outputs(4925));
    layer3_outputs(5551) <= not(layer2_outputs(8178));
    layer3_outputs(5552) <= layer2_outputs(4924);
    layer3_outputs(5553) <= layer2_outputs(3593);
    layer3_outputs(5554) <= (layer2_outputs(9829)) and not (layer2_outputs(8634));
    layer3_outputs(5555) <= (layer2_outputs(5715)) and not (layer2_outputs(2880));
    layer3_outputs(5556) <= not((layer2_outputs(1231)) xor (layer2_outputs(8730)));
    layer3_outputs(5557) <= layer2_outputs(10097);
    layer3_outputs(5558) <= layer2_outputs(7448);
    layer3_outputs(5559) <= '0';
    layer3_outputs(5560) <= not((layer2_outputs(1381)) xor (layer2_outputs(7316)));
    layer3_outputs(5561) <= (layer2_outputs(5439)) and (layer2_outputs(4024));
    layer3_outputs(5562) <= (layer2_outputs(328)) xor (layer2_outputs(9668));
    layer3_outputs(5563) <= (layer2_outputs(3436)) and not (layer2_outputs(1852));
    layer3_outputs(5564) <= (layer2_outputs(5900)) and not (layer2_outputs(8894));
    layer3_outputs(5565) <= not((layer2_outputs(1582)) xor (layer2_outputs(2761)));
    layer3_outputs(5566) <= not((layer2_outputs(243)) xor (layer2_outputs(3417)));
    layer3_outputs(5567) <= not((layer2_outputs(4230)) and (layer2_outputs(7339)));
    layer3_outputs(5568) <= (layer2_outputs(255)) xor (layer2_outputs(2747));
    layer3_outputs(5569) <= not(layer2_outputs(5818));
    layer3_outputs(5570) <= not((layer2_outputs(5128)) xor (layer2_outputs(5506)));
    layer3_outputs(5571) <= not(layer2_outputs(6835));
    layer3_outputs(5572) <= (layer2_outputs(413)) and not (layer2_outputs(6458));
    layer3_outputs(5573) <= not((layer2_outputs(848)) xor (layer2_outputs(6342)));
    layer3_outputs(5574) <= not((layer2_outputs(4972)) and (layer2_outputs(6768)));
    layer3_outputs(5575) <= not(layer2_outputs(9763));
    layer3_outputs(5576) <= layer2_outputs(7747);
    layer3_outputs(5577) <= (layer2_outputs(9454)) or (layer2_outputs(1468));
    layer3_outputs(5578) <= (layer2_outputs(5356)) and (layer2_outputs(5575));
    layer3_outputs(5579) <= layer2_outputs(9918);
    layer3_outputs(5580) <= not(layer2_outputs(6550));
    layer3_outputs(5581) <= (layer2_outputs(5448)) and (layer2_outputs(7738));
    layer3_outputs(5582) <= layer2_outputs(6991);
    layer3_outputs(5583) <= layer2_outputs(5151);
    layer3_outputs(5584) <= not(layer2_outputs(1573));
    layer3_outputs(5585) <= (layer2_outputs(3468)) and (layer2_outputs(6974));
    layer3_outputs(5586) <= not(layer2_outputs(7968));
    layer3_outputs(5587) <= layer2_outputs(839);
    layer3_outputs(5588) <= layer2_outputs(1508);
    layer3_outputs(5589) <= not(layer2_outputs(4463));
    layer3_outputs(5590) <= not(layer2_outputs(1551));
    layer3_outputs(5591) <= '0';
    layer3_outputs(5592) <= layer2_outputs(7562);
    layer3_outputs(5593) <= (layer2_outputs(4999)) or (layer2_outputs(4014));
    layer3_outputs(5594) <= layer2_outputs(9898);
    layer3_outputs(5595) <= not(layer2_outputs(5896));
    layer3_outputs(5596) <= (layer2_outputs(590)) xor (layer2_outputs(386));
    layer3_outputs(5597) <= not(layer2_outputs(4327));
    layer3_outputs(5598) <= layer2_outputs(6570);
    layer3_outputs(5599) <= (layer2_outputs(9552)) or (layer2_outputs(3402));
    layer3_outputs(5600) <= not(layer2_outputs(6482));
    layer3_outputs(5601) <= not(layer2_outputs(9262));
    layer3_outputs(5602) <= not(layer2_outputs(356)) or (layer2_outputs(4130));
    layer3_outputs(5603) <= not(layer2_outputs(5268));
    layer3_outputs(5604) <= (layer2_outputs(155)) or (layer2_outputs(3383));
    layer3_outputs(5605) <= (layer2_outputs(6380)) and (layer2_outputs(8443));
    layer3_outputs(5606) <= (layer2_outputs(3210)) and not (layer2_outputs(188));
    layer3_outputs(5607) <= not(layer2_outputs(9210)) or (layer2_outputs(5135));
    layer3_outputs(5608) <= not(layer2_outputs(3843));
    layer3_outputs(5609) <= not(layer2_outputs(8266));
    layer3_outputs(5610) <= not(layer2_outputs(5198));
    layer3_outputs(5611) <= not(layer2_outputs(10009));
    layer3_outputs(5612) <= layer2_outputs(6848);
    layer3_outputs(5613) <= (layer2_outputs(802)) and not (layer2_outputs(4060));
    layer3_outputs(5614) <= layer2_outputs(8171);
    layer3_outputs(5615) <= not(layer2_outputs(4366)) or (layer2_outputs(6442));
    layer3_outputs(5616) <= not(layer2_outputs(8447));
    layer3_outputs(5617) <= (layer2_outputs(839)) xor (layer2_outputs(10019));
    layer3_outputs(5618) <= (layer2_outputs(9595)) or (layer2_outputs(8818));
    layer3_outputs(5619) <= layer2_outputs(6786);
    layer3_outputs(5620) <= (layer2_outputs(1643)) or (layer2_outputs(1926));
    layer3_outputs(5621) <= layer2_outputs(4347);
    layer3_outputs(5622) <= (layer2_outputs(7668)) and not (layer2_outputs(8094));
    layer3_outputs(5623) <= not((layer2_outputs(3867)) or (layer2_outputs(1874)));
    layer3_outputs(5624) <= (layer2_outputs(9131)) and not (layer2_outputs(9022));
    layer3_outputs(5625) <= not(layer2_outputs(10200));
    layer3_outputs(5626) <= layer2_outputs(941);
    layer3_outputs(5627) <= (layer2_outputs(2460)) and not (layer2_outputs(2053));
    layer3_outputs(5628) <= not(layer2_outputs(2604));
    layer3_outputs(5629) <= not(layer2_outputs(6423));
    layer3_outputs(5630) <= not((layer2_outputs(2869)) xor (layer2_outputs(8334)));
    layer3_outputs(5631) <= (layer2_outputs(10038)) and not (layer2_outputs(8031));
    layer3_outputs(5632) <= (layer2_outputs(2384)) and not (layer2_outputs(4603));
    layer3_outputs(5633) <= '0';
    layer3_outputs(5634) <= not(layer2_outputs(7227)) or (layer2_outputs(3181));
    layer3_outputs(5635) <= not(layer2_outputs(4990));
    layer3_outputs(5636) <= (layer2_outputs(4755)) and (layer2_outputs(3756));
    layer3_outputs(5637) <= not(layer2_outputs(6903));
    layer3_outputs(5638) <= layer2_outputs(9619);
    layer3_outputs(5639) <= (layer2_outputs(9091)) or (layer2_outputs(1565));
    layer3_outputs(5640) <= layer2_outputs(7472);
    layer3_outputs(5641) <= layer2_outputs(7415);
    layer3_outputs(5642) <= '0';
    layer3_outputs(5643) <= not(layer2_outputs(3910));
    layer3_outputs(5644) <= not(layer2_outputs(9891));
    layer3_outputs(5645) <= not((layer2_outputs(7646)) xor (layer2_outputs(10206)));
    layer3_outputs(5646) <= layer2_outputs(6309);
    layer3_outputs(5647) <= not(layer2_outputs(7890));
    layer3_outputs(5648) <= not(layer2_outputs(2519));
    layer3_outputs(5649) <= not((layer2_outputs(8080)) or (layer2_outputs(1760)));
    layer3_outputs(5650) <= not(layer2_outputs(5513));
    layer3_outputs(5651) <= not(layer2_outputs(8063)) or (layer2_outputs(7479));
    layer3_outputs(5652) <= layer2_outputs(9287);
    layer3_outputs(5653) <= (layer2_outputs(2640)) xor (layer2_outputs(1384));
    layer3_outputs(5654) <= (layer2_outputs(6709)) and not (layer2_outputs(2919));
    layer3_outputs(5655) <= not(layer2_outputs(3290)) or (layer2_outputs(7041));
    layer3_outputs(5656) <= not(layer2_outputs(9142));
    layer3_outputs(5657) <= not((layer2_outputs(7499)) and (layer2_outputs(1884)));
    layer3_outputs(5658) <= not((layer2_outputs(6479)) or (layer2_outputs(2922)));
    layer3_outputs(5659) <= (layer2_outputs(6332)) or (layer2_outputs(4427));
    layer3_outputs(5660) <= not(layer2_outputs(8100));
    layer3_outputs(5661) <= not(layer2_outputs(3314)) or (layer2_outputs(4365));
    layer3_outputs(5662) <= layer2_outputs(9571);
    layer3_outputs(5663) <= not(layer2_outputs(1261)) or (layer2_outputs(1553));
    layer3_outputs(5664) <= (layer2_outputs(5735)) or (layer2_outputs(101));
    layer3_outputs(5665) <= (layer2_outputs(1182)) and (layer2_outputs(5631));
    layer3_outputs(5666) <= layer2_outputs(398);
    layer3_outputs(5667) <= not(layer2_outputs(1018));
    layer3_outputs(5668) <= not(layer2_outputs(2678)) or (layer2_outputs(1820));
    layer3_outputs(5669) <= not((layer2_outputs(4936)) or (layer2_outputs(2884)));
    layer3_outputs(5670) <= not(layer2_outputs(3611));
    layer3_outputs(5671) <= not(layer2_outputs(6493)) or (layer2_outputs(1041));
    layer3_outputs(5672) <= (layer2_outputs(6141)) or (layer2_outputs(7550));
    layer3_outputs(5673) <= not(layer2_outputs(5739));
    layer3_outputs(5674) <= layer2_outputs(9149);
    layer3_outputs(5675) <= (layer2_outputs(4343)) or (layer2_outputs(8132));
    layer3_outputs(5676) <= not(layer2_outputs(4905));
    layer3_outputs(5677) <= not(layer2_outputs(5190));
    layer3_outputs(5678) <= (layer2_outputs(7598)) xor (layer2_outputs(5015));
    layer3_outputs(5679) <= not(layer2_outputs(5209));
    layer3_outputs(5680) <= not((layer2_outputs(6069)) and (layer2_outputs(5362)));
    layer3_outputs(5681) <= not(layer2_outputs(794));
    layer3_outputs(5682) <= not(layer2_outputs(10199));
    layer3_outputs(5683) <= layer2_outputs(6847);
    layer3_outputs(5684) <= not(layer2_outputs(5394));
    layer3_outputs(5685) <= (layer2_outputs(9925)) and (layer2_outputs(1700));
    layer3_outputs(5686) <= layer2_outputs(3522);
    layer3_outputs(5687) <= layer2_outputs(1148);
    layer3_outputs(5688) <= layer2_outputs(5854);
    layer3_outputs(5689) <= layer2_outputs(3679);
    layer3_outputs(5690) <= (layer2_outputs(2776)) and not (layer2_outputs(7315));
    layer3_outputs(5691) <= layer2_outputs(3737);
    layer3_outputs(5692) <= not(layer2_outputs(207));
    layer3_outputs(5693) <= layer2_outputs(2738);
    layer3_outputs(5694) <= not((layer2_outputs(3667)) or (layer2_outputs(9239)));
    layer3_outputs(5695) <= (layer2_outputs(2856)) and not (layer2_outputs(4912));
    layer3_outputs(5696) <= not(layer2_outputs(152));
    layer3_outputs(5697) <= (layer2_outputs(6928)) and (layer2_outputs(7538));
    layer3_outputs(5698) <= not(layer2_outputs(7512));
    layer3_outputs(5699) <= not((layer2_outputs(307)) and (layer2_outputs(385)));
    layer3_outputs(5700) <= layer2_outputs(4169);
    layer3_outputs(5701) <= not(layer2_outputs(9298));
    layer3_outputs(5702) <= layer2_outputs(7567);
    layer3_outputs(5703) <= (layer2_outputs(2006)) or (layer2_outputs(4339));
    layer3_outputs(5704) <= not(layer2_outputs(6610)) or (layer2_outputs(4088));
    layer3_outputs(5705) <= layer2_outputs(6763);
    layer3_outputs(5706) <= not(layer2_outputs(6155));
    layer3_outputs(5707) <= (layer2_outputs(8495)) and not (layer2_outputs(1973));
    layer3_outputs(5708) <= not(layer2_outputs(9063));
    layer3_outputs(5709) <= layer2_outputs(7170);
    layer3_outputs(5710) <= (layer2_outputs(5505)) and not (layer2_outputs(1310));
    layer3_outputs(5711) <= layer2_outputs(7595);
    layer3_outputs(5712) <= (layer2_outputs(6307)) and not (layer2_outputs(6137));
    layer3_outputs(5713) <= '1';
    layer3_outputs(5714) <= not(layer2_outputs(2996));
    layer3_outputs(5715) <= (layer2_outputs(9905)) and not (layer2_outputs(5227));
    layer3_outputs(5716) <= (layer2_outputs(4757)) and not (layer2_outputs(7254));
    layer3_outputs(5717) <= not(layer2_outputs(4011));
    layer3_outputs(5718) <= layer2_outputs(745);
    layer3_outputs(5719) <= '0';
    layer3_outputs(5720) <= not(layer2_outputs(7475));
    layer3_outputs(5721) <= (layer2_outputs(3730)) and (layer2_outputs(1819));
    layer3_outputs(5722) <= not(layer2_outputs(4942));
    layer3_outputs(5723) <= not((layer2_outputs(7640)) xor (layer2_outputs(439)));
    layer3_outputs(5724) <= not(layer2_outputs(8890));
    layer3_outputs(5725) <= not((layer2_outputs(5509)) or (layer2_outputs(1847)));
    layer3_outputs(5726) <= not((layer2_outputs(5542)) or (layer2_outputs(6649)));
    layer3_outputs(5727) <= (layer2_outputs(921)) xor (layer2_outputs(3529));
    layer3_outputs(5728) <= not(layer2_outputs(3265));
    layer3_outputs(5729) <= not(layer2_outputs(281));
    layer3_outputs(5730) <= not(layer2_outputs(5604)) or (layer2_outputs(2674));
    layer3_outputs(5731) <= (layer2_outputs(4923)) and not (layer2_outputs(2675));
    layer3_outputs(5732) <= not(layer2_outputs(919));
    layer3_outputs(5733) <= (layer2_outputs(2966)) and not (layer2_outputs(4875));
    layer3_outputs(5734) <= not(layer2_outputs(1858));
    layer3_outputs(5735) <= layer2_outputs(462);
    layer3_outputs(5736) <= not((layer2_outputs(10146)) xor (layer2_outputs(5874)));
    layer3_outputs(5737) <= (layer2_outputs(2281)) and not (layer2_outputs(9757));
    layer3_outputs(5738) <= layer2_outputs(8813);
    layer3_outputs(5739) <= layer2_outputs(4895);
    layer3_outputs(5740) <= (layer2_outputs(2927)) xor (layer2_outputs(3386));
    layer3_outputs(5741) <= (layer2_outputs(2553)) and (layer2_outputs(1122));
    layer3_outputs(5742) <= not((layer2_outputs(7236)) xor (layer2_outputs(8884)));
    layer3_outputs(5743) <= layer2_outputs(9828);
    layer3_outputs(5744) <= not(layer2_outputs(7990)) or (layer2_outputs(5931));
    layer3_outputs(5745) <= not(layer2_outputs(8239));
    layer3_outputs(5746) <= layer2_outputs(9224);
    layer3_outputs(5747) <= not((layer2_outputs(7877)) and (layer2_outputs(1936)));
    layer3_outputs(5748) <= layer2_outputs(3392);
    layer3_outputs(5749) <= not((layer2_outputs(8098)) xor (layer2_outputs(107)));
    layer3_outputs(5750) <= not((layer2_outputs(2618)) and (layer2_outputs(2862)));
    layer3_outputs(5751) <= (layer2_outputs(6370)) and (layer2_outputs(1470));
    layer3_outputs(5752) <= (layer2_outputs(2547)) xor (layer2_outputs(661));
    layer3_outputs(5753) <= not((layer2_outputs(6934)) and (layer2_outputs(1741)));
    layer3_outputs(5754) <= not((layer2_outputs(1521)) xor (layer2_outputs(3747)));
    layer3_outputs(5755) <= not((layer2_outputs(8213)) and (layer2_outputs(6603)));
    layer3_outputs(5756) <= not((layer2_outputs(5238)) and (layer2_outputs(8656)));
    layer3_outputs(5757) <= layer2_outputs(6059);
    layer3_outputs(5758) <= not(layer2_outputs(9225)) or (layer2_outputs(5907));
    layer3_outputs(5759) <= not((layer2_outputs(1917)) and (layer2_outputs(8540)));
    layer3_outputs(5760) <= not(layer2_outputs(5482));
    layer3_outputs(5761) <= not(layer2_outputs(4286));
    layer3_outputs(5762) <= not(layer2_outputs(3807));
    layer3_outputs(5763) <= layer2_outputs(5386);
    layer3_outputs(5764) <= (layer2_outputs(9973)) and not (layer2_outputs(649));
    layer3_outputs(5765) <= (layer2_outputs(41)) xor (layer2_outputs(630));
    layer3_outputs(5766) <= layer2_outputs(7579);
    layer3_outputs(5767) <= not(layer2_outputs(4967));
    layer3_outputs(5768) <= not(layer2_outputs(5387)) or (layer2_outputs(6108));
    layer3_outputs(5769) <= (layer2_outputs(136)) xor (layer2_outputs(1029));
    layer3_outputs(5770) <= layer2_outputs(3056);
    layer3_outputs(5771) <= not(layer2_outputs(10069));
    layer3_outputs(5772) <= layer2_outputs(7012);
    layer3_outputs(5773) <= not((layer2_outputs(1328)) or (layer2_outputs(9411)));
    layer3_outputs(5774) <= (layer2_outputs(3555)) xor (layer2_outputs(9036));
    layer3_outputs(5775) <= (layer2_outputs(10061)) and not (layer2_outputs(2531));
    layer3_outputs(5776) <= layer2_outputs(8911);
    layer3_outputs(5777) <= not(layer2_outputs(7152));
    layer3_outputs(5778) <= '0';
    layer3_outputs(5779) <= not(layer2_outputs(9509));
    layer3_outputs(5780) <= not((layer2_outputs(5912)) and (layer2_outputs(3222)));
    layer3_outputs(5781) <= '1';
    layer3_outputs(5782) <= not(layer2_outputs(6523));
    layer3_outputs(5783) <= (layer2_outputs(5279)) and (layer2_outputs(9877));
    layer3_outputs(5784) <= layer2_outputs(973);
    layer3_outputs(5785) <= (layer2_outputs(145)) xor (layer2_outputs(6883));
    layer3_outputs(5786) <= '1';
    layer3_outputs(5787) <= not(layer2_outputs(6001));
    layer3_outputs(5788) <= (layer2_outputs(2965)) or (layer2_outputs(4722));
    layer3_outputs(5789) <= layer2_outputs(7639);
    layer3_outputs(5790) <= layer2_outputs(2473);
    layer3_outputs(5791) <= (layer2_outputs(9179)) and (layer2_outputs(78));
    layer3_outputs(5792) <= (layer2_outputs(5950)) xor (layer2_outputs(926));
    layer3_outputs(5793) <= not(layer2_outputs(2502));
    layer3_outputs(5794) <= not(layer2_outputs(1649));
    layer3_outputs(5795) <= layer2_outputs(8637);
    layer3_outputs(5796) <= not(layer2_outputs(10097));
    layer3_outputs(5797) <= not(layer2_outputs(3716));
    layer3_outputs(5798) <= (layer2_outputs(6378)) or (layer2_outputs(3777));
    layer3_outputs(5799) <= (layer2_outputs(9640)) and (layer2_outputs(6907));
    layer3_outputs(5800) <= not(layer2_outputs(1343));
    layer3_outputs(5801) <= not(layer2_outputs(10140));
    layer3_outputs(5802) <= not((layer2_outputs(9634)) or (layer2_outputs(3095)));
    layer3_outputs(5803) <= (layer2_outputs(467)) and not (layer2_outputs(9528));
    layer3_outputs(5804) <= '1';
    layer3_outputs(5805) <= layer2_outputs(2822);
    layer3_outputs(5806) <= (layer2_outputs(2167)) or (layer2_outputs(5895));
    layer3_outputs(5807) <= (layer2_outputs(5819)) and not (layer2_outputs(5877));
    layer3_outputs(5808) <= not((layer2_outputs(4667)) xor (layer2_outputs(9902)));
    layer3_outputs(5809) <= (layer2_outputs(10226)) and (layer2_outputs(5883));
    layer3_outputs(5810) <= not((layer2_outputs(7172)) xor (layer2_outputs(7930)));
    layer3_outputs(5811) <= layer2_outputs(1145);
    layer3_outputs(5812) <= (layer2_outputs(4704)) and not (layer2_outputs(8047));
    layer3_outputs(5813) <= not(layer2_outputs(3019));
    layer3_outputs(5814) <= layer2_outputs(3543);
    layer3_outputs(5815) <= not(layer2_outputs(6261));
    layer3_outputs(5816) <= (layer2_outputs(437)) and (layer2_outputs(6400));
    layer3_outputs(5817) <= (layer2_outputs(849)) xor (layer2_outputs(1745));
    layer3_outputs(5818) <= layer2_outputs(5361);
    layer3_outputs(5819) <= (layer2_outputs(5714)) and (layer2_outputs(4558));
    layer3_outputs(5820) <= (layer2_outputs(8018)) or (layer2_outputs(2198));
    layer3_outputs(5821) <= (layer2_outputs(1374)) and (layer2_outputs(4944));
    layer3_outputs(5822) <= layer2_outputs(9727);
    layer3_outputs(5823) <= not(layer2_outputs(958)) or (layer2_outputs(10193));
    layer3_outputs(5824) <= (layer2_outputs(3960)) and (layer2_outputs(8573));
    layer3_outputs(5825) <= not((layer2_outputs(3728)) xor (layer2_outputs(5134)));
    layer3_outputs(5826) <= layer2_outputs(6403);
    layer3_outputs(5827) <= not((layer2_outputs(8075)) xor (layer2_outputs(1940)));
    layer3_outputs(5828) <= not((layer2_outputs(5929)) or (layer2_outputs(2698)));
    layer3_outputs(5829) <= not(layer2_outputs(7606)) or (layer2_outputs(5930));
    layer3_outputs(5830) <= not(layer2_outputs(8926));
    layer3_outputs(5831) <= layer2_outputs(1407);
    layer3_outputs(5832) <= (layer2_outputs(7791)) xor (layer2_outputs(631));
    layer3_outputs(5833) <= not((layer2_outputs(1561)) xor (layer2_outputs(2135)));
    layer3_outputs(5834) <= not(layer2_outputs(941));
    layer3_outputs(5835) <= layer2_outputs(535);
    layer3_outputs(5836) <= layer2_outputs(5007);
    layer3_outputs(5837) <= (layer2_outputs(8396)) or (layer2_outputs(6822));
    layer3_outputs(5838) <= (layer2_outputs(1807)) and not (layer2_outputs(3495));
    layer3_outputs(5839) <= not((layer2_outputs(9740)) and (layer2_outputs(4745)));
    layer3_outputs(5840) <= layer2_outputs(1927);
    layer3_outputs(5841) <= not((layer2_outputs(5522)) xor (layer2_outputs(5281)));
    layer3_outputs(5842) <= not((layer2_outputs(5186)) xor (layer2_outputs(2752)));
    layer3_outputs(5843) <= layer2_outputs(6249);
    layer3_outputs(5844) <= '0';
    layer3_outputs(5845) <= (layer2_outputs(2400)) and not (layer2_outputs(4646));
    layer3_outputs(5846) <= layer2_outputs(6804);
    layer3_outputs(5847) <= not(layer2_outputs(8236));
    layer3_outputs(5848) <= not(layer2_outputs(5914));
    layer3_outputs(5849) <= not(layer2_outputs(3795));
    layer3_outputs(5850) <= not(layer2_outputs(2508));
    layer3_outputs(5851) <= not(layer2_outputs(8761));
    layer3_outputs(5852) <= (layer2_outputs(7921)) and not (layer2_outputs(4069));
    layer3_outputs(5853) <= not(layer2_outputs(2359));
    layer3_outputs(5854) <= not(layer2_outputs(404)) or (layer2_outputs(10085));
    layer3_outputs(5855) <= layer2_outputs(4455);
    layer3_outputs(5856) <= not(layer2_outputs(7505));
    layer3_outputs(5857) <= layer2_outputs(692);
    layer3_outputs(5858) <= not((layer2_outputs(1474)) or (layer2_outputs(6820)));
    layer3_outputs(5859) <= layer2_outputs(2157);
    layer3_outputs(5860) <= layer2_outputs(3642);
    layer3_outputs(5861) <= '1';
    layer3_outputs(5862) <= not(layer2_outputs(10213));
    layer3_outputs(5863) <= layer2_outputs(689);
    layer3_outputs(5864) <= not((layer2_outputs(5821)) and (layer2_outputs(244)));
    layer3_outputs(5865) <= (layer2_outputs(4376)) or (layer2_outputs(3489));
    layer3_outputs(5866) <= '1';
    layer3_outputs(5867) <= not(layer2_outputs(918));
    layer3_outputs(5868) <= (layer2_outputs(4660)) and (layer2_outputs(6112));
    layer3_outputs(5869) <= not(layer2_outputs(2436));
    layer3_outputs(5870) <= not(layer2_outputs(7398));
    layer3_outputs(5871) <= layer2_outputs(9610);
    layer3_outputs(5872) <= '0';
    layer3_outputs(5873) <= layer2_outputs(4670);
    layer3_outputs(5874) <= layer2_outputs(3157);
    layer3_outputs(5875) <= (layer2_outputs(6819)) and not (layer2_outputs(3926));
    layer3_outputs(5876) <= (layer2_outputs(8215)) or (layer2_outputs(6690));
    layer3_outputs(5877) <= not(layer2_outputs(7815));
    layer3_outputs(5878) <= not((layer2_outputs(8362)) or (layer2_outputs(5935)));
    layer3_outputs(5879) <= (layer2_outputs(3699)) and not (layer2_outputs(444));
    layer3_outputs(5880) <= (layer2_outputs(7013)) or (layer2_outputs(4939));
    layer3_outputs(5881) <= not(layer2_outputs(10135));
    layer3_outputs(5882) <= layer2_outputs(4432);
    layer3_outputs(5883) <= not((layer2_outputs(1189)) xor (layer2_outputs(4218)));
    layer3_outputs(5884) <= (layer2_outputs(605)) xor (layer2_outputs(2181));
    layer3_outputs(5885) <= (layer2_outputs(8182)) and (layer2_outputs(972));
    layer3_outputs(5886) <= not(layer2_outputs(466));
    layer3_outputs(5887) <= layer2_outputs(2453);
    layer3_outputs(5888) <= layer2_outputs(2019);
    layer3_outputs(5889) <= (layer2_outputs(9920)) and not (layer2_outputs(8844));
    layer3_outputs(5890) <= not(layer2_outputs(9838));
    layer3_outputs(5891) <= not(layer2_outputs(414));
    layer3_outputs(5892) <= '1';
    layer3_outputs(5893) <= layer2_outputs(8919);
    layer3_outputs(5894) <= not(layer2_outputs(9098));
    layer3_outputs(5895) <= not(layer2_outputs(1285));
    layer3_outputs(5896) <= layer2_outputs(6429);
    layer3_outputs(5897) <= not(layer2_outputs(1720));
    layer3_outputs(5898) <= layer2_outputs(6118);
    layer3_outputs(5899) <= (layer2_outputs(9751)) or (layer2_outputs(2515));
    layer3_outputs(5900) <= '1';
    layer3_outputs(5901) <= not((layer2_outputs(9806)) xor (layer2_outputs(8217)));
    layer3_outputs(5902) <= (layer2_outputs(5914)) and not (layer2_outputs(3330));
    layer3_outputs(5903) <= (layer2_outputs(497)) and not (layer2_outputs(7625));
    layer3_outputs(5904) <= not((layer2_outputs(6203)) xor (layer2_outputs(4812)));
    layer3_outputs(5905) <= not(layer2_outputs(5147));
    layer3_outputs(5906) <= not((layer2_outputs(8838)) or (layer2_outputs(2695)));
    layer3_outputs(5907) <= not(layer2_outputs(9561));
    layer3_outputs(5908) <= (layer2_outputs(8006)) or (layer2_outputs(10119));
    layer3_outputs(5909) <= not((layer2_outputs(3954)) and (layer2_outputs(8392)));
    layer3_outputs(5910) <= layer2_outputs(5944);
    layer3_outputs(5911) <= not(layer2_outputs(419)) or (layer2_outputs(8042));
    layer3_outputs(5912) <= not((layer2_outputs(1369)) xor (layer2_outputs(3002)));
    layer3_outputs(5913) <= layer2_outputs(5675);
    layer3_outputs(5914) <= (layer2_outputs(9478)) or (layer2_outputs(3338));
    layer3_outputs(5915) <= layer2_outputs(1087);
    layer3_outputs(5916) <= (layer2_outputs(3585)) or (layer2_outputs(4221));
    layer3_outputs(5917) <= layer2_outputs(2130);
    layer3_outputs(5918) <= not((layer2_outputs(8379)) xor (layer2_outputs(3892)));
    layer3_outputs(5919) <= not(layer2_outputs(2645));
    layer3_outputs(5920) <= not(layer2_outputs(9767));
    layer3_outputs(5921) <= '1';
    layer3_outputs(5922) <= layer2_outputs(3038);
    layer3_outputs(5923) <= layer2_outputs(4951);
    layer3_outputs(5924) <= not((layer2_outputs(3006)) xor (layer2_outputs(2255)));
    layer3_outputs(5925) <= (layer2_outputs(964)) and not (layer2_outputs(1034));
    layer3_outputs(5926) <= not(layer2_outputs(3151)) or (layer2_outputs(2639));
    layer3_outputs(5927) <= not(layer2_outputs(5376));
    layer3_outputs(5928) <= not((layer2_outputs(5690)) xor (layer2_outputs(4578)));
    layer3_outputs(5929) <= (layer2_outputs(4728)) or (layer2_outputs(5137));
    layer3_outputs(5930) <= not(layer2_outputs(2224)) or (layer2_outputs(6150));
    layer3_outputs(5931) <= not((layer2_outputs(6806)) or (layer2_outputs(1215)));
    layer3_outputs(5932) <= not(layer2_outputs(319));
    layer3_outputs(5933) <= not((layer2_outputs(3925)) xor (layer2_outputs(2914)));
    layer3_outputs(5934) <= not((layer2_outputs(858)) or (layer2_outputs(6845)));
    layer3_outputs(5935) <= not(layer2_outputs(930));
    layer3_outputs(5936) <= not((layer2_outputs(4582)) and (layer2_outputs(8208)));
    layer3_outputs(5937) <= not((layer2_outputs(4416)) xor (layer2_outputs(1866)));
    layer3_outputs(5938) <= not((layer2_outputs(2580)) xor (layer2_outputs(6941)));
    layer3_outputs(5939) <= (layer2_outputs(6224)) and (layer2_outputs(1509));
    layer3_outputs(5940) <= not(layer2_outputs(10189));
    layer3_outputs(5941) <= (layer2_outputs(6606)) or (layer2_outputs(2021));
    layer3_outputs(5942) <= (layer2_outputs(3670)) xor (layer2_outputs(5069));
    layer3_outputs(5943) <= not((layer2_outputs(2030)) and (layer2_outputs(295)));
    layer3_outputs(5944) <= not(layer2_outputs(193));
    layer3_outputs(5945) <= not(layer2_outputs(7676));
    layer3_outputs(5946) <= (layer2_outputs(9106)) or (layer2_outputs(8175));
    layer3_outputs(5947) <= not(layer2_outputs(4224));
    layer3_outputs(5948) <= (layer2_outputs(1832)) or (layer2_outputs(6718));
    layer3_outputs(5949) <= not(layer2_outputs(5428));
    layer3_outputs(5950) <= not(layer2_outputs(2020));
    layer3_outputs(5951) <= layer2_outputs(8341);
    layer3_outputs(5952) <= not(layer2_outputs(9975));
    layer3_outputs(5953) <= (layer2_outputs(5773)) or (layer2_outputs(5157));
    layer3_outputs(5954) <= not(layer2_outputs(7939)) or (layer2_outputs(1423));
    layer3_outputs(5955) <= not(layer2_outputs(8000));
    layer3_outputs(5956) <= (layer2_outputs(1405)) or (layer2_outputs(4137));
    layer3_outputs(5957) <= not((layer2_outputs(312)) xor (layer2_outputs(6565)));
    layer3_outputs(5958) <= not(layer2_outputs(7083));
    layer3_outputs(5959) <= layer2_outputs(6612);
    layer3_outputs(5960) <= not(layer2_outputs(1727)) or (layer2_outputs(7285));
    layer3_outputs(5961) <= (layer2_outputs(10218)) xor (layer2_outputs(4913));
    layer3_outputs(5962) <= (layer2_outputs(2483)) or (layer2_outputs(2534));
    layer3_outputs(5963) <= not((layer2_outputs(4321)) and (layer2_outputs(2686)));
    layer3_outputs(5964) <= not((layer2_outputs(5251)) and (layer2_outputs(1445)));
    layer3_outputs(5965) <= not((layer2_outputs(9821)) xor (layer2_outputs(6348)));
    layer3_outputs(5966) <= not(layer2_outputs(4113));
    layer3_outputs(5967) <= not(layer2_outputs(3295));
    layer3_outputs(5968) <= not(layer2_outputs(2370));
    layer3_outputs(5969) <= not(layer2_outputs(9809)) or (layer2_outputs(2106));
    layer3_outputs(5970) <= layer2_outputs(7692);
    layer3_outputs(5971) <= (layer2_outputs(2584)) and not (layer2_outputs(8592));
    layer3_outputs(5972) <= (layer2_outputs(4946)) and not (layer2_outputs(9637));
    layer3_outputs(5973) <= not((layer2_outputs(1021)) and (layer2_outputs(5152)));
    layer3_outputs(5974) <= (layer2_outputs(2806)) xor (layer2_outputs(1422));
    layer3_outputs(5975) <= layer2_outputs(8537);
    layer3_outputs(5976) <= (layer2_outputs(664)) or (layer2_outputs(7475));
    layer3_outputs(5977) <= (layer2_outputs(6288)) and not (layer2_outputs(2317));
    layer3_outputs(5978) <= not(layer2_outputs(2653));
    layer3_outputs(5979) <= not((layer2_outputs(6361)) or (layer2_outputs(399)));
    layer3_outputs(5980) <= (layer2_outputs(2110)) and not (layer2_outputs(2144));
    layer3_outputs(5981) <= (layer2_outputs(3873)) and not (layer2_outputs(3897));
    layer3_outputs(5982) <= (layer2_outputs(8117)) and (layer2_outputs(6518));
    layer3_outputs(5983) <= layer2_outputs(7142);
    layer3_outputs(5984) <= not(layer2_outputs(8892)) or (layer2_outputs(4500));
    layer3_outputs(5985) <= (layer2_outputs(387)) and (layer2_outputs(8945));
    layer3_outputs(5986) <= (layer2_outputs(7703)) and not (layer2_outputs(2114));
    layer3_outputs(5987) <= not((layer2_outputs(3830)) and (layer2_outputs(3839)));
    layer3_outputs(5988) <= not(layer2_outputs(4777));
    layer3_outputs(5989) <= not(layer2_outputs(4178)) or (layer2_outputs(9895));
    layer3_outputs(5990) <= (layer2_outputs(80)) xor (layer2_outputs(5106));
    layer3_outputs(5991) <= not(layer2_outputs(5871));
    layer3_outputs(5992) <= not(layer2_outputs(2754));
    layer3_outputs(5993) <= not(layer2_outputs(8355));
    layer3_outputs(5994) <= not(layer2_outputs(2128));
    layer3_outputs(5995) <= not(layer2_outputs(9202));
    layer3_outputs(5996) <= not(layer2_outputs(8400));
    layer3_outputs(5997) <= not(layer2_outputs(8478));
    layer3_outputs(5998) <= (layer2_outputs(7633)) and (layer2_outputs(4717));
    layer3_outputs(5999) <= layer2_outputs(6516);
    layer3_outputs(6000) <= not(layer2_outputs(9305));
    layer3_outputs(6001) <= layer2_outputs(4904);
    layer3_outputs(6002) <= layer2_outputs(1318);
    layer3_outputs(6003) <= (layer2_outputs(6758)) or (layer2_outputs(7880));
    layer3_outputs(6004) <= not(layer2_outputs(6549));
    layer3_outputs(6005) <= not(layer2_outputs(623)) or (layer2_outputs(8880));
    layer3_outputs(6006) <= (layer2_outputs(2240)) and not (layer2_outputs(6284));
    layer3_outputs(6007) <= layer2_outputs(2335);
    layer3_outputs(6008) <= not((layer2_outputs(3233)) and (layer2_outputs(7892)));
    layer3_outputs(6009) <= not((layer2_outputs(3725)) or (layer2_outputs(4967)));
    layer3_outputs(6010) <= layer2_outputs(8546);
    layer3_outputs(6011) <= not((layer2_outputs(6103)) or (layer2_outputs(6557)));
    layer3_outputs(6012) <= layer2_outputs(7141);
    layer3_outputs(6013) <= layer2_outputs(1891);
    layer3_outputs(6014) <= not(layer2_outputs(9898)) or (layer2_outputs(9374));
    layer3_outputs(6015) <= (layer2_outputs(1016)) xor (layer2_outputs(5499));
    layer3_outputs(6016) <= layer2_outputs(9865);
    layer3_outputs(6017) <= not(layer2_outputs(8740)) or (layer2_outputs(7496));
    layer3_outputs(6018) <= not((layer2_outputs(2259)) and (layer2_outputs(8224)));
    layer3_outputs(6019) <= layer2_outputs(9654);
    layer3_outputs(6020) <= not((layer2_outputs(1943)) xor (layer2_outputs(7566)));
    layer3_outputs(6021) <= layer2_outputs(3963);
    layer3_outputs(6022) <= not(layer2_outputs(2679));
    layer3_outputs(6023) <= (layer2_outputs(6304)) xor (layer2_outputs(2839));
    layer3_outputs(6024) <= not(layer2_outputs(5211));
    layer3_outputs(6025) <= not(layer2_outputs(2641));
    layer3_outputs(6026) <= not(layer2_outputs(8837)) or (layer2_outputs(786));
    layer3_outputs(6027) <= layer2_outputs(8624);
    layer3_outputs(6028) <= not(layer2_outputs(7514));
    layer3_outputs(6029) <= not((layer2_outputs(5442)) or (layer2_outputs(6252)));
    layer3_outputs(6030) <= layer2_outputs(2728);
    layer3_outputs(6031) <= not(layer2_outputs(4713));
    layer3_outputs(6032) <= (layer2_outputs(8539)) or (layer2_outputs(54));
    layer3_outputs(6033) <= (layer2_outputs(2011)) and not (layer2_outputs(1340));
    layer3_outputs(6034) <= not(layer2_outputs(9527));
    layer3_outputs(6035) <= not(layer2_outputs(8427)) or (layer2_outputs(64));
    layer3_outputs(6036) <= not(layer2_outputs(7157)) or (layer2_outputs(5463));
    layer3_outputs(6037) <= not(layer2_outputs(4871));
    layer3_outputs(6038) <= layer2_outputs(6216);
    layer3_outputs(6039) <= not((layer2_outputs(9857)) and (layer2_outputs(6379)));
    layer3_outputs(6040) <= not((layer2_outputs(1736)) or (layer2_outputs(5588)));
    layer3_outputs(6041) <= not(layer2_outputs(3033));
    layer3_outputs(6042) <= not(layer2_outputs(9919));
    layer3_outputs(6043) <= not(layer2_outputs(730)) or (layer2_outputs(7288));
    layer3_outputs(6044) <= layer2_outputs(7552);
    layer3_outputs(6045) <= layer2_outputs(151);
    layer3_outputs(6046) <= not(layer2_outputs(2818));
    layer3_outputs(6047) <= (layer2_outputs(7102)) and (layer2_outputs(1726));
    layer3_outputs(6048) <= not((layer2_outputs(9362)) or (layer2_outputs(891)));
    layer3_outputs(6049) <= layer2_outputs(1762);
    layer3_outputs(6050) <= (layer2_outputs(7437)) or (layer2_outputs(4652));
    layer3_outputs(6051) <= (layer2_outputs(5269)) and not (layer2_outputs(5095));
    layer3_outputs(6052) <= not(layer2_outputs(2649));
    layer3_outputs(6053) <= layer2_outputs(9670);
    layer3_outputs(6054) <= not(layer2_outputs(8081));
    layer3_outputs(6055) <= not(layer2_outputs(2937));
    layer3_outputs(6056) <= not((layer2_outputs(367)) and (layer2_outputs(4196)));
    layer3_outputs(6057) <= not(layer2_outputs(8044));
    layer3_outputs(6058) <= layer2_outputs(5748);
    layer3_outputs(6059) <= not(layer2_outputs(4042));
    layer3_outputs(6060) <= not(layer2_outputs(4139));
    layer3_outputs(6061) <= not(layer2_outputs(9356)) or (layer2_outputs(9383));
    layer3_outputs(6062) <= not(layer2_outputs(5167));
    layer3_outputs(6063) <= layer2_outputs(2629);
    layer3_outputs(6064) <= layer2_outputs(8750);
    layer3_outputs(6065) <= not(layer2_outputs(6826));
    layer3_outputs(6066) <= not(layer2_outputs(5619));
    layer3_outputs(6067) <= not(layer2_outputs(7594)) or (layer2_outputs(3167));
    layer3_outputs(6068) <= not(layer2_outputs(10187));
    layer3_outputs(6069) <= not((layer2_outputs(2717)) and (layer2_outputs(7749)));
    layer3_outputs(6070) <= layer2_outputs(8312);
    layer3_outputs(6071) <= not(layer2_outputs(5743));
    layer3_outputs(6072) <= not(layer2_outputs(9453));
    layer3_outputs(6073) <= layer2_outputs(4082);
    layer3_outputs(6074) <= (layer2_outputs(1193)) and not (layer2_outputs(10092));
    layer3_outputs(6075) <= (layer2_outputs(1195)) or (layer2_outputs(2825));
    layer3_outputs(6076) <= not(layer2_outputs(6972)) or (layer2_outputs(8952));
    layer3_outputs(6077) <= layer2_outputs(3797);
    layer3_outputs(6078) <= not(layer2_outputs(2938));
    layer3_outputs(6079) <= not((layer2_outputs(3432)) or (layer2_outputs(1389)));
    layer3_outputs(6080) <= (layer2_outputs(3546)) and not (layer2_outputs(948));
    layer3_outputs(6081) <= not(layer2_outputs(9138)) or (layer2_outputs(1895));
    layer3_outputs(6082) <= '0';
    layer3_outputs(6083) <= (layer2_outputs(9281)) xor (layer2_outputs(8200));
    layer3_outputs(6084) <= layer2_outputs(1720);
    layer3_outputs(6085) <= not(layer2_outputs(7740));
    layer3_outputs(6086) <= (layer2_outputs(6360)) xor (layer2_outputs(240));
    layer3_outputs(6087) <= '1';
    layer3_outputs(6088) <= not((layer2_outputs(4345)) and (layer2_outputs(1623)));
    layer3_outputs(6089) <= not((layer2_outputs(2546)) xor (layer2_outputs(1622)));
    layer3_outputs(6090) <= (layer2_outputs(5981)) or (layer2_outputs(4674));
    layer3_outputs(6091) <= (layer2_outputs(9924)) xor (layer2_outputs(9494));
    layer3_outputs(6092) <= layer2_outputs(6755);
    layer3_outputs(6093) <= not(layer2_outputs(9731));
    layer3_outputs(6094) <= not(layer2_outputs(2615));
    layer3_outputs(6095) <= layer2_outputs(1800);
    layer3_outputs(6096) <= (layer2_outputs(3227)) and (layer2_outputs(3133));
    layer3_outputs(6097) <= not((layer2_outputs(605)) or (layer2_outputs(8179)));
    layer3_outputs(6098) <= layer2_outputs(7900);
    layer3_outputs(6099) <= (layer2_outputs(7150)) xor (layer2_outputs(5151));
    layer3_outputs(6100) <= (layer2_outputs(329)) xor (layer2_outputs(9165));
    layer3_outputs(6101) <= (layer2_outputs(3071)) or (layer2_outputs(2904));
    layer3_outputs(6102) <= layer2_outputs(3552);
    layer3_outputs(6103) <= not(layer2_outputs(3818)) or (layer2_outputs(4374));
    layer3_outputs(6104) <= layer2_outputs(2104);
    layer3_outputs(6105) <= not(layer2_outputs(2913));
    layer3_outputs(6106) <= not(layer2_outputs(4153));
    layer3_outputs(6107) <= (layer2_outputs(7310)) and not (layer2_outputs(8902));
    layer3_outputs(6108) <= not((layer2_outputs(7815)) and (layer2_outputs(1362)));
    layer3_outputs(6109) <= not((layer2_outputs(2278)) xor (layer2_outputs(1601)));
    layer3_outputs(6110) <= not(layer2_outputs(5597));
    layer3_outputs(6111) <= (layer2_outputs(9502)) xor (layer2_outputs(9328));
    layer3_outputs(6112) <= not(layer2_outputs(3336));
    layer3_outputs(6113) <= '1';
    layer3_outputs(6114) <= layer2_outputs(4405);
    layer3_outputs(6115) <= layer2_outputs(7700);
    layer3_outputs(6116) <= not(layer2_outputs(219));
    layer3_outputs(6117) <= (layer2_outputs(8279)) and (layer2_outputs(5681));
    layer3_outputs(6118) <= not(layer2_outputs(7093));
    layer3_outputs(6119) <= (layer2_outputs(7569)) xor (layer2_outputs(5105));
    layer3_outputs(6120) <= '0';
    layer3_outputs(6121) <= not(layer2_outputs(840)) or (layer2_outputs(4441));
    layer3_outputs(6122) <= layer2_outputs(75);
    layer3_outputs(6123) <= layer2_outputs(2097);
    layer3_outputs(6124) <= not(layer2_outputs(1787));
    layer3_outputs(6125) <= not(layer2_outputs(626)) or (layer2_outputs(180));
    layer3_outputs(6126) <= (layer2_outputs(7786)) or (layer2_outputs(679));
    layer3_outputs(6127) <= (layer2_outputs(9323)) and (layer2_outputs(5018));
    layer3_outputs(6128) <= layer2_outputs(8452);
    layer3_outputs(6129) <= not(layer2_outputs(4423)) or (layer2_outputs(228));
    layer3_outputs(6130) <= (layer2_outputs(4470)) or (layer2_outputs(1541));
    layer3_outputs(6131) <= layer2_outputs(9207);
    layer3_outputs(6132) <= (layer2_outputs(2524)) or (layer2_outputs(7971));
    layer3_outputs(6133) <= not(layer2_outputs(413));
    layer3_outputs(6134) <= (layer2_outputs(9569)) or (layer2_outputs(636));
    layer3_outputs(6135) <= layer2_outputs(5589);
    layer3_outputs(6136) <= not((layer2_outputs(7432)) or (layer2_outputs(3844)));
    layer3_outputs(6137) <= not((layer2_outputs(5149)) or (layer2_outputs(1461)));
    layer3_outputs(6138) <= not((layer2_outputs(4282)) and (layer2_outputs(2215)));
    layer3_outputs(6139) <= layer2_outputs(4441);
    layer3_outputs(6140) <= not(layer2_outputs(7712)) or (layer2_outputs(7946));
    layer3_outputs(6141) <= layer2_outputs(8998);
    layer3_outputs(6142) <= layer2_outputs(1625);
    layer3_outputs(6143) <= not(layer2_outputs(5004)) or (layer2_outputs(632));
    layer3_outputs(6144) <= not((layer2_outputs(8272)) xor (layer2_outputs(6647)));
    layer3_outputs(6145) <= layer2_outputs(2473);
    layer3_outputs(6146) <= not(layer2_outputs(8938));
    layer3_outputs(6147) <= not(layer2_outputs(10123));
    layer3_outputs(6148) <= not((layer2_outputs(3120)) and (layer2_outputs(680)));
    layer3_outputs(6149) <= not(layer2_outputs(5932));
    layer3_outputs(6150) <= layer2_outputs(8338);
    layer3_outputs(6151) <= layer2_outputs(10187);
    layer3_outputs(6152) <= not((layer2_outputs(2673)) and (layer2_outputs(5097)));
    layer3_outputs(6153) <= not(layer2_outputs(5764)) or (layer2_outputs(5766));
    layer3_outputs(6154) <= layer2_outputs(10013);
    layer3_outputs(6155) <= not(layer2_outputs(6544));
    layer3_outputs(6156) <= not(layer2_outputs(8093));
    layer3_outputs(6157) <= (layer2_outputs(5323)) xor (layer2_outputs(3383));
    layer3_outputs(6158) <= not(layer2_outputs(3563));
    layer3_outputs(6159) <= (layer2_outputs(6879)) and not (layer2_outputs(6308));
    layer3_outputs(6160) <= layer2_outputs(2057);
    layer3_outputs(6161) <= layer2_outputs(4476);
    layer3_outputs(6162) <= (layer2_outputs(7289)) and not (layer2_outputs(245));
    layer3_outputs(6163) <= not((layer2_outputs(3221)) xor (layer2_outputs(9258)));
    layer3_outputs(6164) <= (layer2_outputs(3)) xor (layer2_outputs(1840));
    layer3_outputs(6165) <= not((layer2_outputs(3280)) xor (layer2_outputs(5525)));
    layer3_outputs(6166) <= not((layer2_outputs(9947)) or (layer2_outputs(3242)));
    layer3_outputs(6167) <= (layer2_outputs(8049)) xor (layer2_outputs(5960));
    layer3_outputs(6168) <= not(layer2_outputs(1452));
    layer3_outputs(6169) <= (layer2_outputs(7111)) and not (layer2_outputs(1901));
    layer3_outputs(6170) <= (layer2_outputs(1301)) and not (layer2_outputs(3939));
    layer3_outputs(6171) <= layer2_outputs(4187);
    layer3_outputs(6172) <= (layer2_outputs(1697)) or (layer2_outputs(9461));
    layer3_outputs(6173) <= not(layer2_outputs(6425));
    layer3_outputs(6174) <= (layer2_outputs(1182)) xor (layer2_outputs(3154));
    layer3_outputs(6175) <= not((layer2_outputs(9317)) xor (layer2_outputs(5274)));
    layer3_outputs(6176) <= (layer2_outputs(6368)) and not (layer2_outputs(7407));
    layer3_outputs(6177) <= '1';
    layer3_outputs(6178) <= (layer2_outputs(7933)) and not (layer2_outputs(1273));
    layer3_outputs(6179) <= not(layer2_outputs(8157));
    layer3_outputs(6180) <= layer2_outputs(8695);
    layer3_outputs(6181) <= layer2_outputs(3736);
    layer3_outputs(6182) <= (layer2_outputs(1102)) and not (layer2_outputs(3476));
    layer3_outputs(6183) <= not((layer2_outputs(9762)) or (layer2_outputs(7271)));
    layer3_outputs(6184) <= not(layer2_outputs(3450)) or (layer2_outputs(8880));
    layer3_outputs(6185) <= not(layer2_outputs(1337));
    layer3_outputs(6186) <= not(layer2_outputs(10034));
    layer3_outputs(6187) <= (layer2_outputs(9331)) and (layer2_outputs(859));
    layer3_outputs(6188) <= (layer2_outputs(506)) and not (layer2_outputs(3358));
    layer3_outputs(6189) <= not(layer2_outputs(8026));
    layer3_outputs(6190) <= not(layer2_outputs(4965));
    layer3_outputs(6191) <= not(layer2_outputs(6961)) or (layer2_outputs(5828));
    layer3_outputs(6192) <= layer2_outputs(5300);
    layer3_outputs(6193) <= layer2_outputs(3561);
    layer3_outputs(6194) <= '0';
    layer3_outputs(6195) <= (layer2_outputs(1583)) and not (layer2_outputs(8432));
    layer3_outputs(6196) <= layer2_outputs(3906);
    layer3_outputs(6197) <= layer2_outputs(4130);
    layer3_outputs(6198) <= not((layer2_outputs(248)) and (layer2_outputs(1648)));
    layer3_outputs(6199) <= not(layer2_outputs(5743));
    layer3_outputs(6200) <= layer2_outputs(5784);
    layer3_outputs(6201) <= not(layer2_outputs(4746));
    layer3_outputs(6202) <= not((layer2_outputs(5441)) xor (layer2_outputs(703)));
    layer3_outputs(6203) <= not(layer2_outputs(10016));
    layer3_outputs(6204) <= layer2_outputs(8422);
    layer3_outputs(6205) <= layer2_outputs(3139);
    layer3_outputs(6206) <= layer2_outputs(9519);
    layer3_outputs(6207) <= layer2_outputs(6445);
    layer3_outputs(6208) <= not((layer2_outputs(8848)) or (layer2_outputs(8290)));
    layer3_outputs(6209) <= (layer2_outputs(9067)) and not (layer2_outputs(5539));
    layer3_outputs(6210) <= not(layer2_outputs(929));
    layer3_outputs(6211) <= not(layer2_outputs(1079));
    layer3_outputs(6212) <= not(layer2_outputs(4609));
    layer3_outputs(6213) <= not(layer2_outputs(7861)) or (layer2_outputs(3325));
    layer3_outputs(6214) <= (layer2_outputs(8759)) and not (layer2_outputs(1001));
    layer3_outputs(6215) <= not(layer2_outputs(2742)) or (layer2_outputs(4644));
    layer3_outputs(6216) <= layer2_outputs(8988);
    layer3_outputs(6217) <= layer2_outputs(2391);
    layer3_outputs(6218) <= not(layer2_outputs(1443));
    layer3_outputs(6219) <= layer2_outputs(3779);
    layer3_outputs(6220) <= (layer2_outputs(9493)) and not (layer2_outputs(1099));
    layer3_outputs(6221) <= (layer2_outputs(9349)) and not (layer2_outputs(5502));
    layer3_outputs(6222) <= (layer2_outputs(2634)) or (layer2_outputs(3098));
    layer3_outputs(6223) <= (layer2_outputs(6119)) xor (layer2_outputs(4255));
    layer3_outputs(6224) <= not(layer2_outputs(1084)) or (layer2_outputs(5917));
    layer3_outputs(6225) <= (layer2_outputs(5682)) and (layer2_outputs(8416));
    layer3_outputs(6226) <= not(layer2_outputs(4241));
    layer3_outputs(6227) <= layer2_outputs(10239);
    layer3_outputs(6228) <= layer2_outputs(2387);
    layer3_outputs(6229) <= layer2_outputs(7696);
    layer3_outputs(6230) <= (layer2_outputs(2669)) and not (layer2_outputs(7853));
    layer3_outputs(6231) <= (layer2_outputs(7072)) or (layer2_outputs(5927));
    layer3_outputs(6232) <= '1';
    layer3_outputs(6233) <= not((layer2_outputs(1991)) xor (layer2_outputs(8417)));
    layer3_outputs(6234) <= (layer2_outputs(3224)) and (layer2_outputs(3146));
    layer3_outputs(6235) <= layer2_outputs(9119);
    layer3_outputs(6236) <= (layer2_outputs(9083)) and not (layer2_outputs(3539));
    layer3_outputs(6237) <= (layer2_outputs(8828)) or (layer2_outputs(8419));
    layer3_outputs(6238) <= (layer2_outputs(6648)) and not (layer2_outputs(7526));
    layer3_outputs(6239) <= (layer2_outputs(4131)) xor (layer2_outputs(8292));
    layer3_outputs(6240) <= not(layer2_outputs(5871));
    layer3_outputs(6241) <= layer2_outputs(5745);
    layer3_outputs(6242) <= layer2_outputs(10117);
    layer3_outputs(6243) <= not(layer2_outputs(2283)) or (layer2_outputs(2430));
    layer3_outputs(6244) <= not(layer2_outputs(10101)) or (layer2_outputs(10005));
    layer3_outputs(6245) <= '0';
    layer3_outputs(6246) <= layer2_outputs(6799);
    layer3_outputs(6247) <= not((layer2_outputs(5359)) xor (layer2_outputs(716)));
    layer3_outputs(6248) <= (layer2_outputs(3662)) or (layer2_outputs(9871));
    layer3_outputs(6249) <= layer2_outputs(7651);
    layer3_outputs(6250) <= not(layer2_outputs(7334));
    layer3_outputs(6251) <= not(layer2_outputs(5543));
    layer3_outputs(6252) <= layer2_outputs(139);
    layer3_outputs(6253) <= not(layer2_outputs(6454));
    layer3_outputs(6254) <= (layer2_outputs(9506)) and not (layer2_outputs(8533));
    layer3_outputs(6255) <= not(layer2_outputs(509));
    layer3_outputs(6256) <= not(layer2_outputs(7163)) or (layer2_outputs(8037));
    layer3_outputs(6257) <= not((layer2_outputs(8372)) or (layer2_outputs(8876)));
    layer3_outputs(6258) <= (layer2_outputs(7024)) and not (layer2_outputs(2759));
    layer3_outputs(6259) <= layer2_outputs(9572);
    layer3_outputs(6260) <= layer2_outputs(630);
    layer3_outputs(6261) <= not((layer2_outputs(5670)) xor (layer2_outputs(6573)));
    layer3_outputs(6262) <= not((layer2_outputs(5168)) xor (layer2_outputs(9440)));
    layer3_outputs(6263) <= not((layer2_outputs(369)) and (layer2_outputs(181)));
    layer3_outputs(6264) <= (layer2_outputs(4206)) and not (layer2_outputs(1378));
    layer3_outputs(6265) <= (layer2_outputs(1731)) and not (layer2_outputs(8177));
    layer3_outputs(6266) <= layer2_outputs(9608);
    layer3_outputs(6267) <= layer2_outputs(7868);
    layer3_outputs(6268) <= not(layer2_outputs(6656)) or (layer2_outputs(8882));
    layer3_outputs(6269) <= not((layer2_outputs(8140)) or (layer2_outputs(7229)));
    layer3_outputs(6270) <= layer2_outputs(6947);
    layer3_outputs(6271) <= '0';
    layer3_outputs(6272) <= not(layer2_outputs(7418)) or (layer2_outputs(7947));
    layer3_outputs(6273) <= not((layer2_outputs(4827)) and (layer2_outputs(4023)));
    layer3_outputs(6274) <= (layer2_outputs(172)) or (layer2_outputs(3683));
    layer3_outputs(6275) <= layer2_outputs(8943);
    layer3_outputs(6276) <= not(layer2_outputs(9278));
    layer3_outputs(6277) <= layer2_outputs(7777);
    layer3_outputs(6278) <= not(layer2_outputs(1728)) or (layer2_outputs(1394));
    layer3_outputs(6279) <= '1';
    layer3_outputs(6280) <= not(layer2_outputs(2458)) or (layer2_outputs(5068));
    layer3_outputs(6281) <= '1';
    layer3_outputs(6282) <= (layer2_outputs(5628)) and not (layer2_outputs(4867));
    layer3_outputs(6283) <= not(layer2_outputs(4388));
    layer3_outputs(6284) <= (layer2_outputs(9498)) and (layer2_outputs(6757));
    layer3_outputs(6285) <= layer2_outputs(1608);
    layer3_outputs(6286) <= layer2_outputs(5493);
    layer3_outputs(6287) <= '1';
    layer3_outputs(6288) <= not(layer2_outputs(7010));
    layer3_outputs(6289) <= layer2_outputs(10125);
    layer3_outputs(6290) <= layer2_outputs(2778);
    layer3_outputs(6291) <= not((layer2_outputs(1045)) or (layer2_outputs(1395)));
    layer3_outputs(6292) <= (layer2_outputs(8484)) or (layer2_outputs(4763));
    layer3_outputs(6293) <= not(layer2_outputs(1113)) or (layer2_outputs(5075));
    layer3_outputs(6294) <= '0';
    layer3_outputs(6295) <= not(layer2_outputs(8196)) or (layer2_outputs(10182));
    layer3_outputs(6296) <= layer2_outputs(6086);
    layer3_outputs(6297) <= not((layer2_outputs(3669)) or (layer2_outputs(7666)));
    layer3_outputs(6298) <= not((layer2_outputs(3150)) xor (layer2_outputs(7505)));
    layer3_outputs(6299) <= layer2_outputs(7419);
    layer3_outputs(6300) <= layer2_outputs(9280);
    layer3_outputs(6301) <= not((layer2_outputs(4286)) and (layer2_outputs(1457)));
    layer3_outputs(6302) <= not((layer2_outputs(1593)) or (layer2_outputs(1798)));
    layer3_outputs(6303) <= not((layer2_outputs(6619)) and (layer2_outputs(560)));
    layer3_outputs(6304) <= (layer2_outputs(4962)) and not (layer2_outputs(3510));
    layer3_outputs(6305) <= (layer2_outputs(9407)) xor (layer2_outputs(8332));
    layer3_outputs(6306) <= layer2_outputs(3709);
    layer3_outputs(6307) <= not(layer2_outputs(8305));
    layer3_outputs(6308) <= (layer2_outputs(5780)) and (layer2_outputs(4750));
    layer3_outputs(6309) <= (layer2_outputs(3461)) and not (layer2_outputs(2932));
    layer3_outputs(6310) <= not(layer2_outputs(5599));
    layer3_outputs(6311) <= not((layer2_outputs(2139)) and (layer2_outputs(7424)));
    layer3_outputs(6312) <= not((layer2_outputs(2544)) and (layer2_outputs(8728)));
    layer3_outputs(6313) <= not(layer2_outputs(5984));
    layer3_outputs(6314) <= layer2_outputs(6633);
    layer3_outputs(6315) <= layer2_outputs(5551);
    layer3_outputs(6316) <= not(layer2_outputs(9148));
    layer3_outputs(6317) <= not(layer2_outputs(10148)) or (layer2_outputs(8687));
    layer3_outputs(6318) <= not(layer2_outputs(5830));
    layer3_outputs(6319) <= not(layer2_outputs(9255));
    layer3_outputs(6320) <= layer2_outputs(449);
    layer3_outputs(6321) <= (layer2_outputs(3571)) or (layer2_outputs(4783));
    layer3_outputs(6322) <= not((layer2_outputs(5429)) xor (layer2_outputs(8475)));
    layer3_outputs(6323) <= (layer2_outputs(2288)) or (layer2_outputs(1919));
    layer3_outputs(6324) <= not(layer2_outputs(9275)) or (layer2_outputs(6167));
    layer3_outputs(6325) <= layer2_outputs(3874);
    layer3_outputs(6326) <= (layer2_outputs(4122)) and not (layer2_outputs(2768));
    layer3_outputs(6327) <= layer2_outputs(6542);
    layer3_outputs(6328) <= not(layer2_outputs(5658));
    layer3_outputs(6329) <= layer2_outputs(228);
    layer3_outputs(6330) <= not(layer2_outputs(10186));
    layer3_outputs(6331) <= layer2_outputs(5489);
    layer3_outputs(6332) <= layer2_outputs(7733);
    layer3_outputs(6333) <= not(layer2_outputs(8569)) or (layer2_outputs(9934));
    layer3_outputs(6334) <= layer2_outputs(2322);
    layer3_outputs(6335) <= not(layer2_outputs(5033)) or (layer2_outputs(148));
    layer3_outputs(6336) <= layer2_outputs(121);
    layer3_outputs(6337) <= (layer2_outputs(6281)) and not (layer2_outputs(5094));
    layer3_outputs(6338) <= not(layer2_outputs(4211));
    layer3_outputs(6339) <= layer2_outputs(9435);
    layer3_outputs(6340) <= (layer2_outputs(870)) and not (layer2_outputs(2843));
    layer3_outputs(6341) <= (layer2_outputs(7296)) and not (layer2_outputs(4486));
    layer3_outputs(6342) <= not(layer2_outputs(2645));
    layer3_outputs(6343) <= not((layer2_outputs(3902)) or (layer2_outputs(3132)));
    layer3_outputs(6344) <= layer2_outputs(4072);
    layer3_outputs(6345) <= (layer2_outputs(7247)) and not (layer2_outputs(7063));
    layer3_outputs(6346) <= not(layer2_outputs(6361));
    layer3_outputs(6347) <= not(layer2_outputs(2677));
    layer3_outputs(6348) <= not((layer2_outputs(4050)) xor (layer2_outputs(5149)));
    layer3_outputs(6349) <= not((layer2_outputs(206)) or (layer2_outputs(7026)));
    layer3_outputs(6350) <= (layer2_outputs(8204)) and not (layer2_outputs(2886));
    layer3_outputs(6351) <= not(layer2_outputs(5933));
    layer3_outputs(6352) <= not(layer2_outputs(4527));
    layer3_outputs(6353) <= layer2_outputs(2958);
    layer3_outputs(6354) <= (layer2_outputs(2314)) and (layer2_outputs(9854));
    layer3_outputs(6355) <= not((layer2_outputs(1541)) xor (layer2_outputs(2595)));
    layer3_outputs(6356) <= not(layer2_outputs(3885)) or (layer2_outputs(1177));
    layer3_outputs(6357) <= '0';
    layer3_outputs(6358) <= not((layer2_outputs(4378)) and (layer2_outputs(4839)));
    layer3_outputs(6359) <= not(layer2_outputs(4878)) or (layer2_outputs(4310));
    layer3_outputs(6360) <= not(layer2_outputs(1119)) or (layer2_outputs(4709));
    layer3_outputs(6361) <= layer2_outputs(4160);
    layer3_outputs(6362) <= (layer2_outputs(7818)) xor (layer2_outputs(7657));
    layer3_outputs(6363) <= not(layer2_outputs(8444)) or (layer2_outputs(9735));
    layer3_outputs(6364) <= not(layer2_outputs(9447));
    layer3_outputs(6365) <= (layer2_outputs(2372)) and (layer2_outputs(9920));
    layer3_outputs(6366) <= layer2_outputs(3397);
    layer3_outputs(6367) <= not(layer2_outputs(6278));
    layer3_outputs(6368) <= not((layer2_outputs(977)) xor (layer2_outputs(9261)));
    layer3_outputs(6369) <= layer2_outputs(4557);
    layer3_outputs(6370) <= not(layer2_outputs(7558));
    layer3_outputs(6371) <= layer2_outputs(2760);
    layer3_outputs(6372) <= not(layer2_outputs(6645));
    layer3_outputs(6373) <= not(layer2_outputs(1162));
    layer3_outputs(6374) <= (layer2_outputs(6064)) xor (layer2_outputs(2306));
    layer3_outputs(6375) <= not(layer2_outputs(3041));
    layer3_outputs(6376) <= layer2_outputs(4596);
    layer3_outputs(6377) <= not(layer2_outputs(3772)) or (layer2_outputs(1344));
    layer3_outputs(6378) <= layer2_outputs(615);
    layer3_outputs(6379) <= not((layer2_outputs(973)) xor (layer2_outputs(2088)));
    layer3_outputs(6380) <= (layer2_outputs(821)) xor (layer2_outputs(2193));
    layer3_outputs(6381) <= not(layer2_outputs(4064));
    layer3_outputs(6382) <= not(layer2_outputs(3077));
    layer3_outputs(6383) <= (layer2_outputs(334)) xor (layer2_outputs(1096));
    layer3_outputs(6384) <= layer2_outputs(7399);
    layer3_outputs(6385) <= not(layer2_outputs(1131));
    layer3_outputs(6386) <= layer2_outputs(4483);
    layer3_outputs(6387) <= not(layer2_outputs(132));
    layer3_outputs(6388) <= '0';
    layer3_outputs(6389) <= not(layer2_outputs(7213));
    layer3_outputs(6390) <= not((layer2_outputs(7314)) xor (layer2_outputs(8404)));
    layer3_outputs(6391) <= layer2_outputs(5513);
    layer3_outputs(6392) <= not((layer2_outputs(204)) or (layer2_outputs(1680)));
    layer3_outputs(6393) <= not((layer2_outputs(8360)) or (layer2_outputs(3480)));
    layer3_outputs(6394) <= not(layer2_outputs(6888));
    layer3_outputs(6395) <= (layer2_outputs(2695)) or (layer2_outputs(5992));
    layer3_outputs(6396) <= layer2_outputs(1506);
    layer3_outputs(6397) <= not((layer2_outputs(5283)) or (layer2_outputs(8509)));
    layer3_outputs(6398) <= (layer2_outputs(8014)) or (layer2_outputs(4436));
    layer3_outputs(6399) <= (layer2_outputs(2783)) or (layer2_outputs(8300));
    layer3_outputs(6400) <= layer2_outputs(5253);
    layer3_outputs(6401) <= not(layer2_outputs(8346)) or (layer2_outputs(8438));
    layer3_outputs(6402) <= layer2_outputs(7881);
    layer3_outputs(6403) <= (layer2_outputs(7449)) and (layer2_outputs(9480));
    layer3_outputs(6404) <= layer2_outputs(5245);
    layer3_outputs(6405) <= not(layer2_outputs(6639));
    layer3_outputs(6406) <= '0';
    layer3_outputs(6407) <= (layer2_outputs(5123)) and (layer2_outputs(1688));
    layer3_outputs(6408) <= (layer2_outputs(3122)) and not (layer2_outputs(7376));
    layer3_outputs(6409) <= not(layer2_outputs(2732));
    layer3_outputs(6410) <= not(layer2_outputs(3467)) or (layer2_outputs(2301));
    layer3_outputs(6411) <= (layer2_outputs(9218)) or (layer2_outputs(6118));
    layer3_outputs(6412) <= (layer2_outputs(418)) or (layer2_outputs(1159));
    layer3_outputs(6413) <= layer2_outputs(10127);
    layer3_outputs(6414) <= not(layer2_outputs(9245)) or (layer2_outputs(6393));
    layer3_outputs(6415) <= not(layer2_outputs(9830)) or (layer2_outputs(7385));
    layer3_outputs(6416) <= not(layer2_outputs(4521));
    layer3_outputs(6417) <= layer2_outputs(5401);
    layer3_outputs(6418) <= (layer2_outputs(4662)) or (layer2_outputs(6074));
    layer3_outputs(6419) <= (layer2_outputs(2498)) and not (layer2_outputs(1134));
    layer3_outputs(6420) <= layer2_outputs(6528);
    layer3_outputs(6421) <= layer2_outputs(6805);
    layer3_outputs(6422) <= (layer2_outputs(739)) or (layer2_outputs(9050));
    layer3_outputs(6423) <= not((layer2_outputs(5254)) or (layer2_outputs(9108)));
    layer3_outputs(6424) <= not(layer2_outputs(2667));
    layer3_outputs(6425) <= not(layer2_outputs(6891));
    layer3_outputs(6426) <= (layer2_outputs(9233)) and not (layer2_outputs(8477));
    layer3_outputs(6427) <= (layer2_outputs(9360)) xor (layer2_outputs(9853));
    layer3_outputs(6428) <= layer2_outputs(384);
    layer3_outputs(6429) <= not(layer2_outputs(5640)) or (layer2_outputs(1138));
    layer3_outputs(6430) <= not(layer2_outputs(5578));
    layer3_outputs(6431) <= layer2_outputs(9659);
    layer3_outputs(6432) <= '0';
    layer3_outputs(6433) <= (layer2_outputs(432)) and (layer2_outputs(3545));
    layer3_outputs(6434) <= not((layer2_outputs(1076)) xor (layer2_outputs(3669)));
    layer3_outputs(6435) <= (layer2_outputs(963)) and not (layer2_outputs(8532));
    layer3_outputs(6436) <= '1';
    layer3_outputs(6437) <= (layer2_outputs(1917)) and not (layer2_outputs(6135));
    layer3_outputs(6438) <= not(layer2_outputs(8129));
    layer3_outputs(6439) <= layer2_outputs(5903);
    layer3_outputs(6440) <= not(layer2_outputs(2809));
    layer3_outputs(6441) <= not(layer2_outputs(6329));
    layer3_outputs(6442) <= '0';
    layer3_outputs(6443) <= (layer2_outputs(1680)) or (layer2_outputs(5048));
    layer3_outputs(6444) <= not(layer2_outputs(2995));
    layer3_outputs(6445) <= not(layer2_outputs(742));
    layer3_outputs(6446) <= layer2_outputs(4495);
    layer3_outputs(6447) <= not((layer2_outputs(9248)) and (layer2_outputs(5164)));
    layer3_outputs(6448) <= not(layer2_outputs(4367)) or (layer2_outputs(3016));
    layer3_outputs(6449) <= not((layer2_outputs(8570)) and (layer2_outputs(7424)));
    layer3_outputs(6450) <= (layer2_outputs(2126)) and not (layer2_outputs(4654));
    layer3_outputs(6451) <= (layer2_outputs(2332)) xor (layer2_outputs(7352));
    layer3_outputs(6452) <= not((layer2_outputs(8631)) or (layer2_outputs(5735)));
    layer3_outputs(6453) <= not(layer2_outputs(4132));
    layer3_outputs(6454) <= not(layer2_outputs(3771));
    layer3_outputs(6455) <= not(layer2_outputs(6738));
    layer3_outputs(6456) <= not((layer2_outputs(6300)) xor (layer2_outputs(4233)));
    layer3_outputs(6457) <= not(layer2_outputs(6562));
    layer3_outputs(6458) <= (layer2_outputs(3630)) or (layer2_outputs(7381));
    layer3_outputs(6459) <= not(layer2_outputs(4850)) or (layer2_outputs(2306));
    layer3_outputs(6460) <= (layer2_outputs(7976)) and not (layer2_outputs(4906));
    layer3_outputs(6461) <= layer2_outputs(2912);
    layer3_outputs(6462) <= not(layer2_outputs(6098));
    layer3_outputs(6463) <= not(layer2_outputs(4159)) or (layer2_outputs(92));
    layer3_outputs(6464) <= not(layer2_outputs(6316));
    layer3_outputs(6465) <= not((layer2_outputs(3371)) or (layer2_outputs(8716)));
    layer3_outputs(6466) <= not((layer2_outputs(7661)) xor (layer2_outputs(6898)));
    layer3_outputs(6467) <= not(layer2_outputs(8048));
    layer3_outputs(6468) <= layer2_outputs(8888);
    layer3_outputs(6469) <= (layer2_outputs(8499)) xor (layer2_outputs(6596));
    layer3_outputs(6470) <= (layer2_outputs(4290)) or (layer2_outputs(9573));
    layer3_outputs(6471) <= not((layer2_outputs(5985)) xor (layer2_outputs(146)));
    layer3_outputs(6472) <= not((layer2_outputs(9452)) xor (layer2_outputs(5082)));
    layer3_outputs(6473) <= not(layer2_outputs(2494));
    layer3_outputs(6474) <= (layer2_outputs(3825)) and not (layer2_outputs(7793));
    layer3_outputs(6475) <= (layer2_outputs(3488)) or (layer2_outputs(1822));
    layer3_outputs(6476) <= (layer2_outputs(3692)) or (layer2_outputs(4865));
    layer3_outputs(6477) <= (layer2_outputs(2072)) and (layer2_outputs(4162));
    layer3_outputs(6478) <= not(layer2_outputs(2421));
    layer3_outputs(6479) <= not((layer2_outputs(3014)) xor (layer2_outputs(4501)));
    layer3_outputs(6480) <= layer2_outputs(2653);
    layer3_outputs(6481) <= not(layer2_outputs(6553));
    layer3_outputs(6482) <= '1';
    layer3_outputs(6483) <= not(layer2_outputs(7730));
    layer3_outputs(6484) <= not(layer2_outputs(9300));
    layer3_outputs(6485) <= (layer2_outputs(7684)) xor (layer2_outputs(5707));
    layer3_outputs(6486) <= layer2_outputs(2881);
    layer3_outputs(6487) <= layer2_outputs(4964);
    layer3_outputs(6488) <= (layer2_outputs(957)) and not (layer2_outputs(8608));
    layer3_outputs(6489) <= not(layer2_outputs(9818));
    layer3_outputs(6490) <= not(layer2_outputs(6516));
    layer3_outputs(6491) <= layer2_outputs(7259);
    layer3_outputs(6492) <= (layer2_outputs(1994)) and (layer2_outputs(5410));
    layer3_outputs(6493) <= not(layer2_outputs(7616));
    layer3_outputs(6494) <= not(layer2_outputs(7527)) or (layer2_outputs(2585));
    layer3_outputs(6495) <= layer2_outputs(730);
    layer3_outputs(6496) <= (layer2_outputs(6893)) or (layer2_outputs(842));
    layer3_outputs(6497) <= not(layer2_outputs(7279));
    layer3_outputs(6498) <= (layer2_outputs(2439)) and not (layer2_outputs(4201));
    layer3_outputs(6499) <= not((layer2_outputs(9798)) xor (layer2_outputs(6862)));
    layer3_outputs(6500) <= (layer2_outputs(6469)) and (layer2_outputs(453));
    layer3_outputs(6501) <= not(layer2_outputs(4465)) or (layer2_outputs(3758));
    layer3_outputs(6502) <= not((layer2_outputs(4762)) and (layer2_outputs(7980)));
    layer3_outputs(6503) <= (layer2_outputs(7803)) and (layer2_outputs(1000));
    layer3_outputs(6504) <= not(layer2_outputs(7959));
    layer3_outputs(6505) <= not((layer2_outputs(6640)) and (layer2_outputs(9619)));
    layer3_outputs(6506) <= (layer2_outputs(2750)) and (layer2_outputs(4092));
    layer3_outputs(6507) <= not(layer2_outputs(5972));
    layer3_outputs(6508) <= (layer2_outputs(1997)) xor (layer2_outputs(8692));
    layer3_outputs(6509) <= not((layer2_outputs(10094)) and (layer2_outputs(554)));
    layer3_outputs(6510) <= not(layer2_outputs(8798));
    layer3_outputs(6511) <= not(layer2_outputs(7303));
    layer3_outputs(6512) <= not(layer2_outputs(4538));
    layer3_outputs(6513) <= (layer2_outputs(2518)) and not (layer2_outputs(5446));
    layer3_outputs(6514) <= (layer2_outputs(3381)) or (layer2_outputs(3820));
    layer3_outputs(6515) <= (layer2_outputs(9861)) and (layer2_outputs(9921));
    layer3_outputs(6516) <= (layer2_outputs(3531)) or (layer2_outputs(9033));
    layer3_outputs(6517) <= layer2_outputs(1180);
    layer3_outputs(6518) <= not((layer2_outputs(9783)) xor (layer2_outputs(650)));
    layer3_outputs(6519) <= not(layer2_outputs(6342)) or (layer2_outputs(5512));
    layer3_outputs(6520) <= (layer2_outputs(1010)) or (layer2_outputs(9162));
    layer3_outputs(6521) <= layer2_outputs(3055);
    layer3_outputs(6522) <= (layer2_outputs(6333)) or (layer2_outputs(2872));
    layer3_outputs(6523) <= (layer2_outputs(2047)) and not (layer2_outputs(3229));
    layer3_outputs(6524) <= layer2_outputs(2486);
    layer3_outputs(6525) <= not(layer2_outputs(5405)) or (layer2_outputs(2839));
    layer3_outputs(6526) <= (layer2_outputs(6004)) and not (layer2_outputs(4885));
    layer3_outputs(6527) <= not(layer2_outputs(6857)) or (layer2_outputs(3759));
    layer3_outputs(6528) <= (layer2_outputs(7177)) xor (layer2_outputs(9212));
    layer3_outputs(6529) <= (layer2_outputs(5861)) and not (layer2_outputs(9122));
    layer3_outputs(6530) <= not(layer2_outputs(5521));
    layer3_outputs(6531) <= not(layer2_outputs(9562));
    layer3_outputs(6532) <= not(layer2_outputs(4499));
    layer3_outputs(6533) <= layer2_outputs(8242);
    layer3_outputs(6534) <= layer2_outputs(8103);
    layer3_outputs(6535) <= not(layer2_outputs(4290));
    layer3_outputs(6536) <= not(layer2_outputs(3984));
    layer3_outputs(6537) <= (layer2_outputs(5172)) and not (layer2_outputs(7700));
    layer3_outputs(6538) <= (layer2_outputs(2427)) or (layer2_outputs(9432));
    layer3_outputs(6539) <= not(layer2_outputs(4703));
    layer3_outputs(6540) <= (layer2_outputs(8216)) and not (layer2_outputs(3371));
    layer3_outputs(6541) <= not((layer2_outputs(8809)) and (layer2_outputs(2964)));
    layer3_outputs(6542) <= layer2_outputs(4292);
    layer3_outputs(6543) <= layer2_outputs(7598);
    layer3_outputs(6544) <= (layer2_outputs(1453)) and not (layer2_outputs(4576));
    layer3_outputs(6545) <= layer2_outputs(6172);
    layer3_outputs(6546) <= not(layer2_outputs(1726));
    layer3_outputs(6547) <= layer2_outputs(6825);
    layer3_outputs(6548) <= not(layer2_outputs(4916));
    layer3_outputs(6549) <= (layer2_outputs(7859)) and not (layer2_outputs(8673));
    layer3_outputs(6550) <= not((layer2_outputs(3369)) xor (layer2_outputs(1145)));
    layer3_outputs(6551) <= not(layer2_outputs(8308));
    layer3_outputs(6552) <= (layer2_outputs(9170)) and not (layer2_outputs(9252));
    layer3_outputs(6553) <= not((layer2_outputs(9745)) xor (layer2_outputs(3110)));
    layer3_outputs(6554) <= not(layer2_outputs(5307));
    layer3_outputs(6555) <= not(layer2_outputs(5841));
    layer3_outputs(6556) <= layer2_outputs(6866);
    layer3_outputs(6557) <= not(layer2_outputs(1853));
    layer3_outputs(6558) <= not(layer2_outputs(5385));
    layer3_outputs(6559) <= layer2_outputs(8039);
    layer3_outputs(6560) <= layer2_outputs(5796);
    layer3_outputs(6561) <= layer2_outputs(5087);
    layer3_outputs(6562) <= not(layer2_outputs(2711));
    layer3_outputs(6563) <= layer2_outputs(3304);
    layer3_outputs(6564) <= (layer2_outputs(6353)) or (layer2_outputs(1539));
    layer3_outputs(6565) <= layer2_outputs(7426);
    layer3_outputs(6566) <= not((layer2_outputs(8362)) xor (layer2_outputs(7058)));
    layer3_outputs(6567) <= '1';
    layer3_outputs(6568) <= (layer2_outputs(5345)) xor (layer2_outputs(6352));
    layer3_outputs(6569) <= not((layer2_outputs(6363)) xor (layer2_outputs(6285)));
    layer3_outputs(6570) <= not(layer2_outputs(3220));
    layer3_outputs(6571) <= (layer2_outputs(9182)) and not (layer2_outputs(9508));
    layer3_outputs(6572) <= not(layer2_outputs(9959)) or (layer2_outputs(4174));
    layer3_outputs(6573) <= not((layer2_outputs(8523)) and (layer2_outputs(5742)));
    layer3_outputs(6574) <= not(layer2_outputs(5213));
    layer3_outputs(6575) <= '1';
    layer3_outputs(6576) <= not(layer2_outputs(97)) or (layer2_outputs(4641));
    layer3_outputs(6577) <= layer2_outputs(7387);
    layer3_outputs(6578) <= not(layer2_outputs(1350)) or (layer2_outputs(67));
    layer3_outputs(6579) <= layer2_outputs(568);
    layer3_outputs(6580) <= not(layer2_outputs(5182));
    layer3_outputs(6581) <= not((layer2_outputs(5790)) or (layer2_outputs(9816)));
    layer3_outputs(6582) <= layer2_outputs(4395);
    layer3_outputs(6583) <= layer2_outputs(7175);
    layer3_outputs(6584) <= layer2_outputs(4119);
    layer3_outputs(6585) <= layer2_outputs(6661);
    layer3_outputs(6586) <= layer2_outputs(4951);
    layer3_outputs(6587) <= not(layer2_outputs(4098));
    layer3_outputs(6588) <= not(layer2_outputs(2247));
    layer3_outputs(6589) <= not(layer2_outputs(6854)) or (layer2_outputs(9689));
    layer3_outputs(6590) <= not(layer2_outputs(7631));
    layer3_outputs(6591) <= layer2_outputs(6785);
    layer3_outputs(6592) <= (layer2_outputs(3597)) xor (layer2_outputs(7436));
    layer3_outputs(6593) <= not(layer2_outputs(6024));
    layer3_outputs(6594) <= layer2_outputs(6084);
    layer3_outputs(6595) <= layer2_outputs(4372);
    layer3_outputs(6596) <= layer2_outputs(9536);
    layer3_outputs(6597) <= (layer2_outputs(8310)) and not (layer2_outputs(1300));
    layer3_outputs(6598) <= not(layer2_outputs(264)) or (layer2_outputs(815));
    layer3_outputs(6599) <= layer2_outputs(1698);
    layer3_outputs(6600) <= (layer2_outputs(2214)) xor (layer2_outputs(9646));
    layer3_outputs(6601) <= layer2_outputs(807);
    layer3_outputs(6602) <= '0';
    layer3_outputs(6603) <= (layer2_outputs(9234)) and not (layer2_outputs(8105));
    layer3_outputs(6604) <= not(layer2_outputs(7781));
    layer3_outputs(6605) <= (layer2_outputs(4717)) and (layer2_outputs(6499));
    layer3_outputs(6606) <= not(layer2_outputs(4540)) or (layer2_outputs(2468));
    layer3_outputs(6607) <= layer2_outputs(781);
    layer3_outputs(6608) <= not(layer2_outputs(1559));
    layer3_outputs(6609) <= layer2_outputs(2012);
    layer3_outputs(6610) <= not(layer2_outputs(8900));
    layer3_outputs(6611) <= not(layer2_outputs(2485));
    layer3_outputs(6612) <= not((layer2_outputs(4453)) and (layer2_outputs(7404)));
    layer3_outputs(6613) <= not(layer2_outputs(2806));
    layer3_outputs(6614) <= (layer2_outputs(34)) and not (layer2_outputs(836));
    layer3_outputs(6615) <= not((layer2_outputs(9406)) xor (layer2_outputs(6213)));
    layer3_outputs(6616) <= '1';
    layer3_outputs(6617) <= not(layer2_outputs(724));
    layer3_outputs(6618) <= not(layer2_outputs(2641));
    layer3_outputs(6619) <= (layer2_outputs(8857)) or (layer2_outputs(1272));
    layer3_outputs(6620) <= not(layer2_outputs(5271));
    layer3_outputs(6621) <= not((layer2_outputs(7718)) xor (layer2_outputs(2525)));
    layer3_outputs(6622) <= '0';
    layer3_outputs(6623) <= (layer2_outputs(1886)) and not (layer2_outputs(1396));
    layer3_outputs(6624) <= layer2_outputs(6203);
    layer3_outputs(6625) <= (layer2_outputs(5090)) xor (layer2_outputs(7698));
    layer3_outputs(6626) <= not(layer2_outputs(2156)) or (layer2_outputs(9276));
    layer3_outputs(6627) <= not((layer2_outputs(3801)) xor (layer2_outputs(5032)));
    layer3_outputs(6628) <= not(layer2_outputs(4057)) or (layer2_outputs(7483));
    layer3_outputs(6629) <= layer2_outputs(1822);
    layer3_outputs(6630) <= not(layer2_outputs(8547)) or (layer2_outputs(224));
    layer3_outputs(6631) <= layer2_outputs(4458);
    layer3_outputs(6632) <= (layer2_outputs(1258)) or (layer2_outputs(5627));
    layer3_outputs(6633) <= not(layer2_outputs(7194)) or (layer2_outputs(6607));
    layer3_outputs(6634) <= not((layer2_outputs(229)) and (layer2_outputs(2197)));
    layer3_outputs(6635) <= not(layer2_outputs(8009));
    layer3_outputs(6636) <= layer2_outputs(7491);
    layer3_outputs(6637) <= layer2_outputs(9927);
    layer3_outputs(6638) <= not((layer2_outputs(6348)) and (layer2_outputs(1319)));
    layer3_outputs(6639) <= not(layer2_outputs(8762));
    layer3_outputs(6640) <= not((layer2_outputs(8642)) and (layer2_outputs(5671)));
    layer3_outputs(6641) <= (layer2_outputs(9472)) xor (layer2_outputs(4026));
    layer3_outputs(6642) <= (layer2_outputs(5110)) and not (layer2_outputs(8947));
    layer3_outputs(6643) <= '1';
    layer3_outputs(6644) <= (layer2_outputs(1890)) and not (layer2_outputs(6131));
    layer3_outputs(6645) <= not((layer2_outputs(5074)) and (layer2_outputs(3729)));
    layer3_outputs(6646) <= not((layer2_outputs(7138)) and (layer2_outputs(3340)));
    layer3_outputs(6647) <= not(layer2_outputs(8768));
    layer3_outputs(6648) <= not(layer2_outputs(10108));
    layer3_outputs(6649) <= (layer2_outputs(6518)) and (layer2_outputs(5568));
    layer3_outputs(6650) <= (layer2_outputs(2234)) and not (layer2_outputs(6402));
    layer3_outputs(6651) <= not(layer2_outputs(8511));
    layer3_outputs(6652) <= not(layer2_outputs(118));
    layer3_outputs(6653) <= layer2_outputs(4981);
    layer3_outputs(6654) <= layer2_outputs(5666);
    layer3_outputs(6655) <= not(layer2_outputs(2118));
    layer3_outputs(6656) <= layer2_outputs(1467);
    layer3_outputs(6657) <= layer2_outputs(5065);
    layer3_outputs(6658) <= '0';
    layer3_outputs(6659) <= layer2_outputs(6447);
    layer3_outputs(6660) <= layer2_outputs(5216);
    layer3_outputs(6661) <= '0';
    layer3_outputs(6662) <= not(layer2_outputs(10216)) or (layer2_outputs(2845));
    layer3_outputs(6663) <= layer2_outputs(4274);
    layer3_outputs(6664) <= layer2_outputs(3950);
    layer3_outputs(6665) <= layer2_outputs(4110);
    layer3_outputs(6666) <= not(layer2_outputs(8151)) or (layer2_outputs(6457));
    layer3_outputs(6667) <= not(layer2_outputs(5781));
    layer3_outputs(6668) <= not(layer2_outputs(8926));
    layer3_outputs(6669) <= not(layer2_outputs(1349));
    layer3_outputs(6670) <= not(layer2_outputs(580));
    layer3_outputs(6671) <= (layer2_outputs(6427)) and not (layer2_outputs(1581));
    layer3_outputs(6672) <= (layer2_outputs(9781)) xor (layer2_outputs(9940));
    layer3_outputs(6673) <= not(layer2_outputs(363));
    layer3_outputs(6674) <= not((layer2_outputs(540)) or (layer2_outputs(5540)));
    layer3_outputs(6675) <= not((layer2_outputs(8265)) and (layer2_outputs(559)));
    layer3_outputs(6676) <= not((layer2_outputs(5626)) xor (layer2_outputs(2227)));
    layer3_outputs(6677) <= not(layer2_outputs(6634)) or (layer2_outputs(3290));
    layer3_outputs(6678) <= not(layer2_outputs(195)) or (layer2_outputs(7353));
    layer3_outputs(6679) <= not((layer2_outputs(707)) xor (layer2_outputs(9236)));
    layer3_outputs(6680) <= not(layer2_outputs(6540));
    layer3_outputs(6681) <= not(layer2_outputs(274));
    layer3_outputs(6682) <= not(layer2_outputs(8535));
    layer3_outputs(6683) <= not(layer2_outputs(1718)) or (layer2_outputs(1393));
    layer3_outputs(6684) <= (layer2_outputs(9297)) or (layer2_outputs(1196));
    layer3_outputs(6685) <= not(layer2_outputs(5864));
    layer3_outputs(6686) <= not((layer2_outputs(1717)) xor (layer2_outputs(7099)));
    layer3_outputs(6687) <= not(layer2_outputs(7057));
    layer3_outputs(6688) <= not(layer2_outputs(4580));
    layer3_outputs(6689) <= not((layer2_outputs(2050)) xor (layer2_outputs(9101)));
    layer3_outputs(6690) <= (layer2_outputs(8831)) and (layer2_outputs(8917));
    layer3_outputs(6691) <= layer2_outputs(897);
    layer3_outputs(6692) <= (layer2_outputs(132)) xor (layer2_outputs(9473));
    layer3_outputs(6693) <= layer2_outputs(1606);
    layer3_outputs(6694) <= not((layer2_outputs(4606)) xor (layer2_outputs(3403)));
    layer3_outputs(6695) <= (layer2_outputs(2112)) or (layer2_outputs(5942));
    layer3_outputs(6696) <= not((layer2_outputs(526)) xor (layer2_outputs(9489)));
    layer3_outputs(6697) <= layer2_outputs(6369);
    layer3_outputs(6698) <= (layer2_outputs(4352)) and (layer2_outputs(8148));
    layer3_outputs(6699) <= '1';
    layer3_outputs(6700) <= (layer2_outputs(2970)) and not (layer2_outputs(5352));
    layer3_outputs(6701) <= (layer2_outputs(5893)) and not (layer2_outputs(1838));
    layer3_outputs(6702) <= not(layer2_outputs(5453));
    layer3_outputs(6703) <= not(layer2_outputs(5778));
    layer3_outputs(6704) <= not((layer2_outputs(8594)) and (layer2_outputs(9000)));
    layer3_outputs(6705) <= (layer2_outputs(1736)) and (layer2_outputs(8542));
    layer3_outputs(6706) <= not((layer2_outputs(4944)) or (layer2_outputs(2353)));
    layer3_outputs(6707) <= (layer2_outputs(5798)) and not (layer2_outputs(8563));
    layer3_outputs(6708) <= (layer2_outputs(2266)) xor (layer2_outputs(1654));
    layer3_outputs(6709) <= not(layer2_outputs(1005)) or (layer2_outputs(4293));
    layer3_outputs(6710) <= (layer2_outputs(6154)) and not (layer2_outputs(7828));
    layer3_outputs(6711) <= (layer2_outputs(8915)) and not (layer2_outputs(39));
    layer3_outputs(6712) <= layer2_outputs(5603);
    layer3_outputs(6713) <= not(layer2_outputs(1351));
    layer3_outputs(6714) <= not(layer2_outputs(8601));
    layer3_outputs(6715) <= not((layer2_outputs(1049)) and (layer2_outputs(331)));
    layer3_outputs(6716) <= (layer2_outputs(3997)) and not (layer2_outputs(8199));
    layer3_outputs(6717) <= not((layer2_outputs(6942)) or (layer2_outputs(4695)));
    layer3_outputs(6718) <= layer2_outputs(2644);
    layer3_outputs(6719) <= (layer2_outputs(3192)) xor (layer2_outputs(6102));
    layer3_outputs(6720) <= not(layer2_outputs(288)) or (layer2_outputs(6417));
    layer3_outputs(6721) <= not(layer2_outputs(5661));
    layer3_outputs(6722) <= layer2_outputs(6003);
    layer3_outputs(6723) <= (layer2_outputs(4035)) and not (layer2_outputs(5553));
    layer3_outputs(6724) <= layer2_outputs(7351);
    layer3_outputs(6725) <= layer2_outputs(8621);
    layer3_outputs(6726) <= '0';
    layer3_outputs(6727) <= not((layer2_outputs(9852)) and (layer2_outputs(8791)));
    layer3_outputs(6728) <= not((layer2_outputs(9732)) and (layer2_outputs(3306)));
    layer3_outputs(6729) <= not((layer2_outputs(5946)) or (layer2_outputs(8388)));
    layer3_outputs(6730) <= not(layer2_outputs(8338));
    layer3_outputs(6731) <= not(layer2_outputs(760));
    layer3_outputs(6732) <= '1';
    layer3_outputs(6733) <= (layer2_outputs(7143)) xor (layer2_outputs(8147));
    layer3_outputs(6734) <= layer2_outputs(5520);
    layer3_outputs(6735) <= layer2_outputs(7138);
    layer3_outputs(6736) <= layer2_outputs(3194);
    layer3_outputs(6737) <= (layer2_outputs(8541)) and not (layer2_outputs(4040));
    layer3_outputs(6738) <= (layer2_outputs(4610)) xor (layer2_outputs(5083));
    layer3_outputs(6739) <= layer2_outputs(3116);
    layer3_outputs(6740) <= (layer2_outputs(722)) and not (layer2_outputs(1473));
    layer3_outputs(6741) <= not(layer2_outputs(2612));
    layer3_outputs(6742) <= not((layer2_outputs(964)) xor (layer2_outputs(1197)));
    layer3_outputs(6743) <= not(layer2_outputs(7002));
    layer3_outputs(6744) <= not(layer2_outputs(6359));
    layer3_outputs(6745) <= not(layer2_outputs(4690)) or (layer2_outputs(23));
    layer3_outputs(6746) <= not((layer2_outputs(1962)) and (layer2_outputs(7631)));
    layer3_outputs(6747) <= layer2_outputs(4143);
    layer3_outputs(6748) <= not((layer2_outputs(6965)) or (layer2_outputs(5541)));
    layer3_outputs(6749) <= not((layer2_outputs(831)) xor (layer2_outputs(4601)));
    layer3_outputs(6750) <= not(layer2_outputs(7585));
    layer3_outputs(6751) <= not((layer2_outputs(9201)) or (layer2_outputs(5724)));
    layer3_outputs(6752) <= (layer2_outputs(8352)) and (layer2_outputs(5371));
    layer3_outputs(6753) <= not((layer2_outputs(5282)) xor (layer2_outputs(1524)));
    layer3_outputs(6754) <= not(layer2_outputs(1100));
    layer3_outputs(6755) <= not((layer2_outputs(9954)) or (layer2_outputs(5332)));
    layer3_outputs(6756) <= (layer2_outputs(2642)) and not (layer2_outputs(2952));
    layer3_outputs(6757) <= layer2_outputs(2628);
    layer3_outputs(6758) <= not(layer2_outputs(184)) or (layer2_outputs(1923));
    layer3_outputs(6759) <= not((layer2_outputs(3866)) and (layer2_outputs(8382)));
    layer3_outputs(6760) <= not((layer2_outputs(5147)) and (layer2_outputs(3809)));
    layer3_outputs(6761) <= not(layer2_outputs(3126));
    layer3_outputs(6762) <= not((layer2_outputs(316)) and (layer2_outputs(4362)));
    layer3_outputs(6763) <= layer2_outputs(1207);
    layer3_outputs(6764) <= not(layer2_outputs(2289));
    layer3_outputs(6765) <= not((layer2_outputs(1361)) xor (layer2_outputs(1153)));
    layer3_outputs(6766) <= (layer2_outputs(1237)) and not (layer2_outputs(4586));
    layer3_outputs(6767) <= not(layer2_outputs(485));
    layer3_outputs(6768) <= layer2_outputs(4359);
    layer3_outputs(6769) <= not(layer2_outputs(974));
    layer3_outputs(6770) <= not(layer2_outputs(8586));
    layer3_outputs(6771) <= not(layer2_outputs(6218));
    layer3_outputs(6772) <= not(layer2_outputs(888));
    layer3_outputs(6773) <= not(layer2_outputs(3555)) or (layer2_outputs(1053));
    layer3_outputs(6774) <= not((layer2_outputs(5776)) or (layer2_outputs(246)));
    layer3_outputs(6775) <= layer2_outputs(7237);
    layer3_outputs(6776) <= not(layer2_outputs(635));
    layer3_outputs(6777) <= not((layer2_outputs(7862)) xor (layer2_outputs(9607)));
    layer3_outputs(6778) <= not(layer2_outputs(2400));
    layer3_outputs(6779) <= layer2_outputs(8090);
    layer3_outputs(6780) <= not(layer2_outputs(6672));
    layer3_outputs(6781) <= not(layer2_outputs(5709));
    layer3_outputs(6782) <= not((layer2_outputs(7107)) or (layer2_outputs(493)));
    layer3_outputs(6783) <= (layer2_outputs(643)) and (layer2_outputs(2451));
    layer3_outputs(6784) <= not((layer2_outputs(4599)) xor (layer2_outputs(916)));
    layer3_outputs(6785) <= (layer2_outputs(1796)) and not (layer2_outputs(1580));
    layer3_outputs(6786) <= (layer2_outputs(9935)) xor (layer2_outputs(4844));
    layer3_outputs(6787) <= not(layer2_outputs(5639));
    layer3_outputs(6788) <= layer2_outputs(7453);
    layer3_outputs(6789) <= not(layer2_outputs(332));
    layer3_outputs(6790) <= not(layer2_outputs(1982));
    layer3_outputs(6791) <= (layer2_outputs(4990)) and (layer2_outputs(3560));
    layer3_outputs(6792) <= layer2_outputs(6706);
    layer3_outputs(6793) <= not((layer2_outputs(4129)) or (layer2_outputs(879)));
    layer3_outputs(6794) <= (layer2_outputs(10131)) and (layer2_outputs(4664));
    layer3_outputs(6795) <= (layer2_outputs(6888)) and not (layer2_outputs(8515));
    layer3_outputs(6796) <= not(layer2_outputs(9678)) or (layer2_outputs(2961));
    layer3_outputs(6797) <= not(layer2_outputs(7047)) or (layer2_outputs(2477));
    layer3_outputs(6798) <= (layer2_outputs(5694)) and (layer2_outputs(6989));
    layer3_outputs(6799) <= not((layer2_outputs(3067)) and (layer2_outputs(5305)));
    layer3_outputs(6800) <= layer2_outputs(936);
    layer3_outputs(6801) <= layer2_outputs(7486);
    layer3_outputs(6802) <= not((layer2_outputs(1288)) and (layer2_outputs(5360)));
    layer3_outputs(6803) <= not(layer2_outputs(7588)) or (layer2_outputs(255));
    layer3_outputs(6804) <= not(layer2_outputs(1985));
    layer3_outputs(6805) <= (layer2_outputs(1046)) and not (layer2_outputs(2978));
    layer3_outputs(6806) <= not(layer2_outputs(8380)) or (layer2_outputs(2516));
    layer3_outputs(6807) <= (layer2_outputs(934)) xor (layer2_outputs(3548));
    layer3_outputs(6808) <= (layer2_outputs(4650)) xor (layer2_outputs(5328));
    layer3_outputs(6809) <= not(layer2_outputs(9880)) or (layer2_outputs(9760));
    layer3_outputs(6810) <= not(layer2_outputs(7491));
    layer3_outputs(6811) <= not(layer2_outputs(9476));
    layer3_outputs(6812) <= (layer2_outputs(9422)) xor (layer2_outputs(5276));
    layer3_outputs(6813) <= (layer2_outputs(1050)) or (layer2_outputs(595));
    layer3_outputs(6814) <= (layer2_outputs(10003)) and (layer2_outputs(1165));
    layer3_outputs(6815) <= not(layer2_outputs(8424));
    layer3_outputs(6816) <= layer2_outputs(2697);
    layer3_outputs(6817) <= layer2_outputs(6772);
    layer3_outputs(6818) <= layer2_outputs(9366);
    layer3_outputs(6819) <= (layer2_outputs(293)) xor (layer2_outputs(723));
    layer3_outputs(6820) <= not(layer2_outputs(8927)) or (layer2_outputs(9549));
    layer3_outputs(6821) <= (layer2_outputs(7542)) or (layer2_outputs(3951));
    layer3_outputs(6822) <= not(layer2_outputs(9135));
    layer3_outputs(6823) <= not(layer2_outputs(3992));
    layer3_outputs(6824) <= (layer2_outputs(2005)) and (layer2_outputs(5939));
    layer3_outputs(6825) <= layer2_outputs(10163);
    layer3_outputs(6826) <= not(layer2_outputs(1304));
    layer3_outputs(6827) <= layer2_outputs(3097);
    layer3_outputs(6828) <= not(layer2_outputs(8811)) or (layer2_outputs(9591));
    layer3_outputs(6829) <= not(layer2_outputs(7736));
    layer3_outputs(6830) <= layer2_outputs(3069);
    layer3_outputs(6831) <= not(layer2_outputs(8285));
    layer3_outputs(6832) <= not(layer2_outputs(4867)) or (layer2_outputs(9389));
    layer3_outputs(6833) <= '1';
    layer3_outputs(6834) <= (layer2_outputs(3186)) or (layer2_outputs(1042));
    layer3_outputs(6835) <= not(layer2_outputs(1290));
    layer3_outputs(6836) <= layer2_outputs(6971);
    layer3_outputs(6837) <= layer2_outputs(5256);
    layer3_outputs(6838) <= (layer2_outputs(7051)) or (layer2_outputs(7228));
    layer3_outputs(6839) <= layer2_outputs(1202);
    layer3_outputs(6840) <= not((layer2_outputs(1308)) and (layer2_outputs(344)));
    layer3_outputs(6841) <= not(layer2_outputs(2176));
    layer3_outputs(6842) <= not(layer2_outputs(7504));
    layer3_outputs(6843) <= not(layer2_outputs(7394));
    layer3_outputs(6844) <= layer2_outputs(5535);
    layer3_outputs(6845) <= (layer2_outputs(9462)) and not (layer2_outputs(7386));
    layer3_outputs(6846) <= not(layer2_outputs(3276)) or (layer2_outputs(5265));
    layer3_outputs(6847) <= layer2_outputs(8185);
    layer3_outputs(6848) <= not(layer2_outputs(6838));
    layer3_outputs(6849) <= not(layer2_outputs(5363));
    layer3_outputs(6850) <= not(layer2_outputs(1166));
    layer3_outputs(6851) <= layer2_outputs(7305);
    layer3_outputs(6852) <= (layer2_outputs(7756)) xor (layer2_outputs(7029));
    layer3_outputs(6853) <= layer2_outputs(6767);
    layer3_outputs(6854) <= (layer2_outputs(7361)) or (layer2_outputs(1914));
    layer3_outputs(6855) <= layer2_outputs(389);
    layer3_outputs(6856) <= layer2_outputs(8061);
    layer3_outputs(6857) <= not(layer2_outputs(136)) or (layer2_outputs(8111));
    layer3_outputs(6858) <= not(layer2_outputs(6025)) or (layer2_outputs(5327));
    layer3_outputs(6859) <= not((layer2_outputs(6079)) and (layer2_outputs(5929)));
    layer3_outputs(6860) <= layer2_outputs(6703);
    layer3_outputs(6861) <= (layer2_outputs(7681)) and not (layer2_outputs(2791));
    layer3_outputs(6862) <= not(layer2_outputs(8008));
    layer3_outputs(6863) <= not((layer2_outputs(366)) or (layer2_outputs(520)));
    layer3_outputs(6864) <= not(layer2_outputs(2780)) or (layer2_outputs(6473));
    layer3_outputs(6865) <= layer2_outputs(2637);
    layer3_outputs(6866) <= layer2_outputs(7024);
    layer3_outputs(6867) <= not(layer2_outputs(3229)) or (layer2_outputs(9842));
    layer3_outputs(6868) <= layer2_outputs(409);
    layer3_outputs(6869) <= (layer2_outputs(2293)) xor (layer2_outputs(6320));
    layer3_outputs(6870) <= '0';
    layer3_outputs(6871) <= (layer2_outputs(7943)) and not (layer2_outputs(9215));
    layer3_outputs(6872) <= not(layer2_outputs(8159));
    layer3_outputs(6873) <= '0';
    layer3_outputs(6874) <= '0';
    layer3_outputs(6875) <= (layer2_outputs(2424)) or (layer2_outputs(4599));
    layer3_outputs(6876) <= not(layer2_outputs(6896));
    layer3_outputs(6877) <= (layer2_outputs(5354)) and (layer2_outputs(10238));
    layer3_outputs(6878) <= not((layer2_outputs(5610)) or (layer2_outputs(8836)));
    layer3_outputs(6879) <= not((layer2_outputs(9765)) xor (layer2_outputs(3470)));
    layer3_outputs(6880) <= not(layer2_outputs(4660));
    layer3_outputs(6881) <= layer2_outputs(6297);
    layer3_outputs(6882) <= (layer2_outputs(5080)) or (layer2_outputs(5440));
    layer3_outputs(6883) <= not(layer2_outputs(10080));
    layer3_outputs(6884) <= not(layer2_outputs(5235));
    layer3_outputs(6885) <= not(layer2_outputs(3121));
    layer3_outputs(6886) <= layer2_outputs(5373);
    layer3_outputs(6887) <= not(layer2_outputs(7403));
    layer3_outputs(6888) <= (layer2_outputs(616)) and (layer2_outputs(3526));
    layer3_outputs(6889) <= not(layer2_outputs(9073));
    layer3_outputs(6890) <= (layer2_outputs(1141)) and not (layer2_outputs(5223));
    layer3_outputs(6891) <= not(layer2_outputs(7618)) or (layer2_outputs(8994));
    layer3_outputs(6892) <= not(layer2_outputs(10026));
    layer3_outputs(6893) <= not((layer2_outputs(1479)) and (layer2_outputs(9387)));
    layer3_outputs(6894) <= layer2_outputs(4072);
    layer3_outputs(6895) <= not(layer2_outputs(5584));
    layer3_outputs(6896) <= not(layer2_outputs(3776));
    layer3_outputs(6897) <= layer2_outputs(1298);
    layer3_outputs(6898) <= not((layer2_outputs(6650)) xor (layer2_outputs(7789)));
    layer3_outputs(6899) <= not(layer2_outputs(6031));
    layer3_outputs(6900) <= (layer2_outputs(5622)) or (layer2_outputs(7279));
    layer3_outputs(6901) <= layer2_outputs(4953);
    layer3_outputs(6902) <= not(layer2_outputs(10107));
    layer3_outputs(6903) <= not(layer2_outputs(4665));
    layer3_outputs(6904) <= not(layer2_outputs(4775));
    layer3_outputs(6905) <= layer2_outputs(951);
    layer3_outputs(6906) <= (layer2_outputs(2847)) or (layer2_outputs(5105));
    layer3_outputs(6907) <= not((layer2_outputs(1516)) and (layer2_outputs(4009)));
    layer3_outputs(6908) <= not(layer2_outputs(7834));
    layer3_outputs(6909) <= (layer2_outputs(7872)) or (layer2_outputs(3021));
    layer3_outputs(6910) <= not(layer2_outputs(2358));
    layer3_outputs(6911) <= not(layer2_outputs(8576));
    layer3_outputs(6912) <= layer2_outputs(9817);
    layer3_outputs(6913) <= layer2_outputs(4707);
    layer3_outputs(6914) <= not(layer2_outputs(2499)) or (layer2_outputs(6656));
    layer3_outputs(6915) <= layer2_outputs(2561);
    layer3_outputs(6916) <= layer2_outputs(6394);
    layer3_outputs(6917) <= not(layer2_outputs(1345)) or (layer2_outputs(3917));
    layer3_outputs(6918) <= (layer2_outputs(3436)) xor (layer2_outputs(5331));
    layer3_outputs(6919) <= not((layer2_outputs(6849)) and (layer2_outputs(9864)));
    layer3_outputs(6920) <= not((layer2_outputs(7871)) xor (layer2_outputs(10105)));
    layer3_outputs(6921) <= not(layer2_outputs(7523));
    layer3_outputs(6922) <= not((layer2_outputs(6806)) xor (layer2_outputs(5053)));
    layer3_outputs(6923) <= (layer2_outputs(9732)) and not (layer2_outputs(1588));
    layer3_outputs(6924) <= not((layer2_outputs(10065)) or (layer2_outputs(2240)));
    layer3_outputs(6925) <= (layer2_outputs(5939)) and not (layer2_outputs(224));
    layer3_outputs(6926) <= (layer2_outputs(3621)) and not (layer2_outputs(9710));
    layer3_outputs(6927) <= not(layer2_outputs(9495)) or (layer2_outputs(9534));
    layer3_outputs(6928) <= layer2_outputs(348);
    layer3_outputs(6929) <= not(layer2_outputs(4472));
    layer3_outputs(6930) <= not(layer2_outputs(6677));
    layer3_outputs(6931) <= not(layer2_outputs(5117));
    layer3_outputs(6932) <= (layer2_outputs(4425)) xor (layer2_outputs(113));
    layer3_outputs(6933) <= not((layer2_outputs(4894)) xor (layer2_outputs(4961)));
    layer3_outputs(6934) <= '1';
    layer3_outputs(6935) <= '1';
    layer3_outputs(6936) <= layer2_outputs(1045);
    layer3_outputs(6937) <= not((layer2_outputs(3124)) or (layer2_outputs(6577)));
    layer3_outputs(6938) <= layer2_outputs(4834);
    layer3_outputs(6939) <= layer2_outputs(6037);
    layer3_outputs(6940) <= layer2_outputs(8790);
    layer3_outputs(6941) <= not((layer2_outputs(7302)) and (layer2_outputs(2651)));
    layer3_outputs(6942) <= (layer2_outputs(908)) or (layer2_outputs(9822));
    layer3_outputs(6943) <= layer2_outputs(798);
    layer3_outputs(6944) <= layer2_outputs(355);
    layer3_outputs(6945) <= not(layer2_outputs(756));
    layer3_outputs(6946) <= layer2_outputs(9693);
    layer3_outputs(6947) <= not(layer2_outputs(1088)) or (layer2_outputs(3532));
    layer3_outputs(6948) <= (layer2_outputs(185)) and not (layer2_outputs(6456));
    layer3_outputs(6949) <= not(layer2_outputs(7099)) or (layer2_outputs(5349));
    layer3_outputs(6950) <= not(layer2_outputs(9486));
    layer3_outputs(6951) <= not(layer2_outputs(6193));
    layer3_outputs(6952) <= layer2_outputs(4146);
    layer3_outputs(6953) <= (layer2_outputs(8346)) xor (layer2_outputs(2440));
    layer3_outputs(6954) <= not(layer2_outputs(8646));
    layer3_outputs(6955) <= not(layer2_outputs(2910));
    layer3_outputs(6956) <= layer2_outputs(2734);
    layer3_outputs(6957) <= not((layer2_outputs(9296)) xor (layer2_outputs(4871)));
    layer3_outputs(6958) <= not(layer2_outputs(3148));
    layer3_outputs(6959) <= not(layer2_outputs(1233));
    layer3_outputs(6960) <= not((layer2_outputs(10023)) xor (layer2_outputs(8493)));
    layer3_outputs(6961) <= not(layer2_outputs(1156)) or (layer2_outputs(5438));
    layer3_outputs(6962) <= (layer2_outputs(4374)) and not (layer2_outputs(8992));
    layer3_outputs(6963) <= (layer2_outputs(3128)) xor (layer2_outputs(8531));
    layer3_outputs(6964) <= not((layer2_outputs(5375)) xor (layer2_outputs(7674)));
    layer3_outputs(6965) <= not((layer2_outputs(2606)) or (layer2_outputs(57)));
    layer3_outputs(6966) <= layer2_outputs(1140);
    layer3_outputs(6967) <= '0';
    layer3_outputs(6968) <= '1';
    layer3_outputs(6969) <= not(layer2_outputs(4684));
    layer3_outputs(6970) <= layer2_outputs(8449);
    layer3_outputs(6971) <= (layer2_outputs(6217)) xor (layer2_outputs(433));
    layer3_outputs(6972) <= layer2_outputs(5119);
    layer3_outputs(6973) <= not(layer2_outputs(4909));
    layer3_outputs(6974) <= layer2_outputs(6723);
    layer3_outputs(6975) <= layer2_outputs(3113);
    layer3_outputs(6976) <= (layer2_outputs(6492)) or (layer2_outputs(2376));
    layer3_outputs(6977) <= not(layer2_outputs(6959));
    layer3_outputs(6978) <= layer2_outputs(8189);
    layer3_outputs(6979) <= not((layer2_outputs(9165)) and (layer2_outputs(699)));
    layer3_outputs(6980) <= not(layer2_outputs(7349)) or (layer2_outputs(7123));
    layer3_outputs(6981) <= not(layer2_outputs(3534));
    layer3_outputs(6982) <= not((layer2_outputs(9808)) and (layer2_outputs(4714)));
    layer3_outputs(6983) <= not(layer2_outputs(4047));
    layer3_outputs(6984) <= layer2_outputs(6957);
    layer3_outputs(6985) <= not(layer2_outputs(7687));
    layer3_outputs(6986) <= not((layer2_outputs(6561)) and (layer2_outputs(2307)));
    layer3_outputs(6987) <= not(layer2_outputs(7619));
    layer3_outputs(6988) <= layer2_outputs(3901);
    layer3_outputs(6989) <= not(layer2_outputs(7428)) or (layer2_outputs(7145));
    layer3_outputs(6990) <= not(layer2_outputs(4152));
    layer3_outputs(6991) <= not(layer2_outputs(8561)) or (layer2_outputs(7672));
    layer3_outputs(6992) <= (layer2_outputs(9467)) and (layer2_outputs(17));
    layer3_outputs(6993) <= layer2_outputs(9164);
    layer3_outputs(6994) <= (layer2_outputs(335)) xor (layer2_outputs(388));
    layer3_outputs(6995) <= layer2_outputs(3372);
    layer3_outputs(6996) <= not(layer2_outputs(381));
    layer3_outputs(6997) <= (layer2_outputs(5953)) and (layer2_outputs(1415));
    layer3_outputs(6998) <= not(layer2_outputs(4140));
    layer3_outputs(6999) <= not(layer2_outputs(2071)) or (layer2_outputs(1513));
    layer3_outputs(7000) <= not((layer2_outputs(8311)) or (layer2_outputs(4845)));
    layer3_outputs(7001) <= (layer2_outputs(1453)) and not (layer2_outputs(4750));
    layer3_outputs(7002) <= (layer2_outputs(1351)) and not (layer2_outputs(7064));
    layer3_outputs(7003) <= layer2_outputs(7730);
    layer3_outputs(7004) <= not(layer2_outputs(5915));
    layer3_outputs(7005) <= not((layer2_outputs(3244)) and (layer2_outputs(1892)));
    layer3_outputs(7006) <= layer2_outputs(10105);
    layer3_outputs(7007) <= not((layer2_outputs(9061)) xor (layer2_outputs(1228)));
    layer3_outputs(7008) <= not(layer2_outputs(3894));
    layer3_outputs(7009) <= (layer2_outputs(5519)) and not (layer2_outputs(3685));
    layer3_outputs(7010) <= not(layer2_outputs(246));
    layer3_outputs(7011) <= not(layer2_outputs(6115));
    layer3_outputs(7012) <= layer2_outputs(8238);
    layer3_outputs(7013) <= layer2_outputs(2387);
    layer3_outputs(7014) <= not(layer2_outputs(60));
    layer3_outputs(7015) <= layer2_outputs(5423);
    layer3_outputs(7016) <= not(layer2_outputs(2748)) or (layer2_outputs(1256));
    layer3_outputs(7017) <= (layer2_outputs(6912)) xor (layer2_outputs(6050));
    layer3_outputs(7018) <= (layer2_outputs(6531)) and not (layer2_outputs(6381));
    layer3_outputs(7019) <= (layer2_outputs(1623)) or (layer2_outputs(5991));
    layer3_outputs(7020) <= not(layer2_outputs(5738));
    layer3_outputs(7021) <= not(layer2_outputs(738)) or (layer2_outputs(845));
    layer3_outputs(7022) <= (layer2_outputs(3117)) and not (layer2_outputs(7189));
    layer3_outputs(7023) <= not(layer2_outputs(9033));
    layer3_outputs(7024) <= layer2_outputs(1755);
    layer3_outputs(7025) <= (layer2_outputs(6288)) and (layer2_outputs(9460));
    layer3_outputs(7026) <= (layer2_outputs(4564)) and not (layer2_outputs(1519));
    layer3_outputs(7027) <= layer2_outputs(8434);
    layer3_outputs(7028) <= layer2_outputs(3236);
    layer3_outputs(7029) <= not(layer2_outputs(4856));
    layer3_outputs(7030) <= layer2_outputs(2456);
    layer3_outputs(7031) <= (layer2_outputs(5034)) and (layer2_outputs(3907));
    layer3_outputs(7032) <= not(layer2_outputs(9567));
    layer3_outputs(7033) <= layer2_outputs(7328);
    layer3_outputs(7034) <= not(layer2_outputs(1698));
    layer3_outputs(7035) <= (layer2_outputs(3629)) or (layer2_outputs(8959));
    layer3_outputs(7036) <= not(layer2_outputs(7717));
    layer3_outputs(7037) <= not((layer2_outputs(9667)) or (layer2_outputs(2688)));
    layer3_outputs(7038) <= layer2_outputs(7228);
    layer3_outputs(7039) <= (layer2_outputs(5004)) and not (layer2_outputs(3969));
    layer3_outputs(7040) <= not(layer2_outputs(5638)) or (layer2_outputs(167));
    layer3_outputs(7041) <= '1';
    layer3_outputs(7042) <= not(layer2_outputs(6745));
    layer3_outputs(7043) <= layer2_outputs(9685);
    layer3_outputs(7044) <= layer2_outputs(6021);
    layer3_outputs(7045) <= layer2_outputs(2636);
    layer3_outputs(7046) <= layer2_outputs(3684);
    layer3_outputs(7047) <= (layer2_outputs(10128)) and not (layer2_outputs(5474));
    layer3_outputs(7048) <= not(layer2_outputs(3660));
    layer3_outputs(7049) <= layer2_outputs(3536);
    layer3_outputs(7050) <= layer2_outputs(9630);
    layer3_outputs(7051) <= not(layer2_outputs(251));
    layer3_outputs(7052) <= (layer2_outputs(7813)) xor (layer2_outputs(3214));
    layer3_outputs(7053) <= layer2_outputs(1223);
    layer3_outputs(7054) <= layer2_outputs(1993);
    layer3_outputs(7055) <= layer2_outputs(778);
    layer3_outputs(7056) <= layer2_outputs(845);
    layer3_outputs(7057) <= not(layer2_outputs(3896));
    layer3_outputs(7058) <= not(layer2_outputs(8691));
    layer3_outputs(7059) <= not((layer2_outputs(3208)) or (layer2_outputs(8834)));
    layer3_outputs(7060) <= '1';
    layer3_outputs(7061) <= not((layer2_outputs(8076)) or (layer2_outputs(9404)));
    layer3_outputs(7062) <= not(layer2_outputs(5087));
    layer3_outputs(7063) <= not(layer2_outputs(1913)) or (layer2_outputs(2836));
    layer3_outputs(7064) <= not(layer2_outputs(5554));
    layer3_outputs(7065) <= not(layer2_outputs(7253));
    layer3_outputs(7066) <= layer2_outputs(1451);
    layer3_outputs(7067) <= (layer2_outputs(6253)) or (layer2_outputs(8143));
    layer3_outputs(7068) <= not((layer2_outputs(10041)) or (layer2_outputs(10126)));
    layer3_outputs(7069) <= (layer2_outputs(2087)) xor (layer2_outputs(2469));
    layer3_outputs(7070) <= (layer2_outputs(8011)) and not (layer2_outputs(7581));
    layer3_outputs(7071) <= not((layer2_outputs(1068)) or (layer2_outputs(8282)));
    layer3_outputs(7072) <= not((layer2_outputs(9126)) or (layer2_outputs(1724)));
    layer3_outputs(7073) <= not((layer2_outputs(959)) or (layer2_outputs(1522)));
    layer3_outputs(7074) <= (layer2_outputs(5130)) or (layer2_outputs(3710));
    layer3_outputs(7075) <= layer2_outputs(7352);
    layer3_outputs(7076) <= not(layer2_outputs(8806));
    layer3_outputs(7077) <= not(layer2_outputs(4235));
    layer3_outputs(7078) <= (layer2_outputs(7366)) and (layer2_outputs(6762));
    layer3_outputs(7079) <= (layer2_outputs(1446)) and not (layer2_outputs(3609));
    layer3_outputs(7080) <= layer2_outputs(3235);
    layer3_outputs(7081) <= (layer2_outputs(8414)) or (layer2_outputs(4080));
    layer3_outputs(7082) <= '0';
    layer3_outputs(7083) <= (layer2_outputs(6438)) or (layer2_outputs(9145));
    layer3_outputs(7084) <= not((layer2_outputs(9620)) and (layer2_outputs(7993)));
    layer3_outputs(7085) <= not(layer2_outputs(235)) or (layer2_outputs(572));
    layer3_outputs(7086) <= (layer2_outputs(6443)) xor (layer2_outputs(8760));
    layer3_outputs(7087) <= not((layer2_outputs(3233)) and (layer2_outputs(9040)));
    layer3_outputs(7088) <= not((layer2_outputs(3013)) xor (layer2_outputs(7242)));
    layer3_outputs(7089) <= not((layer2_outputs(2255)) or (layer2_outputs(6057)));
    layer3_outputs(7090) <= not(layer2_outputs(6629));
    layer3_outputs(7091) <= not(layer2_outputs(864));
    layer3_outputs(7092) <= not(layer2_outputs(8781));
    layer3_outputs(7093) <= not(layer2_outputs(9104));
    layer3_outputs(7094) <= not(layer2_outputs(7388)) or (layer2_outputs(9545));
    layer3_outputs(7095) <= layer2_outputs(564);
    layer3_outputs(7096) <= not(layer2_outputs(404));
    layer3_outputs(7097) <= not((layer2_outputs(3087)) or (layer2_outputs(3837)));
    layer3_outputs(7098) <= not((layer2_outputs(2358)) xor (layer2_outputs(1722)));
    layer3_outputs(7099) <= (layer2_outputs(3803)) and not (layer2_outputs(4921));
    layer3_outputs(7100) <= not(layer2_outputs(2350));
    layer3_outputs(7101) <= not((layer2_outputs(5515)) xor (layer2_outputs(4316)));
    layer3_outputs(7102) <= not((layer2_outputs(4773)) and (layer2_outputs(9279)));
    layer3_outputs(7103) <= (layer2_outputs(4445)) and not (layer2_outputs(3388));
    layer3_outputs(7104) <= not((layer2_outputs(8657)) or (layer2_outputs(9390)));
    layer3_outputs(7105) <= (layer2_outputs(4551)) and (layer2_outputs(8958));
    layer3_outputs(7106) <= not(layer2_outputs(2916));
    layer3_outputs(7107) <= not((layer2_outputs(7950)) and (layer2_outputs(7101)));
    layer3_outputs(7108) <= not(layer2_outputs(6009));
    layer3_outputs(7109) <= (layer2_outputs(8063)) and (layer2_outputs(7785));
    layer3_outputs(7110) <= not((layer2_outputs(8315)) xor (layer2_outputs(275)));
    layer3_outputs(7111) <= not(layer2_outputs(8742));
    layer3_outputs(7112) <= not(layer2_outputs(3433));
    layer3_outputs(7113) <= (layer2_outputs(4149)) xor (layer2_outputs(532));
    layer3_outputs(7114) <= (layer2_outputs(3262)) and not (layer2_outputs(6661));
    layer3_outputs(7115) <= layer2_outputs(5669);
    layer3_outputs(7116) <= (layer2_outputs(4260)) xor (layer2_outputs(1637));
    layer3_outputs(7117) <= not(layer2_outputs(6523));
    layer3_outputs(7118) <= not(layer2_outputs(4380));
    layer3_outputs(7119) <= not(layer2_outputs(1517));
    layer3_outputs(7120) <= layer2_outputs(1911);
    layer3_outputs(7121) <= (layer2_outputs(10165)) or (layer2_outputs(854));
    layer3_outputs(7122) <= (layer2_outputs(1259)) or (layer2_outputs(6526));
    layer3_outputs(7123) <= not(layer2_outputs(2385));
    layer3_outputs(7124) <= not((layer2_outputs(5348)) or (layer2_outputs(1928)));
    layer3_outputs(7125) <= not(layer2_outputs(8355));
    layer3_outputs(7126) <= not(layer2_outputs(9539));
    layer3_outputs(7127) <= not(layer2_outputs(9660));
    layer3_outputs(7128) <= not(layer2_outputs(1433)) or (layer2_outputs(3077));
    layer3_outputs(7129) <= not((layer2_outputs(3333)) or (layer2_outputs(4482)));
    layer3_outputs(7130) <= not(layer2_outputs(8807));
    layer3_outputs(7131) <= not(layer2_outputs(2662));
    layer3_outputs(7132) <= not(layer2_outputs(2627));
    layer3_outputs(7133) <= not(layer2_outputs(9179));
    layer3_outputs(7134) <= layer2_outputs(2734);
    layer3_outputs(7135) <= layer2_outputs(7578);
    layer3_outputs(7136) <= not(layer2_outputs(3915));
    layer3_outputs(7137) <= not((layer2_outputs(1783)) or (layer2_outputs(234)));
    layer3_outputs(7138) <= not(layer2_outputs(9142));
    layer3_outputs(7139) <= '1';
    layer3_outputs(7140) <= not((layer2_outputs(11)) or (layer2_outputs(371)));
    layer3_outputs(7141) <= (layer2_outputs(1543)) xor (layer2_outputs(2461));
    layer3_outputs(7142) <= layer2_outputs(9390);
    layer3_outputs(7143) <= (layer2_outputs(8748)) or (layer2_outputs(1485));
    layer3_outputs(7144) <= not(layer2_outputs(3592));
    layer3_outputs(7145) <= (layer2_outputs(880)) and not (layer2_outputs(5683));
    layer3_outputs(7146) <= (layer2_outputs(357)) and not (layer2_outputs(4853));
    layer3_outputs(7147) <= (layer2_outputs(7264)) or (layer2_outputs(2029));
    layer3_outputs(7148) <= not(layer2_outputs(9079));
    layer3_outputs(7149) <= layer2_outputs(2928);
    layer3_outputs(7150) <= not(layer2_outputs(6852));
    layer3_outputs(7151) <= not(layer2_outputs(5451));
    layer3_outputs(7152) <= layer2_outputs(1982);
    layer3_outputs(7153) <= not(layer2_outputs(2969));
    layer3_outputs(7154) <= not(layer2_outputs(2603));
    layer3_outputs(7155) <= layer2_outputs(9593);
    layer3_outputs(7156) <= (layer2_outputs(3718)) and (layer2_outputs(8524));
    layer3_outputs(7157) <= not(layer2_outputs(629));
    layer3_outputs(7158) <= (layer2_outputs(1660)) and not (layer2_outputs(7167));
    layer3_outputs(7159) <= layer2_outputs(2999);
    layer3_outputs(7160) <= not(layer2_outputs(1030)) or (layer2_outputs(7780));
    layer3_outputs(7161) <= (layer2_outputs(5058)) xor (layer2_outputs(8692));
    layer3_outputs(7162) <= (layer2_outputs(8115)) and (layer2_outputs(749));
    layer3_outputs(7163) <= layer2_outputs(7845);
    layer3_outputs(7164) <= (layer2_outputs(2894)) and (layer2_outputs(7240));
    layer3_outputs(7165) <= layer2_outputs(492);
    layer3_outputs(7166) <= not(layer2_outputs(7983)) or (layer2_outputs(7416));
    layer3_outputs(7167) <= (layer2_outputs(392)) or (layer2_outputs(1239));
    layer3_outputs(7168) <= not(layer2_outputs(7243)) or (layer2_outputs(3977));
    layer3_outputs(7169) <= (layer2_outputs(4614)) or (layer2_outputs(8625));
    layer3_outputs(7170) <= not(layer2_outputs(4339));
    layer3_outputs(7171) <= (layer2_outputs(9484)) and not (layer2_outputs(4390));
    layer3_outputs(7172) <= not(layer2_outputs(8106));
    layer3_outputs(7173) <= (layer2_outputs(6986)) and (layer2_outputs(1194));
    layer3_outputs(7174) <= layer2_outputs(7850);
    layer3_outputs(7175) <= (layer2_outputs(7266)) or (layer2_outputs(3420));
    layer3_outputs(7176) <= layer2_outputs(1324);
    layer3_outputs(7177) <= (layer2_outputs(7129)) and not (layer2_outputs(6110));
    layer3_outputs(7178) <= not(layer2_outputs(525));
    layer3_outputs(7179) <= (layer2_outputs(6895)) or (layer2_outputs(6862));
    layer3_outputs(7180) <= (layer2_outputs(5008)) and not (layer2_outputs(9200));
    layer3_outputs(7181) <= not(layer2_outputs(3744));
    layer3_outputs(7182) <= not(layer2_outputs(10171));
    layer3_outputs(7183) <= (layer2_outputs(10219)) or (layer2_outputs(3448));
    layer3_outputs(7184) <= not(layer2_outputs(6648));
    layer3_outputs(7185) <= not(layer2_outputs(7969)) or (layer2_outputs(3474));
    layer3_outputs(7186) <= not((layer2_outputs(800)) or (layer2_outputs(1380)));
    layer3_outputs(7187) <= not(layer2_outputs(4466));
    layer3_outputs(7188) <= not(layer2_outputs(4729));
    layer3_outputs(7189) <= layer2_outputs(3451);
    layer3_outputs(7190) <= not(layer2_outputs(5239));
    layer3_outputs(7191) <= not(layer2_outputs(8786));
    layer3_outputs(7192) <= (layer2_outputs(3740)) and not (layer2_outputs(5624));
    layer3_outputs(7193) <= (layer2_outputs(2820)) or (layer2_outputs(1948));
    layer3_outputs(7194) <= not(layer2_outputs(5064));
    layer3_outputs(7195) <= not((layer2_outputs(9326)) xor (layer2_outputs(8342)));
    layer3_outputs(7196) <= not(layer2_outputs(774));
    layer3_outputs(7197) <= (layer2_outputs(7430)) and not (layer2_outputs(3327));
    layer3_outputs(7198) <= not(layer2_outputs(5273));
    layer3_outputs(7199) <= (layer2_outputs(8867)) or (layer2_outputs(2159));
    layer3_outputs(7200) <= not(layer2_outputs(743));
    layer3_outputs(7201) <= (layer2_outputs(8439)) and (layer2_outputs(1562));
    layer3_outputs(7202) <= layer2_outputs(3185);
    layer3_outputs(7203) <= not(layer2_outputs(3071));
    layer3_outputs(7204) <= (layer2_outputs(8939)) and not (layer2_outputs(4409));
    layer3_outputs(7205) <= (layer2_outputs(6066)) xor (layer2_outputs(2340));
    layer3_outputs(7206) <= not((layer2_outputs(7970)) and (layer2_outputs(5284)));
    layer3_outputs(7207) <= not(layer2_outputs(6901));
    layer3_outputs(7208) <= layer2_outputs(7595);
    layer3_outputs(7209) <= layer2_outputs(4899);
    layer3_outputs(7210) <= not(layer2_outputs(2450));
    layer3_outputs(7211) <= layer2_outputs(6783);
    layer3_outputs(7212) <= (layer2_outputs(9201)) xor (layer2_outputs(7712));
    layer3_outputs(7213) <= not(layer2_outputs(8881));
    layer3_outputs(7214) <= (layer2_outputs(318)) xor (layer2_outputs(3995));
    layer3_outputs(7215) <= not(layer2_outputs(3030));
    layer3_outputs(7216) <= not((layer2_outputs(3114)) or (layer2_outputs(2917)));
    layer3_outputs(7217) <= '1';
    layer3_outputs(7218) <= layer2_outputs(7143);
    layer3_outputs(7219) <= not((layer2_outputs(1356)) or (layer2_outputs(9402)));
    layer3_outputs(7220) <= layer2_outputs(7554);
    layer3_outputs(7221) <= not((layer2_outputs(4914)) xor (layer2_outputs(965)));
    layer3_outputs(7222) <= (layer2_outputs(416)) and (layer2_outputs(5855));
    layer3_outputs(7223) <= not((layer2_outputs(9913)) and (layer2_outputs(5262)));
    layer3_outputs(7224) <= not(layer2_outputs(2234));
    layer3_outputs(7225) <= layer2_outputs(6065);
    layer3_outputs(7226) <= layer2_outputs(4298);
    layer3_outputs(7227) <= not(layer2_outputs(2066)) or (layer2_outputs(7993));
    layer3_outputs(7228) <= layer2_outputs(2877);
    layer3_outputs(7229) <= layer2_outputs(3783);
    layer3_outputs(7230) <= layer2_outputs(3559);
    layer3_outputs(7231) <= not(layer2_outputs(3372));
    layer3_outputs(7232) <= not(layer2_outputs(6044));
    layer3_outputs(7233) <= not((layer2_outputs(1815)) or (layer2_outputs(418)));
    layer3_outputs(7234) <= (layer2_outputs(4262)) or (layer2_outputs(6920));
    layer3_outputs(7235) <= not(layer2_outputs(8651));
    layer3_outputs(7236) <= layer2_outputs(2483);
    layer3_outputs(7237) <= layer2_outputs(4353);
    layer3_outputs(7238) <= not(layer2_outputs(7852));
    layer3_outputs(7239) <= (layer2_outputs(2083)) or (layer2_outputs(6822));
    layer3_outputs(7240) <= not((layer2_outputs(3918)) or (layer2_outputs(4031)));
    layer3_outputs(7241) <= not(layer2_outputs(6011)) or (layer2_outputs(1055));
    layer3_outputs(7242) <= (layer2_outputs(52)) xor (layer2_outputs(2190));
    layer3_outputs(7243) <= layer2_outputs(3872);
    layer3_outputs(7244) <= (layer2_outputs(7823)) xor (layer2_outputs(7084));
    layer3_outputs(7245) <= (layer2_outputs(4307)) and not (layer2_outputs(4798));
    layer3_outputs(7246) <= not(layer2_outputs(982));
    layer3_outputs(7247) <= not((layer2_outputs(7654)) and (layer2_outputs(4000)));
    layer3_outputs(7248) <= layer2_outputs(3708);
    layer3_outputs(7249) <= '0';
    layer3_outputs(7250) <= not((layer2_outputs(9312)) or (layer2_outputs(1609)));
    layer3_outputs(7251) <= (layer2_outputs(9960)) xor (layer2_outputs(6197));
    layer3_outputs(7252) <= layer2_outputs(4704);
    layer3_outputs(7253) <= layer2_outputs(1353);
    layer3_outputs(7254) <= (layer2_outputs(1374)) and (layer2_outputs(5444));
    layer3_outputs(7255) <= (layer2_outputs(812)) and not (layer2_outputs(6602));
    layer3_outputs(7256) <= not(layer2_outputs(5429)) or (layer2_outputs(2471));
    layer3_outputs(7257) <= layer2_outputs(8016);
    layer3_outputs(7258) <= not(layer2_outputs(6892));
    layer3_outputs(7259) <= not(layer2_outputs(8804));
    layer3_outputs(7260) <= not(layer2_outputs(7224));
    layer3_outputs(7261) <= (layer2_outputs(4278)) and not (layer2_outputs(9064));
    layer3_outputs(7262) <= (layer2_outputs(5233)) and not (layer2_outputs(5846));
    layer3_outputs(7263) <= not(layer2_outputs(9606));
    layer3_outputs(7264) <= layer2_outputs(7864);
    layer3_outputs(7265) <= not(layer2_outputs(5202));
    layer3_outputs(7266) <= not(layer2_outputs(7259));
    layer3_outputs(7267) <= not((layer2_outputs(6185)) xor (layer2_outputs(6583)));
    layer3_outputs(7268) <= not(layer2_outputs(2635)) or (layer2_outputs(9614));
    layer3_outputs(7269) <= (layer2_outputs(1702)) xor (layer2_outputs(1154));
    layer3_outputs(7270) <= (layer2_outputs(3692)) and not (layer2_outputs(2106));
    layer3_outputs(7271) <= (layer2_outputs(6364)) or (layer2_outputs(8877));
    layer3_outputs(7272) <= layer2_outputs(8245);
    layer3_outputs(7273) <= layer2_outputs(6679);
    layer3_outputs(7274) <= layer2_outputs(8812);
    layer3_outputs(7275) <= not(layer2_outputs(4052));
    layer3_outputs(7276) <= (layer2_outputs(7521)) and (layer2_outputs(4812));
    layer3_outputs(7277) <= layer2_outputs(5600);
    layer3_outputs(7278) <= (layer2_outputs(10213)) or (layer2_outputs(3678));
    layer3_outputs(7279) <= (layer2_outputs(6967)) or (layer2_outputs(2898));
    layer3_outputs(7280) <= (layer2_outputs(2879)) xor (layer2_outputs(2095));
    layer3_outputs(7281) <= (layer2_outputs(4329)) and not (layer2_outputs(1587));
    layer3_outputs(7282) <= layer2_outputs(9501);
    layer3_outputs(7283) <= not(layer2_outputs(5232));
    layer3_outputs(7284) <= layer2_outputs(7820);
    layer3_outputs(7285) <= layer2_outputs(4028);
    layer3_outputs(7286) <= not(layer2_outputs(4036)) or (layer2_outputs(3001));
    layer3_outputs(7287) <= not(layer2_outputs(8924));
    layer3_outputs(7288) <= not((layer2_outputs(3791)) and (layer2_outputs(4095)));
    layer3_outputs(7289) <= (layer2_outputs(9957)) or (layer2_outputs(6728));
    layer3_outputs(7290) <= layer2_outputs(2023);
    layer3_outputs(7291) <= layer2_outputs(2659);
    layer3_outputs(7292) <= layer2_outputs(5922);
    layer3_outputs(7293) <= layer2_outputs(9208);
    layer3_outputs(7294) <= (layer2_outputs(5495)) and not (layer2_outputs(5912));
    layer3_outputs(7295) <= not(layer2_outputs(9896)) or (layer2_outputs(1630));
    layer3_outputs(7296) <= not(layer2_outputs(10177));
    layer3_outputs(7297) <= (layer2_outputs(5517)) and not (layer2_outputs(2494));
    layer3_outputs(7298) <= layer2_outputs(9591);
    layer3_outputs(7299) <= (layer2_outputs(7025)) and not (layer2_outputs(6663));
    layer3_outputs(7300) <= (layer2_outputs(8237)) and not (layer2_outputs(9082));
    layer3_outputs(7301) <= (layer2_outputs(4124)) and (layer2_outputs(4267));
    layer3_outputs(7302) <= layer2_outputs(8683);
    layer3_outputs(7303) <= not((layer2_outputs(9717)) or (layer2_outputs(5776)));
    layer3_outputs(7304) <= layer2_outputs(181);
    layer3_outputs(7305) <= layer2_outputs(3572);
    layer3_outputs(7306) <= not(layer2_outputs(402)) or (layer2_outputs(8414));
    layer3_outputs(7307) <= not((layer2_outputs(1114)) or (layer2_outputs(4605)));
    layer3_outputs(7308) <= layer2_outputs(1851);
    layer3_outputs(7309) <= not((layer2_outputs(3963)) xor (layer2_outputs(8762)));
    layer3_outputs(7310) <= layer2_outputs(3827);
    layer3_outputs(7311) <= layer2_outputs(9307);
    layer3_outputs(7312) <= not(layer2_outputs(4608)) or (layer2_outputs(5971));
    layer3_outputs(7313) <= (layer2_outputs(1670)) and not (layer2_outputs(4034));
    layer3_outputs(7314) <= not(layer2_outputs(9054));
    layer3_outputs(7315) <= not(layer2_outputs(7236));
    layer3_outputs(7316) <= not(layer2_outputs(2935));
    layer3_outputs(7317) <= '0';
    layer3_outputs(7318) <= not((layer2_outputs(3198)) or (layer2_outputs(399)));
    layer3_outputs(7319) <= not(layer2_outputs(1373));
    layer3_outputs(7320) <= not((layer2_outputs(8180)) and (layer2_outputs(4654)));
    layer3_outputs(7321) <= layer2_outputs(4600);
    layer3_outputs(7322) <= layer2_outputs(9673);
    layer3_outputs(7323) <= (layer2_outputs(3022)) or (layer2_outputs(347));
    layer3_outputs(7324) <= (layer2_outputs(9808)) and not (layer2_outputs(7875));
    layer3_outputs(7325) <= not(layer2_outputs(86));
    layer3_outputs(7326) <= (layer2_outputs(8122)) or (layer2_outputs(9938));
    layer3_outputs(7327) <= not(layer2_outputs(9901));
    layer3_outputs(7328) <= not(layer2_outputs(5880)) or (layer2_outputs(1723));
    layer3_outputs(7329) <= (layer2_outputs(5726)) and not (layer2_outputs(7162));
    layer3_outputs(7330) <= layer2_outputs(7030);
    layer3_outputs(7331) <= not(layer2_outputs(8814));
    layer3_outputs(7332) <= (layer2_outputs(8981)) and not (layer2_outputs(10145));
    layer3_outputs(7333) <= (layer2_outputs(3930)) and not (layer2_outputs(8559));
    layer3_outputs(7334) <= (layer2_outputs(1196)) and not (layer2_outputs(1969));
    layer3_outputs(7335) <= (layer2_outputs(9336)) and (layer2_outputs(98));
    layer3_outputs(7336) <= layer2_outputs(3478);
    layer3_outputs(7337) <= layer2_outputs(1584);
    layer3_outputs(7338) <= not(layer2_outputs(3353));
    layer3_outputs(7339) <= not(layer2_outputs(7901));
    layer3_outputs(7340) <= (layer2_outputs(5625)) and not (layer2_outputs(3707));
    layer3_outputs(7341) <= (layer2_outputs(5761)) and (layer2_outputs(4930));
    layer3_outputs(7342) <= not(layer2_outputs(6938));
    layer3_outputs(7343) <= not((layer2_outputs(5188)) and (layer2_outputs(5769)));
    layer3_outputs(7344) <= layer2_outputs(3981);
    layer3_outputs(7345) <= (layer2_outputs(9267)) xor (layer2_outputs(6808));
    layer3_outputs(7346) <= '1';
    layer3_outputs(7347) <= layer2_outputs(7200);
    layer3_outputs(7348) <= not((layer2_outputs(7495)) xor (layer2_outputs(6091)));
    layer3_outputs(7349) <= not(layer2_outputs(1870)) or (layer2_outputs(7977));
    layer3_outputs(7350) <= not(layer2_outputs(6699));
    layer3_outputs(7351) <= not((layer2_outputs(4772)) xor (layer2_outputs(3485)));
    layer3_outputs(7352) <= (layer2_outputs(766)) or (layer2_outputs(6853));
    layer3_outputs(7353) <= layer2_outputs(2910);
    layer3_outputs(7354) <= not(layer2_outputs(9555));
    layer3_outputs(7355) <= (layer2_outputs(6689)) and not (layer2_outputs(2975));
    layer3_outputs(7356) <= not((layer2_outputs(9685)) and (layer2_outputs(3967)));
    layer3_outputs(7357) <= (layer2_outputs(1281)) and not (layer2_outputs(5557));
    layer3_outputs(7358) <= not(layer2_outputs(1866)) or (layer2_outputs(5319));
    layer3_outputs(7359) <= not((layer2_outputs(267)) or (layer2_outputs(9055)));
    layer3_outputs(7360) <= not(layer2_outputs(10096));
    layer3_outputs(7361) <= not(layer2_outputs(3720));
    layer3_outputs(7362) <= layer2_outputs(5681);
    layer3_outputs(7363) <= (layer2_outputs(894)) xor (layer2_outputs(9918));
    layer3_outputs(7364) <= not(layer2_outputs(6959));
    layer3_outputs(7365) <= (layer2_outputs(9415)) and not (layer2_outputs(2477));
    layer3_outputs(7366) <= layer2_outputs(2973);
    layer3_outputs(7367) <= layer2_outputs(536);
    layer3_outputs(7368) <= not(layer2_outputs(1896));
    layer3_outputs(7369) <= not((layer2_outputs(4797)) or (layer2_outputs(9900)));
    layer3_outputs(7370) <= not(layer2_outputs(340));
    layer3_outputs(7371) <= layer2_outputs(4792);
    layer3_outputs(7372) <= (layer2_outputs(365)) and not (layer2_outputs(3156));
    layer3_outputs(7373) <= (layer2_outputs(325)) and not (layer2_outputs(6367));
    layer3_outputs(7374) <= not(layer2_outputs(8281)) or (layer2_outputs(284));
    layer3_outputs(7375) <= layer2_outputs(5921);
    layer3_outputs(7376) <= layer2_outputs(95);
    layer3_outputs(7377) <= not(layer2_outputs(4006));
    layer3_outputs(7378) <= not(layer2_outputs(259));
    layer3_outputs(7379) <= (layer2_outputs(2561)) and not (layer2_outputs(7435));
    layer3_outputs(7380) <= not((layer2_outputs(3471)) or (layer2_outputs(2023)));
    layer3_outputs(7381) <= (layer2_outputs(3399)) or (layer2_outputs(3561));
    layer3_outputs(7382) <= layer2_outputs(6559);
    layer3_outputs(7383) <= not(layer2_outputs(7536)) or (layer2_outputs(10075));
    layer3_outputs(7384) <= not((layer2_outputs(7945)) xor (layer2_outputs(7317)));
    layer3_outputs(7385) <= (layer2_outputs(8662)) and not (layer2_outputs(4419));
    layer3_outputs(7386) <= '1';
    layer3_outputs(7387) <= not((layer2_outputs(2327)) and (layer2_outputs(2326)));
    layer3_outputs(7388) <= not((layer2_outputs(7211)) xor (layer2_outputs(2328)));
    layer3_outputs(7389) <= not(layer2_outputs(817)) or (layer2_outputs(3887));
    layer3_outputs(7390) <= (layer2_outputs(8756)) and not (layer2_outputs(3088));
    layer3_outputs(7391) <= (layer2_outputs(9121)) and not (layer2_outputs(8965));
    layer3_outputs(7392) <= (layer2_outputs(5311)) or (layer2_outputs(5548));
    layer3_outputs(7393) <= (layer2_outputs(9890)) and (layer2_outputs(8042));
    layer3_outputs(7394) <= not(layer2_outputs(9951));
    layer3_outputs(7395) <= not(layer2_outputs(8921));
    layer3_outputs(7396) <= not((layer2_outputs(6511)) or (layer2_outputs(4307)));
    layer3_outputs(7397) <= not((layer2_outputs(10196)) xor (layer2_outputs(4417)));
    layer3_outputs(7398) <= layer2_outputs(8595);
    layer3_outputs(7399) <= '1';
    layer3_outputs(7400) <= (layer2_outputs(1286)) xor (layer2_outputs(3671));
    layer3_outputs(7401) <= not(layer2_outputs(2763));
    layer3_outputs(7402) <= layer2_outputs(7281);
    layer3_outputs(7403) <= layer2_outputs(3596);
    layer3_outputs(7404) <= not(layer2_outputs(5718)) or (layer2_outputs(5233));
    layer3_outputs(7405) <= not(layer2_outputs(8023)) or (layer2_outputs(2396));
    layer3_outputs(7406) <= not(layer2_outputs(7059));
    layer3_outputs(7407) <= layer2_outputs(1256);
    layer3_outputs(7408) <= layer2_outputs(259);
    layer3_outputs(7409) <= layer2_outputs(7645);
    layer3_outputs(7410) <= not(layer2_outputs(5800));
    layer3_outputs(7411) <= (layer2_outputs(2352)) or (layer2_outputs(7750));
    layer3_outputs(7412) <= (layer2_outputs(3956)) and not (layer2_outputs(2976));
    layer3_outputs(7413) <= not(layer2_outputs(771));
    layer3_outputs(7414) <= not((layer2_outputs(3526)) and (layer2_outputs(4568)));
    layer3_outputs(7415) <= not(layer2_outputs(10068)) or (layer2_outputs(2313));
    layer3_outputs(7416) <= layer2_outputs(4811);
    layer3_outputs(7417) <= (layer2_outputs(6315)) and (layer2_outputs(3394));
    layer3_outputs(7418) <= layer2_outputs(5259);
    layer3_outputs(7419) <= (layer2_outputs(5616)) and not (layer2_outputs(4526));
    layer3_outputs(7420) <= not(layer2_outputs(3936));
    layer3_outputs(7421) <= not(layer2_outputs(6395));
    layer3_outputs(7422) <= not(layer2_outputs(8884));
    layer3_outputs(7423) <= layer2_outputs(2751);
    layer3_outputs(7424) <= layer2_outputs(6264);
    layer3_outputs(7425) <= not(layer2_outputs(10099));
    layer3_outputs(7426) <= layer2_outputs(8526);
    layer3_outputs(7427) <= not(layer2_outputs(4969));
    layer3_outputs(7428) <= not((layer2_outputs(3286)) and (layer2_outputs(1439)));
    layer3_outputs(7429) <= (layer2_outputs(9746)) and not (layer2_outputs(3584));
    layer3_outputs(7430) <= (layer2_outputs(521)) or (layer2_outputs(8877));
    layer3_outputs(7431) <= layer2_outputs(6951);
    layer3_outputs(7432) <= (layer2_outputs(5035)) or (layer2_outputs(2132));
    layer3_outputs(7433) <= not(layer2_outputs(232));
    layer3_outputs(7434) <= not(layer2_outputs(1338));
    layer3_outputs(7435) <= (layer2_outputs(4954)) and not (layer2_outputs(6966));
    layer3_outputs(7436) <= layer2_outputs(7420);
    layer3_outputs(7437) <= (layer2_outputs(7845)) xor (layer2_outputs(4645));
    layer3_outputs(7438) <= not(layer2_outputs(8294));
    layer3_outputs(7439) <= layer2_outputs(9203);
    layer3_outputs(7440) <= layer2_outputs(6874);
    layer3_outputs(7441) <= layer2_outputs(182);
    layer3_outputs(7442) <= layer2_outputs(6708);
    layer3_outputs(7443) <= not(layer2_outputs(5133)) or (layer2_outputs(4043));
    layer3_outputs(7444) <= layer2_outputs(7497);
    layer3_outputs(7445) <= not(layer2_outputs(9954));
    layer3_outputs(7446) <= (layer2_outputs(5777)) and not (layer2_outputs(5646));
    layer3_outputs(7447) <= layer2_outputs(3091);
    layer3_outputs(7448) <= not(layer2_outputs(2271));
    layer3_outputs(7449) <= not(layer2_outputs(9259));
    layer3_outputs(7450) <= layer2_outputs(1943);
    layer3_outputs(7451) <= (layer2_outputs(5388)) and not (layer2_outputs(1979));
    layer3_outputs(7452) <= layer2_outputs(661);
    layer3_outputs(7453) <= (layer2_outputs(4329)) and not (layer2_outputs(6372));
    layer3_outputs(7454) <= (layer2_outputs(8705)) or (layer2_outputs(6196));
    layer3_outputs(7455) <= not(layer2_outputs(2201));
    layer3_outputs(7456) <= not(layer2_outputs(6409)) or (layer2_outputs(1885));
    layer3_outputs(7457) <= (layer2_outputs(3228)) and (layer2_outputs(5260));
    layer3_outputs(7458) <= layer2_outputs(3314);
    layer3_outputs(7459) <= (layer2_outputs(5968)) and not (layer2_outputs(1209));
    layer3_outputs(7460) <= (layer2_outputs(5977)) and (layer2_outputs(4724));
    layer3_outputs(7461) <= not(layer2_outputs(4893)) or (layer2_outputs(8398));
    layer3_outputs(7462) <= (layer2_outputs(5070)) or (layer2_outputs(2656));
    layer3_outputs(7463) <= not(layer2_outputs(2002));
    layer3_outputs(7464) <= (layer2_outputs(9066)) xor (layer2_outputs(10199));
    layer3_outputs(7465) <= not(layer2_outputs(6351));
    layer3_outputs(7466) <= not(layer2_outputs(4832));
    layer3_outputs(7467) <= not((layer2_outputs(1998)) or (layer2_outputs(12)));
    layer3_outputs(7468) <= not(layer2_outputs(4229));
    layer3_outputs(7469) <= layer2_outputs(2707);
    layer3_outputs(7470) <= (layer2_outputs(3373)) and not (layer2_outputs(5314));
    layer3_outputs(7471) <= (layer2_outputs(8409)) and not (layer2_outputs(79));
    layer3_outputs(7472) <= not(layer2_outputs(1176)) or (layer2_outputs(5457));
    layer3_outputs(7473) <= not((layer2_outputs(9306)) or (layer2_outputs(8354)));
    layer3_outputs(7474) <= (layer2_outputs(2924)) xor (layer2_outputs(2664));
    layer3_outputs(7475) <= not((layer2_outputs(3063)) xor (layer2_outputs(2635)));
    layer3_outputs(7476) <= not(layer2_outputs(2209));
    layer3_outputs(7477) <= not(layer2_outputs(2598));
    layer3_outputs(7478) <= not(layer2_outputs(8905));
    layer3_outputs(7479) <= (layer2_outputs(539)) and (layer2_outputs(3708));
    layer3_outputs(7480) <= not(layer2_outputs(9832));
    layer3_outputs(7481) <= not((layer2_outputs(4732)) xor (layer2_outputs(8131)));
    layer3_outputs(7482) <= (layer2_outputs(6228)) and not (layer2_outputs(3790));
    layer3_outputs(7483) <= (layer2_outputs(803)) xor (layer2_outputs(5609));
    layer3_outputs(7484) <= layer2_outputs(3299);
    layer3_outputs(7485) <= not(layer2_outputs(1816));
    layer3_outputs(7486) <= layer2_outputs(3745);
    layer3_outputs(7487) <= layer2_outputs(3492);
    layer3_outputs(7488) <= not(layer2_outputs(425));
    layer3_outputs(7489) <= not(layer2_outputs(2538));
    layer3_outputs(7490) <= not((layer2_outputs(8886)) xor (layer2_outputs(4229)));
    layer3_outputs(7491) <= not(layer2_outputs(1267));
    layer3_outputs(7492) <= (layer2_outputs(5704)) or (layer2_outputs(2673));
    layer3_outputs(7493) <= not((layer2_outputs(4351)) xor (layer2_outputs(1357)));
    layer3_outputs(7494) <= not(layer2_outputs(4291));
    layer3_outputs(7495) <= (layer2_outputs(2258)) and (layer2_outputs(5394));
    layer3_outputs(7496) <= '1';
    layer3_outputs(7497) <= not(layer2_outputs(2798)) or (layer2_outputs(8956));
    layer3_outputs(7498) <= '0';
    layer3_outputs(7499) <= not(layer2_outputs(903)) or (layer2_outputs(1254));
    layer3_outputs(7500) <= layer2_outputs(4467);
    layer3_outputs(7501) <= layer2_outputs(3957);
    layer3_outputs(7502) <= layer2_outputs(7643);
    layer3_outputs(7503) <= layer2_outputs(3315);
    layer3_outputs(7504) <= layer2_outputs(1732);
    layer3_outputs(7505) <= not(layer2_outputs(4007)) or (layer2_outputs(8322));
    layer3_outputs(7506) <= not((layer2_outputs(9961)) or (layer2_outputs(5479)));
    layer3_outputs(7507) <= not(layer2_outputs(4208));
    layer3_outputs(7508) <= layer2_outputs(9127);
    layer3_outputs(7509) <= not(layer2_outputs(102));
    layer3_outputs(7510) <= not((layer2_outputs(6331)) xor (layer2_outputs(2468)));
    layer3_outputs(7511) <= not(layer2_outputs(805));
    layer3_outputs(7512) <= not(layer2_outputs(5816));
    layer3_outputs(7513) <= not(layer2_outputs(2108));
    layer3_outputs(7514) <= not(layer2_outputs(1187));
    layer3_outputs(7515) <= not(layer2_outputs(10082));
    layer3_outputs(7516) <= (layer2_outputs(9026)) or (layer2_outputs(2729));
    layer3_outputs(7517) <= not(layer2_outputs(5642));
    layer3_outputs(7518) <= not(layer2_outputs(4550));
    layer3_outputs(7519) <= '0';
    layer3_outputs(7520) <= not((layer2_outputs(2926)) and (layer2_outputs(5482)));
    layer3_outputs(7521) <= not(layer2_outputs(9301));
    layer3_outputs(7522) <= '1';
    layer3_outputs(7523) <= not(layer2_outputs(1023)) or (layer2_outputs(265));
    layer3_outputs(7524) <= (layer2_outputs(1401)) xor (layer2_outputs(6399));
    layer3_outputs(7525) <= not((layer2_outputs(9972)) and (layer2_outputs(6188)));
    layer3_outputs(7526) <= not((layer2_outputs(6048)) or (layer2_outputs(2006)));
    layer3_outputs(7527) <= not(layer2_outputs(6389)) or (layer2_outputs(8685));
    layer3_outputs(7528) <= not((layer2_outputs(4305)) xor (layer2_outputs(553)));
    layer3_outputs(7529) <= not((layer2_outputs(4511)) or (layer2_outputs(2646)));
    layer3_outputs(7530) <= (layer2_outputs(2081)) or (layer2_outputs(8121));
    layer3_outputs(7531) <= layer2_outputs(4340);
    layer3_outputs(7532) <= not(layer2_outputs(4298)) or (layer2_outputs(1532));
    layer3_outputs(7533) <= layer2_outputs(3296);
    layer3_outputs(7534) <= (layer2_outputs(2699)) or (layer2_outputs(8643));
    layer3_outputs(7535) <= not(layer2_outputs(4858));
    layer3_outputs(7536) <= (layer2_outputs(6651)) xor (layer2_outputs(9183));
    layer3_outputs(7537) <= not(layer2_outputs(867));
    layer3_outputs(7538) <= layer2_outputs(7727);
    layer3_outputs(7539) <= layer2_outputs(144);
    layer3_outputs(7540) <= (layer2_outputs(993)) and not (layer2_outputs(2408));
    layer3_outputs(7541) <= layer2_outputs(4238);
    layer3_outputs(7542) <= layer2_outputs(9284);
    layer3_outputs(7543) <= layer2_outputs(7594);
    layer3_outputs(7544) <= not(layer2_outputs(7018));
    layer3_outputs(7545) <= layer2_outputs(6599);
    layer3_outputs(7546) <= not((layer2_outputs(9337)) or (layer2_outputs(7590)));
    layer3_outputs(7547) <= not(layer2_outputs(2594)) or (layer2_outputs(4354));
    layer3_outputs(7548) <= not(layer2_outputs(3868));
    layer3_outputs(7549) <= not(layer2_outputs(5697)) or (layer2_outputs(4477));
    layer3_outputs(7550) <= (layer2_outputs(3427)) xor (layer2_outputs(7795));
    layer3_outputs(7551) <= not((layer2_outputs(6526)) xor (layer2_outputs(6055)));
    layer3_outputs(7552) <= not(layer2_outputs(2507));
    layer3_outputs(7553) <= layer2_outputs(1491);
    layer3_outputs(7554) <= not(layer2_outputs(10118)) or (layer2_outputs(6312));
    layer3_outputs(7555) <= not(layer2_outputs(1776)) or (layer2_outputs(7623));
    layer3_outputs(7556) <= (layer2_outputs(8735)) and (layer2_outputs(1750));
    layer3_outputs(7557) <= '1';
    layer3_outputs(7558) <= layer2_outputs(7157);
    layer3_outputs(7559) <= layer2_outputs(4318);
    layer3_outputs(7560) <= layer2_outputs(8564);
    layer3_outputs(7561) <= not((layer2_outputs(3497)) xor (layer2_outputs(5978)));
    layer3_outputs(7562) <= layer2_outputs(847);
    layer3_outputs(7563) <= not(layer2_outputs(2320)) or (layer2_outputs(6383));
    layer3_outputs(7564) <= not(layer2_outputs(3504));
    layer3_outputs(7565) <= layer2_outputs(7142);
    layer3_outputs(7566) <= layer2_outputs(10007);
    layer3_outputs(7567) <= not(layer2_outputs(7676));
    layer3_outputs(7568) <= (layer2_outputs(9958)) and not (layer2_outputs(8337));
    layer3_outputs(7569) <= not(layer2_outputs(1621));
    layer3_outputs(7570) <= not(layer2_outputs(1534));
    layer3_outputs(7571) <= not(layer2_outputs(3628)) or (layer2_outputs(1148));
    layer3_outputs(7572) <= layer2_outputs(5738);
    layer3_outputs(7573) <= layer2_outputs(5558);
    layer3_outputs(7574) <= not(layer2_outputs(587)) or (layer2_outputs(4269));
    layer3_outputs(7575) <= layer2_outputs(5393);
    layer3_outputs(7576) <= layer2_outputs(6881);
    layer3_outputs(7577) <= layer2_outputs(7057);
    layer3_outputs(7578) <= layer2_outputs(4879);
    layer3_outputs(7579) <= layer2_outputs(726);
    layer3_outputs(7580) <= layer2_outputs(7004);
    layer3_outputs(7581) <= layer2_outputs(8849);
    layer3_outputs(7582) <= not(layer2_outputs(8152));
    layer3_outputs(7583) <= (layer2_outputs(6068)) and not (layer2_outputs(8320));
    layer3_outputs(7584) <= layer2_outputs(7628);
    layer3_outputs(7585) <= not(layer2_outputs(4776));
    layer3_outputs(7586) <= (layer2_outputs(2919)) or (layer2_outputs(4161));
    layer3_outputs(7587) <= layer2_outputs(8680);
    layer3_outputs(7588) <= not(layer2_outputs(8804));
    layer3_outputs(7589) <= not((layer2_outputs(4014)) and (layer2_outputs(2633)));
    layer3_outputs(7590) <= (layer2_outputs(4597)) or (layer2_outputs(6157));
    layer3_outputs(7591) <= not(layer2_outputs(2028));
    layer3_outputs(7592) <= (layer2_outputs(643)) xor (layer2_outputs(8597));
    layer3_outputs(7593) <= layer2_outputs(7709);
    layer3_outputs(7594) <= '0';
    layer3_outputs(7595) <= (layer2_outputs(151)) and not (layer2_outputs(3500));
    layer3_outputs(7596) <= not((layer2_outputs(1096)) or (layer2_outputs(4595)));
    layer3_outputs(7597) <= not((layer2_outputs(4718)) and (layer2_outputs(5199)));
    layer3_outputs(7598) <= layer2_outputs(8256);
    layer3_outputs(7599) <= not(layer2_outputs(1229));
    layer3_outputs(7600) <= not((layer2_outputs(3067)) or (layer2_outputs(2293)));
    layer3_outputs(7601) <= not(layer2_outputs(2324));
    layer3_outputs(7602) <= (layer2_outputs(1806)) and not (layer2_outputs(4552));
    layer3_outputs(7603) <= layer2_outputs(3089);
    layer3_outputs(7604) <= not((layer2_outputs(6982)) xor (layer2_outputs(463)));
    layer3_outputs(7605) <= not(layer2_outputs(7751));
    layer3_outputs(7606) <= not(layer2_outputs(2551));
    layer3_outputs(7607) <= layer2_outputs(7395);
    layer3_outputs(7608) <= not(layer2_outputs(9430));
    layer3_outputs(7609) <= not(layer2_outputs(9598));
    layer3_outputs(7610) <= layer2_outputs(5015);
    layer3_outputs(7611) <= layer2_outputs(5176);
    layer3_outputs(7612) <= not((layer2_outputs(8240)) or (layer2_outputs(438)));
    layer3_outputs(7613) <= layer2_outputs(2805);
    layer3_outputs(7614) <= not(layer2_outputs(5487)) or (layer2_outputs(803));
    layer3_outputs(7615) <= layer2_outputs(3496);
    layer3_outputs(7616) <= not((layer2_outputs(5678)) xor (layer2_outputs(7592)));
    layer3_outputs(7617) <= (layer2_outputs(7037)) and not (layer2_outputs(6714));
    layer3_outputs(7618) <= not(layer2_outputs(6555));
    layer3_outputs(7619) <= layer2_outputs(2410);
    layer3_outputs(7620) <= (layer2_outputs(5254)) and not (layer2_outputs(1947));
    layer3_outputs(7621) <= layer2_outputs(9867);
    layer3_outputs(7622) <= not(layer2_outputs(5470));
    layer3_outputs(7623) <= layer2_outputs(8060);
    layer3_outputs(7624) <= (layer2_outputs(3344)) and not (layer2_outputs(9436));
    layer3_outputs(7625) <= not((layer2_outputs(2018)) and (layer2_outputs(202)));
    layer3_outputs(7626) <= not((layer2_outputs(7301)) xor (layer2_outputs(1004)));
    layer3_outputs(7627) <= layer2_outputs(1265);
    layer3_outputs(7628) <= layer2_outputs(116);
    layer3_outputs(7629) <= not(layer2_outputs(310));
    layer3_outputs(7630) <= not(layer2_outputs(4107));
    layer3_outputs(7631) <= not(layer2_outputs(287)) or (layer2_outputs(1782));
    layer3_outputs(7632) <= '1';
    layer3_outputs(7633) <= layer2_outputs(7286);
    layer3_outputs(7634) <= (layer2_outputs(7364)) and not (layer2_outputs(7734));
    layer3_outputs(7635) <= (layer2_outputs(9561)) and not (layer2_outputs(4673));
    layer3_outputs(7636) <= layer2_outputs(8473);
    layer3_outputs(7637) <= (layer2_outputs(9385)) xor (layer2_outputs(8341));
    layer3_outputs(7638) <= layer2_outputs(5883);
    layer3_outputs(7639) <= layer2_outputs(6065);
    layer3_outputs(7640) <= not((layer2_outputs(7113)) or (layer2_outputs(4069)));
    layer3_outputs(7641) <= not(layer2_outputs(8643));
    layer3_outputs(7642) <= layer2_outputs(3254);
    layer3_outputs(7643) <= (layer2_outputs(8676)) xor (layer2_outputs(7109));
    layer3_outputs(7644) <= not(layer2_outputs(3324)) or (layer2_outputs(3505));
    layer3_outputs(7645) <= (layer2_outputs(5837)) and (layer2_outputs(3169));
    layer3_outputs(7646) <= (layer2_outputs(2794)) and (layer2_outputs(3399));
    layer3_outputs(7647) <= not((layer2_outputs(8292)) or (layer2_outputs(3819)));
    layer3_outputs(7648) <= '1';
    layer3_outputs(7649) <= not((layer2_outputs(1514)) and (layer2_outputs(2925)));
    layer3_outputs(7650) <= not((layer2_outputs(2682)) and (layer2_outputs(2553)));
    layer3_outputs(7651) <= (layer2_outputs(4305)) xor (layer2_outputs(5579));
    layer3_outputs(7652) <= layer2_outputs(1703);
    layer3_outputs(7653) <= not((layer2_outputs(8972)) and (layer2_outputs(5774)));
    layer3_outputs(7654) <= not((layer2_outputs(3046)) or (layer2_outputs(7979)));
    layer3_outputs(7655) <= (layer2_outputs(2979)) or (layer2_outputs(373));
    layer3_outputs(7656) <= not(layer2_outputs(829)) or (layer2_outputs(8027));
    layer3_outputs(7657) <= (layer2_outputs(5990)) and not (layer2_outputs(3384));
    layer3_outputs(7658) <= (layer2_outputs(8261)) and not (layer2_outputs(8957));
    layer3_outputs(7659) <= not(layer2_outputs(1729));
    layer3_outputs(7660) <= layer2_outputs(3633);
    layer3_outputs(7661) <= not(layer2_outputs(3033)) or (layer2_outputs(2159));
    layer3_outputs(7662) <= layer2_outputs(4985);
    layer3_outputs(7663) <= not(layer2_outputs(10056)) or (layer2_outputs(449));
    layer3_outputs(7664) <= not((layer2_outputs(9359)) xor (layer2_outputs(3131)));
    layer3_outputs(7665) <= (layer2_outputs(701)) xor (layer2_outputs(6078));
    layer3_outputs(7666) <= not(layer2_outputs(2107));
    layer3_outputs(7667) <= layer2_outputs(4048);
    layer3_outputs(7668) <= layer2_outputs(6475);
    layer3_outputs(7669) <= (layer2_outputs(2364)) and (layer2_outputs(2266));
    layer3_outputs(7670) <= '0';
    layer3_outputs(7671) <= (layer2_outputs(3979)) and not (layer2_outputs(8174));
    layer3_outputs(7672) <= not(layer2_outputs(10018)) or (layer2_outputs(3147));
    layer3_outputs(7673) <= not(layer2_outputs(7174));
    layer3_outputs(7674) <= layer2_outputs(9804);
    layer3_outputs(7675) <= not((layer2_outputs(4638)) and (layer2_outputs(8605)));
    layer3_outputs(7676) <= (layer2_outputs(101)) and not (layer2_outputs(2444));
    layer3_outputs(7677) <= layer2_outputs(5153);
    layer3_outputs(7678) <= layer2_outputs(6340);
    layer3_outputs(7679) <= not((layer2_outputs(4898)) xor (layer2_outputs(7302)));
    layer3_outputs(7680) <= (layer2_outputs(8894)) xor (layer2_outputs(6440));
    layer3_outputs(7681) <= not(layer2_outputs(6039));
    layer3_outputs(7682) <= layer2_outputs(9382);
    layer3_outputs(7683) <= not((layer2_outputs(2875)) or (layer2_outputs(359)));
    layer3_outputs(7684) <= not((layer2_outputs(5804)) or (layer2_outputs(7956)));
    layer3_outputs(7685) <= not(layer2_outputs(6462));
    layer3_outputs(7686) <= not(layer2_outputs(3066));
    layer3_outputs(7687) <= (layer2_outputs(9610)) and not (layer2_outputs(9764));
    layer3_outputs(7688) <= layer2_outputs(1689);
    layer3_outputs(7689) <= layer2_outputs(6132);
    layer3_outputs(7690) <= layer2_outputs(1893);
    layer3_outputs(7691) <= (layer2_outputs(1372)) xor (layer2_outputs(539));
    layer3_outputs(7692) <= (layer2_outputs(9906)) and not (layer2_outputs(5552));
    layer3_outputs(7693) <= (layer2_outputs(7673)) and not (layer2_outputs(8416));
    layer3_outputs(7694) <= layer2_outputs(5644);
    layer3_outputs(7695) <= not((layer2_outputs(5508)) or (layer2_outputs(1158)));
    layer3_outputs(7696) <= (layer2_outputs(1366)) and not (layer2_outputs(5881));
    layer3_outputs(7697) <= layer2_outputs(2655);
    layer3_outputs(7698) <= not(layer2_outputs(9444));
    layer3_outputs(7699) <= '1';
    layer3_outputs(7700) <= not(layer2_outputs(5378));
    layer3_outputs(7701) <= not(layer2_outputs(3976));
    layer3_outputs(7702) <= (layer2_outputs(6085)) and not (layer2_outputs(9833));
    layer3_outputs(7703) <= not(layer2_outputs(5987));
    layer3_outputs(7704) <= not(layer2_outputs(7039));
    layer3_outputs(7705) <= layer2_outputs(2144);
    layer3_outputs(7706) <= layer2_outputs(1675);
    layer3_outputs(7707) <= not(layer2_outputs(1583));
    layer3_outputs(7708) <= not(layer2_outputs(3363));
    layer3_outputs(7709) <= (layer2_outputs(2476)) xor (layer2_outputs(2052));
    layer3_outputs(7710) <= layer2_outputs(5419);
    layer3_outputs(7711) <= layer2_outputs(4754);
    layer3_outputs(7712) <= (layer2_outputs(8987)) and not (layer2_outputs(3828));
    layer3_outputs(7713) <= (layer2_outputs(9970)) and not (layer2_outputs(4103));
    layer3_outputs(7714) <= '0';
    layer3_outputs(7715) <= (layer2_outputs(10098)) and (layer2_outputs(5045));
    layer3_outputs(7716) <= not(layer2_outputs(4786));
    layer3_outputs(7717) <= layer2_outputs(5949);
    layer3_outputs(7718) <= (layer2_outputs(2454)) and not (layer2_outputs(3857));
    layer3_outputs(7719) <= not((layer2_outputs(4389)) and (layer2_outputs(1706)));
    layer3_outputs(7720) <= (layer2_outputs(2165)) and (layer2_outputs(2840));
    layer3_outputs(7721) <= layer2_outputs(4027);
    layer3_outputs(7722) <= not(layer2_outputs(6929));
    layer3_outputs(7723) <= not((layer2_outputs(843)) or (layer2_outputs(8462)));
    layer3_outputs(7724) <= not(layer2_outputs(3529));
    layer3_outputs(7725) <= not(layer2_outputs(1903)) or (layer2_outputs(4970));
    layer3_outputs(7726) <= layer2_outputs(4818);
    layer3_outputs(7727) <= layer2_outputs(909);
    layer3_outputs(7728) <= not((layer2_outputs(501)) or (layer2_outputs(10155)));
    layer3_outputs(7729) <= not(layer2_outputs(7865));
    layer3_outputs(7730) <= (layer2_outputs(5612)) and not (layer2_outputs(534));
    layer3_outputs(7731) <= (layer2_outputs(1766)) and (layer2_outputs(5201));
    layer3_outputs(7732) <= not(layer2_outputs(552));
    layer3_outputs(7733) <= '1';
    layer3_outputs(7734) <= not(layer2_outputs(4390));
    layer3_outputs(7735) <= not((layer2_outputs(9077)) xor (layer2_outputs(71)));
    layer3_outputs(7736) <= (layer2_outputs(2821)) and not (layer2_outputs(9246));
    layer3_outputs(7737) <= not(layer2_outputs(7061)) or (layer2_outputs(5705));
    layer3_outputs(7738) <= not(layer2_outputs(4434)) or (layer2_outputs(4992));
    layer3_outputs(7739) <= layer2_outputs(6748);
    layer3_outputs(7740) <= layer2_outputs(8800);
    layer3_outputs(7741) <= not(layer2_outputs(3483)) or (layer2_outputs(6883));
    layer3_outputs(7742) <= (layer2_outputs(2550)) and not (layer2_outputs(8040));
    layer3_outputs(7743) <= layer2_outputs(6151);
    layer3_outputs(7744) <= not(layer2_outputs(463)) or (layer2_outputs(4569));
    layer3_outputs(7745) <= (layer2_outputs(8445)) and not (layer2_outputs(9379));
    layer3_outputs(7746) <= '0';
    layer3_outputs(7747) <= layer2_outputs(321);
    layer3_outputs(7748) <= not(layer2_outputs(937));
    layer3_outputs(7749) <= not(layer2_outputs(3651));
    layer3_outputs(7750) <= (layer2_outputs(6008)) or (layer2_outputs(9010));
    layer3_outputs(7751) <= not(layer2_outputs(6612));
    layer3_outputs(7752) <= (layer2_outputs(7539)) and not (layer2_outputs(1482));
    layer3_outputs(7753) <= not(layer2_outputs(5026));
    layer3_outputs(7754) <= (layer2_outputs(2316)) and not (layer2_outputs(1404));
    layer3_outputs(7755) <= not((layer2_outputs(9032)) and (layer2_outputs(8446)));
    layer3_outputs(7756) <= '0';
    layer3_outputs(7757) <= (layer2_outputs(530)) or (layer2_outputs(2300));
    layer3_outputs(7758) <= not(layer2_outputs(5418));
    layer3_outputs(7759) <= (layer2_outputs(2488)) and not (layer2_outputs(1230));
    layer3_outputs(7760) <= layer2_outputs(9708);
    layer3_outputs(7761) <= not(layer2_outputs(5043));
    layer3_outputs(7762) <= not((layer2_outputs(1725)) xor (layer2_outputs(9101)));
    layer3_outputs(7763) <= layer2_outputs(1174);
    layer3_outputs(7764) <= not(layer2_outputs(4627)) or (layer2_outputs(5496));
    layer3_outputs(7765) <= layer2_outputs(3522);
    layer3_outputs(7766) <= layer2_outputs(8603);
    layer3_outputs(7767) <= not((layer2_outputs(6811)) or (layer2_outputs(5291)));
    layer3_outputs(7768) <= layer2_outputs(3003);
    layer3_outputs(7769) <= layer2_outputs(1139);
    layer3_outputs(7770) <= (layer2_outputs(3430)) xor (layer2_outputs(3343));
    layer3_outputs(7771) <= not(layer2_outputs(7498)) or (layer2_outputs(6926));
    layer3_outputs(7772) <= layer2_outputs(3931);
    layer3_outputs(7773) <= not((layer2_outputs(1605)) or (layer2_outputs(8263)));
    layer3_outputs(7774) <= layer2_outputs(9027);
    layer3_outputs(7775) <= layer2_outputs(9096);
    layer3_outputs(7776) <= layer2_outputs(5949);
    layer3_outputs(7777) <= layer2_outputs(3169);
    layer3_outputs(7778) <= layer2_outputs(1627);
    layer3_outputs(7779) <= not((layer2_outputs(8146)) or (layer2_outputs(5652)));
    layer3_outputs(7780) <= (layer2_outputs(3427)) xor (layer2_outputs(9845));
    layer3_outputs(7781) <= not(layer2_outputs(308)) or (layer2_outputs(3278));
    layer3_outputs(7782) <= not(layer2_outputs(8386));
    layer3_outputs(7783) <= (layer2_outputs(9940)) or (layer2_outputs(2378));
    layer3_outputs(7784) <= layer2_outputs(25);
    layer3_outputs(7785) <= layer2_outputs(6386);
    layer3_outputs(7786) <= (layer2_outputs(6488)) xor (layer2_outputs(1530));
    layer3_outputs(7787) <= layer2_outputs(5214);
    layer3_outputs(7788) <= (layer2_outputs(3241)) and not (layer2_outputs(8087));
    layer3_outputs(7789) <= not((layer2_outputs(8732)) or (layer2_outputs(4502)));
    layer3_outputs(7790) <= layer2_outputs(4085);
    layer3_outputs(7791) <= layer2_outputs(5509);
    layer3_outputs(7792) <= not(layer2_outputs(3893));
    layer3_outputs(7793) <= (layer2_outputs(3956)) or (layer2_outputs(820));
    layer3_outputs(7794) <= not((layer2_outputs(1739)) and (layer2_outputs(1211)));
    layer3_outputs(7795) <= not(layer2_outputs(5167));
    layer3_outputs(7796) <= layer2_outputs(6750);
    layer3_outputs(7797) <= not((layer2_outputs(2951)) xor (layer2_outputs(8183)));
    layer3_outputs(7798) <= layer2_outputs(160);
    layer3_outputs(7799) <= not(layer2_outputs(7363));
    layer3_outputs(7800) <= (layer2_outputs(2838)) and not (layer2_outputs(3814));
    layer3_outputs(7801) <= not(layer2_outputs(2896));
    layer3_outputs(7802) <= layer2_outputs(9776);
    layer3_outputs(7803) <= not((layer2_outputs(3917)) or (layer2_outputs(4847)));
    layer3_outputs(7804) <= not(layer2_outputs(1269));
    layer3_outputs(7805) <= layer2_outputs(6156);
    layer3_outputs(7806) <= not(layer2_outputs(8141));
    layer3_outputs(7807) <= not((layer2_outputs(642)) or (layer2_outputs(8280)));
    layer3_outputs(7808) <= not((layer2_outputs(2347)) xor (layer2_outputs(7069)));
    layer3_outputs(7809) <= layer2_outputs(7379);
    layer3_outputs(7810) <= not((layer2_outputs(8901)) xor (layer2_outputs(3476)));
    layer3_outputs(7811) <= not((layer2_outputs(7711)) and (layer2_outputs(1302)));
    layer3_outputs(7812) <= layer2_outputs(4431);
    layer3_outputs(7813) <= not(layer2_outputs(3115));
    layer3_outputs(7814) <= '0';
    layer3_outputs(7815) <= not(layer2_outputs(876));
    layer3_outputs(7816) <= layer2_outputs(3235);
    layer3_outputs(7817) <= layer2_outputs(6220);
    layer3_outputs(7818) <= '1';
    layer3_outputs(7819) <= not(layer2_outputs(1223));
    layer3_outputs(7820) <= (layer2_outputs(2185)) and (layer2_outputs(6659));
    layer3_outputs(7821) <= (layer2_outputs(10008)) or (layer2_outputs(5397));
    layer3_outputs(7822) <= not((layer2_outputs(2265)) xor (layer2_outputs(5160)));
    layer3_outputs(7823) <= not(layer2_outputs(1319)) or (layer2_outputs(8829));
    layer3_outputs(7824) <= layer2_outputs(4341);
    layer3_outputs(7825) <= layer2_outputs(8554);
    layer3_outputs(7826) <= layer2_outputs(7907);
    layer3_outputs(7827) <= (layer2_outputs(8090)) xor (layer2_outputs(7719));
    layer3_outputs(7828) <= (layer2_outputs(901)) xor (layer2_outputs(5380));
    layer3_outputs(7829) <= (layer2_outputs(7469)) and not (layer2_outputs(6346));
    layer3_outputs(7830) <= not(layer2_outputs(2476));
    layer3_outputs(7831) <= not(layer2_outputs(5994));
    layer3_outputs(7832) <= not((layer2_outputs(4596)) or (layer2_outputs(7762)));
    layer3_outputs(7833) <= not(layer2_outputs(2972));
    layer3_outputs(7834) <= (layer2_outputs(846)) and not (layer2_outputs(3618));
    layer3_outputs(7835) <= layer2_outputs(1900);
    layer3_outputs(7836) <= (layer2_outputs(8024)) and not (layer2_outputs(459));
    layer3_outputs(7837) <= (layer2_outputs(3292)) or (layer2_outputs(9119));
    layer3_outputs(7838) <= not(layer2_outputs(9992));
    layer3_outputs(7839) <= '1';
    layer3_outputs(7840) <= (layer2_outputs(5919)) or (layer2_outputs(9877));
    layer3_outputs(7841) <= not(layer2_outputs(2449));
    layer3_outputs(7842) <= layer2_outputs(627);
    layer3_outputs(7843) <= not(layer2_outputs(9));
    layer3_outputs(7844) <= not(layer2_outputs(6296));
    layer3_outputs(7845) <= (layer2_outputs(4337)) and not (layer2_outputs(3845));
    layer3_outputs(7846) <= layer2_outputs(9381);
    layer3_outputs(7847) <= (layer2_outputs(2657)) and not (layer2_outputs(4084));
    layer3_outputs(7848) <= not(layer2_outputs(361));
    layer3_outputs(7849) <= not(layer2_outputs(6864));
    layer3_outputs(7850) <= (layer2_outputs(1435)) xor (layer2_outputs(6655));
    layer3_outputs(7851) <= layer2_outputs(7547);
    layer3_outputs(7852) <= layer2_outputs(3241);
    layer3_outputs(7853) <= not(layer2_outputs(81));
    layer3_outputs(7854) <= '1';
    layer3_outputs(7855) <= not((layer2_outputs(5617)) and (layer2_outputs(9754)));
    layer3_outputs(7856) <= not((layer2_outputs(6044)) xor (layer2_outputs(4294)));
    layer3_outputs(7857) <= not(layer2_outputs(723)) or (layer2_outputs(2557));
    layer3_outputs(7858) <= not(layer2_outputs(7124));
    layer3_outputs(7859) <= not(layer2_outputs(8192));
    layer3_outputs(7860) <= not(layer2_outputs(6415));
    layer3_outputs(7861) <= not(layer2_outputs(5849)) or (layer2_outputs(8917));
    layer3_outputs(7862) <= not(layer2_outputs(9328));
    layer3_outputs(7863) <= not((layer2_outputs(283)) or (layer2_outputs(6945)));
    layer3_outputs(7864) <= layer2_outputs(9796);
    layer3_outputs(7865) <= not(layer2_outputs(1079));
    layer3_outputs(7866) <= layer2_outputs(5598);
    layer3_outputs(7867) <= layer2_outputs(2230);
    layer3_outputs(7868) <= (layer2_outputs(8840)) xor (layer2_outputs(6796));
    layer3_outputs(7869) <= not((layer2_outputs(191)) and (layer2_outputs(3490)));
    layer3_outputs(7870) <= not(layer2_outputs(134));
    layer3_outputs(7871) <= (layer2_outputs(5705)) and (layer2_outputs(9106));
    layer3_outputs(7872) <= layer2_outputs(1867);
    layer3_outputs(7873) <= (layer2_outputs(1119)) and not (layer2_outputs(3202));
    layer3_outputs(7874) <= not(layer2_outputs(7110));
    layer3_outputs(7875) <= layer2_outputs(1062);
    layer3_outputs(7876) <= (layer2_outputs(2793)) and not (layer2_outputs(10030));
    layer3_outputs(7877) <= (layer2_outputs(8276)) xor (layer2_outputs(1833));
    layer3_outputs(7878) <= (layer2_outputs(8398)) and not (layer2_outputs(2510));
    layer3_outputs(7879) <= (layer2_outputs(10178)) xor (layer2_outputs(427));
    layer3_outputs(7880) <= not(layer2_outputs(1682)) or (layer2_outputs(7074));
    layer3_outputs(7881) <= not((layer2_outputs(1249)) or (layer2_outputs(4850)));
    layer3_outputs(7882) <= layer2_outputs(6541);
    layer3_outputs(7883) <= not(layer2_outputs(10225)) or (layer2_outputs(8116));
    layer3_outputs(7884) <= (layer2_outputs(351)) and not (layer2_outputs(8118));
    layer3_outputs(7885) <= (layer2_outputs(32)) and (layer2_outputs(8385));
    layer3_outputs(7886) <= (layer2_outputs(6424)) xor (layer2_outputs(4254));
    layer3_outputs(7887) <= not((layer2_outputs(5325)) and (layer2_outputs(4144)));
    layer3_outputs(7888) <= layer2_outputs(8683);
    layer3_outputs(7889) <= not((layer2_outputs(5751)) xor (layer2_outputs(9157)));
    layer3_outputs(7890) <= not(layer2_outputs(5431));
    layer3_outputs(7891) <= not(layer2_outputs(72));
    layer3_outputs(7892) <= not(layer2_outputs(2549));
    layer3_outputs(7893) <= not(layer2_outputs(3366)) or (layer2_outputs(6890));
    layer3_outputs(7894) <= (layer2_outputs(2631)) and not (layer2_outputs(3382));
    layer3_outputs(7895) <= (layer2_outputs(1127)) or (layer2_outputs(3962));
    layer3_outputs(7896) <= not(layer2_outputs(6912));
    layer3_outputs(7897) <= not((layer2_outputs(1809)) or (layer2_outputs(9094)));
    layer3_outputs(7898) <= (layer2_outputs(9355)) and not (layer2_outputs(1434));
    layer3_outputs(7899) <= layer2_outputs(10009);
    layer3_outputs(7900) <= not((layer2_outputs(1778)) or (layer2_outputs(1429)));
    layer3_outputs(7901) <= layer2_outputs(7293);
    layer3_outputs(7902) <= not(layer2_outputs(10029));
    layer3_outputs(7903) <= layer2_outputs(6884);
    layer3_outputs(7904) <= '1';
    layer3_outputs(7905) <= layer2_outputs(666);
    layer3_outputs(7906) <= (layer2_outputs(9018)) or (layer2_outputs(6687));
    layer3_outputs(7907) <= (layer2_outputs(5498)) and (layer2_outputs(4738));
    layer3_outputs(7908) <= not((layer2_outputs(1762)) or (layer2_outputs(947)));
    layer3_outputs(7909) <= layer2_outputs(787);
    layer3_outputs(7910) <= layer2_outputs(7605);
    layer3_outputs(7911) <= not(layer2_outputs(3989));
    layer3_outputs(7912) <= (layer2_outputs(6621)) and (layer2_outputs(9952));
    layer3_outputs(7913) <= layer2_outputs(6717);
    layer3_outputs(7914) <= layer2_outputs(2795);
    layer3_outputs(7915) <= layer2_outputs(9151);
    layer3_outputs(7916) <= (layer2_outputs(9915)) and not (layer2_outputs(345));
    layer3_outputs(7917) <= (layer2_outputs(2242)) and not (layer2_outputs(8576));
    layer3_outputs(7918) <= not((layer2_outputs(7235)) xor (layer2_outputs(9040)));
    layer3_outputs(7919) <= not(layer2_outputs(7450));
    layer3_outputs(7920) <= (layer2_outputs(3908)) xor (layer2_outputs(9791));
    layer3_outputs(7921) <= not((layer2_outputs(8407)) and (layer2_outputs(2732)));
    layer3_outputs(7922) <= (layer2_outputs(5333)) and not (layer2_outputs(1610));
    layer3_outputs(7923) <= layer2_outputs(8266);
    layer3_outputs(7924) <= layer2_outputs(3757);
    layer3_outputs(7925) <= '1';
    layer3_outputs(7926) <= (layer2_outputs(7038)) and not (layer2_outputs(6890));
    layer3_outputs(7927) <= layer2_outputs(5492);
    layer3_outputs(7928) <= not(layer2_outputs(6452)) or (layer2_outputs(8557));
    layer3_outputs(7929) <= layer2_outputs(3652);
    layer3_outputs(7930) <= '1';
    layer3_outputs(7931) <= layer2_outputs(8774);
    layer3_outputs(7932) <= layer2_outputs(363);
    layer3_outputs(7933) <= (layer2_outputs(7118)) and not (layer2_outputs(10093));
    layer3_outputs(7934) <= (layer2_outputs(4731)) and not (layer2_outputs(3792));
    layer3_outputs(7935) <= layer2_outputs(7515);
    layer3_outputs(7936) <= not(layer2_outputs(4386)) or (layer2_outputs(9399));
    layer3_outputs(7937) <= not((layer2_outputs(178)) and (layer2_outputs(8000)));
    layer3_outputs(7938) <= not(layer2_outputs(9250));
    layer3_outputs(7939) <= not((layer2_outputs(5816)) or (layer2_outputs(4406)));
    layer3_outputs(7940) <= (layer2_outputs(1289)) or (layer2_outputs(6152));
    layer3_outputs(7941) <= not((layer2_outputs(4803)) or (layer2_outputs(4753)));
    layer3_outputs(7942) <= not(layer2_outputs(3986));
    layer3_outputs(7943) <= (layer2_outputs(5782)) and not (layer2_outputs(2349));
    layer3_outputs(7944) <= not(layer2_outputs(9030)) or (layer2_outputs(808));
    layer3_outputs(7945) <= layer2_outputs(7757);
    layer3_outputs(7946) <= layer2_outputs(9681);
    layer3_outputs(7947) <= layer2_outputs(394);
    layer3_outputs(7948) <= not(layer2_outputs(2510));
    layer3_outputs(7949) <= (layer2_outputs(6450)) xor (layer2_outputs(8275));
    layer3_outputs(7950) <= layer2_outputs(7474);
    layer3_outputs(7951) <= not(layer2_outputs(2134));
    layer3_outputs(7952) <= not(layer2_outputs(2435)) or (layer2_outputs(176));
    layer3_outputs(7953) <= layer2_outputs(9421);
    layer3_outputs(7954) <= not(layer2_outputs(997));
    layer3_outputs(7955) <= not((layer2_outputs(3318)) and (layer2_outputs(3281)));
    layer3_outputs(7956) <= not(layer2_outputs(109));
    layer3_outputs(7957) <= layer2_outputs(9524);
    layer3_outputs(7958) <= not((layer2_outputs(7677)) and (layer2_outputs(5009)));
    layer3_outputs(7959) <= not(layer2_outputs(3664));
    layer3_outputs(7960) <= not((layer2_outputs(3544)) xor (layer2_outputs(8912)));
    layer3_outputs(7961) <= not(layer2_outputs(8534));
    layer3_outputs(7962) <= not((layer2_outputs(220)) xor (layer2_outputs(4707)));
    layer3_outputs(7963) <= not((layer2_outputs(9135)) xor (layer2_outputs(5855)));
    layer3_outputs(7964) <= (layer2_outputs(1142)) and not (layer2_outputs(7792));
    layer3_outputs(7965) <= (layer2_outputs(7761)) and (layer2_outputs(734));
    layer3_outputs(7966) <= not(layer2_outputs(7695));
    layer3_outputs(7967) <= not(layer2_outputs(3407)) or (layer2_outputs(860));
    layer3_outputs(7968) <= not((layer2_outputs(104)) or (layer2_outputs(4381)));
    layer3_outputs(7969) <= '1';
    layer3_outputs(7970) <= not(layer2_outputs(5674));
    layer3_outputs(7971) <= layer2_outputs(6365);
    layer3_outputs(7972) <= (layer2_outputs(9019)) or (layer2_outputs(3899));
    layer3_outputs(7973) <= not(layer2_outputs(9414));
    layer3_outputs(7974) <= not((layer2_outputs(4079)) or (layer2_outputs(7551)));
    layer3_outputs(7975) <= not(layer2_outputs(6368));
    layer3_outputs(7976) <= not((layer2_outputs(9204)) xor (layer2_outputs(1130)));
    layer3_outputs(7977) <= (layer2_outputs(1125)) and not (layer2_outputs(360));
    layer3_outputs(7978) <= layer2_outputs(7420);
    layer3_outputs(7979) <= (layer2_outputs(10235)) or (layer2_outputs(5876));
    layer3_outputs(7980) <= (layer2_outputs(19)) and not (layer2_outputs(1434));
    layer3_outputs(7981) <= (layer2_outputs(1880)) and not (layer2_outputs(3922));
    layer3_outputs(7982) <= not(layer2_outputs(9269));
    layer3_outputs(7983) <= layer2_outputs(8719);
    layer3_outputs(7984) <= (layer2_outputs(7361)) and not (layer2_outputs(9213));
    layer3_outputs(7985) <= layer2_outputs(6422);
    layer3_outputs(7986) <= layer2_outputs(2146);
    layer3_outputs(7987) <= not((layer2_outputs(1754)) or (layer2_outputs(5959)));
    layer3_outputs(7988) <= not(layer2_outputs(856));
    layer3_outputs(7989) <= '1';
    layer3_outputs(7990) <= not((layer2_outputs(6545)) and (layer2_outputs(1008)));
    layer3_outputs(7991) <= not((layer2_outputs(4074)) and (layer2_outputs(3048)));
    layer3_outputs(7992) <= not(layer2_outputs(9741));
    layer3_outputs(7993) <= (layer2_outputs(6437)) and (layer2_outputs(2603));
    layer3_outputs(7994) <= (layer2_outputs(142)) and not (layer2_outputs(5664));
    layer3_outputs(7995) <= not(layer2_outputs(4183));
    layer3_outputs(7996) <= not((layer2_outputs(7250)) xor (layer2_outputs(8784)));
    layer3_outputs(7997) <= (layer2_outputs(8569)) and (layer2_outputs(8295));
    layer3_outputs(7998) <= not((layer2_outputs(8073)) xor (layer2_outputs(6073)));
    layer3_outputs(7999) <= layer2_outputs(2658);
    layer3_outputs(8000) <= not((layer2_outputs(8206)) xor (layer2_outputs(7582)));
    layer3_outputs(8001) <= (layer2_outputs(8480)) or (layer2_outputs(7934));
    layer3_outputs(8002) <= layer2_outputs(9098);
    layer3_outputs(8003) <= not(layer2_outputs(7728));
    layer3_outputs(8004) <= not(layer2_outputs(5447));
    layer3_outputs(8005) <= (layer2_outputs(2701)) xor (layer2_outputs(2905));
    layer3_outputs(8006) <= (layer2_outputs(1795)) or (layer2_outputs(2990));
    layer3_outputs(8007) <= not((layer2_outputs(5112)) and (layer2_outputs(6914)));
    layer3_outputs(8008) <= layer2_outputs(7094);
    layer3_outputs(8009) <= not(layer2_outputs(9059));
    layer3_outputs(8010) <= not((layer2_outputs(6682)) or (layer2_outputs(1936)));
    layer3_outputs(8011) <= layer2_outputs(6362);
    layer3_outputs(8012) <= (layer2_outputs(6455)) xor (layer2_outputs(4774));
    layer3_outputs(8013) <= (layer2_outputs(7546)) and not (layer2_outputs(6418));
    layer3_outputs(8014) <= layer2_outputs(8014);
    layer3_outputs(8015) <= not(layer2_outputs(8028)) or (layer2_outputs(7928));
    layer3_outputs(8016) <= layer2_outputs(2591);
    layer3_outputs(8017) <= (layer2_outputs(6407)) or (layer2_outputs(1497));
    layer3_outputs(8018) <= not(layer2_outputs(3217));
    layer3_outputs(8019) <= layer2_outputs(6355);
    layer3_outputs(8020) <= not(layer2_outputs(6167)) or (layer2_outputs(9557));
    layer3_outputs(8021) <= not(layer2_outputs(8803)) or (layer2_outputs(1879));
    layer3_outputs(8022) <= not((layer2_outputs(5618)) xor (layer2_outputs(4953)));
    layer3_outputs(8023) <= layer2_outputs(10184);
    layer3_outputs(8024) <= layer2_outputs(6234);
    layer3_outputs(8025) <= not(layer2_outputs(8095)) or (layer2_outputs(6950));
    layer3_outputs(8026) <= not((layer2_outputs(2830)) xor (layer2_outputs(2652)));
    layer3_outputs(8027) <= (layer2_outputs(9682)) and not (layer2_outputs(1463));
    layer3_outputs(8028) <= layer2_outputs(3583);
    layer3_outputs(8029) <= (layer2_outputs(3521)) and not (layer2_outputs(5382));
    layer3_outputs(8030) <= '1';
    layer3_outputs(8031) <= layer2_outputs(8184);
    layer3_outputs(8032) <= not(layer2_outputs(8581));
    layer3_outputs(8033) <= not(layer2_outputs(4287));
    layer3_outputs(8034) <= layer2_outputs(4176);
    layer3_outputs(8035) <= (layer2_outputs(6256)) and not (layer2_outputs(9338));
    layer3_outputs(8036) <= (layer2_outputs(5729)) and not (layer2_outputs(7207));
    layer3_outputs(8037) <= not(layer2_outputs(8715));
    layer3_outputs(8038) <= not((layer2_outputs(7190)) xor (layer2_outputs(7759)));
    layer3_outputs(8039) <= layer2_outputs(369);
    layer3_outputs(8040) <= not(layer2_outputs(7966));
    layer3_outputs(8041) <= not(layer2_outputs(946));
    layer3_outputs(8042) <= not(layer2_outputs(5806));
    layer3_outputs(8043) <= not((layer2_outputs(4033)) xor (layer2_outputs(4272)));
    layer3_outputs(8044) <= not(layer2_outputs(8472));
    layer3_outputs(8045) <= (layer2_outputs(7454)) or (layer2_outputs(8140));
    layer3_outputs(8046) <= not(layer2_outputs(9628));
    layer3_outputs(8047) <= not(layer2_outputs(3559));
    layer3_outputs(8048) <= layer2_outputs(9558);
    layer3_outputs(8049) <= layer2_outputs(9763);
    layer3_outputs(8050) <= not(layer2_outputs(7744));
    layer3_outputs(8051) <= not((layer2_outputs(7497)) xor (layer2_outputs(6547)));
    layer3_outputs(8052) <= not(layer2_outputs(517));
    layer3_outputs(8053) <= (layer2_outputs(7611)) and (layer2_outputs(1578));
    layer3_outputs(8054) <= (layer2_outputs(688)) xor (layer2_outputs(8076));
    layer3_outputs(8055) <= layer2_outputs(6464);
    layer3_outputs(8056) <= not(layer2_outputs(1619));
    layer3_outputs(8057) <= (layer2_outputs(6607)) and not (layer2_outputs(4016));
    layer3_outputs(8058) <= layer2_outputs(6754);
    layer3_outputs(8059) <= layer2_outputs(8558);
    layer3_outputs(8060) <= (layer2_outputs(7371)) or (layer2_outputs(5537));
    layer3_outputs(8061) <= '0';
    layer3_outputs(8062) <= (layer2_outputs(8372)) and not (layer2_outputs(7570));
    layer3_outputs(8063) <= not(layer2_outputs(4700));
    layer3_outputs(8064) <= not(layer2_outputs(4285));
    layer3_outputs(8065) <= layer2_outputs(1956);
    layer3_outputs(8066) <= not(layer2_outputs(2778));
    layer3_outputs(8067) <= not(layer2_outputs(8108));
    layer3_outputs(8068) <= not((layer2_outputs(1116)) or (layer2_outputs(6184)));
    layer3_outputs(8069) <= not(layer2_outputs(4056));
    layer3_outputs(8070) <= not((layer2_outputs(9513)) xor (layer2_outputs(7004)));
    layer3_outputs(8071) <= layer2_outputs(1881);
    layer3_outputs(8072) <= '1';
    layer3_outputs(8073) <= not((layer2_outputs(1057)) and (layer2_outputs(1597)));
    layer3_outputs(8074) <= not(layer2_outputs(1334));
    layer3_outputs(8075) <= not(layer2_outputs(7339));
    layer3_outputs(8076) <= not(layer2_outputs(6032));
    layer3_outputs(8077) <= not(layer2_outputs(3369));
    layer3_outputs(8078) <= layer2_outputs(1906);
    layer3_outputs(8079) <= layer2_outputs(780);
    layer3_outputs(8080) <= (layer2_outputs(1836)) and (layer2_outputs(1988));
    layer3_outputs(8081) <= layer2_outputs(3182);
    layer3_outputs(8082) <= not(layer2_outputs(6023));
    layer3_outputs(8083) <= not(layer2_outputs(3331));
    layer3_outputs(8084) <= (layer2_outputs(5391)) or (layer2_outputs(1781));
    layer3_outputs(8085) <= (layer2_outputs(3359)) or (layer2_outputs(7348));
    layer3_outputs(8086) <= not(layer2_outputs(2033));
    layer3_outputs(8087) <= not(layer2_outputs(1359)) or (layer2_outputs(8340));
    layer3_outputs(8088) <= layer2_outputs(7806);
    layer3_outputs(8089) <= not(layer2_outputs(7918));
    layer3_outputs(8090) <= not(layer2_outputs(188));
    layer3_outputs(8091) <= not((layer2_outputs(10046)) xor (layer2_outputs(8933)));
    layer3_outputs(8092) <= not(layer2_outputs(468));
    layer3_outputs(8093) <= (layer2_outputs(7970)) or (layer2_outputs(9971));
    layer3_outputs(8094) <= not(layer2_outputs(1056));
    layer3_outputs(8095) <= not(layer2_outputs(1417));
    layer3_outputs(8096) <= not((layer2_outputs(7769)) xor (layer2_outputs(2779)));
    layer3_outputs(8097) <= '0';
    layer3_outputs(8098) <= not((layer2_outputs(6201)) and (layer2_outputs(9428)));
    layer3_outputs(8099) <= not((layer2_outputs(3256)) xor (layer2_outputs(5098)));
    layer3_outputs(8100) <= layer2_outputs(1137);
    layer3_outputs(8101) <= (layer2_outputs(4861)) xor (layer2_outputs(3288));
    layer3_outputs(8102) <= not(layer2_outputs(11));
    layer3_outputs(8103) <= '1';
    layer3_outputs(8104) <= (layer2_outputs(6111)) and not (layer2_outputs(1166));
    layer3_outputs(8105) <= not((layer2_outputs(2459)) xor (layer2_outputs(7964)));
    layer3_outputs(8106) <= layer2_outputs(10107);
    layer3_outputs(8107) <= (layer2_outputs(3552)) or (layer2_outputs(525));
    layer3_outputs(8108) <= (layer2_outputs(1759)) xor (layer2_outputs(4008));
    layer3_outputs(8109) <= not(layer2_outputs(4283)) or (layer2_outputs(7796));
    layer3_outputs(8110) <= '1';
    layer3_outputs(8111) <= (layer2_outputs(9659)) and not (layer2_outputs(2907));
    layer3_outputs(8112) <= not((layer2_outputs(8044)) or (layer2_outputs(1051)));
    layer3_outputs(8113) <= layer2_outputs(7250);
    layer3_outputs(8114) <= (layer2_outputs(4770)) and not (layer2_outputs(831));
    layer3_outputs(8115) <= layer2_outputs(7492);
    layer3_outputs(8116) <= (layer2_outputs(837)) xor (layer2_outputs(4846));
    layer3_outputs(8117) <= '1';
    layer3_outputs(8118) <= not((layer2_outputs(2200)) xor (layer2_outputs(9626)));
    layer3_outputs(8119) <= layer2_outputs(7389);
    layer3_outputs(8120) <= layer2_outputs(8786);
    layer3_outputs(8121) <= not((layer2_outputs(10192)) or (layer2_outputs(5950)));
    layer3_outputs(8122) <= not(layer2_outputs(4310));
    layer3_outputs(8123) <= not((layer2_outputs(6756)) or (layer2_outputs(5754)));
    layer3_outputs(8124) <= layer2_outputs(3980);
    layer3_outputs(8125) <= not(layer2_outputs(2690));
    layer3_outputs(8126) <= layer2_outputs(1338);
    layer3_outputs(8127) <= not(layer2_outputs(8795));
    layer3_outputs(8128) <= not((layer2_outputs(3431)) or (layer2_outputs(9146)));
    layer3_outputs(8129) <= not(layer2_outputs(9559));
    layer3_outputs(8130) <= (layer2_outputs(5050)) xor (layer2_outputs(3506));
    layer3_outputs(8131) <= (layer2_outputs(4768)) and (layer2_outputs(9261));
    layer3_outputs(8132) <= (layer2_outputs(6563)) and not (layer2_outputs(6285));
    layer3_outputs(8133) <= layer2_outputs(168);
    layer3_outputs(8134) <= not((layer2_outputs(9576)) and (layer2_outputs(9773)));
    layer3_outputs(8135) <= (layer2_outputs(8113)) and not (layer2_outputs(5279));
    layer3_outputs(8136) <= (layer2_outputs(3072)) xor (layer2_outputs(6212));
    layer3_outputs(8137) <= not((layer2_outputs(5823)) and (layer2_outputs(6685)));
    layer3_outputs(8138) <= (layer2_outputs(7766)) and not (layer2_outputs(5721));
    layer3_outputs(8139) <= not(layer2_outputs(9530));
    layer3_outputs(8140) <= '1';
    layer3_outputs(8141) <= (layer2_outputs(2156)) and not (layer2_outputs(238));
    layer3_outputs(8142) <= not(layer2_outputs(8718));
    layer3_outputs(8143) <= not(layer2_outputs(1538));
    layer3_outputs(8144) <= layer2_outputs(9066);
    layer3_outputs(8145) <= (layer2_outputs(6420)) and (layer2_outputs(3079));
    layer3_outputs(8146) <= not((layer2_outputs(1035)) or (layer2_outputs(4364)));
    layer3_outputs(8147) <= layer2_outputs(2370);
    layer3_outputs(8148) <= not(layer2_outputs(7035));
    layer3_outputs(8149) <= not((layer2_outputs(3913)) or (layer2_outputs(528)));
    layer3_outputs(8150) <= not(layer2_outputs(2096));
    layer3_outputs(8151) <= not((layer2_outputs(9373)) or (layer2_outputs(7490)));
    layer3_outputs(8152) <= not(layer2_outputs(5251)) or (layer2_outputs(9850));
    layer3_outputs(8153) <= layer2_outputs(1996);
    layer3_outputs(8154) <= not(layer2_outputs(5084));
    layer3_outputs(8155) <= not(layer2_outputs(6089)) or (layer2_outputs(9700));
    layer3_outputs(8156) <= not((layer2_outputs(4451)) xor (layer2_outputs(4123)));
    layer3_outputs(8157) <= not((layer2_outputs(6664)) or (layer2_outputs(2070)));
    layer3_outputs(8158) <= not((layer2_outputs(2945)) xor (layer2_outputs(3368)));
    layer3_outputs(8159) <= not(layer2_outputs(7892));
    layer3_outputs(8160) <= not((layer2_outputs(7590)) or (layer2_outputs(1739)));
    layer3_outputs(8161) <= '1';
    layer3_outputs(8162) <= (layer2_outputs(9631)) and not (layer2_outputs(4037));
    layer3_outputs(8163) <= (layer2_outputs(753)) and not (layer2_outputs(9184));
    layer3_outputs(8164) <= not((layer2_outputs(3410)) xor (layer2_outputs(6508)));
    layer3_outputs(8165) <= (layer2_outputs(5563)) and (layer2_outputs(1306));
    layer3_outputs(8166) <= layer2_outputs(3052);
    layer3_outputs(8167) <= not(layer2_outputs(8226));
    layer3_outputs(8168) <= (layer2_outputs(1251)) and (layer2_outputs(3824));
    layer3_outputs(8169) <= (layer2_outputs(5898)) and (layer2_outputs(8254));
    layer3_outputs(8170) <= layer2_outputs(4834);
    layer3_outputs(8171) <= (layer2_outputs(7819)) and not (layer2_outputs(3451));
    layer3_outputs(8172) <= layer2_outputs(408);
    layer3_outputs(8173) <= '1';
    layer3_outputs(8174) <= (layer2_outputs(4811)) and not (layer2_outputs(2338));
    layer3_outputs(8175) <= layer2_outputs(1520);
    layer3_outputs(8176) <= not(layer2_outputs(511));
    layer3_outputs(8177) <= not(layer2_outputs(1298));
    layer3_outputs(8178) <= not(layer2_outputs(793));
    layer3_outputs(8179) <= (layer2_outputs(9520)) and not (layer2_outputs(714));
    layer3_outputs(8180) <= not(layer2_outputs(2219)) or (layer2_outputs(7149));
    layer3_outputs(8181) <= '0';
    layer3_outputs(8182) <= layer2_outputs(4526);
    layer3_outputs(8183) <= layer2_outputs(10081);
    layer3_outputs(8184) <= layer2_outputs(4313);
    layer3_outputs(8185) <= not(layer2_outputs(7537));
    layer3_outputs(8186) <= not(layer2_outputs(5049)) or (layer2_outputs(3219));
    layer3_outputs(8187) <= (layer2_outputs(5080)) xor (layer2_outputs(4590));
    layer3_outputs(8188) <= not((layer2_outputs(4328)) or (layer2_outputs(330)));
    layer3_outputs(8189) <= not((layer2_outputs(9046)) or (layer2_outputs(2795)));
    layer3_outputs(8190) <= not(layer2_outputs(7376));
    layer3_outputs(8191) <= not((layer2_outputs(6766)) and (layer2_outputs(7379)));
    layer3_outputs(8192) <= (layer2_outputs(194)) and not (layer2_outputs(3443));
    layer3_outputs(8193) <= layer2_outputs(8453);
    layer3_outputs(8194) <= not(layer2_outputs(4700)) or (layer2_outputs(6430));
    layer3_outputs(8195) <= not(layer2_outputs(9305));
    layer3_outputs(8196) <= layer2_outputs(1317);
    layer3_outputs(8197) <= not(layer2_outputs(9547)) or (layer2_outputs(6246));
    layer3_outputs(8198) <= layer2_outputs(6297);
    layer3_outputs(8199) <= layer2_outputs(2821);
    layer3_outputs(8200) <= not(layer2_outputs(7148));
    layer3_outputs(8201) <= (layer2_outputs(3027)) or (layer2_outputs(6554));
    layer3_outputs(8202) <= layer2_outputs(8403);
    layer3_outputs(8203) <= (layer2_outputs(5798)) and (layer2_outputs(8913));
    layer3_outputs(8204) <= layer2_outputs(9745);
    layer3_outputs(8205) <= (layer2_outputs(1250)) or (layer2_outputs(3933));
    layer3_outputs(8206) <= not(layer2_outputs(8260));
    layer3_outputs(8207) <= not(layer2_outputs(7596));
    layer3_outputs(8208) <= not(layer2_outputs(5179));
    layer3_outputs(8209) <= layer2_outputs(8423);
    layer3_outputs(8210) <= layer2_outputs(5586);
    layer3_outputs(8211) <= not((layer2_outputs(9986)) or (layer2_outputs(2459)));
    layer3_outputs(8212) <= layer2_outputs(6421);
    layer3_outputs(8213) <= not((layer2_outputs(8648)) and (layer2_outputs(1727)));
    layer3_outputs(8214) <= (layer2_outputs(391)) xor (layer2_outputs(4785));
    layer3_outputs(8215) <= not(layer2_outputs(4215));
    layer3_outputs(8216) <= (layer2_outputs(8245)) and not (layer2_outputs(7612));
    layer3_outputs(8217) <= layer2_outputs(3096);
    layer3_outputs(8218) <= (layer2_outputs(1412)) and not (layer2_outputs(6887));
    layer3_outputs(8219) <= layer2_outputs(3700);
    layer3_outputs(8220) <= not(layer2_outputs(6827));
    layer3_outputs(8221) <= (layer2_outputs(8477)) and (layer2_outputs(6922));
    layer3_outputs(8222) <= not(layer2_outputs(104));
    layer3_outputs(8223) <= layer2_outputs(9750);
    layer3_outputs(8224) <= not(layer2_outputs(4403));
    layer3_outputs(8225) <= not((layer2_outputs(3259)) and (layer2_outputs(2356)));
    layer3_outputs(8226) <= not(layer2_outputs(6793)) or (layer2_outputs(4734));
    layer3_outputs(8227) <= not((layer2_outputs(7192)) xor (layer2_outputs(4306)));
    layer3_outputs(8228) <= not((layer2_outputs(4785)) xor (layer2_outputs(6660)));
    layer3_outputs(8229) <= layer2_outputs(4287);
    layer3_outputs(8230) <= layer2_outputs(1460);
    layer3_outputs(8231) <= (layer2_outputs(6202)) and not (layer2_outputs(8768));
    layer3_outputs(8232) <= not(layer2_outputs(10209)) or (layer2_outputs(3537));
    layer3_outputs(8233) <= not(layer2_outputs(597));
    layer3_outputs(8234) <= not((layer2_outputs(1964)) and (layer2_outputs(9522)));
    layer3_outputs(8235) <= not(layer2_outputs(7622));
    layer3_outputs(8236) <= not(layer2_outputs(2149)) or (layer2_outputs(569));
    layer3_outputs(8237) <= layer2_outputs(8386);
    layer3_outputs(8238) <= layer2_outputs(4681);
    layer3_outputs(8239) <= not(layer2_outputs(4215));
    layer3_outputs(8240) <= layer2_outputs(3061);
    layer3_outputs(8241) <= not((layer2_outputs(1845)) and (layer2_outputs(7171)));
    layer3_outputs(8242) <= not((layer2_outputs(1411)) and (layer2_outputs(3641)));
    layer3_outputs(8243) <= not(layer2_outputs(5545));
    layer3_outputs(8244) <= not(layer2_outputs(6886));
    layer3_outputs(8245) <= '1';
    layer3_outputs(8246) <= not(layer2_outputs(2617));
    layer3_outputs(8247) <= not((layer2_outputs(3175)) xor (layer2_outputs(8146)));
    layer3_outputs(8248) <= not((layer2_outputs(4477)) xor (layer2_outputs(634)));
    layer3_outputs(8249) <= not(layer2_outputs(4643));
    layer3_outputs(8250) <= not(layer2_outputs(10018));
    layer3_outputs(8251) <= not(layer2_outputs(6192));
    layer3_outputs(8252) <= layer2_outputs(1371);
    layer3_outputs(8253) <= layer2_outputs(6940);
    layer3_outputs(8254) <= (layer2_outputs(8963)) xor (layer2_outputs(9639));
    layer3_outputs(8255) <= not(layer2_outputs(9690)) or (layer2_outputs(2663));
    layer3_outputs(8256) <= layer2_outputs(3409);
    layer3_outputs(8257) <= layer2_outputs(7417);
    layer3_outputs(8258) <= not(layer2_outputs(4962)) or (layer2_outputs(4439));
    layer3_outputs(8259) <= layer2_outputs(1855);
    layer3_outputs(8260) <= not((layer2_outputs(3107)) xor (layer2_outputs(2088)));
    layer3_outputs(8261) <= layer2_outputs(5029);
    layer3_outputs(8262) <= not(layer2_outputs(7622));
    layer3_outputs(8263) <= (layer2_outputs(10001)) and not (layer2_outputs(7693));
    layer3_outputs(8264) <= (layer2_outputs(3591)) or (layer2_outputs(69));
    layer3_outputs(8265) <= not(layer2_outputs(9585)) or (layer2_outputs(30));
    layer3_outputs(8266) <= not(layer2_outputs(3318));
    layer3_outputs(8267) <= (layer2_outputs(961)) and (layer2_outputs(4881));
    layer3_outputs(8268) <= '1';
    layer3_outputs(8269) <= not(layer2_outputs(9307));
    layer3_outputs(8270) <= (layer2_outputs(8826)) and not (layer2_outputs(4336));
    layer3_outputs(8271) <= (layer2_outputs(1602)) or (layer2_outputs(588));
    layer3_outputs(8272) <= not(layer2_outputs(9037));
    layer3_outputs(8273) <= layer2_outputs(1922);
    layer3_outputs(8274) <= (layer2_outputs(3150)) or (layer2_outputs(8502));
    layer3_outputs(8275) <= not((layer2_outputs(4338)) or (layer2_outputs(2435)));
    layer3_outputs(8276) <= layer2_outputs(7274);
    layer3_outputs(8277) <= layer2_outputs(9936);
    layer3_outputs(8278) <= layer2_outputs(239);
    layer3_outputs(8279) <= layer2_outputs(5996);
    layer3_outputs(8280) <= not(layer2_outputs(5857));
    layer3_outputs(8281) <= not(layer2_outputs(3632)) or (layer2_outputs(8314));
    layer3_outputs(8282) <= layer2_outputs(4053);
    layer3_outputs(8283) <= (layer2_outputs(8905)) and (layer2_outputs(7329));
    layer3_outputs(8284) <= (layer2_outputs(5438)) and not (layer2_outputs(5007));
    layer3_outputs(8285) <= layer2_outputs(3711);
    layer3_outputs(8286) <= (layer2_outputs(8330)) or (layer2_outputs(2458));
    layer3_outputs(8287) <= not(layer2_outputs(222));
    layer3_outputs(8288) <= not((layer2_outputs(9419)) xor (layer2_outputs(5689)));
    layer3_outputs(8289) <= not((layer2_outputs(5418)) xor (layer2_outputs(5176)));
    layer3_outputs(8290) <= (layer2_outputs(6391)) and not (layer2_outputs(8728));
    layer3_outputs(8291) <= layer2_outputs(8225);
    layer3_outputs(8292) <= layer2_outputs(6668);
    layer3_outputs(8293) <= not((layer2_outputs(7253)) and (layer2_outputs(4199)));
    layer3_outputs(8294) <= layer2_outputs(3042);
    layer3_outputs(8295) <= (layer2_outputs(2620)) xor (layer2_outputs(3330));
    layer3_outputs(8296) <= not(layer2_outputs(3620));
    layer3_outputs(8297) <= not(layer2_outputs(5788)) or (layer2_outputs(4041));
    layer3_outputs(8298) <= not(layer2_outputs(5667));
    layer3_outputs(8299) <= not((layer2_outputs(5793)) xor (layer2_outputs(7169)));
    layer3_outputs(8300) <= not(layer2_outputs(8269));
    layer3_outputs(8301) <= layer2_outputs(9653);
    layer3_outputs(8302) <= layer2_outputs(2403);
    layer3_outputs(8303) <= not(layer2_outputs(216));
    layer3_outputs(8304) <= not(layer2_outputs(8989)) or (layer2_outputs(2164));
    layer3_outputs(8305) <= layer2_outputs(9733);
    layer3_outputs(8306) <= layer2_outputs(7848);
    layer3_outputs(8307) <= (layer2_outputs(6823)) and (layer2_outputs(334));
    layer3_outputs(8308) <= not(layer2_outputs(7330));
    layer3_outputs(8309) <= not(layer2_outputs(2681)) or (layer2_outputs(4919));
    layer3_outputs(8310) <= layer2_outputs(73);
    layer3_outputs(8311) <= not(layer2_outputs(4862)) or (layer2_outputs(758));
    layer3_outputs(8312) <= not(layer2_outputs(2046));
    layer3_outputs(8313) <= not(layer2_outputs(1147));
    layer3_outputs(8314) <= not(layer2_outputs(5676));
    layer3_outputs(8315) <= not(layer2_outputs(1639));
    layer3_outputs(8316) <= not(layer2_outputs(7790));
    layer3_outputs(8317) <= not(layer2_outputs(1156)) or (layer2_outputs(8636));
    layer3_outputs(8318) <= not(layer2_outputs(698));
    layer3_outputs(8319) <= (layer2_outputs(1673)) and not (layer2_outputs(6891));
    layer3_outputs(8320) <= not((layer2_outputs(5069)) or (layer2_outputs(5467)));
    layer3_outputs(8321) <= '0';
    layer3_outputs(8322) <= layer2_outputs(5414);
    layer3_outputs(8323) <= layer2_outputs(1058);
    layer3_outputs(8324) <= not(layer2_outputs(1769));
    layer3_outputs(8325) <= not((layer2_outputs(2091)) xor (layer2_outputs(4002)));
    layer3_outputs(8326) <= '0';
    layer3_outputs(8327) <= (layer2_outputs(8787)) xor (layer2_outputs(1577));
    layer3_outputs(8328) <= not(layer2_outputs(2539));
    layer3_outputs(8329) <= (layer2_outputs(1844)) and not (layer2_outputs(8521));
    layer3_outputs(8330) <= '1';
    layer3_outputs(8331) <= (layer2_outputs(2348)) and (layer2_outputs(8732));
    layer3_outputs(8332) <= not((layer2_outputs(7182)) and (layer2_outputs(481)));
    layer3_outputs(8333) <= layer2_outputs(9990);
    layer3_outputs(8334) <= not(layer2_outputs(6241));
    layer3_outputs(8335) <= not(layer2_outputs(5917)) or (layer2_outputs(2450));
    layer3_outputs(8336) <= not(layer2_outputs(2277));
    layer3_outputs(8337) <= layer2_outputs(4497);
    layer3_outputs(8338) <= layer2_outputs(8155);
    layer3_outputs(8339) <= (layer2_outputs(8377)) and not (layer2_outputs(8521));
    layer3_outputs(8340) <= not((layer2_outputs(6328)) and (layer2_outputs(3203)));
    layer3_outputs(8341) <= not(layer2_outputs(757)) or (layer2_outputs(3892));
    layer3_outputs(8342) <= not(layer2_outputs(2310));
    layer3_outputs(8343) <= (layer2_outputs(3656)) and (layer2_outputs(2482));
    layer3_outputs(8344) <= layer2_outputs(5806);
    layer3_outputs(8345) <= layer2_outputs(9413);
    layer3_outputs(8346) <= not(layer2_outputs(483)) or (layer2_outputs(7069));
    layer3_outputs(8347) <= not(layer2_outputs(6576));
    layer3_outputs(8348) <= (layer2_outputs(6729)) or (layer2_outputs(362));
    layer3_outputs(8349) <= not(layer2_outputs(2102));
    layer3_outputs(8350) <= (layer2_outputs(5222)) or (layer2_outputs(2712));
    layer3_outputs(8351) <= not((layer2_outputs(8394)) xor (layer2_outputs(1251)));
    layer3_outputs(8352) <= not(layer2_outputs(8517));
    layer3_outputs(8353) <= '0';
    layer3_outputs(8354) <= (layer2_outputs(485)) and not (layer2_outputs(2703));
    layer3_outputs(8355) <= not(layer2_outputs(4573));
    layer3_outputs(8356) <= not(layer2_outputs(536));
    layer3_outputs(8357) <= '0';
    layer3_outputs(8358) <= (layer2_outputs(4213)) and not (layer2_outputs(1477));
    layer3_outputs(8359) <= layer2_outputs(1414);
    layer3_outputs(8360) <= (layer2_outputs(6674)) xor (layer2_outputs(7048));
    layer3_outputs(8361) <= (layer2_outputs(7931)) and not (layer2_outputs(4788));
    layer3_outputs(8362) <= not(layer2_outputs(1379)) or (layer2_outputs(7788));
    layer3_outputs(8363) <= layer2_outputs(634);
    layer3_outputs(8364) <= layer2_outputs(270);
    layer3_outputs(8365) <= not((layer2_outputs(8097)) or (layer2_outputs(7953)));
    layer3_outputs(8366) <= not((layer2_outputs(3161)) or (layer2_outputs(7205)));
    layer3_outputs(8367) <= not(layer2_outputs(3911)) or (layer2_outputs(406));
    layer3_outputs(8368) <= (layer2_outputs(15)) and (layer2_outputs(10012));
    layer3_outputs(8369) <= not(layer2_outputs(6637));
    layer3_outputs(8370) <= not(layer2_outputs(8706));
    layer3_outputs(8371) <= layer2_outputs(189);
    layer3_outputs(8372) <= not(layer2_outputs(8228));
    layer3_outputs(8373) <= not((layer2_outputs(9728)) or (layer2_outputs(3408)));
    layer3_outputs(8374) <= not(layer2_outputs(7719));
    layer3_outputs(8375) <= (layer2_outputs(2788)) and (layer2_outputs(8806));
    layer3_outputs(8376) <= not(layer2_outputs(4481));
    layer3_outputs(8377) <= (layer2_outputs(8987)) or (layer2_outputs(5399));
    layer3_outputs(8378) <= layer2_outputs(2858);
    layer3_outputs(8379) <= layer2_outputs(3309);
    layer3_outputs(8380) <= (layer2_outputs(5902)) and (layer2_outputs(1764));
    layer3_outputs(8381) <= layer2_outputs(5999);
    layer3_outputs(8382) <= not((layer2_outputs(5979)) xor (layer2_outputs(3923)));
    layer3_outputs(8383) <= (layer2_outputs(7882)) xor (layer2_outputs(548));
    layer3_outputs(8384) <= not(layer2_outputs(5258));
    layer3_outputs(8385) <= layer2_outputs(9074);
    layer3_outputs(8386) <= (layer2_outputs(1773)) or (layer2_outputs(3523));
    layer3_outputs(8387) <= layer2_outputs(6129);
    layer3_outputs(8388) <= not(layer2_outputs(8991));
    layer3_outputs(8389) <= not(layer2_outputs(6090));
    layer3_outputs(8390) <= not(layer2_outputs(7431));
    layer3_outputs(8391) <= not(layer2_outputs(4747)) or (layer2_outputs(9837));
    layer3_outputs(8392) <= not((layer2_outputs(652)) xor (layer2_outputs(7156)));
    layer3_outputs(8393) <= not(layer2_outputs(9256)) or (layer2_outputs(2779));
    layer3_outputs(8394) <= not(layer2_outputs(6215)) or (layer2_outputs(3328));
    layer3_outputs(8395) <= not(layer2_outputs(7390)) or (layer2_outputs(9016));
    layer3_outputs(8396) <= (layer2_outputs(8422)) xor (layer2_outputs(10048));
    layer3_outputs(8397) <= layer2_outputs(5324);
    layer3_outputs(8398) <= (layer2_outputs(4513)) or (layer2_outputs(7170));
    layer3_outputs(8399) <= (layer2_outputs(2067)) and not (layer2_outputs(6475));
    layer3_outputs(8400) <= not(layer2_outputs(3785)) or (layer2_outputs(632));
    layer3_outputs(8401) <= (layer2_outputs(7326)) xor (layer2_outputs(8783));
    layer3_outputs(8402) <= not((layer2_outputs(3903)) and (layer2_outputs(9956)));
    layer3_outputs(8403) <= layer2_outputs(3889);
    layer3_outputs(8404) <= (layer2_outputs(2427)) and (layer2_outputs(9829));
    layer3_outputs(8405) <= (layer2_outputs(920)) xor (layer2_outputs(8326));
    layer3_outputs(8406) <= not(layer2_outputs(442)) or (layer2_outputs(4908));
    layer3_outputs(8407) <= not((layer2_outputs(7119)) and (layer2_outputs(4005)));
    layer3_outputs(8408) <= not(layer2_outputs(3333)) or (layer2_outputs(1112));
    layer3_outputs(8409) <= not(layer2_outputs(5443));
    layer3_outputs(8410) <= layer2_outputs(144);
    layer3_outputs(8411) <= layer2_outputs(9151);
    layer3_outputs(8412) <= not(layer2_outputs(5299));
    layer3_outputs(8413) <= (layer2_outputs(7689)) xor (layer2_outputs(4099));
    layer3_outputs(8414) <= not(layer2_outputs(8147));
    layer3_outputs(8415) <= not((layer2_outputs(4823)) xor (layer2_outputs(1907)));
    layer3_outputs(8416) <= not(layer2_outputs(3370)) or (layer2_outputs(2415));
    layer3_outputs(8417) <= layer2_outputs(9454);
    layer3_outputs(8418) <= layer2_outputs(2355);
    layer3_outputs(8419) <= not(layer2_outputs(695));
    layer3_outputs(8420) <= not((layer2_outputs(2735)) xor (layer2_outputs(6552)));
    layer3_outputs(8421) <= not(layer2_outputs(3489));
    layer3_outputs(8422) <= not(layer2_outputs(1448)) or (layer2_outputs(1418));
    layer3_outputs(8423) <= (layer2_outputs(4715)) and (layer2_outputs(5884));
    layer3_outputs(8424) <= not((layer2_outputs(6828)) or (layer2_outputs(2339)));
    layer3_outputs(8425) <= (layer2_outputs(1998)) and not (layer2_outputs(8191));
    layer3_outputs(8426) <= not(layer2_outputs(7969));
    layer3_outputs(8427) <= (layer2_outputs(881)) xor (layer2_outputs(9262));
    layer3_outputs(8428) <= not(layer2_outputs(9576)) or (layer2_outputs(9488));
    layer3_outputs(8429) <= not(layer2_outputs(1270)) or (layer2_outputs(3701));
    layer3_outputs(8430) <= layer2_outputs(350);
    layer3_outputs(8431) <= layer2_outputs(3179);
    layer3_outputs(8432) <= '0';
    layer3_outputs(8433) <= layer2_outputs(2564);
    layer3_outputs(8434) <= (layer2_outputs(6803)) and not (layer2_outputs(382));
    layer3_outputs(8435) <= not((layer2_outputs(4246)) xor (layer2_outputs(9892)));
    layer3_outputs(8436) <= not(layer2_outputs(9123));
    layer3_outputs(8437) <= not(layer2_outputs(4888));
    layer3_outputs(8438) <= not(layer2_outputs(448)) or (layer2_outputs(9715));
    layer3_outputs(8439) <= not(layer2_outputs(920)) or (layer2_outputs(9770));
    layer3_outputs(8440) <= layer2_outputs(3119);
    layer3_outputs(8441) <= layer2_outputs(7977);
    layer3_outputs(8442) <= layer2_outputs(1352);
    layer3_outputs(8443) <= '0';
    layer3_outputs(8444) <= not(layer2_outputs(928));
    layer3_outputs(8445) <= (layer2_outputs(3023)) or (layer2_outputs(8866));
    layer3_outputs(8446) <= not((layer2_outputs(9612)) xor (layer2_outputs(7686)));
    layer3_outputs(8447) <= (layer2_outputs(5490)) or (layer2_outputs(4790));
    layer3_outputs(8448) <= not(layer2_outputs(7307));
    layer3_outputs(8449) <= not(layer2_outputs(7345));
    layer3_outputs(8450) <= not(layer2_outputs(1691));
    layer3_outputs(8451) <= '1';
    layer3_outputs(8452) <= (layer2_outputs(6791)) or (layer2_outputs(3741));
    layer3_outputs(8453) <= layer2_outputs(7866);
    layer3_outputs(8454) <= not((layer2_outputs(5891)) or (layer2_outputs(6016)));
    layer3_outputs(8455) <= '1';
    layer3_outputs(8456) <= layer2_outputs(1937);
    layer3_outputs(8457) <= not(layer2_outputs(3657));
    layer3_outputs(8458) <= (layer2_outputs(8253)) xor (layer2_outputs(1039));
    layer3_outputs(8459) <= layer2_outputs(1436);
    layer3_outputs(8460) <= not(layer2_outputs(5965)) or (layer2_outputs(1275));
    layer3_outputs(8461) <= not((layer2_outputs(325)) or (layer2_outputs(4127)));
    layer3_outputs(8462) <= layer2_outputs(3838);
    layer3_outputs(8463) <= '1';
    layer3_outputs(8464) <= not((layer2_outputs(7211)) or (layer2_outputs(8862)));
    layer3_outputs(8465) <= not(layer2_outputs(6522));
    layer3_outputs(8466) <= (layer2_outputs(7438)) or (layer2_outputs(169));
    layer3_outputs(8467) <= not(layer2_outputs(4342)) or (layer2_outputs(6089));
    layer3_outputs(8468) <= not(layer2_outputs(3136));
    layer3_outputs(8469) <= (layer2_outputs(1585)) and not (layer2_outputs(8460));
    layer3_outputs(8470) <= layer2_outputs(6460);
    layer3_outputs(8471) <= '0';
    layer3_outputs(8472) <= not((layer2_outputs(9800)) or (layer2_outputs(8766)));
    layer3_outputs(8473) <= not(layer2_outputs(8485));
    layer3_outputs(8474) <= not((layer2_outputs(1897)) or (layer2_outputs(9034)));
    layer3_outputs(8475) <= layer2_outputs(8111);
    layer3_outputs(8476) <= (layer2_outputs(6735)) and not (layer2_outputs(4993));
    layer3_outputs(8477) <= not(layer2_outputs(755));
    layer3_outputs(8478) <= not(layer2_outputs(9819));
    layer3_outputs(8479) <= (layer2_outputs(9640)) or (layer2_outputs(3306));
    layer3_outputs(8480) <= (layer2_outputs(6712)) and not (layer2_outputs(7119));
    layer3_outputs(8481) <= (layer2_outputs(5042)) and not (layer2_outputs(9546));
    layer3_outputs(8482) <= not(layer2_outputs(9372));
    layer3_outputs(8483) <= (layer2_outputs(3581)) and not (layer2_outputs(2462));
    layer3_outputs(8484) <= not(layer2_outputs(9316)) or (layer2_outputs(9746));
    layer3_outputs(8485) <= not(layer2_outputs(4873));
    layer3_outputs(8486) <= not((layer2_outputs(8505)) or (layer2_outputs(9950)));
    layer3_outputs(8487) <= layer2_outputs(3623);
    layer3_outputs(8488) <= layer2_outputs(5436);
    layer3_outputs(8489) <= not((layer2_outputs(6274)) and (layer2_outputs(8889)));
    layer3_outputs(8490) <= layer2_outputs(4150);
    layer3_outputs(8491) <= layer2_outputs(8462);
    layer3_outputs(8492) <= layer2_outputs(2518);
    layer3_outputs(8493) <= layer2_outputs(2188);
    layer3_outputs(8494) <= layer2_outputs(7357);
    layer3_outputs(8495) <= not(layer2_outputs(4595));
    layer3_outputs(8496) <= layer2_outputs(5163);
    layer3_outputs(8497) <= (layer2_outputs(1656)) and not (layer2_outputs(6434));
    layer3_outputs(8498) <= (layer2_outputs(5343)) xor (layer2_outputs(7462));
    layer3_outputs(8499) <= (layer2_outputs(8400)) and not (layer2_outputs(5171));
    layer3_outputs(8500) <= layer2_outputs(6989);
    layer3_outputs(8501) <= not(layer2_outputs(8190)) or (layer2_outputs(9878));
    layer3_outputs(8502) <= not((layer2_outputs(3719)) xor (layer2_outputs(6952)));
    layer3_outputs(8503) <= layer2_outputs(7023);
    layer3_outputs(8504) <= (layer2_outputs(2383)) and (layer2_outputs(5396));
    layer3_outputs(8505) <= (layer2_outputs(5515)) or (layer2_outputs(1132));
    layer3_outputs(8506) <= not((layer2_outputs(6731)) or (layer2_outputs(10015)));
    layer3_outputs(8507) <= layer2_outputs(3985);
    layer3_outputs(8508) <= (layer2_outputs(103)) or (layer2_outputs(4607));
    layer3_outputs(8509) <= layer2_outputs(6720);
    layer3_outputs(8510) <= not(layer2_outputs(4449)) or (layer2_outputs(1511));
    layer3_outputs(8511) <= layer2_outputs(6481);
    layer3_outputs(8512) <= not((layer2_outputs(5500)) xor (layer2_outputs(3677)));
    layer3_outputs(8513) <= layer2_outputs(2848);
    layer3_outputs(8514) <= not(layer2_outputs(5145));
    layer3_outputs(8515) <= '1';
    layer3_outputs(8516) <= layer2_outputs(7574);
    layer3_outputs(8517) <= not((layer2_outputs(177)) xor (layer2_outputs(3395)));
    layer3_outputs(8518) <= layer2_outputs(1829);
    layer3_outputs(8519) <= (layer2_outputs(7906)) and (layer2_outputs(9470));
    layer3_outputs(8520) <= (layer2_outputs(475)) xor (layer2_outputs(7829));
    layer3_outputs(8521) <= (layer2_outputs(7765)) and not (layer2_outputs(6461));
    layer3_outputs(8522) <= not(layer2_outputs(8303));
    layer3_outputs(8523) <= layer2_outputs(620);
    layer3_outputs(8524) <= not(layer2_outputs(140));
    layer3_outputs(8525) <= not(layer2_outputs(7646));
    layer3_outputs(8526) <= (layer2_outputs(9543)) and not (layer2_outputs(6620));
    layer3_outputs(8527) <= not((layer2_outputs(905)) and (layer2_outputs(2196)));
    layer3_outputs(8528) <= layer2_outputs(118);
    layer3_outputs(8529) <= not(layer2_outputs(8606)) or (layer2_outputs(2751));
    layer3_outputs(8530) <= layer2_outputs(777);
    layer3_outputs(8531) <= (layer2_outputs(140)) xor (layer2_outputs(1144));
    layer3_outputs(8532) <= (layer2_outputs(10153)) and (layer2_outputs(7363));
    layer3_outputs(8533) <= not((layer2_outputs(10042)) or (layer2_outputs(4907)));
    layer3_outputs(8534) <= layer2_outputs(8077);
    layer3_outputs(8535) <= layer2_outputs(8899);
    layer3_outputs(8536) <= not((layer2_outputs(3819)) and (layer2_outputs(6116)));
    layer3_outputs(8537) <= not(layer2_outputs(4545)) or (layer2_outputs(7684));
    layer3_outputs(8538) <= not(layer2_outputs(2498)) or (layer2_outputs(6149));
    layer3_outputs(8539) <= not(layer2_outputs(5404)) or (layer2_outputs(9483));
    layer3_outputs(8540) <= not(layer2_outputs(3260));
    layer3_outputs(8541) <= '0';
    layer3_outputs(8542) <= not(layer2_outputs(1665)) or (layer2_outputs(8301));
    layer3_outputs(8543) <= not(layer2_outputs(3172));
    layer3_outputs(8544) <= not(layer2_outputs(2057));
    layer3_outputs(8545) <= layer2_outputs(10038);
    layer3_outputs(8546) <= (layer2_outputs(1650)) and not (layer2_outputs(7470));
    layer3_outputs(8547) <= layer2_outputs(3590);
    layer3_outputs(8548) <= not(layer2_outputs(5278));
    layer3_outputs(8549) <= '0';
    layer3_outputs(8550) <= not(layer2_outputs(7103));
    layer3_outputs(8551) <= (layer2_outputs(6590)) and not (layer2_outputs(8333));
    layer3_outputs(8552) <= layer2_outputs(8468);
    layer3_outputs(8553) <= layer2_outputs(2565);
    layer3_outputs(8554) <= not(layer2_outputs(8206)) or (layer2_outputs(4913));
    layer3_outputs(8555) <= (layer2_outputs(9618)) or (layer2_outputs(5809));
    layer3_outputs(8556) <= not(layer2_outputs(9789));
    layer3_outputs(8557) <= not(layer2_outputs(1954));
    layer3_outputs(8558) <= layer2_outputs(7277);
    layer3_outputs(8559) <= (layer2_outputs(8918)) and (layer2_outputs(2132));
    layer3_outputs(8560) <= (layer2_outputs(7460)) and not (layer2_outputs(3018));
    layer3_outputs(8561) <= layer2_outputs(674);
    layer3_outputs(8562) <= layer2_outputs(3651);
    layer3_outputs(8563) <= not(layer2_outputs(7952)) or (layer2_outputs(8195));
    layer3_outputs(8564) <= (layer2_outputs(6861)) and (layer2_outputs(9517));
    layer3_outputs(8565) <= (layer2_outputs(10110)) or (layer2_outputs(2618));
    layer3_outputs(8566) <= not(layer2_outputs(4658)) or (layer2_outputs(10022));
    layer3_outputs(8567) <= (layer2_outputs(4878)) and not (layer2_outputs(8715));
    layer3_outputs(8568) <= (layer2_outputs(797)) and (layer2_outputs(10194));
    layer3_outputs(8569) <= layer2_outputs(3031);
    layer3_outputs(8570) <= layer2_outputs(9222);
    layer3_outputs(8571) <= (layer2_outputs(3984)) and not (layer2_outputs(1655));
    layer3_outputs(8572) <= (layer2_outputs(7246)) and not (layer2_outputs(1658));
    layer3_outputs(8573) <= layer2_outputs(5592);
    layer3_outputs(8574) <= '0';
    layer3_outputs(8575) <= not(layer2_outputs(3263));
    layer3_outputs(8576) <= (layer2_outputs(7072)) and (layer2_outputs(2215));
    layer3_outputs(8577) <= (layer2_outputs(4456)) or (layer2_outputs(2581));
    layer3_outputs(8578) <= layer2_outputs(663);
    layer3_outputs(8579) <= not(layer2_outputs(520)) or (layer2_outputs(7284));
    layer3_outputs(8580) <= layer2_outputs(8778);
    layer3_outputs(8581) <= not((layer2_outputs(4209)) or (layer2_outputs(2287)));
    layer3_outputs(8582) <= not(layer2_outputs(1515));
    layer3_outputs(8583) <= not((layer2_outputs(1289)) xor (layer2_outputs(5628)));
    layer3_outputs(8584) <= layer2_outputs(713);
    layer3_outputs(8585) <= layer2_outputs(4674);
    layer3_outputs(8586) <= not(layer2_outputs(6319));
    layer3_outputs(8587) <= (layer2_outputs(3473)) or (layer2_outputs(9866));
    layer3_outputs(8588) <= not((layer2_outputs(5765)) and (layer2_outputs(3271)));
    layer3_outputs(8589) <= not((layer2_outputs(4308)) xor (layer2_outputs(9730)));
    layer3_outputs(8590) <= layer2_outputs(2186);
    layer3_outputs(8591) <= layer2_outputs(7950);
    layer3_outputs(8592) <= not((layer2_outputs(7140)) xor (layer2_outputs(1898)));
    layer3_outputs(8593) <= not(layer2_outputs(1009));
    layer3_outputs(8594) <= (layer2_outputs(6911)) and (layer2_outputs(991));
    layer3_outputs(8595) <= not((layer2_outputs(2469)) and (layer2_outputs(7368)));
    layer3_outputs(8596) <= not((layer2_outputs(8828)) or (layer2_outputs(10195)));
    layer3_outputs(8597) <= not(layer2_outputs(9100));
    layer3_outputs(8598) <= layer2_outputs(1580);
    layer3_outputs(8599) <= not((layer2_outputs(7647)) and (layer2_outputs(1106)));
    layer3_outputs(8600) <= (layer2_outputs(2661)) or (layer2_outputs(5107));
    layer3_outputs(8601) <= not(layer2_outputs(461));
    layer3_outputs(8602) <= (layer2_outputs(5173)) or (layer2_outputs(2127));
    layer3_outputs(8603) <= layer2_outputs(5483);
    layer3_outputs(8604) <= not(layer2_outputs(5518)) or (layer2_outputs(4111));
    layer3_outputs(8605) <= not(layer2_outputs(5852)) or (layer2_outputs(7266));
    layer3_outputs(8606) <= layer2_outputs(10206);
    layer3_outputs(8607) <= '1';
    layer3_outputs(8608) <= (layer2_outputs(3663)) and (layer2_outputs(6404));
    layer3_outputs(8609) <= layer2_outputs(1513);
    layer3_outputs(8610) <= not((layer2_outputs(2803)) and (layer2_outputs(1364)));
    layer3_outputs(8611) <= not(layer2_outputs(6131));
    layer3_outputs(8612) <= not(layer2_outputs(639)) or (layer2_outputs(8007));
    layer3_outputs(8613) <= layer2_outputs(4941);
    layer3_outputs(8614) <= (layer2_outputs(6144)) or (layer2_outputs(7534));
    layer3_outputs(8615) <= layer2_outputs(1394);
    layer3_outputs(8616) <= layer2_outputs(4809);
    layer3_outputs(8617) <= (layer2_outputs(4302)) xor (layer2_outputs(1293));
    layer3_outputs(8618) <= not((layer2_outputs(3163)) or (layer2_outputs(2817)));
    layer3_outputs(8619) <= (layer2_outputs(3039)) or (layer2_outputs(2394));
    layer3_outputs(8620) <= not(layer2_outputs(6513));
    layer3_outputs(8621) <= not(layer2_outputs(8859));
    layer3_outputs(8622) <= not(layer2_outputs(10214));
    layer3_outputs(8623) <= not(layer2_outputs(3008));
    layer3_outputs(8624) <= (layer2_outputs(4593)) or (layer2_outputs(1827));
    layer3_outputs(8625) <= not((layer2_outputs(3832)) or (layer2_outputs(2765)));
    layer3_outputs(8626) <= layer2_outputs(8426);
    layer3_outputs(8627) <= (layer2_outputs(7791)) or (layer2_outputs(10055));
    layer3_outputs(8628) <= layer2_outputs(1092);
    layer3_outputs(8629) <= (layer2_outputs(8729)) and not (layer2_outputs(8574));
    layer3_outputs(8630) <= layer2_outputs(10081);
    layer3_outputs(8631) <= layer2_outputs(4575);
    layer3_outputs(8632) <= (layer2_outputs(2377)) xor (layer2_outputs(2982));
    layer3_outputs(8633) <= (layer2_outputs(3724)) and not (layer2_outputs(7994));
    layer3_outputs(8634) <= (layer2_outputs(5749)) or (layer2_outputs(4947));
    layer3_outputs(8635) <= (layer2_outputs(1451)) or (layer2_outputs(1756));
    layer3_outputs(8636) <= not(layer2_outputs(1035));
    layer3_outputs(8637) <= layer2_outputs(9548);
    layer3_outputs(8638) <= (layer2_outputs(5081)) and not (layer2_outputs(8193));
    layer3_outputs(8639) <= layer2_outputs(8003);
    layer3_outputs(8640) <= layer2_outputs(3231);
    layer3_outputs(8641) <= layer2_outputs(9196);
    layer3_outputs(8642) <= not((layer2_outputs(4822)) or (layer2_outputs(90)));
    layer3_outputs(8643) <= not((layer2_outputs(7601)) xor (layer2_outputs(3501)));
    layer3_outputs(8644) <= not(layer2_outputs(4177));
    layer3_outputs(8645) <= (layer2_outputs(5756)) and (layer2_outputs(3964));
    layer3_outputs(8646) <= not((layer2_outputs(996)) xor (layer2_outputs(1267)));
    layer3_outputs(8647) <= layer2_outputs(3957);
    layer3_outputs(8648) <= not(layer2_outputs(3734));
    layer3_outputs(8649) <= not(layer2_outputs(4767)) or (layer2_outputs(5751));
    layer3_outputs(8650) <= not(layer2_outputs(4976));
    layer3_outputs(8651) <= layer2_outputs(217);
    layer3_outputs(8652) <= (layer2_outputs(4267)) and not (layer2_outputs(199));
    layer3_outputs(8653) <= layer2_outputs(6187);
    layer3_outputs(8654) <= not((layer2_outputs(9123)) and (layer2_outputs(8611)));
    layer3_outputs(8655) <= not((layer2_outputs(945)) xor (layer2_outputs(3727)));
    layer3_outputs(8656) <= (layer2_outputs(3836)) and (layer2_outputs(4473));
    layer3_outputs(8657) <= not(layer2_outputs(3885));
    layer3_outputs(8658) <= not((layer2_outputs(9559)) and (layer2_outputs(3255)));
    layer3_outputs(8659) <= not((layer2_outputs(4364)) or (layer2_outputs(1560)));
    layer3_outputs(8660) <= not((layer2_outputs(80)) xor (layer2_outputs(645)));
    layer3_outputs(8661) <= not((layer2_outputs(9203)) and (layer2_outputs(5826)));
    layer3_outputs(8662) <= (layer2_outputs(6659)) xor (layer2_outputs(2610));
    layer3_outputs(8663) <= layer2_outputs(9596);
    layer3_outputs(8664) <= not(layer2_outputs(8577));
    layer3_outputs(8665) <= not((layer2_outputs(8013)) or (layer2_outputs(3822)));
    layer3_outputs(8666) <= layer2_outputs(8789);
    layer3_outputs(8667) <= (layer2_outputs(6928)) or (layer2_outputs(8765));
    layer3_outputs(8668) <= not(layer2_outputs(3066));
    layer3_outputs(8669) <= layer2_outputs(7318);
    layer3_outputs(8670) <= not(layer2_outputs(1544));
    layer3_outputs(8671) <= (layer2_outputs(2568)) and not (layer2_outputs(4194));
    layer3_outputs(8672) <= layer2_outputs(7688);
    layer3_outputs(8673) <= not(layer2_outputs(8545)) or (layer2_outputs(9051));
    layer3_outputs(8674) <= not((layer2_outputs(8168)) and (layer2_outputs(989)));
    layer3_outputs(8675) <= (layer2_outputs(9888)) and not (layer2_outputs(9072));
    layer3_outputs(8676) <= layer2_outputs(3566);
    layer3_outputs(8677) <= not(layer2_outputs(2903)) or (layer2_outputs(3038));
    layer3_outputs(8678) <= (layer2_outputs(739)) or (layer2_outputs(9278));
    layer3_outputs(8679) <= (layer2_outputs(4686)) and not (layer2_outputs(195));
    layer3_outputs(8680) <= layer2_outputs(3622);
    layer3_outputs(8681) <= layer2_outputs(9057);
    layer3_outputs(8682) <= not(layer2_outputs(4837));
    layer3_outputs(8683) <= not(layer2_outputs(3176)) or (layer2_outputs(6053));
    layer3_outputs(8684) <= not(layer2_outputs(58)) or (layer2_outputs(9823));
    layer3_outputs(8685) <= not(layer2_outputs(1438));
    layer3_outputs(8686) <= (layer2_outputs(7453)) and not (layer2_outputs(4916));
    layer3_outputs(8687) <= not(layer2_outputs(9294));
    layer3_outputs(8688) <= not(layer2_outputs(7911)) or (layer2_outputs(7586));
    layer3_outputs(8689) <= not(layer2_outputs(6079));
    layer3_outputs(8690) <= (layer2_outputs(6485)) or (layer2_outputs(4381));
    layer3_outputs(8691) <= layer2_outputs(984);
    layer3_outputs(8692) <= layer2_outputs(6035);
    layer3_outputs(8693) <= layer2_outputs(7060);
    layer3_outputs(8694) <= not(layer2_outputs(2080));
    layer3_outputs(8695) <= (layer2_outputs(7660)) and not (layer2_outputs(5450));
    layer3_outputs(8696) <= not(layer2_outputs(7912));
    layer3_outputs(8697) <= not(layer2_outputs(287));
    layer3_outputs(8698) <= layer2_outputs(3486);
    layer3_outputs(8699) <= not(layer2_outputs(8572)) or (layer2_outputs(673));
    layer3_outputs(8700) <= not(layer2_outputs(6275));
    layer3_outputs(8701) <= not(layer2_outputs(170));
    layer3_outputs(8702) <= layer2_outputs(7608);
    layer3_outputs(8703) <= layer2_outputs(906);
    layer3_outputs(8704) <= layer2_outputs(2773);
    layer3_outputs(8705) <= not((layer2_outputs(2491)) xor (layer2_outputs(5368)));
    layer3_outputs(8706) <= not(layer2_outputs(1871));
    layer3_outputs(8707) <= layer2_outputs(1234);
    layer3_outputs(8708) <= (layer2_outputs(4496)) and (layer2_outputs(8470));
    layer3_outputs(8709) <= not(layer2_outputs(1801));
    layer3_outputs(8710) <= layer2_outputs(9045);
    layer3_outputs(8711) <= (layer2_outputs(1235)) xor (layer2_outputs(5982));
    layer3_outputs(8712) <= '1';
    layer3_outputs(8713) <= (layer2_outputs(8584)) xor (layer2_outputs(4455));
    layer3_outputs(8714) <= not(layer2_outputs(3778));
    layer3_outputs(8715) <= not((layer2_outputs(5555)) and (layer2_outputs(9195)));
    layer3_outputs(8716) <= not(layer2_outputs(1073)) or (layer2_outputs(8980));
    layer3_outputs(8717) <= layer2_outputs(4789);
    layer3_outputs(8718) <= not(layer2_outputs(5037));
    layer3_outputs(8719) <= layer2_outputs(4928);
    layer3_outputs(8720) <= not((layer2_outputs(6017)) and (layer2_outputs(8947)));
    layer3_outputs(8721) <= layer2_outputs(9075);
    layer3_outputs(8722) <= not(layer2_outputs(1398));
    layer3_outputs(8723) <= not(layer2_outputs(2583));
    layer3_outputs(8724) <= not((layer2_outputs(7703)) and (layer2_outputs(9699)));
    layer3_outputs(8725) <= not(layer2_outputs(2784));
    layer3_outputs(8726) <= not(layer2_outputs(5126));
    layer3_outputs(8727) <= not(layer2_outputs(3412));
    layer3_outputs(8728) <= layer2_outputs(3256);
    layer3_outputs(8729) <= (layer2_outputs(2860)) and not (layer2_outputs(3551));
    layer3_outputs(8730) <= layer2_outputs(10106);
    layer3_outputs(8731) <= not(layer2_outputs(6129));
    layer3_outputs(8732) <= (layer2_outputs(5533)) and not (layer2_outputs(8780));
    layer3_outputs(8733) <= layer2_outputs(4463);
    layer3_outputs(8734) <= (layer2_outputs(1241)) and not (layer2_outputs(12));
    layer3_outputs(8735) <= layer2_outputs(2892);
    layer3_outputs(8736) <= (layer2_outputs(5772)) and (layer2_outputs(6969));
    layer3_outputs(8737) <= not(layer2_outputs(52)) or (layer2_outputs(3570));
    layer3_outputs(8738) <= not((layer2_outputs(5219)) xor (layer2_outputs(4017)));
    layer3_outputs(8739) <= '0';
    layer3_outputs(8740) <= (layer2_outputs(3742)) xor (layer2_outputs(7905));
    layer3_outputs(8741) <= not(layer2_outputs(4313));
    layer3_outputs(8742) <= layer2_outputs(8371);
    layer3_outputs(8743) <= not(layer2_outputs(9219)) or (layer2_outputs(939));
    layer3_outputs(8744) <= (layer2_outputs(7484)) and (layer2_outputs(1176));
    layer3_outputs(8745) <= (layer2_outputs(9271)) or (layer2_outputs(1431));
    layer3_outputs(8746) <= (layer2_outputs(62)) and (layer2_outputs(2908));
    layer3_outputs(8747) <= (layer2_outputs(3725)) or (layer2_outputs(5052));
    layer3_outputs(8748) <= not(layer2_outputs(8937));
    layer3_outputs(8749) <= (layer2_outputs(6608)) and not (layer2_outputs(6346));
    layer3_outputs(8750) <= not(layer2_outputs(3516));
    layer3_outputs(8751) <= layer2_outputs(1356);
    layer3_outputs(8752) <= '1';
    layer3_outputs(8753) <= layer2_outputs(7348);
    layer3_outputs(8754) <= not((layer2_outputs(6395)) xor (layer2_outputs(6537)));
    layer3_outputs(8755) <= layer2_outputs(7725);
    layer3_outputs(8756) <= not(layer2_outputs(2582));
    layer3_outputs(8757) <= (layer2_outputs(4833)) xor (layer2_outputs(370));
    layer3_outputs(8758) <= layer2_outputs(5761);
    layer3_outputs(8759) <= not((layer2_outputs(4575)) xor (layer2_outputs(7311)));
    layer3_outputs(8760) <= not(layer2_outputs(3291));
    layer3_outputs(8761) <= layer2_outputs(5592);
    layer3_outputs(8762) <= not((layer2_outputs(262)) xor (layer2_outputs(6779)));
    layer3_outputs(8763) <= layer2_outputs(8585);
    layer3_outputs(8764) <= (layer2_outputs(10236)) and not (layer2_outputs(3838));
    layer3_outputs(8765) <= layer2_outputs(935);
    layer3_outputs(8766) <= (layer2_outputs(4533)) xor (layer2_outputs(3937));
    layer3_outputs(8767) <= layer2_outputs(9186);
    layer3_outputs(8768) <= not((layer2_outputs(3461)) xor (layer2_outputs(5152)));
    layer3_outputs(8769) <= not((layer2_outputs(1814)) and (layer2_outputs(813)));
    layer3_outputs(8770) <= (layer2_outputs(5135)) xor (layer2_outputs(1770));
    layer3_outputs(8771) <= not(layer2_outputs(5115)) or (layer2_outputs(6377));
    layer3_outputs(8772) <= (layer2_outputs(7372)) and not (layer2_outputs(6711));
    layer3_outputs(8773) <= layer2_outputs(1017);
    layer3_outputs(8774) <= not(layer2_outputs(1854));
    layer3_outputs(8775) <= (layer2_outputs(8639)) xor (layer2_outputs(2700));
    layer3_outputs(8776) <= not(layer2_outputs(8690));
    layer3_outputs(8777) <= (layer2_outputs(3174)) or (layer2_outputs(5755));
    layer3_outputs(8778) <= not(layer2_outputs(3598));
    layer3_outputs(8779) <= (layer2_outputs(9627)) and (layer2_outputs(5136));
    layer3_outputs(8780) <= not((layer2_outputs(5531)) or (layer2_outputs(5249)));
    layer3_outputs(8781) <= not((layer2_outputs(6493)) and (layer2_outputs(6054)));
    layer3_outputs(8782) <= (layer2_outputs(5995)) and not (layer2_outputs(2007));
    layer3_outputs(8783) <= (layer2_outputs(5901)) and (layer2_outputs(6507));
    layer3_outputs(8784) <= (layer2_outputs(1909)) and not (layer2_outputs(6821));
    layer3_outputs(8785) <= layer2_outputs(278);
    layer3_outputs(8786) <= not((layer2_outputs(864)) and (layer2_outputs(4150)));
    layer3_outputs(8787) <= not(layer2_outputs(1612)) or (layer2_outputs(4108));
    layer3_outputs(8788) <= '0';
    layer3_outputs(8789) <= not((layer2_outputs(6754)) and (layer2_outputs(8929)));
    layer3_outputs(8790) <= layer2_outputs(7442);
    layer3_outputs(8791) <= layer2_outputs(1109);
    layer3_outputs(8792) <= not((layer2_outputs(2891)) or (layer2_outputs(8411)));
    layer3_outputs(8793) <= layer2_outputs(4419);
    layer3_outputs(8794) <= layer2_outputs(4641);
    layer3_outputs(8795) <= (layer2_outputs(7239)) xor (layer2_outputs(1332));
    layer3_outputs(8796) <= layer2_outputs(560);
    layer3_outputs(8797) <= layer2_outputs(7287);
    layer3_outputs(8798) <= not(layer2_outputs(311));
    layer3_outputs(8799) <= not(layer2_outputs(9853));
    layer3_outputs(8800) <= not(layer2_outputs(8834));
    layer3_outputs(8801) <= not((layer2_outputs(220)) and (layer2_outputs(428)));
    layer3_outputs(8802) <= (layer2_outputs(8015)) and (layer2_outputs(6462));
    layer3_outputs(8803) <= not((layer2_outputs(2272)) xor (layer2_outputs(4434)));
    layer3_outputs(8804) <= layer2_outputs(7196);
    layer3_outputs(8805) <= not(layer2_outputs(9363));
    layer3_outputs(8806) <= not(layer2_outputs(8));
    layer3_outputs(8807) <= layer2_outputs(3934);
    layer3_outputs(8808) <= (layer2_outputs(3269)) xor (layer2_outputs(6062));
    layer3_outputs(8809) <= (layer2_outputs(2572)) and not (layer2_outputs(2908));
    layer3_outputs(8810) <= not(layer2_outputs(2957));
    layer3_outputs(8811) <= '0';
    layer3_outputs(8812) <= not(layer2_outputs(2560));
    layer3_outputs(8813) <= not(layer2_outputs(2744));
    layer3_outputs(8814) <= not((layer2_outputs(3084)) or (layer2_outputs(2587)));
    layer3_outputs(8815) <= (layer2_outputs(7125)) and not (layer2_outputs(8529));
    layer3_outputs(8816) <= layer2_outputs(6582);
    layer3_outputs(8817) <= layer2_outputs(5989);
    layer3_outputs(8818) <= not(layer2_outputs(1159)) or (layer2_outputs(1817));
    layer3_outputs(8819) <= (layer2_outputs(7218)) and (layer2_outputs(6293));
    layer3_outputs(8820) <= (layer2_outputs(2436)) and not (layer2_outputs(1042));
    layer3_outputs(8821) <= not(layer2_outputs(8579)) or (layer2_outputs(2554));
    layer3_outputs(8822) <= not((layer2_outputs(7891)) and (layer2_outputs(2533)));
    layer3_outputs(8823) <= not(layer2_outputs(1201));
    layer3_outputs(8824) <= layer2_outputs(6072);
    layer3_outputs(8825) <= not(layer2_outputs(10225)) or (layer2_outputs(5687));
    layer3_outputs(8826) <= not(layer2_outputs(8704)) or (layer2_outputs(4196));
    layer3_outputs(8827) <= not(layer2_outputs(9137));
    layer3_outputs(8828) <= not((layer2_outputs(2312)) xor (layer2_outputs(8018)));
    layer3_outputs(8829) <= not(layer2_outputs(3715)) or (layer2_outputs(8339));
    layer3_outputs(8830) <= not(layer2_outputs(1536)) or (layer2_outputs(5989));
    layer3_outputs(8831) <= layer2_outputs(3356);
    layer3_outputs(8832) <= '0';
    layer3_outputs(8833) <= not(layer2_outputs(9478));
    layer3_outputs(8834) <= (layer2_outputs(6064)) and (layer2_outputs(2632));
    layer3_outputs(8835) <= (layer2_outputs(1324)) and not (layer2_outputs(4901));
    layer3_outputs(8836) <= (layer2_outputs(4214)) and not (layer2_outputs(8725));
    layer3_outputs(8837) <= layer2_outputs(4204);
    layer3_outputs(8838) <= layer2_outputs(10111);
    layer3_outputs(8839) <= layer2_outputs(6704);
    layer3_outputs(8840) <= not(layer2_outputs(5347));
    layer3_outputs(8841) <= (layer2_outputs(1636)) and not (layer2_outputs(7117));
    layer3_outputs(8842) <= (layer2_outputs(2674)) and (layer2_outputs(9871));
    layer3_outputs(8843) <= layer2_outputs(5600);
    layer3_outputs(8844) <= not(layer2_outputs(538));
    layer3_outputs(8845) <= (layer2_outputs(8650)) xor (layer2_outputs(9551));
    layer3_outputs(8846) <= layer2_outputs(3965);
    layer3_outputs(8847) <= not((layer2_outputs(4516)) and (layer2_outputs(1263)));
    layer3_outputs(8848) <= not(layer2_outputs(7144)) or (layer2_outputs(8393));
    layer3_outputs(8849) <= not(layer2_outputs(9839));
    layer3_outputs(8850) <= not(layer2_outputs(6719));
    layer3_outputs(8851) <= not(layer2_outputs(1627));
    layer3_outputs(8852) <= not(layer2_outputs(2271));
    layer3_outputs(8853) <= (layer2_outputs(8722)) and (layer2_outputs(5270));
    layer3_outputs(8854) <= not(layer2_outputs(8478));
    layer3_outputs(8855) <= layer2_outputs(2048);
    layer3_outputs(8856) <= not(layer2_outputs(4220));
    layer3_outputs(8857) <= layer2_outputs(7151);
    layer3_outputs(8858) <= not(layer2_outputs(7932));
    layer3_outputs(8859) <= not(layer2_outputs(6040));
    layer3_outputs(8860) <= (layer2_outputs(7763)) or (layer2_outputs(5756));
    layer3_outputs(8861) <= not(layer2_outputs(7743));
    layer3_outputs(8862) <= not(layer2_outputs(7568));
    layer3_outputs(8863) <= '1';
    layer3_outputs(8864) <= (layer2_outputs(7476)) or (layer2_outputs(5571));
    layer3_outputs(8865) <= not((layer2_outputs(9037)) or (layer2_outputs(7771)));
    layer3_outputs(8866) <= (layer2_outputs(439)) or (layer2_outputs(5273));
    layer3_outputs(8867) <= (layer2_outputs(4347)) and not (layer2_outputs(1242));
    layer3_outputs(8868) <= not((layer2_outputs(9694)) or (layer2_outputs(2004)));
    layer3_outputs(8869) <= not(layer2_outputs(1873));
    layer3_outputs(8870) <= not(layer2_outputs(5753));
    layer3_outputs(8871) <= not(layer2_outputs(795));
    layer3_outputs(8872) <= layer2_outputs(4793);
    layer3_outputs(8873) <= (layer2_outputs(4922)) xor (layer2_outputs(8761));
    layer3_outputs(8874) <= not(layer2_outputs(6090)) or (layer2_outputs(5433));
    layer3_outputs(8875) <= (layer2_outputs(7803)) and not (layer2_outputs(3852));
    layer3_outputs(8876) <= layer2_outputs(6292);
    layer3_outputs(8877) <= not((layer2_outputs(8667)) xor (layer2_outputs(4710)));
    layer3_outputs(8878) <= layer2_outputs(8900);
    layer3_outputs(8879) <= layer2_outputs(9192);
    layer3_outputs(8880) <= layer2_outputs(6799);
    layer3_outputs(8881) <= layer2_outputs(7261);
    layer3_outputs(8882) <= (layer2_outputs(6357)) and not (layer2_outputs(4584));
    layer3_outputs(8883) <= not((layer2_outputs(5538)) xor (layer2_outputs(5134)));
    layer3_outputs(8884) <= not(layer2_outputs(2221));
    layer3_outputs(8885) <= not((layer2_outputs(355)) xor (layer2_outputs(324)));
    layer3_outputs(8886) <= not((layer2_outputs(5148)) or (layer2_outputs(5097)));
    layer3_outputs(8887) <= layer2_outputs(4701);
    layer3_outputs(8888) <= layer2_outputs(8056);
    layer3_outputs(8889) <= (layer2_outputs(2741)) and not (layer2_outputs(7461));
    layer3_outputs(8890) <= not((layer2_outputs(6275)) or (layer2_outputs(3738)));
    layer3_outputs(8891) <= not(layer2_outputs(10164)) or (layer2_outputs(2624));
    layer3_outputs(8892) <= not(layer2_outputs(6363));
    layer3_outputs(8893) <= (layer2_outputs(1305)) or (layer2_outputs(6473));
    layer3_outputs(8894) <= (layer2_outputs(8191)) and (layer2_outputs(5966));
    layer3_outputs(8895) <= not(layer2_outputs(6779));
    layer3_outputs(8896) <= not(layer2_outputs(5629));
    layer3_outputs(8897) <= layer2_outputs(2770);
    layer3_outputs(8898) <= (layer2_outputs(2198)) and (layer2_outputs(9505));
    layer3_outputs(8899) <= '0';
    layer3_outputs(8900) <= (layer2_outputs(562)) xor (layer2_outputs(5034));
    layer3_outputs(8901) <= (layer2_outputs(672)) and not (layer2_outputs(2169));
    layer3_outputs(8902) <= not(layer2_outputs(420)) or (layer2_outputs(8356));
    layer3_outputs(8903) <= '1';
    layer3_outputs(8904) <= not(layer2_outputs(9653));
    layer3_outputs(8905) <= not((layer2_outputs(426)) xor (layer2_outputs(9737)));
    layer3_outputs(8906) <= not(layer2_outputs(3397));
    layer3_outputs(8907) <= (layer2_outputs(2843)) and (layer2_outputs(1807));
    layer3_outputs(8908) <= not((layer2_outputs(4143)) or (layer2_outputs(4505)));
    layer3_outputs(8909) <= layer2_outputs(8901);
    layer3_outputs(8910) <= layer2_outputs(7855);
    layer3_outputs(8911) <= layer2_outputs(7174);
    layer3_outputs(8912) <= (layer2_outputs(1923)) or (layer2_outputs(4862));
    layer3_outputs(8913) <= layer2_outputs(1868);
    layer3_outputs(8914) <= (layer2_outputs(1331)) and not (layer2_outputs(3626));
    layer3_outputs(8915) <= not(layer2_outputs(6147));
    layer3_outputs(8916) <= not(layer2_outputs(2329));
    layer3_outputs(8917) <= layer2_outputs(4261);
    layer3_outputs(8918) <= layer2_outputs(1472);
    layer3_outputs(8919) <= (layer2_outputs(897)) and (layer2_outputs(2536));
    layer3_outputs(8920) <= not(layer2_outputs(5258));
    layer3_outputs(8921) <= not(layer2_outputs(205));
    layer3_outputs(8922) <= not((layer2_outputs(9691)) xor (layer2_outputs(264)));
    layer3_outputs(8923) <= layer2_outputs(3627);
    layer3_outputs(8924) <= not((layer2_outputs(3860)) and (layer2_outputs(2894)));
    layer3_outputs(8925) <= (layer2_outputs(5267)) and not (layer2_outputs(2337));
    layer3_outputs(8926) <= (layer2_outputs(5842)) xor (layer2_outputs(949));
    layer3_outputs(8927) <= not((layer2_outputs(5088)) and (layer2_outputs(3462)));
    layer3_outputs(8928) <= (layer2_outputs(2274)) or (layer2_outputs(8589));
    layer3_outputs(8929) <= (layer2_outputs(4225)) xor (layer2_outputs(3751));
    layer3_outputs(8930) <= not(layer2_outputs(2320)) or (layer2_outputs(5885));
    layer3_outputs(8931) <= not(layer2_outputs(1240));
    layer3_outputs(8932) <= not(layer2_outputs(8307));
    layer3_outputs(8933) <= '1';
    layer3_outputs(8934) <= not(layer2_outputs(6128));
    layer3_outputs(8935) <= not(layer2_outputs(274));
    layer3_outputs(8936) <= (layer2_outputs(1217)) and not (layer2_outputs(6265));
    layer3_outputs(8937) <= layer2_outputs(2329);
    layer3_outputs(8938) <= not(layer2_outputs(806));
    layer3_outputs(8939) <= not(layer2_outputs(6134));
    layer3_outputs(8940) <= (layer2_outputs(130)) or (layer2_outputs(6305));
    layer3_outputs(8941) <= layer2_outputs(6385);
    layer3_outputs(8942) <= not(layer2_outputs(6949));
    layer3_outputs(8943) <= not((layer2_outputs(3326)) xor (layer2_outputs(3653)));
    layer3_outputs(8944) <= not(layer2_outputs(2022)) or (layer2_outputs(7501));
    layer3_outputs(8945) <= layer2_outputs(2109);
    layer3_outputs(8946) <= layer2_outputs(100);
    layer3_outputs(8947) <= (layer2_outputs(2062)) and not (layer2_outputs(9526));
    layer3_outputs(8948) <= not(layer2_outputs(296));
    layer3_outputs(8949) <= layer2_outputs(7974);
    layer3_outputs(8950) <= not((layer2_outputs(4184)) or (layer2_outputs(4771)));
    layer3_outputs(8951) <= not(layer2_outputs(216));
    layer3_outputs(8952) <= (layer2_outputs(3947)) or (layer2_outputs(797));
    layer3_outputs(8953) <= not(layer2_outputs(9112)) or (layer2_outputs(2223));
    layer3_outputs(8954) <= (layer2_outputs(1198)) or (layer2_outputs(5320));
    layer3_outputs(8955) <= (layer2_outputs(1449)) xor (layer2_outputs(7725));
    layer3_outputs(8956) <= layer2_outputs(5870);
    layer3_outputs(8957) <= (layer2_outputs(5491)) and not (layer2_outputs(7477));
    layer3_outputs(8958) <= not(layer2_outputs(2557));
    layer3_outputs(8959) <= layer2_outputs(170);
    layer3_outputs(8960) <= not((layer2_outputs(7511)) and (layer2_outputs(257)));
    layer3_outputs(8961) <= (layer2_outputs(2953)) and not (layer2_outputs(6066));
    layer3_outputs(8962) <= (layer2_outputs(546)) and not (layer2_outputs(365));
    layer3_outputs(8963) <= not(layer2_outputs(3523));
    layer3_outputs(8964) <= not(layer2_outputs(4062));
    layer3_outputs(8965) <= (layer2_outputs(208)) xor (layer2_outputs(7656));
    layer3_outputs(8966) <= not(layer2_outputs(7943)) or (layer2_outputs(1719));
    layer3_outputs(8967) <= not(layer2_outputs(2439)) or (layer2_outputs(1274));
    layer3_outputs(8968) <= (layer2_outputs(5275)) and (layer2_outputs(8883));
    layer3_outputs(8969) <= '1';
    layer3_outputs(8970) <= layer2_outputs(2442);
    layer3_outputs(8971) <= not(layer2_outputs(2646)) or (layer2_outputs(3641));
    layer3_outputs(8972) <= (layer2_outputs(5538)) xor (layer2_outputs(9398));
    layer3_outputs(8973) <= not((layer2_outputs(5372)) xor (layer2_outputs(9830)));
    layer3_outputs(8974) <= layer2_outputs(2824);
    layer3_outputs(8975) <= not((layer2_outputs(6931)) and (layer2_outputs(1381)));
    layer3_outputs(8976) <= not(layer2_outputs(4407));
    layer3_outputs(8977) <= not(layer2_outputs(9648)) or (layer2_outputs(7097));
    layer3_outputs(8978) <= not(layer2_outputs(10109)) or (layer2_outputs(3377));
    layer3_outputs(8979) <= layer2_outputs(6410);
    layer3_outputs(8980) <= (layer2_outputs(4911)) and not (layer2_outputs(3994));
    layer3_outputs(8981) <= (layer2_outputs(10065)) and not (layer2_outputs(4554));
    layer3_outputs(8982) <= (layer2_outputs(8899)) and not (layer2_outputs(9602));
    layer3_outputs(8983) <= (layer2_outputs(9866)) and (layer2_outputs(2209));
    layer3_outputs(8984) <= not(layer2_outputs(2369));
    layer3_outputs(8985) <= not((layer2_outputs(8738)) and (layer2_outputs(8649)));
    layer3_outputs(8986) <= layer2_outputs(894);
    layer3_outputs(8987) <= (layer2_outputs(2729)) and (layer2_outputs(1336));
    layer3_outputs(8988) <= not((layer2_outputs(6917)) and (layer2_outputs(1280)));
    layer3_outputs(8989) <= not(layer2_outputs(10224));
    layer3_outputs(8990) <= not(layer2_outputs(1));
    layer3_outputs(8991) <= (layer2_outputs(1286)) xor (layer2_outputs(9088));
    layer3_outputs(8992) <= (layer2_outputs(6005)) and not (layer2_outputs(9070));
    layer3_outputs(8993) <= layer2_outputs(7873);
    layer3_outputs(8994) <= layer2_outputs(3323);
    layer3_outputs(8995) <= not((layer2_outputs(3894)) and (layer2_outputs(3185)));
    layer3_outputs(8996) <= layer2_outputs(5308);
    layer3_outputs(8997) <= layer2_outputs(5779);
    layer3_outputs(8998) <= not((layer2_outputs(8738)) and (layer2_outputs(9176)));
    layer3_outputs(8999) <= not((layer2_outputs(9039)) xor (layer2_outputs(1886)));
    layer3_outputs(9000) <= layer2_outputs(3341);
    layer3_outputs(9001) <= not(layer2_outputs(5198)) or (layer2_outputs(2217));
    layer3_outputs(9002) <= not(layer2_outputs(5413)) or (layer2_outputs(3681));
    layer3_outputs(9003) <= (layer2_outputs(981)) and not (layer2_outputs(4772));
    layer3_outputs(9004) <= not(layer2_outputs(6653));
    layer3_outputs(9005) <= layer2_outputs(3524);
    layer3_outputs(9006) <= layer2_outputs(7731);
    layer3_outputs(9007) <= (layer2_outputs(2552)) and not (layer2_outputs(558));
    layer3_outputs(9008) <= not(layer2_outputs(6673));
    layer3_outputs(9009) <= layer2_outputs(10083);
    layer3_outputs(9010) <= not(layer2_outputs(9587));
    layer3_outputs(9011) <= layer2_outputs(5022);
    layer3_outputs(9012) <= (layer2_outputs(2541)) and not (layer2_outputs(5530));
    layer3_outputs(9013) <= layer2_outputs(396);
    layer3_outputs(9014) <= (layer2_outputs(9351)) and not (layer2_outputs(3733));
    layer3_outputs(9015) <= not(layer2_outputs(4635));
    layer3_outputs(9016) <= layer2_outputs(9094);
    layer3_outputs(9017) <= not(layer2_outputs(3927));
    layer3_outputs(9018) <= (layer2_outputs(9921)) and not (layer2_outputs(8220));
    layer3_outputs(9019) <= not(layer2_outputs(6669));
    layer3_outputs(9020) <= (layer2_outputs(5588)) or (layer2_outputs(1972));
    layer3_outputs(9021) <= (layer2_outputs(2355)) and not (layer2_outputs(10203));
    layer3_outputs(9022) <= not((layer2_outputs(3130)) xor (layer2_outputs(10042)));
    layer3_outputs(9023) <= (layer2_outputs(599)) and not (layer2_outputs(8650));
    layer3_outputs(9024) <= layer2_outputs(9250);
    layer3_outputs(9025) <= (layer2_outputs(2346)) or (layer2_outputs(6338));
    layer3_outputs(9026) <= not(layer2_outputs(4604));
    layer3_outputs(9027) <= not((layer2_outputs(3205)) and (layer2_outputs(9716)));
    layer3_outputs(9028) <= not(layer2_outputs(8805));
    layer3_outputs(9029) <= not((layer2_outputs(6596)) or (layer2_outputs(15)));
    layer3_outputs(9030) <= not(layer2_outputs(346)) or (layer2_outputs(5008));
    layer3_outputs(9031) <= (layer2_outputs(3023)) and (layer2_outputs(200));
    layer3_outputs(9032) <= layer2_outputs(6849);
    layer3_outputs(9033) <= not(layer2_outputs(5623));
    layer3_outputs(9034) <= '1';
    layer3_outputs(9035) <= (layer2_outputs(6936)) or (layer2_outputs(7766));
    layer3_outputs(9036) <= layer2_outputs(1591);
    layer3_outputs(9037) <= not(layer2_outputs(6875));
    layer3_outputs(9038) <= not((layer2_outputs(8409)) and (layer2_outputs(6741)));
    layer3_outputs(9039) <= (layer2_outputs(1897)) xor (layer2_outputs(9044));
    layer3_outputs(9040) <= not(layer2_outputs(5020));
    layer3_outputs(9041) <= not((layer2_outputs(2042)) or (layer2_outputs(1904)));
    layer3_outputs(9042) <= not((layer2_outputs(9837)) xor (layer2_outputs(2911)));
    layer3_outputs(9043) <= not(layer2_outputs(3129));
    layer3_outputs(9044) <= layer2_outputs(4322);
    layer3_outputs(9045) <= (layer2_outputs(4855)) or (layer2_outputs(3682));
    layer3_outputs(9046) <= layer2_outputs(3697);
    layer3_outputs(9047) <= not(layer2_outputs(6952));
    layer3_outputs(9048) <= (layer2_outputs(1092)) and (layer2_outputs(4233));
    layer3_outputs(9049) <= (layer2_outputs(7005)) or (layer2_outputs(6905));
    layer3_outputs(9050) <= layer2_outputs(9676);
    layer3_outputs(9051) <= layer2_outputs(6039);
    layer3_outputs(9052) <= layer2_outputs(6171);
    layer3_outputs(9053) <= not(layer2_outputs(3540));
    layer3_outputs(9054) <= not(layer2_outputs(8577)) or (layer2_outputs(2558));
    layer3_outputs(9055) <= layer2_outputs(9429);
    layer3_outputs(9056) <= not(layer2_outputs(9231));
    layer3_outputs(9057) <= (layer2_outputs(799)) or (layer2_outputs(1942));
    layer3_outputs(9058) <= not(layer2_outputs(4362)) or (layer2_outputs(3945));
    layer3_outputs(9059) <= not(layer2_outputs(729));
    layer3_outputs(9060) <= (layer2_outputs(9805)) xor (layer2_outputs(2044));
    layer3_outputs(9061) <= layer2_outputs(4573);
    layer3_outputs(9062) <= not(layer2_outputs(7886));
    layer3_outputs(9063) <= (layer2_outputs(7878)) or (layer2_outputs(5622));
    layer3_outputs(9064) <= not((layer2_outputs(4020)) and (layer2_outputs(3661)));
    layer3_outputs(9065) <= layer2_outputs(6394);
    layer3_outputs(9066) <= not(layer2_outputs(5734)) or (layer2_outputs(6953));
    layer3_outputs(9067) <= (layer2_outputs(2262)) and (layer2_outputs(940));
    layer3_outputs(9068) <= layer2_outputs(1492);
    layer3_outputs(9069) <= (layer2_outputs(7472)) or (layer2_outputs(6217));
    layer3_outputs(9070) <= (layer2_outputs(1873)) or (layer2_outputs(2084));
    layer3_outputs(9071) <= layer2_outputs(8036);
    layer3_outputs(9072) <= not(layer2_outputs(3481));
    layer3_outputs(9073) <= not(layer2_outputs(2556));
    layer3_outputs(9074) <= not(layer2_outputs(4698));
    layer3_outputs(9075) <= (layer2_outputs(1440)) xor (layer2_outputs(1719));
    layer3_outputs(9076) <= not((layer2_outputs(7565)) xor (layer2_outputs(5651)));
    layer3_outputs(9077) <= not((layer2_outputs(8006)) or (layer2_outputs(5491)));
    layer3_outputs(9078) <= not((layer2_outputs(6606)) xor (layer2_outputs(3974)));
    layer3_outputs(9079) <= layer2_outputs(3921);
    layer3_outputs(9080) <= (layer2_outputs(6983)) and not (layer2_outputs(4799));
    layer3_outputs(9081) <= not(layer2_outputs(7284)) or (layer2_outputs(8983));
    layer3_outputs(9082) <= not(layer2_outputs(2408));
    layer3_outputs(9083) <= (layer2_outputs(5645)) or (layer2_outputs(8518));
    layer3_outputs(9084) <= not(layer2_outputs(10222)) or (layer2_outputs(2175));
    layer3_outputs(9085) <= '0';
    layer3_outputs(9086) <= (layer2_outputs(899)) and (layer2_outputs(4758));
    layer3_outputs(9087) <= not((layer2_outputs(1883)) or (layer2_outputs(1244)));
    layer3_outputs(9088) <= (layer2_outputs(2543)) and not (layer2_outputs(4915));
    layer3_outputs(9089) <= not(layer2_outputs(3003));
    layer3_outputs(9090) <= not(layer2_outputs(1701));
    layer3_outputs(9091) <= (layer2_outputs(4624)) and not (layer2_outputs(8137));
    layer3_outputs(9092) <= not(layer2_outputs(7481));
    layer3_outputs(9093) <= (layer2_outputs(8407)) xor (layer2_outputs(1383));
    layer3_outputs(9094) <= layer2_outputs(2251);
    layer3_outputs(9095) <= not(layer2_outputs(1071));
    layer3_outputs(9096) <= '0';
    layer3_outputs(9097) <= not(layer2_outputs(9718));
    layer3_outputs(9098) <= not((layer2_outputs(9529)) and (layer2_outputs(1930)));
    layer3_outputs(9099) <= (layer2_outputs(881)) and (layer2_outputs(2978));
    layer3_outputs(9100) <= not(layer2_outputs(57));
    layer3_outputs(9101) <= (layer2_outputs(1878)) and (layer2_outputs(5462));
    layer3_outputs(9102) <= layer2_outputs(9952);
    layer3_outputs(9103) <= (layer2_outputs(112)) and not (layer2_outputs(225));
    layer3_outputs(9104) <= '1';
    layer3_outputs(9105) <= layer2_outputs(150);
    layer3_outputs(9106) <= not(layer2_outputs(657));
    layer3_outputs(9107) <= not((layer2_outputs(2492)) and (layer2_outputs(997)));
    layer3_outputs(9108) <= (layer2_outputs(5089)) or (layer2_outputs(2692));
    layer3_outputs(9109) <= not(layer2_outputs(9996));
    layer3_outputs(9110) <= not((layer2_outputs(9406)) or (layer2_outputs(9210)));
    layer3_outputs(9111) <= not(layer2_outputs(8839));
    layer3_outputs(9112) <= not((layer2_outputs(9398)) or (layer2_outputs(5035)));
    layer3_outputs(9113) <= not(layer2_outputs(6409));
    layer3_outputs(9114) <= not((layer2_outputs(4963)) and (layer2_outputs(3117)));
    layer3_outputs(9115) <= not(layer2_outputs(4956));
    layer3_outputs(9116) <= not((layer2_outputs(7179)) or (layer2_outputs(4551)));
    layer3_outputs(9117) <= not(layer2_outputs(8981));
    layer3_outputs(9118) <= not(layer2_outputs(2441));
    layer3_outputs(9119) <= layer2_outputs(5403);
    layer3_outputs(9120) <= '0';
    layer3_outputs(9121) <= (layer2_outputs(9961)) and (layer2_outputs(8154));
    layer3_outputs(9122) <= layer2_outputs(7644);
    layer3_outputs(9123) <= not(layer2_outputs(5432));
    layer3_outputs(9124) <= not(layer2_outputs(4219)) or (layer2_outputs(7121));
    layer3_outputs(9125) <= not((layer2_outputs(4200)) and (layer2_outputs(6996)));
    layer3_outputs(9126) <= not(layer2_outputs(769));
    layer3_outputs(9127) <= not((layer2_outputs(6663)) or (layer2_outputs(9671)));
    layer3_outputs(9128) <= (layer2_outputs(9310)) and (layer2_outputs(1404));
    layer3_outputs(9129) <= (layer2_outputs(7423)) or (layer2_outputs(9253));
    layer3_outputs(9130) <= not(layer2_outputs(5787));
    layer3_outputs(9131) <= layer2_outputs(687);
    layer3_outputs(9132) <= not(layer2_outputs(1575)) or (layer2_outputs(2041));
    layer3_outputs(9133) <= layer2_outputs(4450);
    layer3_outputs(9134) <= (layer2_outputs(8805)) and (layer2_outputs(4442));
    layer3_outputs(9135) <= not((layer2_outputs(9099)) or (layer2_outputs(1102)));
    layer3_outputs(9136) <= not(layer2_outputs(276)) or (layer2_outputs(4265));
    layer3_outputs(9137) <= not((layer2_outputs(4971)) and (layer2_outputs(9638)));
    layer3_outputs(9138) <= not(layer2_outputs(2880)) or (layer2_outputs(7327));
    layer3_outputs(9139) <= not(layer2_outputs(9017));
    layer3_outputs(9140) <= not((layer2_outputs(6654)) and (layer2_outputs(1386)));
    layer3_outputs(9141) <= (layer2_outputs(1710)) and not (layer2_outputs(9217));
    layer3_outputs(9142) <= not(layer2_outputs(811));
    layer3_outputs(9143) <= not(layer2_outputs(9223));
    layer3_outputs(9144) <= not(layer2_outputs(9202));
    layer3_outputs(9145) <= layer2_outputs(6491);
    layer3_outputs(9146) <= (layer2_outputs(8224)) or (layer2_outputs(618));
    layer3_outputs(9147) <= '1';
    layer3_outputs(9148) <= not((layer2_outputs(1283)) xor (layer2_outputs(9322)));
    layer3_outputs(9149) <= layer2_outputs(63);
    layer3_outputs(9150) <= layer2_outputs(8620);
    layer3_outputs(9151) <= not(layer2_outputs(8212));
    layer3_outputs(9152) <= not((layer2_outputs(2702)) xor (layer2_outputs(6311)));
    layer3_outputs(9153) <= (layer2_outputs(6856)) and not (layer2_outputs(9480));
    layer3_outputs(9154) <= not((layer2_outputs(2835)) or (layer2_outputs(4494)));
    layer3_outputs(9155) <= (layer2_outputs(7235)) xor (layer2_outputs(742));
    layer3_outputs(9156) <= layer2_outputs(271);
    layer3_outputs(9157) <= (layer2_outputs(1171)) and not (layer2_outputs(6517));
    layer3_outputs(9158) <= not(layer2_outputs(5694));
    layer3_outputs(9159) <= (layer2_outputs(7870)) xor (layer2_outputs(1278));
    layer3_outputs(9160) <= '1';
    layer3_outputs(9161) <= (layer2_outputs(4068)) xor (layer2_outputs(9177));
    layer3_outputs(9162) <= (layer2_outputs(4804)) and not (layer2_outputs(7513));
    layer3_outputs(9163) <= layer2_outputs(122);
    layer3_outputs(9164) <= (layer2_outputs(2624)) and not (layer2_outputs(7001));
    layer3_outputs(9165) <= layer2_outputs(7557);
    layer3_outputs(9166) <= (layer2_outputs(9481)) or (layer2_outputs(9999));
    layer3_outputs(9167) <= layer2_outputs(3007);
    layer3_outputs(9168) <= layer2_outputs(7378);
    layer3_outputs(9169) <= (layer2_outputs(579)) or (layer2_outputs(3514));
    layer3_outputs(9170) <= (layer2_outputs(7843)) or (layer2_outputs(8846));
    layer3_outputs(9171) <= layer2_outputs(2062);
    layer3_outputs(9172) <= (layer2_outputs(1971)) and (layer2_outputs(10046));
    layer3_outputs(9173) <= (layer2_outputs(7249)) or (layer2_outputs(9554));
    layer3_outputs(9174) <= not(layer2_outputs(9093));
    layer3_outputs(9175) <= layer2_outputs(3698);
    layer3_outputs(9176) <= (layer2_outputs(6674)) and not (layer2_outputs(236));
    layer3_outputs(9177) <= not((layer2_outputs(10166)) and (layer2_outputs(6858)));
    layer3_outputs(9178) <= (layer2_outputs(3658)) and not (layer2_outputs(2893));
    layer3_outputs(9179) <= not((layer2_outputs(3125)) and (layer2_outputs(2200)));
    layer3_outputs(9180) <= layer2_outputs(9052);
    layer3_outputs(9181) <= not(layer2_outputs(8666));
    layer3_outputs(9182) <= not(layer2_outputs(7814));
    layer3_outputs(9183) <= not(layer2_outputs(10025));
    layer3_outputs(9184) <= (layer2_outputs(2001)) or (layer2_outputs(5266));
    layer3_outputs(9185) <= not(layer2_outputs(7234));
    layer3_outputs(9186) <= not(layer2_outputs(2508)) or (layer2_outputs(7245));
    layer3_outputs(9187) <= (layer2_outputs(7413)) and not (layer2_outputs(838));
    layer3_outputs(9188) <= not(layer2_outputs(5301));
    layer3_outputs(9189) <= not(layer2_outputs(4741));
    layer3_outputs(9190) <= not((layer2_outputs(5459)) or (layer2_outputs(5356)));
    layer3_outputs(9191) <= (layer2_outputs(1110)) xor (layer2_outputs(6266));
    layer3_outputs(9192) <= not(layer2_outputs(2103));
    layer3_outputs(9193) <= not((layer2_outputs(2698)) xor (layer2_outputs(8887)));
    layer3_outputs(9194) <= not(layer2_outputs(2876)) or (layer2_outputs(8086));
    layer3_outputs(9195) <= not(layer2_outputs(10091));
    layer3_outputs(9196) <= '1';
    layer3_outputs(9197) <= not(layer2_outputs(4539));
    layer3_outputs(9198) <= layer2_outputs(5873);
    layer3_outputs(9199) <= not(layer2_outputs(3898));
    layer3_outputs(9200) <= not(layer2_outputs(2716));
    layer3_outputs(9201) <= not(layer2_outputs(5858));
    layer3_outputs(9202) <= (layer2_outputs(5447)) and not (layer2_outputs(9922));
    layer3_outputs(9203) <= not(layer2_outputs(9180));
    layer3_outputs(9204) <= '0';
    layer3_outputs(9205) <= (layer2_outputs(3414)) and (layer2_outputs(1112));
    layer3_outputs(9206) <= not((layer2_outputs(3411)) and (layer2_outputs(6861)));
    layer3_outputs(9207) <= not(layer2_outputs(4540)) or (layer2_outputs(7346));
    layer3_outputs(9208) <= not((layer2_outputs(3509)) xor (layer2_outputs(6745)));
    layer3_outputs(9209) <= (layer2_outputs(3525)) and not (layer2_outputs(9057));
    layer3_outputs(9210) <= not(layer2_outputs(9395));
    layer3_outputs(9211) <= layer2_outputs(4629);
    layer3_outputs(9212) <= (layer2_outputs(6650)) xor (layer2_outputs(5546));
    layer3_outputs(9213) <= not(layer2_outputs(9720));
    layer3_outputs(9214) <= not(layer2_outputs(8940));
    layer3_outputs(9215) <= layer2_outputs(2333);
    layer3_outputs(9216) <= not(layer2_outputs(1224));
    layer3_outputs(9217) <= (layer2_outputs(6601)) or (layer2_outputs(5357));
    layer3_outputs(9218) <= (layer2_outputs(1117)) and not (layer2_outputs(3553));
    layer3_outputs(9219) <= (layer2_outputs(6354)) and (layer2_outputs(1067));
    layer3_outputs(9220) <= not(layer2_outputs(9426)) or (layer2_outputs(10210));
    layer3_outputs(9221) <= not(layer2_outputs(7774)) or (layer2_outputs(4076));
    layer3_outputs(9222) <= layer2_outputs(8847);
    layer3_outputs(9223) <= not(layer2_outputs(9824));
    layer3_outputs(9224) <= not(layer2_outputs(8875)) or (layer2_outputs(2815));
    layer3_outputs(9225) <= not(layer2_outputs(5237));
    layer3_outputs(9226) <= (layer2_outputs(2145)) xor (layer2_outputs(933));
    layer3_outputs(9227) <= layer2_outputs(7397);
    layer3_outputs(9228) <= not(layer2_outputs(6872)) or (layer2_outputs(6691));
    layer3_outputs(9229) <= not(layer2_outputs(5737));
    layer3_outputs(9230) <= not(layer2_outputs(2464));
    layer3_outputs(9231) <= (layer2_outputs(1456)) xor (layer2_outputs(3171));
    layer3_outputs(9232) <= layer2_outputs(4876);
    layer3_outputs(9233) <= not((layer2_outputs(99)) and (layer2_outputs(1512)));
    layer3_outputs(9234) <= not(layer2_outputs(6914)) or (layer2_outputs(6784));
    layer3_outputs(9235) <= (layer2_outputs(2929)) and (layer2_outputs(6916));
    layer3_outputs(9236) <= not((layer2_outputs(6308)) xor (layer2_outputs(3379)));
    layer3_outputs(9237) <= not((layer2_outputs(8072)) or (layer2_outputs(1353)));
    layer3_outputs(9238) <= not(layer2_outputs(8552));
    layer3_outputs(9239) <= not((layer2_outputs(2118)) and (layer2_outputs(7830)));
    layer3_outputs(9240) <= layer2_outputs(5586);
    layer3_outputs(9241) <= not((layer2_outputs(4393)) and (layer2_outputs(2212)));
    layer3_outputs(9242) <= layer2_outputs(4405);
    layer3_outputs(9243) <= not((layer2_outputs(7350)) xor (layer2_outputs(4431)));
    layer3_outputs(9244) <= not(layer2_outputs(9874));
    layer3_outputs(9245) <= layer2_outputs(6686);
    layer3_outputs(9246) <= layer2_outputs(978);
    layer3_outputs(9247) <= not(layer2_outputs(426)) or (layer2_outputs(783));
    layer3_outputs(9248) <= not(layer2_outputs(5371));
    layer3_outputs(9249) <= (layer2_outputs(2540)) and not (layer2_outputs(1549));
    layer3_outputs(9250) <= layer2_outputs(212);
    layer3_outputs(9251) <= not(layer2_outputs(8229));
    layer3_outputs(9252) <= not(layer2_outputs(3553));
    layer3_outputs(9253) <= not(layer2_outputs(4484)) or (layer2_outputs(4918));
    layer3_outputs(9254) <= not(layer2_outputs(4950)) or (layer2_outputs(7130));
    layer3_outputs(9255) <= layer2_outputs(2104);
    layer3_outputs(9256) <= (layer2_outputs(7670)) or (layer2_outputs(8512));
    layer3_outputs(9257) <= layer2_outputs(5763);
    layer3_outputs(9258) <= (layer2_outputs(1113)) xor (layer2_outputs(4679));
    layer3_outputs(9259) <= (layer2_outputs(4253)) and not (layer2_outputs(9137));
    layer3_outputs(9260) <= not(layer2_outputs(8358));
    layer3_outputs(9261) <= layer2_outputs(9587);
    layer3_outputs(9262) <= not(layer2_outputs(3111));
    layer3_outputs(9263) <= not(layer2_outputs(3474));
    layer3_outputs(9264) <= not(layer2_outputs(9198));
    layer3_outputs(9265) <= not(layer2_outputs(8522));
    layer3_outputs(9266) <= not(layer2_outputs(5821));
    layer3_outputs(9267) <= not(layer2_outputs(5383));
    layer3_outputs(9268) <= not((layer2_outputs(2311)) and (layer2_outputs(6681)));
    layer3_outputs(9269) <= not(layer2_outputs(7449)) or (layer2_outputs(7234));
    layer3_outputs(9270) <= not(layer2_outputs(858));
    layer3_outputs(9271) <= not(layer2_outputs(7081));
    layer3_outputs(9272) <= not(layer2_outputs(1269));
    layer3_outputs(9273) <= not(layer2_outputs(9231)) or (layer2_outputs(8030));
    layer3_outputs(9274) <= not(layer2_outputs(5020)) or (layer2_outputs(1372));
    layer3_outputs(9275) <= (layer2_outputs(6018)) xor (layer2_outputs(3527));
    layer3_outputs(9276) <= (layer2_outputs(9062)) and (layer2_outputs(5553));
    layer3_outputs(9277) <= layer2_outputs(4487);
    layer3_outputs(9278) <= not(layer2_outputs(2224)) or (layer2_outputs(5290));
    layer3_outputs(9279) <= layer2_outputs(7294);
    layer3_outputs(9280) <= not(layer2_outputs(3491));
    layer3_outputs(9281) <= layer2_outputs(2117);
    layer3_outputs(9282) <= layer2_outputs(1302);
    layer3_outputs(9283) <= (layer2_outputs(1094)) and not (layer2_outputs(9349));
    layer3_outputs(9284) <= not(layer2_outputs(682));
    layer3_outputs(9285) <= not((layer2_outputs(8166)) and (layer2_outputs(6582)));
    layer3_outputs(9286) <= not(layer2_outputs(5795)) or (layer2_outputs(7454));
    layer3_outputs(9287) <= not(layer2_outputs(3325));
    layer3_outputs(9288) <= (layer2_outputs(2069)) and not (layer2_outputs(7251));
    layer3_outputs(9289) <= layer2_outputs(6702);
    layer3_outputs(9290) <= '0';
    layer3_outputs(9291) <= not(layer2_outputs(7312));
    layer3_outputs(9292) <= not(layer2_outputs(5974)) or (layer2_outputs(8700));
    layer3_outputs(9293) <= layer2_outputs(4025);
    layer3_outputs(9294) <= (layer2_outputs(3206)) and not (layer2_outputs(96));
    layer3_outputs(9295) <= not(layer2_outputs(9728));
    layer3_outputs(9296) <= not(layer2_outputs(9260)) or (layer2_outputs(4112));
    layer3_outputs(9297) <= layer2_outputs(127);
    layer3_outputs(9298) <= (layer2_outputs(500)) xor (layer2_outputs(2285));
    layer3_outputs(9299) <= layer2_outputs(1333);
    layer3_outputs(9300) <= not(layer2_outputs(7265)) or (layer2_outputs(1502));
    layer3_outputs(9301) <= layer2_outputs(1718);
    layer3_outputs(9302) <= layer2_outputs(1246);
    layer3_outputs(9303) <= (layer2_outputs(8175)) and not (layer2_outputs(4355));
    layer3_outputs(9304) <= not(layer2_outputs(3148));
    layer3_outputs(9305) <= (layer2_outputs(1619)) and not (layer2_outputs(7127));
    layer3_outputs(9306) <= layer2_outputs(1227);
    layer3_outputs(9307) <= (layer2_outputs(8134)) and not (layer2_outputs(3327));
    layer3_outputs(9308) <= not((layer2_outputs(9310)) and (layer2_outputs(2135)));
    layer3_outputs(9309) <= not(layer2_outputs(6148)) or (layer2_outputs(719));
    layer3_outputs(9310) <= (layer2_outputs(8725)) and (layer2_outputs(3285));
    layer3_outputs(9311) <= layer2_outputs(4775);
    layer3_outputs(9312) <= not(layer2_outputs(1357));
    layer3_outputs(9313) <= layer2_outputs(8029);
    layer3_outputs(9314) <= (layer2_outputs(4835)) and not (layer2_outputs(8137));
    layer3_outputs(9315) <= not(layer2_outputs(356));
    layer3_outputs(9316) <= (layer2_outputs(8133)) and not (layer2_outputs(8001));
    layer3_outputs(9317) <= not(layer2_outputs(8247));
    layer3_outputs(9318) <= (layer2_outputs(1907)) and (layer2_outputs(2573));
    layer3_outputs(9319) <= not(layer2_outputs(10095));
    layer3_outputs(9320) <= not((layer2_outputs(10146)) or (layer2_outputs(5557)));
    layer3_outputs(9321) <= (layer2_outputs(2750)) and not (layer2_outputs(4623));
    layer3_outputs(9322) <= (layer2_outputs(4679)) and (layer2_outputs(4903));
    layer3_outputs(9323) <= '0';
    layer3_outputs(9324) <= layer2_outputs(1550);
    layer3_outputs(9325) <= not(layer2_outputs(4264));
    layer3_outputs(9326) <= (layer2_outputs(4158)) or (layer2_outputs(1352));
    layer3_outputs(9327) <= (layer2_outputs(3829)) or (layer2_outputs(7846));
    layer3_outputs(9328) <= (layer2_outputs(8483)) or (layer2_outputs(10025));
    layer3_outputs(9329) <= layer2_outputs(9687);
    layer3_outputs(9330) <= layer2_outputs(5469);
    layer3_outputs(9331) <= (layer2_outputs(4787)) or (layer2_outputs(3400));
    layer3_outputs(9332) <= layer2_outputs(882);
    layer3_outputs(9333) <= layer2_outputs(8054);
    layer3_outputs(9334) <= not((layer2_outputs(5142)) and (layer2_outputs(2078)));
    layer3_outputs(9335) <= layer2_outputs(5992);
    layer3_outputs(9336) <= layer2_outputs(497);
    layer3_outputs(9337) <= layer2_outputs(9809);
    layer3_outputs(9338) <= layer2_outputs(4845);
    layer3_outputs(9339) <= '1';
    layer3_outputs(9340) <= (layer2_outputs(6721)) or (layer2_outputs(6525));
    layer3_outputs(9341) <= (layer2_outputs(1530)) or (layer2_outputs(4355));
    layer3_outputs(9342) <= layer2_outputs(9003);
    layer3_outputs(9343) <= layer2_outputs(1813);
    layer3_outputs(9344) <= (layer2_outputs(5120)) and (layer2_outputs(3530));
    layer3_outputs(9345) <= '0';
    layer3_outputs(9346) <= layer2_outputs(6979);
    layer3_outputs(9347) <= not(layer2_outputs(9985));
    layer3_outputs(9348) <= layer2_outputs(8713);
    layer3_outputs(9349) <= not(layer2_outputs(2250));
    layer3_outputs(9350) <= (layer2_outputs(9941)) xor (layer2_outputs(6843));
    layer3_outputs(9351) <= layer2_outputs(8914);
    layer3_outputs(9352) <= layer2_outputs(1586);
    layer3_outputs(9353) <= (layer2_outputs(6558)) or (layer2_outputs(9696));
    layer3_outputs(9354) <= not(layer2_outputs(7435));
    layer3_outputs(9355) <= not(layer2_outputs(7798));
    layer3_outputs(9356) <= not(layer2_outputs(3520));
    layer3_outputs(9357) <= not((layer2_outputs(9139)) and (layer2_outputs(6953)));
    layer3_outputs(9358) <= not(layer2_outputs(4371));
    layer3_outputs(9359) <= not((layer2_outputs(5893)) or (layer2_outputs(9988)));
    layer3_outputs(9360) <= (layer2_outputs(5353)) or (layer2_outputs(983));
    layer3_outputs(9361) <= not((layer2_outputs(727)) and (layer2_outputs(4518)));
    layer3_outputs(9362) <= (layer2_outputs(1327)) and (layer2_outputs(7964));
    layer3_outputs(9363) <= not(layer2_outputs(3193));
    layer3_outputs(9364) <= not((layer2_outputs(9909)) and (layer2_outputs(4528)));
    layer3_outputs(9365) <= not(layer2_outputs(360)) or (layer2_outputs(6838));
    layer3_outputs(9366) <= layer2_outputs(9221);
    layer3_outputs(9367) <= not(layer2_outputs(7207));
    layer3_outputs(9368) <= layer2_outputs(3744);
    layer3_outputs(9369) <= (layer2_outputs(4003)) or (layer2_outputs(6345));
    layer3_outputs(9370) <= layer2_outputs(1805);
    layer3_outputs(9371) <= layer2_outputs(275);
    layer3_outputs(9372) <= not(layer2_outputs(5879));
    layer3_outputs(9373) <= (layer2_outputs(9581)) and (layer2_outputs(1789));
    layer3_outputs(9374) <= not(layer2_outputs(8323));
    layer3_outputs(9375) <= layer2_outputs(7155);
    layer3_outputs(9376) <= (layer2_outputs(6837)) and not (layer2_outputs(3830));
    layer3_outputs(9377) <= layer2_outputs(5633);
    layer3_outputs(9378) <= (layer2_outputs(1039)) and (layer2_outputs(5717));
    layer3_outputs(9379) <= (layer2_outputs(464)) xor (layer2_outputs(10064));
    layer3_outputs(9380) <= not(layer2_outputs(5615));
    layer3_outputs(9381) <= not(layer2_outputs(4203));
    layer3_outputs(9382) <= (layer2_outputs(5111)) xor (layer2_outputs(7903));
    layer3_outputs(9383) <= not(layer2_outputs(6179));
    layer3_outputs(9384) <= (layer2_outputs(8543)) and not (layer2_outputs(8666));
    layer3_outputs(9385) <= not((layer2_outputs(6324)) and (layer2_outputs(3864)));
    layer3_outputs(9386) <= not((layer2_outputs(4949)) or (layer2_outputs(3741)));
    layer3_outputs(9387) <= not(layer2_outputs(8490)) or (layer2_outputs(7634));
    layer3_outputs(9388) <= not(layer2_outputs(9420));
    layer3_outputs(9389) <= not(layer2_outputs(6142)) or (layer2_outputs(6032));
    layer3_outputs(9390) <= not(layer2_outputs(8145));
    layer3_outputs(9391) <= not(layer2_outputs(7152)) or (layer2_outputs(2616));
    layer3_outputs(9392) <= layer2_outputs(7412);
    layer3_outputs(9393) <= not((layer2_outputs(318)) xor (layer2_outputs(8731)));
    layer3_outputs(9394) <= (layer2_outputs(8101)) or (layer2_outputs(10173));
    layer3_outputs(9395) <= (layer2_outputs(996)) and (layer2_outputs(7827));
    layer3_outputs(9396) <= layer2_outputs(988);
    layer3_outputs(9397) <= layer2_outputs(6332);
    layer3_outputs(9398) <= layer2_outputs(9834);
    layer3_outputs(9399) <= (layer2_outputs(4621)) xor (layer2_outputs(10231));
    layer3_outputs(9400) <= layer2_outputs(2243);
    layer3_outputs(9401) <= layer2_outputs(8595);
    layer3_outputs(9402) <= layer2_outputs(2367);
    layer3_outputs(9403) <= not(layer2_outputs(4244));
    layer3_outputs(9404) <= not(layer2_outputs(2970)) or (layer2_outputs(5910));
    layer3_outputs(9405) <= layer2_outputs(1272);
    layer3_outputs(9406) <= layer2_outputs(7570);
    layer3_outputs(9407) <= not(layer2_outputs(4242));
    layer3_outputs(9408) <= not((layer2_outputs(2440)) or (layer2_outputs(1248)));
    layer3_outputs(9409) <= layer2_outputs(8236);
    layer3_outputs(9410) <= not(layer2_outputs(1691));
    layer3_outputs(9411) <= layer2_outputs(5190);
    layer3_outputs(9412) <= layer2_outputs(7490);
    layer3_outputs(9413) <= not(layer2_outputs(6258));
    layer3_outputs(9414) <= layer2_outputs(3801);
    layer3_outputs(9415) <= layer2_outputs(1487);
    layer3_outputs(9416) <= (layer2_outputs(7366)) and not (layer2_outputs(8608));
    layer3_outputs(9417) <= '1';
    layer3_outputs(9418) <= not(layer2_outputs(5303));
    layer3_outputs(9419) <= not(layer2_outputs(7637));
    layer3_outputs(9420) <= (layer2_outputs(1070)) and (layer2_outputs(293));
    layer3_outputs(9421) <= not(layer2_outputs(7465)) or (layer2_outputs(9734));
    layer3_outputs(9422) <= layer2_outputs(1803);
    layer3_outputs(9423) <= layer2_outputs(8401);
    layer3_outputs(9424) <= not(layer2_outputs(7278)) or (layer2_outputs(6860));
    layer3_outputs(9425) <= not((layer2_outputs(1153)) and (layer2_outputs(4223)));
    layer3_outputs(9426) <= (layer2_outputs(63)) and not (layer2_outputs(6287));
    layer3_outputs(9427) <= (layer2_outputs(2428)) and not (layer2_outputs(1548));
    layer3_outputs(9428) <= (layer2_outputs(4860)) and not (layer2_outputs(884));
    layer3_outputs(9429) <= (layer2_outputs(7273)) and not (layer2_outputs(1622));
    layer3_outputs(9430) <= not(layer2_outputs(9019)) or (layer2_outputs(10039));
    layer3_outputs(9431) <= layer2_outputs(3126);
    layer3_outputs(9432) <= not(layer2_outputs(1578));
    layer3_outputs(9433) <= layer2_outputs(7747);
    layer3_outputs(9434) <= not(layer2_outputs(5305)) or (layer2_outputs(7608));
    layer3_outputs(9435) <= (layer2_outputs(8455)) xor (layer2_outputs(4544));
    layer3_outputs(9436) <= not((layer2_outputs(2828)) xor (layer2_outputs(8511)));
    layer3_outputs(9437) <= (layer2_outputs(8202)) and not (layer2_outputs(8142));
    layer3_outputs(9438) <= '1';
    layer3_outputs(9439) <= not(layer2_outputs(5833));
    layer3_outputs(9440) <= not((layer2_outputs(6049)) xor (layer2_outputs(3420)));
    layer3_outputs(9441) <= not((layer2_outputs(9998)) and (layer2_outputs(7525)));
    layer3_outputs(9442) <= not((layer2_outputs(1047)) and (layer2_outputs(3068)));
    layer3_outputs(9443) <= not(layer2_outputs(5978));
    layer3_outputs(9444) <= not(layer2_outputs(5746));
    layer3_outputs(9445) <= (layer2_outputs(6717)) and (layer2_outputs(8124));
    layer3_outputs(9446) <= layer2_outputs(7071);
    layer3_outputs(9447) <= layer2_outputs(2623);
    layer3_outputs(9448) <= not(layer2_outputs(8281));
    layer3_outputs(9449) <= (layer2_outputs(6387)) xor (layer2_outputs(7384));
    layer3_outputs(9450) <= layer2_outputs(3660);
    layer3_outputs(9451) <= not(layer2_outputs(9645));
    layer3_outputs(9452) <= not((layer2_outputs(1348)) or (layer2_outputs(528)));
    layer3_outputs(9453) <= not(layer2_outputs(6931)) or (layer2_outputs(6007));
    layer3_outputs(9454) <= (layer2_outputs(2909)) and not (layer2_outputs(6250));
    layer3_outputs(9455) <= layer2_outputs(3253);
    layer3_outputs(9456) <= (layer2_outputs(7693)) and not (layer2_outputs(4937));
    layer3_outputs(9457) <= (layer2_outputs(2189)) and not (layer2_outputs(460));
    layer3_outputs(9458) <= (layer2_outputs(2755)) and not (layer2_outputs(1284));
    layer3_outputs(9459) <= (layer2_outputs(6998)) and not (layer2_outputs(8889));
    layer3_outputs(9460) <= (layer2_outputs(4243)) and not (layer2_outputs(4782));
    layer3_outputs(9461) <= (layer2_outputs(2270)) and (layer2_outputs(460));
    layer3_outputs(9462) <= not(layer2_outputs(8744)) or (layer2_outputs(3159));
    layer3_outputs(9463) <= not(layer2_outputs(9329));
    layer3_outputs(9464) <= not(layer2_outputs(3811));
    layer3_outputs(9465) <= layer2_outputs(4758);
    layer3_outputs(9466) <= not(layer2_outputs(604)) or (layer2_outputs(628));
    layer3_outputs(9467) <= not(layer2_outputs(7360));
    layer3_outputs(9468) <= (layer2_outputs(3062)) xor (layer2_outputs(59));
    layer3_outputs(9469) <= layer2_outputs(6052);
    layer3_outputs(9470) <= not((layer2_outputs(4379)) and (layer2_outputs(7023)));
    layer3_outputs(9471) <= layer2_outputs(9194);
    layer3_outputs(9472) <= not(layer2_outputs(2063));
    layer3_outputs(9473) <= (layer2_outputs(352)) and not (layer2_outputs(9815));
    layer3_outputs(9474) <= not(layer2_outputs(8244));
    layer3_outputs(9475) <= layer2_outputs(1771);
    layer3_outputs(9476) <= not(layer2_outputs(7955));
    layer3_outputs(9477) <= layer2_outputs(26);
    layer3_outputs(9478) <= not((layer2_outputs(642)) xor (layer2_outputs(773)));
    layer3_outputs(9479) <= layer2_outputs(7902);
    layer3_outputs(9480) <= '1';
    layer3_outputs(9481) <= not(layer2_outputs(5887));
    layer3_outputs(9482) <= not((layer2_outputs(7809)) xor (layer2_outputs(9442)));
    layer3_outputs(9483) <= not((layer2_outputs(6530)) or (layer2_outputs(4179)));
    layer3_outputs(9484) <= not(layer2_outputs(5287)) or (layer2_outputs(2431));
    layer3_outputs(9485) <= not(layer2_outputs(3355));
    layer3_outputs(9486) <= not(layer2_outputs(7508));
    layer3_outputs(9487) <= not(layer2_outputs(493));
    layer3_outputs(9488) <= not(layer2_outputs(5583));
    layer3_outputs(9489) <= not(layer2_outputs(4010));
    layer3_outputs(9490) <= not(layer2_outputs(2581));
    layer3_outputs(9491) <= layer2_outputs(9655);
    layer3_outputs(9492) <= not((layer2_outputs(2223)) or (layer2_outputs(5671)));
    layer3_outputs(9493) <= not(layer2_outputs(7197));
    layer3_outputs(9494) <= not((layer2_outputs(2954)) or (layer2_outputs(7324)));
    layer3_outputs(9495) <= not(layer2_outputs(9914));
    layer3_outputs(9496) <= layer2_outputs(1599);
    layer3_outputs(9497) <= not((layer2_outputs(9704)) xor (layer2_outputs(2479)));
    layer3_outputs(9498) <= (layer2_outputs(2140)) xor (layer2_outputs(5570));
    layer3_outputs(9499) <= layer2_outputs(8771);
    layer3_outputs(9500) <= not(layer2_outputs(7513)) or (layer2_outputs(2050));
    layer3_outputs(9501) <= layer2_outputs(7847);
    layer3_outputs(9502) <= not(layer2_outputs(4814));
    layer3_outputs(9503) <= not(layer2_outputs(6730));
    layer3_outputs(9504) <= (layer2_outputs(2754)) and (layer2_outputs(8423));
    layer3_outputs(9505) <= '0';
    layer3_outputs(9506) <= not(layer2_outputs(8037)) or (layer2_outputs(7858));
    layer3_outputs(9507) <= layer2_outputs(1642);
    layer3_outputs(9508) <= (layer2_outputs(7445)) xor (layer2_outputs(1919));
    layer3_outputs(9509) <= not(layer2_outputs(7375));
    layer3_outputs(9510) <= (layer2_outputs(3795)) and not (layer2_outputs(3347));
    layer3_outputs(9511) <= not(layer2_outputs(6405));
    layer3_outputs(9512) <= not(layer2_outputs(2011)) or (layer2_outputs(3128));
    layer3_outputs(9513) <= not(layer2_outputs(5932)) or (layer2_outputs(3527));
    layer3_outputs(9514) <= not((layer2_outputs(3785)) or (layer2_outputs(7455)));
    layer3_outputs(9515) <= (layer2_outputs(8788)) xor (layer2_outputs(7183));
    layer3_outputs(9516) <= (layer2_outputs(8747)) and (layer2_outputs(5036));
    layer3_outputs(9517) <= (layer2_outputs(980)) and not (layer2_outputs(7670));
    layer3_outputs(9518) <= layer2_outputs(5472);
    layer3_outputs(9519) <= not((layer2_outputs(9321)) or (layer2_outputs(3667)));
    layer3_outputs(9520) <= (layer2_outputs(3606)) and not (layer2_outputs(4480));
    layer3_outputs(9521) <= (layer2_outputs(2514)) and not (layer2_outputs(4864));
    layer3_outputs(9522) <= not(layer2_outputs(5275));
    layer3_outputs(9523) <= layer2_outputs(4375);
    layer3_outputs(9524) <= not(layer2_outputs(8170));
    layer3_outputs(9525) <= not(layer2_outputs(2100));
    layer3_outputs(9526) <= (layer2_outputs(8937)) and not (layer2_outputs(8536));
    layer3_outputs(9527) <= not(layer2_outputs(2157)) or (layer2_outputs(6502));
    layer3_outputs(9528) <= not((layer2_outputs(1830)) and (layer2_outputs(9652)));
    layer3_outputs(9529) <= (layer2_outputs(3663)) and (layer2_outputs(5925));
    layer3_outputs(9530) <= (layer2_outputs(1097)) and (layer2_outputs(4737));
    layer3_outputs(9531) <= (layer2_outputs(10133)) and (layer2_outputs(10069));
    layer3_outputs(9532) <= not((layer2_outputs(6199)) or (layer2_outputs(9812)));
    layer3_outputs(9533) <= not(layer2_outputs(3605));
    layer3_outputs(9534) <= layer2_outputs(2974);
    layer3_outputs(9535) <= layer2_outputs(8638);
    layer3_outputs(9536) <= not((layer2_outputs(4220)) and (layer2_outputs(5261)));
    layer3_outputs(9537) <= not(layer2_outputs(829));
    layer3_outputs(9538) <= (layer2_outputs(6233)) xor (layer2_outputs(5928));
    layer3_outputs(9539) <= '1';
    layer3_outputs(9540) <= '1';
    layer3_outputs(9541) <= not(layer2_outputs(7960));
    layer3_outputs(9542) <= not(layer2_outputs(9769));
    layer3_outputs(9543) <= not(layer2_outputs(3216)) or (layer2_outputs(8591));
    layer3_outputs(9544) <= (layer2_outputs(8998)) and not (layer2_outputs(6104));
    layer3_outputs(9545) <= (layer2_outputs(1006)) xor (layer2_outputs(753));
    layer3_outputs(9546) <= not((layer2_outputs(1474)) and (layer2_outputs(2996)));
    layer3_outputs(9547) <= not(layer2_outputs(2380));
    layer3_outputs(9548) <= (layer2_outputs(8556)) or (layer2_outputs(6193));
    layer3_outputs(9549) <= not(layer2_outputs(1202));
    layer3_outputs(9550) <= not(layer2_outputs(6037));
    layer3_outputs(9551) <= (layer2_outputs(3347)) and not (layer2_outputs(6900));
    layer3_outputs(9552) <= not(layer2_outputs(4180));
    layer3_outputs(9553) <= (layer2_outputs(9723)) or (layer2_outputs(1402));
    layer3_outputs(9554) <= layer2_outputs(7507);
    layer3_outputs(9555) <= layer2_outputs(773);
    layer3_outputs(9556) <= not((layer2_outputs(7378)) or (layer2_outputs(7312)));
    layer3_outputs(9557) <= not(layer2_outputs(1441));
    layer3_outputs(9558) <= not(layer2_outputs(2246));
    layer3_outputs(9559) <= layer2_outputs(8287);
    layer3_outputs(9560) <= not(layer2_outputs(7530));
    layer3_outputs(9561) <= layer2_outputs(1487);
    layer3_outputs(9562) <= '0';
    layer3_outputs(9563) <= (layer2_outputs(4685)) or (layer2_outputs(6591));
    layer3_outputs(9564) <= layer2_outputs(1864);
    layer3_outputs(9565) <= not(layer2_outputs(5550));
    layer3_outputs(9566) <= not(layer2_outputs(9544));
    layer3_outputs(9567) <= not(layer2_outputs(6630));
    layer3_outputs(9568) <= layer2_outputs(4243);
    layer3_outputs(9569) <= not(layer2_outputs(1268)) or (layer2_outputs(3168));
    layer3_outputs(9570) <= (layer2_outputs(2906)) and (layer2_outputs(7079));
    layer3_outputs(9571) <= layer2_outputs(5139);
    layer3_outputs(9572) <= not((layer2_outputs(2926)) xor (layer2_outputs(91)));
    layer3_outputs(9573) <= layer2_outputs(1808);
    layer3_outputs(9574) <= layer2_outputs(4560);
    layer3_outputs(9575) <= not(layer2_outputs(2597));
    layer3_outputs(9576) <= layer2_outputs(2666);
    layer3_outputs(9577) <= layer2_outputs(5536);
    layer3_outputs(9578) <= not(layer2_outputs(6430));
    layer3_outputs(9579) <= not(layer2_outputs(8633));
    layer3_outputs(9580) <= layer2_outputs(4504);
    layer3_outputs(9581) <= not(layer2_outputs(3699));
    layer3_outputs(9582) <= layer2_outputs(4304);
    layer3_outputs(9583) <= not(layer2_outputs(4022));
    layer3_outputs(9584) <= not(layer2_outputs(10168));
    layer3_outputs(9585) <= not(layer2_outputs(4011));
    layer3_outputs(9586) <= not(layer2_outputs(6083));
    layer3_outputs(9587) <= not(layer2_outputs(6817));
    layer3_outputs(9588) <= not(layer2_outputs(8587));
    layer3_outputs(9589) <= layer2_outputs(123);
    layer3_outputs(9590) <= (layer2_outputs(6049)) and not (layer2_outputs(7037));
    layer3_outputs(9591) <= layer2_outputs(2178);
    layer3_outputs(9592) <= not(layer2_outputs(2513));
    layer3_outputs(9593) <= not((layer2_outputs(6471)) and (layer2_outputs(9132)));
    layer3_outputs(9594) <= not(layer2_outputs(3729));
    layer3_outputs(9595) <= layer2_outputs(3201);
    layer3_outputs(9596) <= layer2_outputs(7274);
    layer3_outputs(9597) <= not(layer2_outputs(3632));
    layer3_outputs(9598) <= not(layer2_outputs(8210));
    layer3_outputs(9599) <= not(layer2_outputs(5779));
    layer3_outputs(9600) <= not(layer2_outputs(4565));
    layer3_outputs(9601) <= not(layer2_outputs(3122));
    layer3_outputs(9602) <= layer2_outputs(5437);
    layer3_outputs(9603) <= (layer2_outputs(1313)) xor (layer2_outputs(7260));
    layer3_outputs(9604) <= not(layer2_outputs(610));
    layer3_outputs(9605) <= layer2_outputs(2327);
    layer3_outputs(9606) <= not(layer2_outputs(3407));
    layer3_outputs(9607) <= (layer2_outputs(9103)) xor (layer2_outputs(9844));
    layer3_outputs(9608) <= not(layer2_outputs(2229));
    layer3_outputs(9609) <= not(layer2_outputs(6063));
    layer3_outputs(9610) <= layer2_outputs(7269);
    layer3_outputs(9611) <= not(layer2_outputs(9508)) or (layer2_outputs(10114));
    layer3_outputs(9612) <= not(layer2_outputs(1254)) or (layer2_outputs(1385));
    layer3_outputs(9613) <= layer2_outputs(6943);
    layer3_outputs(9614) <= not(layer2_outputs(1184));
    layer3_outputs(9615) <= not((layer2_outputs(6765)) xor (layer2_outputs(8885)));
    layer3_outputs(9616) <= layer2_outputs(7035);
    layer3_outputs(9617) <= not(layer2_outputs(7370));
    layer3_outputs(9618) <= not(layer2_outputs(4498));
    layer3_outputs(9619) <= layer2_outputs(1227);
    layer3_outputs(9620) <= not((layer2_outputs(8220)) xor (layer2_outputs(10182)));
    layer3_outputs(9621) <= layer2_outputs(7772);
    layer3_outputs(9622) <= (layer2_outputs(45)) and not (layer2_outputs(10181));
    layer3_outputs(9623) <= not(layer2_outputs(1965)) or (layer2_outputs(8408));
    layer3_outputs(9624) <= layer2_outputs(9869);
    layer3_outputs(9625) <= not(layer2_outputs(9188)) or (layer2_outputs(8026));
    layer3_outputs(9626) <= (layer2_outputs(4648)) xor (layer2_outputs(3969));
    layer3_outputs(9627) <= (layer2_outputs(7582)) and not (layer2_outputs(332));
    layer3_outputs(9628) <= '1';
    layer3_outputs(9629) <= (layer2_outputs(6142)) xor (layer2_outputs(9113));
    layer3_outputs(9630) <= (layer2_outputs(5702)) and not (layer2_outputs(10075));
    layer3_outputs(9631) <= layer2_outputs(6003);
    layer3_outputs(9632) <= not((layer2_outputs(3900)) and (layer2_outputs(6903)));
    layer3_outputs(9633) <= not(layer2_outputs(7894));
    layer3_outputs(9634) <= not(layer2_outputs(1564));
    layer3_outputs(9635) <= layer2_outputs(9091);
    layer3_outputs(9636) <= '1';
    layer3_outputs(9637) <= not((layer2_outputs(2147)) and (layer2_outputs(3958)));
    layer3_outputs(9638) <= not(layer2_outputs(106)) or (layer2_outputs(1475));
    layer3_outputs(9639) <= layer2_outputs(1528);
    layer3_outputs(9640) <= not(layer2_outputs(6451)) or (layer2_outputs(2232));
    layer3_outputs(9641) <= (layer2_outputs(2495)) or (layer2_outputs(7241));
    layer3_outputs(9642) <= not(layer2_outputs(7533));
    layer3_outputs(9643) <= (layer2_outputs(1105)) and not (layer2_outputs(4972));
    layer3_outputs(9644) <= (layer2_outputs(2784)) xor (layer2_outputs(4490));
    layer3_outputs(9645) <= not(layer2_outputs(6927)) or (layer2_outputs(6146));
    layer3_outputs(9646) <= not(layer2_outputs(5603)) or (layer2_outputs(1010));
    layer3_outputs(9647) <= (layer2_outputs(1243)) xor (layer2_outputs(4824));
    layer3_outputs(9648) <= not(layer2_outputs(641));
    layer3_outputs(9649) <= (layer2_outputs(6678)) or (layer2_outputs(10062));
    layer3_outputs(9650) <= '0';
    layer3_outputs(9651) <= layer2_outputs(4120);
    layer3_outputs(9652) <= not(layer2_outputs(5510));
    layer3_outputs(9653) <= layer2_outputs(9714);
    layer3_outputs(9654) <= not(layer2_outputs(9282));
    layer3_outputs(9655) <= not((layer2_outputs(3186)) or (layer2_outputs(5560)));
    layer3_outputs(9656) <= not(layer2_outputs(1636)) or (layer2_outputs(5434));
    layer3_outputs(9657) <= (layer2_outputs(10190)) and not (layer2_outputs(9445));
    layer3_outputs(9658) <= not(layer2_outputs(2952));
    layer3_outputs(9659) <= layer2_outputs(2532);
    layer3_outputs(9660) <= not((layer2_outputs(2226)) xor (layer2_outputs(6103)));
    layer3_outputs(9661) <= not(layer2_outputs(2133)) or (layer2_outputs(7658));
    layer3_outputs(9662) <= not(layer2_outputs(2937));
    layer3_outputs(9663) <= layer2_outputs(1586);
    layer3_outputs(9664) <= layer2_outputs(4123);
    layer3_outputs(9665) <= layer2_outputs(3445);
    layer3_outputs(9666) <= layer2_outputs(3055);
    layer3_outputs(9667) <= not(layer2_outputs(3793));
    layer3_outputs(9668) <= not(layer2_outputs(7893)) or (layer2_outputs(2767));
    layer3_outputs(9669) <= (layer2_outputs(8883)) and not (layer2_outputs(551));
    layer3_outputs(9670) <= (layer2_outputs(3857)) and not (layer2_outputs(6855));
    layer3_outputs(9671) <= '1';
    layer3_outputs(9672) <= (layer2_outputs(2563)) and (layer2_outputs(5583));
    layer3_outputs(9673) <= (layer2_outputs(8350)) or (layer2_outputs(5599));
    layer3_outputs(9674) <= (layer2_outputs(9024)) or (layer2_outputs(927));
    layer3_outputs(9675) <= '0';
    layer3_outputs(9676) <= layer2_outputs(8590);
    layer3_outputs(9677) <= layer2_outputs(6884);
    layer3_outputs(9678) <= not((layer2_outputs(9507)) and (layer2_outputs(8332)));
    layer3_outputs(9679) <= not((layer2_outputs(4598)) xor (layer2_outputs(5006)));
    layer3_outputs(9680) <= not((layer2_outputs(3702)) and (layer2_outputs(2921)));
    layer3_outputs(9681) <= not(layer2_outputs(9301));
    layer3_outputs(9682) <= layer2_outputs(7690);
    layer3_outputs(9683) <= not(layer2_outputs(1849));
    layer3_outputs(9684) <= not(layer2_outputs(3262));
    layer3_outputs(9685) <= (layer2_outputs(2868)) and not (layer2_outputs(8466));
    layer3_outputs(9686) <= (layer2_outputs(6747)) and not (layer2_outputs(1804));
    layer3_outputs(9687) <= (layer2_outputs(1393)) and not (layer2_outputs(2164));
    layer3_outputs(9688) <= not((layer2_outputs(8193)) and (layer2_outputs(3465)));
    layer3_outputs(9689) <= (layer2_outputs(6243)) and not (layer2_outputs(7411));
    layer3_outputs(9690) <= (layer2_outputs(2448)) and (layer2_outputs(1674));
    layer3_outputs(9691) <= (layer2_outputs(4100)) and (layer2_outputs(8139));
    layer3_outputs(9692) <= not(layer2_outputs(10201)) or (layer2_outputs(9209));
    layer3_outputs(9693) <= layer2_outputs(9980);
    layer3_outputs(9694) <= not(layer2_outputs(5826));
    layer3_outputs(9695) <= layer2_outputs(7849);
    layer3_outputs(9696) <= (layer2_outputs(6732)) and not (layer2_outputs(9107));
    layer3_outputs(9697) <= not(layer2_outputs(4564)) or (layer2_outputs(4712));
    layer3_outputs(9698) <= not(layer2_outputs(7188));
    layer3_outputs(9699) <= not(layer2_outputs(7070));
    layer3_outputs(9700) <= not(layer2_outputs(7344));
    layer3_outputs(9701) <= '1';
    layer3_outputs(9702) <= '1';
    layer3_outputs(9703) <= not(layer2_outputs(9343));
    layer3_outputs(9704) <= not((layer2_outputs(7126)) xor (layer2_outputs(9987)));
    layer3_outputs(9705) <= not(layer2_outputs(3415));
    layer3_outputs(9706) <= layer2_outputs(1881);
    layer3_outputs(9707) <= layer2_outputs(3507);
    layer3_outputs(9708) <= not(layer2_outputs(4226));
    layer3_outputs(9709) <= (layer2_outputs(4001)) or (layer2_outputs(8248));
    layer3_outputs(9710) <= not(layer2_outputs(675));
    layer3_outputs(9711) <= '1';
    layer3_outputs(9712) <= not(layer2_outputs(3662));
    layer3_outputs(9713) <= (layer2_outputs(8486)) and not (layer2_outputs(384));
    layer3_outputs(9714) <= (layer2_outputs(9251)) and (layer2_outputs(3789));
    layer3_outputs(9715) <= layer2_outputs(4495);
    layer3_outputs(9716) <= not((layer2_outputs(3141)) xor (layer2_outputs(8475)));
    layer3_outputs(9717) <= not(layer2_outputs(1529));
    layer3_outputs(9718) <= layer2_outputs(8566);
    layer3_outputs(9719) <= layer2_outputs(5764);
    layer3_outputs(9720) <= not(layer2_outputs(10158));
    layer3_outputs(9721) <= layer2_outputs(3960);
    layer3_outputs(9722) <= not(layer2_outputs(5762)) or (layer2_outputs(2579));
    layer3_outputs(9723) <= layer2_outputs(3953);
    layer3_outputs(9724) <= not(layer2_outputs(2604)) or (layer2_outputs(4966));
    layer3_outputs(9725) <= not(layer2_outputs(4047));
    layer3_outputs(9726) <= not(layer2_outputs(898)) or (layer2_outputs(8524));
    layer3_outputs(9727) <= not((layer2_outputs(8389)) and (layer2_outputs(592)));
    layer3_outputs(9728) <= layer2_outputs(5471);
    layer3_outputs(9729) <= not((layer2_outputs(10157)) or (layer2_outputs(5397)));
    layer3_outputs(9730) <= layer2_outputs(9308);
    layer3_outputs(9731) <= (layer2_outputs(4459)) or (layer2_outputs(6623));
    layer3_outputs(9732) <= (layer2_outputs(9277)) and (layer2_outputs(2650));
    layer3_outputs(9733) <= not(layer2_outputs(1918)) or (layer2_outputs(510));
    layer3_outputs(9734) <= not(layer2_outputs(9197));
    layer3_outputs(9735) <= layer2_outputs(3769);
    layer3_outputs(9736) <= not(layer2_outputs(4331));
    layer3_outputs(9737) <= not((layer2_outputs(158)) and (layer2_outputs(3503)));
    layer3_outputs(9738) <= not((layer2_outputs(3940)) or (layer2_outputs(9044)));
    layer3_outputs(9739) <= layer2_outputs(4198);
    layer3_outputs(9740) <= not(layer2_outputs(7051));
    layer3_outputs(9741) <= (layer2_outputs(3252)) and (layer2_outputs(4853));
    layer3_outputs(9742) <= layer2_outputs(5840);
    layer3_outputs(9743) <= layer2_outputs(7860);
    layer3_outputs(9744) <= not(layer2_outputs(7863));
    layer3_outputs(9745) <= not(layer2_outputs(5517));
    layer3_outputs(9746) <= (layer2_outputs(2788)) and not (layer2_outputs(2897));
    layer3_outputs(9747) <= layer2_outputs(6719);
    layer3_outputs(9748) <= not(layer2_outputs(2985));
    layer3_outputs(9749) <= not(layer2_outputs(2040));
    layer3_outputs(9750) <= layer2_outputs(1206);
    layer3_outputs(9751) <= not((layer2_outputs(3762)) and (layer2_outputs(34)));
    layer3_outputs(9752) <= '1';
    layer3_outputs(9753) <= (layer2_outputs(6601)) or (layer2_outputs(10121));
    layer3_outputs(9754) <= not(layer2_outputs(6949));
    layer3_outputs(9755) <= (layer2_outputs(8799)) or (layer2_outputs(8668));
    layer3_outputs(9756) <= not((layer2_outputs(5122)) or (layer2_outputs(8420)));
    layer3_outputs(9757) <= not((layer2_outputs(5792)) or (layer2_outputs(8925)));
    layer3_outputs(9758) <= (layer2_outputs(379)) xor (layer2_outputs(4120));
    layer3_outputs(9759) <= layer2_outputs(479);
    layer3_outputs(9760) <= not(layer2_outputs(7265));
    layer3_outputs(9761) <= layer2_outputs(5752);
    layer3_outputs(9762) <= layer2_outputs(10166);
    layer3_outputs(9763) <= layer2_outputs(6192);
    layer3_outputs(9764) <= layer2_outputs(4324);
    layer3_outputs(9765) <= (layer2_outputs(6696)) or (layer2_outputs(4549));
    layer3_outputs(9766) <= not(layer2_outputs(3058));
    layer3_outputs(9767) <= not(layer2_outputs(8823));
    layer3_outputs(9768) <= (layer2_outputs(9889)) and not (layer2_outputs(4256));
    layer3_outputs(9769) <= not((layer2_outputs(8027)) xor (layer2_outputs(679)));
    layer3_outputs(9770) <= not(layer2_outputs(6510)) or (layer2_outputs(7780));
    layer3_outputs(9771) <= not(layer2_outputs(3354));
    layer3_outputs(9772) <= not((layer2_outputs(5899)) xor (layer2_outputs(2865)));
    layer3_outputs(9773) <= (layer2_outputs(1491)) and (layer2_outputs(3294));
    layer3_outputs(9774) <= layer2_outputs(532);
    layer3_outputs(9775) <= layer2_outputs(6786);
    layer3_outputs(9776) <= layer2_outputs(571);
    layer3_outputs(9777) <= (layer2_outputs(3659)) xor (layer2_outputs(1772));
    layer3_outputs(9778) <= '0';
    layer3_outputs(9779) <= not(layer2_outputs(3804)) or (layer2_outputs(1455));
    layer3_outputs(9780) <= layer2_outputs(4230);
    layer3_outputs(9781) <= (layer2_outputs(8055)) and not (layer2_outputs(8041));
    layer3_outputs(9782) <= not(layer2_outputs(9095));
    layer3_outputs(9783) <= not((layer2_outputs(8045)) or (layer2_outputs(3267)));
    layer3_outputs(9784) <= layer2_outputs(1609);
    layer3_outputs(9785) <= layer2_outputs(2368);
    layer3_outputs(9786) <= '1';
    layer3_outputs(9787) <= layer2_outputs(4550);
    layer3_outputs(9788) <= not(layer2_outputs(1476));
    layer3_outputs(9789) <= not(layer2_outputs(3548));
    layer3_outputs(9790) <= (layer2_outputs(9968)) or (layer2_outputs(82));
    layer3_outputs(9791) <= not((layer2_outputs(8855)) and (layer2_outputs(2021)));
    layer3_outputs(9792) <= '0';
    layer3_outputs(9793) <= (layer2_outputs(1758)) xor (layer2_outputs(5632));
    layer3_outputs(9794) <= (layer2_outputs(5580)) and (layer2_outputs(2622));
    layer3_outputs(9795) <= not(layer2_outputs(9358));
    layer3_outputs(9796) <= not(layer2_outputs(5969)) or (layer2_outputs(3693));
    layer3_outputs(9797) <= not((layer2_outputs(3562)) xor (layer2_outputs(4659)));
    layer3_outputs(9798) <= (layer2_outputs(6164)) and not (layer2_outputs(4581));
    layer3_outputs(9799) <= '1';
    layer3_outputs(9800) <= (layer2_outputs(2172)) and (layer2_outputs(6147));
    layer3_outputs(9801) <= (layer2_outputs(2416)) xor (layer2_outputs(1291));
    layer3_outputs(9802) <= not((layer2_outputs(7978)) or (layer2_outputs(7580)));
    layer3_outputs(9803) <= (layer2_outputs(5475)) and not (layer2_outputs(940));
    layer3_outputs(9804) <= layer2_outputs(3991);
    layer3_outputs(9805) <= layer2_outputs(7200);
    layer3_outputs(9806) <= not((layer2_outputs(4461)) or (layer2_outputs(9886)));
    layer3_outputs(9807) <= not(layer2_outputs(1214));
    layer3_outputs(9808) <= (layer2_outputs(6615)) and not (layer2_outputs(4144));
    layer3_outputs(9809) <= not(layer2_outputs(8067));
    layer3_outputs(9810) <= not((layer2_outputs(3790)) and (layer2_outputs(5866)));
    layer3_outputs(9811) <= '0';
    layer3_outputs(9812) <= (layer2_outputs(612)) and not (layer2_outputs(3953));
    layer3_outputs(9813) <= not(layer2_outputs(4858));
    layer3_outputs(9814) <= (layer2_outputs(1171)) xor (layer2_outputs(5904));
    layer3_outputs(9815) <= layer2_outputs(8963);
    layer3_outputs(9816) <= layer2_outputs(8348);
    layer3_outputs(9817) <= layer2_outputs(2230);
    layer3_outputs(9818) <= not((layer2_outputs(9434)) or (layer2_outputs(1220)));
    layer3_outputs(9819) <= layer2_outputs(9289);
    layer3_outputs(9820) <= not((layer2_outputs(4398)) or (layer2_outputs(1258)));
    layer3_outputs(9821) <= layer2_outputs(1469);
    layer3_outputs(9822) <= (layer2_outputs(7665)) or (layer2_outputs(9332));
    layer3_outputs(9823) <= (layer2_outputs(2998)) or (layer2_outputs(7395));
    layer3_outputs(9824) <= '1';
    layer3_outputs(9825) <= layer2_outputs(508);
    layer3_outputs(9826) <= layer2_outputs(7782);
    layer3_outputs(9827) <= layer2_outputs(2076);
    layer3_outputs(9828) <= not(layer2_outputs(8940));
    layer3_outputs(9829) <= layer2_outputs(9903);
    layer3_outputs(9830) <= layer2_outputs(5549);
    layer3_outputs(9831) <= (layer2_outputs(2873)) xor (layer2_outputs(3268));
    layer3_outputs(9832) <= not(layer2_outputs(9402));
    layer3_outputs(9833) <= not(layer2_outputs(307));
    layer3_outputs(9834) <= layer2_outputs(8047);
    layer3_outputs(9835) <= not(layer2_outputs(7411)) or (layer2_outputs(1411));
    layer3_outputs(9836) <= not((layer2_outputs(5379)) and (layer2_outputs(1604)));
    layer3_outputs(9837) <= not((layer2_outputs(6325)) and (layer2_outputs(8198)));
    layer3_outputs(9838) <= not((layer2_outputs(503)) xor (layer2_outputs(7331)));
    layer3_outputs(9839) <= layer2_outputs(9126);
    layer3_outputs(9840) <= not(layer2_outputs(5001)) or (layer2_outputs(875));
    layer3_outputs(9841) <= not(layer2_outputs(6303));
    layer3_outputs(9842) <= not(layer2_outputs(7984));
    layer3_outputs(9843) <= not(layer2_outputs(4299));
    layer3_outputs(9844) <= (layer2_outputs(9011)) or (layer2_outputs(4236));
    layer3_outputs(9845) <= layer2_outputs(9024);
    layer3_outputs(9846) <= (layer2_outputs(3999)) or (layer2_outputs(1225));
    layer3_outputs(9847) <= not((layer2_outputs(2971)) and (layer2_outputs(10079)));
    layer3_outputs(9848) <= (layer2_outputs(3988)) and (layer2_outputs(5689));
    layer3_outputs(9849) <= layer2_outputs(9951);
    layer3_outputs(9850) <= not(layer2_outputs(676));
    layer3_outputs(9851) <= not(layer2_outputs(5633));
    layer3_outputs(9852) <= not(layer2_outputs(543));
    layer3_outputs(9853) <= layer2_outputs(3284);
    layer3_outputs(9854) <= not(layer2_outputs(4792)) or (layer2_outputs(5351));
    layer3_outputs(9855) <= layer2_outputs(2772);
    layer3_outputs(9856) <= '0';
    layer3_outputs(9857) <= not(layer2_outputs(8942)) or (layer2_outputs(3770));
    layer3_outputs(9858) <= not(layer2_outputs(3683));
    layer3_outputs(9859) <= (layer2_outputs(1554)) and not (layer2_outputs(4655));
    layer3_outputs(9860) <= layer2_outputs(7223);
    layer3_outputs(9861) <= (layer2_outputs(8916)) and (layer2_outputs(6483));
    layer3_outputs(9862) <= layer2_outputs(8077);
    layer3_outputs(9863) <= layer2_outputs(1791);
    layer3_outputs(9864) <= not(layer2_outputs(1481));
    layer3_outputs(9865) <= '1';
    layer3_outputs(9866) <= layer2_outputs(10122);
    layer3_outputs(9867) <= not(layer2_outputs(6153)) or (layer2_outputs(7770));
    layer3_outputs(9868) <= (layer2_outputs(7181)) xor (layer2_outputs(2225));
    layer3_outputs(9869) <= not(layer2_outputs(2724));
    layer3_outputs(9870) <= not(layer2_outputs(4191));
    layer3_outputs(9871) <= not(layer2_outputs(682));
    layer3_outputs(9872) <= not(layer2_outputs(8207));
    layer3_outputs(9873) <= not(layer2_outputs(10133)) or (layer2_outputs(4223));
    layer3_outputs(9874) <= layer2_outputs(8158);
    layer3_outputs(9875) <= not(layer2_outputs(892));
    layer3_outputs(9876) <= not((layer2_outputs(8180)) or (layer2_outputs(5719)));
    layer3_outputs(9877) <= (layer2_outputs(3851)) and not (layer2_outputs(7842));
    layer3_outputs(9878) <= '1';
    layer3_outputs(9879) <= layer2_outputs(10190);
    layer3_outputs(9880) <= not((layer2_outputs(6200)) or (layer2_outputs(1667)));
    layer3_outputs(9881) <= not(layer2_outputs(9744));
    layer3_outputs(9882) <= '0';
    layer3_outputs(9883) <= layer2_outputs(431);
    layer3_outputs(9884) <= not(layer2_outputs(7017));
    layer3_outputs(9885) <= layer2_outputs(5065);
    layer3_outputs(9886) <= (layer2_outputs(3391)) and (layer2_outputs(6091));
    layer3_outputs(9887) <= layer2_outputs(3197);
    layer3_outputs(9888) <= layer2_outputs(8444);
    layer3_outputs(9889) <= (layer2_outputs(4849)) and (layer2_outputs(8573));
    layer3_outputs(9890) <= not((layer2_outputs(9723)) and (layer2_outputs(2497)));
    layer3_outputs(9891) <= layer2_outputs(826);
    layer3_outputs(9892) <= layer2_outputs(3078);
    layer3_outputs(9893) <= not((layer2_outputs(6122)) and (layer2_outputs(8437)));
    layer3_outputs(9894) <= not(layer2_outputs(163));
    layer3_outputs(9895) <= not(layer2_outputs(29));
    layer3_outputs(9896) <= (layer2_outputs(6842)) or (layer2_outputs(10174));
    layer3_outputs(9897) <= not(layer2_outputs(7162));
    layer3_outputs(9898) <= layer2_outputs(6706);
    layer3_outputs(9899) <= not(layer2_outputs(3821));
    layer3_outputs(9900) <= layer2_outputs(9187);
    layer3_outputs(9901) <= (layer2_outputs(640)) and not (layer2_outputs(7466));
    layer3_outputs(9902) <= layer2_outputs(5056);
    layer3_outputs(9903) <= layer2_outputs(8494);
    layer3_outputs(9904) <= not(layer2_outputs(2799)) or (layer2_outputs(1400));
    layer3_outputs(9905) <= (layer2_outputs(154)) and not (layer2_outputs(174));
    layer3_outputs(9906) <= (layer2_outputs(4062)) and not (layer2_outputs(9880));
    layer3_outputs(9907) <= layer2_outputs(10185);
    layer3_outputs(9908) <= not(layer2_outputs(9152)) or (layer2_outputs(3028));
    layer3_outputs(9909) <= layer2_outputs(1140);
    layer3_outputs(9910) <= layer2_outputs(5203);
    layer3_outputs(9911) <= not((layer2_outputs(696)) or (layer2_outputs(4669)));
    layer3_outputs(9912) <= not(layer2_outputs(8417)) or (layer2_outputs(992));
    layer3_outputs(9913) <= (layer2_outputs(3249)) and (layer2_outputs(681));
    layer3_outputs(9914) <= not(layer2_outputs(4126));
    layer3_outputs(9915) <= layer2_outputs(4372);
    layer3_outputs(9916) <= not(layer2_outputs(2748));
    layer3_outputs(9917) <= not(layer2_outputs(9664)) or (layer2_outputs(5562));
    layer3_outputs(9918) <= layer2_outputs(2889);
    layer3_outputs(9919) <= layer2_outputs(624);
    layer3_outputs(9920) <= layer2_outputs(6265);
    layer3_outputs(9921) <= not(layer2_outputs(5499));
    layer3_outputs(9922) <= layer2_outputs(8489);
    layer3_outputs(9923) <= layer2_outputs(7246);
    layer3_outputs(9924) <= (layer2_outputs(3891)) and not (layer2_outputs(3510));
    layer3_outputs(9925) <= not(layer2_outputs(5921));
    layer3_outputs(9926) <= not(layer2_outputs(211));
    layer3_outputs(9927) <= '1';
    layer3_outputs(9928) <= layer2_outputs(4360);
    layer3_outputs(9929) <= not((layer2_outputs(6870)) and (layer2_outputs(2420)));
    layer3_outputs(9930) <= not(layer2_outputs(4124)) or (layer2_outputs(5314));
    layer3_outputs(9931) <= (layer2_outputs(2651)) or (layer2_outputs(5232));
    layer3_outputs(9932) <= not(layer2_outputs(4802));
    layer3_outputs(9933) <= layer2_outputs(1895);
    layer3_outputs(9934) <= not(layer2_outputs(1347));
    layer3_outputs(9935) <= layer2_outputs(6796);
    layer3_outputs(9936) <= layer2_outputs(9450);
    layer3_outputs(9937) <= not(layer2_outputs(4190));
    layer3_outputs(9938) <= not((layer2_outputs(367)) xor (layer2_outputs(7091)));
    layer3_outputs(9939) <= not((layer2_outputs(8849)) xor (layer2_outputs(9635)));
    layer3_outputs(9940) <= layer2_outputs(1274);
    layer3_outputs(9941) <= not(layer2_outputs(7830));
    layer3_outputs(9942) <= layer2_outputs(146);
    layer3_outputs(9943) <= (layer2_outputs(4997)) or (layer2_outputs(5988));
    layer3_outputs(9944) <= layer2_outputs(4773);
    layer3_outputs(9945) <= not(layer2_outputs(7034));
    layer3_outputs(9946) <= not(layer2_outputs(3761));
    layer3_outputs(9947) <= layer2_outputs(5808);
    layer3_outputs(9948) <= '1';
    layer3_outputs(9949) <= (layer2_outputs(5573)) and not (layer2_outputs(4005));
    layer3_outputs(9950) <= layer2_outputs(5660);
    layer3_outputs(9951) <= not((layer2_outputs(1388)) and (layer2_outputs(5877)));
    layer3_outputs(9952) <= not(layer2_outputs(9497));
    layer3_outputs(9953) <= (layer2_outputs(9219)) xor (layer2_outputs(2092));
    layer3_outputs(9954) <= not((layer2_outputs(8153)) xor (layer2_outputs(5104)));
    layer3_outputs(9955) <= not(layer2_outputs(4952));
    layer3_outputs(9956) <= layer2_outputs(8359);
    layer3_outputs(9957) <= not(layer2_outputs(3174));
    layer3_outputs(9958) <= (layer2_outputs(2283)) and not (layer2_outputs(1549));
    layer3_outputs(9959) <= not(layer2_outputs(9919));
    layer3_outputs(9960) <= not(layer2_outputs(8872));
    layer3_outputs(9961) <= layer2_outputs(42);
    layer3_outputs(9962) <= layer2_outputs(6997);
    layer3_outputs(9963) <= not(layer2_outputs(9520));
    layer3_outputs(9964) <= not(layer2_outputs(5969));
    layer3_outputs(9965) <= layer2_outputs(2082);
    layer3_outputs(9966) <= (layer2_outputs(5725)) or (layer2_outputs(8225));
    layer3_outputs(9967) <= not(layer2_outputs(2143));
    layer3_outputs(9968) <= not(layer2_outputs(4304));
    layer3_outputs(9969) <= '1';
    layer3_outputs(9970) <= layer2_outputs(8119);
    layer3_outputs(9971) <= layer2_outputs(4820);
    layer3_outputs(9972) <= (layer2_outputs(2174)) xor (layer2_outputs(7916));
    layer3_outputs(9973) <= not(layer2_outputs(4909));
    layer3_outputs(9974) <= layer2_outputs(1713);
    layer3_outputs(9975) <= not(layer2_outputs(9955));
    layer3_outputs(9976) <= not(layer2_outputs(1852));
    layer3_outputs(9977) <= not(layer2_outputs(5508));
    layer3_outputs(9978) <= (layer2_outputs(3690)) and not (layer2_outputs(6556));
    layer3_outputs(9979) <= (layer2_outputs(617)) and not (layer2_outputs(8326));
    layer3_outputs(9980) <= layer2_outputs(6555);
    layer3_outputs(9981) <= layer2_outputs(8247);
    layer3_outputs(9982) <= not((layer2_outputs(4719)) xor (layer2_outputs(9188)));
    layer3_outputs(9983) <= not(layer2_outputs(3852));
    layer3_outputs(9984) <= not(layer2_outputs(3639));
    layer3_outputs(9985) <= layer2_outputs(4604);
    layer3_outputs(9986) <= not(layer2_outputs(3155));
    layer3_outputs(9987) <= not(layer2_outputs(6001));
    layer3_outputs(9988) <= '1';
    layer3_outputs(9989) <= layer2_outputs(953);
    layer3_outputs(9990) <= (layer2_outputs(3479)) or (layer2_outputs(4251));
    layer3_outputs(9991) <= layer2_outputs(1132);
    layer3_outputs(9992) <= layer2_outputs(2013);
    layer3_outputs(9993) <= layer2_outputs(7180);
    layer3_outputs(9994) <= layer2_outputs(5778);
    layer3_outputs(9995) <= not(layer2_outputs(8997));
    layer3_outputs(9996) <= (layer2_outputs(6986)) or (layer2_outputs(7369));
    layer3_outputs(9997) <= layer2_outputs(5617);
    layer3_outputs(9998) <= layer2_outputs(6973);
    layer3_outputs(9999) <= not((layer2_outputs(4536)) and (layer2_outputs(4524)));
    layer3_outputs(10000) <= (layer2_outputs(9158)) or (layer2_outputs(2341));
    layer3_outputs(10001) <= not(layer2_outputs(4869)) or (layer2_outputs(3195));
    layer3_outputs(10002) <= (layer2_outputs(3060)) and (layer2_outputs(9687));
    layer3_outputs(10003) <= not((layer2_outputs(2819)) xor (layer2_outputs(1966)));
    layer3_outputs(10004) <= '0';
    layer3_outputs(10005) <= layer2_outputs(5309);
    layer3_outputs(10006) <= (layer2_outputs(7816)) or (layer2_outputs(6826));
    layer3_outputs(10007) <= not(layer2_outputs(1389));
    layer3_outputs(10008) <= (layer2_outputs(3648)) and (layer2_outputs(447));
    layer3_outputs(10009) <= not(layer2_outputs(2601));
    layer3_outputs(10010) <= layer2_outputs(7148);
    layer3_outputs(10011) <= not(layer2_outputs(6502)) or (layer2_outputs(282));
    layer3_outputs(10012) <= (layer2_outputs(6290)) xor (layer2_outputs(4093));
    layer3_outputs(10013) <= layer2_outputs(4854);
    layer3_outputs(10014) <= not(layer2_outputs(6453));
    layer3_outputs(10015) <= not((layer2_outputs(2109)) and (layer2_outputs(2726)));
    layer3_outputs(10016) <= not(layer2_outputs(9828));
    layer3_outputs(10017) <= not((layer2_outputs(3454)) and (layer2_outputs(8445)));
    layer3_outputs(10018) <= not(layer2_outputs(3105));
    layer3_outputs(10019) <= not((layer2_outputs(6392)) xor (layer2_outputs(476)));
    layer3_outputs(10020) <= not(layer2_outputs(8305));
    layer3_outputs(10021) <= not((layer2_outputs(5862)) xor (layer2_outputs(10092)));
    layer3_outputs(10022) <= '1';
    layer3_outputs(10023) <= layer2_outputs(9992);
    layer3_outputs(10024) <= not(layer2_outputs(4566));
    layer3_outputs(10025) <= layer2_outputs(1595);
    layer3_outputs(10026) <= not((layer2_outputs(1503)) and (layer2_outputs(6399)));
    layer3_outputs(10027) <= layer2_outputs(8187);
    layer3_outputs(10028) <= not(layer2_outputs(3616));
    layer3_outputs(10029) <= layer2_outputs(1425);
    layer3_outputs(10030) <= layer2_outputs(1018);
    layer3_outputs(10031) <= layer2_outputs(8955);
    layer3_outputs(10032) <= not(layer2_outputs(6658));
    layer3_outputs(10033) <= layer2_outputs(5810);
    layer3_outputs(10034) <= layer2_outputs(7095);
    layer3_outputs(10035) <= (layer2_outputs(7021)) xor (layer2_outputs(8859));
    layer3_outputs(10036) <= not((layer2_outputs(4759)) or (layer2_outputs(1342)));
    layer3_outputs(10037) <= layer2_outputs(2207);
    layer3_outputs(10038) <= layer2_outputs(8594);
    layer3_outputs(10039) <= (layer2_outputs(8543)) and (layer2_outputs(5206));
    layer3_outputs(10040) <= layer2_outputs(1566);
    layer3_outputs(10041) <= not(layer2_outputs(7802)) or (layer2_outputs(6252));
    layer3_outputs(10042) <= not(layer2_outputs(7966));
    layer3_outputs(10043) <= not(layer2_outputs(2328)) or (layer2_outputs(3907));
    layer3_outputs(10044) <= not(layer2_outputs(8603));
    layer3_outputs(10045) <= '0';
    layer3_outputs(10046) <= not(layer2_outputs(245)) or (layer2_outputs(7226));
    layer3_outputs(10047) <= not(layer2_outputs(2244)) or (layer2_outputs(1812));
    layer3_outputs(10048) <= not((layer2_outputs(6721)) and (layer2_outputs(9324)));
    layer3_outputs(10049) <= not(layer2_outputs(4798)) or (layer2_outputs(8735));
    layer3_outputs(10050) <= (layer2_outputs(4469)) and not (layer2_outputs(6266));
    layer3_outputs(10051) <= layer2_outputs(5123);
    layer3_outputs(10052) <= layer2_outputs(9253);
    layer3_outputs(10053) <= not((layer2_outputs(3164)) or (layer2_outputs(4471)));
    layer3_outputs(10054) <= not(layer2_outputs(7003));
    layer3_outputs(10055) <= not(layer2_outputs(6031)) or (layer2_outputs(9193));
    layer3_outputs(10056) <= layer2_outputs(7015);
    layer3_outputs(10057) <= not(layer2_outputs(7522)) or (layer2_outputs(564));
    layer3_outputs(10058) <= not((layer2_outputs(4926)) and (layer2_outputs(9688)));
    layer3_outputs(10059) <= (layer2_outputs(445)) xor (layer2_outputs(986));
    layer3_outputs(10060) <= not(layer2_outputs(686));
    layer3_outputs(10061) <= not(layer2_outputs(10227));
    layer3_outputs(10062) <= layer2_outputs(1672);
    layer3_outputs(10063) <= layer2_outputs(1724);
    layer3_outputs(10064) <= layer2_outputs(2942);
    layer3_outputs(10065) <= not((layer2_outputs(7640)) xor (layer2_outputs(6970)));
    layer3_outputs(10066) <= (layer2_outputs(9522)) and not (layer2_outputs(5127));
    layer3_outputs(10067) <= (layer2_outputs(5267)) and not (layer2_outputs(4784));
    layer3_outputs(10068) <= not(layer2_outputs(3219)) or (layer2_outputs(7859));
    layer3_outputs(10069) <= not((layer2_outputs(8874)) xor (layer2_outputs(990)));
    layer3_outputs(10070) <= not((layer2_outputs(1224)) or (layer2_outputs(6187)));
    layer3_outputs(10071) <= not(layer2_outputs(4911)) or (layer2_outputs(8234));
    layer3_outputs(10072) <= not((layer2_outputs(5446)) or (layer2_outputs(4965)));
    layer3_outputs(10073) <= layer2_outputs(9299);
    layer3_outputs(10074) <= not(layer2_outputs(8742));
    layer3_outputs(10075) <= layer2_outputs(5138);
    layer3_outputs(10076) <= layer2_outputs(9387);
    layer3_outputs(10077) <= layer2_outputs(257);
    layer3_outputs(10078) <= (layer2_outputs(10228)) or (layer2_outputs(1103));
    layer3_outputs(10079) <= not(layer2_outputs(10047)) or (layer2_outputs(2148));
    layer3_outputs(10080) <= layer2_outputs(261);
    layer3_outputs(10081) <= not(layer2_outputs(8179));
    layer3_outputs(10082) <= '1';
    layer3_outputs(10083) <= not(layer2_outputs(1063));
    layer3_outputs(10084) <= not((layer2_outputs(9353)) or (layer2_outputs(6802)));
    layer3_outputs(10085) <= not((layer2_outputs(2534)) and (layer2_outputs(3538)));
    layer3_outputs(10086) <= not((layer2_outputs(3334)) and (layer2_outputs(6561)));
    layer3_outputs(10087) <= (layer2_outputs(6289)) xor (layer2_outputs(8916));
    layer3_outputs(10088) <= layer2_outputs(3446);
    layer3_outputs(10089) <= (layer2_outputs(4687)) xor (layer2_outputs(1708));
    layer3_outputs(10090) <= '0';
    layer3_outputs(10091) <= not(layer2_outputs(8336));
    layer3_outputs(10092) <= not((layer2_outputs(4330)) xor (layer2_outputs(9761)));
    layer3_outputs(10093) <= not(layer2_outputs(2472));
    layer3_outputs(10094) <= not(layer2_outputs(7223));
    layer3_outputs(10095) <= not(layer2_outputs(6134)) or (layer2_outputs(6141));
    layer3_outputs(10096) <= '0';
    layer3_outputs(10097) <= layer2_outputs(3676);
    layer3_outputs(10098) <= not((layer2_outputs(6540)) and (layer2_outputs(4991)));
    layer3_outputs(10099) <= not((layer2_outputs(9978)) and (layer2_outputs(3170)));
    layer3_outputs(10100) <= layer2_outputs(3916);
    layer3_outputs(10101) <= not(layer2_outputs(7495));
    layer3_outputs(10102) <= not(layer2_outputs(5865));
    layer3_outputs(10103) <= '1';
    layer3_outputs(10104) <= not(layer2_outputs(10208));
    layer3_outputs(10105) <= not(layer2_outputs(336));
    layer3_outputs(10106) <= not((layer2_outputs(556)) and (layer2_outputs(1918)));
    layer3_outputs(10107) <= not(layer2_outputs(9333));
    layer3_outputs(10108) <= layer2_outputs(3146);
    layer3_outputs(10109) <= layer2_outputs(6446);
    layer3_outputs(10110) <= not(layer2_outputs(6583));
    layer3_outputs(10111) <= not(layer2_outputs(4030));
    layer3_outputs(10112) <= (layer2_outputs(6237)) or (layer2_outputs(9532));
    layer3_outputs(10113) <= layer2_outputs(1033);
    layer3_outputs(10114) <= (layer2_outputs(502)) and (layer2_outputs(6834));
    layer3_outputs(10115) <= (layer2_outputs(6117)) and not (layer2_outputs(9145));
    layer3_outputs(10116) <= not(layer2_outputs(5103)) or (layer2_outputs(5410));
    layer3_outputs(10117) <= (layer2_outputs(9438)) xor (layer2_outputs(7271));
    layer3_outputs(10118) <= not(layer2_outputs(8618));
    layer3_outputs(10119) <= not((layer2_outputs(592)) and (layer2_outputs(8698)));
    layer3_outputs(10120) <= (layer2_outputs(3528)) and not (layer2_outputs(4629));
    layer3_outputs(10121) <= (layer2_outputs(6565)) and (layer2_outputs(10090));
    layer3_outputs(10122) <= layer2_outputs(4543);
    layer3_outputs(10123) <= layer2_outputs(9690);
    layer3_outputs(10124) <= (layer2_outputs(1656)) and not (layer2_outputs(3746));
    layer3_outputs(10125) <= not(layer2_outputs(2323));
    layer3_outputs(10126) <= (layer2_outputs(4325)) and (layer2_outputs(1961));
    layer3_outputs(10127) <= not(layer2_outputs(637));
    layer3_outputs(10128) <= not((layer2_outputs(6020)) xor (layer2_outputs(1409)));
    layer3_outputs(10129) <= not(layer2_outputs(1564));
    layer3_outputs(10130) <= not(layer2_outputs(8912));
    layer3_outputs(10131) <= not(layer2_outputs(6692));
    layer3_outputs(10132) <= not(layer2_outputs(10021));
    layer3_outputs(10133) <= not(layer2_outputs(7370));
    layer3_outputs(10134) <= layer2_outputs(4708);
    layer3_outputs(10135) <= layer2_outputs(4649);
    layer3_outputs(10136) <= (layer2_outputs(2535)) or (layer2_outputs(7244));
    layer3_outputs(10137) <= layer2_outputs(5299);
    layer3_outputs(10138) <= not(layer2_outputs(3109)) or (layer2_outputs(9894));
    layer3_outputs(10139) <= layer2_outputs(4491);
    layer3_outputs(10140) <= layer2_outputs(962);
    layer3_outputs(10141) <= (layer2_outputs(1606)) and not (layer2_outputs(9635));
    layer3_outputs(10142) <= (layer2_outputs(5533)) or (layer2_outputs(3296));
    layer3_outputs(10143) <= layer2_outputs(5996);
    layer3_outputs(10144) <= (layer2_outputs(8686)) or (layer2_outputs(5967));
    layer3_outputs(10145) <= not((layer2_outputs(8746)) and (layer2_outputs(6736)));
    layer3_outputs(10146) <= layer2_outputs(5302);
    layer3_outputs(10147) <= layer2_outputs(7022);
    layer3_outputs(10148) <= not(layer2_outputs(2338));
    layer3_outputs(10149) <= not(layer2_outputs(7098));
    layer3_outputs(10150) <= not(layer2_outputs(2236)) or (layer2_outputs(1376));
    layer3_outputs(10151) <= not(layer2_outputs(9532));
    layer3_outputs(10152) <= not((layer2_outputs(2452)) and (layer2_outputs(4280)));
    layer3_outputs(10153) <= not(layer2_outputs(4092));
    layer3_outputs(10154) <= (layer2_outputs(5608)) or (layer2_outputs(3232));
    layer3_outputs(10155) <= not(layer2_outputs(5402));
    layer3_outputs(10156) <= layer2_outputs(4661);
    layer3_outputs(10157) <= not(layer2_outputs(6441));
    layer3_outputs(10158) <= not(layer2_outputs(6537));
    layer3_outputs(10159) <= layer2_outputs(3922);
    layer3_outputs(10160) <= layer2_outputs(6594);
    layer3_outputs(10161) <= not(layer2_outputs(5373));
    layer3_outputs(10162) <= not((layer2_outputs(3396)) or (layer2_outputs(1234)));
    layer3_outputs(10163) <= layer2_outputs(7334);
    layer3_outputs(10164) <= not(layer2_outputs(551)) or (layer2_outputs(9618));
    layer3_outputs(10165) <= not(layer2_outputs(7209));
    layer3_outputs(10166) <= layer2_outputs(6562);
    layer3_outputs(10167) <= '1';
    layer3_outputs(10168) <= layer2_outputs(3351);
    layer3_outputs(10169) <= (layer2_outputs(9437)) xor (layer2_outputs(3008));
    layer3_outputs(10170) <= not(layer2_outputs(10063));
    layer3_outputs(10171) <= not((layer2_outputs(4826)) or (layer2_outputs(4048)));
    layer3_outputs(10172) <= '1';
    layer3_outputs(10173) <= (layer2_outputs(7851)) and not (layer2_outputs(1069));
    layer3_outputs(10174) <= layer2_outputs(9244);
    layer3_outputs(10175) <= not((layer2_outputs(3817)) or (layer2_outputs(5062)));
    layer3_outputs(10176) <= (layer2_outputs(2352)) and not (layer2_outputs(9496));
    layer3_outputs(10177) <= not(layer2_outputs(5788));
    layer3_outputs(10178) <= not(layer2_outputs(1809));
    layer3_outputs(10179) <= layer2_outputs(6581);
    layer3_outputs(10180) <= not((layer2_outputs(9022)) and (layer2_outputs(827)));
    layer3_outputs(10181) <= not((layer2_outputs(1475)) xor (layer2_outputs(7305)));
    layer3_outputs(10182) <= not(layer2_outputs(4941));
    layer3_outputs(10183) <= not(layer2_outputs(1026));
    layer3_outputs(10184) <= not(layer2_outputs(7817)) or (layer2_outputs(8944));
    layer3_outputs(10185) <= not(layer2_outputs(547)) or (layer2_outputs(9686));
    layer3_outputs(10186) <= (layer2_outputs(3884)) and not (layer2_outputs(5125));
    layer3_outputs(10187) <= layer2_outputs(6418);
    layer3_outputs(10188) <= (layer2_outputs(883)) and not (layer2_outputs(7116));
    layer3_outputs(10189) <= layer2_outputs(5393);
    layer3_outputs(10190) <= not(layer2_outputs(2121));
    layer3_outputs(10191) <= not(layer2_outputs(6705));
    layer3_outputs(10192) <= '1';
    layer3_outputs(10193) <= (layer2_outputs(5443)) and (layer2_outputs(2256));
    layer3_outputs(10194) <= '0';
    layer3_outputs(10195) <= not((layer2_outputs(6178)) xor (layer2_outputs(431)));
    layer3_outputs(10196) <= not((layer2_outputs(10193)) xor (layer2_outputs(3458)));
    layer3_outputs(10197) <= layer2_outputs(8322);
    layer3_outputs(10198) <= layer2_outputs(1151);
    layer3_outputs(10199) <= not(layer2_outputs(5819));
    layer3_outputs(10200) <= (layer2_outputs(3924)) or (layer2_outputs(7262));
    layer3_outputs(10201) <= not((layer2_outputs(3361)) and (layer2_outputs(1465)));
    layer3_outputs(10202) <= not(layer2_outputs(4881));
    layer3_outputs(10203) <= (layer2_outputs(4212)) xor (layer2_outputs(2801));
    layer3_outputs(10204) <= not(layer2_outputs(8599));
    layer3_outputs(10205) <= not(layer2_outputs(150));
    layer3_outputs(10206) <= not((layer2_outputs(573)) and (layer2_outputs(8348)));
    layer3_outputs(10207) <= not(layer2_outputs(693));
    layer3_outputs(10208) <= layer2_outputs(1309);
    layer3_outputs(10209) <= layer2_outputs(7948);
    layer3_outputs(10210) <= not(layer2_outputs(9166));
    layer3_outputs(10211) <= (layer2_outputs(5713)) xor (layer2_outputs(7076));
    layer3_outputs(10212) <= (layer2_outputs(9257)) xor (layer2_outputs(9516));
    layer3_outputs(10213) <= not(layer2_outputs(277));
    layer3_outputs(10214) <= (layer2_outputs(10074)) and not (layer2_outputs(8831));
    layer3_outputs(10215) <= (layer2_outputs(5962)) or (layer2_outputs(2579));
    layer3_outputs(10216) <= not(layer2_outputs(462));
    layer3_outputs(10217) <= layer2_outputs(8578);
    layer3_outputs(10218) <= (layer2_outputs(3534)) or (layer2_outputs(6400));
    layer3_outputs(10219) <= layer2_outputs(2150);
    layer3_outputs(10220) <= not(layer2_outputs(9669)) or (layer2_outputs(5383));
    layer3_outputs(10221) <= '1';
    layer3_outputs(10222) <= (layer2_outputs(9166)) or (layer2_outputs(5486));
    layer3_outputs(10223) <= not(layer2_outputs(7883));
    layer3_outputs(10224) <= (layer2_outputs(2201)) and not (layer2_outputs(9739));
    layer3_outputs(10225) <= not(layer2_outputs(5218));
    layer3_outputs(10226) <= '1';
    layer3_outputs(10227) <= not(layer2_outputs(1143));
    layer3_outputs(10228) <= (layer2_outputs(10005)) xor (layer2_outputs(3681));
    layer3_outputs(10229) <= (layer2_outputs(6776)) and not (layer2_outputs(1437));
    layer3_outputs(10230) <= layer2_outputs(5293);
    layer3_outputs(10231) <= (layer2_outputs(1554)) and (layer2_outputs(9421));
    layer3_outputs(10232) <= layer2_outputs(3002);
    layer3_outputs(10233) <= not((layer2_outputs(298)) or (layer2_outputs(6384)));
    layer3_outputs(10234) <= not((layer2_outputs(516)) or (layer2_outputs(5607)));
    layer3_outputs(10235) <= (layer2_outputs(8677)) and not (layer2_outputs(180));
    layer3_outputs(10236) <= not(layer2_outputs(2670)) or (layer2_outputs(7256));
    layer3_outputs(10237) <= layer2_outputs(3385);
    layer3_outputs(10238) <= (layer2_outputs(7554)) and (layer2_outputs(4166));
    layer3_outputs(10239) <= (layer2_outputs(2864)) and not (layer2_outputs(2600));
    layer4_outputs(0) <= '1';
    layer4_outputs(1) <= (layer3_outputs(1421)) xor (layer3_outputs(4009));
    layer4_outputs(2) <= not(layer3_outputs(6633)) or (layer3_outputs(10006));
    layer4_outputs(3) <= not(layer3_outputs(2386));
    layer4_outputs(4) <= not(layer3_outputs(1797));
    layer4_outputs(5) <= (layer3_outputs(5197)) xor (layer3_outputs(2739));
    layer4_outputs(6) <= not(layer3_outputs(9078));
    layer4_outputs(7) <= layer3_outputs(6334);
    layer4_outputs(8) <= not(layer3_outputs(8897)) or (layer3_outputs(6524));
    layer4_outputs(9) <= not(layer3_outputs(7008));
    layer4_outputs(10) <= (layer3_outputs(9751)) and not (layer3_outputs(357));
    layer4_outputs(11) <= not(layer3_outputs(5156));
    layer4_outputs(12) <= layer3_outputs(1579);
    layer4_outputs(13) <= layer3_outputs(2674);
    layer4_outputs(14) <= not(layer3_outputs(6343));
    layer4_outputs(15) <= not((layer3_outputs(2923)) xor (layer3_outputs(8753)));
    layer4_outputs(16) <= not(layer3_outputs(1798));
    layer4_outputs(17) <= layer3_outputs(2490);
    layer4_outputs(18) <= (layer3_outputs(6289)) xor (layer3_outputs(9136));
    layer4_outputs(19) <= '1';
    layer4_outputs(20) <= not(layer3_outputs(8518));
    layer4_outputs(21) <= not((layer3_outputs(6942)) xor (layer3_outputs(5949)));
    layer4_outputs(22) <= not(layer3_outputs(5422)) or (layer3_outputs(434));
    layer4_outputs(23) <= not(layer3_outputs(7297));
    layer4_outputs(24) <= layer3_outputs(5973);
    layer4_outputs(25) <= (layer3_outputs(3992)) xor (layer3_outputs(3789));
    layer4_outputs(26) <= layer3_outputs(6795);
    layer4_outputs(27) <= not(layer3_outputs(7205));
    layer4_outputs(28) <= not(layer3_outputs(2293));
    layer4_outputs(29) <= not(layer3_outputs(8314));
    layer4_outputs(30) <= layer3_outputs(5587);
    layer4_outputs(31) <= not(layer3_outputs(6980));
    layer4_outputs(32) <= layer3_outputs(6828);
    layer4_outputs(33) <= (layer3_outputs(4480)) xor (layer3_outputs(5523));
    layer4_outputs(34) <= (layer3_outputs(8099)) and not (layer3_outputs(5072));
    layer4_outputs(35) <= layer3_outputs(7151);
    layer4_outputs(36) <= (layer3_outputs(8087)) and (layer3_outputs(7586));
    layer4_outputs(37) <= layer3_outputs(8215);
    layer4_outputs(38) <= layer3_outputs(7288);
    layer4_outputs(39) <= not(layer3_outputs(2779));
    layer4_outputs(40) <= layer3_outputs(3106);
    layer4_outputs(41) <= not(layer3_outputs(9057));
    layer4_outputs(42) <= not(layer3_outputs(4731));
    layer4_outputs(43) <= not(layer3_outputs(2044));
    layer4_outputs(44) <= '0';
    layer4_outputs(45) <= (layer3_outputs(4937)) and not (layer3_outputs(425));
    layer4_outputs(46) <= not((layer3_outputs(382)) xor (layer3_outputs(4789)));
    layer4_outputs(47) <= not(layer3_outputs(9658));
    layer4_outputs(48) <= not((layer3_outputs(5936)) xor (layer3_outputs(4396)));
    layer4_outputs(49) <= not(layer3_outputs(259));
    layer4_outputs(50) <= '0';
    layer4_outputs(51) <= not(layer3_outputs(8536));
    layer4_outputs(52) <= not(layer3_outputs(7232));
    layer4_outputs(53) <= (layer3_outputs(1637)) xor (layer3_outputs(9218));
    layer4_outputs(54) <= not((layer3_outputs(5328)) and (layer3_outputs(9032)));
    layer4_outputs(55) <= not(layer3_outputs(2616));
    layer4_outputs(56) <= layer3_outputs(5108);
    layer4_outputs(57) <= not((layer3_outputs(5528)) xor (layer3_outputs(8517)));
    layer4_outputs(58) <= not(layer3_outputs(5487));
    layer4_outputs(59) <= (layer3_outputs(7799)) xor (layer3_outputs(9749));
    layer4_outputs(60) <= not(layer3_outputs(4410)) or (layer3_outputs(6256));
    layer4_outputs(61) <= not(layer3_outputs(2761));
    layer4_outputs(62) <= not(layer3_outputs(10112));
    layer4_outputs(63) <= layer3_outputs(3319);
    layer4_outputs(64) <= not(layer3_outputs(7998)) or (layer3_outputs(1891));
    layer4_outputs(65) <= not(layer3_outputs(9038)) or (layer3_outputs(9669));
    layer4_outputs(66) <= (layer3_outputs(5948)) and not (layer3_outputs(9546));
    layer4_outputs(67) <= not((layer3_outputs(4810)) or (layer3_outputs(8095)));
    layer4_outputs(68) <= '0';
    layer4_outputs(69) <= not(layer3_outputs(5077));
    layer4_outputs(70) <= not((layer3_outputs(9092)) xor (layer3_outputs(5015)));
    layer4_outputs(71) <= not(layer3_outputs(2342));
    layer4_outputs(72) <= layer3_outputs(6257);
    layer4_outputs(73) <= (layer3_outputs(4371)) and (layer3_outputs(5358));
    layer4_outputs(74) <= not(layer3_outputs(1395));
    layer4_outputs(75) <= not(layer3_outputs(7387));
    layer4_outputs(76) <= not(layer3_outputs(681));
    layer4_outputs(77) <= (layer3_outputs(7608)) and (layer3_outputs(773));
    layer4_outputs(78) <= layer3_outputs(5259);
    layer4_outputs(79) <= layer3_outputs(7942);
    layer4_outputs(80) <= not(layer3_outputs(5503)) or (layer3_outputs(524));
    layer4_outputs(81) <= (layer3_outputs(8741)) or (layer3_outputs(2207));
    layer4_outputs(82) <= not(layer3_outputs(5388)) or (layer3_outputs(356));
    layer4_outputs(83) <= not((layer3_outputs(2549)) xor (layer3_outputs(6167)));
    layer4_outputs(84) <= not(layer3_outputs(8785));
    layer4_outputs(85) <= (layer3_outputs(4470)) and (layer3_outputs(8102));
    layer4_outputs(86) <= not(layer3_outputs(4724));
    layer4_outputs(87) <= not((layer3_outputs(7652)) xor (layer3_outputs(742)));
    layer4_outputs(88) <= not(layer3_outputs(9992));
    layer4_outputs(89) <= (layer3_outputs(6800)) xor (layer3_outputs(8180));
    layer4_outputs(90) <= (layer3_outputs(1727)) xor (layer3_outputs(1487));
    layer4_outputs(91) <= (layer3_outputs(362)) or (layer3_outputs(6796));
    layer4_outputs(92) <= not(layer3_outputs(5963));
    layer4_outputs(93) <= not(layer3_outputs(3482));
    layer4_outputs(94) <= (layer3_outputs(2627)) and not (layer3_outputs(1376));
    layer4_outputs(95) <= not(layer3_outputs(9005));
    layer4_outputs(96) <= layer3_outputs(3340);
    layer4_outputs(97) <= not(layer3_outputs(2769));
    layer4_outputs(98) <= layer3_outputs(7773);
    layer4_outputs(99) <= layer3_outputs(8145);
    layer4_outputs(100) <= (layer3_outputs(7647)) xor (layer3_outputs(9876));
    layer4_outputs(101) <= (layer3_outputs(7088)) and not (layer3_outputs(2461));
    layer4_outputs(102) <= (layer3_outputs(2933)) and not (layer3_outputs(4048));
    layer4_outputs(103) <= not(layer3_outputs(4391));
    layer4_outputs(104) <= not((layer3_outputs(7217)) or (layer3_outputs(2130)));
    layer4_outputs(105) <= layer3_outputs(5214);
    layer4_outputs(106) <= layer3_outputs(1205);
    layer4_outputs(107) <= layer3_outputs(1677);
    layer4_outputs(108) <= not(layer3_outputs(10205)) or (layer3_outputs(3408));
    layer4_outputs(109) <= (layer3_outputs(8834)) and not (layer3_outputs(7866));
    layer4_outputs(110) <= (layer3_outputs(6672)) or (layer3_outputs(6493));
    layer4_outputs(111) <= not(layer3_outputs(10150));
    layer4_outputs(112) <= (layer3_outputs(7614)) and not (layer3_outputs(5047));
    layer4_outputs(113) <= not((layer3_outputs(4117)) xor (layer3_outputs(3472)));
    layer4_outputs(114) <= not((layer3_outputs(9794)) xor (layer3_outputs(5625)));
    layer4_outputs(115) <= layer3_outputs(8040);
    layer4_outputs(116) <= not((layer3_outputs(9612)) xor (layer3_outputs(9563)));
    layer4_outputs(117) <= not((layer3_outputs(8157)) xor (layer3_outputs(7617)));
    layer4_outputs(118) <= layer3_outputs(4800);
    layer4_outputs(119) <= layer3_outputs(997);
    layer4_outputs(120) <= (layer3_outputs(6140)) xor (layer3_outputs(3308));
    layer4_outputs(121) <= not((layer3_outputs(4243)) xor (layer3_outputs(3815)));
    layer4_outputs(122) <= layer3_outputs(1329);
    layer4_outputs(123) <= not(layer3_outputs(6639)) or (layer3_outputs(9548));
    layer4_outputs(124) <= not(layer3_outputs(7122)) or (layer3_outputs(1082));
    layer4_outputs(125) <= layer3_outputs(6600);
    layer4_outputs(126) <= not((layer3_outputs(383)) xor (layer3_outputs(3310)));
    layer4_outputs(127) <= '1';
    layer4_outputs(128) <= not(layer3_outputs(1264)) or (layer3_outputs(7385));
    layer4_outputs(129) <= layer3_outputs(177);
    layer4_outputs(130) <= not(layer3_outputs(2566));
    layer4_outputs(131) <= not(layer3_outputs(258));
    layer4_outputs(132) <= (layer3_outputs(9148)) and (layer3_outputs(8960));
    layer4_outputs(133) <= not(layer3_outputs(3074)) or (layer3_outputs(2520));
    layer4_outputs(134) <= not(layer3_outputs(2465));
    layer4_outputs(135) <= not(layer3_outputs(8516));
    layer4_outputs(136) <= (layer3_outputs(5939)) xor (layer3_outputs(262));
    layer4_outputs(137) <= not(layer3_outputs(6828));
    layer4_outputs(138) <= layer3_outputs(505);
    layer4_outputs(139) <= not(layer3_outputs(4495)) or (layer3_outputs(2112));
    layer4_outputs(140) <= (layer3_outputs(3120)) and (layer3_outputs(10181));
    layer4_outputs(141) <= (layer3_outputs(3335)) or (layer3_outputs(2330));
    layer4_outputs(142) <= not(layer3_outputs(3460));
    layer4_outputs(143) <= (layer3_outputs(10131)) xor (layer3_outputs(3716));
    layer4_outputs(144) <= (layer3_outputs(5468)) xor (layer3_outputs(6681));
    layer4_outputs(145) <= layer3_outputs(5594);
    layer4_outputs(146) <= not((layer3_outputs(7271)) xor (layer3_outputs(9360)));
    layer4_outputs(147) <= not(layer3_outputs(4501)) or (layer3_outputs(3815));
    layer4_outputs(148) <= (layer3_outputs(7325)) and (layer3_outputs(9940));
    layer4_outputs(149) <= (layer3_outputs(751)) and not (layer3_outputs(7506));
    layer4_outputs(150) <= (layer3_outputs(9769)) and not (layer3_outputs(5061));
    layer4_outputs(151) <= layer3_outputs(2806);
    layer4_outputs(152) <= (layer3_outputs(1494)) xor (layer3_outputs(10118));
    layer4_outputs(153) <= layer3_outputs(6821);
    layer4_outputs(154) <= (layer3_outputs(1467)) or (layer3_outputs(178));
    layer4_outputs(155) <= not(layer3_outputs(4313));
    layer4_outputs(156) <= layer3_outputs(3472);
    layer4_outputs(157) <= not((layer3_outputs(8663)) xor (layer3_outputs(5415)));
    layer4_outputs(158) <= not(layer3_outputs(3075));
    layer4_outputs(159) <= (layer3_outputs(8501)) and not (layer3_outputs(5352));
    layer4_outputs(160) <= (layer3_outputs(4211)) xor (layer3_outputs(7409));
    layer4_outputs(161) <= not(layer3_outputs(4361));
    layer4_outputs(162) <= not((layer3_outputs(8597)) xor (layer3_outputs(48)));
    layer4_outputs(163) <= layer3_outputs(3025);
    layer4_outputs(164) <= not((layer3_outputs(4014)) and (layer3_outputs(2358)));
    layer4_outputs(165) <= not((layer3_outputs(6521)) and (layer3_outputs(6567)));
    layer4_outputs(166) <= not(layer3_outputs(6404));
    layer4_outputs(167) <= not(layer3_outputs(8760));
    layer4_outputs(168) <= (layer3_outputs(6682)) and (layer3_outputs(4278));
    layer4_outputs(169) <= (layer3_outputs(3553)) and not (layer3_outputs(3271));
    layer4_outputs(170) <= layer3_outputs(1024);
    layer4_outputs(171) <= not(layer3_outputs(7940)) or (layer3_outputs(3326));
    layer4_outputs(172) <= not(layer3_outputs(4476));
    layer4_outputs(173) <= (layer3_outputs(9335)) or (layer3_outputs(5243));
    layer4_outputs(174) <= layer3_outputs(9573);
    layer4_outputs(175) <= not(layer3_outputs(1380));
    layer4_outputs(176) <= (layer3_outputs(2065)) or (layer3_outputs(2197));
    layer4_outputs(177) <= not(layer3_outputs(4022));
    layer4_outputs(178) <= layer3_outputs(7126);
    layer4_outputs(179) <= (layer3_outputs(6682)) and (layer3_outputs(1009));
    layer4_outputs(180) <= (layer3_outputs(2733)) xor (layer3_outputs(63));
    layer4_outputs(181) <= not(layer3_outputs(6094));
    layer4_outputs(182) <= not(layer3_outputs(151));
    layer4_outputs(183) <= not(layer3_outputs(2568));
    layer4_outputs(184) <= not((layer3_outputs(183)) xor (layer3_outputs(3606)));
    layer4_outputs(185) <= layer3_outputs(7423);
    layer4_outputs(186) <= layer3_outputs(1337);
    layer4_outputs(187) <= not(layer3_outputs(3039)) or (layer3_outputs(5006));
    layer4_outputs(188) <= (layer3_outputs(4412)) and not (layer3_outputs(4366));
    layer4_outputs(189) <= layer3_outputs(7176);
    layer4_outputs(190) <= layer3_outputs(7675);
    layer4_outputs(191) <= not(layer3_outputs(6668));
    layer4_outputs(192) <= not((layer3_outputs(4214)) or (layer3_outputs(9325)));
    layer4_outputs(193) <= layer3_outputs(6707);
    layer4_outputs(194) <= (layer3_outputs(619)) xor (layer3_outputs(4301));
    layer4_outputs(195) <= not(layer3_outputs(3037));
    layer4_outputs(196) <= not(layer3_outputs(3009));
    layer4_outputs(197) <= layer3_outputs(1850);
    layer4_outputs(198) <= layer3_outputs(4191);
    layer4_outputs(199) <= not(layer3_outputs(5429));
    layer4_outputs(200) <= not(layer3_outputs(6491));
    layer4_outputs(201) <= not((layer3_outputs(3877)) or (layer3_outputs(1037)));
    layer4_outputs(202) <= not((layer3_outputs(6642)) xor (layer3_outputs(7162)));
    layer4_outputs(203) <= layer3_outputs(4048);
    layer4_outputs(204) <= layer3_outputs(9242);
    layer4_outputs(205) <= (layer3_outputs(3563)) or (layer3_outputs(8981));
    layer4_outputs(206) <= (layer3_outputs(5942)) and not (layer3_outputs(7696));
    layer4_outputs(207) <= (layer3_outputs(2075)) and (layer3_outputs(2678));
    layer4_outputs(208) <= not((layer3_outputs(3628)) and (layer3_outputs(4294)));
    layer4_outputs(209) <= not(layer3_outputs(7321));
    layer4_outputs(210) <= not(layer3_outputs(2938));
    layer4_outputs(211) <= layer3_outputs(3239);
    layer4_outputs(212) <= (layer3_outputs(8826)) xor (layer3_outputs(9611));
    layer4_outputs(213) <= layer3_outputs(5300);
    layer4_outputs(214) <= not((layer3_outputs(1623)) or (layer3_outputs(466)));
    layer4_outputs(215) <= '0';
    layer4_outputs(216) <= not(layer3_outputs(3511));
    layer4_outputs(217) <= (layer3_outputs(6249)) and not (layer3_outputs(6610));
    layer4_outputs(218) <= not(layer3_outputs(2287));
    layer4_outputs(219) <= not(layer3_outputs(2170)) or (layer3_outputs(4681));
    layer4_outputs(220) <= layer3_outputs(725);
    layer4_outputs(221) <= not(layer3_outputs(931)) or (layer3_outputs(1839));
    layer4_outputs(222) <= not(layer3_outputs(865));
    layer4_outputs(223) <= layer3_outputs(86);
    layer4_outputs(224) <= (layer3_outputs(4392)) and not (layer3_outputs(1164));
    layer4_outputs(225) <= not(layer3_outputs(5444));
    layer4_outputs(226) <= not(layer3_outputs(3973));
    layer4_outputs(227) <= layer3_outputs(2570);
    layer4_outputs(228) <= not(layer3_outputs(4500)) or (layer3_outputs(3083));
    layer4_outputs(229) <= not(layer3_outputs(8050));
    layer4_outputs(230) <= not(layer3_outputs(9549));
    layer4_outputs(231) <= (layer3_outputs(3793)) and not (layer3_outputs(6310));
    layer4_outputs(232) <= not(layer3_outputs(7484));
    layer4_outputs(233) <= layer3_outputs(4473);
    layer4_outputs(234) <= not(layer3_outputs(9849));
    layer4_outputs(235) <= (layer3_outputs(6497)) xor (layer3_outputs(5082));
    layer4_outputs(236) <= not(layer3_outputs(2995));
    layer4_outputs(237) <= (layer3_outputs(49)) and (layer3_outputs(7860));
    layer4_outputs(238) <= not(layer3_outputs(9293)) or (layer3_outputs(837));
    layer4_outputs(239) <= not(layer3_outputs(9018));
    layer4_outputs(240) <= layer3_outputs(7424);
    layer4_outputs(241) <= layer3_outputs(4405);
    layer4_outputs(242) <= (layer3_outputs(10225)) and not (layer3_outputs(9081));
    layer4_outputs(243) <= (layer3_outputs(9211)) xor (layer3_outputs(2125));
    layer4_outputs(244) <= not(layer3_outputs(7016));
    layer4_outputs(245) <= not(layer3_outputs(8090));
    layer4_outputs(246) <= layer3_outputs(729);
    layer4_outputs(247) <= not(layer3_outputs(7195));
    layer4_outputs(248) <= not((layer3_outputs(1945)) or (layer3_outputs(9382)));
    layer4_outputs(249) <= (layer3_outputs(8725)) and not (layer3_outputs(4684));
    layer4_outputs(250) <= not(layer3_outputs(8626)) or (layer3_outputs(782));
    layer4_outputs(251) <= not((layer3_outputs(5613)) xor (layer3_outputs(8181)));
    layer4_outputs(252) <= not(layer3_outputs(8241));
    layer4_outputs(253) <= layer3_outputs(1735);
    layer4_outputs(254) <= (layer3_outputs(8337)) and (layer3_outputs(3309));
    layer4_outputs(255) <= not((layer3_outputs(9929)) and (layer3_outputs(6913)));
    layer4_outputs(256) <= not(layer3_outputs(472));
    layer4_outputs(257) <= not(layer3_outputs(7535)) or (layer3_outputs(4849));
    layer4_outputs(258) <= not((layer3_outputs(2828)) and (layer3_outputs(5011)));
    layer4_outputs(259) <= (layer3_outputs(6938)) and (layer3_outputs(7648));
    layer4_outputs(260) <= (layer3_outputs(7882)) xor (layer3_outputs(7900));
    layer4_outputs(261) <= not(layer3_outputs(9617));
    layer4_outputs(262) <= layer3_outputs(6842);
    layer4_outputs(263) <= not(layer3_outputs(2811));
    layer4_outputs(264) <= (layer3_outputs(911)) xor (layer3_outputs(9237));
    layer4_outputs(265) <= layer3_outputs(4762);
    layer4_outputs(266) <= layer3_outputs(3013);
    layer4_outputs(267) <= layer3_outputs(5463);
    layer4_outputs(268) <= not(layer3_outputs(7997));
    layer4_outputs(269) <= not(layer3_outputs(7909)) or (layer3_outputs(4351));
    layer4_outputs(270) <= (layer3_outputs(2415)) and not (layer3_outputs(4783));
    layer4_outputs(271) <= (layer3_outputs(7785)) and (layer3_outputs(10155));
    layer4_outputs(272) <= (layer3_outputs(1197)) and not (layer3_outputs(1286));
    layer4_outputs(273) <= layer3_outputs(6711);
    layer4_outputs(274) <= layer3_outputs(514);
    layer4_outputs(275) <= layer3_outputs(516);
    layer4_outputs(276) <= not(layer3_outputs(1453)) or (layer3_outputs(3954));
    layer4_outputs(277) <= (layer3_outputs(2461)) or (layer3_outputs(8894));
    layer4_outputs(278) <= not((layer3_outputs(9026)) and (layer3_outputs(375)));
    layer4_outputs(279) <= not(layer3_outputs(1671));
    layer4_outputs(280) <= not(layer3_outputs(3283));
    layer4_outputs(281) <= not((layer3_outputs(5248)) or (layer3_outputs(6128)));
    layer4_outputs(282) <= not(layer3_outputs(996)) or (layer3_outputs(2040));
    layer4_outputs(283) <= not(layer3_outputs(1070));
    layer4_outputs(284) <= not(layer3_outputs(3313));
    layer4_outputs(285) <= (layer3_outputs(6669)) and not (layer3_outputs(4840));
    layer4_outputs(286) <= not(layer3_outputs(2005)) or (layer3_outputs(1920));
    layer4_outputs(287) <= layer3_outputs(7854);
    layer4_outputs(288) <= not((layer3_outputs(7715)) and (layer3_outputs(8300)));
    layer4_outputs(289) <= not((layer3_outputs(4218)) and (layer3_outputs(8003)));
    layer4_outputs(290) <= (layer3_outputs(9921)) and (layer3_outputs(3679));
    layer4_outputs(291) <= (layer3_outputs(4775)) and not (layer3_outputs(4158));
    layer4_outputs(292) <= (layer3_outputs(8643)) xor (layer3_outputs(4349));
    layer4_outputs(293) <= layer3_outputs(9698);
    layer4_outputs(294) <= layer3_outputs(6879);
    layer4_outputs(295) <= (layer3_outputs(3163)) xor (layer3_outputs(5908));
    layer4_outputs(296) <= (layer3_outputs(7979)) and not (layer3_outputs(5880));
    layer4_outputs(297) <= (layer3_outputs(3438)) xor (layer3_outputs(9802));
    layer4_outputs(298) <= not(layer3_outputs(7419));
    layer4_outputs(299) <= layer3_outputs(3222);
    layer4_outputs(300) <= not(layer3_outputs(7550));
    layer4_outputs(301) <= not((layer3_outputs(3908)) and (layer3_outputs(1402)));
    layer4_outputs(302) <= layer3_outputs(9692);
    layer4_outputs(303) <= (layer3_outputs(4164)) and not (layer3_outputs(666));
    layer4_outputs(304) <= not(layer3_outputs(5303));
    layer4_outputs(305) <= not((layer3_outputs(5033)) xor (layer3_outputs(134)));
    layer4_outputs(306) <= not(layer3_outputs(1442));
    layer4_outputs(307) <= not((layer3_outputs(9471)) or (layer3_outputs(2273)));
    layer4_outputs(308) <= layer3_outputs(8556);
    layer4_outputs(309) <= layer3_outputs(10142);
    layer4_outputs(310) <= not(layer3_outputs(8296)) or (layer3_outputs(6734));
    layer4_outputs(311) <= layer3_outputs(6401);
    layer4_outputs(312) <= not(layer3_outputs(9870));
    layer4_outputs(313) <= not(layer3_outputs(9621));
    layer4_outputs(314) <= layer3_outputs(9980);
    layer4_outputs(315) <= layer3_outputs(9569);
    layer4_outputs(316) <= not(layer3_outputs(9880));
    layer4_outputs(317) <= not(layer3_outputs(6554)) or (layer3_outputs(10013));
    layer4_outputs(318) <= layer3_outputs(3365);
    layer4_outputs(319) <= (layer3_outputs(4438)) xor (layer3_outputs(1030));
    layer4_outputs(320) <= (layer3_outputs(3699)) and not (layer3_outputs(322));
    layer4_outputs(321) <= (layer3_outputs(5212)) and not (layer3_outputs(4786));
    layer4_outputs(322) <= not(layer3_outputs(4068));
    layer4_outputs(323) <= not(layer3_outputs(8365));
    layer4_outputs(324) <= layer3_outputs(2384);
    layer4_outputs(325) <= not(layer3_outputs(516));
    layer4_outputs(326) <= (layer3_outputs(761)) xor (layer3_outputs(7902));
    layer4_outputs(327) <= not(layer3_outputs(7229)) or (layer3_outputs(2234));
    layer4_outputs(328) <= not((layer3_outputs(7349)) xor (layer3_outputs(8156)));
    layer4_outputs(329) <= not(layer3_outputs(5597));
    layer4_outputs(330) <= layer3_outputs(1832);
    layer4_outputs(331) <= not(layer3_outputs(5562));
    layer4_outputs(332) <= not(layer3_outputs(951));
    layer4_outputs(333) <= not(layer3_outputs(9214)) or (layer3_outputs(4743));
    layer4_outputs(334) <= not(layer3_outputs(3973)) or (layer3_outputs(6513));
    layer4_outputs(335) <= not(layer3_outputs(9933));
    layer4_outputs(336) <= not((layer3_outputs(4006)) and (layer3_outputs(1894)));
    layer4_outputs(337) <= (layer3_outputs(7189)) and not (layer3_outputs(8083));
    layer4_outputs(338) <= not(layer3_outputs(2845)) or (layer3_outputs(7605));
    layer4_outputs(339) <= layer3_outputs(3049);
    layer4_outputs(340) <= not(layer3_outputs(3531));
    layer4_outputs(341) <= layer3_outputs(507);
    layer4_outputs(342) <= not((layer3_outputs(7658)) xor (layer3_outputs(8860)));
    layer4_outputs(343) <= not(layer3_outputs(5142));
    layer4_outputs(344) <= layer3_outputs(6937);
    layer4_outputs(345) <= not(layer3_outputs(600));
    layer4_outputs(346) <= layer3_outputs(8258);
    layer4_outputs(347) <= (layer3_outputs(6297)) and (layer3_outputs(2647));
    layer4_outputs(348) <= not((layer3_outputs(276)) xor (layer3_outputs(502)));
    layer4_outputs(349) <= not(layer3_outputs(259));
    layer4_outputs(350) <= (layer3_outputs(3736)) xor (layer3_outputs(5296));
    layer4_outputs(351) <= (layer3_outputs(2628)) xor (layer3_outputs(5751));
    layer4_outputs(352) <= not((layer3_outputs(1796)) xor (layer3_outputs(4628)));
    layer4_outputs(353) <= (layer3_outputs(9264)) and (layer3_outputs(6432));
    layer4_outputs(354) <= layer3_outputs(8747);
    layer4_outputs(355) <= (layer3_outputs(8602)) and (layer3_outputs(213));
    layer4_outputs(356) <= layer3_outputs(9908);
    layer4_outputs(357) <= layer3_outputs(1645);
    layer4_outputs(358) <= (layer3_outputs(7221)) xor (layer3_outputs(6811));
    layer4_outputs(359) <= not(layer3_outputs(7064));
    layer4_outputs(360) <= not(layer3_outputs(2945));
    layer4_outputs(361) <= layer3_outputs(9222);
    layer4_outputs(362) <= not((layer3_outputs(9927)) xor (layer3_outputs(2267)));
    layer4_outputs(363) <= (layer3_outputs(8195)) and (layer3_outputs(4747));
    layer4_outputs(364) <= layer3_outputs(6003);
    layer4_outputs(365) <= not(layer3_outputs(5023));
    layer4_outputs(366) <= not((layer3_outputs(5653)) xor (layer3_outputs(3920)));
    layer4_outputs(367) <= layer3_outputs(6055);
    layer4_outputs(368) <= (layer3_outputs(3676)) xor (layer3_outputs(6001));
    layer4_outputs(369) <= not(layer3_outputs(7410));
    layer4_outputs(370) <= not(layer3_outputs(1946));
    layer4_outputs(371) <= layer3_outputs(6783);
    layer4_outputs(372) <= not((layer3_outputs(7499)) xor (layer3_outputs(3319)));
    layer4_outputs(373) <= layer3_outputs(3297);
    layer4_outputs(374) <= not(layer3_outputs(3866));
    layer4_outputs(375) <= not((layer3_outputs(9997)) xor (layer3_outputs(8541)));
    layer4_outputs(376) <= not(layer3_outputs(442));
    layer4_outputs(377) <= not(layer3_outputs(9124));
    layer4_outputs(378) <= not((layer3_outputs(1448)) xor (layer3_outputs(2061)));
    layer4_outputs(379) <= not(layer3_outputs(1419));
    layer4_outputs(380) <= not(layer3_outputs(9410));
    layer4_outputs(381) <= layer3_outputs(2242);
    layer4_outputs(382) <= layer3_outputs(7427);
    layer4_outputs(383) <= (layer3_outputs(6422)) or (layer3_outputs(2644));
    layer4_outputs(384) <= layer3_outputs(126);
    layer4_outputs(385) <= (layer3_outputs(9802)) or (layer3_outputs(1643));
    layer4_outputs(386) <= layer3_outputs(1054);
    layer4_outputs(387) <= not(layer3_outputs(6886));
    layer4_outputs(388) <= not((layer3_outputs(8569)) or (layer3_outputs(10192)));
    layer4_outputs(389) <= (layer3_outputs(8500)) and (layer3_outputs(599));
    layer4_outputs(390) <= layer3_outputs(1726);
    layer4_outputs(391) <= layer3_outputs(65);
    layer4_outputs(392) <= layer3_outputs(6306);
    layer4_outputs(393) <= layer3_outputs(5540);
    layer4_outputs(394) <= not(layer3_outputs(3509));
    layer4_outputs(395) <= (layer3_outputs(10053)) xor (layer3_outputs(8970));
    layer4_outputs(396) <= not(layer3_outputs(1524));
    layer4_outputs(397) <= (layer3_outputs(8304)) and not (layer3_outputs(1022));
    layer4_outputs(398) <= layer3_outputs(1372);
    layer4_outputs(399) <= not(layer3_outputs(2139));
    layer4_outputs(400) <= not(layer3_outputs(2721));
    layer4_outputs(401) <= not(layer3_outputs(1092));
    layer4_outputs(402) <= not(layer3_outputs(8843));
    layer4_outputs(403) <= layer3_outputs(5022);
    layer4_outputs(404) <= layer3_outputs(2990);
    layer4_outputs(405) <= layer3_outputs(10016);
    layer4_outputs(406) <= layer3_outputs(8186);
    layer4_outputs(407) <= (layer3_outputs(10024)) and (layer3_outputs(7857));
    layer4_outputs(408) <= layer3_outputs(8867);
    layer4_outputs(409) <= not((layer3_outputs(1699)) xor (layer3_outputs(7051)));
    layer4_outputs(410) <= not(layer3_outputs(7892));
    layer4_outputs(411) <= not((layer3_outputs(870)) and (layer3_outputs(2024)));
    layer4_outputs(412) <= layer3_outputs(7944);
    layer4_outputs(413) <= not((layer3_outputs(5809)) xor (layer3_outputs(589)));
    layer4_outputs(414) <= (layer3_outputs(6832)) xor (layer3_outputs(2113));
    layer4_outputs(415) <= (layer3_outputs(8181)) and (layer3_outputs(512));
    layer4_outputs(416) <= not(layer3_outputs(8895));
    layer4_outputs(417) <= layer3_outputs(467);
    layer4_outputs(418) <= (layer3_outputs(98)) xor (layer3_outputs(4474));
    layer4_outputs(419) <= not(layer3_outputs(2512));
    layer4_outputs(420) <= not(layer3_outputs(115));
    layer4_outputs(421) <= not(layer3_outputs(3613)) or (layer3_outputs(4874));
    layer4_outputs(422) <= not(layer3_outputs(7778));
    layer4_outputs(423) <= not(layer3_outputs(5731)) or (layer3_outputs(4281));
    layer4_outputs(424) <= not(layer3_outputs(934));
    layer4_outputs(425) <= (layer3_outputs(2550)) xor (layer3_outputs(1045));
    layer4_outputs(426) <= not((layer3_outputs(7833)) or (layer3_outputs(3716)));
    layer4_outputs(427) <= (layer3_outputs(4464)) xor (layer3_outputs(10074));
    layer4_outputs(428) <= (layer3_outputs(2379)) and (layer3_outputs(5577));
    layer4_outputs(429) <= not(layer3_outputs(1958));
    layer4_outputs(430) <= not((layer3_outputs(5093)) xor (layer3_outputs(2548)));
    layer4_outputs(431) <= not(layer3_outputs(6544));
    layer4_outputs(432) <= not((layer3_outputs(1724)) xor (layer3_outputs(3481)));
    layer4_outputs(433) <= layer3_outputs(6711);
    layer4_outputs(434) <= not(layer3_outputs(1038));
    layer4_outputs(435) <= not(layer3_outputs(2744)) or (layer3_outputs(8724));
    layer4_outputs(436) <= not((layer3_outputs(7662)) xor (layer3_outputs(5350)));
    layer4_outputs(437) <= (layer3_outputs(8078)) and (layer3_outputs(8588));
    layer4_outputs(438) <= not(layer3_outputs(81));
    layer4_outputs(439) <= not((layer3_outputs(6875)) xor (layer3_outputs(9326)));
    layer4_outputs(440) <= layer3_outputs(10153);
    layer4_outputs(441) <= not(layer3_outputs(2051));
    layer4_outputs(442) <= layer3_outputs(2613);
    layer4_outputs(443) <= not(layer3_outputs(495));
    layer4_outputs(444) <= layer3_outputs(9427);
    layer4_outputs(445) <= not((layer3_outputs(7870)) xor (layer3_outputs(2690)));
    layer4_outputs(446) <= not(layer3_outputs(5831));
    layer4_outputs(447) <= layer3_outputs(9620);
    layer4_outputs(448) <= layer3_outputs(2662);
    layer4_outputs(449) <= '0';
    layer4_outputs(450) <= not(layer3_outputs(7830));
    layer4_outputs(451) <= layer3_outputs(1349);
    layer4_outputs(452) <= (layer3_outputs(4157)) and not (layer3_outputs(6583));
    layer4_outputs(453) <= layer3_outputs(7819);
    layer4_outputs(454) <= not(layer3_outputs(5625)) or (layer3_outputs(4469));
    layer4_outputs(455) <= not(layer3_outputs(9051));
    layer4_outputs(456) <= (layer3_outputs(5130)) and (layer3_outputs(10046));
    layer4_outputs(457) <= not(layer3_outputs(5941)) or (layer3_outputs(6918));
    layer4_outputs(458) <= not((layer3_outputs(9504)) xor (layer3_outputs(4294)));
    layer4_outputs(459) <= layer3_outputs(8940);
    layer4_outputs(460) <= (layer3_outputs(10062)) and not (layer3_outputs(9016));
    layer4_outputs(461) <= (layer3_outputs(5690)) or (layer3_outputs(6270));
    layer4_outputs(462) <= not(layer3_outputs(991));
    layer4_outputs(463) <= not(layer3_outputs(4939));
    layer4_outputs(464) <= layer3_outputs(8691);
    layer4_outputs(465) <= (layer3_outputs(7072)) or (layer3_outputs(6713));
    layer4_outputs(466) <= not((layer3_outputs(4144)) xor (layer3_outputs(2450)));
    layer4_outputs(467) <= not(layer3_outputs(8138));
    layer4_outputs(468) <= (layer3_outputs(238)) and not (layer3_outputs(219));
    layer4_outputs(469) <= not(layer3_outputs(3431));
    layer4_outputs(470) <= not(layer3_outputs(7182));
    layer4_outputs(471) <= layer3_outputs(5551);
    layer4_outputs(472) <= layer3_outputs(4812);
    layer4_outputs(473) <= (layer3_outputs(5639)) and not (layer3_outputs(1720));
    layer4_outputs(474) <= layer3_outputs(6574);
    layer4_outputs(475) <= not(layer3_outputs(3167));
    layer4_outputs(476) <= not(layer3_outputs(8584));
    layer4_outputs(477) <= layer3_outputs(5524);
    layer4_outputs(478) <= layer3_outputs(6855);
    layer4_outputs(479) <= layer3_outputs(8794);
    layer4_outputs(480) <= not((layer3_outputs(7876)) and (layer3_outputs(10068)));
    layer4_outputs(481) <= (layer3_outputs(7096)) and (layer3_outputs(3698));
    layer4_outputs(482) <= (layer3_outputs(8682)) xor (layer3_outputs(9858));
    layer4_outputs(483) <= (layer3_outputs(1875)) and (layer3_outputs(338));
    layer4_outputs(484) <= (layer3_outputs(2518)) xor (layer3_outputs(8456));
    layer4_outputs(485) <= not(layer3_outputs(3268));
    layer4_outputs(486) <= (layer3_outputs(895)) xor (layer3_outputs(874));
    layer4_outputs(487) <= not(layer3_outputs(7147)) or (layer3_outputs(6744));
    layer4_outputs(488) <= not(layer3_outputs(1908));
    layer4_outputs(489) <= not(layer3_outputs(2495)) or (layer3_outputs(6187));
    layer4_outputs(490) <= not(layer3_outputs(4210));
    layer4_outputs(491) <= not(layer3_outputs(6087)) or (layer3_outputs(5207));
    layer4_outputs(492) <= not(layer3_outputs(7100));
    layer4_outputs(493) <= (layer3_outputs(9110)) xor (layer3_outputs(6552));
    layer4_outputs(494) <= not(layer3_outputs(9791));
    layer4_outputs(495) <= not((layer3_outputs(197)) or (layer3_outputs(6486)));
    layer4_outputs(496) <= (layer3_outputs(2533)) xor (layer3_outputs(5547));
    layer4_outputs(497) <= not(layer3_outputs(9687)) or (layer3_outputs(9138));
    layer4_outputs(498) <= not(layer3_outputs(8671));
    layer4_outputs(499) <= not(layer3_outputs(7951));
    layer4_outputs(500) <= not(layer3_outputs(9695));
    layer4_outputs(501) <= (layer3_outputs(5956)) and not (layer3_outputs(359));
    layer4_outputs(502) <= (layer3_outputs(680)) xor (layer3_outputs(6012));
    layer4_outputs(503) <= (layer3_outputs(9446)) xor (layer3_outputs(9473));
    layer4_outputs(504) <= layer3_outputs(9965);
    layer4_outputs(505) <= not(layer3_outputs(5767));
    layer4_outputs(506) <= layer3_outputs(5060);
    layer4_outputs(507) <= (layer3_outputs(8792)) xor (layer3_outputs(9632));
    layer4_outputs(508) <= layer3_outputs(9300);
    layer4_outputs(509) <= '0';
    layer4_outputs(510) <= layer3_outputs(10177);
    layer4_outputs(511) <= (layer3_outputs(2567)) xor (layer3_outputs(7149));
    layer4_outputs(512) <= (layer3_outputs(5251)) xor (layer3_outputs(9497));
    layer4_outputs(513) <= (layer3_outputs(9678)) and (layer3_outputs(3897));
    layer4_outputs(514) <= not((layer3_outputs(6338)) xor (layer3_outputs(8960)));
    layer4_outputs(515) <= layer3_outputs(648);
    layer4_outputs(516) <= layer3_outputs(9987);
    layer4_outputs(517) <= layer3_outputs(3505);
    layer4_outputs(518) <= layer3_outputs(8147);
    layer4_outputs(519) <= layer3_outputs(7272);
    layer4_outputs(520) <= not(layer3_outputs(7008));
    layer4_outputs(521) <= '0';
    layer4_outputs(522) <= layer3_outputs(4324);
    layer4_outputs(523) <= layer3_outputs(2602);
    layer4_outputs(524) <= layer3_outputs(3276);
    layer4_outputs(525) <= layer3_outputs(6092);
    layer4_outputs(526) <= layer3_outputs(6375);
    layer4_outputs(527) <= not(layer3_outputs(3198)) or (layer3_outputs(7504));
    layer4_outputs(528) <= layer3_outputs(7135);
    layer4_outputs(529) <= not(layer3_outputs(9918));
    layer4_outputs(530) <= (layer3_outputs(8529)) and not (layer3_outputs(7416));
    layer4_outputs(531) <= not((layer3_outputs(5725)) or (layer3_outputs(3678)));
    layer4_outputs(532) <= '1';
    layer4_outputs(533) <= layer3_outputs(9996);
    layer4_outputs(534) <= layer3_outputs(3090);
    layer4_outputs(535) <= not(layer3_outputs(9871));
    layer4_outputs(536) <= not((layer3_outputs(5323)) xor (layer3_outputs(2526)));
    layer4_outputs(537) <= layer3_outputs(2250);
    layer4_outputs(538) <= not((layer3_outputs(4193)) and (layer3_outputs(1213)));
    layer4_outputs(539) <= layer3_outputs(1538);
    layer4_outputs(540) <= not(layer3_outputs(3028));
    layer4_outputs(541) <= '0';
    layer4_outputs(542) <= layer3_outputs(1823);
    layer4_outputs(543) <= (layer3_outputs(737)) xor (layer3_outputs(7017));
    layer4_outputs(544) <= not(layer3_outputs(9311));
    layer4_outputs(545) <= not(layer3_outputs(3635)) or (layer3_outputs(582));
    layer4_outputs(546) <= (layer3_outputs(2329)) and not (layer3_outputs(7803));
    layer4_outputs(547) <= not(layer3_outputs(9503));
    layer4_outputs(548) <= layer3_outputs(9396);
    layer4_outputs(549) <= not(layer3_outputs(8339));
    layer4_outputs(550) <= not(layer3_outputs(2904)) or (layer3_outputs(8788));
    layer4_outputs(551) <= (layer3_outputs(1721)) xor (layer3_outputs(8655));
    layer4_outputs(552) <= not(layer3_outputs(5173));
    layer4_outputs(553) <= layer3_outputs(1984);
    layer4_outputs(554) <= not(layer3_outputs(3972));
    layer4_outputs(555) <= not(layer3_outputs(4365)) or (layer3_outputs(7797));
    layer4_outputs(556) <= (layer3_outputs(739)) and (layer3_outputs(7147));
    layer4_outputs(557) <= not(layer3_outputs(5721)) or (layer3_outputs(7312));
    layer4_outputs(558) <= layer3_outputs(2634);
    layer4_outputs(559) <= layer3_outputs(7796);
    layer4_outputs(560) <= (layer3_outputs(6506)) xor (layer3_outputs(771));
    layer4_outputs(561) <= not(layer3_outputs(2422)) or (layer3_outputs(727));
    layer4_outputs(562) <= not((layer3_outputs(7767)) xor (layer3_outputs(2918)));
    layer4_outputs(563) <= (layer3_outputs(631)) and not (layer3_outputs(1970));
    layer4_outputs(564) <= layer3_outputs(2518);
    layer4_outputs(565) <= (layer3_outputs(5148)) xor (layer3_outputs(2993));
    layer4_outputs(566) <= not(layer3_outputs(1310)) or (layer3_outputs(7453));
    layer4_outputs(567) <= not(layer3_outputs(7827));
    layer4_outputs(568) <= not(layer3_outputs(2964)) or (layer3_outputs(5790));
    layer4_outputs(569) <= layer3_outputs(9071);
    layer4_outputs(570) <= not(layer3_outputs(6953)) or (layer3_outputs(8459));
    layer4_outputs(571) <= not(layer3_outputs(4582));
    layer4_outputs(572) <= not(layer3_outputs(7137));
    layer4_outputs(573) <= not((layer3_outputs(5472)) xor (layer3_outputs(375)));
    layer4_outputs(574) <= not(layer3_outputs(8976));
    layer4_outputs(575) <= (layer3_outputs(4044)) xor (layer3_outputs(8773));
    layer4_outputs(576) <= not(layer3_outputs(7573));
    layer4_outputs(577) <= not(layer3_outputs(9095)) or (layer3_outputs(8292));
    layer4_outputs(578) <= not(layer3_outputs(6799));
    layer4_outputs(579) <= not(layer3_outputs(4259)) or (layer3_outputs(6856));
    layer4_outputs(580) <= not((layer3_outputs(5272)) or (layer3_outputs(3970)));
    layer4_outputs(581) <= not(layer3_outputs(1281)) or (layer3_outputs(2052));
    layer4_outputs(582) <= not((layer3_outputs(7653)) xor (layer3_outputs(4171)));
    layer4_outputs(583) <= not(layer3_outputs(3289));
    layer4_outputs(584) <= layer3_outputs(5668);
    layer4_outputs(585) <= (layer3_outputs(9645)) and not (layer3_outputs(81));
    layer4_outputs(586) <= not(layer3_outputs(1425)) or (layer3_outputs(6540));
    layer4_outputs(587) <= not((layer3_outputs(368)) or (layer3_outputs(3759)));
    layer4_outputs(588) <= not(layer3_outputs(8498));
    layer4_outputs(589) <= not(layer3_outputs(668));
    layer4_outputs(590) <= layer3_outputs(4897);
    layer4_outputs(591) <= not(layer3_outputs(449));
    layer4_outputs(592) <= not((layer3_outputs(8366)) or (layer3_outputs(6422)));
    layer4_outputs(593) <= not(layer3_outputs(2326));
    layer4_outputs(594) <= not(layer3_outputs(6613));
    layer4_outputs(595) <= layer3_outputs(3002);
    layer4_outputs(596) <= (layer3_outputs(6006)) xor (layer3_outputs(5933));
    layer4_outputs(597) <= not(layer3_outputs(1076));
    layer4_outputs(598) <= (layer3_outputs(1348)) and not (layer3_outputs(9079));
    layer4_outputs(599) <= (layer3_outputs(3232)) and (layer3_outputs(8266));
    layer4_outputs(600) <= layer3_outputs(5331);
    layer4_outputs(601) <= layer3_outputs(802);
    layer4_outputs(602) <= layer3_outputs(5329);
    layer4_outputs(603) <= (layer3_outputs(3669)) xor (layer3_outputs(3417));
    layer4_outputs(604) <= not((layer3_outputs(6988)) xor (layer3_outputs(8587)));
    layer4_outputs(605) <= layer3_outputs(7782);
    layer4_outputs(606) <= layer3_outputs(6751);
    layer4_outputs(607) <= (layer3_outputs(2586)) or (layer3_outputs(5797));
    layer4_outputs(608) <= not(layer3_outputs(9474));
    layer4_outputs(609) <= not(layer3_outputs(2751));
    layer4_outputs(610) <= layer3_outputs(3033);
    layer4_outputs(611) <= not(layer3_outputs(6715)) or (layer3_outputs(9396));
    layer4_outputs(612) <= not((layer3_outputs(8604)) xor (layer3_outputs(1392)));
    layer4_outputs(613) <= (layer3_outputs(5471)) xor (layer3_outputs(8508));
    layer4_outputs(614) <= not((layer3_outputs(6556)) or (layer3_outputs(2974)));
    layer4_outputs(615) <= not((layer3_outputs(1987)) and (layer3_outputs(185)));
    layer4_outputs(616) <= not(layer3_outputs(699));
    layer4_outputs(617) <= not((layer3_outputs(7885)) xor (layer3_outputs(2675)));
    layer4_outputs(618) <= not(layer3_outputs(8151));
    layer4_outputs(619) <= not(layer3_outputs(4330));
    layer4_outputs(620) <= (layer3_outputs(10154)) and not (layer3_outputs(6503));
    layer4_outputs(621) <= not((layer3_outputs(7891)) xor (layer3_outputs(2013)));
    layer4_outputs(622) <= (layer3_outputs(8209)) xor (layer3_outputs(3088));
    layer4_outputs(623) <= not(layer3_outputs(3922));
    layer4_outputs(624) <= (layer3_outputs(8782)) or (layer3_outputs(2612));
    layer4_outputs(625) <= '0';
    layer4_outputs(626) <= not(layer3_outputs(2447));
    layer4_outputs(627) <= not((layer3_outputs(1595)) and (layer3_outputs(970)));
    layer4_outputs(628) <= not(layer3_outputs(9971));
    layer4_outputs(629) <= (layer3_outputs(4353)) xor (layer3_outputs(9657));
    layer4_outputs(630) <= (layer3_outputs(1470)) and (layer3_outputs(474));
    layer4_outputs(631) <= not((layer3_outputs(2086)) xor (layer3_outputs(1464)));
    layer4_outputs(632) <= (layer3_outputs(1617)) and not (layer3_outputs(1085));
    layer4_outputs(633) <= not((layer3_outputs(687)) or (layer3_outputs(7576)));
    layer4_outputs(634) <= not(layer3_outputs(4755)) or (layer3_outputs(1354));
    layer4_outputs(635) <= layer3_outputs(2412);
    layer4_outputs(636) <= (layer3_outputs(966)) or (layer3_outputs(4533));
    layer4_outputs(637) <= (layer3_outputs(431)) xor (layer3_outputs(957));
    layer4_outputs(638) <= layer3_outputs(2838);
    layer4_outputs(639) <= not((layer3_outputs(5546)) xor (layer3_outputs(3585)));
    layer4_outputs(640) <= not(layer3_outputs(6416)) or (layer3_outputs(180));
    layer4_outputs(641) <= not(layer3_outputs(6929));
    layer4_outputs(642) <= not(layer3_outputs(1188));
    layer4_outputs(643) <= not(layer3_outputs(4844));
    layer4_outputs(644) <= layer3_outputs(330);
    layer4_outputs(645) <= not(layer3_outputs(8965));
    layer4_outputs(646) <= (layer3_outputs(5113)) xor (layer3_outputs(5791));
    layer4_outputs(647) <= not(layer3_outputs(9987));
    layer4_outputs(648) <= not(layer3_outputs(2704));
    layer4_outputs(649) <= layer3_outputs(5380);
    layer4_outputs(650) <= (layer3_outputs(838)) xor (layer3_outputs(3514));
    layer4_outputs(651) <= not(layer3_outputs(6370));
    layer4_outputs(652) <= layer3_outputs(749);
    layer4_outputs(653) <= (layer3_outputs(7554)) or (layer3_outputs(5812));
    layer4_outputs(654) <= (layer3_outputs(7308)) and not (layer3_outputs(9827));
    layer4_outputs(655) <= not((layer3_outputs(9720)) xor (layer3_outputs(7964)));
    layer4_outputs(656) <= not(layer3_outputs(9230)) or (layer3_outputs(782));
    layer4_outputs(657) <= layer3_outputs(8764);
    layer4_outputs(658) <= layer3_outputs(5256);
    layer4_outputs(659) <= not(layer3_outputs(8447));
    layer4_outputs(660) <= not(layer3_outputs(7210)) or (layer3_outputs(6532));
    layer4_outputs(661) <= layer3_outputs(4567);
    layer4_outputs(662) <= not(layer3_outputs(4716));
    layer4_outputs(663) <= layer3_outputs(4926);
    layer4_outputs(664) <= layer3_outputs(1427);
    layer4_outputs(665) <= (layer3_outputs(5076)) and not (layer3_outputs(3831));
    layer4_outputs(666) <= not((layer3_outputs(7043)) xor (layer3_outputs(7094)));
    layer4_outputs(667) <= not((layer3_outputs(184)) xor (layer3_outputs(2252)));
    layer4_outputs(668) <= (layer3_outputs(4712)) and (layer3_outputs(8932));
    layer4_outputs(669) <= (layer3_outputs(1280)) and not (layer3_outputs(4534));
    layer4_outputs(670) <= not((layer3_outputs(6846)) xor (layer3_outputs(10227)));
    layer4_outputs(671) <= not(layer3_outputs(6404)) or (layer3_outputs(8283));
    layer4_outputs(672) <= layer3_outputs(5478);
    layer4_outputs(673) <= not((layer3_outputs(7930)) xor (layer3_outputs(4841)));
    layer4_outputs(674) <= not(layer3_outputs(4813));
    layer4_outputs(675) <= not((layer3_outputs(3367)) xor (layer3_outputs(6610)));
    layer4_outputs(676) <= not(layer3_outputs(6391)) or (layer3_outputs(9619));
    layer4_outputs(677) <= layer3_outputs(4880);
    layer4_outputs(678) <= not(layer3_outputs(2897));
    layer4_outputs(679) <= not(layer3_outputs(8431));
    layer4_outputs(680) <= not(layer3_outputs(9754));
    layer4_outputs(681) <= layer3_outputs(3259);
    layer4_outputs(682) <= not(layer3_outputs(1102)) or (layer3_outputs(2896));
    layer4_outputs(683) <= not((layer3_outputs(9438)) and (layer3_outputs(1282)));
    layer4_outputs(684) <= not((layer3_outputs(137)) xor (layer3_outputs(7650)));
    layer4_outputs(685) <= not((layer3_outputs(6211)) or (layer3_outputs(7823)));
    layer4_outputs(686) <= (layer3_outputs(6399)) or (layer3_outputs(6076));
    layer4_outputs(687) <= not(layer3_outputs(3603));
    layer4_outputs(688) <= layer3_outputs(7289);
    layer4_outputs(689) <= not(layer3_outputs(7892));
    layer4_outputs(690) <= not(layer3_outputs(932));
    layer4_outputs(691) <= not(layer3_outputs(3041));
    layer4_outputs(692) <= not(layer3_outputs(3931));
    layer4_outputs(693) <= not(layer3_outputs(4924));
    layer4_outputs(694) <= (layer3_outputs(2212)) and (layer3_outputs(6496));
    layer4_outputs(695) <= layer3_outputs(3015);
    layer4_outputs(696) <= not((layer3_outputs(5611)) and (layer3_outputs(5157)));
    layer4_outputs(697) <= not((layer3_outputs(5669)) and (layer3_outputs(503)));
    layer4_outputs(698) <= not((layer3_outputs(6696)) and (layer3_outputs(8542)));
    layer4_outputs(699) <= (layer3_outputs(10036)) and not (layer3_outputs(6407));
    layer4_outputs(700) <= layer3_outputs(3704);
    layer4_outputs(701) <= not((layer3_outputs(2765)) and (layer3_outputs(4121)));
    layer4_outputs(702) <= (layer3_outputs(4896)) and (layer3_outputs(1951));
    layer4_outputs(703) <= layer3_outputs(4295);
    layer4_outputs(704) <= not(layer3_outputs(315));
    layer4_outputs(705) <= not((layer3_outputs(7209)) xor (layer3_outputs(3323)));
    layer4_outputs(706) <= not((layer3_outputs(1513)) xor (layer3_outputs(4482)));
    layer4_outputs(707) <= not((layer3_outputs(3690)) or (layer3_outputs(4231)));
    layer4_outputs(708) <= not(layer3_outputs(8118));
    layer4_outputs(709) <= layer3_outputs(6884);
    layer4_outputs(710) <= layer3_outputs(8223);
    layer4_outputs(711) <= not(layer3_outputs(1488));
    layer4_outputs(712) <= not(layer3_outputs(4644));
    layer4_outputs(713) <= not(layer3_outputs(4443));
    layer4_outputs(714) <= not(layer3_outputs(5133));
    layer4_outputs(715) <= (layer3_outputs(2574)) and (layer3_outputs(9045));
    layer4_outputs(716) <= not((layer3_outputs(3828)) xor (layer3_outputs(4832)));
    layer4_outputs(717) <= not((layer3_outputs(6148)) xor (layer3_outputs(3741)));
    layer4_outputs(718) <= layer3_outputs(6794);
    layer4_outputs(719) <= not(layer3_outputs(3133));
    layer4_outputs(720) <= (layer3_outputs(8255)) and not (layer3_outputs(9984));
    layer4_outputs(721) <= layer3_outputs(3515);
    layer4_outputs(722) <= layer3_outputs(8814);
    layer4_outputs(723) <= layer3_outputs(9537);
    layer4_outputs(724) <= (layer3_outputs(4479)) and (layer3_outputs(3684));
    layer4_outputs(725) <= not((layer3_outputs(9126)) or (layer3_outputs(1584)));
    layer4_outputs(726) <= layer3_outputs(1559);
    layer4_outputs(727) <= not(layer3_outputs(8449)) or (layer3_outputs(3517));
    layer4_outputs(728) <= not((layer3_outputs(7725)) and (layer3_outputs(7343)));
    layer4_outputs(729) <= not(layer3_outputs(1634));
    layer4_outputs(730) <= (layer3_outputs(9903)) or (layer3_outputs(1121));
    layer4_outputs(731) <= not((layer3_outputs(948)) and (layer3_outputs(4126)));
    layer4_outputs(732) <= not(layer3_outputs(8507)) or (layer3_outputs(6223));
    layer4_outputs(733) <= not((layer3_outputs(6405)) xor (layer3_outputs(4834)));
    layer4_outputs(734) <= not(layer3_outputs(5034));
    layer4_outputs(735) <= not(layer3_outputs(1185));
    layer4_outputs(736) <= layer3_outputs(563);
    layer4_outputs(737) <= not((layer3_outputs(344)) xor (layer3_outputs(2271)));
    layer4_outputs(738) <= not(layer3_outputs(1676));
    layer4_outputs(739) <= not((layer3_outputs(943)) xor (layer3_outputs(4901)));
    layer4_outputs(740) <= (layer3_outputs(9931)) and not (layer3_outputs(5424));
    layer4_outputs(741) <= not(layer3_outputs(1977));
    layer4_outputs(742) <= not(layer3_outputs(3361));
    layer4_outputs(743) <= not(layer3_outputs(1369));
    layer4_outputs(744) <= (layer3_outputs(2379)) and (layer3_outputs(305));
    layer4_outputs(745) <= not(layer3_outputs(6111));
    layer4_outputs(746) <= not(layer3_outputs(6932)) or (layer3_outputs(2108));
    layer4_outputs(747) <= layer3_outputs(2418);
    layer4_outputs(748) <= not(layer3_outputs(1910));
    layer4_outputs(749) <= not(layer3_outputs(3530));
    layer4_outputs(750) <= '1';
    layer4_outputs(751) <= (layer3_outputs(1711)) or (layer3_outputs(839));
    layer4_outputs(752) <= layer3_outputs(7407);
    layer4_outputs(753) <= (layer3_outputs(8576)) and (layer3_outputs(7738));
    layer4_outputs(754) <= layer3_outputs(8068);
    layer4_outputs(755) <= (layer3_outputs(891)) and not (layer3_outputs(8882));
    layer4_outputs(756) <= layer3_outputs(2838);
    layer4_outputs(757) <= layer3_outputs(264);
    layer4_outputs(758) <= not(layer3_outputs(3257));
    layer4_outputs(759) <= not(layer3_outputs(8383)) or (layer3_outputs(6499));
    layer4_outputs(760) <= not((layer3_outputs(4341)) and (layer3_outputs(8268)));
    layer4_outputs(761) <= layer3_outputs(952);
    layer4_outputs(762) <= (layer3_outputs(8093)) and not (layer3_outputs(10214));
    layer4_outputs(763) <= (layer3_outputs(410)) or (layer3_outputs(7855));
    layer4_outputs(764) <= layer3_outputs(930);
    layer4_outputs(765) <= (layer3_outputs(6930)) xor (layer3_outputs(3513));
    layer4_outputs(766) <= (layer3_outputs(6580)) xor (layer3_outputs(4996));
    layer4_outputs(767) <= not((layer3_outputs(7686)) xor (layer3_outputs(9805)));
    layer4_outputs(768) <= not(layer3_outputs(10177));
    layer4_outputs(769) <= not(layer3_outputs(6733));
    layer4_outputs(770) <= layer3_outputs(1498);
    layer4_outputs(771) <= (layer3_outputs(347)) and not (layer3_outputs(3646));
    layer4_outputs(772) <= layer3_outputs(5168);
    layer4_outputs(773) <= layer3_outputs(3488);
    layer4_outputs(774) <= layer3_outputs(7825);
    layer4_outputs(775) <= layer3_outputs(7481);
    layer4_outputs(776) <= not(layer3_outputs(9209));
    layer4_outputs(777) <= not(layer3_outputs(2843));
    layer4_outputs(778) <= not((layer3_outputs(3758)) and (layer3_outputs(7785)));
    layer4_outputs(779) <= layer3_outputs(4144);
    layer4_outputs(780) <= layer3_outputs(7477);
    layer4_outputs(781) <= (layer3_outputs(3138)) xor (layer3_outputs(4180));
    layer4_outputs(782) <= (layer3_outputs(6891)) xor (layer3_outputs(9521));
    layer4_outputs(783) <= (layer3_outputs(1603)) and (layer3_outputs(7120));
    layer4_outputs(784) <= '0';
    layer4_outputs(785) <= not(layer3_outputs(3024));
    layer4_outputs(786) <= (layer3_outputs(7311)) xor (layer3_outputs(2157));
    layer4_outputs(787) <= layer3_outputs(504);
    layer4_outputs(788) <= not(layer3_outputs(2041));
    layer4_outputs(789) <= not((layer3_outputs(2689)) and (layer3_outputs(5599)));
    layer4_outputs(790) <= (layer3_outputs(1954)) xor (layer3_outputs(8108));
    layer4_outputs(791) <= not(layer3_outputs(3224)) or (layer3_outputs(5802));
    layer4_outputs(792) <= layer3_outputs(6163);
    layer4_outputs(793) <= '0';
    layer4_outputs(794) <= (layer3_outputs(5321)) and not (layer3_outputs(4941));
    layer4_outputs(795) <= not((layer3_outputs(6768)) xor (layer3_outputs(6465)));
    layer4_outputs(796) <= not((layer3_outputs(1167)) and (layer3_outputs(7684)));
    layer4_outputs(797) <= not((layer3_outputs(1648)) xor (layer3_outputs(14)));
    layer4_outputs(798) <= layer3_outputs(7036);
    layer4_outputs(799) <= (layer3_outputs(6028)) xor (layer3_outputs(8014));
    layer4_outputs(800) <= not(layer3_outputs(2711));
    layer4_outputs(801) <= not((layer3_outputs(6822)) xor (layer3_outputs(9672)));
    layer4_outputs(802) <= not(layer3_outputs(8760)) or (layer3_outputs(4170));
    layer4_outputs(803) <= not(layer3_outputs(10225));
    layer4_outputs(804) <= not(layer3_outputs(7067));
    layer4_outputs(805) <= not((layer3_outputs(796)) xor (layer3_outputs(8748)));
    layer4_outputs(806) <= not((layer3_outputs(2350)) and (layer3_outputs(1731)));
    layer4_outputs(807) <= not((layer3_outputs(3103)) xor (layer3_outputs(1049)));
    layer4_outputs(808) <= not(layer3_outputs(1533)) or (layer3_outputs(668));
    layer4_outputs(809) <= not(layer3_outputs(10073));
    layer4_outputs(810) <= layer3_outputs(2369);
    layer4_outputs(811) <= layer3_outputs(69);
    layer4_outputs(812) <= not(layer3_outputs(3103));
    layer4_outputs(813) <= layer3_outputs(8392);
    layer4_outputs(814) <= not(layer3_outputs(4027));
    layer4_outputs(815) <= layer3_outputs(8175);
    layer4_outputs(816) <= not(layer3_outputs(5165));
    layer4_outputs(817) <= (layer3_outputs(4640)) and (layer3_outputs(9913));
    layer4_outputs(818) <= layer3_outputs(5031);
    layer4_outputs(819) <= not(layer3_outputs(5799));
    layer4_outputs(820) <= not(layer3_outputs(8728)) or (layer3_outputs(7207));
    layer4_outputs(821) <= not((layer3_outputs(3564)) xor (layer3_outputs(7976)));
    layer4_outputs(822) <= not(layer3_outputs(9313));
    layer4_outputs(823) <= (layer3_outputs(705)) and not (layer3_outputs(4526));
    layer4_outputs(824) <= layer3_outputs(2036);
    layer4_outputs(825) <= '1';
    layer4_outputs(826) <= (layer3_outputs(4096)) and (layer3_outputs(5664));
    layer4_outputs(827) <= not(layer3_outputs(8524));
    layer4_outputs(828) <= not(layer3_outputs(9922));
    layer4_outputs(829) <= layer3_outputs(6623);
    layer4_outputs(830) <= not((layer3_outputs(318)) xor (layer3_outputs(10186)));
    layer4_outputs(831) <= (layer3_outputs(3376)) or (layer3_outputs(6623));
    layer4_outputs(832) <= (layer3_outputs(2256)) xor (layer3_outputs(6811));
    layer4_outputs(833) <= not(layer3_outputs(7810));
    layer4_outputs(834) <= not(layer3_outputs(8352)) or (layer3_outputs(8801));
    layer4_outputs(835) <= not((layer3_outputs(7236)) and (layer3_outputs(8511)));
    layer4_outputs(836) <= not((layer3_outputs(9828)) and (layer3_outputs(9139)));
    layer4_outputs(837) <= not(layer3_outputs(4161)) or (layer3_outputs(2119));
    layer4_outputs(838) <= not((layer3_outputs(7237)) xor (layer3_outputs(2429)));
    layer4_outputs(839) <= (layer3_outputs(3379)) and not (layer3_outputs(3833));
    layer4_outputs(840) <= not((layer3_outputs(929)) or (layer3_outputs(1755)));
    layer4_outputs(841) <= not(layer3_outputs(170));
    layer4_outputs(842) <= not(layer3_outputs(1842)) or (layer3_outputs(2561));
    layer4_outputs(843) <= (layer3_outputs(9707)) and (layer3_outputs(334));
    layer4_outputs(844) <= not(layer3_outputs(5396));
    layer4_outputs(845) <= (layer3_outputs(5833)) and not (layer3_outputs(6553));
    layer4_outputs(846) <= not(layer3_outputs(3821));
    layer4_outputs(847) <= not(layer3_outputs(8585));
    layer4_outputs(848) <= not(layer3_outputs(9559)) or (layer3_outputs(6502));
    layer4_outputs(849) <= layer3_outputs(7042);
    layer4_outputs(850) <= not(layer3_outputs(5246));
    layer4_outputs(851) <= not(layer3_outputs(7810));
    layer4_outputs(852) <= layer3_outputs(4438);
    layer4_outputs(853) <= not(layer3_outputs(2668));
    layer4_outputs(854) <= (layer3_outputs(2496)) and not (layer3_outputs(10));
    layer4_outputs(855) <= not((layer3_outputs(8913)) xor (layer3_outputs(5646)));
    layer4_outputs(856) <= layer3_outputs(5801);
    layer4_outputs(857) <= not(layer3_outputs(2428));
    layer4_outputs(858) <= (layer3_outputs(9766)) and not (layer3_outputs(8484));
    layer4_outputs(859) <= layer3_outputs(4015);
    layer4_outputs(860) <= not((layer3_outputs(5181)) xor (layer3_outputs(5224)));
    layer4_outputs(861) <= layer3_outputs(5539);
    layer4_outputs(862) <= (layer3_outputs(9279)) and (layer3_outputs(8479));
    layer4_outputs(863) <= layer3_outputs(1555);
    layer4_outputs(864) <= layer3_outputs(9998);
    layer4_outputs(865) <= layer3_outputs(10077);
    layer4_outputs(866) <= not((layer3_outputs(349)) xor (layer3_outputs(7624)));
    layer4_outputs(867) <= not(layer3_outputs(7669));
    layer4_outputs(868) <= layer3_outputs(4997);
    layer4_outputs(869) <= (layer3_outputs(5518)) xor (layer3_outputs(4159));
    layer4_outputs(870) <= '1';
    layer4_outputs(871) <= not(layer3_outputs(7795));
    layer4_outputs(872) <= layer3_outputs(541);
    layer4_outputs(873) <= layer3_outputs(9923);
    layer4_outputs(874) <= (layer3_outputs(2601)) and not (layer3_outputs(3912));
    layer4_outputs(875) <= not(layer3_outputs(10105));
    layer4_outputs(876) <= (layer3_outputs(9970)) and (layer3_outputs(6244));
    layer4_outputs(877) <= not(layer3_outputs(7865));
    layer4_outputs(878) <= layer3_outputs(4396);
    layer4_outputs(879) <= not((layer3_outputs(6522)) xor (layer3_outputs(1293)));
    layer4_outputs(880) <= layer3_outputs(6349);
    layer4_outputs(881) <= not(layer3_outputs(8064));
    layer4_outputs(882) <= layer3_outputs(10151);
    layer4_outputs(883) <= not(layer3_outputs(9428));
    layer4_outputs(884) <= layer3_outputs(10159);
    layer4_outputs(885) <= not(layer3_outputs(6680));
    layer4_outputs(886) <= not(layer3_outputs(7035));
    layer4_outputs(887) <= (layer3_outputs(2524)) xor (layer3_outputs(8387));
    layer4_outputs(888) <= not(layer3_outputs(5438)) or (layer3_outputs(5096));
    layer4_outputs(889) <= not(layer3_outputs(10040));
    layer4_outputs(890) <= not(layer3_outputs(7310));
    layer4_outputs(891) <= not(layer3_outputs(7980));
    layer4_outputs(892) <= layer3_outputs(8739);
    layer4_outputs(893) <= '1';
    layer4_outputs(894) <= not(layer3_outputs(1660)) or (layer3_outputs(6299));
    layer4_outputs(895) <= not(layer3_outputs(7251));
    layer4_outputs(896) <= not(layer3_outputs(4567));
    layer4_outputs(897) <= not(layer3_outputs(5247));
    layer4_outputs(898) <= not((layer3_outputs(7260)) and (layer3_outputs(240)));
    layer4_outputs(899) <= not((layer3_outputs(3303)) or (layer3_outputs(1895)));
    layer4_outputs(900) <= not((layer3_outputs(7525)) xor (layer3_outputs(6871)));
    layer4_outputs(901) <= (layer3_outputs(2805)) and (layer3_outputs(1965));
    layer4_outputs(902) <= not(layer3_outputs(8500));
    layer4_outputs(903) <= not(layer3_outputs(2244));
    layer4_outputs(904) <= not(layer3_outputs(6057));
    layer4_outputs(905) <= not((layer3_outputs(1265)) xor (layer3_outputs(5263)));
    layer4_outputs(906) <= not(layer3_outputs(3508));
    layer4_outputs(907) <= not((layer3_outputs(1874)) xor (layer3_outputs(2902)));
    layer4_outputs(908) <= not(layer3_outputs(1156)) or (layer3_outputs(2042));
    layer4_outputs(909) <= not(layer3_outputs(4094)) or (layer3_outputs(8629));
    layer4_outputs(910) <= not(layer3_outputs(8513));
    layer4_outputs(911) <= (layer3_outputs(1144)) xor (layer3_outputs(5109));
    layer4_outputs(912) <= (layer3_outputs(1475)) xor (layer3_outputs(8767));
    layer4_outputs(913) <= not((layer3_outputs(8011)) or (layer3_outputs(1330)));
    layer4_outputs(914) <= not(layer3_outputs(1949)) or (layer3_outputs(1162));
    layer4_outputs(915) <= not(layer3_outputs(8397));
    layer4_outputs(916) <= layer3_outputs(7596);
    layer4_outputs(917) <= not(layer3_outputs(2455));
    layer4_outputs(918) <= (layer3_outputs(7524)) or (layer3_outputs(86));
    layer4_outputs(919) <= layer3_outputs(4620);
    layer4_outputs(920) <= (layer3_outputs(4424)) or (layer3_outputs(9635));
    layer4_outputs(921) <= not((layer3_outputs(8164)) or (layer3_outputs(3930)));
    layer4_outputs(922) <= not(layer3_outputs(6393)) or (layer3_outputs(4225));
    layer4_outputs(923) <= layer3_outputs(1318);
    layer4_outputs(924) <= layer3_outputs(9475);
    layer4_outputs(925) <= not(layer3_outputs(9368));
    layer4_outputs(926) <= not(layer3_outputs(4033)) or (layer3_outputs(9208));
    layer4_outputs(927) <= not(layer3_outputs(552));
    layer4_outputs(928) <= not(layer3_outputs(8273));
    layer4_outputs(929) <= layer3_outputs(7485);
    layer4_outputs(930) <= not((layer3_outputs(2867)) xor (layer3_outputs(5909)));
    layer4_outputs(931) <= (layer3_outputs(10231)) and not (layer3_outputs(2940));
    layer4_outputs(932) <= not(layer3_outputs(8807));
    layer4_outputs(933) <= (layer3_outputs(788)) or (layer3_outputs(9163));
    layer4_outputs(934) <= layer3_outputs(501);
    layer4_outputs(935) <= layer3_outputs(3528);
    layer4_outputs(936) <= layer3_outputs(2943);
    layer4_outputs(937) <= layer3_outputs(4187);
    layer4_outputs(938) <= not(layer3_outputs(982));
    layer4_outputs(939) <= (layer3_outputs(9457)) and (layer3_outputs(8893));
    layer4_outputs(940) <= not((layer3_outputs(4986)) xor (layer3_outputs(6653)));
    layer4_outputs(941) <= (layer3_outputs(8911)) and (layer3_outputs(7312));
    layer4_outputs(942) <= not(layer3_outputs(2920));
    layer4_outputs(943) <= (layer3_outputs(7537)) and not (layer3_outputs(5809));
    layer4_outputs(944) <= layer3_outputs(5560);
    layer4_outputs(945) <= not(layer3_outputs(7403));
    layer4_outputs(946) <= (layer3_outputs(6856)) xor (layer3_outputs(994));
    layer4_outputs(947) <= (layer3_outputs(9985)) and not (layer3_outputs(4705));
    layer4_outputs(948) <= layer3_outputs(9167);
    layer4_outputs(949) <= not(layer3_outputs(5344));
    layer4_outputs(950) <= layer3_outputs(3658);
    layer4_outputs(951) <= (layer3_outputs(6285)) xor (layer3_outputs(8772));
    layer4_outputs(952) <= not(layer3_outputs(6636));
    layer4_outputs(953) <= not(layer3_outputs(5854));
    layer4_outputs(954) <= '0';
    layer4_outputs(955) <= not(layer3_outputs(8350));
    layer4_outputs(956) <= (layer3_outputs(1125)) xor (layer3_outputs(6830));
    layer4_outputs(957) <= not(layer3_outputs(8066));
    layer4_outputs(958) <= not((layer3_outputs(5653)) xor (layer3_outputs(5067)));
    layer4_outputs(959) <= not(layer3_outputs(3057)) or (layer3_outputs(6752));
    layer4_outputs(960) <= (layer3_outputs(3360)) and not (layer3_outputs(2911));
    layer4_outputs(961) <= layer3_outputs(2378);
    layer4_outputs(962) <= not((layer3_outputs(50)) and (layer3_outputs(3425)));
    layer4_outputs(963) <= layer3_outputs(1925);
    layer4_outputs(964) <= not((layer3_outputs(5563)) xor (layer3_outputs(4295)));
    layer4_outputs(965) <= (layer3_outputs(8931)) and not (layer3_outputs(3021));
    layer4_outputs(966) <= (layer3_outputs(3745)) and (layer3_outputs(4748));
    layer4_outputs(967) <= (layer3_outputs(10145)) and (layer3_outputs(1701));
    layer4_outputs(968) <= not(layer3_outputs(6760));
    layer4_outputs(969) <= (layer3_outputs(3402)) and not (layer3_outputs(6439));
    layer4_outputs(970) <= not(layer3_outputs(627));
    layer4_outputs(971) <= layer3_outputs(4646);
    layer4_outputs(972) <= not(layer3_outputs(168));
    layer4_outputs(973) <= not(layer3_outputs(7352));
    layer4_outputs(974) <= layer3_outputs(1590);
    layer4_outputs(975) <= not(layer3_outputs(7494));
    layer4_outputs(976) <= (layer3_outputs(9851)) xor (layer3_outputs(1606));
    layer4_outputs(977) <= not((layer3_outputs(2810)) or (layer3_outputs(3959)));
    layer4_outputs(978) <= not((layer3_outputs(6655)) and (layer3_outputs(2459)));
    layer4_outputs(979) <= not((layer3_outputs(5106)) xor (layer3_outputs(3454)));
    layer4_outputs(980) <= not(layer3_outputs(9968));
    layer4_outputs(981) <= not(layer3_outputs(6100));
    layer4_outputs(982) <= (layer3_outputs(8703)) and (layer3_outputs(5020));
    layer4_outputs(983) <= layer3_outputs(1652);
    layer4_outputs(984) <= (layer3_outputs(1655)) or (layer3_outputs(8424));
    layer4_outputs(985) <= layer3_outputs(1924);
    layer4_outputs(986) <= not(layer3_outputs(5218)) or (layer3_outputs(2685));
    layer4_outputs(987) <= not(layer3_outputs(3622));
    layer4_outputs(988) <= not(layer3_outputs(236));
    layer4_outputs(989) <= not((layer3_outputs(1166)) or (layer3_outputs(4155)));
    layer4_outputs(990) <= layer3_outputs(129);
    layer4_outputs(991) <= (layer3_outputs(731)) and (layer3_outputs(8148));
    layer4_outputs(992) <= (layer3_outputs(8788)) xor (layer3_outputs(5409));
    layer4_outputs(993) <= not((layer3_outputs(5966)) and (layer3_outputs(8813)));
    layer4_outputs(994) <= not((layer3_outputs(6640)) xor (layer3_outputs(9447)));
    layer4_outputs(995) <= (layer3_outputs(2005)) and not (layer3_outputs(8051));
    layer4_outputs(996) <= not(layer3_outputs(5042)) or (layer3_outputs(695));
    layer4_outputs(997) <= not((layer3_outputs(1433)) and (layer3_outputs(879)));
    layer4_outputs(998) <= layer3_outputs(5874);
    layer4_outputs(999) <= not(layer3_outputs(963));
    layer4_outputs(1000) <= layer3_outputs(4803);
    layer4_outputs(1001) <= not(layer3_outputs(4603));
    layer4_outputs(1002) <= not(layer3_outputs(10056));
    layer4_outputs(1003) <= (layer3_outputs(8143)) xor (layer3_outputs(5301));
    layer4_outputs(1004) <= not((layer3_outputs(8002)) xor (layer3_outputs(9780)));
    layer4_outputs(1005) <= layer3_outputs(1413);
    layer4_outputs(1006) <= layer3_outputs(6922);
    layer4_outputs(1007) <= not(layer3_outputs(6820));
    layer4_outputs(1008) <= not(layer3_outputs(196)) or (layer3_outputs(5096));
    layer4_outputs(1009) <= (layer3_outputs(575)) xor (layer3_outputs(9219));
    layer4_outputs(1010) <= layer3_outputs(6219);
    layer4_outputs(1011) <= not(layer3_outputs(9390)) or (layer3_outputs(979));
    layer4_outputs(1012) <= not(layer3_outputs(7496)) or (layer3_outputs(6844));
    layer4_outputs(1013) <= layer3_outputs(7424);
    layer4_outputs(1014) <= not(layer3_outputs(2166));
    layer4_outputs(1015) <= not(layer3_outputs(744));
    layer4_outputs(1016) <= not((layer3_outputs(8650)) xor (layer3_outputs(2235)));
    layer4_outputs(1017) <= layer3_outputs(607);
    layer4_outputs(1018) <= not((layer3_outputs(9150)) xor (layer3_outputs(5737)));
    layer4_outputs(1019) <= '0';
    layer4_outputs(1020) <= not((layer3_outputs(2859)) or (layer3_outputs(9319)));
    layer4_outputs(1021) <= not(layer3_outputs(7918));
    layer4_outputs(1022) <= layer3_outputs(2770);
    layer4_outputs(1023) <= layer3_outputs(3978);
    layer4_outputs(1024) <= not(layer3_outputs(9041));
    layer4_outputs(1025) <= layer3_outputs(8857);
    layer4_outputs(1026) <= layer3_outputs(7656);
    layer4_outputs(1027) <= layer3_outputs(9052);
    layer4_outputs(1028) <= (layer3_outputs(3486)) xor (layer3_outputs(613));
    layer4_outputs(1029) <= (layer3_outputs(2505)) and (layer3_outputs(1705));
    layer4_outputs(1030) <= layer3_outputs(3791);
    layer4_outputs(1031) <= (layer3_outputs(6193)) and (layer3_outputs(6654));
    layer4_outputs(1032) <= not(layer3_outputs(2143));
    layer4_outputs(1033) <= (layer3_outputs(4941)) xor (layer3_outputs(2592));
    layer4_outputs(1034) <= not((layer3_outputs(2834)) and (layer3_outputs(5628)));
    layer4_outputs(1035) <= (layer3_outputs(2240)) xor (layer3_outputs(1575));
    layer4_outputs(1036) <= layer3_outputs(2776);
    layer4_outputs(1037) <= not(layer3_outputs(6370));
    layer4_outputs(1038) <= not(layer3_outputs(9509));
    layer4_outputs(1039) <= (layer3_outputs(6381)) or (layer3_outputs(915));
    layer4_outputs(1040) <= not((layer3_outputs(3398)) and (layer3_outputs(467)));
    layer4_outputs(1041) <= not(layer3_outputs(440)) or (layer3_outputs(6631));
    layer4_outputs(1042) <= not(layer3_outputs(8778));
    layer4_outputs(1043) <= not(layer3_outputs(5962));
    layer4_outputs(1044) <= layer3_outputs(9164);
    layer4_outputs(1045) <= layer3_outputs(1570);
    layer4_outputs(1046) <= layer3_outputs(9023);
    layer4_outputs(1047) <= layer3_outputs(5575);
    layer4_outputs(1048) <= layer3_outputs(5371);
    layer4_outputs(1049) <= not(layer3_outputs(1412)) or (layer3_outputs(8821));
    layer4_outputs(1050) <= not((layer3_outputs(3876)) xor (layer3_outputs(5975)));
    layer4_outputs(1051) <= (layer3_outputs(8287)) xor (layer3_outputs(8989));
    layer4_outputs(1052) <= not(layer3_outputs(3671));
    layer4_outputs(1053) <= '0';
    layer4_outputs(1054) <= not((layer3_outputs(1168)) xor (layer3_outputs(1530)));
    layer4_outputs(1055) <= not((layer3_outputs(4719)) xor (layer3_outputs(2763)));
    layer4_outputs(1056) <= (layer3_outputs(4925)) xor (layer3_outputs(522));
    layer4_outputs(1057) <= layer3_outputs(7111);
    layer4_outputs(1058) <= layer3_outputs(4218);
    layer4_outputs(1059) <= (layer3_outputs(4613)) or (layer3_outputs(8120));
    layer4_outputs(1060) <= not((layer3_outputs(696)) xor (layer3_outputs(10144)));
    layer4_outputs(1061) <= not((layer3_outputs(9901)) xor (layer3_outputs(7875)));
    layer4_outputs(1062) <= (layer3_outputs(2851)) and not (layer3_outputs(1801));
    layer4_outputs(1063) <= not((layer3_outputs(8230)) xor (layer3_outputs(4728)));
    layer4_outputs(1064) <= (layer3_outputs(4011)) and (layer3_outputs(269));
    layer4_outputs(1065) <= layer3_outputs(4073);
    layer4_outputs(1066) <= (layer3_outputs(1152)) and (layer3_outputs(3935));
    layer4_outputs(1067) <= (layer3_outputs(6254)) and (layer3_outputs(520));
    layer4_outputs(1068) <= (layer3_outputs(4820)) xor (layer3_outputs(143));
    layer4_outputs(1069) <= not((layer3_outputs(2795)) or (layer3_outputs(5715)));
    layer4_outputs(1070) <= not((layer3_outputs(586)) xor (layer3_outputs(1641)));
    layer4_outputs(1071) <= (layer3_outputs(2977)) and not (layer3_outputs(3907));
    layer4_outputs(1072) <= layer3_outputs(2965);
    layer4_outputs(1073) <= layer3_outputs(3932);
    layer4_outputs(1074) <= layer3_outputs(935);
    layer4_outputs(1075) <= not(layer3_outputs(2637));
    layer4_outputs(1076) <= not((layer3_outputs(2165)) xor (layer3_outputs(5517)));
    layer4_outputs(1077) <= not(layer3_outputs(1412)) or (layer3_outputs(6537));
    layer4_outputs(1078) <= not(layer3_outputs(2681));
    layer4_outputs(1079) <= not(layer3_outputs(1625)) or (layer3_outputs(8855));
    layer4_outputs(1080) <= not(layer3_outputs(8866)) or (layer3_outputs(9524));
    layer4_outputs(1081) <= not(layer3_outputs(2996)) or (layer3_outputs(2434));
    layer4_outputs(1082) <= layer3_outputs(3117);
    layer4_outputs(1083) <= layer3_outputs(222);
    layer4_outputs(1084) <= not((layer3_outputs(6261)) or (layer3_outputs(6033)));
    layer4_outputs(1085) <= (layer3_outputs(9387)) and not (layer3_outputs(2662));
    layer4_outputs(1086) <= layer3_outputs(5035);
    layer4_outputs(1087) <= layer3_outputs(113);
    layer4_outputs(1088) <= not(layer3_outputs(10043));
    layer4_outputs(1089) <= (layer3_outputs(9755)) xor (layer3_outputs(3090));
    layer4_outputs(1090) <= (layer3_outputs(7529)) xor (layer3_outputs(8399));
    layer4_outputs(1091) <= not(layer3_outputs(7706));
    layer4_outputs(1092) <= layer3_outputs(1367);
    layer4_outputs(1093) <= not(layer3_outputs(4640));
    layer4_outputs(1094) <= (layer3_outputs(3093)) and not (layer3_outputs(1245));
    layer4_outputs(1095) <= layer3_outputs(5596);
    layer4_outputs(1096) <= not(layer3_outputs(890));
    layer4_outputs(1097) <= not(layer3_outputs(2476));
    layer4_outputs(1098) <= (layer3_outputs(364)) xor (layer3_outputs(7822));
    layer4_outputs(1099) <= (layer3_outputs(10045)) and not (layer3_outputs(2022));
    layer4_outputs(1100) <= not((layer3_outputs(6355)) or (layer3_outputs(2987)));
    layer4_outputs(1101) <= not(layer3_outputs(6260)) or (layer3_outputs(9344));
    layer4_outputs(1102) <= (layer3_outputs(8199)) and (layer3_outputs(9902));
    layer4_outputs(1103) <= layer3_outputs(1889);
    layer4_outputs(1104) <= layer3_outputs(4738);
    layer4_outputs(1105) <= layer3_outputs(10051);
    layer4_outputs(1106) <= layer3_outputs(9508);
    layer4_outputs(1107) <= not(layer3_outputs(3607));
    layer4_outputs(1108) <= '0';
    layer4_outputs(1109) <= not(layer3_outputs(5979));
    layer4_outputs(1110) <= layer3_outputs(1729);
    layer4_outputs(1111) <= not(layer3_outputs(3893));
    layer4_outputs(1112) <= (layer3_outputs(4445)) and (layer3_outputs(1344));
    layer4_outputs(1113) <= (layer3_outputs(5229)) or (layer3_outputs(4511));
    layer4_outputs(1114) <= '1';
    layer4_outputs(1115) <= not(layer3_outputs(6634));
    layer4_outputs(1116) <= not((layer3_outputs(2752)) xor (layer3_outputs(5541)));
    layer4_outputs(1117) <= (layer3_outputs(2818)) or (layer3_outputs(233));
    layer4_outputs(1118) <= (layer3_outputs(8383)) xor (layer3_outputs(8240));
    layer4_outputs(1119) <= (layer3_outputs(5390)) and not (layer3_outputs(4334));
    layer4_outputs(1120) <= not(layer3_outputs(430));
    layer4_outputs(1121) <= layer3_outputs(4418);
    layer4_outputs(1122) <= not(layer3_outputs(3943));
    layer4_outputs(1123) <= (layer3_outputs(17)) and not (layer3_outputs(8534));
    layer4_outputs(1124) <= layer3_outputs(9242);
    layer4_outputs(1125) <= not((layer3_outputs(5310)) xor (layer3_outputs(1600)));
    layer4_outputs(1126) <= layer3_outputs(2171);
    layer4_outputs(1127) <= layer3_outputs(4120);
    layer4_outputs(1128) <= not((layer3_outputs(4836)) or (layer3_outputs(6887)));
    layer4_outputs(1129) <= (layer3_outputs(7212)) xor (layer3_outputs(8027));
    layer4_outputs(1130) <= layer3_outputs(2354);
    layer4_outputs(1131) <= layer3_outputs(8947);
    layer4_outputs(1132) <= layer3_outputs(5702);
    layer4_outputs(1133) <= not(layer3_outputs(7768));
    layer4_outputs(1134) <= not(layer3_outputs(1062)) or (layer3_outputs(2658));
    layer4_outputs(1135) <= not((layer3_outputs(1183)) and (layer3_outputs(3075)));
    layer4_outputs(1136) <= layer3_outputs(1928);
    layer4_outputs(1137) <= not(layer3_outputs(2277));
    layer4_outputs(1138) <= not((layer3_outputs(8464)) xor (layer3_outputs(4961)));
    layer4_outputs(1139) <= layer3_outputs(6031);
    layer4_outputs(1140) <= layer3_outputs(4220);
    layer4_outputs(1141) <= (layer3_outputs(1608)) and (layer3_outputs(9466));
    layer4_outputs(1142) <= (layer3_outputs(7286)) or (layer3_outputs(8909));
    layer4_outputs(1143) <= layer3_outputs(8968);
    layer4_outputs(1144) <= not((layer3_outputs(3987)) xor (layer3_outputs(7832)));
    layer4_outputs(1145) <= (layer3_outputs(5880)) and not (layer3_outputs(7460));
    layer4_outputs(1146) <= (layer3_outputs(1825)) or (layer3_outputs(395));
    layer4_outputs(1147) <= not((layer3_outputs(195)) xor (layer3_outputs(4167)));
    layer4_outputs(1148) <= not((layer3_outputs(2815)) and (layer3_outputs(715)));
    layer4_outputs(1149) <= layer3_outputs(8902);
    layer4_outputs(1150) <= (layer3_outputs(3950)) xor (layer3_outputs(4468));
    layer4_outputs(1151) <= layer3_outputs(8286);
    layer4_outputs(1152) <= not(layer3_outputs(7283));
    layer4_outputs(1153) <= not(layer3_outputs(9587));
    layer4_outputs(1154) <= layer3_outputs(2578);
    layer4_outputs(1155) <= not((layer3_outputs(713)) or (layer3_outputs(8452)));
    layer4_outputs(1156) <= layer3_outputs(550);
    layer4_outputs(1157) <= not(layer3_outputs(7192));
    layer4_outputs(1158) <= not(layer3_outputs(5126)) or (layer3_outputs(1117));
    layer4_outputs(1159) <= (layer3_outputs(5671)) xor (layer3_outputs(6453));
    layer4_outputs(1160) <= layer3_outputs(6147);
    layer4_outputs(1161) <= layer3_outputs(5354);
    layer4_outputs(1162) <= layer3_outputs(6578);
    layer4_outputs(1163) <= not(layer3_outputs(1432));
    layer4_outputs(1164) <= not((layer3_outputs(961)) or (layer3_outputs(8157)));
    layer4_outputs(1165) <= layer3_outputs(6693);
    layer4_outputs(1166) <= not((layer3_outputs(7845)) or (layer3_outputs(6963)));
    layer4_outputs(1167) <= not((layer3_outputs(2457)) xor (layer3_outputs(4699)));
    layer4_outputs(1168) <= '0';
    layer4_outputs(1169) <= (layer3_outputs(326)) and not (layer3_outputs(3110));
    layer4_outputs(1170) <= not(layer3_outputs(2270)) or (layer3_outputs(2509));
    layer4_outputs(1171) <= (layer3_outputs(6792)) and not (layer3_outputs(6492));
    layer4_outputs(1172) <= (layer3_outputs(9222)) and not (layer3_outputs(7912));
    layer4_outputs(1173) <= (layer3_outputs(5199)) and not (layer3_outputs(3213));
    layer4_outputs(1174) <= layer3_outputs(6066);
    layer4_outputs(1175) <= layer3_outputs(7853);
    layer4_outputs(1176) <= layer3_outputs(7472);
    layer4_outputs(1177) <= not((layer3_outputs(2355)) and (layer3_outputs(9104)));
    layer4_outputs(1178) <= layer3_outputs(9581);
    layer4_outputs(1179) <= not(layer3_outputs(593));
    layer4_outputs(1180) <= not((layer3_outputs(2268)) xor (layer3_outputs(10162)));
    layer4_outputs(1181) <= (layer3_outputs(3574)) or (layer3_outputs(9250));
    layer4_outputs(1182) <= (layer3_outputs(7710)) and (layer3_outputs(5688));
    layer4_outputs(1183) <= (layer3_outputs(5443)) or (layer3_outputs(2290));
    layer4_outputs(1184) <= (layer3_outputs(169)) and (layer3_outputs(3480));
    layer4_outputs(1185) <= not((layer3_outputs(7077)) and (layer3_outputs(4200)));
    layer4_outputs(1186) <= not(layer3_outputs(992));
    layer4_outputs(1187) <= not((layer3_outputs(7712)) and (layer3_outputs(818)));
    layer4_outputs(1188) <= layer3_outputs(2046);
    layer4_outputs(1189) <= (layer3_outputs(8974)) and (layer3_outputs(5588));
    layer4_outputs(1190) <= not(layer3_outputs(1632));
    layer4_outputs(1191) <= layer3_outputs(8155);
    layer4_outputs(1192) <= layer3_outputs(4626);
    layer4_outputs(1193) <= not(layer3_outputs(8387)) or (layer3_outputs(10137));
    layer4_outputs(1194) <= layer3_outputs(9649);
    layer4_outputs(1195) <= layer3_outputs(731);
    layer4_outputs(1196) <= (layer3_outputs(8244)) and not (layer3_outputs(6717));
    layer4_outputs(1197) <= layer3_outputs(10094);
    layer4_outputs(1198) <= layer3_outputs(9260);
    layer4_outputs(1199) <= (layer3_outputs(4478)) or (layer3_outputs(831));
    layer4_outputs(1200) <= not((layer3_outputs(738)) and (layer3_outputs(5044)));
    layer4_outputs(1201) <= layer3_outputs(6098);
    layer4_outputs(1202) <= layer3_outputs(8396);
    layer4_outputs(1203) <= (layer3_outputs(2150)) or (layer3_outputs(7766));
    layer4_outputs(1204) <= not((layer3_outputs(980)) or (layer3_outputs(6095)));
    layer4_outputs(1205) <= (layer3_outputs(7531)) xor (layer3_outputs(6529));
    layer4_outputs(1206) <= not((layer3_outputs(5169)) xor (layer3_outputs(4766)));
    layer4_outputs(1207) <= (layer3_outputs(2718)) or (layer3_outputs(1070));
    layer4_outputs(1208) <= '1';
    layer4_outputs(1209) <= layer3_outputs(3102);
    layer4_outputs(1210) <= not(layer3_outputs(1468));
    layer4_outputs(1211) <= not(layer3_outputs(9048)) or (layer3_outputs(1662));
    layer4_outputs(1212) <= (layer3_outputs(7567)) and not (layer3_outputs(7059));
    layer4_outputs(1213) <= not((layer3_outputs(2002)) or (layer3_outputs(9783)));
    layer4_outputs(1214) <= not(layer3_outputs(3105));
    layer4_outputs(1215) <= layer3_outputs(4128);
    layer4_outputs(1216) <= not(layer3_outputs(6206));
    layer4_outputs(1217) <= not((layer3_outputs(9118)) or (layer3_outputs(5372)));
    layer4_outputs(1218) <= (layer3_outputs(4003)) or (layer3_outputs(270));
    layer4_outputs(1219) <= not(layer3_outputs(8681));
    layer4_outputs(1220) <= not(layer3_outputs(4141));
    layer4_outputs(1221) <= layer3_outputs(2154);
    layer4_outputs(1222) <= not(layer3_outputs(6829)) or (layer3_outputs(2701));
    layer4_outputs(1223) <= (layer3_outputs(9857)) xor (layer3_outputs(9469));
    layer4_outputs(1224) <= not(layer3_outputs(6262)) or (layer3_outputs(1384));
    layer4_outputs(1225) <= not(layer3_outputs(9873));
    layer4_outputs(1226) <= (layer3_outputs(9819)) and (layer3_outputs(3769));
    layer4_outputs(1227) <= not((layer3_outputs(7788)) or (layer3_outputs(5186)));
    layer4_outputs(1228) <= (layer3_outputs(671)) and not (layer3_outputs(5100));
    layer4_outputs(1229) <= layer3_outputs(5739);
    layer4_outputs(1230) <= not(layer3_outputs(1146));
    layer4_outputs(1231) <= '0';
    layer4_outputs(1232) <= (layer3_outputs(3331)) and not (layer3_outputs(2318));
    layer4_outputs(1233) <= not(layer3_outputs(4865));
    layer4_outputs(1234) <= layer3_outputs(5275);
    layer4_outputs(1235) <= not((layer3_outputs(6332)) or (layer3_outputs(1306)));
    layer4_outputs(1236) <= layer3_outputs(3439);
    layer4_outputs(1237) <= not(layer3_outputs(6350));
    layer4_outputs(1238) <= not(layer3_outputs(8804));
    layer4_outputs(1239) <= not(layer3_outputs(2189));
    layer4_outputs(1240) <= not(layer3_outputs(10012));
    layer4_outputs(1241) <= layer3_outputs(9910);
    layer4_outputs(1242) <= not(layer3_outputs(6883));
    layer4_outputs(1243) <= (layer3_outputs(7597)) and not (layer3_outputs(4818));
    layer4_outputs(1244) <= (layer3_outputs(7435)) or (layer3_outputs(8496));
    layer4_outputs(1245) <= not(layer3_outputs(1264));
    layer4_outputs(1246) <= not((layer3_outputs(7091)) xor (layer3_outputs(4500)));
    layer4_outputs(1247) <= layer3_outputs(4524);
    layer4_outputs(1248) <= (layer3_outputs(6596)) and (layer3_outputs(4898));
    layer4_outputs(1249) <= not(layer3_outputs(8233));
    layer4_outputs(1250) <= not(layer3_outputs(403));
    layer4_outputs(1251) <= not(layer3_outputs(9910)) or (layer3_outputs(6419));
    layer4_outputs(1252) <= (layer3_outputs(9951)) and not (layer3_outputs(9965));
    layer4_outputs(1253) <= layer3_outputs(3770);
    layer4_outputs(1254) <= layer3_outputs(6073);
    layer4_outputs(1255) <= not((layer3_outputs(331)) xor (layer3_outputs(714)));
    layer4_outputs(1256) <= '1';
    layer4_outputs(1257) <= not(layer3_outputs(8192));
    layer4_outputs(1258) <= layer3_outputs(4355);
    layer4_outputs(1259) <= not(layer3_outputs(7180));
    layer4_outputs(1260) <= (layer3_outputs(889)) xor (layer3_outputs(4439));
    layer4_outputs(1261) <= layer3_outputs(9351);
    layer4_outputs(1262) <= not(layer3_outputs(798));
    layer4_outputs(1263) <= layer3_outputs(7730);
    layer4_outputs(1264) <= not(layer3_outputs(2807));
    layer4_outputs(1265) <= not((layer3_outputs(4894)) xor (layer3_outputs(684)));
    layer4_outputs(1266) <= layer3_outputs(2202);
    layer4_outputs(1267) <= (layer3_outputs(4836)) xor (layer3_outputs(546));
    layer4_outputs(1268) <= not(layer3_outputs(3679)) or (layer3_outputs(3280));
    layer4_outputs(1269) <= (layer3_outputs(2733)) and (layer3_outputs(7001));
    layer4_outputs(1270) <= not(layer3_outputs(9151));
    layer4_outputs(1271) <= not(layer3_outputs(2012)) or (layer3_outputs(7528));
    layer4_outputs(1272) <= not(layer3_outputs(6227)) or (layer3_outputs(896));
    layer4_outputs(1273) <= (layer3_outputs(9385)) and not (layer3_outputs(6484));
    layer4_outputs(1274) <= not((layer3_outputs(2195)) and (layer3_outputs(4917)));
    layer4_outputs(1275) <= not((layer3_outputs(1184)) xor (layer3_outputs(4310)));
    layer4_outputs(1276) <= not(layer3_outputs(1001));
    layer4_outputs(1277) <= (layer3_outputs(5105)) and not (layer3_outputs(6549));
    layer4_outputs(1278) <= not(layer3_outputs(5583));
    layer4_outputs(1279) <= not(layer3_outputs(8075));
    layer4_outputs(1280) <= not(layer3_outputs(753));
    layer4_outputs(1281) <= (layer3_outputs(8264)) and not (layer3_outputs(5364));
    layer4_outputs(1282) <= (layer3_outputs(6746)) xor (layer3_outputs(9135));
    layer4_outputs(1283) <= layer3_outputs(6577);
    layer4_outputs(1284) <= not((layer3_outputs(7769)) xor (layer3_outputs(52)));
    layer4_outputs(1285) <= not(layer3_outputs(7610));
    layer4_outputs(1286) <= not(layer3_outputs(5631));
    layer4_outputs(1287) <= layer3_outputs(3643);
    layer4_outputs(1288) <= layer3_outputs(5228);
    layer4_outputs(1289) <= not(layer3_outputs(2490));
    layer4_outputs(1290) <= (layer3_outputs(8752)) and not (layer3_outputs(6686));
    layer4_outputs(1291) <= layer3_outputs(3443);
    layer4_outputs(1292) <= (layer3_outputs(2524)) and not (layer3_outputs(1153));
    layer4_outputs(1293) <= not(layer3_outputs(5640));
    layer4_outputs(1294) <= layer3_outputs(4877);
    layer4_outputs(1295) <= (layer3_outputs(880)) xor (layer3_outputs(8060));
    layer4_outputs(1296) <= (layer3_outputs(4990)) and not (layer3_outputs(4795));
    layer4_outputs(1297) <= not(layer3_outputs(6228));
    layer4_outputs(1298) <= layer3_outputs(23);
    layer4_outputs(1299) <= not(layer3_outputs(1478));
    layer4_outputs(1300) <= not((layer3_outputs(4574)) xor (layer3_outputs(1833)));
    layer4_outputs(1301) <= layer3_outputs(5666);
    layer4_outputs(1302) <= not(layer3_outputs(3755));
    layer4_outputs(1303) <= not(layer3_outputs(70));
    layer4_outputs(1304) <= layer3_outputs(8047);
    layer4_outputs(1305) <= not((layer3_outputs(3847)) xor (layer3_outputs(3753)));
    layer4_outputs(1306) <= layer3_outputs(8088);
    layer4_outputs(1307) <= not(layer3_outputs(7568));
    layer4_outputs(1308) <= layer3_outputs(2841);
    layer4_outputs(1309) <= layer3_outputs(1128);
    layer4_outputs(1310) <= (layer3_outputs(1252)) and not (layer3_outputs(10106));
    layer4_outputs(1311) <= not(layer3_outputs(2776));
    layer4_outputs(1312) <= not(layer3_outputs(5131));
    layer4_outputs(1313) <= layer3_outputs(2257);
    layer4_outputs(1314) <= not(layer3_outputs(2987));
    layer4_outputs(1315) <= not(layer3_outputs(6827));
    layer4_outputs(1316) <= not(layer3_outputs(887));
    layer4_outputs(1317) <= not(layer3_outputs(6588));
    layer4_outputs(1318) <= (layer3_outputs(6673)) or (layer3_outputs(2443));
    layer4_outputs(1319) <= not(layer3_outputs(1922)) or (layer3_outputs(5225));
    layer4_outputs(1320) <= not((layer3_outputs(6239)) xor (layer3_outputs(9898)));
    layer4_outputs(1321) <= not(layer3_outputs(1020)) or (layer3_outputs(5341));
    layer4_outputs(1322) <= (layer3_outputs(7888)) or (layer3_outputs(7065));
    layer4_outputs(1323) <= not(layer3_outputs(5147));
    layer4_outputs(1324) <= not(layer3_outputs(9834));
    layer4_outputs(1325) <= layer3_outputs(9061);
    layer4_outputs(1326) <= (layer3_outputs(497)) and not (layer3_outputs(4318));
    layer4_outputs(1327) <= layer3_outputs(8203);
    layer4_outputs(1328) <= '1';
    layer4_outputs(1329) <= not(layer3_outputs(5628));
    layer4_outputs(1330) <= layer3_outputs(9014);
    layer4_outputs(1331) <= layer3_outputs(8411);
    layer4_outputs(1332) <= (layer3_outputs(5065)) xor (layer3_outputs(9326));
    layer4_outputs(1333) <= not(layer3_outputs(8344)) or (layer3_outputs(2720));
    layer4_outputs(1334) <= layer3_outputs(2691);
    layer4_outputs(1335) <= layer3_outputs(9527);
    layer4_outputs(1336) <= layer3_outputs(7142);
    layer4_outputs(1337) <= not(layer3_outputs(1176));
    layer4_outputs(1338) <= layer3_outputs(3992);
    layer4_outputs(1339) <= layer3_outputs(3099);
    layer4_outputs(1340) <= not(layer3_outputs(6535));
    layer4_outputs(1341) <= (layer3_outputs(2668)) xor (layer3_outputs(7538));
    layer4_outputs(1342) <= layer3_outputs(2277);
    layer4_outputs(1343) <= not((layer3_outputs(421)) and (layer3_outputs(6354)));
    layer4_outputs(1344) <= not(layer3_outputs(7534));
    layer4_outputs(1345) <= not(layer3_outputs(3799));
    layer4_outputs(1346) <= layer3_outputs(8805);
    layer4_outputs(1347) <= not(layer3_outputs(9064)) or (layer3_outputs(1239));
    layer4_outputs(1348) <= (layer3_outputs(128)) xor (layer3_outputs(2962));
    layer4_outputs(1349) <= layer3_outputs(6903);
    layer4_outputs(1350) <= layer3_outputs(9667);
    layer4_outputs(1351) <= layer3_outputs(6530);
    layer4_outputs(1352) <= not(layer3_outputs(9853));
    layer4_outputs(1353) <= (layer3_outputs(7574)) xor (layer3_outputs(3264));
    layer4_outputs(1354) <= (layer3_outputs(1576)) xor (layer3_outputs(2762));
    layer4_outputs(1355) <= not(layer3_outputs(6061)) or (layer3_outputs(1392));
    layer4_outputs(1356) <= layer3_outputs(2200);
    layer4_outputs(1357) <= not(layer3_outputs(8222)) or (layer3_outputs(908));
    layer4_outputs(1358) <= layer3_outputs(3295);
    layer4_outputs(1359) <= (layer3_outputs(8566)) or (layer3_outputs(4177));
    layer4_outputs(1360) <= not((layer3_outputs(5920)) or (layer3_outputs(1532)));
    layer4_outputs(1361) <= not((layer3_outputs(7868)) and (layer3_outputs(8511)));
    layer4_outputs(1362) <= not(layer3_outputs(529));
    layer4_outputs(1363) <= not(layer3_outputs(4817));
    layer4_outputs(1364) <= not((layer3_outputs(2966)) xor (layer3_outputs(9207)));
    layer4_outputs(1365) <= not((layer3_outputs(9962)) or (layer3_outputs(9958)));
    layer4_outputs(1366) <= not(layer3_outputs(9682)) or (layer3_outputs(1334));
    layer4_outputs(1367) <= not(layer3_outputs(7395));
    layer4_outputs(1368) <= layer3_outputs(3947);
    layer4_outputs(1369) <= layer3_outputs(529);
    layer4_outputs(1370) <= not((layer3_outputs(6710)) and (layer3_outputs(9028)));
    layer4_outputs(1371) <= not(layer3_outputs(58)) or (layer3_outputs(7742));
    layer4_outputs(1372) <= (layer3_outputs(8227)) and not (layer3_outputs(9487));
    layer4_outputs(1373) <= not(layer3_outputs(4345));
    layer4_outputs(1374) <= layer3_outputs(2878);
    layer4_outputs(1375) <= not((layer3_outputs(4921)) and (layer3_outputs(4244)));
    layer4_outputs(1376) <= (layer3_outputs(7116)) xor (layer3_outputs(6212));
    layer4_outputs(1377) <= not((layer3_outputs(7604)) and (layer3_outputs(8293)));
    layer4_outputs(1378) <= (layer3_outputs(4043)) and not (layer3_outputs(7703));
    layer4_outputs(1379) <= not((layer3_outputs(4991)) xor (layer3_outputs(2266)));
    layer4_outputs(1380) <= (layer3_outputs(2297)) and not (layer3_outputs(6981));
    layer4_outputs(1381) <= (layer3_outputs(904)) xor (layer3_outputs(9855));
    layer4_outputs(1382) <= not(layer3_outputs(4550)) or (layer3_outputs(5785));
    layer4_outputs(1383) <= (layer3_outputs(26)) or (layer3_outputs(813));
    layer4_outputs(1384) <= (layer3_outputs(763)) and not (layer3_outputs(8474));
    layer4_outputs(1385) <= not(layer3_outputs(804));
    layer4_outputs(1386) <= not(layer3_outputs(7067));
    layer4_outputs(1387) <= not(layer3_outputs(9959)) or (layer3_outputs(1283));
    layer4_outputs(1388) <= (layer3_outputs(5243)) and (layer3_outputs(6109));
    layer4_outputs(1389) <= not((layer3_outputs(6867)) or (layer3_outputs(3527)));
    layer4_outputs(1390) <= layer3_outputs(22);
    layer4_outputs(1391) <= not(layer3_outputs(2077));
    layer4_outputs(1392) <= not(layer3_outputs(1756)) or (layer3_outputs(6688));
    layer4_outputs(1393) <= not((layer3_outputs(8117)) xor (layer3_outputs(6416)));
    layer4_outputs(1394) <= layer3_outputs(460);
    layer4_outputs(1395) <= (layer3_outputs(5906)) xor (layer3_outputs(5454));
    layer4_outputs(1396) <= (layer3_outputs(7712)) xor (layer3_outputs(350));
    layer4_outputs(1397) <= (layer3_outputs(302)) or (layer3_outputs(1724));
    layer4_outputs(1398) <= layer3_outputs(10070);
    layer4_outputs(1399) <= not(layer3_outputs(5521));
    layer4_outputs(1400) <= not(layer3_outputs(640));
    layer4_outputs(1401) <= not(layer3_outputs(4702));
    layer4_outputs(1402) <= not(layer3_outputs(3042)) or (layer3_outputs(6052));
    layer4_outputs(1403) <= layer3_outputs(6857);
    layer4_outputs(1404) <= layer3_outputs(3434);
    layer4_outputs(1405) <= not(layer3_outputs(2806));
    layer4_outputs(1406) <= not(layer3_outputs(7620));
    layer4_outputs(1407) <= not((layer3_outputs(1552)) xor (layer3_outputs(1081)));
    layer4_outputs(1408) <= layer3_outputs(7780);
    layer4_outputs(1409) <= (layer3_outputs(9641)) and not (layer3_outputs(5228));
    layer4_outputs(1410) <= (layer3_outputs(8166)) xor (layer3_outputs(364));
    layer4_outputs(1411) <= layer3_outputs(5874);
    layer4_outputs(1412) <= not(layer3_outputs(9008));
    layer4_outputs(1413) <= not(layer3_outputs(5735));
    layer4_outputs(1414) <= not((layer3_outputs(6371)) and (layer3_outputs(1032)));
    layer4_outputs(1415) <= layer3_outputs(7958);
    layer4_outputs(1416) <= (layer3_outputs(7552)) and not (layer3_outputs(1170));
    layer4_outputs(1417) <= (layer3_outputs(5810)) xor (layer3_outputs(8221));
    layer4_outputs(1418) <= not((layer3_outputs(8961)) or (layer3_outputs(553)));
    layer4_outputs(1419) <= not((layer3_outputs(3436)) xor (layer3_outputs(6164)));
    layer4_outputs(1420) <= not(layer3_outputs(1557)) or (layer3_outputs(4267));
    layer4_outputs(1421) <= (layer3_outputs(3457)) xor (layer3_outputs(4415));
    layer4_outputs(1422) <= not(layer3_outputs(9287));
    layer4_outputs(1423) <= not(layer3_outputs(652));
    layer4_outputs(1424) <= layer3_outputs(4147);
    layer4_outputs(1425) <= (layer3_outputs(6976)) or (layer3_outputs(5988));
    layer4_outputs(1426) <= layer3_outputs(6637);
    layer4_outputs(1427) <= (layer3_outputs(3422)) and (layer3_outputs(5554));
    layer4_outputs(1428) <= not(layer3_outputs(508));
    layer4_outputs(1429) <= layer3_outputs(4982);
    layer4_outputs(1430) <= not(layer3_outputs(5370));
    layer4_outputs(1431) <= layer3_outputs(5295);
    layer4_outputs(1432) <= layer3_outputs(12);
    layer4_outputs(1433) <= layer3_outputs(2206);
    layer4_outputs(1434) <= (layer3_outputs(2513)) and not (layer3_outputs(4766));
    layer4_outputs(1435) <= not((layer3_outputs(7469)) and (layer3_outputs(2760)));
    layer4_outputs(1436) <= not(layer3_outputs(2498));
    layer4_outputs(1437) <= not(layer3_outputs(204)) or (layer3_outputs(1819));
    layer4_outputs(1438) <= not((layer3_outputs(4948)) and (layer3_outputs(8779)));
    layer4_outputs(1439) <= not(layer3_outputs(9203));
    layer4_outputs(1440) <= (layer3_outputs(1994)) and not (layer3_outputs(7413));
    layer4_outputs(1441) <= not(layer3_outputs(1518));
    layer4_outputs(1442) <= not(layer3_outputs(1441));
    layer4_outputs(1443) <= not((layer3_outputs(8941)) and (layer3_outputs(9304)));
    layer4_outputs(1444) <= not(layer3_outputs(3743));
    layer4_outputs(1445) <= (layer3_outputs(6983)) and not (layer3_outputs(6079));
    layer4_outputs(1446) <= (layer3_outputs(5193)) xor (layer3_outputs(4352));
    layer4_outputs(1447) <= (layer3_outputs(3442)) and (layer3_outputs(8683));
    layer4_outputs(1448) <= not(layer3_outputs(5954)) or (layer3_outputs(7077));
    layer4_outputs(1449) <= layer3_outputs(5100);
    layer4_outputs(1450) <= (layer3_outputs(7863)) or (layer3_outputs(9472));
    layer4_outputs(1451) <= layer3_outputs(4261);
    layer4_outputs(1452) <= (layer3_outputs(2893)) and not (layer3_outputs(9893));
    layer4_outputs(1453) <= not((layer3_outputs(4571)) xor (layer3_outputs(1133)));
    layer4_outputs(1454) <= not(layer3_outputs(2925));
    layer4_outputs(1455) <= not(layer3_outputs(9399));
    layer4_outputs(1456) <= not((layer3_outputs(10199)) or (layer3_outputs(3566)));
    layer4_outputs(1457) <= not(layer3_outputs(6044)) or (layer3_outputs(9010));
    layer4_outputs(1458) <= not(layer3_outputs(6383)) or (layer3_outputs(5805));
    layer4_outputs(1459) <= not((layer3_outputs(2196)) and (layer3_outputs(5538)));
    layer4_outputs(1460) <= '1';
    layer4_outputs(1461) <= not((layer3_outputs(9376)) and (layer3_outputs(6179)));
    layer4_outputs(1462) <= not(layer3_outputs(3657));
    layer4_outputs(1463) <= (layer3_outputs(2997)) xor (layer3_outputs(4796));
    layer4_outputs(1464) <= not(layer3_outputs(400));
    layer4_outputs(1465) <= not(layer3_outputs(6572)) or (layer3_outputs(9532));
    layer4_outputs(1466) <= layer3_outputs(4665);
    layer4_outputs(1467) <= not(layer3_outputs(6591));
    layer4_outputs(1468) <= not(layer3_outputs(8131));
    layer4_outputs(1469) <= not(layer3_outputs(3779));
    layer4_outputs(1470) <= layer3_outputs(4816);
    layer4_outputs(1471) <= not((layer3_outputs(5413)) xor (layer3_outputs(9709)));
    layer4_outputs(1472) <= layer3_outputs(6645);
    layer4_outputs(1473) <= layer3_outputs(7007);
    layer4_outputs(1474) <= layer3_outputs(8874);
    layer4_outputs(1475) <= (layer3_outputs(9556)) and (layer3_outputs(4751));
    layer4_outputs(1476) <= layer3_outputs(6617);
    layer4_outputs(1477) <= not(layer3_outputs(10081));
    layer4_outputs(1478) <= not(layer3_outputs(9770));
    layer4_outputs(1479) <= not((layer3_outputs(7186)) or (layer3_outputs(9454)));
    layer4_outputs(1480) <= layer3_outputs(5607);
    layer4_outputs(1481) <= (layer3_outputs(917)) or (layer3_outputs(4556));
    layer4_outputs(1482) <= not(layer3_outputs(8713));
    layer4_outputs(1483) <= not((layer3_outputs(3594)) xor (layer3_outputs(7922)));
    layer4_outputs(1484) <= not((layer3_outputs(9252)) and (layer3_outputs(1917)));
    layer4_outputs(1485) <= not((layer3_outputs(7473)) or (layer3_outputs(4037)));
    layer4_outputs(1486) <= (layer3_outputs(133)) xor (layer3_outputs(3236));
    layer4_outputs(1487) <= layer3_outputs(6136);
    layer4_outputs(1488) <= not(layer3_outputs(10081));
    layer4_outputs(1489) <= not(layer3_outputs(4525));
    layer4_outputs(1490) <= layer3_outputs(10109);
    layer4_outputs(1491) <= not(layer3_outputs(9202));
    layer4_outputs(1492) <= layer3_outputs(613);
    layer4_outputs(1493) <= not(layer3_outputs(7259));
    layer4_outputs(1494) <= layer3_outputs(5043);
    layer4_outputs(1495) <= (layer3_outputs(9246)) xor (layer3_outputs(8977));
    layer4_outputs(1496) <= not(layer3_outputs(8793));
    layer4_outputs(1497) <= (layer3_outputs(8862)) xor (layer3_outputs(3639));
    layer4_outputs(1498) <= layer3_outputs(3087);
    layer4_outputs(1499) <= (layer3_outputs(4749)) and not (layer3_outputs(9973));
    layer4_outputs(1500) <= not(layer3_outputs(2710));
    layer4_outputs(1501) <= '0';
    layer4_outputs(1502) <= not(layer3_outputs(4952)) or (layer3_outputs(4777));
    layer4_outputs(1503) <= layer3_outputs(5955);
    layer4_outputs(1504) <= not(layer3_outputs(6590));
    layer4_outputs(1505) <= layer3_outputs(1142);
    layer4_outputs(1506) <= (layer3_outputs(3554)) or (layer3_outputs(426));
    layer4_outputs(1507) <= layer3_outputs(8363);
    layer4_outputs(1508) <= not((layer3_outputs(27)) or (layer3_outputs(315)));
    layer4_outputs(1509) <= not(layer3_outputs(9703));
    layer4_outputs(1510) <= layer3_outputs(3442);
    layer4_outputs(1511) <= layer3_outputs(6642);
    layer4_outputs(1512) <= layer3_outputs(8091);
    layer4_outputs(1513) <= not(layer3_outputs(58)) or (layer3_outputs(7117));
    layer4_outputs(1514) <= not(layer3_outputs(8688)) or (layer3_outputs(2748));
    layer4_outputs(1515) <= not(layer3_outputs(6849));
    layer4_outputs(1516) <= not((layer3_outputs(4070)) or (layer3_outputs(8246)));
    layer4_outputs(1517) <= not(layer3_outputs(6831)) or (layer3_outputs(7250));
    layer4_outputs(1518) <= not(layer3_outputs(5730)) or (layer3_outputs(9420));
    layer4_outputs(1519) <= not(layer3_outputs(13)) or (layer3_outputs(2103));
    layer4_outputs(1520) <= layer3_outputs(5092);
    layer4_outputs(1521) <= not((layer3_outputs(6861)) xor (layer3_outputs(9694)));
    layer4_outputs(1522) <= (layer3_outputs(7488)) and not (layer3_outputs(7071));
    layer4_outputs(1523) <= not(layer3_outputs(8830));
    layer4_outputs(1524) <= not(layer3_outputs(3165)) or (layer3_outputs(9484));
    layer4_outputs(1525) <= layer3_outputs(3301);
    layer4_outputs(1526) <= layer3_outputs(8701);
    layer4_outputs(1527) <= not(layer3_outputs(3697));
    layer4_outputs(1528) <= (layer3_outputs(4591)) and not (layer3_outputs(2484));
    layer4_outputs(1529) <= not(layer3_outputs(4505));
    layer4_outputs(1530) <= layer3_outputs(327);
    layer4_outputs(1531) <= not((layer3_outputs(1260)) and (layer3_outputs(6250)));
    layer4_outputs(1532) <= not((layer3_outputs(5905)) and (layer3_outputs(9369)));
    layer4_outputs(1533) <= not(layer3_outputs(5691));
    layer4_outputs(1534) <= not((layer3_outputs(2082)) or (layer3_outputs(7703)));
    layer4_outputs(1535) <= layer3_outputs(9539);
    layer4_outputs(1536) <= (layer3_outputs(1197)) and not (layer3_outputs(2232));
    layer4_outputs(1537) <= (layer3_outputs(2716)) or (layer3_outputs(3910));
    layer4_outputs(1538) <= layer3_outputs(6680);
    layer4_outputs(1539) <= not(layer3_outputs(3179));
    layer4_outputs(1540) <= not((layer3_outputs(10017)) or (layer3_outputs(7636)));
    layer4_outputs(1541) <= (layer3_outputs(5856)) or (layer3_outputs(5758));
    layer4_outputs(1542) <= layer3_outputs(2618);
    layer4_outputs(1543) <= not((layer3_outputs(2159)) xor (layer3_outputs(3920)));
    layer4_outputs(1544) <= not((layer3_outputs(1874)) xor (layer3_outputs(10183)));
    layer4_outputs(1545) <= (layer3_outputs(7011)) and not (layer3_outputs(2923));
    layer4_outputs(1546) <= not((layer3_outputs(4377)) xor (layer3_outputs(8933)));
    layer4_outputs(1547) <= not((layer3_outputs(4597)) and (layer3_outputs(3963)));
    layer4_outputs(1548) <= (layer3_outputs(7786)) xor (layer3_outputs(2519));
    layer4_outputs(1549) <= not(layer3_outputs(5706));
    layer4_outputs(1550) <= not((layer3_outputs(9906)) or (layer3_outputs(1591)));
    layer4_outputs(1551) <= (layer3_outputs(7641)) xor (layer3_outputs(4317));
    layer4_outputs(1552) <= (layer3_outputs(5079)) and (layer3_outputs(5030));
    layer4_outputs(1553) <= not(layer3_outputs(9130));
    layer4_outputs(1554) <= not((layer3_outputs(2497)) or (layer3_outputs(4587)));
    layer4_outputs(1555) <= not(layer3_outputs(6427));
    layer4_outputs(1556) <= not((layer3_outputs(1552)) xor (layer3_outputs(2778)));
    layer4_outputs(1557) <= not(layer3_outputs(5700));
    layer4_outputs(1558) <= not((layer3_outputs(8219)) xor (layer3_outputs(5208)));
    layer4_outputs(1559) <= layer3_outputs(6074);
    layer4_outputs(1560) <= not(layer3_outputs(4390)) or (layer3_outputs(3242));
    layer4_outputs(1561) <= not(layer3_outputs(3884));
    layer4_outputs(1562) <= layer3_outputs(7606);
    layer4_outputs(1563) <= not(layer3_outputs(7429));
    layer4_outputs(1564) <= not(layer3_outputs(6539));
    layer4_outputs(1565) <= (layer3_outputs(5992)) or (layer3_outputs(8872));
    layer4_outputs(1566) <= not((layer3_outputs(8942)) xor (layer3_outputs(514)));
    layer4_outputs(1567) <= not((layer3_outputs(7938)) xor (layer3_outputs(3594)));
    layer4_outputs(1568) <= not((layer3_outputs(6649)) and (layer3_outputs(8618)));
    layer4_outputs(1569) <= not(layer3_outputs(7031));
    layer4_outputs(1570) <= layer3_outputs(829);
    layer4_outputs(1571) <= layer3_outputs(556);
    layer4_outputs(1572) <= not((layer3_outputs(7220)) xor (layer3_outputs(1541)));
    layer4_outputs(1573) <= layer3_outputs(5438);
    layer4_outputs(1574) <= not(layer3_outputs(1368)) or (layer3_outputs(1262));
    layer4_outputs(1575) <= layer3_outputs(2757);
    layer4_outputs(1576) <= (layer3_outputs(9798)) xor (layer3_outputs(7395));
    layer4_outputs(1577) <= layer3_outputs(4717);
    layer4_outputs(1578) <= not(layer3_outputs(8313));
    layer4_outputs(1579) <= not(layer3_outputs(3193));
    layer4_outputs(1580) <= (layer3_outputs(9948)) and (layer3_outputs(2539));
    layer4_outputs(1581) <= layer3_outputs(1650);
    layer4_outputs(1582) <= not(layer3_outputs(6948));
    layer4_outputs(1583) <= '0';
    layer4_outputs(1584) <= (layer3_outputs(6668)) and not (layer3_outputs(10120));
    layer4_outputs(1585) <= not(layer3_outputs(9394));
    layer4_outputs(1586) <= not((layer3_outputs(6177)) xor (layer3_outputs(3113)));
    layer4_outputs(1587) <= layer3_outputs(8824);
    layer4_outputs(1588) <= not((layer3_outputs(1862)) or (layer3_outputs(4414)));
    layer4_outputs(1589) <= not((layer3_outputs(4430)) or (layer3_outputs(7531)));
    layer4_outputs(1590) <= layer3_outputs(5346);
    layer4_outputs(1591) <= layer3_outputs(9388);
    layer4_outputs(1592) <= not((layer3_outputs(5493)) or (layer3_outputs(785)));
    layer4_outputs(1593) <= layer3_outputs(1312);
    layer4_outputs(1594) <= layer3_outputs(2374);
    layer4_outputs(1595) <= not(layer3_outputs(4217));
    layer4_outputs(1596) <= not(layer3_outputs(9309));
    layer4_outputs(1597) <= (layer3_outputs(9489)) and (layer3_outputs(2686));
    layer4_outputs(1598) <= not(layer3_outputs(6601));
    layer4_outputs(1599) <= not(layer3_outputs(4914));
    layer4_outputs(1600) <= not(layer3_outputs(5508));
    layer4_outputs(1601) <= (layer3_outputs(7388)) and (layer3_outputs(4058));
    layer4_outputs(1602) <= not(layer3_outputs(9950));
    layer4_outputs(1603) <= not((layer3_outputs(7774)) xor (layer3_outputs(7281)));
    layer4_outputs(1604) <= layer3_outputs(10027);
    layer4_outputs(1605) <= not(layer3_outputs(7595));
    layer4_outputs(1606) <= (layer3_outputs(3392)) and not (layer3_outputs(4105));
    layer4_outputs(1607) <= not(layer3_outputs(4257)) or (layer3_outputs(7980));
    layer4_outputs(1608) <= layer3_outputs(8533);
    layer4_outputs(1609) <= not((layer3_outputs(6650)) xor (layer3_outputs(7642)));
    layer4_outputs(1610) <= (layer3_outputs(2771)) or (layer3_outputs(8570));
    layer4_outputs(1611) <= (layer3_outputs(5747)) xor (layer3_outputs(7323));
    layer4_outputs(1612) <= not((layer3_outputs(4170)) xor (layer3_outputs(7054)));
    layer4_outputs(1613) <= layer3_outputs(56);
    layer4_outputs(1614) <= (layer3_outputs(2257)) and not (layer3_outputs(4427));
    layer4_outputs(1615) <= layer3_outputs(5209);
    layer4_outputs(1616) <= not(layer3_outputs(9683));
    layer4_outputs(1617) <= layer3_outputs(1684);
    layer4_outputs(1618) <= not((layer3_outputs(4757)) and (layer3_outputs(9413)));
    layer4_outputs(1619) <= not(layer3_outputs(960));
    layer4_outputs(1620) <= (layer3_outputs(161)) and not (layer3_outputs(1007));
    layer4_outputs(1621) <= not(layer3_outputs(4262));
    layer4_outputs(1622) <= (layer3_outputs(4530)) xor (layer3_outputs(5782));
    layer4_outputs(1623) <= not(layer3_outputs(6487));
    layer4_outputs(1624) <= layer3_outputs(8657);
    layer4_outputs(1625) <= not((layer3_outputs(9845)) or (layer3_outputs(1261)));
    layer4_outputs(1626) <= (layer3_outputs(8738)) or (layer3_outputs(10031));
    layer4_outputs(1627) <= layer3_outputs(3143);
    layer4_outputs(1628) <= (layer3_outputs(88)) and (layer3_outputs(3588));
    layer4_outputs(1629) <= not(layer3_outputs(3765));
    layer4_outputs(1630) <= not(layer3_outputs(2392)) or (layer3_outputs(9007));
    layer4_outputs(1631) <= not(layer3_outputs(4106));
    layer4_outputs(1632) <= not(layer3_outputs(5992));
    layer4_outputs(1633) <= not(layer3_outputs(3097));
    layer4_outputs(1634) <= not(layer3_outputs(819));
    layer4_outputs(1635) <= not((layer3_outputs(3194)) and (layer3_outputs(1702)));
    layer4_outputs(1636) <= not(layer3_outputs(1146));
    layer4_outputs(1637) <= not(layer3_outputs(4568));
    layer4_outputs(1638) <= layer3_outputs(1692);
    layer4_outputs(1639) <= not(layer3_outputs(9008));
    layer4_outputs(1640) <= not(layer3_outputs(3972));
    layer4_outputs(1641) <= not((layer3_outputs(3925)) xor (layer3_outputs(192)));
    layer4_outputs(1642) <= not((layer3_outputs(369)) xor (layer3_outputs(2390)));
    layer4_outputs(1643) <= not(layer3_outputs(1506));
    layer4_outputs(1644) <= not(layer3_outputs(6154)) or (layer3_outputs(1106));
    layer4_outputs(1645) <= not(layer3_outputs(388)) or (layer3_outputs(8758));
    layer4_outputs(1646) <= not((layer3_outputs(3581)) or (layer3_outputs(9818)));
    layer4_outputs(1647) <= layer3_outputs(3552);
    layer4_outputs(1648) <= not(layer3_outputs(9226));
    layer4_outputs(1649) <= layer3_outputs(4473);
    layer4_outputs(1650) <= (layer3_outputs(1081)) and (layer3_outputs(43));
    layer4_outputs(1651) <= layer3_outputs(61);
    layer4_outputs(1652) <= (layer3_outputs(6877)) and (layer3_outputs(4078));
    layer4_outputs(1653) <= not(layer3_outputs(2293));
    layer4_outputs(1654) <= layer3_outputs(6367);
    layer4_outputs(1655) <= (layer3_outputs(3022)) xor (layer3_outputs(6209));
    layer4_outputs(1656) <= not(layer3_outputs(3890));
    layer4_outputs(1657) <= not(layer3_outputs(728));
    layer4_outputs(1658) <= (layer3_outputs(1297)) and not (layer3_outputs(6540));
    layer4_outputs(1659) <= not(layer3_outputs(1709));
    layer4_outputs(1660) <= not(layer3_outputs(526)) or (layer3_outputs(1312));
    layer4_outputs(1661) <= not(layer3_outputs(2100)) or (layer3_outputs(361));
    layer4_outputs(1662) <= not(layer3_outputs(7929));
    layer4_outputs(1663) <= layer3_outputs(8428);
    layer4_outputs(1664) <= not(layer3_outputs(6981));
    layer4_outputs(1665) <= layer3_outputs(6579);
    layer4_outputs(1666) <= layer3_outputs(7062);
    layer4_outputs(1667) <= layer3_outputs(186);
    layer4_outputs(1668) <= not(layer3_outputs(6173));
    layer4_outputs(1669) <= layer3_outputs(3713);
    layer4_outputs(1670) <= (layer3_outputs(9337)) xor (layer3_outputs(5306));
    layer4_outputs(1671) <= not(layer3_outputs(7005)) or (layer3_outputs(4391));
    layer4_outputs(1672) <= not(layer3_outputs(8554));
    layer4_outputs(1673) <= layer3_outputs(4919);
    layer4_outputs(1674) <= layer3_outputs(6745);
    layer4_outputs(1675) <= (layer3_outputs(3844)) xor (layer3_outputs(8390));
    layer4_outputs(1676) <= not(layer3_outputs(9520));
    layer4_outputs(1677) <= layer3_outputs(7963);
    layer4_outputs(1678) <= (layer3_outputs(4956)) xor (layer3_outputs(4401));
    layer4_outputs(1679) <= not(layer3_outputs(8129));
    layer4_outputs(1680) <= not((layer3_outputs(3474)) xor (layer3_outputs(9254)));
    layer4_outputs(1681) <= layer3_outputs(4756);
    layer4_outputs(1682) <= not(layer3_outputs(7588));
    layer4_outputs(1683) <= not(layer3_outputs(5106));
    layer4_outputs(1684) <= layer3_outputs(5902);
    layer4_outputs(1685) <= layer3_outputs(1296);
    layer4_outputs(1686) <= not(layer3_outputs(7607));
    layer4_outputs(1687) <= layer3_outputs(6785);
    layer4_outputs(1688) <= not((layer3_outputs(7577)) xor (layer3_outputs(5524)));
    layer4_outputs(1689) <= layer3_outputs(9528);
    layer4_outputs(1690) <= not(layer3_outputs(8263));
    layer4_outputs(1691) <= layer3_outputs(1922);
    layer4_outputs(1692) <= not((layer3_outputs(3324)) xor (layer3_outputs(4429)));
    layer4_outputs(1693) <= layer3_outputs(1498);
    layer4_outputs(1694) <= not(layer3_outputs(8345));
    layer4_outputs(1695) <= not((layer3_outputs(8773)) xor (layer3_outputs(54)));
    layer4_outputs(1696) <= (layer3_outputs(1562)) or (layer3_outputs(1104));
    layer4_outputs(1697) <= (layer3_outputs(2833)) xor (layer3_outputs(701));
    layer4_outputs(1698) <= layer3_outputs(2413);
    layer4_outputs(1699) <= not(layer3_outputs(9228));
    layer4_outputs(1700) <= layer3_outputs(8844);
    layer4_outputs(1701) <= layer3_outputs(6085);
    layer4_outputs(1702) <= layer3_outputs(4251);
    layer4_outputs(1703) <= not((layer3_outputs(3700)) or (layer3_outputs(9460)));
    layer4_outputs(1704) <= layer3_outputs(7408);
    layer4_outputs(1705) <= layer3_outputs(7602);
    layer4_outputs(1706) <= (layer3_outputs(8490)) or (layer3_outputs(6418));
    layer4_outputs(1707) <= layer3_outputs(2224);
    layer4_outputs(1708) <= (layer3_outputs(3147)) and not (layer3_outputs(1880));
    layer4_outputs(1709) <= layer3_outputs(5806);
    layer4_outputs(1710) <= layer3_outputs(4633);
    layer4_outputs(1711) <= not(layer3_outputs(7142));
    layer4_outputs(1712) <= (layer3_outputs(6684)) or (layer3_outputs(571));
    layer4_outputs(1713) <= (layer3_outputs(9454)) or (layer3_outputs(5126));
    layer4_outputs(1714) <= not((layer3_outputs(1311)) and (layer3_outputs(6114)));
    layer4_outputs(1715) <= layer3_outputs(3823);
    layer4_outputs(1716) <= not(layer3_outputs(5231));
    layer4_outputs(1717) <= not(layer3_outputs(6703));
    layer4_outputs(1718) <= not((layer3_outputs(323)) and (layer3_outputs(5708)));
    layer4_outputs(1719) <= not(layer3_outputs(9105));
    layer4_outputs(1720) <= (layer3_outputs(8022)) and not (layer3_outputs(5859));
    layer4_outputs(1721) <= (layer3_outputs(3246)) and not (layer3_outputs(7634));
    layer4_outputs(1722) <= not((layer3_outputs(4696)) xor (layer3_outputs(433)));
    layer4_outputs(1723) <= not(layer3_outputs(2563));
    layer4_outputs(1724) <= (layer3_outputs(3312)) xor (layer3_outputs(4185));
    layer4_outputs(1725) <= not(layer3_outputs(6490));
    layer4_outputs(1726) <= (layer3_outputs(2930)) xor (layer3_outputs(2814));
    layer4_outputs(1727) <= layer3_outputs(9824);
    layer4_outputs(1728) <= layer3_outputs(8662);
    layer4_outputs(1729) <= layer3_outputs(2999);
    layer4_outputs(1730) <= not(layer3_outputs(7174));
    layer4_outputs(1731) <= layer3_outputs(2500);
    layer4_outputs(1732) <= (layer3_outputs(6501)) and (layer3_outputs(4387));
    layer4_outputs(1733) <= layer3_outputs(959);
    layer4_outputs(1734) <= (layer3_outputs(10140)) and not (layer3_outputs(8301));
    layer4_outputs(1735) <= layer3_outputs(6890);
    layer4_outputs(1736) <= (layer3_outputs(8527)) and not (layer3_outputs(678));
    layer4_outputs(1737) <= (layer3_outputs(1668)) and (layer3_outputs(1675));
    layer4_outputs(1738) <= layer3_outputs(9685);
    layer4_outputs(1739) <= not(layer3_outputs(5312)) or (layer3_outputs(6388));
    layer4_outputs(1740) <= not(layer3_outputs(234));
    layer4_outputs(1741) <= not((layer3_outputs(6315)) xor (layer3_outputs(1353)));
    layer4_outputs(1742) <= not((layer3_outputs(1809)) or (layer3_outputs(814)));
    layer4_outputs(1743) <= not(layer3_outputs(2191));
    layer4_outputs(1744) <= (layer3_outputs(5468)) and not (layer3_outputs(7448));
    layer4_outputs(1745) <= layer3_outputs(4848);
    layer4_outputs(1746) <= not((layer3_outputs(164)) or (layer3_outputs(2559)));
    layer4_outputs(1747) <= (layer3_outputs(9455)) and (layer3_outputs(8945));
    layer4_outputs(1748) <= not((layer3_outputs(4821)) and (layer3_outputs(8614)));
    layer4_outputs(1749) <= (layer3_outputs(5110)) or (layer3_outputs(1566));
    layer4_outputs(1750) <= not((layer3_outputs(2676)) or (layer3_outputs(9514)));
    layer4_outputs(1751) <= not(layer3_outputs(3731)) or (layer3_outputs(4474));
    layer4_outputs(1752) <= not(layer3_outputs(6709));
    layer4_outputs(1753) <= layer3_outputs(10020);
    layer4_outputs(1754) <= not(layer3_outputs(2827));
    layer4_outputs(1755) <= not((layer3_outputs(1131)) xor (layer3_outputs(1897)));
    layer4_outputs(1756) <= (layer3_outputs(36)) xor (layer3_outputs(3976));
    layer4_outputs(1757) <= not((layer3_outputs(4529)) xor (layer3_outputs(4266)));
    layer4_outputs(1758) <= (layer3_outputs(2438)) and not (layer3_outputs(3986));
    layer4_outputs(1759) <= layer3_outputs(3720);
    layer4_outputs(1760) <= (layer3_outputs(8906)) and not (layer3_outputs(8273));
    layer4_outputs(1761) <= not((layer3_outputs(5092)) xor (layer3_outputs(4536)));
    layer4_outputs(1762) <= layer3_outputs(6864);
    layer4_outputs(1763) <= layer3_outputs(4957);
    layer4_outputs(1764) <= not(layer3_outputs(1316));
    layer4_outputs(1765) <= not((layer3_outputs(3763)) xor (layer3_outputs(3962)));
    layer4_outputs(1766) <= (layer3_outputs(738)) and (layer3_outputs(6463));
    layer4_outputs(1767) <= not(layer3_outputs(7480));
    layer4_outputs(1768) <= layer3_outputs(8450);
    layer4_outputs(1769) <= not(layer3_outputs(3750));
    layer4_outputs(1770) <= (layer3_outputs(5001)) and not (layer3_outputs(3771));
    layer4_outputs(1771) <= not(layer3_outputs(8646));
    layer4_outputs(1772) <= (layer3_outputs(5268)) or (layer3_outputs(442));
    layer4_outputs(1773) <= layer3_outputs(3521);
    layer4_outputs(1774) <= (layer3_outputs(7202)) and (layer3_outputs(8041));
    layer4_outputs(1775) <= not(layer3_outputs(8764));
    layer4_outputs(1776) <= (layer3_outputs(6862)) and (layer3_outputs(2931));
    layer4_outputs(1777) <= not(layer3_outputs(7360));
    layer4_outputs(1778) <= not(layer3_outputs(6555));
    layer4_outputs(1779) <= not(layer3_outputs(4906));
    layer4_outputs(1780) <= (layer3_outputs(8731)) and not (layer3_outputs(8937));
    layer4_outputs(1781) <= layer3_outputs(6073);
    layer4_outputs(1782) <= layer3_outputs(7310);
    layer4_outputs(1783) <= not(layer3_outputs(6821));
    layer4_outputs(1784) <= not(layer3_outputs(4481));
    layer4_outputs(1785) <= not((layer3_outputs(4466)) xor (layer3_outputs(2248)));
    layer4_outputs(1786) <= not(layer3_outputs(10147));
    layer4_outputs(1787) <= (layer3_outputs(8302)) and (layer3_outputs(2109));
    layer4_outputs(1788) <= (layer3_outputs(4652)) and not (layer3_outputs(4014));
    layer4_outputs(1789) <= not(layer3_outputs(5857));
    layer4_outputs(1790) <= layer3_outputs(7455);
    layer4_outputs(1791) <= not(layer3_outputs(173));
    layer4_outputs(1792) <= not(layer3_outputs(3057));
    layer4_outputs(1793) <= not(layer3_outputs(4946));
    layer4_outputs(1794) <= not((layer3_outputs(6082)) xor (layer3_outputs(3498)));
    layer4_outputs(1795) <= layer3_outputs(6977);
    layer4_outputs(1796) <= not(layer3_outputs(245)) or (layer3_outputs(521));
    layer4_outputs(1797) <= (layer3_outputs(4738)) or (layer3_outputs(579));
    layer4_outputs(1798) <= (layer3_outputs(9018)) and not (layer3_outputs(3677));
    layer4_outputs(1799) <= (layer3_outputs(7522)) and not (layer3_outputs(3724));
    layer4_outputs(1800) <= (layer3_outputs(4007)) xor (layer3_outputs(6704));
    layer4_outputs(1801) <= not(layer3_outputs(2349));
    layer4_outputs(1802) <= (layer3_outputs(593)) or (layer3_outputs(3939));
    layer4_outputs(1803) <= not((layer3_outputs(5614)) xor (layer3_outputs(6493)));
    layer4_outputs(1804) <= layer3_outputs(4486);
    layer4_outputs(1805) <= not(layer3_outputs(4994));
    layer4_outputs(1806) <= layer3_outputs(18);
    layer4_outputs(1807) <= (layer3_outputs(5703)) and not (layer3_outputs(8675));
    layer4_outputs(1808) <= layer3_outputs(3618);
    layer4_outputs(1809) <= not(layer3_outputs(8578));
    layer4_outputs(1810) <= (layer3_outputs(2208)) and not (layer3_outputs(2584));
    layer4_outputs(1811) <= not(layer3_outputs(6757)) or (layer3_outputs(31));
    layer4_outputs(1812) <= (layer3_outputs(6506)) xor (layer3_outputs(7042));
    layer4_outputs(1813) <= not((layer3_outputs(8732)) or (layer3_outputs(3545)));
    layer4_outputs(1814) <= (layer3_outputs(3985)) and (layer3_outputs(8197));
    layer4_outputs(1815) <= not(layer3_outputs(6110));
    layer4_outputs(1816) <= not(layer3_outputs(7331));
    layer4_outputs(1817) <= not(layer3_outputs(7541));
    layer4_outputs(1818) <= (layer3_outputs(1296)) and not (layer3_outputs(7838));
    layer4_outputs(1819) <= not(layer3_outputs(653)) or (layer3_outputs(10180));
    layer4_outputs(1820) <= not(layer3_outputs(7968));
    layer4_outputs(1821) <= layer3_outputs(6214);
    layer4_outputs(1822) <= (layer3_outputs(7200)) and not (layer3_outputs(4358));
    layer4_outputs(1823) <= (layer3_outputs(5604)) xor (layer3_outputs(3932));
    layer4_outputs(1824) <= not(layer3_outputs(4255));
    layer4_outputs(1825) <= not(layer3_outputs(7757));
    layer4_outputs(1826) <= (layer3_outputs(96)) xor (layer3_outputs(6791));
    layer4_outputs(1827) <= layer3_outputs(140);
    layer4_outputs(1828) <= not((layer3_outputs(3394)) xor (layer3_outputs(9680)));
    layer4_outputs(1829) <= (layer3_outputs(325)) xor (layer3_outputs(7605));
    layer4_outputs(1830) <= (layer3_outputs(3673)) and not (layer3_outputs(5174));
    layer4_outputs(1831) <= (layer3_outputs(8428)) and (layer3_outputs(5677));
    layer4_outputs(1832) <= (layer3_outputs(1467)) xor (layer3_outputs(1943));
    layer4_outputs(1833) <= not((layer3_outputs(5534)) and (layer3_outputs(7906)));
    layer4_outputs(1834) <= layer3_outputs(9470);
    layer4_outputs(1835) <= not(layer3_outputs(5542));
    layer4_outputs(1836) <= layer3_outputs(7759);
    layer4_outputs(1837) <= not((layer3_outputs(5960)) xor (layer3_outputs(4486)));
    layer4_outputs(1838) <= not(layer3_outputs(1525)) or (layer3_outputs(7269));
    layer4_outputs(1839) <= layer3_outputs(1987);
    layer4_outputs(1840) <= layer3_outputs(7054);
    layer4_outputs(1841) <= layer3_outputs(2085);
    layer4_outputs(1842) <= not(layer3_outputs(154));
    layer4_outputs(1843) <= (layer3_outputs(9750)) and (layer3_outputs(3730));
    layer4_outputs(1844) <= not(layer3_outputs(1882)) or (layer3_outputs(3803));
    layer4_outputs(1845) <= not(layer3_outputs(3292));
    layer4_outputs(1846) <= not((layer3_outputs(8600)) xor (layer3_outputs(5457)));
    layer4_outputs(1847) <= not(layer3_outputs(5660)) or (layer3_outputs(3206));
    layer4_outputs(1848) <= (layer3_outputs(1340)) and not (layer3_outputs(5835));
    layer4_outputs(1849) <= not((layer3_outputs(3759)) and (layer3_outputs(2116)));
    layer4_outputs(1850) <= layer3_outputs(1588);
    layer4_outputs(1851) <= (layer3_outputs(954)) xor (layer3_outputs(4449));
    layer4_outputs(1852) <= layer3_outputs(6494);
    layer4_outputs(1853) <= layer3_outputs(6627);
    layer4_outputs(1854) <= not(layer3_outputs(6892));
    layer4_outputs(1855) <= not(layer3_outputs(398));
    layer4_outputs(1856) <= (layer3_outputs(4152)) or (layer3_outputs(9087));
    layer4_outputs(1857) <= not((layer3_outputs(7891)) xor (layer3_outputs(5838)));
    layer4_outputs(1858) <= not(layer3_outputs(7337));
    layer4_outputs(1859) <= layer3_outputs(9618);
    layer4_outputs(1860) <= not((layer3_outputs(2266)) xor (layer3_outputs(9481)));
    layer4_outputs(1861) <= not(layer3_outputs(5296));
    layer4_outputs(1862) <= (layer3_outputs(5111)) and (layer3_outputs(2597));
    layer4_outputs(1863) <= not((layer3_outputs(2156)) xor (layer3_outputs(2857)));
    layer4_outputs(1864) <= not(layer3_outputs(677)) or (layer3_outputs(8294));
    layer4_outputs(1865) <= not((layer3_outputs(2625)) xor (layer3_outputs(6721)));
    layer4_outputs(1866) <= layer3_outputs(4277);
    layer4_outputs(1867) <= (layer3_outputs(2453)) or (layer3_outputs(3067));
    layer4_outputs(1868) <= layer3_outputs(8210);
    layer4_outputs(1869) <= not(layer3_outputs(7021));
    layer4_outputs(1870) <= layer3_outputs(3245);
    layer4_outputs(1871) <= not(layer3_outputs(1165));
    layer4_outputs(1872) <= not(layer3_outputs(6536));
    layer4_outputs(1873) <= not(layer3_outputs(2090));
    layer4_outputs(1874) <= not(layer3_outputs(2941));
    layer4_outputs(1875) <= layer3_outputs(3795);
    layer4_outputs(1876) <= layer3_outputs(8049);
    layer4_outputs(1877) <= not((layer3_outputs(182)) and (layer3_outputs(7704)));
    layer4_outputs(1878) <= not(layer3_outputs(8053));
    layer4_outputs(1879) <= layer3_outputs(4172);
    layer4_outputs(1880) <= not((layer3_outputs(8512)) xor (layer3_outputs(9867)));
    layer4_outputs(1881) <= (layer3_outputs(9261)) and (layer3_outputs(2369));
    layer4_outputs(1882) <= layer3_outputs(5476);
    layer4_outputs(1883) <= not((layer3_outputs(7557)) or (layer3_outputs(7844)));
    layer4_outputs(1884) <= layer3_outputs(5638);
    layer4_outputs(1885) <= not(layer3_outputs(8954));
    layer4_outputs(1886) <= not((layer3_outputs(165)) and (layer3_outputs(3602)));
    layer4_outputs(1887) <= not((layer3_outputs(7183)) or (layer3_outputs(2489)));
    layer4_outputs(1888) <= not(layer3_outputs(4845));
    layer4_outputs(1889) <= layer3_outputs(6365);
    layer4_outputs(1890) <= (layer3_outputs(3581)) and (layer3_outputs(7914));
    layer4_outputs(1891) <= layer3_outputs(6300);
    layer4_outputs(1892) <= '0';
    layer4_outputs(1893) <= not(layer3_outputs(463));
    layer4_outputs(1894) <= not((layer3_outputs(3457)) xor (layer3_outputs(279)));
    layer4_outputs(1895) <= not(layer3_outputs(2059));
    layer4_outputs(1896) <= layer3_outputs(4697);
    layer4_outputs(1897) <= not((layer3_outputs(4667)) xor (layer3_outputs(420)));
    layer4_outputs(1898) <= (layer3_outputs(2443)) xor (layer3_outputs(1499));
    layer4_outputs(1899) <= not(layer3_outputs(4876));
    layer4_outputs(1900) <= not(layer3_outputs(9239));
    layer4_outputs(1901) <= not((layer3_outputs(7454)) xor (layer3_outputs(10222)));
    layer4_outputs(1902) <= (layer3_outputs(1805)) or (layer3_outputs(9650));
    layer4_outputs(1903) <= not(layer3_outputs(4925));
    layer4_outputs(1904) <= (layer3_outputs(8191)) and (layer3_outputs(6907));
    layer4_outputs(1905) <= not((layer3_outputs(3623)) xor (layer3_outputs(6753)));
    layer4_outputs(1906) <= not(layer3_outputs(8279));
    layer4_outputs(1907) <= layer3_outputs(2871);
    layer4_outputs(1908) <= not(layer3_outputs(6471));
    layer4_outputs(1909) <= (layer3_outputs(29)) or (layer3_outputs(7814));
    layer4_outputs(1910) <= (layer3_outputs(390)) xor (layer3_outputs(2594));
    layer4_outputs(1911) <= (layer3_outputs(4693)) or (layer3_outputs(3883));
    layer4_outputs(1912) <= not((layer3_outputs(5206)) and (layer3_outputs(41)));
    layer4_outputs(1913) <= not(layer3_outputs(9519));
    layer4_outputs(1914) <= not(layer3_outputs(5385));
    layer4_outputs(1915) <= (layer3_outputs(3265)) xor (layer3_outputs(2809));
    layer4_outputs(1916) <= layer3_outputs(1115);
    layer4_outputs(1917) <= not((layer3_outputs(5155)) xor (layer3_outputs(9716)));
    layer4_outputs(1918) <= not(layer3_outputs(7025));
    layer4_outputs(1919) <= not(layer3_outputs(9840));
    layer4_outputs(1920) <= (layer3_outputs(8736)) xor (layer3_outputs(3601));
    layer4_outputs(1921) <= layer3_outputs(5579);
    layer4_outputs(1922) <= not(layer3_outputs(7560));
    layer4_outputs(1923) <= (layer3_outputs(4009)) and not (layer3_outputs(3516));
    layer4_outputs(1924) <= '0';
    layer4_outputs(1925) <= layer3_outputs(2236);
    layer4_outputs(1926) <= not(layer3_outputs(19));
    layer4_outputs(1927) <= not((layer3_outputs(9092)) xor (layer3_outputs(8213)));
    layer4_outputs(1928) <= not(layer3_outputs(794)) or (layer3_outputs(3598));
    layer4_outputs(1929) <= (layer3_outputs(8471)) xor (layer3_outputs(3845));
    layer4_outputs(1930) <= not(layer3_outputs(2210));
    layer4_outputs(1931) <= layer3_outputs(69);
    layer4_outputs(1932) <= '1';
    layer4_outputs(1933) <= layer3_outputs(9817);
    layer4_outputs(1934) <= not(layer3_outputs(910)) or (layer3_outputs(4487));
    layer4_outputs(1935) <= layer3_outputs(7447);
    layer4_outputs(1936) <= layer3_outputs(2392);
    layer4_outputs(1937) <= (layer3_outputs(3274)) xor (layer3_outputs(2924));
    layer4_outputs(1938) <= not(layer3_outputs(2072));
    layer4_outputs(1939) <= layer3_outputs(4843);
    layer4_outputs(1940) <= not(layer3_outputs(7386));
    layer4_outputs(1941) <= (layer3_outputs(3981)) and not (layer3_outputs(9662));
    layer4_outputs(1942) <= (layer3_outputs(3095)) xor (layer3_outputs(7211));
    layer4_outputs(1943) <= layer3_outputs(9889);
    layer4_outputs(1944) <= not(layer3_outputs(6124));
    layer4_outputs(1945) <= layer3_outputs(5040);
    layer4_outputs(1946) <= layer3_outputs(6240);
    layer4_outputs(1947) <= not(layer3_outputs(5056));
    layer4_outputs(1948) <= (layer3_outputs(7847)) and not (layer3_outputs(2973));
    layer4_outputs(1949) <= not(layer3_outputs(5188)) or (layer3_outputs(5488));
    layer4_outputs(1950) <= (layer3_outputs(9149)) and not (layer3_outputs(8007));
    layer4_outputs(1951) <= (layer3_outputs(1335)) or (layer3_outputs(7618));
    layer4_outputs(1952) <= layer3_outputs(2185);
    layer4_outputs(1953) <= not((layer3_outputs(9556)) or (layer3_outputs(2298)));
    layer4_outputs(1954) <= not(layer3_outputs(9004)) or (layer3_outputs(9155));
    layer4_outputs(1955) <= not(layer3_outputs(7244));
    layer4_outputs(1956) <= not((layer3_outputs(9905)) and (layer3_outputs(1619)));
    layer4_outputs(1957) <= not(layer3_outputs(998)) or (layer3_outputs(1306));
    layer4_outputs(1958) <= not(layer3_outputs(2881));
    layer4_outputs(1959) <= layer3_outputs(7515);
    layer4_outputs(1960) <= not(layer3_outputs(7127));
    layer4_outputs(1961) <= not((layer3_outputs(4413)) xor (layer3_outputs(7020)));
    layer4_outputs(1962) <= not(layer3_outputs(6004));
    layer4_outputs(1963) <= layer3_outputs(161);
    layer4_outputs(1964) <= not((layer3_outputs(2865)) and (layer3_outputs(9625)));
    layer4_outputs(1965) <= not(layer3_outputs(8821));
    layer4_outputs(1966) <= (layer3_outputs(3035)) and not (layer3_outputs(287));
    layer4_outputs(1967) <= layer3_outputs(5692);
    layer4_outputs(1968) <= (layer3_outputs(1929)) and not (layer3_outputs(6426));
    layer4_outputs(1969) <= not((layer3_outputs(692)) and (layer3_outputs(3816)));
    layer4_outputs(1970) <= (layer3_outputs(8969)) and (layer3_outputs(7381));
    layer4_outputs(1971) <= layer3_outputs(6646);
    layer4_outputs(1972) <= (layer3_outputs(4463)) and (layer3_outputs(5571));
    layer4_outputs(1973) <= not(layer3_outputs(4258));
    layer4_outputs(1974) <= not(layer3_outputs(3313));
    layer4_outputs(1975) <= layer3_outputs(6268);
    layer4_outputs(1976) <= not(layer3_outputs(4553)) or (layer3_outputs(1561));
    layer4_outputs(1977) <= not((layer3_outputs(2074)) xor (layer3_outputs(5267)));
    layer4_outputs(1978) <= layer3_outputs(6143);
    layer4_outputs(1979) <= not(layer3_outputs(3735)) or (layer3_outputs(5093));
    layer4_outputs(1980) <= not((layer3_outputs(6955)) or (layer3_outputs(6139)));
    layer4_outputs(1981) <= (layer3_outputs(1989)) and (layer3_outputs(9238));
    layer4_outputs(1982) <= (layer3_outputs(5615)) xor (layer3_outputs(7840));
    layer4_outputs(1983) <= layer3_outputs(7178);
    layer4_outputs(1984) <= not(layer3_outputs(5659));
    layer4_outputs(1985) <= (layer3_outputs(5485)) xor (layer3_outputs(1491));
    layer4_outputs(1986) <= not((layer3_outputs(3391)) and (layer3_outputs(3647)));
    layer4_outputs(1987) <= (layer3_outputs(8482)) or (layer3_outputs(4655));
    layer4_outputs(1988) <= not(layer3_outputs(2029));
    layer4_outputs(1989) <= not(layer3_outputs(9982));
    layer4_outputs(1990) <= layer3_outputs(7544);
    layer4_outputs(1991) <= not(layer3_outputs(7004));
    layer4_outputs(1992) <= (layer3_outputs(4462)) and not (layer3_outputs(9500));
    layer4_outputs(1993) <= layer3_outputs(5217);
    layer4_outputs(1994) <= not(layer3_outputs(540));
    layer4_outputs(1995) <= layer3_outputs(2708);
    layer4_outputs(1996) <= layer3_outputs(9194);
    layer4_outputs(1997) <= layer3_outputs(5171);
    layer4_outputs(1998) <= not(layer3_outputs(7760));
    layer4_outputs(1999) <= layer3_outputs(1966);
    layer4_outputs(2000) <= layer3_outputs(76);
    layer4_outputs(2001) <= layer3_outputs(7532);
    layer4_outputs(2002) <= not(layer3_outputs(1209));
    layer4_outputs(2003) <= not(layer3_outputs(972)) or (layer3_outputs(4695));
    layer4_outputs(2004) <= (layer3_outputs(49)) or (layer3_outputs(2425));
    layer4_outputs(2005) <= not(layer3_outputs(5704));
    layer4_outputs(2006) <= layer3_outputs(3014);
    layer4_outputs(2007) <= (layer3_outputs(1463)) and (layer3_outputs(139));
    layer4_outputs(2008) <= not((layer3_outputs(5068)) and (layer3_outputs(5182)));
    layer4_outputs(2009) <= layer3_outputs(7431);
    layer4_outputs(2010) <= (layer3_outputs(4026)) xor (layer3_outputs(723));
    layer4_outputs(2011) <= (layer3_outputs(2201)) and not (layer3_outputs(1554));
    layer4_outputs(2012) <= layer3_outputs(7355);
    layer4_outputs(2013) <= not((layer3_outputs(6144)) xor (layer3_outputs(4115)));
    layer4_outputs(2014) <= not((layer3_outputs(5309)) or (layer3_outputs(20)));
    layer4_outputs(2015) <= not((layer3_outputs(4115)) xor (layer3_outputs(8797)));
    layer4_outputs(2016) <= (layer3_outputs(5884)) and not (layer3_outputs(3074));
    layer4_outputs(2017) <= not((layer3_outputs(8733)) or (layer3_outputs(6323)));
    layer4_outputs(2018) <= layer3_outputs(8178);
    layer4_outputs(2019) <= layer3_outputs(4321);
    layer4_outputs(2020) <= (layer3_outputs(1403)) and not (layer3_outputs(2991));
    layer4_outputs(2021) <= not(layer3_outputs(929));
    layer4_outputs(2022) <= not((layer3_outputs(8755)) xor (layer3_outputs(9274)));
    layer4_outputs(2023) <= layer3_outputs(7677);
    layer4_outputs(2024) <= not(layer3_outputs(2324));
    layer4_outputs(2025) <= not((layer3_outputs(6685)) and (layer3_outputs(537)));
    layer4_outputs(2026) <= (layer3_outputs(1787)) or (layer3_outputs(4705));
    layer4_outputs(2027) <= layer3_outputs(2713);
    layer4_outputs(2028) <= not((layer3_outputs(9927)) xor (layer3_outputs(37)));
    layer4_outputs(2029) <= (layer3_outputs(8912)) xor (layer3_outputs(3924));
    layer4_outputs(2030) <= not((layer3_outputs(4353)) xor (layer3_outputs(6412)));
    layer4_outputs(2031) <= not(layer3_outputs(1593));
    layer4_outputs(2032) <= not(layer3_outputs(2653));
    layer4_outputs(2033) <= (layer3_outputs(8338)) and not (layer3_outputs(2265));
    layer4_outputs(2034) <= layer3_outputs(2963);
    layer4_outputs(2035) <= layer3_outputs(3675);
    layer4_outputs(2036) <= (layer3_outputs(1443)) and not (layer3_outputs(8990));
    layer4_outputs(2037) <= layer3_outputs(9216);
    layer4_outputs(2038) <= not(layer3_outputs(9515));
    layer4_outputs(2039) <= not((layer3_outputs(1447)) xor (layer3_outputs(3246)));
    layer4_outputs(2040) <= not(layer3_outputs(7370));
    layer4_outputs(2041) <= (layer3_outputs(2812)) and (layer3_outputs(8509));
    layer4_outputs(2042) <= not(layer3_outputs(985));
    layer4_outputs(2043) <= (layer3_outputs(10121)) xor (layer3_outputs(8978));
    layer4_outputs(2044) <= layer3_outputs(5763);
    layer4_outputs(2045) <= (layer3_outputs(10136)) and not (layer3_outputs(6105));
    layer4_outputs(2046) <= layer3_outputs(5619);
    layer4_outputs(2047) <= not(layer3_outputs(2580)) or (layer3_outputs(1965));
    layer4_outputs(2048) <= (layer3_outputs(6347)) xor (layer3_outputs(890));
    layer4_outputs(2049) <= '0';
    layer4_outputs(2050) <= layer3_outputs(7257);
    layer4_outputs(2051) <= (layer3_outputs(10182)) xor (layer3_outputs(8973));
    layer4_outputs(2052) <= (layer3_outputs(3216)) or (layer3_outputs(2331));
    layer4_outputs(2053) <= layer3_outputs(1388);
    layer4_outputs(2054) <= not(layer3_outputs(7491));
    layer4_outputs(2055) <= layer3_outputs(9490);
    layer4_outputs(2056) <= not(layer3_outputs(9673));
    layer4_outputs(2057) <= not(layer3_outputs(5027));
    layer4_outputs(2058) <= (layer3_outputs(8188)) xor (layer3_outputs(4527));
    layer4_outputs(2059) <= layer3_outputs(4367);
    layer4_outputs(2060) <= not((layer3_outputs(1757)) or (layer3_outputs(9182)));
    layer4_outputs(2061) <= not((layer3_outputs(6386)) or (layer3_outputs(5934)));
    layer4_outputs(2062) <= not(layer3_outputs(2469));
    layer4_outputs(2063) <= not(layer3_outputs(3726));
    layer4_outputs(2064) <= (layer3_outputs(8451)) and (layer3_outputs(3517));
    layer4_outputs(2065) <= not(layer3_outputs(9790));
    layer4_outputs(2066) <= layer3_outputs(2114);
    layer4_outputs(2067) <= not((layer3_outputs(5022)) or (layer3_outputs(7324)));
    layer4_outputs(2068) <= (layer3_outputs(570)) and (layer3_outputs(7851));
    layer4_outputs(2069) <= not(layer3_outputs(4182));
    layer4_outputs(2070) <= layer3_outputs(3456);
    layer4_outputs(2071) <= not(layer3_outputs(3363));
    layer4_outputs(2072) <= layer3_outputs(719);
    layer4_outputs(2073) <= not(layer3_outputs(7295));
    layer4_outputs(2074) <= not((layer3_outputs(5389)) xor (layer3_outputs(2483)));
    layer4_outputs(2075) <= (layer3_outputs(8872)) and not (layer3_outputs(97));
    layer4_outputs(2076) <= not(layer3_outputs(2421));
    layer4_outputs(2077) <= layer3_outputs(1964);
    layer4_outputs(2078) <= not(layer3_outputs(9187));
    layer4_outputs(2079) <= not(layer3_outputs(9367));
    layer4_outputs(2080) <= (layer3_outputs(3709)) or (layer3_outputs(6690));
    layer4_outputs(2081) <= not((layer3_outputs(8702)) or (layer3_outputs(9057)));
    layer4_outputs(2082) <= (layer3_outputs(4220)) and not (layer3_outputs(9943));
    layer4_outputs(2083) <= layer3_outputs(5940);
    layer4_outputs(2084) <= not((layer3_outputs(2445)) or (layer3_outputs(4779)));
    layer4_outputs(2085) <= (layer3_outputs(8838)) and not (layer3_outputs(446));
    layer4_outputs(2086) <= layer3_outputs(7612);
    layer4_outputs(2087) <= not(layer3_outputs(8850));
    layer4_outputs(2088) <= layer3_outputs(5138);
    layer4_outputs(2089) <= not(layer3_outputs(4955));
    layer4_outputs(2090) <= not(layer3_outputs(1405));
    layer4_outputs(2091) <= not(layer3_outputs(1533));
    layer4_outputs(2092) <= (layer3_outputs(5062)) xor (layer3_outputs(523));
    layer4_outputs(2093) <= layer3_outputs(3951);
    layer4_outputs(2094) <= (layer3_outputs(4288)) or (layer3_outputs(3936));
    layer4_outputs(2095) <= not((layer3_outputs(276)) or (layer3_outputs(3272)));
    layer4_outputs(2096) <= not(layer3_outputs(7717));
    layer4_outputs(2097) <= layer3_outputs(8185);
    layer4_outputs(2098) <= layer3_outputs(697);
    layer4_outputs(2099) <= not(layer3_outputs(9091));
    layer4_outputs(2100) <= not(layer3_outputs(4274));
    layer4_outputs(2101) <= not((layer3_outputs(5693)) xor (layer3_outputs(6995)));
    layer4_outputs(2102) <= not(layer3_outputs(3400));
    layer4_outputs(2103) <= not(layer3_outputs(5314));
    layer4_outputs(2104) <= '0';
    layer4_outputs(2105) <= layer3_outputs(6554);
    layer4_outputs(2106) <= layer3_outputs(6121);
    layer4_outputs(2107) <= layer3_outputs(2868);
    layer4_outputs(2108) <= layer3_outputs(4515);
    layer4_outputs(2109) <= not((layer3_outputs(6689)) xor (layer3_outputs(4238)));
    layer4_outputs(2110) <= (layer3_outputs(3674)) xor (layer3_outputs(5127));
    layer4_outputs(2111) <= '1';
    layer4_outputs(2112) <= not(layer3_outputs(3352));
    layer4_outputs(2113) <= not(layer3_outputs(9729)) or (layer3_outputs(6476));
    layer4_outputs(2114) <= (layer3_outputs(6377)) and not (layer3_outputs(5259));
    layer4_outputs(2115) <= layer3_outputs(5932);
    layer4_outputs(2116) <= layer3_outputs(5851);
    layer4_outputs(2117) <= layer3_outputs(2516);
    layer4_outputs(2118) <= layer3_outputs(8168);
    layer4_outputs(2119) <= layer3_outputs(3541);
    layer4_outputs(2120) <= layer3_outputs(938);
    layer4_outputs(2121) <= not(layer3_outputs(762));
    layer4_outputs(2122) <= layer3_outputs(3636);
    layer4_outputs(2123) <= not(layer3_outputs(2555));
    layer4_outputs(2124) <= not(layer3_outputs(2863));
    layer4_outputs(2125) <= layer3_outputs(8665);
    layer4_outputs(2126) <= not(layer3_outputs(6171));
    layer4_outputs(2127) <= layer3_outputs(7919);
    layer4_outputs(2128) <= layer3_outputs(8694);
    layer4_outputs(2129) <= not(layer3_outputs(920));
    layer4_outputs(2130) <= not((layer3_outputs(6328)) or (layer3_outputs(1668)));
    layer4_outputs(2131) <= (layer3_outputs(3140)) and not (layer3_outputs(4927));
    layer4_outputs(2132) <= not(layer3_outputs(8355)) or (layer3_outputs(676));
    layer4_outputs(2133) <= not(layer3_outputs(4135));
    layer4_outputs(2134) <= not(layer3_outputs(2539));
    layer4_outputs(2135) <= (layer3_outputs(4771)) and not (layer3_outputs(797));
    layer4_outputs(2136) <= (layer3_outputs(8307)) and not (layer3_outputs(5672));
    layer4_outputs(2137) <= layer3_outputs(2183);
    layer4_outputs(2138) <= layer3_outputs(2175);
    layer4_outputs(2139) <= (layer3_outputs(3919)) xor (layer3_outputs(1574));
    layer4_outputs(2140) <= layer3_outputs(8272);
    layer4_outputs(2141) <= (layer3_outputs(8759)) or (layer3_outputs(7708));
    layer4_outputs(2142) <= layer3_outputs(3788);
    layer4_outputs(2143) <= not(layer3_outputs(1142));
    layer4_outputs(2144) <= not(layer3_outputs(28)) or (layer3_outputs(2302));
    layer4_outputs(2145) <= not(layer3_outputs(5967));
    layer4_outputs(2146) <= (layer3_outputs(7108)) xor (layer3_outputs(3053));
    layer4_outputs(2147) <= (layer3_outputs(9191)) or (layer3_outputs(8944));
    layer4_outputs(2148) <= layer3_outputs(716);
    layer4_outputs(2149) <= (layer3_outputs(6883)) and not (layer3_outputs(250));
    layer4_outputs(2150) <= not((layer3_outputs(2492)) or (layer3_outputs(7990)));
    layer4_outputs(2151) <= not(layer3_outputs(7778));
    layer4_outputs(2152) <= not(layer3_outputs(5548));
    layer4_outputs(2153) <= not((layer3_outputs(5378)) xor (layer3_outputs(7106)));
    layer4_outputs(2154) <= not(layer3_outputs(1053));
    layer4_outputs(2155) <= not((layer3_outputs(1939)) and (layer3_outputs(2464)));
    layer4_outputs(2156) <= not(layer3_outputs(9159)) or (layer3_outputs(5055));
    layer4_outputs(2157) <= not(layer3_outputs(3842));
    layer4_outputs(2158) <= (layer3_outputs(1749)) and not (layer3_outputs(5781));
    layer4_outputs(2159) <= not(layer3_outputs(1718));
    layer4_outputs(2160) <= not((layer3_outputs(8564)) and (layer3_outputs(6401)));
    layer4_outputs(2161) <= not(layer3_outputs(3360));
    layer4_outputs(2162) <= not(layer3_outputs(9994));
    layer4_outputs(2163) <= not((layer3_outputs(39)) and (layer3_outputs(9717)));
    layer4_outputs(2164) <= layer3_outputs(4393);
    layer4_outputs(2165) <= not((layer3_outputs(3065)) and (layer3_outputs(1012)));
    layer4_outputs(2166) <= layer3_outputs(6629);
    layer4_outputs(2167) <= (layer3_outputs(7070)) or (layer3_outputs(3841));
    layer4_outputs(2168) <= layer3_outputs(3511);
    layer4_outputs(2169) <= not(layer3_outputs(1061));
    layer4_outputs(2170) <= (layer3_outputs(2551)) xor (layer3_outputs(7453));
    layer4_outputs(2171) <= not((layer3_outputs(4465)) or (layer3_outputs(8320)));
    layer4_outputs(2172) <= layer3_outputs(727);
    layer4_outputs(2173) <= (layer3_outputs(1585)) xor (layer3_outputs(9655));
    layer4_outputs(2174) <= (layer3_outputs(8935)) or (layer3_outputs(3676));
    layer4_outputs(2175) <= (layer3_outputs(1613)) xor (layer3_outputs(8674));
    layer4_outputs(2176) <= not(layer3_outputs(7100));
    layer4_outputs(2177) <= not(layer3_outputs(683));
    layer4_outputs(2178) <= not((layer3_outputs(1463)) xor (layer3_outputs(4065)));
    layer4_outputs(2179) <= layer3_outputs(6456);
    layer4_outputs(2180) <= not((layer3_outputs(8465)) and (layer3_outputs(5393)));
    layer4_outputs(2181) <= layer3_outputs(8067);
    layer4_outputs(2182) <= (layer3_outputs(269)) and (layer3_outputs(8829));
    layer4_outputs(2183) <= not(layer3_outputs(5150));
    layer4_outputs(2184) <= (layer3_outputs(9478)) or (layer3_outputs(5913));
    layer4_outputs(2185) <= layer3_outputs(7020);
    layer4_outputs(2186) <= layer3_outputs(4559);
    layer4_outputs(2187) <= not((layer3_outputs(1319)) xor (layer3_outputs(7673)));
    layer4_outputs(2188) <= layer3_outputs(1084);
    layer4_outputs(2189) <= layer3_outputs(1898);
    layer4_outputs(2190) <= not(layer3_outputs(7533));
    layer4_outputs(2191) <= (layer3_outputs(7152)) and not (layer3_outputs(5355));
    layer4_outputs(2192) <= not(layer3_outputs(3033)) or (layer3_outputs(7872));
    layer4_outputs(2193) <= layer3_outputs(7048);
    layer4_outputs(2194) <= not(layer3_outputs(8783));
    layer4_outputs(2195) <= layer3_outputs(8675);
    layer4_outputs(2196) <= not(layer3_outputs(3529));
    layer4_outputs(2197) <= (layer3_outputs(6643)) or (layer3_outputs(9630));
    layer4_outputs(2198) <= not(layer3_outputs(5101)) or (layer3_outputs(9411));
    layer4_outputs(2199) <= layer3_outputs(9604);
    layer4_outputs(2200) <= not(layer3_outputs(6594));
    layer4_outputs(2201) <= layer3_outputs(3463);
    layer4_outputs(2202) <= layer3_outputs(5187);
    layer4_outputs(2203) <= not(layer3_outputs(6495));
    layer4_outputs(2204) <= not((layer3_outputs(9693)) xor (layer3_outputs(2632)));
    layer4_outputs(2205) <= not((layer3_outputs(445)) xor (layer3_outputs(493)));
    layer4_outputs(2206) <= not(layer3_outputs(268)) or (layer3_outputs(7722));
    layer4_outputs(2207) <= not(layer3_outputs(9703));
    layer4_outputs(2208) <= (layer3_outputs(1343)) xor (layer3_outputs(5392));
    layer4_outputs(2209) <= not(layer3_outputs(3060));
    layer4_outputs(2210) <= layer3_outputs(9584);
    layer4_outputs(2211) <= (layer3_outputs(1508)) xor (layer3_outputs(5922));
    layer4_outputs(2212) <= layer3_outputs(1995);
    layer4_outputs(2213) <= layer3_outputs(5076);
    layer4_outputs(2214) <= not(layer3_outputs(9941));
    layer4_outputs(2215) <= layer3_outputs(5976);
    layer4_outputs(2216) <= not(layer3_outputs(8256));
    layer4_outputs(2217) <= not(layer3_outputs(5280));
    layer4_outputs(2218) <= (layer3_outputs(500)) and not (layer3_outputs(6675));
    layer4_outputs(2219) <= layer3_outputs(7629);
    layer4_outputs(2220) <= layer3_outputs(951);
    layer4_outputs(2221) <= (layer3_outputs(2317)) and (layer3_outputs(8364));
    layer4_outputs(2222) <= not(layer3_outputs(9684));
    layer4_outputs(2223) <= not(layer3_outputs(9307));
    layer4_outputs(2224) <= not(layer3_outputs(9626));
    layer4_outputs(2225) <= layer3_outputs(4320);
    layer4_outputs(2226) <= not(layer3_outputs(5699)) or (layer3_outputs(3848));
    layer4_outputs(2227) <= not((layer3_outputs(7916)) or (layer3_outputs(1445)));
    layer4_outputs(2228) <= layer3_outputs(4122);
    layer4_outputs(2229) <= not(layer3_outputs(557));
    layer4_outputs(2230) <= not(layer3_outputs(162)) or (layer3_outputs(7358));
    layer4_outputs(2231) <= (layer3_outputs(7687)) xor (layer3_outputs(9796));
    layer4_outputs(2232) <= (layer3_outputs(9331)) xor (layer3_outputs(4181));
    layer4_outputs(2233) <= layer3_outputs(5736);
    layer4_outputs(2234) <= (layer3_outputs(2620)) xor (layer3_outputs(8685));
    layer4_outputs(2235) <= not(layer3_outputs(6804));
    layer4_outputs(2236) <= layer3_outputs(8751);
    layer4_outputs(2237) <= not(layer3_outputs(3));
    layer4_outputs(2238) <= not((layer3_outputs(6005)) and (layer3_outputs(3882)));
    layer4_outputs(2239) <= not(layer3_outputs(5091));
    layer4_outputs(2240) <= not(layer3_outputs(9161));
    layer4_outputs(2241) <= not(layer3_outputs(6496)) or (layer3_outputs(901));
    layer4_outputs(2242) <= not((layer3_outputs(2444)) or (layer3_outputs(2566)));
    layer4_outputs(2243) <= layer3_outputs(6413);
    layer4_outputs(2244) <= (layer3_outputs(9706)) and (layer3_outputs(5041));
    layer4_outputs(2245) <= layer3_outputs(10126);
    layer4_outputs(2246) <= '1';
    layer4_outputs(2247) <= not(layer3_outputs(9850));
    layer4_outputs(2248) <= layer3_outputs(9015);
    layer4_outputs(2249) <= not((layer3_outputs(459)) or (layer3_outputs(4815)));
    layer4_outputs(2250) <= not(layer3_outputs(6829)) or (layer3_outputs(2349));
    layer4_outputs(2251) <= not(layer3_outputs(1251));
    layer4_outputs(2252) <= not(layer3_outputs(56));
    layer4_outputs(2253) <= layer3_outputs(5135);
    layer4_outputs(2254) <= (layer3_outputs(5802)) or (layer3_outputs(9347));
    layer4_outputs(2255) <= layer3_outputs(16);
    layer4_outputs(2256) <= not(layer3_outputs(8231));
    layer4_outputs(2257) <= (layer3_outputs(3440)) xor (layer3_outputs(8402));
    layer4_outputs(2258) <= (layer3_outputs(7942)) and not (layer3_outputs(7377));
    layer4_outputs(2259) <= (layer3_outputs(1936)) and (layer3_outputs(2089));
    layer4_outputs(2260) <= not(layer3_outputs(2670));
    layer4_outputs(2261) <= layer3_outputs(6336);
    layer4_outputs(2262) <= layer3_outputs(7226);
    layer4_outputs(2263) <= not(layer3_outputs(5886));
    layer4_outputs(2264) <= not(layer3_outputs(6619)) or (layer3_outputs(1089));
    layer4_outputs(2265) <= not((layer3_outputs(1148)) xor (layer3_outputs(4687)));
    layer4_outputs(2266) <= not(layer3_outputs(9946));
    layer4_outputs(2267) <= (layer3_outputs(7940)) and (layer3_outputs(3721));
    layer4_outputs(2268) <= not(layer3_outputs(485));
    layer4_outputs(2269) <= not(layer3_outputs(8762));
    layer4_outputs(2270) <= layer3_outputs(8079);
    layer4_outputs(2271) <= not(layer3_outputs(2398));
    layer4_outputs(2272) <= not((layer3_outputs(690)) or (layer3_outputs(8441)));
    layer4_outputs(2273) <= layer3_outputs(2401);
    layer4_outputs(2274) <= (layer3_outputs(3492)) and not (layer3_outputs(4958));
    layer4_outputs(2275) <= (layer3_outputs(7530)) or (layer3_outputs(5410));
    layer4_outputs(2276) <= (layer3_outputs(3813)) or (layer3_outputs(8262));
    layer4_outputs(2277) <= (layer3_outputs(413)) and not (layer3_outputs(7138));
    layer4_outputs(2278) <= '1';
    layer4_outputs(2279) <= (layer3_outputs(9815)) or (layer3_outputs(743));
    layer4_outputs(2280) <= not(layer3_outputs(9053));
    layer4_outputs(2281) <= (layer3_outputs(5109)) xor (layer3_outputs(1174));
    layer4_outputs(2282) <= layer3_outputs(1838);
    layer4_outputs(2283) <= not(layer3_outputs(4176));
    layer4_outputs(2284) <= layer3_outputs(1773);
    layer4_outputs(2285) <= not((layer3_outputs(450)) xor (layer3_outputs(7260)));
    layer4_outputs(2286) <= not(layer3_outputs(2786));
    layer4_outputs(2287) <= (layer3_outputs(3653)) xor (layer3_outputs(1358));
    layer4_outputs(2288) <= layer3_outputs(10110);
    layer4_outputs(2289) <= layer3_outputs(3928);
    layer4_outputs(2290) <= not((layer3_outputs(6719)) or (layer3_outputs(4621)));
    layer4_outputs(2291) <= not((layer3_outputs(2041)) or (layer3_outputs(9586)));
    layer4_outputs(2292) <= not(layer3_outputs(6123));
    layer4_outputs(2293) <= not(layer3_outputs(2162));
    layer4_outputs(2294) <= layer3_outputs(623);
    layer4_outputs(2295) <= layer3_outputs(3161);
    layer4_outputs(2296) <= not(layer3_outputs(5672));
    layer4_outputs(2297) <= (layer3_outputs(7141)) and not (layer3_outputs(3638));
    layer4_outputs(2298) <= not((layer3_outputs(3583)) and (layer3_outputs(6216)));
    layer4_outputs(2299) <= (layer3_outputs(3019)) or (layer3_outputs(9303));
    layer4_outputs(2300) <= '0';
    layer4_outputs(2301) <= (layer3_outputs(7104)) and not (layer3_outputs(3937));
    layer4_outputs(2302) <= not(layer3_outputs(5533));
    layer4_outputs(2303) <= layer3_outputs(4673);
    layer4_outputs(2304) <= (layer3_outputs(4798)) xor (layer3_outputs(6769));
    layer4_outputs(2305) <= layer3_outputs(10127);
    layer4_outputs(2306) <= (layer3_outputs(5910)) and (layer3_outputs(8242));
    layer4_outputs(2307) <= not((layer3_outputs(3537)) or (layer3_outputs(4303)));
    layer4_outputs(2308) <= layer3_outputs(6122);
    layer4_outputs(2309) <= not(layer3_outputs(8557));
    layer4_outputs(2310) <= not(layer3_outputs(7843));
    layer4_outputs(2311) <= layer3_outputs(3448);
    layer4_outputs(2312) <= (layer3_outputs(4056)) or (layer3_outputs(7510));
    layer4_outputs(2313) <= (layer3_outputs(102)) or (layer3_outputs(2940));
    layer4_outputs(2314) <= not(layer3_outputs(8407)) or (layer3_outputs(9589));
    layer4_outputs(2315) <= not(layer3_outputs(4614));
    layer4_outputs(2316) <= layer3_outputs(1923);
    layer4_outputs(2317) <= layer3_outputs(8873);
    layer4_outputs(2318) <= layer3_outputs(6298);
    layer4_outputs(2319) <= not(layer3_outputs(3559));
    layer4_outputs(2320) <= not(layer3_outputs(6729));
    layer4_outputs(2321) <= layer3_outputs(10232);
    layer4_outputs(2322) <= layer3_outputs(1273);
    layer4_outputs(2323) <= not(layer3_outputs(2399));
    layer4_outputs(2324) <= not(layer3_outputs(2052));
    layer4_outputs(2325) <= not((layer3_outputs(5025)) xor (layer3_outputs(2887)));
    layer4_outputs(2326) <= not(layer3_outputs(7762));
    layer4_outputs(2327) <= not((layer3_outputs(4685)) xor (layer3_outputs(6063)));
    layer4_outputs(2328) <= (layer3_outputs(1358)) and not (layer3_outputs(3569));
    layer4_outputs(2329) <= (layer3_outputs(1504)) and (layer3_outputs(6329));
    layer4_outputs(2330) <= not((layer3_outputs(883)) and (layer3_outputs(3833)));
    layer4_outputs(2331) <= not(layer3_outputs(9302));
    layer4_outputs(2332) <= (layer3_outputs(3438)) xor (layer3_outputs(3429));
    layer4_outputs(2333) <= (layer3_outputs(1379)) xor (layer3_outputs(374));
    layer4_outputs(2334) <= (layer3_outputs(1738)) and not (layer3_outputs(5433));
    layer4_outputs(2335) <= not(layer3_outputs(2523));
    layer4_outputs(2336) <= layer3_outputs(5520);
    layer4_outputs(2337) <= (layer3_outputs(7438)) xor (layer3_outputs(6091));
    layer4_outputs(2338) <= not((layer3_outputs(288)) or (layer3_outputs(5222)));
    layer4_outputs(2339) <= (layer3_outputs(4767)) and not (layer3_outputs(6912));
    layer4_outputs(2340) <= not(layer3_outputs(1204));
    layer4_outputs(2341) <= not(layer3_outputs(10086));
    layer4_outputs(2342) <= not((layer3_outputs(2909)) xor (layer3_outputs(5370)));
    layer4_outputs(2343) <= not((layer3_outputs(10091)) xor (layer3_outputs(883)));
    layer4_outputs(2344) <= layer3_outputs(8373);
    layer4_outputs(2345) <= not(layer3_outputs(7834)) or (layer3_outputs(8081));
    layer4_outputs(2346) <= (layer3_outputs(4712)) xor (layer3_outputs(4882));
    layer4_outputs(2347) <= '0';
    layer4_outputs(2348) <= not(layer3_outputs(8770));
    layer4_outputs(2349) <= not(layer3_outputs(345));
    layer4_outputs(2350) <= (layer3_outputs(6575)) and not (layer3_outputs(9009));
    layer4_outputs(2351) <= (layer3_outputs(1060)) or (layer3_outputs(5180));
    layer4_outputs(2352) <= not((layer3_outputs(3116)) xor (layer3_outputs(7240)));
    layer4_outputs(2353) <= not((layer3_outputs(7752)) or (layer3_outputs(7957)));
    layer4_outputs(2354) <= not(layer3_outputs(9024));
    layer4_outputs(2355) <= (layer3_outputs(2508)) and not (layer3_outputs(4609));
    layer4_outputs(2356) <= (layer3_outputs(5053)) xor (layer3_outputs(9345));
    layer4_outputs(2357) <= not((layer3_outputs(3349)) or (layer3_outputs(9491)));
    layer4_outputs(2358) <= (layer3_outputs(6667)) xor (layer3_outputs(1573));
    layer4_outputs(2359) <= layer3_outputs(1755);
    layer4_outputs(2360) <= layer3_outputs(8717);
    layer4_outputs(2361) <= layer3_outputs(4196);
    layer4_outputs(2362) <= layer3_outputs(1609);
    layer4_outputs(2363) <= not((layer3_outputs(9801)) and (layer3_outputs(2220)));
    layer4_outputs(2364) <= (layer3_outputs(1115)) or (layer3_outputs(198));
    layer4_outputs(2365) <= not((layer3_outputs(2533)) and (layer3_outputs(1796)));
    layer4_outputs(2366) <= (layer3_outputs(7044)) xor (layer3_outputs(9886));
    layer4_outputs(2367) <= (layer3_outputs(6812)) xor (layer3_outputs(2720));
    layer4_outputs(2368) <= (layer3_outputs(10127)) or (layer3_outputs(997));
    layer4_outputs(2369) <= layer3_outputs(7168);
    layer4_outputs(2370) <= layer3_outputs(101);
    layer4_outputs(2371) <= (layer3_outputs(7510)) and not (layer3_outputs(376));
    layer4_outputs(2372) <= not((layer3_outputs(2834)) xor (layer3_outputs(1878)));
    layer4_outputs(2373) <= not(layer3_outputs(4201));
    layer4_outputs(2374) <= not(layer3_outputs(6582));
    layer4_outputs(2375) <= not(layer3_outputs(8974));
    layer4_outputs(2376) <= (layer3_outputs(1898)) xor (layer3_outputs(8158));
    layer4_outputs(2377) <= (layer3_outputs(8961)) and not (layer3_outputs(3769));
    layer4_outputs(2378) <= (layer3_outputs(1534)) xor (layer3_outputs(7646));
    layer4_outputs(2379) <= (layer3_outputs(4504)) and (layer3_outputs(7684));
    layer4_outputs(2380) <= layer3_outputs(8327);
    layer4_outputs(2381) <= not(layer3_outputs(5334)) or (layer3_outputs(8739));
    layer4_outputs(2382) <= layer3_outputs(8768);
    layer4_outputs(2383) <= not(layer3_outputs(9732)) or (layer3_outputs(6369));
    layer4_outputs(2384) <= (layer3_outputs(5274)) and (layer3_outputs(8908));
    layer4_outputs(2385) <= layer3_outputs(3673);
    layer4_outputs(2386) <= not(layer3_outputs(4093));
    layer4_outputs(2387) <= (layer3_outputs(2420)) and (layer3_outputs(2011));
    layer4_outputs(2388) <= layer3_outputs(7950);
    layer4_outputs(2389) <= (layer3_outputs(5959)) or (layer3_outputs(5230));
    layer4_outputs(2390) <= layer3_outputs(1953);
    layer4_outputs(2391) <= '0';
    layer4_outputs(2392) <= not(layer3_outputs(7592)) or (layer3_outputs(2576));
    layer4_outputs(2393) <= not(layer3_outputs(8547)) or (layer3_outputs(7383));
    layer4_outputs(2394) <= layer3_outputs(4937);
    layer4_outputs(2395) <= layer3_outputs(4867);
    layer4_outputs(2396) <= '0';
    layer4_outputs(2397) <= not(layer3_outputs(7988));
    layer4_outputs(2398) <= layer3_outputs(5794);
    layer4_outputs(2399) <= not(layer3_outputs(6458)) or (layer3_outputs(2687));
    layer4_outputs(2400) <= layer3_outputs(673);
    layer4_outputs(2401) <= not((layer3_outputs(3234)) and (layer3_outputs(7953)));
    layer4_outputs(2402) <= not(layer3_outputs(3429));
    layer4_outputs(2403) <= (layer3_outputs(1080)) and not (layer3_outputs(3347));
    layer4_outputs(2404) <= not(layer3_outputs(6185));
    layer4_outputs(2405) <= not(layer3_outputs(10156));
    layer4_outputs(2406) <= not((layer3_outputs(6537)) and (layer3_outputs(8611)));
    layer4_outputs(2407) <= (layer3_outputs(5892)) and not (layer3_outputs(6780));
    layer4_outputs(2408) <= not(layer3_outputs(3875)) or (layer3_outputs(219));
    layer4_outputs(2409) <= not(layer3_outputs(7342));
    layer4_outputs(2410) <= not(layer3_outputs(1138));
    layer4_outputs(2411) <= not(layer3_outputs(8071));
    layer4_outputs(2412) <= layer3_outputs(7570);
    layer4_outputs(2413) <= not((layer3_outputs(148)) xor (layer3_outputs(5112)));
    layer4_outputs(2414) <= not(layer3_outputs(346));
    layer4_outputs(2415) <= not(layer3_outputs(6565));
    layer4_outputs(2416) <= (layer3_outputs(10186)) or (layer3_outputs(9065));
    layer4_outputs(2417) <= not(layer3_outputs(4548));
    layer4_outputs(2418) <= (layer3_outputs(1837)) xor (layer3_outputs(8939));
    layer4_outputs(2419) <= not((layer3_outputs(9740)) xor (layer3_outputs(3364)));
    layer4_outputs(2420) <= (layer3_outputs(6089)) xor (layer3_outputs(3124));
    layer4_outputs(2421) <= not(layer3_outputs(7805));
    layer4_outputs(2422) <= not((layer3_outputs(9096)) xor (layer3_outputs(647)));
    layer4_outputs(2423) <= layer3_outputs(2299);
    layer4_outputs(2424) <= (layer3_outputs(581)) and (layer3_outputs(9266));
    layer4_outputs(2425) <= not((layer3_outputs(8907)) xor (layer3_outputs(1267)));
    layer4_outputs(2426) <= not(layer3_outputs(7806));
    layer4_outputs(2427) <= layer3_outputs(1386);
    layer4_outputs(2428) <= layer3_outputs(3963);
    layer4_outputs(2429) <= not((layer3_outputs(9100)) or (layer3_outputs(8568)));
    layer4_outputs(2430) <= (layer3_outputs(3527)) and not (layer3_outputs(7938));
    layer4_outputs(2431) <= (layer3_outputs(7698)) xor (layer3_outputs(8245));
    layer4_outputs(2432) <= not(layer3_outputs(4648));
    layer4_outputs(2433) <= not(layer3_outputs(1816));
    layer4_outputs(2434) <= layer3_outputs(4098);
    layer4_outputs(2435) <= not(layer3_outputs(7242));
    layer4_outputs(2436) <= not((layer3_outputs(3591)) or (layer3_outputs(8034)));
    layer4_outputs(2437) <= not(layer3_outputs(1589));
    layer4_outputs(2438) <= '1';
    layer4_outputs(2439) <= (layer3_outputs(6975)) or (layer3_outputs(2798));
    layer4_outputs(2440) <= not(layer3_outputs(102));
    layer4_outputs(2441) <= not((layer3_outputs(10034)) xor (layer3_outputs(3952)));
    layer4_outputs(2442) <= not((layer3_outputs(7953)) and (layer3_outputs(492)));
    layer4_outputs(2443) <= (layer3_outputs(3713)) and not (layer3_outputs(2654));
    layer4_outputs(2444) <= layer3_outputs(1835);
    layer4_outputs(2445) <= not(layer3_outputs(7971));
    layer4_outputs(2446) <= not(layer3_outputs(6605));
    layer4_outputs(2447) <= layer3_outputs(1399);
    layer4_outputs(2448) <= not(layer3_outputs(4306)) or (layer3_outputs(9025));
    layer4_outputs(2449) <= not(layer3_outputs(8747));
    layer4_outputs(2450) <= not(layer3_outputs(7214));
    layer4_outputs(2451) <= not(layer3_outputs(9924));
    layer4_outputs(2452) <= layer3_outputs(2698);
    layer4_outputs(2453) <= layer3_outputs(786);
    layer4_outputs(2454) <= (layer3_outputs(3375)) and (layer3_outputs(9601));
    layer4_outputs(2455) <= (layer3_outputs(4632)) or (layer3_outputs(1981));
    layer4_outputs(2456) <= layer3_outputs(5689);
    layer4_outputs(2457) <= layer3_outputs(8165);
    layer4_outputs(2458) <= not((layer3_outputs(9926)) xor (layer3_outputs(2695)));
    layer4_outputs(2459) <= layer3_outputs(7709);
    layer4_outputs(2460) <= (layer3_outputs(5078)) xor (layer3_outputs(2832));
    layer4_outputs(2461) <= (layer3_outputs(4241)) xor (layer3_outputs(379));
    layer4_outputs(2462) <= layer3_outputs(5787);
    layer4_outputs(2463) <= not((layer3_outputs(5989)) and (layer3_outputs(3062)));
    layer4_outputs(2464) <= not((layer3_outputs(679)) xor (layer3_outputs(8630)));
    layer4_outputs(2465) <= (layer3_outputs(7058)) and not (layer3_outputs(3278));
    layer4_outputs(2466) <= not((layer3_outputs(9836)) or (layer3_outputs(5812)));
    layer4_outputs(2467) <= not((layer3_outputs(7839)) or (layer3_outputs(9966)));
    layer4_outputs(2468) <= layer3_outputs(3031);
    layer4_outputs(2469) <= not((layer3_outputs(1223)) or (layer3_outputs(3475)));
    layer4_outputs(2470) <= not(layer3_outputs(5351));
    layer4_outputs(2471) <= layer3_outputs(4951);
    layer4_outputs(2472) <= not(layer3_outputs(3849));
    layer4_outputs(2473) <= (layer3_outputs(5650)) xor (layer3_outputs(5742));
    layer4_outputs(2474) <= not(layer3_outputs(4901)) or (layer3_outputs(7867));
    layer4_outputs(2475) <= not(layer3_outputs(6655)) or (layer3_outputs(2177));
    layer4_outputs(2476) <= not((layer3_outputs(7917)) xor (layer3_outputs(1728)));
    layer4_outputs(2477) <= layer3_outputs(5114);
    layer4_outputs(2478) <= not(layer3_outputs(7583));
    layer4_outputs(2479) <= not((layer3_outputs(881)) xor (layer3_outputs(4784)));
    layer4_outputs(2480) <= not(layer3_outputs(4488));
    layer4_outputs(2481) <= layer3_outputs(7219);
    layer4_outputs(2482) <= not(layer3_outputs(9917));
    layer4_outputs(2483) <= not(layer3_outputs(5382));
    layer4_outputs(2484) <= not(layer3_outputs(9881)) or (layer3_outputs(5862));
    layer4_outputs(2485) <= not((layer3_outputs(7264)) xor (layer3_outputs(3269)));
    layer4_outputs(2486) <= not((layer3_outputs(8090)) xor (layer3_outputs(10202)));
    layer4_outputs(2487) <= (layer3_outputs(9183)) and not (layer3_outputs(1411));
    layer4_outputs(2488) <= layer3_outputs(1670);
    layer4_outputs(2489) <= (layer3_outputs(4125)) xor (layer3_outputs(4428));
    layer4_outputs(2490) <= not((layer3_outputs(5037)) and (layer3_outputs(3378)));
    layer4_outputs(2491) <= not((layer3_outputs(608)) xor (layer3_outputs(5733)));
    layer4_outputs(2492) <= (layer3_outputs(3593)) and (layer3_outputs(8139));
    layer4_outputs(2493) <= not((layer3_outputs(4873)) xor (layer3_outputs(2722)));
    layer4_outputs(2494) <= not((layer3_outputs(10022)) or (layer3_outputs(6622)));
    layer4_outputs(2495) <= layer3_outputs(215);
    layer4_outputs(2496) <= not((layer3_outputs(6139)) xor (layer3_outputs(1924)));
    layer4_outputs(2497) <= layer3_outputs(6261);
    layer4_outputs(2498) <= not(layer3_outputs(9854)) or (layer3_outputs(6062));
    layer4_outputs(2499) <= layer3_outputs(258);
    layer4_outputs(2500) <= (layer3_outputs(9193)) xor (layer3_outputs(7660));
    layer4_outputs(2501) <= layer3_outputs(257);
    layer4_outputs(2502) <= (layer3_outputs(1807)) and not (layer3_outputs(2577));
    layer4_outputs(2503) <= layer3_outputs(1882);
    layer4_outputs(2504) <= not((layer3_outputs(6299)) xor (layer3_outputs(7335)));
    layer4_outputs(2505) <= not(layer3_outputs(5443));
    layer4_outputs(2506) <= not(layer3_outputs(9883));
    layer4_outputs(2507) <= (layer3_outputs(8700)) or (layer3_outputs(7763));
    layer4_outputs(2508) <= (layer3_outputs(2332)) or (layer3_outputs(4205));
    layer4_outputs(2509) <= not(layer3_outputs(5058));
    layer4_outputs(2510) <= not(layer3_outputs(9493));
    layer4_outputs(2511) <= '0';
    layer4_outputs(2512) <= layer3_outputs(1906);
    layer4_outputs(2513) <= not(layer3_outputs(2308));
    layer4_outputs(2514) <= not(layer3_outputs(7301));
    layer4_outputs(2515) <= not((layer3_outputs(32)) xor (layer3_outputs(6356)));
    layer4_outputs(2516) <= (layer3_outputs(2657)) and not (layer3_outputs(4881));
    layer4_outputs(2517) <= not(layer3_outputs(4531));
    layer4_outputs(2518) <= not(layer3_outputs(10010));
    layer4_outputs(2519) <= layer3_outputs(2132);
    layer4_outputs(2520) <= layer3_outputs(991);
    layer4_outputs(2521) <= layer3_outputs(3009);
    layer4_outputs(2522) <= not(layer3_outputs(229));
    layer4_outputs(2523) <= not((layer3_outputs(1846)) xor (layer3_outputs(5637)));
    layer4_outputs(2524) <= not(layer3_outputs(301)) or (layer3_outputs(4840));
    layer4_outputs(2525) <= not((layer3_outputs(2567)) xor (layer3_outputs(642)));
    layer4_outputs(2526) <= not((layer3_outputs(2350)) and (layer3_outputs(89)));
    layer4_outputs(2527) <= not(layer3_outputs(754)) or (layer3_outputs(4934));
    layer4_outputs(2528) <= not((layer3_outputs(2556)) xor (layer3_outputs(5077)));
    layer4_outputs(2529) <= not(layer3_outputs(10224));
    layer4_outputs(2530) <= not(layer3_outputs(4970));
    layer4_outputs(2531) <= (layer3_outputs(4334)) or (layer3_outputs(8927));
    layer4_outputs(2532) <= layer3_outputs(9861);
    layer4_outputs(2533) <= not(layer3_outputs(7000));
    layer4_outputs(2534) <= layer3_outputs(6550);
    layer4_outputs(2535) <= not((layer3_outputs(6738)) and (layer3_outputs(3399)));
    layer4_outputs(2536) <= layer3_outputs(5610);
    layer4_outputs(2537) <= not((layer3_outputs(5241)) or (layer3_outputs(9529)));
    layer4_outputs(2538) <= layer3_outputs(8696);
    layer4_outputs(2539) <= layer3_outputs(3439);
    layer4_outputs(2540) <= (layer3_outputs(1694)) and not (layer3_outputs(2156));
    layer4_outputs(2541) <= '1';
    layer4_outputs(2542) <= not(layer3_outputs(7087));
    layer4_outputs(2543) <= (layer3_outputs(1535)) and not (layer3_outputs(6646));
    layer4_outputs(2544) <= not((layer3_outputs(8322)) xor (layer3_outputs(9235)));
    layer4_outputs(2545) <= not((layer3_outputs(6254)) or (layer3_outputs(5778)));
    layer4_outputs(2546) <= not((layer3_outputs(9281)) xor (layer3_outputs(10188)));
    layer4_outputs(2547) <= layer3_outputs(9592);
    layer4_outputs(2548) <= not(layer3_outputs(5080));
    layer4_outputs(2549) <= not(layer3_outputs(3629));
    layer4_outputs(2550) <= layer3_outputs(2553);
    layer4_outputs(2551) <= layer3_outputs(2596);
    layer4_outputs(2552) <= not(layer3_outputs(186));
    layer4_outputs(2553) <= not((layer3_outputs(8583)) xor (layer3_outputs(1592)));
    layer4_outputs(2554) <= not(layer3_outputs(6972));
    layer4_outputs(2555) <= (layer3_outputs(7074)) and not (layer3_outputs(2263));
    layer4_outputs(2556) <= layer3_outputs(354);
    layer4_outputs(2557) <= not(layer3_outputs(5614)) or (layer3_outputs(82));
    layer4_outputs(2558) <= layer3_outputs(7705);
    layer4_outputs(2559) <= not((layer3_outputs(2272)) and (layer3_outputs(7969)));
    layer4_outputs(2560) <= layer3_outputs(7414);
    layer4_outputs(2561) <= layer3_outputs(2315);
    layer4_outputs(2562) <= not(layer3_outputs(10143));
    layer4_outputs(2563) <= not(layer3_outputs(2433));
    layer4_outputs(2564) <= not((layer3_outputs(5605)) xor (layer3_outputs(8284)));
    layer4_outputs(2565) <= not(layer3_outputs(618));
    layer4_outputs(2566) <= not(layer3_outputs(9244));
    layer4_outputs(2567) <= not(layer3_outputs(628));
    layer4_outputs(2568) <= (layer3_outputs(1631)) and (layer3_outputs(4091));
    layer4_outputs(2569) <= layer3_outputs(5461);
    layer4_outputs(2570) <= layer3_outputs(7671);
    layer4_outputs(2571) <= layer3_outputs(5822);
    layer4_outputs(2572) <= not(layer3_outputs(3993));
    layer4_outputs(2573) <= not(layer3_outputs(4140));
    layer4_outputs(2574) <= not(layer3_outputs(5702));
    layer4_outputs(2575) <= (layer3_outputs(6722)) and not (layer3_outputs(4195));
    layer4_outputs(2576) <= not((layer3_outputs(484)) xor (layer3_outputs(4452)));
    layer4_outputs(2577) <= not((layer3_outputs(5514)) or (layer3_outputs(2404)));
    layer4_outputs(2578) <= not(layer3_outputs(7748));
    layer4_outputs(2579) <= not(layer3_outputs(6608));
    layer4_outputs(2580) <= not(layer3_outputs(1893));
    layer4_outputs(2581) <= layer3_outputs(5048);
    layer4_outputs(2582) <= layer3_outputs(2807);
    layer4_outputs(2583) <= not(layer3_outputs(1005));
    layer4_outputs(2584) <= not(layer3_outputs(3476));
    layer4_outputs(2585) <= layer3_outputs(334);
    layer4_outputs(2586) <= not((layer3_outputs(7848)) xor (layer3_outputs(7517)));
    layer4_outputs(2587) <= layer3_outputs(6594);
    layer4_outputs(2588) <= (layer3_outputs(6787)) or (layer3_outputs(3584));
    layer4_outputs(2589) <= (layer3_outputs(2400)) and (layer3_outputs(9582));
    layer4_outputs(2590) <= (layer3_outputs(9619)) and not (layer3_outputs(6350));
    layer4_outputs(2591) <= not((layer3_outputs(2864)) and (layer3_outputs(9431)));
    layer4_outputs(2592) <= (layer3_outputs(7811)) and (layer3_outputs(751));
    layer4_outputs(2593) <= (layer3_outputs(694)) and (layer3_outputs(8881));
    layer4_outputs(2594) <= layer3_outputs(10007);
    layer4_outputs(2595) <= not((layer3_outputs(6528)) and (layer3_outputs(5780)));
    layer4_outputs(2596) <= (layer3_outputs(2071)) and not (layer3_outputs(1501));
    layer4_outputs(2597) <= (layer3_outputs(1029)) and not (layer3_outputs(8416));
    layer4_outputs(2598) <= layer3_outputs(8731);
    layer4_outputs(2599) <= layer3_outputs(8723);
    layer4_outputs(2600) <= layer3_outputs(9994);
    layer4_outputs(2601) <= not(layer3_outputs(4800));
    layer4_outputs(2602) <= not(layer3_outputs(2382)) or (layer3_outputs(1873));
    layer4_outputs(2603) <= not(layer3_outputs(5324));
    layer4_outputs(2604) <= layer3_outputs(5835);
    layer4_outputs(2605) <= layer3_outputs(1831);
    layer4_outputs(2606) <= (layer3_outputs(1390)) xor (layer3_outputs(6489));
    layer4_outputs(2607) <= not((layer3_outputs(5046)) xor (layer3_outputs(8320)));
    layer4_outputs(2608) <= layer3_outputs(3515);
    layer4_outputs(2609) <= (layer3_outputs(4594)) and not (layer3_outputs(7045));
    layer4_outputs(2610) <= (layer3_outputs(4439)) and not (layer3_outputs(7451));
    layer4_outputs(2611) <= not(layer3_outputs(3503));
    layer4_outputs(2612) <= (layer3_outputs(5718)) or (layer3_outputs(3736));
    layer4_outputs(2613) <= layer3_outputs(7829);
    layer4_outputs(2614) <= (layer3_outputs(10088)) and (layer3_outputs(7166));
    layer4_outputs(2615) <= (layer3_outputs(8666)) xor (layer3_outputs(7613));
    layer4_outputs(2616) <= not(layer3_outputs(4465));
    layer4_outputs(2617) <= layer3_outputs(2711);
    layer4_outputs(2618) <= not(layer3_outputs(4899));
    layer4_outputs(2619) <= layer3_outputs(6389);
    layer4_outputs(2620) <= (layer3_outputs(7562)) and not (layer3_outputs(7302));
    layer4_outputs(2621) <= layer3_outputs(3682);
    layer4_outputs(2622) <= layer3_outputs(1057);
    layer4_outputs(2623) <= not(layer3_outputs(8376));
    layer4_outputs(2624) <= (layer3_outputs(3705)) and not (layer3_outputs(9585));
    layer4_outputs(2625) <= not(layer3_outputs(3357));
    layer4_outputs(2626) <= not(layer3_outputs(1575));
    layer4_outputs(2627) <= not(layer3_outputs(90)) or (layer3_outputs(9146));
    layer4_outputs(2628) <= not(layer3_outputs(2095));
    layer4_outputs(2629) <= not(layer3_outputs(1114));
    layer4_outputs(2630) <= not(layer3_outputs(5969));
    layer4_outputs(2631) <= not(layer3_outputs(6729));
    layer4_outputs(2632) <= not(layer3_outputs(3702));
    layer4_outputs(2633) <= layer3_outputs(3784);
    layer4_outputs(2634) <= not(layer3_outputs(8084)) or (layer3_outputs(2229));
    layer4_outputs(2635) <= not(layer3_outputs(7634));
    layer4_outputs(2636) <= (layer3_outputs(9154)) xor (layer3_outputs(2903));
    layer4_outputs(2637) <= (layer3_outputs(4489)) and not (layer3_outputs(780));
    layer4_outputs(2638) <= layer3_outputs(5720);
    layer4_outputs(2639) <= layer3_outputs(8730);
    layer4_outputs(2640) <= (layer3_outputs(2371)) xor (layer3_outputs(8740));
    layer4_outputs(2641) <= not(layer3_outputs(692)) or (layer3_outputs(4318));
    layer4_outputs(2642) <= layer3_outputs(8318);
    layer4_outputs(2643) <= not(layer3_outputs(5558));
    layer4_outputs(2644) <= layer3_outputs(1766);
    layer4_outputs(2645) <= (layer3_outputs(3209)) or (layer3_outputs(2742));
    layer4_outputs(2646) <= not(layer3_outputs(4029)) or (layer3_outputs(164));
    layer4_outputs(2647) <= (layer3_outputs(6032)) xor (layer3_outputs(5760));
    layer4_outputs(2648) <= '0';
    layer4_outputs(2649) <= not((layer3_outputs(3504)) or (layer3_outputs(4285)));
    layer4_outputs(2650) <= not(layer3_outputs(3348)) or (layer3_outputs(580));
    layer4_outputs(2651) <= layer3_outputs(8308);
    layer4_outputs(2652) <= not((layer3_outputs(2530)) and (layer3_outputs(4827)));
    layer4_outputs(2653) <= '0';
    layer4_outputs(2654) <= (layer3_outputs(1974)) xor (layer3_outputs(3974));
    layer4_outputs(2655) <= not(layer3_outputs(9894));
    layer4_outputs(2656) <= (layer3_outputs(2516)) xor (layer3_outputs(3947));
    layer4_outputs(2657) <= (layer3_outputs(10092)) and not (layer3_outputs(2403));
    layer4_outputs(2658) <= not(layer3_outputs(5643));
    layer4_outputs(2659) <= not(layer3_outputs(5));
    layer4_outputs(2660) <= not(layer3_outputs(6454));
    layer4_outputs(2661) <= layer3_outputs(8598);
    layer4_outputs(2662) <= not(layer3_outputs(1101));
    layer4_outputs(2663) <= (layer3_outputs(6789)) and (layer3_outputs(2844));
    layer4_outputs(2664) <= layer3_outputs(2229);
    layer4_outputs(2665) <= layer3_outputs(714);
    layer4_outputs(2666) <= not(layer3_outputs(7320));
    layer4_outputs(2667) <= layer3_outputs(7549);
    layer4_outputs(2668) <= layer3_outputs(40);
    layer4_outputs(2669) <= layer3_outputs(8217);
    layer4_outputs(2670) <= not(layer3_outputs(7992));
    layer4_outputs(2671) <= (layer3_outputs(8055)) and not (layer3_outputs(7218));
    layer4_outputs(2672) <= not(layer3_outputs(2313)) or (layer3_outputs(4632));
    layer4_outputs(2673) <= not((layer3_outputs(8808)) or (layer3_outputs(7086)));
    layer4_outputs(2674) <= not((layer3_outputs(10232)) xor (layer3_outputs(7386)));
    layer4_outputs(2675) <= not((layer3_outputs(122)) xor (layer3_outputs(9739)));
    layer4_outputs(2676) <= layer3_outputs(3299);
    layer4_outputs(2677) <= layer3_outputs(995);
    layer4_outputs(2678) <= not(layer3_outputs(5877));
    layer4_outputs(2679) <= layer3_outputs(1065);
    layer4_outputs(2680) <= layer3_outputs(652);
    layer4_outputs(2681) <= layer3_outputs(8404);
    layer4_outputs(2682) <= layer3_outputs(5571);
    layer4_outputs(2683) <= layer3_outputs(8937);
    layer4_outputs(2684) <= (layer3_outputs(1928)) xor (layer3_outputs(1942));
    layer4_outputs(2685) <= (layer3_outputs(828)) xor (layer3_outputs(3805));
    layer4_outputs(2686) <= layer3_outputs(4538);
    layer4_outputs(2687) <= '0';
    layer4_outputs(2688) <= not(layer3_outputs(2820));
    layer4_outputs(2689) <= not(layer3_outputs(1935));
    layer4_outputs(2690) <= layer3_outputs(10216);
    layer4_outputs(2691) <= not((layer3_outputs(4077)) or (layer3_outputs(5307)));
    layer4_outputs(2692) <= not(layer3_outputs(1004));
    layer4_outputs(2693) <= (layer3_outputs(2641)) and not (layer3_outputs(2655));
    layer4_outputs(2694) <= layer3_outputs(10148);
    layer4_outputs(2695) <= not(layer3_outputs(4255));
    layer4_outputs(2696) <= (layer3_outputs(6133)) and not (layer3_outputs(9364));
    layer4_outputs(2697) <= layer3_outputs(3241);
    layer4_outputs(2698) <= not(layer3_outputs(5112));
    layer4_outputs(2699) <= (layer3_outputs(4879)) and not (layer3_outputs(5189));
    layer4_outputs(2700) <= not(layer3_outputs(1624));
    layer4_outputs(2701) <= layer3_outputs(803);
    layer4_outputs(2702) <= not(layer3_outputs(4200));
    layer4_outputs(2703) <= not((layer3_outputs(7263)) or (layer3_outputs(1321)));
    layer4_outputs(2704) <= layer3_outputs(3995);
    layer4_outputs(2705) <= not((layer3_outputs(4561)) and (layer3_outputs(2891)));
    layer4_outputs(2706) <= not(layer3_outputs(9212));
    layer4_outputs(2707) <= (layer3_outputs(5277)) and not (layer3_outputs(2187));
    layer4_outputs(2708) <= not(layer3_outputs(1164));
    layer4_outputs(2709) <= layer3_outputs(7462);
    layer4_outputs(2710) <= not(layer3_outputs(596)) or (layer3_outputs(2614));
    layer4_outputs(2711) <= layer3_outputs(7682);
    layer4_outputs(2712) <= layer3_outputs(4071);
    layer4_outputs(2713) <= (layer3_outputs(3538)) or (layer3_outputs(1349));
    layer4_outputs(2714) <= not(layer3_outputs(2199));
    layer4_outputs(2715) <= layer3_outputs(9433);
    layer4_outputs(2716) <= not(layer3_outputs(9501));
    layer4_outputs(2717) <= layer3_outputs(5336);
    layer4_outputs(2718) <= not(layer3_outputs(7224));
    layer4_outputs(2719) <= not(layer3_outputs(7417));
    layer4_outputs(2720) <= not((layer3_outputs(8616)) xor (layer3_outputs(5442)));
    layer4_outputs(2721) <= layer3_outputs(1907);
    layer4_outputs(2722) <= layer3_outputs(1598);
    layer4_outputs(2723) <= (layer3_outputs(5445)) xor (layer3_outputs(253));
    layer4_outputs(2724) <= layer3_outputs(2323);
    layer4_outputs(2725) <= not(layer3_outputs(4372));
    layer4_outputs(2726) <= not(layer3_outputs(791));
    layer4_outputs(2727) <= not(layer3_outputs(5624)) or (layer3_outputs(4891));
    layer4_outputs(2728) <= not(layer3_outputs(5264)) or (layer3_outputs(1544));
    layer4_outputs(2729) <= not(layer3_outputs(9633));
    layer4_outputs(2730) <= layer3_outputs(7543);
    layer4_outputs(2731) <= layer3_outputs(2637);
    layer4_outputs(2732) <= not(layer3_outputs(2798));
    layer4_outputs(2733) <= not(layer3_outputs(4002));
    layer4_outputs(2734) <= layer3_outputs(5997);
    layer4_outputs(2735) <= (layer3_outputs(4780)) xor (layer3_outputs(3337));
    layer4_outputs(2736) <= not(layer3_outputs(8646));
    layer4_outputs(2737) <= (layer3_outputs(4883)) and not (layer3_outputs(8407));
    layer4_outputs(2738) <= not((layer3_outputs(1542)) xor (layer3_outputs(8330)));
    layer4_outputs(2739) <= not(layer3_outputs(6595));
    layer4_outputs(2740) <= layer3_outputs(1523);
    layer4_outputs(2741) <= (layer3_outputs(9090)) xor (layer3_outputs(3575));
    layer4_outputs(2742) <= not(layer3_outputs(6628));
    layer4_outputs(2743) <= layer3_outputs(2869);
    layer4_outputs(2744) <= layer3_outputs(4246);
    layer4_outputs(2745) <= (layer3_outputs(4945)) or (layer3_outputs(9281));
    layer4_outputs(2746) <= layer3_outputs(4454);
    layer4_outputs(2747) <= not(layer3_outputs(4204));
    layer4_outputs(2748) <= not(layer3_outputs(109));
    layer4_outputs(2749) <= not((layer3_outputs(8684)) and (layer3_outputs(3899)));
    layer4_outputs(2750) <= layer3_outputs(1761);
    layer4_outputs(2751) <= layer3_outputs(4801);
    layer4_outputs(2752) <= (layer3_outputs(7664)) xor (layer3_outputs(7498));
    layer4_outputs(2753) <= layer3_outputs(817);
    layer4_outputs(2754) <= not(layer3_outputs(1073));
    layer4_outputs(2755) <= not(layer3_outputs(5013));
    layer4_outputs(2756) <= not(layer3_outputs(596));
    layer4_outputs(2757) <= layer3_outputs(2514);
    layer4_outputs(2758) <= (layer3_outputs(2136)) xor (layer3_outputs(7309));
    layer4_outputs(2759) <= not(layer3_outputs(5158)) or (layer3_outputs(9265));
    layer4_outputs(2760) <= not(layer3_outputs(3362)) or (layer3_outputs(5896));
    layer4_outputs(2761) <= (layer3_outputs(8827)) and not (layer3_outputs(8858));
    layer4_outputs(2762) <= (layer3_outputs(8721)) and not (layer3_outputs(4655));
    layer4_outputs(2763) <= layer3_outputs(5902);
    layer4_outputs(2764) <= not(layer3_outputs(6932));
    layer4_outputs(2765) <= layer3_outputs(5458);
    layer4_outputs(2766) <= layer3_outputs(7593);
    layer4_outputs(2767) <= (layer3_outputs(7348)) xor (layer3_outputs(6459));
    layer4_outputs(2768) <= not((layer3_outputs(4522)) xor (layer3_outputs(6895)));
    layer4_outputs(2769) <= layer3_outputs(9859);
    layer4_outputs(2770) <= layer3_outputs(8334);
    layer4_outputs(2771) <= not(layer3_outputs(4988));
    layer4_outputs(2772) <= not(layer3_outputs(1337)) or (layer3_outputs(9650));
    layer4_outputs(2773) <= layer3_outputs(298);
    layer4_outputs(2774) <= (layer3_outputs(1785)) xor (layer3_outputs(2863));
    layer4_outputs(2775) <= (layer3_outputs(6528)) xor (layer3_outputs(1596));
    layer4_outputs(2776) <= not(layer3_outputs(6049));
    layer4_outputs(2777) <= layer3_outputs(515);
    layer4_outputs(2778) <= not(layer3_outputs(5447));
    layer4_outputs(2779) <= not(layer3_outputs(964)) or (layer3_outputs(8258));
    layer4_outputs(2780) <= not(layer3_outputs(7873));
    layer4_outputs(2781) <= not(layer3_outputs(4276));
    layer4_outputs(2782) <= not(layer3_outputs(7252));
    layer4_outputs(2783) <= not(layer3_outputs(6337));
    layer4_outputs(2784) <= (layer3_outputs(6575)) and not (layer3_outputs(4657));
    layer4_outputs(2785) <= not(layer3_outputs(4021));
    layer4_outputs(2786) <= not(layer3_outputs(527));
    layer4_outputs(2787) <= (layer3_outputs(7201)) xor (layer3_outputs(8734));
    layer4_outputs(2788) <= not((layer3_outputs(10211)) and (layer3_outputs(4875)));
    layer4_outputs(2789) <= layer3_outputs(1313);
    layer4_outputs(2790) <= layer3_outputs(7096);
    layer4_outputs(2791) <= layer3_outputs(1047);
    layer4_outputs(2792) <= (layer3_outputs(7617)) and not (layer3_outputs(4205));
    layer4_outputs(2793) <= not(layer3_outputs(9024));
    layer4_outputs(2794) <= (layer3_outputs(5903)) or (layer3_outputs(445));
    layer4_outputs(2795) <= not((layer3_outputs(6017)) xor (layer3_outputs(7952)));
    layer4_outputs(2796) <= layer3_outputs(8453);
    layer4_outputs(2797) <= not(layer3_outputs(419));
    layer4_outputs(2798) <= layer3_outputs(3067);
    layer4_outputs(2799) <= not(layer3_outputs(8947));
    layer4_outputs(2800) <= (layer3_outputs(2846)) or (layer3_outputs(1322));
    layer4_outputs(2801) <= not((layer3_outputs(9082)) xor (layer3_outputs(1375)));
    layer4_outputs(2802) <= not((layer3_outputs(1014)) or (layer3_outputs(8364)));
    layer4_outputs(2803) <= layer3_outputs(3696);
    layer4_outputs(2804) <= layer3_outputs(1139);
    layer4_outputs(2805) <= (layer3_outputs(1701)) and not (layer3_outputs(1567));
    layer4_outputs(2806) <= not(layer3_outputs(1350));
    layer4_outputs(2807) <= layer3_outputs(9341);
    layer4_outputs(2808) <= not(layer3_outputs(7385));
    layer4_outputs(2809) <= (layer3_outputs(6739)) and not (layer3_outputs(5361));
    layer4_outputs(2810) <= (layer3_outputs(6941)) xor (layer3_outputs(1829));
    layer4_outputs(2811) <= not(layer3_outputs(4390));
    layer4_outputs(2812) <= not(layer3_outputs(9280));
    layer4_outputs(2813) <= layer3_outputs(2578);
    layer4_outputs(2814) <= not(layer3_outputs(7666));
    layer4_outputs(2815) <= not(layer3_outputs(1803));
    layer4_outputs(2816) <= not(layer3_outputs(9277));
    layer4_outputs(2817) <= layer3_outputs(6960);
    layer4_outputs(2818) <= (layer3_outputs(4733)) xor (layer3_outputs(1556));
    layer4_outputs(2819) <= layer3_outputs(251);
    layer4_outputs(2820) <= not(layer3_outputs(1932));
    layer4_outputs(2821) <= not(layer3_outputs(8107));
    layer4_outputs(2822) <= (layer3_outputs(9204)) or (layer3_outputs(8077));
    layer4_outputs(2823) <= not(layer3_outputs(6498)) or (layer3_outputs(8952));
    layer4_outputs(2824) <= layer3_outputs(735);
    layer4_outputs(2825) <= (layer3_outputs(5788)) and not (layer3_outputs(7470));
    layer4_outputs(2826) <= not((layer3_outputs(7421)) xor (layer3_outputs(1973)));
    layer4_outputs(2827) <= layer3_outputs(8391);
    layer4_outputs(2828) <= not(layer3_outputs(491));
    layer4_outputs(2829) <= layer3_outputs(6573);
    layer4_outputs(2830) <= not(layer3_outputs(7553));
    layer4_outputs(2831) <= (layer3_outputs(10163)) and (layer3_outputs(6612));
    layer4_outputs(2832) <= (layer3_outputs(8389)) and (layer3_outputs(8868));
    layer4_outputs(2833) <= layer3_outputs(6979);
    layer4_outputs(2834) <= not(layer3_outputs(6834));
    layer4_outputs(2835) <= (layer3_outputs(3748)) and not (layer3_outputs(4378));
    layer4_outputs(2836) <= (layer3_outputs(5923)) and not (layer3_outputs(7595));
    layer4_outputs(2837) <= not(layer3_outputs(7862));
    layer4_outputs(2838) <= layer3_outputs(8880);
    layer4_outputs(2839) <= not((layer3_outputs(5381)) and (layer3_outputs(8757)));
    layer4_outputs(2840) <= not(layer3_outputs(6838)) or (layer3_outputs(7164));
    layer4_outputs(2841) <= not(layer3_outputs(1820));
    layer4_outputs(2842) <= (layer3_outputs(6021)) and (layer3_outputs(1460));
    layer4_outputs(2843) <= not((layer3_outputs(2824)) xor (layer3_outputs(4338)));
    layer4_outputs(2844) <= not((layer3_outputs(859)) and (layer3_outputs(8172)));
    layer4_outputs(2845) <= layer3_outputs(174);
    layer4_outputs(2846) <= '0';
    layer4_outputs(2847) <= (layer3_outputs(3470)) xor (layer3_outputs(3688));
    layer4_outputs(2848) <= not((layer3_outputs(2237)) or (layer3_outputs(903)));
    layer4_outputs(2849) <= (layer3_outputs(5479)) xor (layer3_outputs(582));
    layer4_outputs(2850) <= not(layer3_outputs(10161));
    layer4_outputs(2851) <= not(layer3_outputs(4572));
    layer4_outputs(2852) <= layer3_outputs(9757);
    layer4_outputs(2853) <= layer3_outputs(5382);
    layer4_outputs(2854) <= layer3_outputs(748);
    layer4_outputs(2855) <= not(layer3_outputs(3109));
    layer4_outputs(2856) <= (layer3_outputs(9952)) xor (layer3_outputs(6726));
    layer4_outputs(2857) <= layer3_outputs(6366);
    layer4_outputs(2858) <= not(layer3_outputs(1736));
    layer4_outputs(2859) <= (layer3_outputs(8837)) and (layer3_outputs(5276));
    layer4_outputs(2860) <= layer3_outputs(6577);
    layer4_outputs(2861) <= not(layer3_outputs(7697));
    layer4_outputs(2862) <= not(layer3_outputs(9316)) or (layer3_outputs(1878));
    layer4_outputs(2863) <= not(layer3_outputs(9140));
    layer4_outputs(2864) <= not((layer3_outputs(6590)) and (layer3_outputs(8941)));
    layer4_outputs(2865) <= not(layer3_outputs(2245));
    layer4_outputs(2866) <= not(layer3_outputs(5308));
    layer4_outputs(2867) <= not((layer3_outputs(6761)) and (layer3_outputs(3784)));
    layer4_outputs(2868) <= not(layer3_outputs(2891));
    layer4_outputs(2869) <= (layer3_outputs(4841)) and not (layer3_outputs(6781));
    layer4_outputs(2870) <= not(layer3_outputs(2281));
    layer4_outputs(2871) <= not(layer3_outputs(7852));
    layer4_outputs(2872) <= (layer3_outputs(9513)) or (layer3_outputs(6744));
    layer4_outputs(2873) <= (layer3_outputs(6841)) and not (layer3_outputs(7018));
    layer4_outputs(2874) <= (layer3_outputs(2669)) xor (layer3_outputs(8550));
    layer4_outputs(2875) <= layer3_outputs(9366);
    layer4_outputs(2876) <= (layer3_outputs(8579)) and not (layer3_outputs(4395));
    layer4_outputs(2877) <= not(layer3_outputs(3094)) or (layer3_outputs(2525));
    layer4_outputs(2878) <= not(layer3_outputs(6986));
    layer4_outputs(2879) <= not(layer3_outputs(9991));
    layer4_outputs(2880) <= layer3_outputs(9099);
    layer4_outputs(2881) <= not(layer3_outputs(4323));
    layer4_outputs(2882) <= layer3_outputs(5326);
    layer4_outputs(2883) <= not(layer3_outputs(2236));
    layer4_outputs(2884) <= layer3_outputs(6135);
    layer4_outputs(2885) <= layer3_outputs(6902);
    layer4_outputs(2886) <= not(layer3_outputs(8171));
    layer4_outputs(2887) <= not(layer3_outputs(8321));
    layer4_outputs(2888) <= not(layer3_outputs(1387)) or (layer3_outputs(3661));
    layer4_outputs(2889) <= not(layer3_outputs(1021));
    layer4_outputs(2890) <= not(layer3_outputs(4292));
    layer4_outputs(2891) <= layer3_outputs(2381);
    layer4_outputs(2892) <= not(layer3_outputs(8280));
    layer4_outputs(2893) <= not(layer3_outputs(6510));
    layer4_outputs(2894) <= '0';
    layer4_outputs(2895) <= (layer3_outputs(1194)) and not (layer3_outputs(10168));
    layer4_outputs(2896) <= not(layer3_outputs(627));
    layer4_outputs(2897) <= layer3_outputs(10196);
    layer4_outputs(2898) <= layer3_outputs(7154);
    layer4_outputs(2899) <= layer3_outputs(615);
    layer4_outputs(2900) <= (layer3_outputs(1725)) and (layer3_outputs(2442));
    layer4_outputs(2901) <= layer3_outputs(2499);
    layer4_outputs(2902) <= (layer3_outputs(3458)) xor (layer3_outputs(5670));
    layer4_outputs(2903) <= layer3_outputs(4368);
    layer4_outputs(2904) <= not(layer3_outputs(7853));
    layer4_outputs(2905) <= (layer3_outputs(4459)) and (layer3_outputs(3827));
    layer4_outputs(2906) <= (layer3_outputs(7907)) and not (layer3_outputs(9761));
    layer4_outputs(2907) <= not(layer3_outputs(6481));
    layer4_outputs(2908) <= layer3_outputs(1892);
    layer4_outputs(2909) <= layer3_outputs(4519);
    layer4_outputs(2910) <= layer3_outputs(6258);
    layer4_outputs(2911) <= not(layer3_outputs(9357));
    layer4_outputs(2912) <= not((layer3_outputs(3222)) xor (layer3_outputs(470)));
    layer4_outputs(2913) <= layer3_outputs(3808);
    layer4_outputs(2914) <= layer3_outputs(1722);
    layer4_outputs(2915) <= layer3_outputs(5135);
    layer4_outputs(2916) <= not(layer3_outputs(8171));
    layer4_outputs(2917) <= (layer3_outputs(9693)) xor (layer3_outputs(9819));
    layer4_outputs(2918) <= (layer3_outputs(6914)) and not (layer3_outputs(9570));
    layer4_outputs(2919) <= (layer3_outputs(3507)) and not (layer3_outputs(2573));
    layer4_outputs(2920) <= not(layer3_outputs(852)) or (layer3_outputs(5962));
    layer4_outputs(2921) <= not((layer3_outputs(2998)) xor (layer3_outputs(3181)));
    layer4_outputs(2922) <= (layer3_outputs(4546)) and not (layer3_outputs(8106));
    layer4_outputs(2923) <= (layer3_outputs(2391)) xor (layer3_outputs(2871));
    layer4_outputs(2924) <= layer3_outputs(7185);
    layer4_outputs(2925) <= layer3_outputs(3064);
    layer4_outputs(2926) <= layer3_outputs(1536);
    layer4_outputs(2927) <= (layer3_outputs(5603)) xor (layer3_outputs(6737));
    layer4_outputs(2928) <= not(layer3_outputs(8100));
    layer4_outputs(2929) <= not((layer3_outputs(6736)) xor (layer3_outputs(8750)));
    layer4_outputs(2930) <= not(layer3_outputs(7753));
    layer4_outputs(2931) <= (layer3_outputs(6878)) and (layer3_outputs(3756));
    layer4_outputs(2932) <= not(layer3_outputs(4025));
    layer4_outputs(2933) <= (layer3_outputs(9308)) and not (layer3_outputs(7040));
    layer4_outputs(2934) <= not(layer3_outputs(7886));
    layer4_outputs(2935) <= not((layer3_outputs(1160)) xor (layer3_outputs(9569)));
    layer4_outputs(2936) <= layer3_outputs(5198);
    layer4_outputs(2937) <= not(layer3_outputs(2679));
    layer4_outputs(2938) <= (layer3_outputs(6440)) xor (layer3_outputs(5358));
    layer4_outputs(2939) <= layer3_outputs(8601);
    layer4_outputs(2940) <= not(layer3_outputs(3706));
    layer4_outputs(2941) <= (layer3_outputs(7046)) and not (layer3_outputs(2828));
    layer4_outputs(2942) <= not(layer3_outputs(5907));
    layer4_outputs(2943) <= not(layer3_outputs(1990));
    layer4_outputs(2944) <= layer3_outputs(6255);
    layer4_outputs(2945) <= not(layer3_outputs(1573));
    layer4_outputs(2946) <= not((layer3_outputs(9852)) or (layer3_outputs(7486)));
    layer4_outputs(2947) <= not(layer3_outputs(4442)) or (layer3_outputs(3861));
    layer4_outputs(2948) <= (layer3_outputs(2609)) and not (layer3_outputs(6578));
    layer4_outputs(2949) <= not((layer3_outputs(3178)) and (layer3_outputs(4461)));
    layer4_outputs(2950) <= layer3_outputs(2897);
    layer4_outputs(2951) <= not(layer3_outputs(8372));
    layer4_outputs(2952) <= (layer3_outputs(4726)) xor (layer3_outputs(5062));
    layer4_outputs(2953) <= (layer3_outputs(71)) or (layer3_outputs(2814));
    layer4_outputs(2954) <= not((layer3_outputs(2340)) and (layer3_outputs(949)));
    layer4_outputs(2955) <= not(layer3_outputs(2684));
    layer4_outputs(2956) <= not((layer3_outputs(369)) and (layer3_outputs(8745)));
    layer4_outputs(2957) <= (layer3_outputs(5690)) xor (layer3_outputs(9477));
    layer4_outputs(2958) <= layer3_outputs(6633);
    layer4_outputs(2959) <= (layer3_outputs(9405)) or (layer3_outputs(5711));
    layer4_outputs(2960) <= not((layer3_outputs(8340)) and (layer3_outputs(3050)));
    layer4_outputs(2961) <= layer3_outputs(3436);
    layer4_outputs(2962) <= not(layer3_outputs(5467));
    layer4_outputs(2963) <= (layer3_outputs(9027)) and not (layer3_outputs(10157));
    layer4_outputs(2964) <= not(layer3_outputs(1222));
    layer4_outputs(2965) <= layer3_outputs(3011);
    layer4_outputs(2966) <= not(layer3_outputs(3520));
    layer4_outputs(2967) <= not(layer3_outputs(8412));
    layer4_outputs(2968) <= layer3_outputs(5833);
    layer4_outputs(2969) <= (layer3_outputs(4169)) xor (layer3_outputs(6053));
    layer4_outputs(2970) <= layer3_outputs(8410);
    layer4_outputs(2971) <= not((layer3_outputs(5769)) or (layer3_outputs(8324)));
    layer4_outputs(2972) <= not(layer3_outputs(587));
    layer4_outputs(2973) <= layer3_outputs(6734);
    layer4_outputs(2974) <= layer3_outputs(3541);
    layer4_outputs(2975) <= not(layer3_outputs(8994)) or (layer3_outputs(2294));
    layer4_outputs(2976) <= layer3_outputs(2812);
    layer4_outputs(2977) <= (layer3_outputs(4870)) and (layer3_outputs(5999));
    layer4_outputs(2978) <= not((layer3_outputs(9838)) and (layer3_outputs(6971)));
    layer4_outputs(2979) <= layer3_outputs(2296);
    layer4_outputs(2980) <= not((layer3_outputs(3859)) or (layer3_outputs(5694)));
    layer4_outputs(2981) <= (layer3_outputs(9914)) or (layer3_outputs(4533));
    layer4_outputs(2982) <= not(layer3_outputs(3757));
    layer4_outputs(2983) <= not(layer3_outputs(6236));
    layer4_outputs(2984) <= not(layer3_outputs(7284)) or (layer3_outputs(3367));
    layer4_outputs(2985) <= layer3_outputs(4191);
    layer4_outputs(2986) <= not(layer3_outputs(4991)) or (layer3_outputs(2474));
    layer4_outputs(2987) <= not((layer3_outputs(6657)) or (layer3_outputs(4656)));
    layer4_outputs(2988) <= not(layer3_outputs(9419));
    layer4_outputs(2989) <= layer3_outputs(5836);
    layer4_outputs(2990) <= not(layer3_outputs(2402));
    layer4_outputs(2991) <= not(layer3_outputs(2795));
    layer4_outputs(2992) <= not(layer3_outputs(7428));
    layer4_outputs(2993) <= (layer3_outputs(4082)) xor (layer3_outputs(1384));
    layer4_outputs(2994) <= not((layer3_outputs(3752)) and (layer3_outputs(10064)));
    layer4_outputs(2995) <= not(layer3_outputs(1611));
    layer4_outputs(2996) <= not(layer3_outputs(10075));
    layer4_outputs(2997) <= not(layer3_outputs(3449));
    layer4_outputs(2998) <= not((layer3_outputs(2441)) xor (layer3_outputs(1266)));
    layer4_outputs(2999) <= not(layer3_outputs(8420));
    layer4_outputs(3000) <= not(layer3_outputs(2640));
    layer4_outputs(3001) <= layer3_outputs(7243);
    layer4_outputs(3002) <= (layer3_outputs(3047)) xor (layer3_outputs(8061));
    layer4_outputs(3003) <= not((layer3_outputs(6183)) and (layer3_outputs(7927)));
    layer4_outputs(3004) <= not(layer3_outputs(9131));
    layer4_outputs(3005) <= (layer3_outputs(299)) and not (layer3_outputs(4750));
    layer4_outputs(3006) <= not((layer3_outputs(801)) xor (layer3_outputs(5484)));
    layer4_outputs(3007) <= (layer3_outputs(4231)) and not (layer3_outputs(9699));
    layer4_outputs(3008) <= (layer3_outputs(2651)) and not (layer3_outputs(7485));
    layer4_outputs(3009) <= layer3_outputs(9479);
    layer4_outputs(3010) <= not((layer3_outputs(3576)) xor (layer3_outputs(8774)));
    layer4_outputs(3011) <= (layer3_outputs(5792)) and (layer3_outputs(8955));
    layer4_outputs(3012) <= (layer3_outputs(1729)) xor (layer3_outputs(7784));
    layer4_outputs(3013) <= not((layer3_outputs(4198)) xor (layer3_outputs(5295)));
    layer4_outputs(3014) <= not((layer3_outputs(9677)) and (layer3_outputs(4357)));
    layer4_outputs(3015) <= not(layer3_outputs(9371)) or (layer3_outputs(2633));
    layer4_outputs(3016) <= layer3_outputs(5770);
    layer4_outputs(3017) <= not(layer3_outputs(9735));
    layer4_outputs(3018) <= not(layer3_outputs(5085));
    layer4_outputs(3019) <= not(layer3_outputs(215));
    layer4_outputs(3020) <= layer3_outputs(5291);
    layer4_outputs(3021) <= not((layer3_outputs(9544)) and (layer3_outputs(1851)));
    layer4_outputs(3022) <= (layer3_outputs(7494)) or (layer3_outputs(9259));
    layer4_outputs(3023) <= layer3_outputs(2423);
    layer4_outputs(3024) <= not((layer3_outputs(2718)) and (layer3_outputs(8823)));
    layer4_outputs(3025) <= not(layer3_outputs(7521));
    layer4_outputs(3026) <= (layer3_outputs(8657)) or (layer3_outputs(4942));
    layer4_outputs(3027) <= layer3_outputs(314);
    layer4_outputs(3028) <= layer3_outputs(8546);
    layer4_outputs(3029) <= not((layer3_outputs(7169)) and (layer3_outputs(3526)));
    layer4_outputs(3030) <= (layer3_outputs(4422)) or (layer3_outputs(2694));
    layer4_outputs(3031) <= (layer3_outputs(3393)) xor (layer3_outputs(432));
    layer4_outputs(3032) <= (layer3_outputs(3791)) and not (layer3_outputs(8279));
    layer4_outputs(3033) <= not((layer3_outputs(1484)) xor (layer3_outputs(6295)));
    layer4_outputs(3034) <= not((layer3_outputs(5039)) and (layer3_outputs(4001)));
    layer4_outputs(3035) <= (layer3_outputs(7190)) xor (layer3_outputs(3490));
    layer4_outputs(3036) <= (layer3_outputs(3407)) and not (layer3_outputs(8990));
    layer4_outputs(3037) <= not(layer3_outputs(9425)) or (layer3_outputs(5830));
    layer4_outputs(3038) <= not((layer3_outputs(4199)) xor (layer3_outputs(887)));
    layer4_outputs(3039) <= not((layer3_outputs(8146)) xor (layer3_outputs(453)));
    layer4_outputs(3040) <= layer3_outputs(5189);
    layer4_outputs(3041) <= not(layer3_outputs(8349));
    layer4_outputs(3042) <= not((layer3_outputs(7099)) and (layer3_outputs(4961)));
    layer4_outputs(3043) <= layer3_outputs(5891);
    layer4_outputs(3044) <= not(layer3_outputs(995)) or (layer3_outputs(8611));
    layer4_outputs(3045) <= not(layer3_outputs(6543)) or (layer3_outputs(7931));
    layer4_outputs(3046) <= (layer3_outputs(9539)) xor (layer3_outputs(6037));
    layer4_outputs(3047) <= (layer3_outputs(7501)) xor (layer3_outputs(6779));
    layer4_outputs(3048) <= not(layer3_outputs(8694));
    layer4_outputs(3049) <= (layer3_outputs(3738)) xor (layer3_outputs(55));
    layer4_outputs(3050) <= layer3_outputs(3900);
    layer4_outputs(3051) <= layer3_outputs(9710);
    layer4_outputs(3052) <= layer3_outputs(1775);
    layer4_outputs(3053) <= (layer3_outputs(5815)) and (layer3_outputs(3739));
    layer4_outputs(3054) <= not(layer3_outputs(560));
    layer4_outputs(3055) <= not((layer3_outputs(3259)) and (layer3_outputs(6249)));
    layer4_outputs(3056) <= not(layer3_outputs(3446));
    layer4_outputs(3057) <= layer3_outputs(4421);
    layer4_outputs(3058) <= not(layer3_outputs(1546));
    layer4_outputs(3059) <= layer3_outputs(9974);
    layer4_outputs(3060) <= (layer3_outputs(6581)) xor (layer3_outputs(7198));
    layer4_outputs(3061) <= not(layer3_outputs(786));
    layer4_outputs(3062) <= not(layer3_outputs(8846));
    layer4_outputs(3063) <= '1';
    layer4_outputs(3064) <= layer3_outputs(5964);
    layer4_outputs(3065) <= not((layer3_outputs(5739)) xor (layer3_outputs(9510)));
    layer4_outputs(3066) <= not(layer3_outputs(4736));
    layer4_outputs(3067) <= not(layer3_outputs(4551));
    layer4_outputs(3068) <= (layer3_outputs(1255)) xor (layer3_outputs(8631));
    layer4_outputs(3069) <= (layer3_outputs(506)) and not (layer3_outputs(1723));
    layer4_outputs(3070) <= not(layer3_outputs(528));
    layer4_outputs(3071) <= (layer3_outputs(8195)) and not (layer3_outputs(5149));
    layer4_outputs(3072) <= layer3_outputs(3578);
    layer4_outputs(3073) <= not(layer3_outputs(5602)) or (layer3_outputs(5317));
    layer4_outputs(3074) <= not(layer3_outputs(3855));
    layer4_outputs(3075) <= not((layer3_outputs(1793)) or (layer3_outputs(7330)));
    layer4_outputs(3076) <= not(layer3_outputs(2120));
    layer4_outputs(3077) <= not(layer3_outputs(3172));
    layer4_outputs(3078) <= not(layer3_outputs(9256));
    layer4_outputs(3079) <= layer3_outputs(7905);
    layer4_outputs(3080) <= not(layer3_outputs(2135));
    layer4_outputs(3081) <= not((layer3_outputs(2954)) and (layer3_outputs(3685)));
    layer4_outputs(3082) <= (layer3_outputs(8109)) and not (layer3_outputs(9332));
    layer4_outputs(3083) <= not(layer3_outputs(5500));
    layer4_outputs(3084) <= not(layer3_outputs(620)) or (layer3_outputs(6825));
    layer4_outputs(3085) <= layer3_outputs(7995);
    layer4_outputs(3086) <= not(layer3_outputs(1451));
    layer4_outputs(3087) <= not(layer3_outputs(9125));
    layer4_outputs(3088) <= layer3_outputs(3189);
    layer4_outputs(3089) <= layer3_outputs(3256);
    layer4_outputs(3090) <= not(layer3_outputs(5757));
    layer4_outputs(3091) <= layer3_outputs(10094);
    layer4_outputs(3092) <= layer3_outputs(8008);
    layer4_outputs(3093) <= not((layer3_outputs(5641)) xor (layer3_outputs(3646)));
    layer4_outputs(3094) <= not(layer3_outputs(2247));
    layer4_outputs(3095) <= layer3_outputs(2072);
    layer4_outputs(3096) <= layer3_outputs(7095);
    layer4_outputs(3097) <= not((layer3_outputs(1275)) or (layer3_outputs(4183)));
    layer4_outputs(3098) <= layer3_outputs(8489);
    layer4_outputs(3099) <= layer3_outputs(5733);
    layer4_outputs(3100) <= not((layer3_outputs(2949)) xor (layer3_outputs(3134)));
    layer4_outputs(3101) <= layer3_outputs(8741);
    layer4_outputs(3102) <= not(layer3_outputs(7991));
    layer4_outputs(3103) <= not(layer3_outputs(9374));
    layer4_outputs(3104) <= (layer3_outputs(2035)) and (layer3_outputs(1955));
    layer4_outputs(3105) <= not(layer3_outputs(1752));
    layer4_outputs(3106) <= (layer3_outputs(5035)) xor (layer3_outputs(7895));
    layer4_outputs(3107) <= not(layer3_outputs(8472));
    layer4_outputs(3108) <= layer3_outputs(7231);
    layer4_outputs(3109) <= (layer3_outputs(6727)) xor (layer3_outputs(8724));
    layer4_outputs(3110) <= layer3_outputs(9060);
    layer4_outputs(3111) <= layer3_outputs(4794);
    layer4_outputs(3112) <= layer3_outputs(2781);
    layer4_outputs(3113) <= layer3_outputs(9450);
    layer4_outputs(3114) <= not(layer3_outputs(10068));
    layer4_outputs(3115) <= not((layer3_outputs(946)) xor (layer3_outputs(3597)));
    layer4_outputs(3116) <= (layer3_outputs(8460)) and not (layer3_outputs(4298));
    layer4_outputs(3117) <= layer3_outputs(4552);
    layer4_outputs(3118) <= layer3_outputs(1318);
    layer4_outputs(3119) <= not((layer3_outputs(4192)) and (layer3_outputs(6253)));
    layer4_outputs(3120) <= not((layer3_outputs(7425)) xor (layer3_outputs(4782)));
    layer4_outputs(3121) <= '1';
    layer4_outputs(3122) <= not(layer3_outputs(4964));
    layer4_outputs(3123) <= not(layer3_outputs(1764));
    layer4_outputs(3124) <= not((layer3_outputs(4883)) and (layer3_outputs(8476)));
    layer4_outputs(3125) <= layer3_outputs(6966);
    layer4_outputs(3126) <= (layer3_outputs(1959)) xor (layer3_outputs(4986));
    layer4_outputs(3127) <= not(layer3_outputs(9568));
    layer4_outputs(3128) <= not(layer3_outputs(3818));
    layer4_outputs(3129) <= layer3_outputs(9206);
    layer4_outputs(3130) <= layer3_outputs(3137);
    layer4_outputs(3131) <= layer3_outputs(3086);
    layer4_outputs(3132) <= layer3_outputs(2393);
    layer4_outputs(3133) <= layer3_outputs(3116);
    layer4_outputs(3134) <= not(layer3_outputs(584));
    layer4_outputs(3135) <= layer3_outputs(6851);
    layer4_outputs(3136) <= not(layer3_outputs(5609));
    layer4_outputs(3137) <= layer3_outputs(2994);
    layer4_outputs(3138) <= layer3_outputs(9468);
    layer4_outputs(3139) <= layer3_outputs(6742);
    layer4_outputs(3140) <= not(layer3_outputs(4136));
    layer4_outputs(3141) <= layer3_outputs(3983);
    layer4_outputs(3142) <= (layer3_outputs(9652)) and (layer3_outputs(8433));
    layer4_outputs(3143) <= (layer3_outputs(4929)) or (layer3_outputs(2999));
    layer4_outputs(3144) <= not(layer3_outputs(8286));
    layer4_outputs(3145) <= (layer3_outputs(4673)) and not (layer3_outputs(2975));
    layer4_outputs(3146) <= not(layer3_outputs(5563));
    layer4_outputs(3147) <= layer3_outputs(1391);
    layer4_outputs(3148) <= not((layer3_outputs(3174)) xor (layer3_outputs(96)));
    layer4_outputs(3149) <= not((layer3_outputs(8893)) xor (layer3_outputs(122)));
    layer4_outputs(3150) <= layer3_outputs(552);
    layer4_outputs(3151) <= not(layer3_outputs(805)) or (layer3_outputs(3995));
    layer4_outputs(3152) <= not(layer3_outputs(8727));
    layer4_outputs(3153) <= not(layer3_outputs(10231));
    layer4_outputs(3154) <= not(layer3_outputs(6815));
    layer4_outputs(3155) <= not(layer3_outputs(4063));
    layer4_outputs(3156) <= layer3_outputs(5235);
    layer4_outputs(3157) <= (layer3_outputs(8607)) and (layer3_outputs(5170));
    layer4_outputs(3158) <= (layer3_outputs(363)) or (layer3_outputs(5147));
    layer4_outputs(3159) <= (layer3_outputs(4116)) xor (layer3_outputs(5019));
    layer4_outputs(3160) <= not(layer3_outputs(8735)) or (layer3_outputs(7159));
    layer4_outputs(3161) <= not((layer3_outputs(8112)) xor (layer3_outputs(9059)));
    layer4_outputs(3162) <= not(layer3_outputs(8620)) or (layer3_outputs(6046));
    layer4_outputs(3163) <= (layer3_outputs(6344)) or (layer3_outputs(6194));
    layer4_outputs(3164) <= not((layer3_outputs(9423)) xor (layer3_outputs(5411)));
    layer4_outputs(3165) <= (layer3_outputs(10158)) or (layer3_outputs(7418));
    layer4_outputs(3166) <= layer3_outputs(1527);
    layer4_outputs(3167) <= layer3_outputs(3016);
    layer4_outputs(3168) <= not(layer3_outputs(2755));
    layer4_outputs(3169) <= not(layer3_outputs(4092));
    layer4_outputs(3170) <= not(layer3_outputs(2014));
    layer4_outputs(3171) <= not(layer3_outputs(218));
    layer4_outputs(3172) <= not(layer3_outputs(2167));
    layer4_outputs(3173) <= layer3_outputs(1845);
    layer4_outputs(3174) <= (layer3_outputs(6683)) xor (layer3_outputs(7568));
    layer4_outputs(3175) <= not(layer3_outputs(9507));
    layer4_outputs(3176) <= (layer3_outputs(1097)) and (layer3_outputs(7432));
    layer4_outputs(3177) <= not((layer3_outputs(2296)) xor (layer3_outputs(1818)));
    layer4_outputs(3178) <= layer3_outputs(7848);
    layer4_outputs(3179) <= not(layer3_outputs(7959));
    layer4_outputs(3180) <= not((layer3_outputs(7315)) xor (layer3_outputs(4337)));
    layer4_outputs(3181) <= not(layer3_outputs(8959));
    layer4_outputs(3182) <= layer3_outputs(9954);
    layer4_outputs(3183) <= not(layer3_outputs(5242));
    layer4_outputs(3184) <= not(layer3_outputs(741));
    layer4_outputs(3185) <= not(layer3_outputs(10013));
    layer4_outputs(3186) <= layer3_outputs(3447);
    layer4_outputs(3187) <= not((layer3_outputs(6670)) or (layer3_outputs(5834)));
    layer4_outputs(3188) <= not(layer3_outputs(5000)) or (layer3_outputs(578));
    layer4_outputs(3189) <= (layer3_outputs(7740)) and not (layer3_outputs(1398));
    layer4_outputs(3190) <= (layer3_outputs(209)) and (layer3_outputs(1416));
    layer4_outputs(3191) <= '0';
    layer4_outputs(3192) <= layer3_outputs(3980);
    layer4_outputs(3193) <= not((layer3_outputs(3144)) xor (layer3_outputs(6485)));
    layer4_outputs(3194) <= not(layer3_outputs(705));
    layer4_outputs(3195) <= (layer3_outputs(10238)) or (layer3_outputs(7053));
    layer4_outputs(3196) <= layer3_outputs(3878);
    layer4_outputs(3197) <= layer3_outputs(1919);
    layer4_outputs(3198) <= (layer3_outputs(9794)) or (layer3_outputs(202));
    layer4_outputs(3199) <= not(layer3_outputs(8798));
    layer4_outputs(3200) <= not(layer3_outputs(7924));
    layer4_outputs(3201) <= (layer3_outputs(8009)) and not (layer3_outputs(1179));
    layer4_outputs(3202) <= not((layer3_outputs(696)) and (layer3_outputs(3702)));
    layer4_outputs(3203) <= layer3_outputs(6156);
    layer4_outputs(3204) <= not(layer3_outputs(4818));
    layer4_outputs(3205) <= not(layer3_outputs(7257));
    layer4_outputs(3206) <= not((layer3_outputs(4541)) xor (layer3_outputs(1116)));
    layer4_outputs(3207) <= not(layer3_outputs(4573));
    layer4_outputs(3208) <= not(layer3_outputs(4604));
    layer4_outputs(3209) <= not(layer3_outputs(8672));
    layer4_outputs(3210) <= layer3_outputs(1208);
    layer4_outputs(3211) <= layer3_outputs(5064);
    layer4_outputs(3212) <= layer3_outputs(6213);
    layer4_outputs(3213) <= (layer3_outputs(2519)) and (layer3_outputs(1661));
    layer4_outputs(3214) <= not((layer3_outputs(4053)) and (layer3_outputs(6138)));
    layer4_outputs(3215) <= layer3_outputs(9885);
    layer4_outputs(3216) <= not(layer3_outputs(3996));
    layer4_outputs(3217) <= not(layer3_outputs(9261));
    layer4_outputs(3218) <= (layer3_outputs(10206)) and not (layer3_outputs(5738));
    layer4_outputs(3219) <= not(layer3_outputs(9707));
    layer4_outputs(3220) <= layer3_outputs(3921);
    layer4_outputs(3221) <= layer3_outputs(7636);
    layer4_outputs(3222) <= not((layer3_outputs(271)) or (layer3_outputs(7359)));
    layer4_outputs(3223) <= not(layer3_outputs(6072));
    layer4_outputs(3224) <= layer3_outputs(6908);
    layer4_outputs(3225) <= layer3_outputs(9338);
    layer4_outputs(3226) <= (layer3_outputs(9739)) xor (layer3_outputs(6752));
    layer4_outputs(3227) <= not(layer3_outputs(2622));
    layer4_outputs(3228) <= layer3_outputs(1238);
    layer4_outputs(3229) <= not(layer3_outputs(7831));
    layer4_outputs(3230) <= (layer3_outputs(6435)) or (layer3_outputs(4019));
    layer4_outputs(3231) <= not(layer3_outputs(7193));
    layer4_outputs(3232) <= layer3_outputs(6657);
    layer4_outputs(3233) <= not(layer3_outputs(6090));
    layer4_outputs(3234) <= layer3_outputs(8640);
    layer4_outputs(3235) <= not((layer3_outputs(1324)) and (layer3_outputs(9618)));
    layer4_outputs(3236) <= (layer3_outputs(439)) xor (layer3_outputs(10129));
    layer4_outputs(3237) <= not(layer3_outputs(5839));
    layer4_outputs(3238) <= not(layer3_outputs(3346)) or (layer3_outputs(5793));
    layer4_outputs(3239) <= not(layer3_outputs(2023));
    layer4_outputs(3240) <= (layer3_outputs(5094)) and not (layer3_outputs(317));
    layer4_outputs(3241) <= not(layer3_outputs(6620));
    layer4_outputs(3242) <= not((layer3_outputs(9717)) and (layer3_outputs(6278)));
    layer4_outputs(3243) <= (layer3_outputs(1320)) xor (layer3_outputs(4536));
    layer4_outputs(3244) <= '1';
    layer4_outputs(3245) <= layer3_outputs(7131);
    layer4_outputs(3246) <= not(layer3_outputs(8409)) or (layer3_outputs(7773));
    layer4_outputs(3247) <= not(layer3_outputs(6691));
    layer4_outputs(3248) <= not((layer3_outputs(8013)) xor (layer3_outputs(4583)));
    layer4_outputs(3249) <= not(layer3_outputs(1771));
    layer4_outputs(3250) <= not(layer3_outputs(7789)) or (layer3_outputs(267));
    layer4_outputs(3251) <= not((layer3_outputs(1730)) and (layer3_outputs(6989)));
    layer4_outputs(3252) <= layer3_outputs(6813);
    layer4_outputs(3253) <= not(layer3_outputs(5919));
    layer4_outputs(3254) <= (layer3_outputs(8315)) and (layer3_outputs(4635));
    layer4_outputs(3255) <= not(layer3_outputs(5807));
    layer4_outputs(3256) <= not(layer3_outputs(1068));
    layer4_outputs(3257) <= (layer3_outputs(825)) and (layer3_outputs(9387));
    layer4_outputs(3258) <= not(layer3_outputs(8713));
    layer4_outputs(3259) <= (layer3_outputs(4058)) xor (layer3_outputs(9459));
    layer4_outputs(3260) <= (layer3_outputs(1065)) or (layer3_outputs(9551));
    layer4_outputs(3261) <= not(layer3_outputs(5599));
    layer4_outputs(3262) <= layer3_outputs(2233);
    layer4_outputs(3263) <= layer3_outputs(2680);
    layer4_outputs(3264) <= (layer3_outputs(6815)) or (layer3_outputs(857));
    layer4_outputs(3265) <= not(layer3_outputs(6513));
    layer4_outputs(3266) <= (layer3_outputs(7633)) xor (layer3_outputs(7705));
    layer4_outputs(3267) <= layer3_outputs(639);
    layer4_outputs(3268) <= layer3_outputs(3560);
    layer4_outputs(3269) <= (layer3_outputs(2796)) or (layer3_outputs(7822));
    layer4_outputs(3270) <= not(layer3_outputs(9203));
    layer4_outputs(3271) <= not((layer3_outputs(5772)) xor (layer3_outputs(8006)));
    layer4_outputs(3272) <= (layer3_outputs(8729)) and not (layer3_outputs(6360));
    layer4_outputs(3273) <= (layer3_outputs(2665)) or (layer3_outputs(9616));
    layer4_outputs(3274) <= layer3_outputs(7359);
    layer4_outputs(3275) <= layer3_outputs(2472);
    layer4_outputs(3276) <= not(layer3_outputs(9737));
    layer4_outputs(3277) <= layer3_outputs(7983);
    layer4_outputs(3278) <= not(layer3_outputs(5918));
    layer4_outputs(3279) <= not(layer3_outputs(10187));
    layer4_outputs(3280) <= not((layer3_outputs(5504)) and (layer3_outputs(6019)));
    layer4_outputs(3281) <= layer3_outputs(5383);
    layer4_outputs(3282) <= layer3_outputs(7694);
    layer4_outputs(3283) <= not(layer3_outputs(7204));
    layer4_outputs(3284) <= (layer3_outputs(2091)) and not (layer3_outputs(2641));
    layer4_outputs(3285) <= not(layer3_outputs(65));
    layer4_outputs(3286) <= (layer3_outputs(5721)) xor (layer3_outputs(6494));
    layer4_outputs(3287) <= not((layer3_outputs(2364)) xor (layer3_outputs(8358)));
    layer4_outputs(3288) <= not(layer3_outputs(8196)) or (layer3_outputs(1361));
    layer4_outputs(3289) <= layer3_outputs(2895);
    layer4_outputs(3290) <= (layer3_outputs(1608)) xor (layer3_outputs(6344));
    layer4_outputs(3291) <= (layer3_outputs(2576)) xor (layer3_outputs(27));
    layer4_outputs(3292) <= layer3_outputs(4578);
    layer4_outputs(3293) <= not(layer3_outputs(7894)) or (layer3_outputs(9320));
    layer4_outputs(3294) <= layer3_outputs(8900);
    layer4_outputs(3295) <= not((layer3_outputs(3810)) and (layer3_outputs(8722)));
    layer4_outputs(3296) <= not(layer3_outputs(6298));
    layer4_outputs(3297) <= not((layer3_outputs(3649)) xor (layer3_outputs(996)));
    layer4_outputs(3298) <= not(layer3_outputs(2535));
    layer4_outputs(3299) <= not(layer3_outputs(7306)) or (layer3_outputs(744));
    layer4_outputs(3300) <= not(layer3_outputs(8412));
    layer4_outputs(3301) <= layer3_outputs(1493);
    layer4_outputs(3302) <= not((layer3_outputs(8605)) and (layer3_outputs(3690)));
    layer4_outputs(3303) <= not(layer3_outputs(5767)) or (layer3_outputs(6386));
    layer4_outputs(3304) <= not(layer3_outputs(6620));
    layer4_outputs(3305) <= layer3_outputs(2144);
    layer4_outputs(3306) <= layer3_outputs(7238);
    layer4_outputs(3307) <= layer3_outputs(7941);
    layer4_outputs(3308) <= (layer3_outputs(7753)) xor (layer3_outputs(1558));
    layer4_outputs(3309) <= not(layer3_outputs(6429));
    layer4_outputs(3310) <= (layer3_outputs(5210)) or (layer3_outputs(5964));
    layer4_outputs(3311) <= not((layer3_outputs(52)) xor (layer3_outputs(3154)));
    layer4_outputs(3312) <= (layer3_outputs(8067)) and not (layer3_outputs(5435));
    layer4_outputs(3313) <= (layer3_outputs(4515)) and not (layer3_outputs(6342));
    layer4_outputs(3314) <= not(layer3_outputs(4830));
    layer4_outputs(3315) <= layer3_outputs(1352);
    layer4_outputs(3316) <= not(layer3_outputs(5613));
    layer4_outputs(3317) <= layer3_outputs(8329);
    layer4_outputs(3318) <= not(layer3_outputs(1581));
    layer4_outputs(3319) <= layer3_outputs(2466);
    layer4_outputs(3320) <= not((layer3_outputs(4328)) or (layer3_outputs(1202)));
    layer4_outputs(3321) <= '0';
    layer4_outputs(3322) <= (layer3_outputs(7047)) or (layer3_outputs(8855));
    layer4_outputs(3323) <= (layer3_outputs(2173)) and not (layer3_outputs(8109));
    layer4_outputs(3324) <= not((layer3_outputs(2195)) or (layer3_outputs(1300)));
    layer4_outputs(3325) <= (layer3_outputs(1255)) and (layer3_outputs(9430));
    layer4_outputs(3326) <= not(layer3_outputs(746));
    layer4_outputs(3327) <= not((layer3_outputs(7184)) or (layer3_outputs(580)));
    layer4_outputs(3328) <= (layer3_outputs(6806)) and not (layer3_outputs(6851));
    layer4_outputs(3329) <= layer3_outputs(41);
    layer4_outputs(3330) <= not(layer3_outputs(6221)) or (layer3_outputs(6962));
    layer4_outputs(3331) <= (layer3_outputs(6545)) and (layer3_outputs(8659));
    layer4_outputs(3332) <= not(layer3_outputs(3381));
    layer4_outputs(3333) <= layer3_outputs(8690);
    layer4_outputs(3334) <= layer3_outputs(7782);
    layer4_outputs(3335) <= not(layer3_outputs(3835));
    layer4_outputs(3336) <= layer3_outputs(3635);
    layer4_outputs(3337) <= (layer3_outputs(1720)) xor (layer3_outputs(1328));
    layer4_outputs(3338) <= layer3_outputs(4557);
    layer4_outputs(3339) <= (layer3_outputs(2930)) xor (layer3_outputs(108));
    layer4_outputs(3340) <= not(layer3_outputs(6375));
    layer4_outputs(3341) <= layer3_outputs(3967);
    layer4_outputs(3342) <= not(layer3_outputs(5012));
    layer4_outputs(3343) <= not(layer3_outputs(9616));
    layer4_outputs(3344) <= not((layer3_outputs(5465)) and (layer3_outputs(2424)));
    layer4_outputs(3345) <= not((layer3_outputs(9032)) or (layer3_outputs(10090)));
    layer4_outputs(3346) <= layer3_outputs(5283);
    layer4_outputs(3347) <= layer3_outputs(8323);
    layer4_outputs(3348) <= '1';
    layer4_outputs(3349) <= not((layer3_outputs(3621)) xor (layer3_outputs(6863)));
    layer4_outputs(3350) <= not(layer3_outputs(855));
    layer4_outputs(3351) <= not(layer3_outputs(6438)) or (layer3_outputs(5620));
    layer4_outputs(3352) <= not(layer3_outputs(5832));
    layer4_outputs(3353) <= not(layer3_outputs(6635));
    layer4_outputs(3354) <= not(layer3_outputs(3354));
    layer4_outputs(3355) <= layer3_outputs(4777);
    layer4_outputs(3356) <= layer3_outputs(10092);
    layer4_outputs(3357) <= '0';
    layer4_outputs(3358) <= layer3_outputs(264);
    layer4_outputs(3359) <= not(layer3_outputs(3071));
    layer4_outputs(3360) <= not(layer3_outputs(1009)) or (layer3_outputs(352));
    layer4_outputs(3361) <= (layer3_outputs(4475)) and not (layer3_outputs(8101));
    layer4_outputs(3362) <= layer3_outputs(7259);
    layer4_outputs(3363) <= not((layer3_outputs(688)) xor (layer3_outputs(7329)));
    layer4_outputs(3364) <= (layer3_outputs(763)) or (layer3_outputs(1180));
    layer4_outputs(3365) <= (layer3_outputs(1566)) or (layer3_outputs(4974));
    layer4_outputs(3366) <= not((layer3_outputs(2861)) xor (layer3_outputs(4892)));
    layer4_outputs(3367) <= layer3_outputs(10101);
    layer4_outputs(3368) <= (layer3_outputs(1622)) xor (layer3_outputs(3595));
    layer4_outputs(3369) <= '0';
    layer4_outputs(3370) <= (layer3_outputs(916)) and not (layer3_outputs(4685));
    layer4_outputs(3371) <= (layer3_outputs(1876)) xor (layer3_outputs(8059));
    layer4_outputs(3372) <= (layer3_outputs(10117)) and not (layer3_outputs(9131));
    layer4_outputs(3373) <= layer3_outputs(8133);
    layer4_outputs(3374) <= not(layer3_outputs(4448)) or (layer3_outputs(4509));
    layer4_outputs(3375) <= (layer3_outputs(214)) and not (layer3_outputs(4008));
    layer4_outputs(3376) <= not(layer3_outputs(647)) or (layer3_outputs(9674));
    layer4_outputs(3377) <= not((layer3_outputs(3100)) xor (layer3_outputs(795)));
    layer4_outputs(3378) <= not(layer3_outputs(9517)) or (layer3_outputs(813));
    layer4_outputs(3379) <= not(layer3_outputs(6153));
    layer4_outputs(3380) <= layer3_outputs(2890);
    layer4_outputs(3381) <= not(layer3_outputs(3292)) or (layer3_outputs(6538));
    layer4_outputs(3382) <= layer3_outputs(3990);
    layer4_outputs(3383) <= not(layer3_outputs(2200));
    layer4_outputs(3384) <= not(layer3_outputs(4739));
    layer4_outputs(3385) <= not(layer3_outputs(6153));
    layer4_outputs(3386) <= (layer3_outputs(2045)) xor (layer3_outputs(2727));
    layer4_outputs(3387) <= not((layer3_outputs(4538)) xor (layer3_outputs(1823)));
    layer4_outputs(3388) <= not(layer3_outputs(2430));
    layer4_outputs(3389) <= not(layer3_outputs(1980));
    layer4_outputs(3390) <= '1';
    layer4_outputs(3391) <= not(layer3_outputs(5267)) or (layer3_outputs(10009));
    layer4_outputs(3392) <= not(layer3_outputs(2978)) or (layer3_outputs(2895));
    layer4_outputs(3393) <= layer3_outputs(6840);
    layer4_outputs(3394) <= not((layer3_outputs(1543)) and (layer3_outputs(7992)));
    layer4_outputs(3395) <= not(layer3_outputs(4027));
    layer4_outputs(3396) <= not((layer3_outputs(1487)) or (layer3_outputs(6546)));
    layer4_outputs(3397) <= not((layer3_outputs(6589)) and (layer3_outputs(2278)));
    layer4_outputs(3398) <= not(layer3_outputs(7444));
    layer4_outputs(3399) <= layer3_outputs(561);
    layer4_outputs(3400) <= layer3_outputs(5266);
    layer4_outputs(3401) <= not(layer3_outputs(4467)) or (layer3_outputs(1822));
    layer4_outputs(3402) <= not(layer3_outputs(5195));
    layer4_outputs(3403) <= (layer3_outputs(7956)) and (layer3_outputs(2221));
    layer4_outputs(3404) <= layer3_outputs(6007);
    layer4_outputs(3405) <= layer3_outputs(645);
    layer4_outputs(3406) <= not(layer3_outputs(9370));
    layer4_outputs(3407) <= not((layer3_outputs(1783)) xor (layer3_outputs(602)));
    layer4_outputs(3408) <= not((layer3_outputs(8380)) xor (layer3_outputs(4790)));
    layer4_outputs(3409) <= (layer3_outputs(10234)) and not (layer3_outputs(464));
    layer4_outputs(3410) <= not(layer3_outputs(2261));
    layer4_outputs(3411) <= not(layer3_outputs(10132));
    layer4_outputs(3412) <= (layer3_outputs(2247)) xor (layer3_outputs(6532));
    layer4_outputs(3413) <= not(layer3_outputs(381));
    layer4_outputs(3414) <= (layer3_outputs(3852)) or (layer3_outputs(9868));
    layer4_outputs(3415) <= (layer3_outputs(2771)) and not (layer3_outputs(3237));
    layer4_outputs(3416) <= (layer3_outputs(921)) and (layer3_outputs(7283));
    layer4_outputs(3417) <= not(layer3_outputs(207));
    layer4_outputs(3418) <= layer3_outputs(2165);
    layer4_outputs(3419) <= not(layer3_outputs(1634));
    layer4_outputs(3420) <= not(layer3_outputs(6612));
    layer4_outputs(3421) <= not((layer3_outputs(2420)) and (layer3_outputs(2299)));
    layer4_outputs(3422) <= not(layer3_outputs(8183));
    layer4_outputs(3423) <= not(layer3_outputs(745)) or (layer3_outputs(5255));
    layer4_outputs(3424) <= not((layer3_outputs(247)) and (layer3_outputs(3630)));
    layer4_outputs(3425) <= not((layer3_outputs(1935)) or (layer3_outputs(421)));
    layer4_outputs(3426) <= not(layer3_outputs(7));
    layer4_outputs(3427) <= not((layer3_outputs(7982)) xor (layer3_outputs(4450)));
    layer4_outputs(3428) <= (layer3_outputs(2471)) and not (layer3_outputs(8926));
    layer4_outputs(3429) <= (layer3_outputs(7420)) or (layer3_outputs(9082));
    layer4_outputs(3430) <= not((layer3_outputs(4131)) or (layer3_outputs(8373)));
    layer4_outputs(3431) <= not(layer3_outputs(2848));
    layer4_outputs(3432) <= not(layer3_outputs(380));
    layer4_outputs(3433) <= not((layer3_outputs(911)) xor (layer3_outputs(91)));
    layer4_outputs(3434) <= not(layer3_outputs(3253));
    layer4_outputs(3435) <= layer3_outputs(5830);
    layer4_outputs(3436) <= (layer3_outputs(5570)) and (layer3_outputs(6243));
    layer4_outputs(3437) <= (layer3_outputs(9807)) and (layer3_outputs(7217));
    layer4_outputs(3438) <= not((layer3_outputs(1838)) xor (layer3_outputs(1191)));
    layer4_outputs(3439) <= layer3_outputs(2199);
    layer4_outputs(3440) <= not(layer3_outputs(9159));
    layer4_outputs(3441) <= (layer3_outputs(610)) and not (layer3_outputs(4284));
    layer4_outputs(3442) <= not(layer3_outputs(4456)) or (layer3_outputs(978));
    layer4_outputs(3443) <= layer3_outputs(2056);
    layer4_outputs(3444) <= layer3_outputs(1870);
    layer4_outputs(3445) <= not(layer3_outputs(928));
    layer4_outputs(3446) <= not((layer3_outputs(4098)) or (layer3_outputs(5244)));
    layer4_outputs(3447) <= not(layer3_outputs(8379));
    layer4_outputs(3448) <= layer3_outputs(8680);
    layer4_outputs(3449) <= layer3_outputs(456);
    layer4_outputs(3450) <= not(layer3_outputs(2765));
    layer4_outputs(3451) <= not((layer3_outputs(10126)) or (layer3_outputs(9605)));
    layer4_outputs(3452) <= layer3_outputs(8123);
    layer4_outputs(3453) <= (layer3_outputs(1789)) or (layer3_outputs(4893));
    layer4_outputs(3454) <= (layer3_outputs(7446)) or (layer3_outputs(1011));
    layer4_outputs(3455) <= not(layer3_outputs(9736));
    layer4_outputs(3456) <= not((layer3_outputs(6504)) and (layer3_outputs(7)));
    layer4_outputs(3457) <= (layer3_outputs(8207)) xor (layer3_outputs(5596));
    layer4_outputs(3458) <= '1';
    layer4_outputs(3459) <= (layer3_outputs(4695)) or (layer3_outputs(6631));
    layer4_outputs(3460) <= layer3_outputs(7107);
    layer4_outputs(3461) <= not(layer3_outputs(1520));
    layer4_outputs(3462) <= layer3_outputs(5916);
    layer4_outputs(3463) <= layer3_outputs(9923);
    layer4_outputs(3464) <= layer3_outputs(7193);
    layer4_outputs(3465) <= not((layer3_outputs(8324)) or (layer3_outputs(9050)));
    layer4_outputs(3466) <= (layer3_outputs(2211)) xor (layer3_outputs(9820));
    layer4_outputs(3467) <= not(layer3_outputs(2706));
    layer4_outputs(3468) <= not((layer3_outputs(9600)) xor (layer3_outputs(983)));
    layer4_outputs(3469) <= layer3_outputs(2721);
    layer4_outputs(3470) <= layer3_outputs(4759);
    layer4_outputs(3471) <= (layer3_outputs(6791)) xor (layer3_outputs(2478));
    layer4_outputs(3472) <= (layer3_outputs(5600)) and (layer3_outputs(7228));
    layer4_outputs(3473) <= not(layer3_outputs(5743));
    layer4_outputs(3474) <= layer3_outputs(1127);
    layer4_outputs(3475) <= (layer3_outputs(4555)) xor (layer3_outputs(9253));
    layer4_outputs(3476) <= not((layer3_outputs(1417)) or (layer3_outputs(2779)));
    layer4_outputs(3477) <= not(layer3_outputs(9439));
    layer4_outputs(3478) <= layer3_outputs(4989);
    layer4_outputs(3479) <= not(layer3_outputs(1280));
    layer4_outputs(3480) <= (layer3_outputs(2333)) and (layer3_outputs(2617));
    layer4_outputs(3481) <= (layer3_outputs(1952)) and not (layer3_outputs(8890));
    layer4_outputs(3482) <= not((layer3_outputs(2419)) or (layer3_outputs(9045)));
    layer4_outputs(3483) <= not((layer3_outputs(3871)) or (layer3_outputs(6058)));
    layer4_outputs(3484) <= not((layer3_outputs(8348)) or (layer3_outputs(9947)));
    layer4_outputs(3485) <= layer3_outputs(7502);
    layer4_outputs(3486) <= '1';
    layer4_outputs(3487) <= not((layer3_outputs(4492)) and (layer3_outputs(5850)));
    layer4_outputs(3488) <= not((layer3_outputs(6756)) or (layer3_outputs(9353)));
    layer4_outputs(3489) <= not(layer3_outputs(4835)) or (layer3_outputs(6034));
    layer4_outputs(3490) <= layer3_outputs(6936);
    layer4_outputs(3491) <= not(layer3_outputs(7508));
    layer4_outputs(3492) <= layer3_outputs(9631);
    layer4_outputs(3493) <= not(layer3_outputs(6849)) or (layer3_outputs(152));
    layer4_outputs(3494) <= not((layer3_outputs(5245)) xor (layer3_outputs(8419)));
    layer4_outputs(3495) <= not(layer3_outputs(8237));
    layer4_outputs(3496) <= not((layer3_outputs(4397)) and (layer3_outputs(1630)));
    layer4_outputs(3497) <= not(layer3_outputs(5473));
    layer4_outputs(3498) <= layer3_outputs(6770);
    layer4_outputs(3499) <= (layer3_outputs(7969)) xor (layer3_outputs(6685));
    layer4_outputs(3500) <= (layer3_outputs(621)) or (layer3_outputs(9213));
    layer4_outputs(3501) <= '1';
    layer4_outputs(3502) <= not(layer3_outputs(6323));
    layer4_outputs(3503) <= not(layer3_outputs(6137));
    layer4_outputs(3504) <= not((layer3_outputs(7293)) or (layer3_outputs(6027)));
    layer4_outputs(3505) <= layer3_outputs(6810);
    layer4_outputs(3506) <= (layer3_outputs(3243)) and (layer3_outputs(7793));
    layer4_outputs(3507) <= layer3_outputs(3432);
    layer4_outputs(3508) <= not(layer3_outputs(8868));
    layer4_outputs(3509) <= layer3_outputs(1904);
    layer4_outputs(3510) <= (layer3_outputs(6677)) and not (layer3_outputs(6526));
    layer4_outputs(3511) <= layer3_outputs(2773);
    layer4_outputs(3512) <= (layer3_outputs(3169)) xor (layer3_outputs(1210));
    layer4_outputs(3513) <= layer3_outputs(10191);
    layer4_outputs(3514) <= not(layer3_outputs(9832));
    layer4_outputs(3515) <= (layer3_outputs(4665)) xor (layer3_outputs(2262));
    layer4_outputs(3516) <= not(layer3_outputs(2128));
    layer4_outputs(3517) <= (layer3_outputs(7367)) xor (layer3_outputs(9392));
    layer4_outputs(3518) <= not((layer3_outputs(2892)) xor (layer3_outputs(1359)));
    layer4_outputs(3519) <= layer3_outputs(7843);
    layer4_outputs(3520) <= layer3_outputs(6660);
    layer4_outputs(3521) <= layer3_outputs(5345);
    layer4_outputs(3522) <= layer3_outputs(3531);
    layer4_outputs(3523) <= not(layer3_outputs(9526));
    layer4_outputs(3524) <= not(layer3_outputs(7935));
    layer4_outputs(3525) <= not((layer3_outputs(8360)) xor (layer3_outputs(5387)));
    layer4_outputs(3526) <= not(layer3_outputs(1224));
    layer4_outputs(3527) <= not(layer3_outputs(518));
    layer4_outputs(3528) <= not(layer3_outputs(5665));
    layer4_outputs(3529) <= layer3_outputs(9683);
    layer4_outputs(3530) <= layer3_outputs(7743);
    layer4_outputs(3531) <= (layer3_outputs(9915)) and (layer3_outputs(195));
    layer4_outputs(3532) <= not(layer3_outputs(5904)) or (layer3_outputs(5642));
    layer4_outputs(3533) <= not(layer3_outputs(7547)) or (layer3_outputs(1770));
    layer4_outputs(3534) <= not((layer3_outputs(7540)) xor (layer3_outputs(8205)));
    layer4_outputs(3535) <= not(layer3_outputs(2126)) or (layer3_outputs(4418));
    layer4_outputs(3536) <= (layer3_outputs(4985)) or (layer3_outputs(8219));
    layer4_outputs(3537) <= (layer3_outputs(9882)) and not (layer3_outputs(6662));
    layer4_outputs(3538) <= (layer3_outputs(7835)) and (layer3_outputs(7062));
    layer4_outputs(3539) <= (layer3_outputs(4319)) and not (layer3_outputs(3831));
    layer4_outputs(3540) <= layer3_outputs(193);
    layer4_outputs(3541) <= (layer3_outputs(1572)) xor (layer3_outputs(1462));
    layer4_outputs(3542) <= (layer3_outputs(7055)) and not (layer3_outputs(1837));
    layer4_outputs(3543) <= layer3_outputs(4802);
    layer4_outputs(3544) <= layer3_outputs(6321);
    layer4_outputs(3545) <= not(layer3_outputs(4400));
    layer4_outputs(3546) <= not(layer3_outputs(9956));
    layer4_outputs(3547) <= (layer3_outputs(1112)) and not (layer3_outputs(1462));
    layer4_outputs(3548) <= (layer3_outputs(7804)) xor (layer3_outputs(6708));
    layer4_outputs(3549) <= not(layer3_outputs(9723));
    layer4_outputs(3550) <= not((layer3_outputs(4006)) or (layer3_outputs(5853)));
    layer4_outputs(3551) <= not(layer3_outputs(2092)) or (layer3_outputs(1317));
    layer4_outputs(3552) <= (layer3_outputs(6424)) and not (layer3_outputs(7548));
    layer4_outputs(3553) <= layer3_outputs(5688);
    layer4_outputs(3554) <= layer3_outputs(9659);
    layer4_outputs(3555) <= not(layer3_outputs(9574));
    layer4_outputs(3556) <= not(layer3_outputs(235));
    layer4_outputs(3557) <= layer3_outputs(6676);
    layer4_outputs(3558) <= not(layer3_outputs(6572));
    layer4_outputs(3559) <= not(layer3_outputs(3516));
    layer4_outputs(3560) <= not(layer3_outputs(10029));
    layer4_outputs(3561) <= layer3_outputs(1737);
    layer4_outputs(3562) <= (layer3_outputs(9727)) and not (layer3_outputs(9773));
    layer4_outputs(3563) <= layer3_outputs(2152);
    layer4_outputs(3564) <= (layer3_outputs(5745)) and (layer3_outputs(8843));
    layer4_outputs(3565) <= layer3_outputs(6130);
    layer4_outputs(3566) <= layer3_outputs(1695);
    layer4_outputs(3567) <= (layer3_outputs(9230)) and not (layer3_outputs(5652));
    layer4_outputs(3568) <= (layer3_outputs(383)) or (layer3_outputs(8001));
    layer4_outputs(3569) <= not((layer3_outputs(1717)) xor (layer3_outputs(3119)));
    layer4_outputs(3570) <= not((layer3_outputs(609)) or (layer3_outputs(566)));
    layer4_outputs(3571) <= (layer3_outputs(8645)) or (layer3_outputs(9323));
    layer4_outputs(3572) <= layer3_outputs(2758);
    layer4_outputs(3573) <= not(layer3_outputs(10051)) or (layer3_outputs(10173));
    layer4_outputs(3574) <= not(layer3_outputs(6178));
    layer4_outputs(3575) <= not((layer3_outputs(7292)) xor (layer3_outputs(3869)));
    layer4_outputs(3576) <= (layer3_outputs(703)) and not (layer3_outputs(1580));
    layer4_outputs(3577) <= layer3_outputs(4832);
    layer4_outputs(3578) <= layer3_outputs(5664);
    layer4_outputs(3579) <= layer3_outputs(7826);
    layer4_outputs(3580) <= not(layer3_outputs(7844));
    layer4_outputs(3581) <= (layer3_outputs(9356)) and not (layer3_outputs(2582));
    layer4_outputs(3582) <= not(layer3_outputs(2569));
    layer4_outputs(3583) <= (layer3_outputs(6314)) xor (layer3_outputs(9773));
    layer4_outputs(3584) <= (layer3_outputs(6246)) and not (layer3_outputs(5695));
    layer4_outputs(3585) <= not((layer3_outputs(9450)) xor (layer3_outputs(6956)));
    layer4_outputs(3586) <= layer3_outputs(5826);
    layer4_outputs(3587) <= not(layer3_outputs(5340));
    layer4_outputs(3588) <= layer3_outputs(6078);
    layer4_outputs(3589) <= not(layer3_outputs(310)) or (layer3_outputs(9901));
    layer4_outputs(3590) <= not(layer3_outputs(8620));
    layer4_outputs(3591) <= layer3_outputs(2952);
    layer4_outputs(3592) <= not(layer3_outputs(151));
    layer4_outputs(3593) <= not((layer3_outputs(10050)) or (layer3_outputs(2498)));
    layer4_outputs(3594) <= (layer3_outputs(3252)) xor (layer3_outputs(7092));
    layer4_outputs(3595) <= (layer3_outputs(1314)) and not (layer3_outputs(3290));
    layer4_outputs(3596) <= not((layer3_outputs(2083)) or (layer3_outputs(9184)));
    layer4_outputs(3597) <= (layer3_outputs(1354)) and not (layer3_outputs(6027));
    layer4_outputs(3598) <= layer3_outputs(3885);
    layer4_outputs(3599) <= not(layer3_outputs(4850)) or (layer3_outputs(7233));
    layer4_outputs(3600) <= not((layer3_outputs(3272)) xor (layer3_outputs(4849)));
    layer4_outputs(3601) <= not(layer3_outputs(3868));
    layer4_outputs(3602) <= not(layer3_outputs(9955));
    layer4_outputs(3603) <= layer3_outputs(7685);
    layer4_outputs(3604) <= not(layer3_outputs(6803));
    layer4_outputs(3605) <= (layer3_outputs(8891)) xor (layer3_outputs(7743));
    layer4_outputs(3606) <= not(layer3_outputs(2252));
    layer4_outputs(3607) <= not((layer3_outputs(7515)) xor (layer3_outputs(2432)));
    layer4_outputs(3608) <= not((layer3_outputs(8097)) xor (layer3_outputs(820)));
    layer4_outputs(3609) <= layer3_outputs(3189);
    layer4_outputs(3610) <= layer3_outputs(4730);
    layer4_outputs(3611) <= (layer3_outputs(1250)) and (layer3_outputs(1143));
    layer4_outputs(3612) <= not(layer3_outputs(2068));
    layer4_outputs(3613) <= not(layer3_outputs(120)) or (layer3_outputs(1484));
    layer4_outputs(3614) <= not(layer3_outputs(976));
    layer4_outputs(3615) <= (layer3_outputs(8813)) and (layer3_outputs(5564));
    layer4_outputs(3616) <= (layer3_outputs(9033)) xor (layer3_outputs(7508));
    layer4_outputs(3617) <= '1';
    layer4_outputs(3618) <= (layer3_outputs(8806)) and not (layer3_outputs(3879));
    layer4_outputs(3619) <= (layer3_outputs(1490)) and (layer3_outputs(8554));
    layer4_outputs(3620) <= not(layer3_outputs(6107));
    layer4_outputs(3621) <= not(layer3_outputs(5698));
    layer4_outputs(3622) <= layer3_outputs(8375);
    layer4_outputs(3623) <= not((layer3_outputs(1785)) and (layer3_outputs(2473)));
    layer4_outputs(3624) <= layer3_outputs(8430);
    layer4_outputs(3625) <= not(layer3_outputs(9350)) or (layer3_outputs(2067));
    layer4_outputs(3626) <= not((layer3_outputs(2363)) xor (layer3_outputs(7949)));
    layer4_outputs(3627) <= not(layer3_outputs(6900)) or (layer3_outputs(6396));
    layer4_outputs(3628) <= (layer3_outputs(2920)) and not (layer3_outputs(1981));
    layer4_outputs(3629) <= not((layer3_outputs(6038)) xor (layer3_outputs(864)));
    layer4_outputs(3630) <= not(layer3_outputs(1777));
    layer4_outputs(3631) <= layer3_outputs(6168);
    layer4_outputs(3632) <= not((layer3_outputs(2168)) or (layer3_outputs(2670)));
    layer4_outputs(3633) <= layer3_outputs(2190);
    layer4_outputs(3634) <= not((layer3_outputs(9477)) and (layer3_outputs(1673)));
    layer4_outputs(3635) <= layer3_outputs(4517);
    layer4_outputs(3636) <= (layer3_outputs(1202)) xor (layer3_outputs(3851));
    layer4_outputs(3637) <= (layer3_outputs(3443)) or (layer3_outputs(416));
    layer4_outputs(3638) <= not((layer3_outputs(2101)) xor (layer3_outputs(6984)));
    layer4_outputs(3639) <= not((layer3_outputs(9552)) xor (layer3_outputs(2529)));
    layer4_outputs(3640) <= layer3_outputs(7682);
    layer4_outputs(3641) <= not(layer3_outputs(10205));
    layer4_outputs(3642) <= layer3_outputs(9464);
    layer4_outputs(3643) <= not(layer3_outputs(3707)) or (layer3_outputs(6474));
    layer4_outputs(3644) <= (layer3_outputs(9067)) and not (layer3_outputs(4797));
    layer4_outputs(3645) <= not((layer3_outputs(1622)) xor (layer3_outputs(5337)));
    layer4_outputs(3646) <= (layer3_outputs(6154)) xor (layer3_outputs(4073));
    layer4_outputs(3647) <= not(layer3_outputs(7017)) or (layer3_outputs(1710));
    layer4_outputs(3648) <= layer3_outputs(1659);
    layer4_outputs(3649) <= layer3_outputs(7970);
    layer4_outputs(3650) <= layer3_outputs(4636);
    layer4_outputs(3651) <= not(layer3_outputs(4586));
    layer4_outputs(3652) <= (layer3_outputs(6126)) xor (layer3_outputs(2496));
    layer4_outputs(3653) <= not(layer3_outputs(5139)) or (layer3_outputs(7169));
    layer4_outputs(3654) <= layer3_outputs(10087);
    layer4_outputs(3655) <= not(layer3_outputs(2154));
    layer4_outputs(3656) <= (layer3_outputs(5309)) xor (layer3_outputs(10184));
    layer4_outputs(3657) <= layer3_outputs(5714);
    layer4_outputs(3658) <= layer3_outputs(439);
    layer4_outputs(3659) <= layer3_outputs(1251);
    layer4_outputs(3660) <= not((layer3_outputs(1696)) xor (layer3_outputs(3066)));
    layer4_outputs(3661) <= not(layer3_outputs(2808));
    layer4_outputs(3662) <= (layer3_outputs(4398)) and not (layer3_outputs(1291));
    layer4_outputs(3663) <= not(layer3_outputs(3350)) or (layer3_outputs(7362));
    layer4_outputs(3664) <= layer3_outputs(2325);
    layer4_outputs(3665) <= not(layer3_outputs(6662));
    layer4_outputs(3666) <= not((layer3_outputs(2274)) and (layer3_outputs(137)));
    layer4_outputs(3667) <= (layer3_outputs(2517)) and not (layer3_outputs(6817));
    layer4_outputs(3668) <= (layer3_outputs(9959)) and not (layer3_outputs(4153));
    layer4_outputs(3669) <= not(layer3_outputs(5776));
    layer4_outputs(3670) <= (layer3_outputs(6012)) and not (layer3_outputs(3775));
    layer4_outputs(3671) <= not(layer3_outputs(7566));
    layer4_outputs(3672) <= not(layer3_outputs(2996));
    layer4_outputs(3673) <= not(layer3_outputs(8884));
    layer4_outputs(3674) <= not(layer3_outputs(4796));
    layer4_outputs(3675) <= (layer3_outputs(6050)) xor (layer3_outputs(5338));
    layer4_outputs(3676) <= layer3_outputs(6778);
    layer4_outputs(3677) <= not(layer3_outputs(907));
    layer4_outputs(3678) <= not((layer3_outputs(6101)) and (layer3_outputs(10134)));
    layer4_outputs(3679) <= layer3_outputs(2079);
    layer4_outputs(3680) <= (layer3_outputs(6707)) and not (layer3_outputs(5585));
    layer4_outputs(3681) <= not((layer3_outputs(3250)) xor (layer3_outputs(1547)));
    layer4_outputs(3682) <= not(layer3_outputs(5005));
    layer4_outputs(3683) <= not((layer3_outputs(2153)) xor (layer3_outputs(189)));
    layer4_outputs(3684) <= layer3_outputs(8689);
    layer4_outputs(3685) <= not((layer3_outputs(6191)) xor (layer3_outputs(7966)));
    layer4_outputs(3686) <= (layer3_outputs(2921)) and not (layer3_outputs(5347));
    layer4_outputs(3687) <= (layer3_outputs(1653)) and not (layer3_outputs(7282));
    layer4_outputs(3688) <= (layer3_outputs(4652)) xor (layer3_outputs(2105));
    layer4_outputs(3689) <= layer3_outputs(2244);
    layer4_outputs(3690) <= not((layer3_outputs(206)) xor (layer3_outputs(9188)));
    layer4_outputs(3691) <= (layer3_outputs(6645)) and not (layer3_outputs(2709));
    layer4_outputs(3692) <= not((layer3_outputs(130)) xor (layer3_outputs(7582)));
    layer4_outputs(3693) <= not(layer3_outputs(9613)) or (layer3_outputs(9215));
    layer4_outputs(3694) <= (layer3_outputs(7000)) and not (layer3_outputs(2098));
    layer4_outputs(3695) <= not((layer3_outputs(7133)) xor (layer3_outputs(279)));
    layer4_outputs(3696) <= layer3_outputs(9787);
    layer4_outputs(3697) <= (layer3_outputs(8699)) xor (layer3_outputs(6907));
    layer4_outputs(3698) <= not((layer3_outputs(6687)) or (layer3_outputs(9224)));
    layer4_outputs(3699) <= layer3_outputs(3095);
    layer4_outputs(3700) <= not(layer3_outputs(1848));
    layer4_outputs(3701) <= not(layer3_outputs(706)) or (layer3_outputs(3227));
    layer4_outputs(3702) <= not(layer3_outputs(1420));
    layer4_outputs(3703) <= not(layer3_outputs(6431));
    layer4_outputs(3704) <= not(layer3_outputs(2014));
    layer4_outputs(3705) <= not(layer3_outputs(9233));
    layer4_outputs(3706) <= not((layer3_outputs(5418)) xor (layer3_outputs(5027)));
    layer4_outputs(3707) <= (layer3_outputs(4202)) and not (layer3_outputs(10215));
    layer4_outputs(3708) <= not(layer3_outputs(5783)) or (layer3_outputs(3477));
    layer4_outputs(3709) <= not((layer3_outputs(5968)) and (layer3_outputs(1357)));
    layer4_outputs(3710) <= not(layer3_outputs(625));
    layer4_outputs(3711) <= '1';
    layer4_outputs(3712) <= (layer3_outputs(3514)) and not (layer3_outputs(5530));
    layer4_outputs(3713) <= (layer3_outputs(1438)) and not (layer3_outputs(8417));
    layer4_outputs(3714) <= '0';
    layer4_outputs(3715) <= not(layer3_outputs(10112));
    layer4_outputs(3716) <= layer3_outputs(1621);
    layer4_outputs(3717) <= not(layer3_outputs(1858));
    layer4_outputs(3718) <= not(layer3_outputs(9742)) or (layer3_outputs(9256));
    layer4_outputs(3719) <= layer3_outputs(1436);
    layer4_outputs(3720) <= (layer3_outputs(6503)) xor (layer3_outputs(8820));
    layer4_outputs(3721) <= (layer3_outputs(1937)) and not (layer3_outputs(2465));
    layer4_outputs(3722) <= layer3_outputs(2319);
    layer4_outputs(3723) <= (layer3_outputs(3481)) and not (layer3_outputs(7670));
    layer4_outputs(3724) <= not(layer3_outputs(9399));
    layer4_outputs(3725) <= layer3_outputs(7468);
    layer4_outputs(3726) <= layer3_outputs(9486);
    layer4_outputs(3727) <= not(layer3_outputs(5471)) or (layer3_outputs(8522));
    layer4_outputs(3728) <= not(layer3_outputs(4784));
    layer4_outputs(3729) <= (layer3_outputs(2437)) and (layer3_outputs(9263));
    layer4_outputs(3730) <= layer3_outputs(7157);
    layer4_outputs(3731) <= not(layer3_outputs(7581));
    layer4_outputs(3732) <= not(layer3_outputs(2804));
    layer4_outputs(3733) <= layer3_outputs(3437);
    layer4_outputs(3734) <= '0';
    layer4_outputs(3735) <= not(layer3_outputs(6076));
    layer4_outputs(3736) <= not((layer3_outputs(266)) xor (layer3_outputs(6534)));
    layer4_outputs(3737) <= not((layer3_outputs(4653)) or (layer3_outputs(5710)));
    layer4_outputs(3738) <= layer3_outputs(8028);
    layer4_outputs(3739) <= layer3_outputs(6959);
    layer4_outputs(3740) <= layer3_outputs(5386);
    layer4_outputs(3741) <= (layer3_outputs(8269)) xor (layer3_outputs(7869));
    layer4_outputs(3742) <= not(layer3_outputs(3610));
    layer4_outputs(3743) <= layer3_outputs(1245);
    layer4_outputs(3744) <= not(layer3_outputs(8369));
    layer4_outputs(3745) <= layer3_outputs(988);
    layer4_outputs(3746) <= not(layer3_outputs(9983));
    layer4_outputs(3747) <= layer3_outputs(8711);
    layer4_outputs(3748) <= not((layer3_outputs(685)) or (layer3_outputs(6614)));
    layer4_outputs(3749) <= not((layer3_outputs(9776)) and (layer3_outputs(9686)));
    layer4_outputs(3750) <= (layer3_outputs(5045)) and not (layer3_outputs(5399));
    layer4_outputs(3751) <= layer3_outputs(1792);
    layer4_outputs(3752) <= not((layer3_outputs(584)) xor (layer3_outputs(5217)));
    layer4_outputs(3753) <= (layer3_outputs(5667)) or (layer3_outputs(3202));
    layer4_outputs(3754) <= (layer3_outputs(6475)) and not (layer3_outputs(2746));
    layer4_outputs(3755) <= (layer3_outputs(5532)) xor (layer3_outputs(10096));
    layer4_outputs(3756) <= not(layer3_outputs(7248));
    layer4_outputs(3757) <= not((layer3_outputs(6889)) and (layer3_outputs(3875)));
    layer4_outputs(3758) <= (layer3_outputs(1407)) and not (layer3_outputs(5087));
    layer4_outputs(3759) <= layer3_outputs(6315);
    layer4_outputs(3760) <= not(layer3_outputs(851));
    layer4_outputs(3761) <= (layer3_outputs(8768)) and (layer3_outputs(7741));
    layer4_outputs(3762) <= layer3_outputs(326);
    layer4_outputs(3763) <= not(layer3_outputs(902));
    layer4_outputs(3764) <= (layer3_outputs(6176)) and (layer3_outputs(3801));
    layer4_outputs(3765) <= (layer3_outputs(275)) xor (layer3_outputs(1624));
    layer4_outputs(3766) <= not(layer3_outputs(7726));
    layer4_outputs(3767) <= not(layer3_outputs(6102)) or (layer3_outputs(1849));
    layer4_outputs(3768) <= not(layer3_outputs(3733));
    layer4_outputs(3769) <= not((layer3_outputs(2073)) xor (layer3_outputs(7701)));
    layer4_outputs(3770) <= layer3_outputs(617);
    layer4_outputs(3771) <= not(layer3_outputs(1105));
    layer4_outputs(3772) <= '1';
    layer4_outputs(3773) <= not(layer3_outputs(6754)) or (layer3_outputs(3523));
    layer4_outputs(3774) <= not(layer3_outputs(8077));
    layer4_outputs(3775) <= not(layer3_outputs(5940));
    layer4_outputs(3776) <= layer3_outputs(5857);
    layer4_outputs(3777) <= not(layer3_outputs(53));
    layer4_outputs(3778) <= not(layer3_outputs(7863));
    layer4_outputs(3779) <= (layer3_outputs(1819)) and not (layer3_outputs(1361));
    layer4_outputs(3780) <= (layer3_outputs(2532)) and (layer3_outputs(5529));
    layer4_outputs(3781) <= (layer3_outputs(5097)) xor (layer3_outputs(1359));
    layer4_outputs(3782) <= (layer3_outputs(9605)) and not (layer3_outputs(6673));
    layer4_outputs(3783) <= not((layer3_outputs(2864)) or (layer3_outputs(1514)));
    layer4_outputs(3784) <= not(layer3_outputs(8492));
    layer4_outputs(3785) <= not((layer3_outputs(5777)) xor (layer3_outputs(4223)));
    layer4_outputs(3786) <= not((layer3_outputs(5729)) or (layer3_outputs(1246)));
    layer4_outputs(3787) <= layer3_outputs(3678);
    layer4_outputs(3788) <= not(layer3_outputs(4363));
    layer4_outputs(3789) <= not(layer3_outputs(5319));
    layer4_outputs(3790) <= not(layer3_outputs(4863)) or (layer3_outputs(9255));
    layer4_outputs(3791) <= not((layer3_outputs(3372)) xor (layer3_outputs(8265)));
    layer4_outputs(3792) <= not(layer3_outputs(4782)) or (layer3_outputs(9655));
    layer4_outputs(3793) <= not(layer3_outputs(8595));
    layer4_outputs(3794) <= layer3_outputs(2777);
    layer4_outputs(3795) <= not(layer3_outputs(6378));
    layer4_outputs(3796) <= not((layer3_outputs(9298)) xor (layer3_outputs(1710)));
    layer4_outputs(3797) <= not(layer3_outputs(7846)) or (layer3_outputs(3064));
    layer4_outputs(3798) <= layer3_outputs(8904);
    layer4_outputs(3799) <= layer3_outputs(2097);
    layer4_outputs(3800) <= not(layer3_outputs(7124));
    layer4_outputs(3801) <= not((layer3_outputs(2274)) and (layer3_outputs(7850)));
    layer4_outputs(3802) <= layer3_outputs(863);
    layer4_outputs(3803) <= (layer3_outputs(1365)) and not (layer3_outputs(1082));
    layer4_outputs(3804) <= layer3_outputs(377);
    layer4_outputs(3805) <= layer3_outputs(3523);
    layer4_outputs(3806) <= (layer3_outputs(4562)) xor (layer3_outputs(5375));
    layer4_outputs(3807) <= layer3_outputs(4270);
    layer4_outputs(3808) <= not((layer3_outputs(6414)) and (layer3_outputs(4156)));
    layer4_outputs(3809) <= layer3_outputs(1674);
    layer4_outputs(3810) <= (layer3_outputs(344)) and not (layer3_outputs(1525));
    layer4_outputs(3811) <= not(layer3_outputs(4364));
    layer4_outputs(3812) <= (layer3_outputs(1459)) xor (layer3_outputs(7241));
    layer4_outputs(3813) <= not((layer3_outputs(7430)) xor (layer3_outputs(6017)));
    layer4_outputs(3814) <= layer3_outputs(2);
    layer4_outputs(3815) <= not(layer3_outputs(9804));
    layer4_outputs(3816) <= not((layer3_outputs(2163)) or (layer3_outputs(397)));
    layer4_outputs(3817) <= layer3_outputs(7102);
    layer4_outputs(3818) <= (layer3_outputs(8170)) xor (layer3_outputs(945));
    layer4_outputs(3819) <= not(layer3_outputs(7984));
    layer4_outputs(3820) <= not(layer3_outputs(1859));
    layer4_outputs(3821) <= layer3_outputs(398);
    layer4_outputs(3822) <= not(layer3_outputs(6509));
    layer4_outputs(3823) <= layer3_outputs(3168);
    layer4_outputs(3824) <= not(layer3_outputs(3114)) or (layer3_outputs(3059));
    layer4_outputs(3825) <= layer3_outputs(8726);
    layer4_outputs(3826) <= layer3_outputs(6899);
    layer4_outputs(3827) <= not(layer3_outputs(8669));
    layer4_outputs(3828) <= not(layer3_outputs(9516));
    layer4_outputs(3829) <= not((layer3_outputs(4254)) xor (layer3_outputs(1284)));
    layer4_outputs(3830) <= not(layer3_outputs(8972));
    layer4_outputs(3831) <= not(layer3_outputs(6433));
    layer4_outputs(3832) <= not(layer3_outputs(260));
    layer4_outputs(3833) <= (layer3_outputs(10121)) and not (layer3_outputs(9459));
    layer4_outputs(3834) <= not((layer3_outputs(265)) xor (layer3_outputs(8268)));
    layer4_outputs(3835) <= layer3_outputs(6674);
    layer4_outputs(3836) <= layer3_outputs(3500);
    layer4_outputs(3837) <= layer3_outputs(8584);
    layer4_outputs(3838) <= (layer3_outputs(490)) or (layer3_outputs(1094));
    layer4_outputs(3839) <= not(layer3_outputs(9154)) or (layer3_outputs(8120));
    layer4_outputs(3840) <= not(layer3_outputs(8621));
    layer4_outputs(3841) <= (layer3_outputs(3629)) or (layer3_outputs(8519));
    layer4_outputs(3842) <= not(layer3_outputs(6797)) or (layer3_outputs(1452));
    layer4_outputs(3843) <= not(layer3_outputs(4143));
    layer4_outputs(3844) <= not((layer3_outputs(4973)) or (layer3_outputs(2196)));
    layer4_outputs(3845) <= not(layer3_outputs(9059));
    layer4_outputs(3846) <= not((layer3_outputs(3782)) xor (layer3_outputs(2831)));
    layer4_outputs(3847) <= (layer3_outputs(10056)) and (layer3_outputs(8405));
    layer4_outputs(3848) <= (layer3_outputs(9881)) and not (layer3_outputs(930));
    layer4_outputs(3849) <= not(layer3_outputs(6947)) or (layer3_outputs(3792));
    layer4_outputs(3850) <= layer3_outputs(8939);
    layer4_outputs(3851) <= not((layer3_outputs(3188)) and (layer3_outputs(2121)));
    layer4_outputs(3852) <= not(layer3_outputs(8986));
    layer4_outputs(3853) <= layer3_outputs(2353);
    layer4_outputs(3854) <= not(layer3_outputs(10093));
    layer4_outputs(3855) <= layer3_outputs(3775);
    layer4_outputs(3856) <= not((layer3_outputs(6507)) or (layer3_outputs(8982)));
    layer4_outputs(3857) <= not((layer3_outputs(4889)) and (layer3_outputs(2504)));
    layer4_outputs(3858) <= not(layer3_outputs(9656));
    layer4_outputs(3859) <= layer3_outputs(9647);
    layer4_outputs(3860) <= layer3_outputs(1110);
    layer4_outputs(3861) <= not(layer3_outputs(8619)) or (layer3_outputs(3166));
    layer4_outputs(3862) <= not(layer3_outputs(2540)) or (layer3_outputs(7340));
    layer4_outputs(3863) <= not((layer3_outputs(5019)) xor (layer3_outputs(9954)));
    layer4_outputs(3864) <= not((layer3_outputs(2179)) xor (layer3_outputs(9571)));
    layer4_outputs(3865) <= layer3_outputs(8992);
    layer4_outputs(3866) <= layer3_outputs(6117);
    layer4_outputs(3867) <= not(layer3_outputs(1396)) or (layer3_outputs(5516));
    layer4_outputs(3868) <= layer3_outputs(4145);
    layer4_outputs(3869) <= layer3_outputs(3433);
    layer4_outputs(3870) <= layer3_outputs(8550);
    layer4_outputs(3871) <= layer3_outputs(2107);
    layer4_outputs(3872) <= layer3_outputs(9588);
    layer4_outputs(3873) <= layer3_outputs(3814);
    layer4_outputs(3874) <= (layer3_outputs(10166)) and not (layer3_outputs(9661));
    layer4_outputs(3875) <= layer3_outputs(6653);
    layer4_outputs(3876) <= (layer3_outputs(355)) and not (layer3_outputs(368));
    layer4_outputs(3877) <= (layer3_outputs(3748)) or (layer3_outputs(4119));
    layer4_outputs(3878) <= layer3_outputs(1788);
    layer4_outputs(3879) <= (layer3_outputs(8126)) and not (layer3_outputs(8275));
    layer4_outputs(3880) <= not(layer3_outputs(9571));
    layer4_outputs(3881) <= layer3_outputs(6917);
    layer4_outputs(3882) <= (layer3_outputs(8274)) and not (layer3_outputs(854));
    layer4_outputs(3883) <= layer3_outputs(6179);
    layer4_outputs(3884) <= not((layer3_outputs(9796)) xor (layer3_outputs(2841)));
    layer4_outputs(3885) <= not(layer3_outputs(607));
    layer4_outputs(3886) <= not((layer3_outputs(3171)) or (layer3_outputs(42)));
    layer4_outputs(3887) <= not(layer3_outputs(4099));
    layer4_outputs(3888) <= not(layer3_outputs(3470));
    layer4_outputs(3889) <= not(layer3_outputs(1744));
    layer4_outputs(3890) <= not((layer3_outputs(3258)) or (layer3_outputs(605)));
    layer4_outputs(3891) <= not(layer3_outputs(4046));
    layer4_outputs(3892) <= not(layer3_outputs(7261));
    layer4_outputs(3893) <= not((layer3_outputs(7226)) xor (layer3_outputs(5237)));
    layer4_outputs(3894) <= (layer3_outputs(9681)) xor (layer3_outputs(8607));
    layer4_outputs(3895) <= (layer3_outputs(9675)) and (layer3_outputs(6376));
    layer4_outputs(3896) <= not(layer3_outputs(10138));
    layer4_outputs(3897) <= not((layer3_outputs(3485)) and (layer3_outputs(9172)));
    layer4_outputs(3898) <= layer3_outputs(7808);
    layer4_outputs(3899) <= (layer3_outputs(5661)) and not (layer3_outputs(1116));
    layer4_outputs(3900) <= not(layer3_outputs(674));
    layer4_outputs(3901) <= (layer3_outputs(10078)) and (layer3_outputs(7821));
    layer4_outputs(3902) <= not(layer3_outputs(3098));
    layer4_outputs(3903) <= (layer3_outputs(6656)) and not (layer3_outputs(9389));
    layer4_outputs(3904) <= (layer3_outputs(541)) and (layer3_outputs(3968));
    layer4_outputs(3905) <= (layer3_outputs(7069)) and (layer3_outputs(391));
    layer4_outputs(3906) <= layer3_outputs(6235);
    layer4_outputs(3907) <= (layer3_outputs(7957)) xor (layer3_outputs(2351));
    layer4_outputs(3908) <= layer3_outputs(3327);
    layer4_outputs(3909) <= layer3_outputs(7612);
    layer4_outputs(3910) <= not((layer3_outputs(2448)) or (layer3_outputs(1043)));
    layer4_outputs(3911) <= (layer3_outputs(4309)) and (layer3_outputs(6743));
    layer4_outputs(3912) <= (layer3_outputs(423)) and not (layer3_outputs(5726));
    layer4_outputs(3913) <= not(layer3_outputs(4659));
    layer4_outputs(3914) <= not(layer3_outputs(5847)) or (layer3_outputs(3654));
    layer4_outputs(3915) <= not(layer3_outputs(3175));
    layer4_outputs(3916) <= (layer3_outputs(6893)) and not (layer3_outputs(4299));
    layer4_outputs(3917) <= layer3_outputs(5937);
    layer4_outputs(3918) <= layer3_outputs(5859);
    layer4_outputs(3919) <= not(layer3_outputs(5687));
    layer4_outputs(3920) <= (layer3_outputs(3351)) and (layer3_outputs(3905));
    layer4_outputs(3921) <= layer3_outputs(7275);
    layer4_outputs(3922) <= (layer3_outputs(5130)) xor (layer3_outputs(2426));
    layer4_outputs(3923) <= not((layer3_outputs(855)) xor (layer3_outputs(5977)));
    layer4_outputs(3924) <= not(layer3_outputs(4104));
    layer4_outputs(3925) <= not(layer3_outputs(18));
    layer4_outputs(3926) <= (layer3_outputs(9292)) and not (layer3_outputs(9006));
    layer4_outputs(3927) <= (layer3_outputs(7586)) or (layer3_outputs(7883));
    layer4_outputs(3928) <= (layer3_outputs(3393)) and (layer3_outputs(5887));
    layer4_outputs(3929) <= not((layer3_outputs(8979)) xor (layer3_outputs(4123)));
    layer4_outputs(3930) <= layer3_outputs(3853);
    layer4_outputs(3931) <= (layer3_outputs(4745)) and not (layer3_outputs(4725));
    layer4_outputs(3932) <= not((layer3_outputs(3451)) or (layer3_outputs(6548)));
    layer4_outputs(3933) <= not(layer3_outputs(5453));
    layer4_outputs(3934) <= layer3_outputs(7200);
    layer4_outputs(3935) <= not(layer3_outputs(7165));
    layer4_outputs(3936) <= not(layer3_outputs(9620));
    layer4_outputs(3937) <= not(layer3_outputs(10160));
    layer4_outputs(3938) <= not((layer3_outputs(1808)) and (layer3_outputs(8687)));
    layer4_outputs(3939) <= not(layer3_outputs(9464));
    layer4_outputs(3940) <= layer3_outputs(7609);
    layer4_outputs(3941) <= (layer3_outputs(3522)) or (layer3_outputs(3925));
    layer4_outputs(3942) <= (layer3_outputs(62)) and (layer3_outputs(2024));
    layer4_outputs(3943) <= not(layer3_outputs(16)) or (layer3_outputs(171));
    layer4_outputs(3944) <= not(layer3_outputs(1811));
    layer4_outputs(3945) <= not(layer3_outputs(2437));
    layer4_outputs(3946) <= layer3_outputs(2460);
    layer4_outputs(3947) <= (layer3_outputs(4897)) xor (layer3_outputs(5078));
    layer4_outputs(3948) <= not(layer3_outputs(9318));
    layer4_outputs(3949) <= not(layer3_outputs(716));
    layer4_outputs(3950) <= '1';
    layer4_outputs(3951) <= '1';
    layer4_outputs(3952) <= layer3_outputs(9582);
    layer4_outputs(3953) <= (layer3_outputs(9719)) or (layer3_outputs(3641));
    layer4_outputs(3954) <= layer3_outputs(1266);
    layer4_outputs(3955) <= (layer3_outputs(3529)) and not (layer3_outputs(4504));
    layer4_outputs(3956) <= (layer3_outputs(1740)) or (layer3_outputs(4509));
    layer4_outputs(3957) <= not(layer3_outputs(10087)) or (layer3_outputs(3395));
    layer4_outputs(3958) <= (layer3_outputs(4769)) and (layer3_outputs(7640));
    layer4_outputs(3959) <= not(layer3_outputs(9740));
    layer4_outputs(3960) <= not(layer3_outputs(68));
    layer4_outputs(3961) <= not(layer3_outputs(3834));
    layer4_outputs(3962) <= not(layer3_outputs(1304));
    layer4_outputs(3963) <= (layer3_outputs(8654)) and not (layer3_outputs(7078));
    layer4_outputs(3964) <= not(layer3_outputs(5446));
    layer4_outputs(3965) <= not((layer3_outputs(4998)) and (layer3_outputs(9076)));
    layer4_outputs(3966) <= (layer3_outputs(9143)) xor (layer3_outputs(10153));
    layer4_outputs(3967) <= layer3_outputs(5972);
    layer4_outputs(3968) <= not((layer3_outputs(3766)) and (layer3_outputs(5624)));
    layer4_outputs(3969) <= layer3_outputs(4036);
    layer4_outputs(3970) <= not(layer3_outputs(1356)) or (layer3_outputs(7437));
    layer4_outputs(3971) <= (layer3_outputs(291)) xor (layer3_outputs(7598));
    layer4_outputs(3972) <= not(layer3_outputs(1881));
    layer4_outputs(3973) <= (layer3_outputs(8842)) and not (layer3_outputs(5036));
    layer4_outputs(3974) <= layer3_outputs(4173);
    layer4_outputs(3975) <= layer3_outputs(2134);
    layer4_outputs(3976) <= not(layer3_outputs(667));
    layer4_outputs(3977) <= (layer3_outputs(6773)) and not (layer3_outputs(6546));
    layer4_outputs(3978) <= layer3_outputs(6755);
    layer4_outputs(3979) <= layer3_outputs(1147);
    layer4_outputs(3980) <= not(layer3_outputs(2191));
    layer4_outputs(3981) <= not(layer3_outputs(5458));
    layer4_outputs(3982) <= (layer3_outputs(8032)) xor (layer3_outputs(8922));
    layer4_outputs(3983) <= not((layer3_outputs(8558)) xor (layer3_outputs(9907)));
    layer4_outputs(3984) <= not(layer3_outputs(8170));
    layer4_outputs(3985) <= layer3_outputs(6714);
    layer4_outputs(3986) <= not(layer3_outputs(3554));
    layer4_outputs(3987) <= not(layer3_outputs(1642)) or (layer3_outputs(9119));
    layer4_outputs(3988) <= (layer3_outputs(4692)) xor (layer3_outputs(7839));
    layer4_outputs(3989) <= not(layer3_outputs(4395));
    layer4_outputs(3990) <= not((layer3_outputs(7830)) or (layer3_outputs(4828)));
    layer4_outputs(3991) <= not(layer3_outputs(3615));
    layer4_outputs(3992) <= not((layer3_outputs(3092)) xor (layer3_outputs(99)));
    layer4_outputs(3993) <= not((layer3_outputs(9689)) or (layer3_outputs(5543)));
    layer4_outputs(3994) <= layer3_outputs(1897);
    layer4_outputs(3995) <= layer3_outputs(2010);
    layer4_outputs(3996) <= not(layer3_outputs(5734));
    layer4_outputs(3997) <= layer3_outputs(966);
    layer4_outputs(3998) <= not((layer3_outputs(9765)) or (layer3_outputs(2415)));
    layer4_outputs(3999) <= (layer3_outputs(7299)) xor (layer3_outputs(572));
    layer4_outputs(4000) <= (layer3_outputs(5427)) or (layer3_outputs(6997));
    layer4_outputs(4001) <= (layer3_outputs(3140)) xor (layer3_outputs(2303));
    layer4_outputs(4002) <= not(layer3_outputs(4089));
    layer4_outputs(4003) <= not((layer3_outputs(5666)) xor (layer3_outputs(7028)));
    layer4_outputs(4004) <= layer3_outputs(2601);
    layer4_outputs(4005) <= not(layer3_outputs(2707));
    layer4_outputs(4006) <= layer3_outputs(1446);
    layer4_outputs(4007) <= not(layer3_outputs(6000));
    layer4_outputs(4008) <= not(layer3_outputs(4276)) or (layer3_outputs(5335));
    layer4_outputs(4009) <= not((layer3_outputs(8156)) or (layer3_outputs(9329)));
    layer4_outputs(4010) <= layer3_outputs(6882);
    layer4_outputs(4011) <= not((layer3_outputs(856)) xor (layer3_outputs(3307)));
    layer4_outputs(4012) <= not((layer3_outputs(922)) or (layer3_outputs(6824)));
    layer4_outputs(4013) <= layer3_outputs(1087);
    layer4_outputs(4014) <= not(layer3_outputs(6408));
    layer4_outputs(4015) <= not(layer3_outputs(8359)) or (layer3_outputs(2292));
    layer4_outputs(4016) <= not(layer3_outputs(6460));
    layer4_outputs(4017) <= layer3_outputs(1458);
    layer4_outputs(4018) <= layer3_outputs(1036);
    layer4_outputs(4019) <= not(layer3_outputs(6175)) or (layer3_outputs(8229));
    layer4_outputs(4020) <= not(layer3_outputs(535));
    layer4_outputs(4021) <= not(layer3_outputs(5239));
    layer4_outputs(4022) <= not((layer3_outputs(2767)) xor (layer3_outputs(2659)));
    layer4_outputs(4023) <= not(layer3_outputs(8327));
    layer4_outputs(4024) <= not(layer3_outputs(1335));
    layer4_outputs(4025) <= not((layer3_outputs(8690)) or (layer3_outputs(6944)));
    layer4_outputs(4026) <= layer3_outputs(1477);
    layer4_outputs(4027) <= not((layer3_outputs(8946)) xor (layer3_outputs(294)));
    layer4_outputs(4028) <= (layer3_outputs(6674)) or (layer3_outputs(2525));
    layer4_outputs(4029) <= not(layer3_outputs(6629)) or (layer3_outputs(6988));
    layer4_outputs(4030) <= layer3_outputs(3746);
    layer4_outputs(4031) <= (layer3_outputs(4166)) and not (layer3_outputs(1493));
    layer4_outputs(4032) <= not((layer3_outputs(5084)) xor (layer3_outputs(10134)));
    layer4_outputs(4033) <= layer3_outputs(5537);
    layer4_outputs(4034) <= not((layer3_outputs(6634)) xor (layer3_outputs(10099)));
    layer4_outputs(4035) <= (layer3_outputs(6872)) and not (layer3_outputs(9055));
    layer4_outputs(4036) <= not((layer3_outputs(709)) and (layer3_outputs(4172)));
    layer4_outputs(4037) <= not((layer3_outputs(6522)) xor (layer3_outputs(4336)));
    layer4_outputs(4038) <= not(layer3_outputs(2438));
    layer4_outputs(4039) <= not(layer3_outputs(2309)) or (layer3_outputs(4472));
    layer4_outputs(4040) <= not(layer3_outputs(9425));
    layer4_outputs(4041) <= layer3_outputs(5319);
    layer4_outputs(4042) <= not((layer3_outputs(4914)) or (layer3_outputs(6901)));
    layer4_outputs(4043) <= (layer3_outputs(3849)) xor (layer3_outputs(937));
    layer4_outputs(4044) <= not(layer3_outputs(2876));
    layer4_outputs(4045) <= layer3_outputs(7433);
    layer4_outputs(4046) <= not(layer3_outputs(222));
    layer4_outputs(4047) <= '0';
    layer4_outputs(4048) <= layer3_outputs(8623);
    layer4_outputs(4049) <= not(layer3_outputs(8834)) or (layer3_outputs(8121));
    layer4_outputs(4050) <= not((layer3_outputs(9586)) or (layer3_outputs(510)));
    layer4_outputs(4051) <= not(layer3_outputs(9673));
    layer4_outputs(4052) <= (layer3_outputs(7520)) or (layer3_outputs(1945));
    layer4_outputs(4053) <= (layer3_outputs(9867)) or (layer3_outputs(923));
    layer4_outputs(4054) <= not((layer3_outputs(8950)) xor (layer3_outputs(1804)));
    layer4_outputs(4055) <= '0';
    layer4_outputs(4056) <= not(layer3_outputs(2076));
    layer4_outputs(4057) <= not((layer3_outputs(3896)) xor (layer3_outputs(8572)));
    layer4_outputs(4058) <= not((layer3_outputs(6406)) and (layer3_outputs(3590)));
    layer4_outputs(4059) <= (layer3_outputs(3873)) xor (layer3_outputs(3445));
    layer4_outputs(4060) <= not((layer3_outputs(1979)) xor (layer3_outputs(5933)));
    layer4_outputs(4061) <= not((layer3_outputs(8978)) xor (layer3_outputs(3198)));
    layer4_outputs(4062) <= not((layer3_outputs(3146)) xor (layer3_outputs(468)));
    layer4_outputs(4063) <= not(layer3_outputs(6924));
    layer4_outputs(4064) <= not(layer3_outputs(4142)) or (layer3_outputs(2816));
    layer4_outputs(4065) <= layer3_outputs(8856);
    layer4_outputs(4066) <= (layer3_outputs(4090)) or (layer3_outputs(7972));
    layer4_outputs(4067) <= '1';
    layer4_outputs(4068) <= layer3_outputs(9639);
    layer4_outputs(4069) <= not((layer3_outputs(3981)) and (layer3_outputs(8176)));
    layer4_outputs(4070) <= layer3_outputs(2961);
    layer4_outputs(4071) <= not(layer3_outputs(5961));
    layer4_outputs(4072) <= layer3_outputs(6843);
    layer4_outputs(4073) <= not((layer3_outputs(898)) xor (layer3_outputs(6009)));
    layer4_outputs(4074) <= not(layer3_outputs(6024));
    layer4_outputs(4075) <= (layer3_outputs(2699)) xor (layer3_outputs(9606));
    layer4_outputs(4076) <= (layer3_outputs(9467)) or (layer3_outputs(3551));
    layer4_outputs(4077) <= (layer3_outputs(2163)) and not (layer3_outputs(5906));
    layer4_outputs(4078) <= (layer3_outputs(6767)) xor (layer3_outputs(6542));
    layer4_outputs(4079) <= layer3_outputs(3829);
    layer4_outputs(4080) <= (layer3_outputs(10067)) xor (layer3_outputs(6638));
    layer4_outputs(4081) <= layer3_outputs(7954);
    layer4_outputs(4082) <= not(layer3_outputs(8786));
    layer4_outputs(4083) <= layer3_outputs(4075);
    layer4_outputs(4084) <= not(layer3_outputs(924));
    layer4_outputs(4085) <= layer3_outputs(3958);
    layer4_outputs(4086) <= layer3_outputs(8246);
    layer4_outputs(4087) <= layer3_outputs(568);
    layer4_outputs(4088) <= not((layer3_outputs(2746)) or (layer3_outputs(1435)));
    layer4_outputs(4089) <= not(layer3_outputs(7954));
    layer4_outputs(4090) <= not(layer3_outputs(8700));
    layer4_outputs(4091) <= not(layer3_outputs(9418)) or (layer3_outputs(7452));
    layer4_outputs(4092) <= not((layer3_outputs(8980)) xor (layer3_outputs(2322)));
    layer4_outputs(4093) <= not(layer3_outputs(6270));
    layer4_outputs(4094) <= not(layer3_outputs(5656));
    layer4_outputs(4095) <= not(layer3_outputs(8010));
    layer4_outputs(4096) <= '0';
    layer4_outputs(4097) <= not(layer3_outputs(8627));
    layer4_outputs(4098) <= not((layer3_outputs(45)) xor (layer3_outputs(8418)));
    layer4_outputs(4099) <= not((layer3_outputs(2214)) and (layer3_outputs(1769)));
    layer4_outputs(4100) <= not(layer3_outputs(2118));
    layer4_outputs(4101) <= (layer3_outputs(3660)) or (layer3_outputs(7309));
    layer4_outputs(4102) <= not(layer3_outputs(4589)) or (layer3_outputs(1099));
    layer4_outputs(4103) <= not(layer3_outputs(4313)) or (layer3_outputs(1274));
    layer4_outputs(4104) <= not(layer3_outputs(7095));
    layer4_outputs(4105) <= not((layer3_outputs(7798)) or (layer3_outputs(7489)));
    layer4_outputs(4106) <= not(layer3_outputs(3571));
    layer4_outputs(4107) <= layer3_outputs(1050);
    layer4_outputs(4108) <= not(layer3_outputs(10055));
    layer4_outputs(4109) <= layer3_outputs(1704);
    layer4_outputs(4110) <= not(layer3_outputs(6430)) or (layer3_outputs(3640));
    layer4_outputs(4111) <= layer3_outputs(6206);
    layer4_outputs(4112) <= (layer3_outputs(9074)) xor (layer3_outputs(9989));
    layer4_outputs(4113) <= not(layer3_outputs(7256));
    layer4_outputs(4114) <= layer3_outputs(664);
    layer4_outputs(4115) <= not(layer3_outputs(4833));
    layer4_outputs(4116) <= not(layer3_outputs(7114));
    layer4_outputs(4117) <= not((layer3_outputs(5470)) xor (layer3_outputs(2372)));
    layer4_outputs(4118) <= not(layer3_outputs(7146));
    layer4_outputs(4119) <= not(layer3_outputs(3020));
    layer4_outputs(4120) <= (layer3_outputs(6178)) and not (layer3_outputs(4155));
    layer4_outputs(4121) <= (layer3_outputs(8709)) and (layer3_outputs(2033));
    layer4_outputs(4122) <= '0';
    layer4_outputs(4123) <= not((layer3_outputs(8009)) xor (layer3_outputs(654)));
    layer4_outputs(4124) <= layer3_outputs(2865);
    layer4_outputs(4125) <= layer3_outputs(4518);
    layer4_outputs(4126) <= layer3_outputs(4275);
    layer4_outputs(4127) <= (layer3_outputs(1708)) and not (layer3_outputs(4195));
    layer4_outputs(4128) <= not(layer3_outputs(9299));
    layer4_outputs(4129) <= not(layer3_outputs(1225));
    layer4_outputs(4130) <= not((layer3_outputs(7437)) xor (layer3_outputs(6801)));
    layer4_outputs(4131) <= not((layer3_outputs(9935)) or (layer3_outputs(9781)));
    layer4_outputs(4132) <= layer3_outputs(8127);
    layer4_outputs(4133) <= not(layer3_outputs(8954)) or (layer3_outputs(4690));
    layer4_outputs(4134) <= layer3_outputs(4926);
    layer4_outputs(4135) <= not(layer3_outputs(4570)) or (layer3_outputs(5793));
    layer4_outputs(4136) <= not(layer3_outputs(1818));
    layer4_outputs(4137) <= not(layer3_outputs(2471));
    layer4_outputs(4138) <= layer3_outputs(1298);
    layer4_outputs(4139) <= not(layer3_outputs(3423));
    layer4_outputs(4140) <= layer3_outputs(4857);
    layer4_outputs(4141) <= not(layer3_outputs(6075));
    layer4_outputs(4142) <= layer3_outputs(5089);
    layer4_outputs(4143) <= (layer3_outputs(6928)) or (layer3_outputs(2564));
    layer4_outputs(4144) <= layer3_outputs(1165);
    layer4_outputs(4145) <= not((layer3_outputs(9841)) or (layer3_outputs(3957)));
    layer4_outputs(4146) <= not(layer3_outputs(9648));
    layer4_outputs(4147) <= layer3_outputs(7478);
    layer4_outputs(4148) <= not(layer3_outputs(8650));
    layer4_outputs(4149) <= (layer3_outputs(6230)) xor (layer3_outputs(7039));
    layer4_outputs(4150) <= layer3_outputs(2563);
    layer4_outputs(4151) <= not(layer3_outputs(9887));
    layer4_outputs(4152) <= not(layer3_outputs(1681)) or (layer3_outputs(5493));
    layer4_outputs(4153) <= not(layer3_outputs(1871)) or (layer3_outputs(8910));
    layer4_outputs(4154) <= not(layer3_outputs(6274)) or (layer3_outputs(1243));
    layer4_outputs(4155) <= not(layer3_outputs(4773));
    layer4_outputs(4156) <= not(layer3_outputs(7858));
    layer4_outputs(4157) <= layer3_outputs(6919);
    layer4_outputs(4158) <= not(layer3_outputs(9442));
    layer4_outputs(4159) <= not(layer3_outputs(3916));
    layer4_outputs(4160) <= layer3_outputs(6797);
    layer4_outputs(4161) <= not(layer3_outputs(578)) or (layer3_outputs(2532));
    layer4_outputs(4162) <= not(layer3_outputs(6326));
    layer4_outputs(4163) <= not(layer3_outputs(5854));
    layer4_outputs(4164) <= (layer3_outputs(5985)) and not (layer3_outputs(6195));
    layer4_outputs(4165) <= not(layer3_outputs(9327)) or (layer3_outputs(8595));
    layer4_outputs(4166) <= layer3_outputs(7973);
    layer4_outputs(4167) <= layer3_outputs(2715);
    layer4_outputs(4168) <= layer3_outputs(2213);
    layer4_outputs(4169) <= not((layer3_outputs(6874)) xor (layer3_outputs(9723)));
    layer4_outputs(4170) <= not(layer3_outputs(1345));
    layer4_outputs(4171) <= layer3_outputs(4963);
    layer4_outputs(4172) <= layer3_outputs(856);
    layer4_outputs(4173) <= layer3_outputs(4910);
    layer4_outputs(4174) <= not(layer3_outputs(6180));
    layer4_outputs(4175) <= layer3_outputs(2002);
    layer4_outputs(4176) <= not((layer3_outputs(7677)) xor (layer3_outputs(5254)));
    layer4_outputs(4177) <= not((layer3_outputs(6688)) and (layer3_outputs(3874)));
    layer4_outputs(4178) <= (layer3_outputs(5876)) xor (layer3_outputs(6041));
    layer4_outputs(4179) <= not((layer3_outputs(9419)) xor (layer3_outputs(5864)));
    layer4_outputs(4180) <= layer3_outputs(3900);
    layer4_outputs(4181) <= not(layer3_outputs(3764));
    layer4_outputs(4182) <= (layer3_outputs(2241)) and (layer3_outputs(9001));
    layer4_outputs(4183) <= (layer3_outputs(8586)) xor (layer3_outputs(6904));
    layer4_outputs(4184) <= not(layer3_outputs(10042));
    layer4_outputs(4185) <= layer3_outputs(8141);
    layer4_outputs(4186) <= (layer3_outputs(8998)) and not (layer3_outputs(1640));
    layer4_outputs(4187) <= not(layer3_outputs(8552));
    layer4_outputs(4188) <= (layer3_outputs(2597)) xor (layer3_outputs(10190));
    layer4_outputs(4189) <= not((layer3_outputs(4576)) xor (layer3_outputs(3030)));
    layer4_outputs(4190) <= '0';
    layer4_outputs(4191) <= not((layer3_outputs(2624)) or (layer3_outputs(2900)));
    layer4_outputs(4192) <= not(layer3_outputs(7689));
    layer4_outputs(4193) <= (layer3_outputs(3401)) and (layer3_outputs(1537));
    layer4_outputs(4194) <= (layer3_outputs(8644)) xor (layer3_outputs(6215));
    layer4_outputs(4195) <= layer3_outputs(5808);
    layer4_outputs(4196) <= '0';
    layer4_outputs(4197) <= not((layer3_outputs(7714)) xor (layer3_outputs(5814)));
    layer4_outputs(4198) <= not((layer3_outputs(3145)) or (layer3_outputs(8484)));
    layer4_outputs(4199) <= not((layer3_outputs(8664)) and (layer3_outputs(5008)));
    layer4_outputs(4200) <= layer3_outputs(7711);
    layer4_outputs(4201) <= (layer3_outputs(6596)) xor (layer3_outputs(4407));
    layer4_outputs(4202) <= not((layer3_outputs(4067)) xor (layer3_outputs(6172)));
    layer4_outputs(4203) <= (layer3_outputs(7454)) xor (layer3_outputs(892));
    layer4_outputs(4204) <= not(layer3_outputs(583)) or (layer3_outputs(6048));
    layer4_outputs(4205) <= not(layer3_outputs(9336));
    layer4_outputs(4206) <= not(layer3_outputs(7630));
    layer4_outputs(4207) <= not(layer3_outputs(5607));
    layer4_outputs(4208) <= not((layer3_outputs(3135)) xor (layer3_outputs(6174)));
    layer4_outputs(4209) <= (layer3_outputs(2047)) xor (layer3_outputs(7128));
    layer4_outputs(4210) <= not(layer3_outputs(3945));
    layer4_outputs(4211) <= not((layer3_outputs(6959)) or (layer3_outputs(2365)));
    layer4_outputs(4212) <= not(layer3_outputs(2881));
    layer4_outputs(4213) <= not((layer3_outputs(6611)) and (layer3_outputs(974)));
    layer4_outputs(4214) <= not(layer3_outputs(1911));
    layer4_outputs(4215) <= not((layer3_outputs(2409)) xor (layer3_outputs(6775)));
    layer4_outputs(4216) <= layer3_outputs(9106);
    layer4_outputs(4217) <= not(layer3_outputs(3284)) or (layer3_outputs(517));
    layer4_outputs(4218) <= not(layer3_outputs(5394));
    layer4_outputs(4219) <= layer3_outputs(7889);
    layer4_outputs(4220) <= not(layer3_outputs(418));
    layer4_outputs(4221) <= not(layer3_outputs(3031));
    layer4_outputs(4222) <= layer3_outputs(6679);
    layer4_outputs(4223) <= not(layer3_outputs(9708));
    layer4_outputs(4224) <= (layer3_outputs(3418)) and (layer3_outputs(2228));
    layer4_outputs(4225) <= (layer3_outputs(3269)) and not (layer3_outputs(8735));
    layer4_outputs(4226) <= layer3_outputs(8667);
    layer4_outputs(4227) <= (layer3_outputs(9418)) and not (layer3_outputs(3322));
    layer4_outputs(4228) <= layer3_outputs(4764);
    layer4_outputs(4229) <= not(layer3_outputs(9880)) or (layer3_outputs(7707));
    layer4_outputs(4230) <= (layer3_outputs(8984)) and not (layer3_outputs(6435));
    layer4_outputs(4231) <= not((layer3_outputs(6233)) or (layer3_outputs(3504)));
    layer4_outputs(4232) <= layer3_outputs(1563);
    layer4_outputs(4233) <= (layer3_outputs(1784)) and (layer3_outputs(844));
    layer4_outputs(4234) <= layer3_outputs(36);
    layer4_outputs(4235) <= (layer3_outputs(5172)) and (layer3_outputs(3210));
    layer4_outputs(4236) <= layer3_outputs(8033);
    layer4_outputs(4237) <= not(layer3_outputs(6471));
    layer4_outputs(4238) <= layer3_outputs(5951);
    layer4_outputs(4239) <= not((layer3_outputs(200)) xor (layer3_outputs(588)));
    layer4_outputs(4240) <= not((layer3_outputs(7341)) and (layer3_outputs(2473)));
    layer4_outputs(4241) <= not((layer3_outputs(1916)) xor (layer3_outputs(2115)));
    layer4_outputs(4242) <= layer3_outputs(544);
    layer4_outputs(4243) <= (layer3_outputs(1046)) and not (layer3_outputs(8012));
    layer4_outputs(4244) <= not((layer3_outputs(2823)) xor (layer3_outputs(9398)));
    layer4_outputs(4245) <= layer3_outputs(6816);
    layer4_outputs(4246) <= layer3_outputs(10185);
    layer4_outputs(4247) <= not(layer3_outputs(3960));
    layer4_outputs(4248) <= not(layer3_outputs(9658));
    layer4_outputs(4249) <= not((layer3_outputs(1228)) xor (layer3_outputs(2671)));
    layer4_outputs(4250) <= layer3_outputs(7493);
    layer4_outputs(4251) <= layer3_outputs(3544);
    layer4_outputs(4252) <= not(layer3_outputs(2055));
    layer4_outputs(4253) <= (layer3_outputs(5683)) and not (layer3_outputs(1113));
    layer4_outputs(4254) <= (layer3_outputs(6459)) and (layer3_outputs(4507));
    layer4_outputs(4255) <= layer3_outputs(3548);
    layer4_outputs(4256) <= '0';
    layer4_outputs(4257) <= not(layer3_outputs(8283));
    layer4_outputs(4258) <= not(layer3_outputs(8230)) or (layer3_outputs(6229));
    layer4_outputs(4259) <= not((layer3_outputs(1992)) xor (layer3_outputs(8076)));
    layer4_outputs(4260) <= not(layer3_outputs(5685));
    layer4_outputs(4261) <= (layer3_outputs(5534)) xor (layer3_outputs(3817));
    layer4_outputs(4262) <= layer3_outputs(6204);
    layer4_outputs(4263) <= not(layer3_outputs(6205));
    layer4_outputs(4264) <= not(layer3_outputs(3136));
    layer4_outputs(4265) <= layer3_outputs(5046);
    layer4_outputs(4266) <= layer3_outputs(6308);
    layer4_outputs(4267) <= not(layer3_outputs(7323));
    layer4_outputs(4268) <= (layer3_outputs(5066)) and not (layer3_outputs(8670));
    layer4_outputs(4269) <= not(layer3_outputs(9484));
    layer4_outputs(4270) <= not(layer3_outputs(6750));
    layer4_outputs(4271) <= not(layer3_outputs(428)) or (layer3_outputs(4732));
    layer4_outputs(4272) <= (layer3_outputs(3374)) xor (layer3_outputs(10234));
    layer4_outputs(4273) <= not(layer3_outputs(1224)) or (layer3_outputs(6586));
    layer4_outputs(4274) <= not(layer3_outputs(7672));
    layer4_outputs(4275) <= (layer3_outputs(550)) or (layer3_outputs(9397));
    layer4_outputs(4276) <= layer3_outputs(2628);
    layer4_outputs(4277) <= '0';
    layer4_outputs(4278) <= (layer3_outputs(7394)) xor (layer3_outputs(1147));
    layer4_outputs(4279) <= not((layer3_outputs(7187)) xor (layer3_outputs(6716)));
    layer4_outputs(4280) <= layer3_outputs(4003);
    layer4_outputs(4281) <= layer3_outputs(4196);
    layer4_outputs(4282) <= (layer3_outputs(4018)) xor (layer3_outputs(3854));
    layer4_outputs(4283) <= not((layer3_outputs(3172)) or (layer3_outputs(6517)));
    layer4_outputs(4284) <= not(layer3_outputs(841));
    layer4_outputs(4285) <= (layer3_outputs(4399)) xor (layer3_outputs(1410));
    layer4_outputs(4286) <= (layer3_outputs(8602)) and not (layer3_outputs(2640));
    layer4_outputs(4287) <= not((layer3_outputs(3283)) or (layer3_outputs(7148)));
    layer4_outputs(4288) <= layer3_outputs(8865);
    layer4_outputs(4289) <= layer3_outputs(3182);
    layer4_outputs(4290) <= not(layer3_outputs(8928));
    layer4_outputs(4291) <= not(layer3_outputs(1781)) or (layer3_outputs(8259));
    layer4_outputs(4292) <= not(layer3_outputs(8881));
    layer4_outputs(4293) <= layer3_outputs(4683);
    layer4_outputs(4294) <= not(layer3_outputs(2708));
    layer4_outputs(4295) <= (layer3_outputs(9549)) and not (layer3_outputs(6635));
    layer4_outputs(4296) <= not((layer3_outputs(8869)) xor (layer3_outputs(2363)));
    layer4_outputs(4297) <= not(layer3_outputs(2448));
    layer4_outputs(4298) <= not((layer3_outputs(2723)) xor (layer3_outputs(9768)));
    layer4_outputs(4299) <= layer3_outputs(2889);
    layer4_outputs(4300) <= not((layer3_outputs(7744)) xor (layer3_outputs(3918)));
    layer4_outputs(4301) <= (layer3_outputs(8335)) and (layer3_outputs(3680));
    layer4_outputs(4302) <= not(layer3_outputs(9992));
    layer4_outputs(4303) <= (layer3_outputs(10175)) xor (layer3_outputs(8670));
    layer4_outputs(4304) <= not(layer3_outputs(5285));
    layer4_outputs(4305) <= not(layer3_outputs(4024));
    layer4_outputs(4306) <= not((layer3_outputs(8101)) xor (layer3_outputs(4907)));
    layer4_outputs(4307) <= not((layer3_outputs(8053)) or (layer3_outputs(665)));
    layer4_outputs(4308) <= not(layer3_outputs(9847));
    layer4_outputs(4309) <= not(layer3_outputs(2329));
    layer4_outputs(4310) <= layer3_outputs(6777);
    layer4_outputs(4311) <= layer3_outputs(6219);
    layer4_outputs(4312) <= not((layer3_outputs(6271)) xor (layer3_outputs(2672)));
    layer4_outputs(4313) <= not(layer3_outputs(8870));
    layer4_outputs(4314) <= '1';
    layer4_outputs(4315) <= layer3_outputs(10028);
    layer4_outputs(4316) <= (layer3_outputs(7845)) and not (layer3_outputs(3085));
    layer4_outputs(4317) <= not((layer3_outputs(10151)) xor (layer3_outputs(591)));
    layer4_outputs(4318) <= not(layer3_outputs(8743));
    layer4_outputs(4319) <= layer3_outputs(9352);
    layer4_outputs(4320) <= not(layer3_outputs(3887)) or (layer3_outputs(513));
    layer4_outputs(4321) <= not(layer3_outputs(8354));
    layer4_outputs(4322) <= (layer3_outputs(733)) and not (layer3_outputs(8809));
    layer4_outputs(4323) <= not(layer3_outputs(1734));
    layer4_outputs(4324) <= not(layer3_outputs(3805));
    layer4_outputs(4325) <= (layer3_outputs(5279)) xor (layer3_outputs(1997));
    layer4_outputs(4326) <= layer3_outputs(9594);
    layer4_outputs(4327) <= '0';
    layer4_outputs(4328) <= not(layer3_outputs(3904)) or (layer3_outputs(6477));
    layer4_outputs(4329) <= not(layer3_outputs(6044));
    layer4_outputs(4330) <= (layer3_outputs(7741)) and not (layer3_outputs(4858));
    layer4_outputs(4331) <= layer3_outputs(2157);
    layer4_outputs(4332) <= not(layer3_outputs(4331));
    layer4_outputs(4333) <= layer3_outputs(8845);
    layer4_outputs(4334) <= not(layer3_outputs(9953));
    layer4_outputs(4335) <= (layer3_outputs(3908)) xor (layer3_outputs(5993));
    layer4_outputs(4336) <= layer3_outputs(5073);
    layer4_outputs(4337) <= layer3_outputs(7313);
    layer4_outputs(4338) <= layer3_outputs(7717);
    layer4_outputs(4339) <= (layer3_outputs(3807)) xor (layer3_outputs(7874));
    layer4_outputs(4340) <= layer3_outputs(7035);
    layer4_outputs(4341) <= layer3_outputs(5242);
    layer4_outputs(4342) <= (layer3_outputs(3378)) and not (layer3_outputs(8787));
    layer4_outputs(4343) <= not((layer3_outputs(4995)) xor (layer3_outputs(8134)));
    layer4_outputs(4344) <= layer3_outputs(7123);
    layer4_outputs(4345) <= not(layer3_outputs(2747)) or (layer3_outputs(6018));
    layer4_outputs(4346) <= not(layer3_outputs(3270));
    layer4_outputs(4347) <= layer3_outputs(3698);
    layer4_outputs(4348) <= (layer3_outputs(6951)) xor (layer3_outputs(3054));
    layer4_outputs(4349) <= not((layer3_outputs(1502)) or (layer3_outputs(8614)));
    layer4_outputs(4350) <= not(layer3_outputs(9145));
    layer4_outputs(4351) <= (layer3_outputs(3466)) xor (layer3_outputs(10000));
    layer4_outputs(4352) <= (layer3_outputs(8845)) and not (layer3_outputs(5251));
    layer4_outputs(4353) <= '0';
    layer4_outputs(4354) <= not((layer3_outputs(110)) xor (layer3_outputs(9170)));
    layer4_outputs(4355) <= not(layer3_outputs(4551));
    layer4_outputs(4356) <= (layer3_outputs(1993)) and not (layer3_outputs(3091));
    layer4_outputs(4357) <= (layer3_outputs(6547)) and not (layer3_outputs(10002));
    layer4_outputs(4358) <= layer3_outputs(3402);
    layer4_outputs(4359) <= not(layer3_outputs(5746)) or (layer3_outputs(5552));
    layer4_outputs(4360) <= not((layer3_outputs(3988)) xor (layer3_outputs(8448)));
    layer4_outputs(4361) <= layer3_outputs(1035);
    layer4_outputs(4362) <= layer3_outputs(802);
    layer4_outputs(4363) <= layer3_outputs(556);
    layer4_outputs(4364) <= layer3_outputs(1106);
    layer4_outputs(4365) <= (layer3_outputs(6288)) xor (layer3_outputs(510));
    layer4_outputs(4366) <= layer3_outputs(5828);
    layer4_outputs(4367) <= not(layer3_outputs(4948));
    layer4_outputs(4368) <= not((layer3_outputs(384)) xor (layer3_outputs(7728)));
    layer4_outputs(4369) <= (layer3_outputs(1276)) or (layer3_outputs(5674));
    layer4_outputs(4370) <= not(layer3_outputs(1140));
    layer4_outputs(4371) <= (layer3_outputs(4618)) or (layer3_outputs(2610));
    layer4_outputs(4372) <= layer3_outputs(9914);
    layer4_outputs(4373) <= (layer3_outputs(4752)) xor (layer3_outputs(976));
    layer4_outputs(4374) <= not((layer3_outputs(8640)) or (layer3_outputs(671)));
    layer4_outputs(4375) <= not(layer3_outputs(7475));
    layer4_outputs(4376) <= layer3_outputs(4002);
    layer4_outputs(4377) <= not(layer3_outputs(6072));
    layer4_outputs(4378) <= (layer3_outputs(4148)) and not (layer3_outputs(9312));
    layer4_outputs(4379) <= not(layer3_outputs(5648));
    layer4_outputs(4380) <= (layer3_outputs(80)) and not (layer3_outputs(4066));
    layer4_outputs(4381) <= (layer3_outputs(8632)) xor (layer3_outputs(1884));
    layer4_outputs(4382) <= layer3_outputs(1284);
    layer4_outputs(4383) <= not(layer3_outputs(1856));
    layer4_outputs(4384) <= not(layer3_outputs(2219));
    layer4_outputs(4385) <= not(layer3_outputs(4993)) or (layer3_outputs(3880));
    layer4_outputs(4386) <= not(layer3_outputs(2543));
    layer4_outputs(4387) <= layer3_outputs(4867);
    layer4_outputs(4388) <= not((layer3_outputs(4876)) and (layer3_outputs(1940)));
    layer4_outputs(4389) <= not(layer3_outputs(5873));
    layer4_outputs(4390) <= not(layer3_outputs(5553));
    layer4_outputs(4391) <= not(layer3_outputs(5594)) or (layer3_outputs(6009));
    layer4_outputs(4392) <= (layer3_outputs(2896)) xor (layer3_outputs(5622));
    layer4_outputs(4393) <= not(layer3_outputs(2137));
    layer4_outputs(4394) <= layer3_outputs(7543);
    layer4_outputs(4395) <= layer3_outputs(1391);
    layer4_outputs(4396) <= not((layer3_outputs(1302)) xor (layer3_outputs(9580)));
    layer4_outputs(4397) <= layer3_outputs(7754);
    layer4_outputs(4398) <= not(layer3_outputs(1150)) or (layer3_outputs(5402));
    layer4_outputs(4399) <= not(layer3_outputs(1758)) or (layer3_outputs(8897));
    layer4_outputs(4400) <= not(layer3_outputs(846)) or (layer3_outputs(8225));
    layer4_outputs(4401) <= layer3_outputs(2883);
    layer4_outputs(4402) <= layer3_outputs(5922);
    layer4_outputs(4403) <= (layer3_outputs(5213)) xor (layer3_outputs(8254));
    layer4_outputs(4404) <= layer3_outputs(1489);
    layer4_outputs(4405) <= (layer3_outputs(5050)) or (layer3_outputs(4772));
    layer4_outputs(4406) <= layer3_outputs(8280);
    layer4_outputs(4407) <= layer3_outputs(9771);
    layer4_outputs(4408) <= layer3_outputs(8095);
    layer4_outputs(4409) <= not((layer3_outputs(9811)) xor (layer3_outputs(6939)));
    layer4_outputs(4410) <= not(layer3_outputs(4498));
    layer4_outputs(4411) <= not((layer3_outputs(5024)) or (layer3_outputs(5740)));
    layer4_outputs(4412) <= (layer3_outputs(4806)) and (layer3_outputs(9537));
    layer4_outputs(4413) <= layer3_outputs(2300);
    layer4_outputs(4414) <= not(layer3_outputs(3175));
    layer4_outputs(4415) <= not(layer3_outputs(9039));
    layer4_outputs(4416) <= layer3_outputs(5502);
    layer4_outputs(4417) <= layer3_outputs(7038);
    layer4_outputs(4418) <= layer3_outputs(7352);
    layer4_outputs(4419) <= not(layer3_outputs(8721));
    layer4_outputs(4420) <= (layer3_outputs(9198)) and not (layer3_outputs(5356));
    layer4_outputs(4421) <= not(layer3_outputs(6307));
    layer4_outputs(4422) <= not((layer3_outputs(2372)) and (layer3_outputs(158)));
    layer4_outputs(4423) <= layer3_outputs(9394);
    layer4_outputs(4424) <= not(layer3_outputs(4005));
    layer4_outputs(4425) <= layer3_outputs(5773);
    layer4_outputs(4426) <= not((layer3_outputs(5713)) or (layer3_outputs(3672)));
    layer4_outputs(4427) <= layer3_outputs(351);
    layer4_outputs(4428) <= not(layer3_outputs(3121));
    layer4_outputs(4429) <= layer3_outputs(8316);
    layer4_outputs(4430) <= not(layer3_outputs(9527)) or (layer3_outputs(4903));
    layer4_outputs(4431) <= layer3_outputs(121);
    layer4_outputs(4432) <= layer3_outputs(9041);
    layer4_outputs(4433) <= layer3_outputs(2354);
    layer4_outputs(4434) <= (layer3_outputs(6320)) or (layer3_outputs(1985));
    layer4_outputs(4435) <= layer3_outputs(3525);
    layer4_outputs(4436) <= (layer3_outputs(661)) and not (layer3_outputs(6520));
    layer4_outputs(4437) <= layer3_outputs(7889);
    layer4_outputs(4438) <= not(layer3_outputs(1079));
    layer4_outputs(4439) <= layer3_outputs(7610);
    layer4_outputs(4440) <= (layer3_outputs(7034)) and (layer3_outputs(8105));
    layer4_outputs(4441) <= layer3_outputs(4120);
    layer4_outputs(4442) <= layer3_outputs(6167);
    layer4_outputs(4443) <= not(layer3_outputs(2997)) or (layer3_outputs(2677));
    layer4_outputs(4444) <= '0';
    layer4_outputs(4445) <= layer3_outputs(3579);
    layer4_outputs(4446) <= not((layer3_outputs(4826)) xor (layer3_outputs(4107)));
    layer4_outputs(4447) <= not((layer3_outputs(977)) and (layer3_outputs(5128)));
    layer4_outputs(4448) <= layer3_outputs(7641);
    layer4_outputs(4449) <= layer3_outputs(6304);
    layer4_outputs(4450) <= not(layer3_outputs(5773));
    layer4_outputs(4451) <= '0';
    layer4_outputs(4452) <= layer3_outputs(9787);
    layer4_outputs(4453) <= layer3_outputs(2750);
    layer4_outputs(4454) <= layer3_outputs(1342);
    layer4_outputs(4455) <= layer3_outputs(7436);
    layer4_outputs(4456) <= (layer3_outputs(307)) xor (layer3_outputs(6348));
    layer4_outputs(4457) <= not(layer3_outputs(8972));
    layer4_outputs(4458) <= (layer3_outputs(7194)) xor (layer3_outputs(5701));
    layer4_outputs(4459) <= not(layer3_outputs(680));
    layer4_outputs(4460) <= layer3_outputs(7740);
    layer4_outputs(4461) <= layer3_outputs(6569);
    layer4_outputs(4462) <= not((layer3_outputs(1107)) xor (layer3_outputs(6984)));
    layer4_outputs(4463) <= not(layer3_outputs(2460));
    layer4_outputs(4464) <= not(layer3_outputs(2034));
    layer4_outputs(4465) <= not(layer3_outputs(7816));
    layer4_outputs(4466) <= not(layer3_outputs(3193));
    layer4_outputs(4467) <= layer3_outputs(6203);
    layer4_outputs(4468) <= (layer3_outputs(4592)) and not (layer3_outputs(3929));
    layer4_outputs(4469) <= not(layer3_outputs(9510));
    layer4_outputs(4470) <= not(layer3_outputs(5703));
    layer4_outputs(4471) <= layer3_outputs(2222);
    layer4_outputs(4472) <= layer3_outputs(4989);
    layer4_outputs(4473) <= (layer3_outputs(6505)) and not (layer3_outputs(1209));
    layer4_outputs(4474) <= (layer3_outputs(471)) and not (layer3_outputs(6220));
    layer4_outputs(4475) <= not(layer3_outputs(859));
    layer4_outputs(4476) <= not(layer3_outputs(687));
    layer4_outputs(4477) <= layer3_outputs(3414);
    layer4_outputs(4478) <= not(layer3_outputs(6050));
    layer4_outputs(4479) <= not((layer3_outputs(118)) and (layer3_outputs(5758)));
    layer4_outputs(4480) <= not(layer3_outputs(5020));
    layer4_outputs(4481) <= not(layer3_outputs(7978));
    layer4_outputs(4482) <= (layer3_outputs(7339)) xor (layer3_outputs(3551));
    layer4_outputs(4483) <= not(layer3_outputs(7278));
    layer4_outputs(4484) <= (layer3_outputs(6647)) xor (layer3_outputs(3610));
    layer4_outputs(4485) <= (layer3_outputs(1471)) and not (layer3_outputs(7253));
    layer4_outputs(4486) <= (layer3_outputs(8597)) xor (layer3_outputs(2538));
    layer4_outputs(4487) <= (layer3_outputs(8233)) xor (layer3_outputs(4608));
    layer4_outputs(4488) <= not(layer3_outputs(5860));
    layer4_outputs(4489) <= not((layer3_outputs(208)) and (layer3_outputs(4698)));
    layer4_outputs(4490) <= not(layer3_outputs(7897));
    layer4_outputs(4491) <= not(layer3_outputs(8774));
    layer4_outputs(4492) <= not(layer3_outputs(1662));
    layer4_outputs(4493) <= '1';
    layer4_outputs(4494) <= layer3_outputs(1075);
    layer4_outputs(4495) <= '1';
    layer4_outputs(4496) <= layer3_outputs(6234);
    layer4_outputs(4497) <= (layer3_outputs(8477)) or (layer3_outputs(8892));
    layer4_outputs(4498) <= not((layer3_outputs(9086)) xor (layer3_outputs(7010)));
    layer4_outputs(4499) <= not(layer3_outputs(943));
    layer4_outputs(4500) <= layer3_outputs(7119);
    layer4_outputs(4501) <= (layer3_outputs(1976)) xor (layer3_outputs(4526));
    layer4_outputs(4502) <= not((layer3_outputs(2837)) xor (layer3_outputs(1055)));
    layer4_outputs(4503) <= (layer3_outputs(4040)) and not (layer3_outputs(3510));
    layer4_outputs(4504) <= not((layer3_outputs(8336)) or (layer3_outputs(7518)));
    layer4_outputs(4505) <= not((layer3_outputs(2215)) and (layer3_outputs(9435)));
    layer4_outputs(4506) <= layer3_outputs(2260);
    layer4_outputs(4507) <= not(layer3_outputs(4204));
    layer4_outputs(4508) <= not(layer3_outputs(2427));
    layer4_outputs(4509) <= not((layer3_outputs(6768)) and (layer3_outputs(851)));
    layer4_outputs(4510) <= (layer3_outputs(8718)) and not (layer3_outputs(6754));
    layer4_outputs(4511) <= layer3_outputs(1393);
    layer4_outputs(4512) <= layer3_outputs(4079);
    layer4_outputs(4513) <= not((layer3_outputs(4987)) or (layer3_outputs(4190)));
    layer4_outputs(4514) <= layer3_outputs(3409);
    layer4_outputs(4515) <= (layer3_outputs(1821)) xor (layer3_outputs(423));
    layer4_outputs(4516) <= (layer3_outputs(4736)) or (layer3_outputs(3909));
    layer4_outputs(4517) <= layer3_outputs(4374);
    layer4_outputs(4518) <= (layer3_outputs(2456)) and not (layer3_outputs(564));
    layer4_outputs(4519) <= not((layer3_outputs(9003)) and (layer3_outputs(4351)));
    layer4_outputs(4520) <= not(layer3_outputs(7455));
    layer4_outputs(4521) <= not(layer3_outputs(832));
    layer4_outputs(4522) <= not(layer3_outputs(1891));
    layer4_outputs(4523) <= not((layer3_outputs(2774)) and (layer3_outputs(3542)));
    layer4_outputs(4524) <= not(layer3_outputs(7127));
    layer4_outputs(4525) <= not(layer3_outputs(6953));
    layer4_outputs(4526) <= not((layer3_outputs(7379)) and (layer3_outputs(197)));
    layer4_outputs(4527) <= layer3_outputs(1999);
    layer4_outputs(4528) <= layer3_outputs(947);
    layer4_outputs(4529) <= layer3_outputs(1519);
    layer4_outputs(4530) <= layer3_outputs(4743);
    layer4_outputs(4531) <= not(layer3_outputs(447)) or (layer3_outputs(5383));
    layer4_outputs(4532) <= not((layer3_outputs(9799)) and (layer3_outputs(9004)));
    layer4_outputs(4533) <= layer3_outputs(4005);
    layer4_outputs(4534) <= (layer3_outputs(8541)) xor (layer3_outputs(8649));
    layer4_outputs(4535) <= not(layer3_outputs(10149));
    layer4_outputs(4536) <= layer3_outputs(4904);
    layer4_outputs(4537) <= not(layer3_outputs(7296)) or (layer3_outputs(3772));
    layer4_outputs(4538) <= (layer3_outputs(9767)) or (layer3_outputs(4983));
    layer4_outputs(4539) <= layer3_outputs(8652);
    layer4_outputs(4540) <= (layer3_outputs(6405)) and (layer3_outputs(8853));
    layer4_outputs(4541) <= not(layer3_outputs(1193)) or (layer3_outputs(5867));
    layer4_outputs(4542) <= (layer3_outputs(2395)) xor (layer3_outputs(6589));
    layer4_outputs(4543) <= not(layer3_outputs(4099)) or (layer3_outputs(3405));
    layer4_outputs(4544) <= not((layer3_outputs(770)) xor (layer3_outputs(746)));
    layer4_outputs(4545) <= layer3_outputs(3522);
    layer4_outputs(4546) <= (layer3_outputs(3809)) xor (layer3_outputs(1620));
    layer4_outputs(4547) <= not(layer3_outputs(7654)) or (layer3_outputs(1780));
    layer4_outputs(4548) <= (layer3_outputs(8079)) and not (layer3_outputs(8444));
    layer4_outputs(4549) <= not(layer3_outputs(6169));
    layer4_outputs(4550) <= not(layer3_outputs(9026));
    layer4_outputs(4551) <= not(layer3_outputs(7761)) or (layer3_outputs(5878));
    layer4_outputs(4552) <= not(layer3_outputs(1907));
    layer4_outputs(4553) <= layer3_outputs(1496);
    layer4_outputs(4554) <= (layer3_outputs(1803)) and (layer3_outputs(6592));
    layer4_outputs(4555) <= layer3_outputs(2348);
    layer4_outputs(4556) <= (layer3_outputs(1095)) or (layer3_outputs(6661));
    layer4_outputs(4557) <= (layer3_outputs(4622)) and (layer3_outputs(3245));
    layer4_outputs(4558) <= not(layer3_outputs(6541));
    layer4_outputs(4559) <= (layer3_outputs(7509)) xor (layer3_outputs(9390));
    layer4_outputs(4560) <= layer3_outputs(1438);
    layer4_outputs(4561) <= (layer3_outputs(2892)) or (layer3_outputs(6312));
    layer4_outputs(4562) <= not(layer3_outputs(6171));
    layer4_outputs(4563) <= (layer3_outputs(2787)) and not (layer3_outputs(7580));
    layer4_outputs(4564) <= layer3_outputs(4693);
    layer4_outputs(4565) <= not((layer3_outputs(3615)) xor (layer3_outputs(8933)));
    layer4_outputs(4566) <= (layer3_outputs(4781)) and (layer3_outputs(682));
    layer4_outputs(4567) <= not(layer3_outputs(8384));
    layer4_outputs(4568) <= (layer3_outputs(8442)) or (layer3_outputs(4250));
    layer4_outputs(4569) <= (layer3_outputs(3106)) and (layer3_outputs(2622));
    layer4_outputs(4570) <= layer3_outputs(2664);
    layer4_outputs(4571) <= not(layer3_outputs(3073)) or (layer3_outputs(3642));
    layer4_outputs(4572) <= not(layer3_outputs(1776)) or (layer3_outputs(8143));
    layer4_outputs(4573) <= (layer3_outputs(8025)) xor (layer3_outputs(6763));
    layer4_outputs(4574) <= not(layer3_outputs(9201)) or (layer3_outputs(8400));
    layer4_outputs(4575) <= not(layer3_outputs(3302)) or (layer3_outputs(8288));
    layer4_outputs(4576) <= (layer3_outputs(9306)) and (layer3_outputs(9955));
    layer4_outputs(4577) <= not(layer3_outputs(8668));
    layer4_outputs(4578) <= layer3_outputs(5627);
    layer4_outputs(4579) <= layer3_outputs(3185);
    layer4_outputs(4580) <= layer3_outputs(9841);
    layer4_outputs(4581) <= not((layer3_outputs(5649)) xor (layer3_outputs(1683)));
    layer4_outputs(4582) <= not((layer3_outputs(3620)) xor (layer3_outputs(1513)));
    layer4_outputs(4583) <= not(layer3_outputs(8687));
    layer4_outputs(4584) <= not(layer3_outputs(1716));
    layer4_outputs(4585) <= not(layer3_outputs(6755));
    layer4_outputs(4586) <= not(layer3_outputs(45));
    layer4_outputs(4587) <= '0';
    layer4_outputs(4588) <= layer3_outputs(5396);
    layer4_outputs(4589) <= layer3_outputs(8561);
    layer4_outputs(4590) <= not((layer3_outputs(6133)) xor (layer3_outputs(612)));
    layer4_outputs(4591) <= layer3_outputs(527);
    layer4_outputs(4592) <= layer3_outputs(5102);
    layer4_outputs(4593) <= (layer3_outputs(1632)) and not (layer3_outputs(5700));
    layer4_outputs(4594) <= not(layer3_outputs(3994));
    layer4_outputs(4595) <= not(layer3_outputs(3539));
    layer4_outputs(4596) <= (layer3_outputs(7456)) and (layer3_outputs(2029));
    layer4_outputs(4597) <= not((layer3_outputs(184)) and (layer3_outputs(5537)));
    layer4_outputs(4598) <= not(layer3_outputs(1814));
    layer4_outputs(4599) <= (layer3_outputs(3192)) xor (layer3_outputs(4680));
    layer4_outputs(4600) <= not(layer3_outputs(7372));
    layer4_outputs(4601) <= layer3_outputs(7024);
    layer4_outputs(4602) <= layer3_outputs(1595);
    layer4_outputs(4603) <= layer3_outputs(937);
    layer4_outputs(4604) <= (layer3_outputs(9816)) xor (layer3_outputs(1580));
    layer4_outputs(4605) <= not(layer3_outputs(4039));
    layer4_outputs(4606) <= not((layer3_outputs(1134)) xor (layer3_outputs(834)));
    layer4_outputs(4607) <= (layer3_outputs(5342)) and (layer3_outputs(7137));
    layer4_outputs(4608) <= not(layer3_outputs(2166));
    layer4_outputs(4609) <= not(layer3_outputs(7465));
    layer4_outputs(4610) <= (layer3_outputs(7776)) and not (layer3_outputs(192));
    layer4_outputs(4611) <= not((layer3_outputs(5676)) and (layer3_outputs(6721)));
    layer4_outputs(4612) <= (layer3_outputs(4382)) and (layer3_outputs(7824));
    layer4_outputs(4613) <= not((layer3_outputs(225)) xor (layer3_outputs(5163)));
    layer4_outputs(4614) <= not(layer3_outputs(2854)) or (layer3_outputs(9088));
    layer4_outputs(4615) <= layer3_outputs(2659);
    layer4_outputs(4616) <= not(layer3_outputs(3672));
    layer4_outputs(4617) <= (layer3_outputs(7040)) and not (layer3_outputs(5996));
    layer4_outputs(4618) <= layer3_outputs(9293);
    layer4_outputs(4619) <= layer3_outputs(4308);
    layer4_outputs(4620) <= '0';
    layer4_outputs(4621) <= not(layer3_outputs(2826)) or (layer3_outputs(3521));
    layer4_outputs(4622) <= not(layer3_outputs(9395));
    layer4_outputs(4623) <= layer3_outputs(4054);
    layer4_outputs(4624) <= not((layer3_outputs(6954)) and (layer3_outputs(2932)));
    layer4_outputs(4625) <= (layer3_outputs(6236)) and not (layer3_outputs(1677));
    layer4_outputs(4626) <= not(layer3_outputs(2218));
    layer4_outputs(4627) <= not(layer3_outputs(712));
    layer4_outputs(4628) <= not((layer3_outputs(8408)) and (layer3_outputs(6266)));
    layer4_outputs(4629) <= layer3_outputs(2458);
    layer4_outputs(4630) <= (layer3_outputs(6708)) and (layer3_outputs(1521));
    layer4_outputs(4631) <= (layer3_outputs(1726)) and not (layer3_outputs(4560));
    layer4_outputs(4632) <= not(layer3_outputs(3463));
    layer4_outputs(4633) <= layer3_outputs(6557);
    layer4_outputs(4634) <= (layer3_outputs(6719)) and not (layer3_outputs(629));
    layer4_outputs(4635) <= (layer3_outputs(399)) xor (layer3_outputs(1049));
    layer4_outputs(4636) <= not(layer3_outputs(6125));
    layer4_outputs(4637) <= layer3_outputs(7156);
    layer4_outputs(4638) <= not(layer3_outputs(3115));
    layer4_outputs(4639) <= not(layer3_outputs(8499));
    layer4_outputs(4640) <= layer3_outputs(9415);
    layer4_outputs(4641) <= layer3_outputs(1866);
    layer4_outputs(4642) <= not(layer3_outputs(1947)) or (layer3_outputs(3018));
    layer4_outputs(4643) <= (layer3_outputs(1191)) and not (layer3_outputs(3251));
    layer4_outputs(4644) <= not((layer3_outputs(640)) or (layer3_outputs(4305)));
    layer4_outputs(4645) <= layer3_outputs(8744);
    layer4_outputs(4646) <= not(layer3_outputs(8126)) or (layer3_outputs(10122));
    layer4_outputs(4647) <= (layer3_outputs(8594)) xor (layer3_outputs(9017));
    layer4_outputs(4648) <= layer3_outputs(9692);
    layer4_outputs(4649) <= (layer3_outputs(6497)) xor (layer3_outputs(9327));
    layer4_outputs(4650) <= not(layer3_outputs(6587));
    layer4_outputs(4651) <= (layer3_outputs(3667)) or (layer3_outputs(8979));
    layer4_outputs(4652) <= (layer3_outputs(3195)) and not (layer3_outputs(7160));
    layer4_outputs(4653) <= not(layer3_outputs(5486));
    layer4_outputs(4654) <= not(layer3_outputs(4237));
    layer4_outputs(4655) <= layer3_outputs(3703);
    layer4_outputs(4656) <= not(layer3_outputs(3729)) or (layer3_outputs(310));
    layer4_outputs(4657) <= not((layer3_outputs(2904)) and (layer3_outputs(9245)));
    layer4_outputs(4658) <= layer3_outputs(2590);
    layer4_outputs(4659) <= not((layer3_outputs(5522)) and (layer3_outputs(630)));
    layer4_outputs(4660) <= layer3_outputs(6077);
    layer4_outputs(4661) <= not((layer3_outputs(2789)) xor (layer3_outputs(1814)));
    layer4_outputs(4662) <= (layer3_outputs(6725)) or (layer3_outputs(9517));
    layer4_outputs(4663) <= (layer3_outputs(4498)) and not (layer3_outputs(9820));
    layer4_outputs(4664) <= (layer3_outputs(6978)) or (layer3_outputs(6724));
    layer4_outputs(4665) <= (layer3_outputs(9269)) and (layer3_outputs(3305));
    layer4_outputs(4666) <= not(layer3_outputs(665));
    layer4_outputs(4667) <= not(layer3_outputs(6559)) or (layer3_outputs(5194));
    layer4_outputs(4668) <= (layer3_outputs(2527)) and not (layer3_outputs(1579));
    layer4_outputs(4669) <= (layer3_outputs(2177)) xor (layer3_outputs(7898));
    layer4_outputs(4670) <= not(layer3_outputs(1738)) or (layer3_outputs(8395));
    layer4_outputs(4671) <= layer3_outputs(5220);
    layer4_outputs(4672) <= layer3_outputs(8777);
    layer4_outputs(4673) <= layer3_outputs(7611);
    layer4_outputs(4674) <= layer3_outputs(7872);
    layer4_outputs(4675) <= layer3_outputs(3590);
    layer4_outputs(4676) <= layer3_outputs(8943);
    layer4_outputs(4677) <= '0';
    layer4_outputs(4678) <= not(layer3_outputs(4485));
    layer4_outputs(4679) <= not(layer3_outputs(7025));
    layer4_outputs(4680) <= not((layer3_outputs(4264)) xor (layer3_outputs(9156)));
    layer4_outputs(4681) <= layer3_outputs(9885);
    layer4_outputs(4682) <= layer3_outputs(8730);
    layer4_outputs(4683) <= layer3_outputs(2900);
    layer4_outputs(4684) <= layer3_outputs(5595);
    layer4_outputs(4685) <= not((layer3_outputs(8078)) or (layer3_outputs(5971)));
    layer4_outputs(4686) <= not((layer3_outputs(8781)) xor (layer3_outputs(10182)));
    layer4_outputs(4687) <= not((layer3_outputs(7817)) xor (layer3_outputs(2253)));
    layer4_outputs(4688) <= not((layer3_outputs(1667)) xor (layer3_outputs(9579)));
    layer4_outputs(4689) <= not(layer3_outputs(9937));
    layer4_outputs(4690) <= layer3_outputs(2743);
    layer4_outputs(4691) <= (layer3_outputs(5567)) and (layer3_outputs(3628));
    layer4_outputs(4692) <= (layer3_outputs(2785)) xor (layer3_outputs(9437));
    layer4_outputs(4693) <= not(layer3_outputs(4727));
    layer4_outputs(4694) <= (layer3_outputs(9171)) and not (layer3_outputs(3032));
    layer4_outputs(4695) <= layer3_outputs(3170);
    layer4_outputs(4696) <= (layer3_outputs(6969)) xor (layer3_outputs(3483));
    layer4_outputs(4697) <= not(layer3_outputs(5587));
    layer4_outputs(4698) <= layer3_outputs(476);
    layer4_outputs(4699) <= not(layer3_outputs(6147)) or (layer3_outputs(4725));
    layer4_outputs(4700) <= layer3_outputs(10190);
    layer4_outputs(4701) <= not((layer3_outputs(8235)) and (layer3_outputs(5325)));
    layer4_outputs(4702) <= layer3_outputs(7251);
    layer4_outputs(4703) <= '1';
    layer4_outputs(4704) <= layer3_outputs(2032);
    layer4_outputs(4705) <= layer3_outputs(5244);
    layer4_outputs(4706) <= (layer3_outputs(8151)) and not (layer3_outputs(4859));
    layer4_outputs(4707) <= (layer3_outputs(9443)) or (layer3_outputs(808));
    layer4_outputs(4708) <= not(layer3_outputs(8608));
    layer4_outputs(4709) <= (layer3_outputs(3446)) and (layer3_outputs(4307));
    layer4_outputs(4710) <= layer3_outputs(6363);
    layer4_outputs(4711) <= layer3_outputs(5202);
    layer4_outputs(4712) <= (layer3_outputs(5404)) and not (layer3_outputs(9262));
    layer4_outputs(4713) <= not(layer3_outputs(247));
    layer4_outputs(4714) <= layer3_outputs(5216);
    layer4_outputs(4715) <= layer3_outputs(9855);
    layer4_outputs(4716) <= not(layer3_outputs(2774));
    layer4_outputs(4717) <= (layer3_outputs(6507)) and not (layer3_outputs(3897));
    layer4_outputs(4718) <= not(layer3_outputs(9798));
    layer4_outputs(4719) <= (layer3_outputs(7055)) or (layer3_outputs(8758));
    layer4_outputs(4720) <= (layer3_outputs(818)) or (layer3_outputs(2362));
    layer4_outputs(4721) <= layer3_outputs(8671);
    layer4_outputs(4722) <= not((layer3_outputs(9217)) xor (layer3_outputs(9331)));
    layer4_outputs(4723) <= layer3_outputs(9294);
    layer4_outputs(4724) <= layer3_outputs(5800);
    layer4_outputs(4725) <= (layer3_outputs(5322)) and not (layer3_outputs(5743));
    layer4_outputs(4726) <= layer3_outputs(9232);
    layer4_outputs(4727) <= layer3_outputs(4775);
    layer4_outputs(4728) <= not(layer3_outputs(2598));
    layer4_outputs(4729) <= not(layer3_outputs(9810));
    layer4_outputs(4730) <= layer3_outputs(7709);
    layer4_outputs(4731) <= not((layer3_outputs(8837)) xor (layer3_outputs(4113)));
    layer4_outputs(4732) <= layer3_outputs(4972);
    layer4_outputs(4733) <= '0';
    layer4_outputs(4734) <= layer3_outputs(7734);
    layer4_outputs(4735) <= (layer3_outputs(7407)) and (layer3_outputs(7243));
    layer4_outputs(4736) <= layer3_outputs(5728);
    layer4_outputs(4737) <= layer3_outputs(6145);
    layer4_outputs(4738) <= not((layer3_outputs(7913)) or (layer3_outputs(7416)));
    layer4_outputs(4739) <= not((layer3_outputs(3861)) xor (layer3_outputs(1896)));
    layer4_outputs(4740) <= layer3_outputs(6431);
    layer4_outputs(4741) <= (layer3_outputs(5033)) and (layer3_outputs(6896));
    layer4_outputs(4742) <= layer3_outputs(2030);
    layer4_outputs(4743) <= not((layer3_outputs(6407)) xor (layer3_outputs(697)));
    layer4_outputs(4744) <= not(layer3_outputs(5421)) or (layer3_outputs(4811));
    layer4_outputs(4745) <= (layer3_outputs(6420)) xor (layer3_outputs(9535));
    layer4_outputs(4746) <= not(layer3_outputs(4506)) or (layer3_outputs(778));
    layer4_outputs(4747) <= (layer3_outputs(181)) and (layer3_outputs(1351));
    layer4_outputs(4748) <= (layer3_outputs(907)) and (layer3_outputs(8701));
    layer4_outputs(4749) <= not(layer3_outputs(5007));
    layer4_outputs(4750) <= not(layer3_outputs(9853)) or (layer3_outputs(1836));
    layer4_outputs(4751) <= (layer3_outputs(6843)) xor (layer3_outputs(5646));
    layer4_outputs(4752) <= (layer3_outputs(5456)) and not (layer3_outputs(7601));
    layer4_outputs(4753) <= (layer3_outputs(9289)) and not (layer3_outputs(2193));
    layer4_outputs(4754) <= not(layer3_outputs(6826));
    layer4_outputs(4755) <= (layer3_outputs(7116)) and not (layer3_outputs(6681));
    layer4_outputs(4756) <= layer3_outputs(4080);
    layer4_outputs(4757) <= not(layer3_outputs(2912)) or (layer3_outputs(100));
    layer4_outputs(4758) <= layer3_outputs(3589);
    layer4_outputs(4759) <= layer3_outputs(1583);
    layer4_outputs(4760) <= layer3_outputs(4263);
    layer4_outputs(4761) <= not(layer3_outputs(5287)) or (layer3_outputs(362));
    layer4_outputs(4762) <= layer3_outputs(4478);
    layer4_outputs(4763) <= not(layer3_outputs(5343)) or (layer3_outputs(7998));
    layer4_outputs(4764) <= not(layer3_outputs(693)) or (layer3_outputs(3256));
    layer4_outputs(4765) <= not((layer3_outputs(5300)) and (layer3_outputs(8651)));
    layer4_outputs(4766) <= not(layer3_outputs(1232));
    layer4_outputs(4767) <= (layer3_outputs(3651)) xor (layer3_outputs(6380));
    layer4_outputs(4768) <= not((layer3_outputs(316)) xor (layer3_outputs(6241)));
    layer4_outputs(4769) <= (layer3_outputs(5845)) xor (layer3_outputs(1568));
    layer4_outputs(4770) <= not((layer3_outputs(1471)) and (layer3_outputs(7179)));
    layer4_outputs(4771) <= layer3_outputs(157);
    layer4_outputs(4772) <= not((layer3_outputs(8103)) xor (layer3_outputs(2405)));
    layer4_outputs(4773) <= not(layer3_outputs(5918)) or (layer3_outputs(9754));
    layer4_outputs(4774) <= not(layer3_outputs(2433));
    layer4_outputs(4775) <= not(layer3_outputs(456));
    layer4_outputs(4776) <= not((layer3_outputs(3296)) xor (layer3_outputs(2945)));
    layer4_outputs(4777) <= not((layer3_outputs(3949)) xor (layer3_outputs(253)));
    layer4_outputs(4778) <= not(layer3_outputs(689));
    layer4_outputs(4779) <= not((layer3_outputs(2560)) or (layer3_outputs(7941)));
    layer4_outputs(4780) <= layer3_outputs(6875);
    layer4_outputs(4781) <= layer3_outputs(3883);
    layer4_outputs(4782) <= not(layer3_outputs(8457)) or (layer3_outputs(5978));
    layer4_outputs(4783) <= (layer3_outputs(296)) and not (layer3_outputs(3656));
    layer4_outputs(4784) <= not(layer3_outputs(4679));
    layer4_outputs(4785) <= not((layer3_outputs(8775)) xor (layer3_outputs(3156)));
    layer4_outputs(4786) <= not(layer3_outputs(7645));
    layer4_outputs(4787) <= not((layer3_outputs(9827)) xor (layer3_outputs(328)));
    layer4_outputs(4788) <= not((layer3_outputs(5038)) xor (layer3_outputs(6314)));
    layer4_outputs(4789) <= not((layer3_outputs(3101)) xor (layer3_outputs(9093)));
    layer4_outputs(4790) <= layer3_outputs(1114);
    layer4_outputs(4791) <= not(layer3_outputs(9990));
    layer4_outputs(4792) <= not((layer3_outputs(1474)) xor (layer3_outputs(1812)));
    layer4_outputs(4793) <= layer3_outputs(3125);
    layer4_outputs(4794) <= (layer3_outputs(1020)) and not (layer3_outputs(5552));
    layer4_outputs(4795) <= (layer3_outputs(7275)) or (layer3_outputs(2994));
    layer4_outputs(4796) <= layer3_outputs(8784);
    layer4_outputs(4797) <= layer3_outputs(8214);
    layer4_outputs(4798) <= layer3_outputs(3703);
    layer4_outputs(4799) <= layer3_outputs(9530);
    layer4_outputs(4800) <= (layer3_outputs(8553)) and (layer3_outputs(10226));
    layer4_outputs(4801) <= not((layer3_outputs(5061)) and (layer3_outputs(9748)));
    layer4_outputs(4802) <= (layer3_outputs(8114)) xor (layer3_outputs(7513));
    layer4_outputs(4803) <= not(layer3_outputs(3867));
    layer4_outputs(4804) <= not((layer3_outputs(9633)) or (layer3_outputs(7910)));
    layer4_outputs(4805) <= not(layer3_outputs(2333));
    layer4_outputs(4806) <= layer3_outputs(9207);
    layer4_outputs(4807) <= not((layer3_outputs(6059)) xor (layer3_outputs(3712)));
    layer4_outputs(4808) <= not(layer3_outputs(9370));
    layer4_outputs(4809) <= not(layer3_outputs(2081)) or (layer3_outputs(7855));
    layer4_outputs(4810) <= not(layer3_outputs(1645));
    layer4_outputs(4811) <= not((layer3_outputs(5372)) or (layer3_outputs(546)));
    layer4_outputs(4812) <= (layer3_outputs(7092)) and (layer3_outputs(4225));
    layer4_outputs(4813) <= (layer3_outputs(5590)) and (layer3_outputs(8691));
    layer4_outputs(4814) <= (layer3_outputs(5302)) and not (layer3_outputs(5190));
    layer4_outputs(4815) <= not(layer3_outputs(8746)) or (layer3_outputs(987));
    layer4_outputs(4816) <= (layer3_outputs(2481)) and not (layer3_outputs(3028));
    layer4_outputs(4817) <= not((layer3_outputs(3662)) xor (layer3_outputs(1056)));
    layer4_outputs(4818) <= not(layer3_outputs(4234));
    layer4_outputs(4819) <= (layer3_outputs(1208)) or (layer3_outputs(7637));
    layer4_outputs(4820) <= not((layer3_outputs(5353)) xor (layer3_outputs(4322)));
    layer4_outputs(4821) <= (layer3_outputs(8761)) and not (layer3_outputs(443));
    layer4_outputs(4822) <= (layer3_outputs(10133)) and (layer3_outputs(2972));
    layer4_outputs(4823) <= layer3_outputs(10028);
    layer4_outputs(4824) <= layer3_outputs(2295);
    layer4_outputs(4825) <= layer3_outputs(812);
    layer4_outputs(4826) <= not((layer3_outputs(135)) xor (layer3_outputs(3426)));
    layer4_outputs(4827) <= layer3_outputs(4978);
    layer4_outputs(4828) <= (layer3_outputs(4004)) and (layer3_outputs(3512));
    layer4_outputs(4829) <= (layer3_outputs(2494)) and (layer3_outputs(8594));
    layer4_outputs(4830) <= not((layer3_outputs(2036)) xor (layer3_outputs(7887)));
    layer4_outputs(4831) <= layer3_outputs(9653);
    layer4_outputs(4832) <= not(layer3_outputs(6443)) or (layer3_outputs(2908));
    layer4_outputs(4833) <= not(layer3_outputs(365)) or (layer3_outputs(6547));
    layer4_outputs(4834) <= not(layer3_outputs(1886));
    layer4_outputs(4835) <= not(layer3_outputs(4570));
    layer4_outputs(4836) <= not(layer3_outputs(4016));
    layer4_outputs(4837) <= not((layer3_outputs(1963)) or (layer3_outputs(2734)));
    layer4_outputs(4838) <= not(layer3_outputs(4326));
    layer4_outputs(4839) <= not(layer3_outputs(2180));
    layer4_outputs(4840) <= not(layer3_outputs(6593));
    layer4_outputs(4841) <= layer3_outputs(8810);
    layer4_outputs(4842) <= not((layer3_outputs(7649)) xor (layer3_outputs(8437)));
    layer4_outputs(4843) <= (layer3_outputs(3461)) and (layer3_outputs(9529));
    layer4_outputs(4844) <= not(layer3_outputs(2440));
    layer4_outputs(4845) <= not(layer3_outputs(1108));
    layer4_outputs(4846) <= (layer3_outputs(9181)) xor (layer3_outputs(8710));
    layer4_outputs(4847) <= layer3_outputs(2435);
    layer4_outputs(4848) <= (layer3_outputs(2766)) and not (layer3_outputs(1553));
    layer4_outputs(4849) <= '1';
    layer4_outputs(4850) <= layer3_outputs(7877);
    layer4_outputs(4851) <= not(layer3_outputs(3298));
    layer4_outputs(4852) <= (layer3_outputs(3982)) and not (layer3_outputs(2464));
    layer4_outputs(4853) <= layer3_outputs(6908);
    layer4_outputs(4854) <= not((layer3_outputs(2436)) or (layer3_outputs(4944)));
    layer4_outputs(4855) <= not((layer3_outputs(722)) xor (layer3_outputs(3370)));
    layer4_outputs(4856) <= not((layer3_outputs(8464)) or (layer3_outputs(4389)));
    layer4_outputs(4857) <= (layer3_outputs(9568)) or (layer3_outputs(2402));
    layer4_outputs(4858) <= (layer3_outputs(3226)) and not (layer3_outputs(7172));
    layer4_outputs(4859) <= (layer3_outputs(8201)) and (layer3_outputs(8723));
    layer4_outputs(4860) <= not((layer3_outputs(8506)) and (layer3_outputs(3295)));
    layer4_outputs(4861) <= (layer3_outputs(3345)) and (layer3_outputs(9101));
    layer4_outputs(4862) <= layer3_outputs(7561);
    layer4_outputs(4863) <= layer3_outputs(3325);
    layer4_outputs(4864) <= not(layer3_outputs(8754));
    layer4_outputs(4865) <= (layer3_outputs(793)) xor (layer3_outputs(807));
    layer4_outputs(4866) <= (layer3_outputs(4281)) and not (layer3_outputs(255));
    layer4_outputs(4867) <= not(layer3_outputs(2605));
    layer4_outputs(4868) <= not((layer3_outputs(8658)) xor (layer3_outputs(1786)));
    layer4_outputs(4869) <= layer3_outputs(6385);
    layer4_outputs(4870) <= not(layer3_outputs(2860)) or (layer3_outputs(7715));
    layer4_outputs(4871) <= not(layer3_outputs(8179));
    layer4_outputs(4872) <= (layer3_outputs(713)) xor (layer3_outputs(4560));
    layer4_outputs(4873) <= not((layer3_outputs(2121)) xor (layer3_outputs(4969)));
    layer4_outputs(4874) <= layer3_outputs(1944);
    layer4_outputs(4875) <= not(layer3_outputs(7602));
    layer4_outputs(4876) <= not((layer3_outputs(2376)) xor (layer3_outputs(6014)));
    layer4_outputs(4877) <= layer3_outputs(4539);
    layer4_outputs(4878) <= (layer3_outputs(1656)) xor (layer3_outputs(3255));
    layer4_outputs(4879) <= not(layer3_outputs(3280));
    layer4_outputs(4880) <= not(layer3_outputs(3217));
    layer4_outputs(4881) <= (layer3_outputs(9964)) xor (layer3_outputs(2738));
    layer4_outputs(4882) <= not(layer3_outputs(1117));
    layer4_outputs(4883) <= '0';
    layer4_outputs(4884) <= (layer3_outputs(1083)) and not (layer3_outputs(5215));
    layer4_outputs(4885) <= not(layer3_outputs(5452));
    layer4_outputs(4886) <= not((layer3_outputs(2283)) xor (layer3_outputs(10212)));
    layer4_outputs(4887) <= not(layer3_outputs(51));
    layer4_outputs(4888) <= not(layer3_outputs(6189));
    layer4_outputs(4889) <= layer3_outputs(3049);
    layer4_outputs(4890) <= not((layer3_outputs(7802)) or (layer3_outputs(9555)));
    layer4_outputs(4891) <= layer3_outputs(3601);
    layer4_outputs(4892) <= not((layer3_outputs(559)) and (layer3_outputs(6597)));
    layer4_outputs(4893) <= not(layer3_outputs(9690));
    layer4_outputs(4894) <= (layer3_outputs(299)) or (layer3_outputs(7106));
    layer4_outputs(4895) <= not((layer3_outputs(8328)) or (layer3_outputs(8489)));
    layer4_outputs(4896) <= layer3_outputs(8565);
    layer4_outputs(4897) <= (layer3_outputs(333)) and (layer3_outputs(6207));
    layer4_outputs(4898) <= (layer3_outputs(6389)) or (layer3_outputs(4960));
    layer4_outputs(4899) <= not((layer3_outputs(4411)) xor (layer3_outputs(2115)));
    layer4_outputs(4900) <= layer3_outputs(2174);
    layer4_outputs(4901) <= (layer3_outputs(3761)) and not (layer3_outputs(4426));
    layer4_outputs(4902) <= not(layer3_outputs(8397));
    layer4_outputs(4903) <= not(layer3_outputs(4404));
    layer4_outputs(4904) <= not(layer3_outputs(4321));
    layer4_outputs(4905) <= not(layer3_outputs(223));
    layer4_outputs(4906) <= layer3_outputs(3643);
    layer4_outputs(4907) <= (layer3_outputs(10179)) and (layer3_outputs(5763));
    layer4_outputs(4908) <= layer3_outputs(9826);
    layer4_outputs(4909) <= layer3_outputs(4247);
    layer4_outputs(4910) <= layer3_outputs(4495);
    layer4_outputs(4911) <= (layer3_outputs(382)) or (layer3_outputs(6353));
    layer4_outputs(4912) <= not(layer3_outputs(2117));
    layer4_outputs(4913) <= not(layer3_outputs(8796));
    layer4_outputs(4914) <= layer3_outputs(7554);
    layer4_outputs(4915) <= not((layer3_outputs(6098)) and (layer3_outputs(5984)));
    layer4_outputs(4916) <= (layer3_outputs(408)) xor (layer3_outputs(5306));
    layer4_outputs(4917) <= (layer3_outputs(6091)) or (layer3_outputs(9483));
    layer4_outputs(4918) <= layer3_outputs(577);
    layer4_outputs(4919) <= not(layer3_outputs(6273));
    layer4_outputs(4920) <= not((layer3_outputs(2754)) and (layer3_outputs(9525)));
    layer4_outputs(4921) <= not(layer3_outputs(1667));
    layer4_outputs(4922) <= not(layer3_outputs(1649)) or (layer3_outputs(6225));
    layer4_outputs(4923) <= not(layer3_outputs(6238)) or (layer3_outputs(6316));
    layer4_outputs(4924) <= not(layer3_outputs(1285));
    layer4_outputs(4925) <= (layer3_outputs(7947)) xor (layer3_outputs(2979));
    layer4_outputs(4926) <= '1';
    layer4_outputs(4927) <= not(layer3_outputs(4828));
    layer4_outputs(4928) <= layer3_outputs(1538);
    layer4_outputs(4929) <= not(layer3_outputs(8385));
    layer4_outputs(4930) <= not(layer3_outputs(6761)) or (layer3_outputs(7220));
    layer4_outputs(4931) <= not(layer3_outputs(5412)) or (layer3_outputs(5271));
    layer4_outputs(4932) <= not(layer3_outputs(9123));
    layer4_outputs(4933) <= '1';
    layer4_outputs(4934) <= layer3_outputs(4734);
    layer4_outputs(4935) <= (layer3_outputs(5170)) and not (layer3_outputs(7719));
    layer4_outputs(4936) <= (layer3_outputs(9531)) or (layer3_outputs(6064));
    layer4_outputs(4937) <= not((layer3_outputs(1591)) or (layer3_outputs(103)));
    layer4_outputs(4938) <= not(layer3_outputs(4352));
    layer4_outputs(4939) <= layer3_outputs(407);
    layer4_outputs(4940) <= not((layer3_outputs(7159)) xor (layer3_outputs(8429)));
    layer4_outputs(4941) <= layer3_outputs(8617);
    layer4_outputs(4942) <= not(layer3_outputs(4799));
    layer4_outputs(4943) <= not(layer3_outputs(468));
    layer4_outputs(4944) <= not(layer3_outputs(4133));
    layer4_outputs(4945) <= (layer3_outputs(4953)) xor (layer3_outputs(2251));
    layer4_outputs(4946) <= (layer3_outputs(286)) and not (layer3_outputs(2265));
    layer4_outputs(4947) <= (layer3_outputs(5470)) xor (layer3_outputs(7959));
    layer4_outputs(4948) <= not(layer3_outputs(7338));
    layer4_outputs(4949) <= layer3_outputs(4584);
    layer4_outputs(4950) <= layer3_outputs(3887);
    layer4_outputs(4951) <= not(layer3_outputs(3785)) or (layer3_outputs(85));
    layer4_outputs(4952) <= layer3_outputs(8314);
    layer4_outputs(4953) <= layer3_outputs(766);
    layer4_outputs(4954) <= not(layer3_outputs(1310));
    layer4_outputs(4955) <= (layer3_outputs(7479)) xor (layer3_outputs(3744));
    layer4_outputs(4956) <= layer3_outputs(4972);
    layer4_outputs(4957) <= not(layer3_outputs(8627));
    layer4_outputs(4958) <= '0';
    layer4_outputs(4959) <= not(layer3_outputs(5226));
    layer4_outputs(4960) <= (layer3_outputs(9076)) and (layer3_outputs(2749));
    layer4_outputs(4961) <= not(layer3_outputs(1088));
    layer4_outputs(4962) <= (layer3_outputs(10048)) and (layer3_outputs(8070));
    layer4_outputs(4963) <= layer3_outputs(5373);
    layer4_outputs(4964) <= (layer3_outputs(2550)) and not (layer3_outputs(3405));
    layer4_outputs(4965) <= layer3_outputs(9976);
    layer4_outputs(4966) <= (layer3_outputs(710)) xor (layer3_outputs(2792));
    layer4_outputs(4967) <= (layer3_outputs(1903)) and not (layer3_outputs(6511));
    layer4_outputs(4968) <= layer3_outputs(6065);
    layer4_outputs(4969) <= layer3_outputs(6309);
    layer4_outputs(4970) <= not((layer3_outputs(3586)) xor (layer3_outputs(885)));
    layer4_outputs(4971) <= not(layer3_outputs(2078)) or (layer3_outputs(10108));
    layer4_outputs(4972) <= not(layer3_outputs(5806));
    layer4_outputs(4973) <= not((layer3_outputs(5392)) xor (layer3_outputs(2979)));
    layer4_outputs(4974) <= not(layer3_outputs(10178)) or (layer3_outputs(1568));
    layer4_outputs(4975) <= (layer3_outputs(10167)) xor (layer3_outputs(4121));
    layer4_outputs(4976) <= not((layer3_outputs(6155)) xor (layer3_outputs(4347)));
    layer4_outputs(4977) <= not(layer3_outputs(5302));
    layer4_outputs(4978) <= (layer3_outputs(9153)) or (layer3_outputs(1254));
    layer4_outputs(4979) <= not((layer3_outputs(261)) xor (layer3_outputs(7131)));
    layer4_outputs(4980) <= (layer3_outputs(4162)) or (layer3_outputs(8829));
    layer4_outputs(4981) <= (layer3_outputs(5448)) and not (layer3_outputs(9660));
    layer4_outputs(4982) <= (layer3_outputs(9661)) and not (layer3_outputs(2790));
    layer4_outputs(4983) <= (layer3_outputs(9557)) xor (layer3_outputs(3385));
    layer4_outputs(4984) <= (layer3_outputs(3070)) and not (layer3_outputs(8625));
    layer4_outputs(4985) <= not((layer3_outputs(193)) and (layer3_outputs(5776)));
    layer4_outputs(4986) <= '0';
    layer4_outputs(4987) <= not((layer3_outputs(7033)) and (layer3_outputs(3239)));
    layer4_outputs(4988) <= (layer3_outputs(3163)) xor (layer3_outputs(10048));
    layer4_outputs(4989) <= (layer3_outputs(5784)) and not (layer3_outputs(3683));
    layer4_outputs(4990) <= not(layer3_outputs(6774));
    layer4_outputs(4991) <= not((layer3_outputs(1309)) xor (layer3_outputs(9520)));
    layer4_outputs(4992) <= '0';
    layer4_outputs(4993) <= layer3_outputs(5073);
    layer4_outputs(4994) <= layer3_outputs(8616);
    layer4_outputs(4995) <= not(layer3_outputs(8023));
    layer4_outputs(4996) <= layer3_outputs(4488);
    layer4_outputs(4997) <= not((layer3_outputs(6400)) xor (layer3_outputs(781)));
    layer4_outputs(4998) <= not(layer3_outputs(787));
    layer4_outputs(4999) <= layer3_outputs(9916);
    layer4_outputs(5000) <= '1';
    layer4_outputs(5001) <= not(layer3_outputs(4778));
    layer4_outputs(5002) <= layer3_outputs(5119);
    layer4_outputs(5003) <= not(layer3_outputs(9806));
    layer4_outputs(5004) <= not(layer3_outputs(8382));
    layer4_outputs(5005) <= not(layer3_outputs(1707));
    layer4_outputs(5006) <= not(layer3_outputs(2521));
    layer4_outputs(5007) <= layer3_outputs(4502);
    layer4_outputs(5008) <= (layer3_outputs(5978)) xor (layer3_outputs(10024));
    layer4_outputs(5009) <= not((layer3_outputs(6533)) or (layer3_outputs(8791)));
    layer4_outputs(5010) <= not((layer3_outputs(4240)) xor (layer3_outputs(7212)));
    layer4_outputs(5011) <= not((layer3_outputs(9274)) and (layer3_outputs(3156)));
    layer4_outputs(5012) <= layer3_outputs(5775);
    layer4_outputs(5013) <= not(layer3_outputs(4435));
    layer4_outputs(5014) <= layer3_outputs(4850);
    layer4_outputs(5015) <= not(layer3_outputs(4793));
    layer4_outputs(5016) <= not(layer3_outputs(3211));
    layer4_outputs(5017) <= not(layer3_outputs(9031));
    layer4_outputs(5018) <= (layer3_outputs(4516)) or (layer3_outputs(3453));
    layer4_outputs(5019) <= not(layer3_outputs(8473));
    layer4_outputs(5020) <= (layer3_outputs(4269)) and not (layer3_outputs(9444));
    layer4_outputs(5021) <= not(layer3_outputs(1120));
    layer4_outputs(5022) <= (layer3_outputs(9084)) and not (layer3_outputs(2207));
    layer4_outputs(5023) <= (layer3_outputs(6793)) and not (layer3_outputs(1733));
    layer4_outputs(5024) <= (layer3_outputs(3935)) xor (layer3_outputs(2468));
    layer4_outputs(5025) <= (layer3_outputs(6455)) or (layer3_outputs(2826));
    layer4_outputs(5026) <= not(layer3_outputs(7604));
    layer4_outputs(5027) <= layer3_outputs(1038);
    layer4_outputs(5028) <= (layer3_outputs(2416)) or (layer3_outputs(526));
    layer4_outputs(5029) <= (layer3_outputs(5965)) and not (layer3_outputs(2388));
    layer4_outputs(5030) <= not((layer3_outputs(2787)) or (layer3_outputs(6158)));
    layer4_outputs(5031) <= (layer3_outputs(5679)) xor (layer3_outputs(1547));
    layer4_outputs(5032) <= (layer3_outputs(3160)) and not (layer3_outputs(8431));
    layer4_outputs(5033) <= (layer3_outputs(7469)) xor (layer3_outputs(7690));
    layer4_outputs(5034) <= not(layer3_outputs(1597));
    layer4_outputs(5035) <= (layer3_outputs(5016)) xor (layer3_outputs(2243));
    layer4_outputs(5036) <= (layer3_outputs(2446)) and not (layer3_outputs(2986));
    layer4_outputs(5037) <= layer3_outputs(9071);
    layer4_outputs(5038) <= layer3_outputs(7502);
    layer4_outputs(5039) <= not(layer3_outputs(1727));
    layer4_outputs(5040) <= (layer3_outputs(7950)) xor (layer3_outputs(1982));
    layer4_outputs(5041) <= (layer3_outputs(2203)) xor (layer3_outputs(7350));
    layer4_outputs(5042) <= not((layer3_outputs(632)) xor (layer3_outputs(8891)));
    layer4_outputs(5043) <= not(layer3_outputs(1696));
    layer4_outputs(5044) <= not(layer3_outputs(2980));
    layer4_outputs(5045) <= (layer3_outputs(7387)) or (layer3_outputs(7879));
    layer4_outputs(5046) <= layer3_outputs(9532);
    layer4_outputs(5047) <= not(layer3_outputs(6302));
    layer4_outputs(5048) <= (layer3_outputs(740)) xor (layer3_outputs(5482));
    layer4_outputs(5049) <= layer3_outputs(3006);
    layer4_outputs(5050) <= layer3_outputs(1864);
    layer4_outputs(5051) <= (layer3_outputs(10104)) and (layer3_outputs(9108));
    layer4_outputs(5052) <= (layer3_outputs(9043)) and not (layer3_outputs(7288));
    layer4_outputs(5053) <= not(layer3_outputs(7676));
    layer4_outputs(5054) <= not((layer3_outputs(7721)) and (layer3_outputs(7079)));
    layer4_outputs(5055) <= (layer3_outputs(8378)) and (layer3_outputs(9543));
    layer4_outputs(5056) <= layer3_outputs(9597);
    layer4_outputs(5057) <= not((layer3_outputs(6915)) xor (layer3_outputs(8886)));
    layer4_outputs(5058) <= layer3_outputs(10057);
    layer4_outputs(5059) <= not(layer3_outputs(5252));
    layer4_outputs(5060) <= not(layer3_outputs(8422)) or (layer3_outputs(405));
    layer4_outputs(5061) <= not(layer3_outputs(2258)) or (layer3_outputs(9866));
    layer4_outputs(5062) <= not(layer3_outputs(7590));
    layer4_outputs(5063) <= layer3_outputs(2837);
    layer4_outputs(5064) <= (layer3_outputs(5774)) xor (layer3_outputs(1638));
    layer4_outputs(5065) <= not((layer3_outputs(6941)) xor (layer3_outputs(10210)));
    layer4_outputs(5066) <= (layer3_outputs(10185)) xor (layer3_outputs(3042));
    layer4_outputs(5067) <= not((layer3_outputs(9813)) or (layer3_outputs(10166)));
    layer4_outputs(5068) <= not(layer3_outputs(7549));
    layer4_outputs(5069) <= not(layer3_outputs(1523)) or (layer3_outputs(2493));
    layer4_outputs(5070) <= not((layer3_outputs(9731)) xor (layer3_outputs(1776)));
    layer4_outputs(5071) <= not(layer3_outputs(4829));
    layer4_outputs(5072) <= not((layer3_outputs(2105)) xor (layer3_outputs(6975)));
    layer4_outputs(5073) <= not((layer3_outputs(5968)) or (layer3_outputs(7792)));
    layer4_outputs(5074) <= not((layer3_outputs(8551)) xor (layer3_outputs(1883)));
    layer4_outputs(5075) <= (layer3_outputs(6258)) xor (layer3_outputs(1048));
    layer4_outputs(5076) <= not((layer3_outputs(2666)) and (layer3_outputs(7073)));
    layer4_outputs(5077) <= not(layer3_outputs(9544));
    layer4_outputs(5078) <= layer3_outputs(4928);
    layer4_outputs(5079) <= layer3_outputs(4323);
    layer4_outputs(5080) <= not((layer3_outputs(4943)) and (layer3_outputs(7380)));
    layer4_outputs(5081) <= not((layer3_outputs(3011)) and (layer3_outputs(9573)));
    layer4_outputs(5082) <= layer3_outputs(3730);
    layer4_outputs(5083) <= not((layer3_outputs(7286)) xor (layer3_outputs(7300)));
    layer4_outputs(5084) <= (layer3_outputs(10125)) and not (layer3_outputs(2385));
    layer4_outputs(5085) <= not((layer3_outputs(1665)) xor (layer3_outputs(417)));
    layer4_outputs(5086) <= not(layer3_outputs(1900)) or (layer3_outputs(1587));
    layer4_outputs(5087) <= (layer3_outputs(5626)) and not (layer3_outputs(9711));
    layer4_outputs(5088) <= layer3_outputs(3993);
    layer4_outputs(5089) <= layer3_outputs(7064);
    layer4_outputs(5090) <= not(layer3_outputs(3224));
    layer4_outputs(5091) <= not(layer3_outputs(449));
    layer4_outputs(5092) <= layer3_outputs(5054);
    layer4_outputs(5093) <= not((layer3_outputs(5200)) xor (layer3_outputs(7665)));
    layer4_outputs(5094) <= layer3_outputs(6198);
    layer4_outputs(5095) <= (layer3_outputs(7210)) xor (layer3_outputs(7027));
    layer4_outputs(5096) <= not(layer3_outputs(1700));
    layer4_outputs(5097) <= layer3_outputs(1759);
    layer4_outputs(5098) <= not(layer3_outputs(3799));
    layer4_outputs(5099) <= (layer3_outputs(847)) and not (layer3_outputs(4975));
    layer4_outputs(5100) <= layer3_outputs(2452);
    layer4_outputs(5101) <= not(layer3_outputs(4934)) or (layer3_outputs(1137));
    layer4_outputs(5102) <= not(layer3_outputs(4111));
    layer4_outputs(5103) <= not(layer3_outputs(1864));
    layer4_outputs(5104) <= layer3_outputs(3214);
    layer4_outputs(5105) <= layer3_outputs(6313);
    layer4_outputs(5106) <= not((layer3_outputs(772)) or (layer3_outputs(5066)));
    layer4_outputs(5107) <= not(layer3_outputs(7662));
    layer4_outputs(5108) <= not(layer3_outputs(5363)) or (layer3_outputs(163));
    layer4_outputs(5109) <= layer3_outputs(4974);
    layer4_outputs(5110) <= not(layer3_outputs(2736));
    layer4_outputs(5111) <= (layer3_outputs(891)) and (layer3_outputs(8048));
    layer4_outputs(5112) <= not((layer3_outputs(257)) xor (layer3_outputs(10193)));
    layer4_outputs(5113) <= not(layer3_outputs(2446));
    layer4_outputs(5114) <= not(layer3_outputs(5548)) or (layer3_outputs(2047));
    layer4_outputs(5115) <= not(layer3_outputs(1450));
    layer4_outputs(5116) <= not((layer3_outputs(1243)) or (layer3_outputs(5937)));
    layer4_outputs(5117) <= '1';
    layer4_outputs(5118) <= not((layer3_outputs(6790)) xor (layer3_outputs(10084)));
    layer4_outputs(5119) <= not(layer3_outputs(9760));
    layer4_outputs(5120) <= (layer3_outputs(2898)) and not (layer3_outputs(1758));
    layer4_outputs(5121) <= not(layer3_outputs(4892));
    layer4_outputs(5122) <= (layer3_outputs(5550)) and not (layer3_outputs(2591));
    layer4_outputs(5123) <= not(layer3_outputs(969));
    layer4_outputs(5124) <= not(layer3_outputs(4615));
    layer4_outputs(5125) <= '0';
    layer4_outputs(5126) <= not((layer3_outputs(9890)) xor (layer3_outputs(2454)));
    layer4_outputs(5127) <= layer3_outputs(1443);
    layer4_outputs(5128) <= not(layer3_outputs(7987));
    layer4_outputs(5129) <= not(layer3_outputs(9072));
    layer4_outputs(5130) <= layer3_outputs(10002);
    layer4_outputs(5131) <= not((layer3_outputs(6698)) xor (layer3_outputs(4831)));
    layer4_outputs(5132) <= (layer3_outputs(2823)) and (layer3_outputs(10115));
    layer4_outputs(5133) <= not((layer3_outputs(3107)) xor (layer3_outputs(6516)));
    layer4_outputs(5134) <= not(layer3_outputs(10133));
    layer4_outputs(5135) <= not(layer3_outputs(3208));
    layer4_outputs(5136) <= (layer3_outputs(7083)) xor (layer3_outputs(7435));
    layer4_outputs(5137) <= '0';
    layer4_outputs(5138) <= (layer3_outputs(6839)) xor (layer3_outputs(3707));
    layer4_outputs(5139) <= (layer3_outputs(5730)) and not (layer3_outputs(5561));
    layer4_outputs(5140) <= (layer3_outputs(5713)) and (layer3_outputs(7326));
    layer4_outputs(5141) <= layer3_outputs(131);
    layer4_outputs(5142) <= layer3_outputs(3783);
    layer4_outputs(5143) <= not(layer3_outputs(8243));
    layer4_outputs(5144) <= layer3_outputs(207);
    layer4_outputs(5145) <= layer3_outputs(7394);
    layer4_outputs(5146) <= not(layer3_outputs(4375));
    layer4_outputs(5147) <= (layer3_outputs(7026)) xor (layer3_outputs(3058));
    layer4_outputs(5148) <= not(layer3_outputs(9524));
    layer4_outputs(5149) <= (layer3_outputs(5337)) or (layer3_outputs(4802));
    layer4_outputs(5150) <= not((layer3_outputs(8012)) xor (layer3_outputs(970)));
    layer4_outputs(5151) <= (layer3_outputs(798)) or (layer3_outputs(9148));
    layer4_outputs(5152) <= not(layer3_outputs(8772));
    layer4_outputs(5153) <= layer3_outputs(6137);
    layer4_outputs(5154) <= layer3_outputs(6237);
    layer4_outputs(5155) <= not(layer3_outputs(9291));
    layer4_outputs(5156) <= (layer3_outputs(2305)) xor (layer3_outputs(3051));
    layer4_outputs(5157) <= not(layer3_outputs(649));
    layer4_outputs(5158) <= not(layer3_outputs(1088));
    layer4_outputs(5159) <= not(layer3_outputs(1111));
    layer4_outputs(5160) <= layer3_outputs(5849);
    layer4_outputs(5161) <= not((layer3_outputs(912)) xor (layer3_outputs(5479)));
    layer4_outputs(5162) <= not((layer3_outputs(4004)) xor (layer3_outputs(6584)));
    layer4_outputs(5163) <= (layer3_outputs(3213)) and not (layer3_outputs(7353));
    layer4_outputs(5164) <= not((layer3_outputs(5499)) or (layer3_outputs(5741)));
    layer4_outputs(5165) <= (layer3_outputs(7305)) and (layer3_outputs(4581));
    layer4_outputs(5166) <= '0';
    layer4_outputs(5167) <= (layer3_outputs(892)) and not (layer3_outputs(2503));
    layer4_outputs(5168) <= layer3_outputs(7087);
    layer4_outputs(5169) <= layer3_outputs(3);
    layer4_outputs(5170) <= not(layer3_outputs(1138));
    layer4_outputs(5171) <= layer3_outputs(3764);
    layer4_outputs(5172) <= not((layer3_outputs(1775)) and (layer3_outputs(950)));
    layer4_outputs(5173) <= not(layer3_outputs(4300));
    layer4_outputs(5174) <= layer3_outputs(8252);
    layer4_outputs(5175) <= layer3_outputs(9282);
    layer4_outputs(5176) <= not((layer3_outputs(8115)) or (layer3_outputs(8994)));
    layer4_outputs(5177) <= (layer3_outputs(8198)) and not (layer3_outputs(7623));
    layer4_outputs(5178) <= not((layer3_outputs(7084)) and (layer3_outputs(8449)));
    layer4_outputs(5179) <= not(layer3_outputs(7363));
    layer4_outputs(5180) <= (layer3_outputs(574)) and not (layer3_outputs(230));
    layer4_outputs(5181) <= not(layer3_outputs(3939));
    layer4_outputs(5182) <= layer3_outputs(3054);
    layer4_outputs(5183) <= not(layer3_outputs(2087)) or (layer3_outputs(3828));
    layer4_outputs(5184) <= layer3_outputs(10099);
    layer4_outputs(5185) <= layer3_outputs(5177);
    layer4_outputs(5186) <= layer3_outputs(9174);
    layer4_outputs(5187) <= (layer3_outputs(5211)) and not (layer3_outputs(9007));
    layer4_outputs(5188) <= not((layer3_outputs(9920)) xor (layer3_outputs(9339)));
    layer4_outputs(5189) <= (layer3_outputs(7205)) or (layer3_outputs(7254));
    layer4_outputs(5190) <= layer3_outputs(6097);
    layer4_outputs(5191) <= not((layer3_outputs(3373)) and (layer3_outputs(9998)));
    layer4_outputs(5192) <= not(layer3_outputs(1300));
    layer4_outputs(5193) <= layer3_outputs(1277);
    layer4_outputs(5194) <= (layer3_outputs(9480)) and not (layer3_outputs(9577));
    layer4_outputs(5195) <= not(layer3_outputs(4186)) or (layer3_outputs(9759));
    layer4_outputs(5196) <= layer3_outputs(6398);
    layer4_outputs(5197) <= not(layer3_outputs(834));
    layer4_outputs(5198) <= not(layer3_outputs(1597));
    layer4_outputs(5199) <= layer3_outputs(6255);
    layer4_outputs(5200) <= (layer3_outputs(9607)) xor (layer3_outputs(749));
    layer4_outputs(5201) <= layer3_outputs(8028);
    layer4_outputs(5202) <= not(layer3_outputs(9830)) or (layer3_outputs(7246));
    layer4_outputs(5203) <= layer3_outputs(8083);
    layer4_outputs(5204) <= (layer3_outputs(4102)) xor (layer3_outputs(6140));
    layer4_outputs(5205) <= (layer3_outputs(1497)) xor (layer3_outputs(9371));
    layer4_outputs(5206) <= layer3_outputs(6145);
    layer4_outputs(5207) <= not(layer3_outputs(1771));
    layer4_outputs(5208) <= not(layer3_outputs(9833)) or (layer3_outputs(8386));
    layer4_outputs(5209) <= layer3_outputs(3561);
    layer4_outputs(5210) <= not(layer3_outputs(8951));
    layer4_outputs(5211) <= not(layer3_outputs(8341));
    layer4_outputs(5212) <= not(layer3_outputs(8849));
    layer4_outputs(5213) <= layer3_outputs(8039);
    layer4_outputs(5214) <= not(layer3_outputs(2071));
    layer4_outputs(5215) <= not(layer3_outputs(8240));
    layer4_outputs(5216) <= layer3_outputs(4814);
    layer4_outputs(5217) <= layer3_outputs(7545);
    layer4_outputs(5218) <= not(layer3_outputs(3023));
    layer4_outputs(5219) <= layer3_outputs(8769);
    layer4_outputs(5220) <= not(layer3_outputs(1760));
    layer4_outputs(5221) <= (layer3_outputs(7411)) xor (layer3_outputs(6949));
    layer4_outputs(5222) <= not(layer3_outputs(8463)) or (layer3_outputs(3599));
    layer4_outputs(5223) <= not(layer3_outputs(3425)) or (layer3_outputs(5846));
    layer4_outputs(5224) <= not(layer3_outputs(7679)) or (layer3_outputs(1432));
    layer4_outputs(5225) <= not((layer3_outputs(6818)) and (layer3_outputs(8494)));
    layer4_outputs(5226) <= layer3_outputs(2107);
    layer4_outputs(5227) <= layer3_outputs(6408);
    layer4_outputs(5228) <= not(layer3_outputs(7932));
    layer4_outputs(5229) <= not(layer3_outputs(93));
    layer4_outputs(5230) <= layer3_outputs(8179);
    layer4_outputs(5231) <= (layer3_outputs(7101)) and (layer3_outputs(8011));
    layer4_outputs(5232) <= not(layer3_outputs(5789)) or (layer3_outputs(9646));
    layer4_outputs(5233) <= (layer3_outputs(903)) xor (layer3_outputs(5526));
    layer4_outputs(5234) <= layer3_outputs(10169);
    layer4_outputs(5235) <= not(layer3_outputs(6300));
    layer4_outputs(5236) <= not(layer3_outputs(4226));
    layer4_outputs(5237) <= not(layer3_outputs(3520));
    layer4_outputs(5238) <= layer3_outputs(2227);
    layer4_outputs(5239) <= not((layer3_outputs(7745)) and (layer3_outputs(5630)));
    layer4_outputs(5240) <= not(layer3_outputs(76));
    layer4_outputs(5241) <= (layer3_outputs(4409)) xor (layer3_outputs(8043));
    layer4_outputs(5242) <= layer3_outputs(2003);
    layer4_outputs(5243) <= layer3_outputs(5266);
    layer4_outputs(5244) <= not((layer3_outputs(7823)) xor (layer3_outputs(8909)));
    layer4_outputs(5245) <= not(layer3_outputs(7332));
    layer4_outputs(5246) <= not(layer3_outputs(9645));
    layer4_outputs(5247) <= layer3_outputs(118);
    layer4_outputs(5248) <= layer3_outputs(1211);
    layer4_outputs(5249) <= not(layer3_outputs(6656));
    layer4_outputs(5250) <= (layer3_outputs(9745)) and not (layer3_outputs(7465));
    layer4_outputs(5251) <= (layer3_outputs(6317)) and (layer3_outputs(7896));
    layer4_outputs(5252) <= not(layer3_outputs(1761));
    layer4_outputs(5253) <= (layer3_outputs(5517)) and not (layer3_outputs(4315));
    layer4_outputs(5254) <= (layer3_outputs(6999)) and (layer3_outputs(9999));
    layer4_outputs(5255) <= not(layer3_outputs(5907));
    layer4_outputs(5256) <= not(layer3_outputs(5820)) or (layer3_outputs(6456));
    layer4_outputs(5257) <= not(layer3_outputs(6242));
    layer4_outputs(5258) <= (layer3_outputs(4531)) xor (layer3_outputs(9388));
    layer4_outputs(5259) <= not((layer3_outputs(6332)) xor (layer3_outputs(1488)));
    layer4_outputs(5260) <= layer3_outputs(9518);
    layer4_outputs(5261) <= layer3_outputs(8323);
    layer4_outputs(5262) <= not(layer3_outputs(1127));
    layer4_outputs(5263) <= (layer3_outputs(9878)) and not (layer3_outputs(384));
    layer4_outputs(5264) <= layer3_outputs(1431);
    layer4_outputs(5265) <= not((layer3_outputs(5095)) and (layer3_outputs(4219)));
    layer4_outputs(5266) <= not(layer3_outputs(8015));
    layer4_outputs(5267) <= '1';
    layer4_outputs(5268) <= layer3_outputs(862);
    layer4_outputs(5269) <= not((layer3_outputs(6088)) xor (layer3_outputs(2491)));
    layer4_outputs(5270) <= not(layer3_outputs(3188));
    layer4_outputs(5271) <= not(layer3_outputs(7181));
    layer4_outputs(5272) <= not(layer3_outputs(6881));
    layer4_outputs(5273) <= not(layer3_outputs(4112));
    layer4_outputs(5274) <= not(layer3_outputs(9359));
    layer4_outputs(5275) <= not(layer3_outputs(1618));
    layer4_outputs(5276) <= not(layer3_outputs(2061));
    layer4_outputs(5277) <= (layer3_outputs(9290)) xor (layer3_outputs(614));
    layer4_outputs(5278) <= (layer3_outputs(3863)) xor (layer3_outputs(3390));
    layer4_outputs(5279) <= not((layer3_outputs(9864)) or (layer3_outputs(2275)));
    layer4_outputs(5280) <= not(layer3_outputs(4686));
    layer4_outputs(5281) <= not(layer3_outputs(7066)) or (layer3_outputs(5616));
    layer4_outputs(5282) <= (layer3_outputs(5182)) and not (layer3_outputs(4394));
    layer4_outputs(5283) <= not(layer3_outputs(7820));
    layer4_outputs(5284) <= not((layer3_outputs(4756)) xor (layer3_outputs(7730)));
    layer4_outputs(5285) <= not(layer3_outputs(9676));
    layer4_outputs(5286) <= (layer3_outputs(4757)) xor (layer3_outputs(2153));
    layer4_outputs(5287) <= layer3_outputs(7043);
    layer4_outputs(5288) <= (layer3_outputs(3998)) or (layer3_outputs(6784));
    layer4_outputs(5289) <= layer3_outputs(6599);
    layer4_outputs(5290) <= not((layer3_outputs(6534)) or (layer3_outputs(6194)));
    layer4_outputs(5291) <= not(layer3_outputs(4217)) or (layer3_outputs(6900));
    layer4_outputs(5292) <= not(layer3_outputs(3353));
    layer4_outputs(5293) <= layer3_outputs(2173);
    layer4_outputs(5294) <= (layer3_outputs(4434)) or (layer3_outputs(2692));
    layer4_outputs(5295) <= (layer3_outputs(9972)) xor (layer3_outputs(8119));
    layer4_outputs(5296) <= not(layer3_outputs(7838));
    layer4_outputs(5297) <= layer3_outputs(10200);
    layer4_outputs(5298) <= not(layer3_outputs(5520));
    layer4_outputs(5299) <= not(layer3_outputs(4935)) or (layer3_outputs(830));
    layer4_outputs(5300) <= (layer3_outputs(6204)) and (layer3_outputs(6382));
    layer4_outputs(5301) <= not(layer3_outputs(3354));
    layer4_outputs(5302) <= not(layer3_outputs(9725));
    layer4_outputs(5303) <= (layer3_outputs(3718)) and (layer3_outputs(2411));
    layer4_outputs(5304) <= not(layer3_outputs(2965));
    layer4_outputs(5305) <= not((layer3_outputs(958)) or (layer3_outputs(9523)));
    layer4_outputs(5306) <= layer3_outputs(8);
    layer4_outputs(5307) <= (layer3_outputs(9664)) xor (layer3_outputs(8344));
    layer4_outputs(5308) <= not(layer3_outputs(3291));
    layer4_outputs(5309) <= not(layer3_outputs(4378));
    layer4_outputs(5310) <= not(layer3_outputs(4698));
    layer4_outputs(5311) <= layer3_outputs(8732);
    layer4_outputs(5312) <= layer3_outputs(1561);
    layer4_outputs(5313) <= not((layer3_outputs(2879)) or (layer3_outputs(4444)));
    layer4_outputs(5314) <= layer3_outputs(2130);
    layer4_outputs(5315) <= layer3_outputs(4767);
    layer4_outputs(5316) <= not(layer3_outputs(5917));
    layer4_outputs(5317) <= layer3_outputs(7686);
    layer4_outputs(5318) <= layer3_outputs(5034);
    layer4_outputs(5319) <= (layer3_outputs(2453)) and not (layer3_outputs(1071));
    layer4_outputs(5320) <= layer3_outputs(72);
    layer4_outputs(5321) <= layer3_outputs(9019);
    layer4_outputs(5322) <= not(layer3_outputs(7666)) or (layer3_outputs(6548));
    layer4_outputs(5323) <= layer3_outputs(6024);
    layer4_outputs(5324) <= (layer3_outputs(8081)) and not (layer3_outputs(5935));
    layer4_outputs(5325) <= not(layer3_outputs(7324));
    layer4_outputs(5326) <= not(layer3_outputs(6115));
    layer4_outputs(5327) <= layer3_outputs(6692);
    layer4_outputs(5328) <= not(layer3_outputs(659));
    layer4_outputs(5329) <= not((layer3_outputs(10139)) or (layer3_outputs(6229)));
    layer4_outputs(5330) <= not(layer3_outputs(9442));
    layer4_outputs(5331) <= layer3_outputs(5755);
    layer4_outputs(5332) <= not(layer3_outputs(7974));
    layer4_outputs(5333) <= layer3_outputs(1813);
    layer4_outputs(5334) <= layer3_outputs(6085);
    layer4_outputs(5335) <= not(layer3_outputs(4411));
    layer4_outputs(5336) <= not((layer3_outputs(8075)) xor (layer3_outputs(10162)));
    layer4_outputs(5337) <= layer3_outputs(2406);
    layer4_outputs(5338) <= not(layer3_outputs(5141));
    layer4_outputs(5339) <= not(layer3_outputs(8159));
    layer4_outputs(5340) <= not(layer3_outputs(9317));
    layer4_outputs(5341) <= layer3_outputs(3104);
    layer4_outputs(5342) <= layer3_outputs(1821);
    layer4_outputs(5343) <= (layer3_outputs(3711)) and not (layer3_outputs(275));
    layer4_outputs(5344) <= not(layer3_outputs(226));
    layer4_outputs(5345) <= (layer3_outputs(5095)) and not (layer3_outputs(2064));
    layer4_outputs(5346) <= layer3_outputs(4362);
    layer4_outputs(5347) <= not(layer3_outputs(7681));
    layer4_outputs(5348) <= not((layer3_outputs(2680)) xor (layer3_outputs(4674)));
    layer4_outputs(5349) <= not(layer3_outputs(1316));
    layer4_outputs(5350) <= (layer3_outputs(9029)) xor (layer3_outputs(4829));
    layer4_outputs(5351) <= not(layer3_outputs(6474));
    layer4_outputs(5352) <= layer3_outputs(6733);
    layer4_outputs(5353) <= not((layer3_outputs(3588)) xor (layer3_outputs(10159)));
    layer4_outputs(5354) <= layer3_outputs(9597);
    layer4_outputs(5355) <= not(layer3_outputs(1256));
    layer4_outputs(5356) <= (layer3_outputs(7861)) and (layer3_outputs(9967));
    layer4_outputs(5357) <= (layer3_outputs(5580)) and not (layer3_outputs(4847));
    layer4_outputs(5358) <= layer3_outputs(9367);
    layer4_outputs(5359) <= layer3_outputs(3415);
    layer4_outputs(5360) <= not(layer3_outputs(7563)) or (layer3_outputs(4108));
    layer4_outputs(5361) <= layer3_outputs(9376);
    layer4_outputs(5362) <= layer3_outputs(8762);
    layer4_outputs(5363) <= not(layer3_outputs(4918));
    layer4_outputs(5364) <= layer3_outputs(6500);
    layer4_outputs(5365) <= (layer3_outputs(4931)) or (layer3_outputs(7461));
    layer4_outputs(5366) <= not((layer3_outputs(5504)) and (layer3_outputs(9993)));
    layer4_outputs(5367) <= layer3_outputs(361);
    layer4_outputs(5368) <= layer3_outputs(1340);
    layer4_outputs(5369) <= layer3_outputs(872);
    layer4_outputs(5370) <= not(layer3_outputs(8146));
    layer4_outputs(5371) <= not(layer3_outputs(2745));
    layer4_outputs(5372) <= not(layer3_outputs(1582)) or (layer3_outputs(5324));
    layer4_outputs(5373) <= (layer3_outputs(7744)) and not (layer3_outputs(6926));
    layer4_outputs(5374) <= layer3_outputs(1217);
    layer4_outputs(5375) <= not((layer3_outputs(10015)) xor (layer3_outputs(8103)));
    layer4_outputs(5376) <= layer3_outputs(3754);
    layer4_outputs(5377) <= (layer3_outputs(3334)) and not (layer3_outputs(2497));
    layer4_outputs(5378) <= layer3_outputs(4142);
    layer4_outputs(5379) <= not((layer3_outputs(3196)) or (layer3_outputs(7332)));
    layer4_outputs(5380) <= not(layer3_outputs(6487)) or (layer3_outputs(9753));
    layer4_outputs(5381) <= layer3_outputs(1626);
    layer4_outputs(5382) <= not(layer3_outputs(8750));
    layer4_outputs(5383) <= (layer3_outputs(1124)) xor (layer3_outputs(7624));
    layer4_outputs(5384) <= not((layer3_outputs(6247)) and (layer3_outputs(2136)));
    layer4_outputs(5385) <= not((layer3_outputs(3882)) and (layer3_outputs(5971)));
    layer4_outputs(5386) <= not(layer3_outputs(5915));
    layer4_outputs(5387) <= not((layer3_outputs(6987)) xor (layer3_outputs(3587)));
    layer4_outputs(5388) <= not((layer3_outputs(509)) or (layer3_outputs(7742)));
    layer4_outputs(5389) <= (layer3_outputs(7071)) or (layer3_outputs(9747));
    layer4_outputs(5390) <= (layer3_outputs(2921)) xor (layer3_outputs(3989));
    layer4_outputs(5391) <= not((layer3_outputs(1326)) or (layer3_outputs(8574)));
    layer4_outputs(5392) <= (layer3_outputs(1370)) or (layer3_outputs(10035));
    layer4_outputs(5393) <= layer3_outputs(1385);
    layer4_outputs(5394) <= not(layer3_outputs(8847)) or (layer3_outputs(5561));
    layer4_outputs(5395) <= not(layer3_outputs(6660)) or (layer3_outputs(8703));
    layer4_outputs(5396) <= not((layer3_outputs(4968)) xor (layer3_outputs(9215)));
    layer4_outputs(5397) <= (layer3_outputs(469)) and not (layer3_outputs(9379));
    layer4_outputs(5398) <= not(layer3_outputs(1207));
    layer4_outputs(5399) <= (layer3_outputs(4814)) and not (layer3_outputs(2149));
    layer4_outputs(5400) <= (layer3_outputs(2373)) and (layer3_outputs(4311));
    layer4_outputs(5401) <= not(layer3_outputs(3197));
    layer4_outputs(5402) <= layer3_outputs(5447);
    layer4_outputs(5403) <= not(layer3_outputs(5667));
    layer4_outputs(5404) <= layer3_outputs(7044);
    layer4_outputs(5405) <= not(layer3_outputs(1436));
    layer4_outputs(5406) <= not(layer3_outputs(2653)) or (layer3_outputs(3797));
    layer4_outputs(5407) <= (layer3_outputs(1216)) or (layer3_outputs(7819));
    layer4_outputs(5408) <= not(layer3_outputs(67));
    layer4_outputs(5409) <= not(layer3_outputs(8190));
    layer4_outputs(5410) <= not(layer3_outputs(469));
    layer4_outputs(5411) <= not(layer3_outputs(922));
    layer4_outputs(5412) <= not(layer3_outputs(1409)) or (layer3_outputs(4580));
    layer4_outputs(5413) <= not(layer3_outputs(3352));
    layer4_outputs(5414) <= not((layer3_outputs(329)) or (layer3_outputs(2008)));
    layer4_outputs(5415) <= layer3_outputs(7364);
    layer4_outputs(5416) <= not(layer3_outputs(9567)) or (layer3_outputs(4227));
    layer4_outputs(5417) <= not(layer3_outputs(2545));
    layer4_outputs(5418) <= not((layer3_outputs(1247)) xor (layer3_outputs(7445)));
    layer4_outputs(5419) <= layer3_outputs(1768);
    layer4_outputs(5420) <= not(layer3_outputs(2766));
    layer4_outputs(5421) <= not((layer3_outputs(480)) and (layer3_outputs(9368)));
    layer4_outputs(5422) <= layer3_outputs(4241);
    layer4_outputs(5423) <= (layer3_outputs(2162)) and not (layer3_outputs(2417));
    layer4_outputs(5424) <= not(layer3_outputs(8297));
    layer4_outputs(5425) <= not((layer3_outputs(8318)) xor (layer3_outputs(5538)));
    layer4_outputs(5426) <= (layer3_outputs(2382)) and not (layer3_outputs(1042));
    layer4_outputs(5427) <= not(layer3_outputs(3991));
    layer4_outputs(5428) <= (layer3_outputs(2935)) or (layer3_outputs(4580));
    layer4_outputs(5429) <= layer3_outputs(9962);
    layer4_outputs(5430) <= not(layer3_outputs(32));
    layer4_outputs(5431) <= not(layer3_outputs(3950)) or (layer3_outputs(2546));
    layer4_outputs(5432) <= layer3_outputs(661);
    layer4_outputs(5433) <= (layer3_outputs(8073)) xor (layer3_outputs(7372));
    layer4_outputs(5434) <= layer3_outputs(8653);
    layer4_outputs(5435) <= layer3_outputs(511);
    layer4_outputs(5436) <= not((layer3_outputs(281)) or (layer3_outputs(2357)));
    layer4_outputs(5437) <= layer3_outputs(2633);
    layer4_outputs(5438) <= layer3_outputs(1389);
    layer4_outputs(5439) <= layer3_outputs(8647);
    layer4_outputs(5440) <= (layer3_outputs(2018)) or (layer3_outputs(7230));
    layer4_outputs(5441) <= (layer3_outputs(4603)) and not (layer3_outputs(4484));
    layer4_outputs(5442) <= not(layer3_outputs(5283));
    layer4_outputs(5443) <= (layer3_outputs(428)) xor (layer3_outputs(3191));
    layer4_outputs(5444) <= not((layer3_outputs(322)) and (layer3_outputs(8863)));
    layer4_outputs(5445) <= not(layer3_outputs(2724));
    layer4_outputs(5446) <= (layer3_outputs(9566)) xor (layer3_outputs(750));
    layer4_outputs(5447) <= (layer3_outputs(4620)) and not (layer3_outputs(3111));
    layer4_outputs(5448) <= (layer3_outputs(6068)) and (layer3_outputs(2305));
    layer4_outputs(5449) <= (layer3_outputs(5954)) and (layer3_outputs(2500));
    layer4_outputs(5450) <= not(layer3_outputs(9405));
    layer4_outputs(5451) <= not((layer3_outputs(9884)) xor (layer3_outputs(6343)));
    layer4_outputs(5452) <= not((layer3_outputs(6278)) and (layer3_outputs(5980)));
    layer4_outputs(5453) <= layer3_outputs(3543);
    layer4_outputs(5454) <= not((layer3_outputs(5361)) and (layer3_outputs(4230)));
    layer4_outputs(5455) <= not(layer3_outputs(9611)) or (layer3_outputs(1253));
    layer4_outputs(5456) <= not(layer3_outputs(1444));
    layer4_outputs(5457) <= layer3_outputs(388);
    layer4_outputs(5458) <= not(layer3_outputs(1291));
    layer4_outputs(5459) <= layer3_outputs(698);
    layer4_outputs(5460) <= not(layer3_outputs(2366));
    layer4_outputs(5461) <= not(layer3_outputs(3836));
    layer4_outputs(5462) <= (layer3_outputs(5980)) or (layer3_outputs(9229));
    layer4_outputs(5463) <= layer3_outputs(10093);
    layer4_outputs(5464) <= layer3_outputs(3878);
    layer4_outputs(5465) <= not((layer3_outputs(7890)) xor (layer3_outputs(7467)));
    layer4_outputs(5466) <= not(layer3_outputs(1782)) or (layer3_outputs(1216));
    layer4_outputs(5467) <= layer3_outputs(9782);
    layer4_outputs(5468) <= (layer3_outputs(3503)) and (layer3_outputs(5254));
    layer4_outputs(5469) <= not(layer3_outputs(4275));
    layer4_outputs(5470) <= layer3_outputs(8906);
    layer4_outputs(5471) <= not((layer3_outputs(1373)) xor (layer3_outputs(1315)));
    layer4_outputs(5472) <= (layer3_outputs(2225)) or (layer3_outputs(781));
    layer4_outputs(5473) <= layer3_outputs(9666);
    layer4_outputs(5474) <= not(layer3_outputs(4346));
    layer4_outputs(5475) <= not((layer3_outputs(3411)) xor (layer3_outputs(9106)));
    layer4_outputs(5476) <= (layer3_outputs(7615)) and not (layer3_outputs(9232));
    layer4_outputs(5477) <= layer3_outputs(1593);
    layer4_outputs(5478) <= (layer3_outputs(2280)) and not (layer3_outputs(3173));
    layer4_outputs(5479) <= (layer3_outputs(3658)) or (layer3_outputs(8434));
    layer4_outputs(5480) <= not(layer3_outputs(6412));
    layer4_outputs(5481) <= (layer3_outputs(6138)) xor (layer3_outputs(6079));
    layer4_outputs(5482) <= (layer3_outputs(51)) and not (layer3_outputs(3722));
    layer4_outputs(5483) <= not(layer3_outputs(9957));
    layer4_outputs(5484) <= not(layer3_outputs(1011));
    layer4_outputs(5485) <= layer3_outputs(1220);
    layer4_outputs(5486) <= not(layer3_outputs(8996));
    layer4_outputs(5487) <= layer3_outputs(6304);
    layer4_outputs(5488) <= layer3_outputs(8461);
    layer4_outputs(5489) <= not(layer3_outputs(4494));
    layer4_outputs(5490) <= not(layer3_outputs(7311));
    layer4_outputs(5491) <= not((layer3_outputs(1866)) or (layer3_outputs(6275)));
    layer4_outputs(5492) <= not(layer3_outputs(5298));
    layer4_outputs(5493) <= not((layer3_outputs(17)) xor (layer3_outputs(2039)));
    layer4_outputs(5494) <= not(layer3_outputs(2094));
    layer4_outputs(5495) <= not(layer3_outputs(190));
    layer4_outputs(5496) <= not(layer3_outputs(2783));
    layer4_outputs(5497) <= not((layer3_outputs(7767)) xor (layer3_outputs(372)));
    layer4_outputs(5498) <= not(layer3_outputs(1678));
    layer4_outputs(5499) <= layer3_outputs(393);
    layer4_outputs(5500) <= layer3_outputs(1134);
    layer4_outputs(5501) <= not(layer3_outputs(6429));
    layer4_outputs(5502) <= (layer3_outputs(1064)) and (layer3_outputs(3008));
    layer4_outputs(5503) <= not(layer3_outputs(1839));
    layer4_outputs(5504) <= not(layer3_outputs(8778));
    layer4_outputs(5505) <= (layer3_outputs(10108)) and not (layer3_outputs(1185));
    layer4_outputs(5506) <= not((layer3_outputs(525)) xor (layer3_outputs(6119)));
    layer4_outputs(5507) <= not(layer3_outputs(2885));
    layer4_outputs(5508) <= layer3_outputs(623);
    layer4_outputs(5509) <= (layer3_outputs(2395)) and (layer3_outputs(3781));
    layer4_outputs(5510) <= layer3_outputs(2062);
    layer4_outputs(5511) <= (layer3_outputs(9177)) and (layer3_outputs(4372));
    layer4_outputs(5512) <= (layer3_outputs(1026)) xor (layer3_outputs(2833));
    layer4_outputs(5513) <= not((layer3_outputs(1016)) xor (layer3_outputs(2276)));
    layer4_outputs(5514) <= layer3_outputs(6841);
    layer4_outputs(5515) <= layer3_outputs(983);
    layer4_outputs(5516) <= not(layer3_outputs(4213)) or (layer3_outputs(8711));
    layer4_outputs(5517) <= not((layer3_outputs(7022)) xor (layer3_outputs(2432)));
    layer4_outputs(5518) <= not(layer3_outputs(4087));
    layer4_outputs(5519) <= layer3_outputs(285);
    layer4_outputs(5520) <= layer3_outputs(827);
    layer4_outputs(5521) <= not(layer3_outputs(10030));
    layer4_outputs(5522) <= not(layer3_outputs(4489));
    layer4_outputs(5523) <= not(layer3_outputs(6970)) or (layer3_outputs(9584));
    layer4_outputs(5524) <= not(layer3_outputs(2462)) or (layer3_outputs(5220));
    layer4_outputs(5525) <= layer3_outputs(10179);
    layer4_outputs(5526) <= layer3_outputs(6621);
    layer4_outputs(5527) <= layer3_outputs(1483);
    layer4_outputs(5528) <= (layer3_outputs(7850)) and (layer3_outputs(2936));
    layer4_outputs(5529) <= (layer3_outputs(2800)) and (layer3_outputs(2353));
    layer4_outputs(5530) <= not(layer3_outputs(1003));
    layer4_outputs(5531) <= not(layer3_outputs(354));
    layer4_outputs(5532) <= not(layer3_outputs(4015));
    layer4_outputs(5533) <= not(layer3_outputs(8401)) or (layer3_outputs(2914));
    layer4_outputs(5534) <= layer3_outputs(3956);
    layer4_outputs(5535) <= not((layer3_outputs(9285)) and (layer3_outputs(5644)));
    layer4_outputs(5536) <= not(layer3_outputs(8742));
    layer4_outputs(5537) <= layer3_outputs(5810);
    layer4_outputs(5538) <= not(layer3_outputs(9981)) or (layer3_outputs(6773));
    layer4_outputs(5539) <= (layer3_outputs(563)) and not (layer3_outputs(2267));
    layer4_outputs(5540) <= not(layer3_outputs(1051));
    layer4_outputs(5541) <= layer3_outputs(4272);
    layer4_outputs(5542) <= not(layer3_outputs(5819)) or (layer3_outputs(8248));
    layer4_outputs(5543) <= layer3_outputs(4256);
    layer4_outputs(5544) <= not(layer3_outputs(145));
    layer4_outputs(5545) <= layer3_outputs(1972);
    layer4_outputs(5546) <= layer3_outputs(2380);
    layer4_outputs(5547) <= not(layer3_outputs(5196)) or (layer3_outputs(9109));
    layer4_outputs(5548) <= layer3_outputs(453);
    layer4_outputs(5549) <= not(layer3_outputs(1123));
    layer4_outputs(5550) <= not(layer3_outputs(6659)) or (layer3_outputs(5454));
    layer4_outputs(5551) <= layer3_outputs(8997);
    layer4_outputs(5552) <= not(layer3_outputs(9784)) or (layer3_outputs(2759));
    layer4_outputs(5553) <= not(layer3_outputs(1233));
    layer4_outputs(5554) <= (layer3_outputs(4884)) or (layer3_outputs(2813));
    layer4_outputs(5555) <= not(layer3_outputs(5645));
    layer4_outputs(5556) <= layer3_outputs(3358);
    layer4_outputs(5557) <= not((layer3_outputs(1)) xor (layer3_outputs(7391)));
    layer4_outputs(5558) <= (layer3_outputs(3901)) and (layer3_outputs(4625));
    layer4_outputs(5559) <= not((layer3_outputs(842)) xor (layer3_outputs(9354)));
    layer4_outputs(5560) <= layer3_outputs(9461);
    layer4_outputs(5561) <= (layer3_outputs(2249)) and not (layer3_outputs(2480));
    layer4_outputs(5562) <= not(layer3_outputs(8065));
    layer4_outputs(5563) <= layer3_outputs(5592);
    layer4_outputs(5564) <= layer3_outputs(268);
    layer4_outputs(5565) <= layer3_outputs(9738);
    layer4_outputs(5566) <= not(layer3_outputs(1449));
    layer4_outputs(5567) <= layer3_outputs(3951);
    layer4_outputs(5568) <= not(layer3_outputs(9741));
    layer4_outputs(5569) <= not(layer3_outputs(6998));
    layer4_outputs(5570) <= not((layer3_outputs(8756)) xor (layer3_outputs(8962)));
    layer4_outputs(5571) <= layer3_outputs(8042);
    layer4_outputs(5572) <= layer3_outputs(6251);
    layer4_outputs(5573) <= (layer3_outputs(2031)) and (layer3_outputs(699));
    layer4_outputs(5574) <= layer3_outputs(4257);
    layer4_outputs(5575) <= layer3_outputs(3311);
    layer4_outputs(5576) <= not(layer3_outputs(7134));
    layer4_outputs(5577) <= layer3_outputs(3240);
    layer4_outputs(5578) <= not((layer3_outputs(8883)) and (layer3_outputs(6208)));
    layer4_outputs(5579) <= not((layer3_outputs(10233)) or (layer3_outputs(3236)));
    layer4_outputs(5580) <= not(layer3_outputs(3809));
    layer4_outputs(5581) <= not(layer3_outputs(10146));
    layer4_outputs(5582) <= layer3_outputs(7119);
    layer4_outputs(5583) <= layer3_outputs(7191);
    layer4_outputs(5584) <= (layer3_outputs(5365)) or (layer3_outputs(7305));
    layer4_outputs(5585) <= (layer3_outputs(3986)) or (layer3_outputs(5117));
    layer4_outputs(5586) <= (layer3_outputs(5632)) xor (layer3_outputs(7884));
    layer4_outputs(5587) <= (layer3_outputs(7728)) xor (layer3_outputs(293));
    layer4_outputs(5588) <= (layer3_outputs(3089)) xor (layer3_outputs(3613));
    layer4_outputs(5589) <= not((layer3_outputs(1440)) and (layer3_outputs(2001)));
    layer4_outputs(5590) <= not((layer3_outputs(3607)) and (layer3_outputs(3727)));
    layer4_outputs(5591) <= not(layer3_outputs(2858)) or (layer3_outputs(5223));
    layer4_outputs(5592) <= (layer3_outputs(1800)) and (layer3_outputs(1908));
    layer4_outputs(5593) <= layer3_outputs(8930);
    layer4_outputs(5594) <= not(layer3_outputs(5497));
    layer4_outputs(5595) <= layer3_outputs(1439);
    layer4_outputs(5596) <= (layer3_outputs(2588)) or (layer3_outputs(9624));
    layer4_outputs(5597) <= not(layer3_outputs(9895));
    layer4_outputs(5598) <= layer3_outputs(7327);
    layer4_outputs(5599) <= (layer3_outputs(10061)) and not (layer3_outputs(6502));
    layer4_outputs(5600) <= not((layer3_outputs(8154)) and (layer3_outputs(8949)));
    layer4_outputs(5601) <= not((layer3_outputs(520)) xor (layer3_outputs(2616)));
    layer4_outputs(5602) <= '0';
    layer4_outputs(5603) <= layer3_outputs(4979);
    layer4_outputs(5604) <= (layer3_outputs(1430)) and (layer3_outputs(339));
    layer4_outputs(5605) <= not((layer3_outputs(10100)) xor (layer3_outputs(9009)));
    layer4_outputs(5606) <= layer3_outputs(9407);
    layer4_outputs(5607) <= not(layer3_outputs(8349));
    layer4_outputs(5608) <= not(layer3_outputs(7487));
    layer4_outputs(5609) <= not(layer3_outputs(9445));
    layer4_outputs(5610) <= (layer3_outputs(3888)) and not (layer3_outputs(1182));
    layer4_outputs(5611) <= (layer3_outputs(9759)) and (layer3_outputs(10210));
    layer4_outputs(5612) <= not(layer3_outputs(3985));
    layer4_outputs(5613) <= not(layer3_outputs(745));
    layer4_outputs(5614) <= not(layer3_outputs(4112));
    layer4_outputs(5615) <= layer3_outputs(2142);
    layer4_outputs(5616) <= not(layer3_outputs(1604)) or (layer3_outputs(4669));
    layer4_outputs(5617) <= not((layer3_outputs(2145)) and (layer3_outputs(7842)));
    layer4_outputs(5618) <= (layer3_outputs(7774)) xor (layer3_outputs(9381));
    layer4_outputs(5619) <= not((layer3_outputs(10059)) or (layer3_outputs(9494)));
    layer4_outputs(5620) <= layer3_outputs(1201);
    layer4_outputs(5621) <= (layer3_outputs(2004)) or (layer3_outputs(9483));
    layer4_outputs(5622) <= (layer3_outputs(7514)) or (layer3_outputs(3476));
    layer4_outputs(5623) <= '0';
    layer4_outputs(5624) <= layer3_outputs(528);
    layer4_outputs(5625) <= (layer3_outputs(4745)) and not (layer3_outputs(6854));
    layer4_outputs(5626) <= not(layer3_outputs(2874));
    layer4_outputs(5627) <= not(layer3_outputs(3123));
    layer4_outputs(5628) <= (layer3_outputs(6341)) and not (layer3_outputs(562));
    layer4_outputs(5629) <= (layer3_outputs(8255)) and (layer3_outputs(3632));
    layer4_outputs(5630) <= (layer3_outputs(2797)) and (layer3_outputs(7175));
    layer4_outputs(5631) <= (layer3_outputs(2910)) and not (layer3_outputs(7540));
    layer4_outputs(5632) <= layer3_outputs(7724);
    layer4_outputs(5633) <= '0';
    layer4_outputs(5634) <= not(layer3_outputs(3452));
    layer4_outputs(5635) <= layer3_outputs(9934);
    layer4_outputs(5636) <= not(layer3_outputs(4035));
    layer4_outputs(5637) <= (layer3_outputs(10237)) xor (layer3_outputs(9856));
    layer4_outputs(5638) <= (layer3_outputs(7378)) and (layer3_outputs(10095));
    layer4_outputs(5639) <= layer3_outputs(789);
    layer4_outputs(5640) <= not(layer3_outputs(4834));
    layer4_outputs(5641) <= (layer3_outputs(8403)) and (layer3_outputs(4734));
    layer4_outputs(5642) <= layer3_outputs(5059);
    layer4_outputs(5643) <= not(layer3_outputs(7707));
    layer4_outputs(5644) <= not(layer3_outputs(5428));
    layer4_outputs(5645) <= layer3_outputs(7873);
    layer4_outputs(5646) <= not(layer3_outputs(5132));
    layer4_outputs(5647) <= (layer3_outputs(2677)) and not (layer3_outputs(4660));
    layer4_outputs(5648) <= layer3_outputs(2441);
    layer4_outputs(5649) <= layer3_outputs(10160);
    layer4_outputs(5650) <= not(layer3_outputs(5967));
    layer4_outputs(5651) <= not(layer3_outputs(3840)) or (layer3_outputs(9409));
    layer4_outputs(5652) <= not(layer3_outputs(8668));
    layer4_outputs(5653) <= not(layer3_outputs(2286));
    layer4_outputs(5654) <= (layer3_outputs(8044)) or (layer3_outputs(6778));
    layer4_outputs(5655) <= not(layer3_outputs(6997));
    layer4_outputs(5656) <= (layer3_outputs(6382)) and not (layer3_outputs(1603));
    layer4_outputs(5657) <= not(layer3_outputs(6667)) or (layer3_outputs(7120));
    layer4_outputs(5658) <= not(layer3_outputs(7287));
    layer4_outputs(5659) <= not(layer3_outputs(6464));
    layer4_outputs(5660) <= not(layer3_outputs(5843));
    layer4_outputs(5661) <= not(layer3_outputs(9873)) or (layer3_outputs(1149));
    layer4_outputs(5662) <= (layer3_outputs(33)) and (layer3_outputs(8394));
    layer4_outputs(5663) <= not(layer3_outputs(2710));
    layer4_outputs(5664) <= not(layer3_outputs(6237));
    layer4_outputs(5665) <= not((layer3_outputs(9248)) xor (layer3_outputs(6213)));
    layer4_outputs(5666) <= not((layer3_outputs(6425)) xor (layer3_outputs(2390)));
    layer4_outputs(5667) <= not(layer3_outputs(9547));
    layer4_outputs(5668) <= not((layer3_outputs(2906)) xor (layer3_outputs(2181)));
    layer4_outputs(5669) <= not(layer3_outputs(7143));
    layer4_outputs(5670) <= layer3_outputs(1782);
    layer4_outputs(5671) <= '1';
    layer4_outputs(5672) <= (layer3_outputs(9280)) xor (layer3_outputs(4629));
    layer4_outputs(5673) <= not(layer3_outputs(7440));
    layer4_outputs(5674) <= layer3_outputs(7827);
    layer4_outputs(5675) <= not(layer3_outputs(9152)) or (layer3_outputs(1064));
    layer4_outputs(5676) <= (layer3_outputs(4935)) and (layer3_outputs(1413));
    layer4_outputs(5677) <= not((layer3_outputs(6648)) and (layer3_outputs(1888)));
    layer4_outputs(5678) <= (layer3_outputs(9670)) and not (layer3_outputs(6906));
    layer4_outputs(5679) <= (layer3_outputs(390)) xor (layer3_outputs(483));
    layer4_outputs(5680) <= (layer3_outputs(3318)) and not (layer3_outputs(3068));
    layer4_outputs(5681) <= (layer3_outputs(451)) or (layer3_outputs(2615));
    layer4_outputs(5682) <= layer3_outputs(9722);
    layer4_outputs(5683) <= not(layer3_outputs(9511)) or (layer3_outputs(8952));
    layer4_outputs(5684) <= layer3_outputs(5765);
    layer4_outputs(5685) <= not(layer3_outputs(7188));
    layer4_outputs(5686) <= not((layer3_outputs(3078)) xor (layer3_outputs(7798)));
    layer4_outputs(5687) <= not(layer3_outputs(6960));
    layer4_outputs(5688) <= (layer3_outputs(8282)) and (layer3_outputs(2215));
    layer4_outputs(5689) <= not(layer3_outputs(839));
    layer4_outputs(5690) <= layer3_outputs(7982);
    layer4_outputs(5691) <= not((layer3_outputs(9561)) or (layer3_outputs(1862)));
    layer4_outputs(5692) <= not(layer3_outputs(7692));
    layer4_outputs(5693) <= not(layer3_outputs(7616));
    layer4_outputs(5694) <= not(layer3_outputs(3420));
    layer4_outputs(5695) <= (layer3_outputs(7726)) and (layer3_outputs(8648));
    layer4_outputs(5696) <= not(layer3_outputs(2262));
    layer4_outputs(5697) <= layer3_outputs(7737);
    layer4_outputs(5698) <= layer3_outputs(3336);
    layer4_outputs(5699) <= not((layer3_outputs(0)) or (layer3_outputs(1883)));
    layer4_outputs(5700) <= layer3_outputs(10219);
    layer4_outputs(5701) <= layer3_outputs(301);
    layer4_outputs(5702) <= layer3_outputs(6097);
    layer4_outputs(5703) <= (layer3_outputs(8340)) and not (layer3_outputs(8816));
    layer4_outputs(5704) <= not((layer3_outputs(6725)) or (layer3_outputs(655)));
    layer4_outputs(5705) <= not(layer3_outputs(108)) or (layer3_outputs(5206));
    layer4_outputs(5706) <= layer3_outputs(5172);
    layer4_outputs(5707) <= not(layer3_outputs(2172));
    layer4_outputs(5708) <= (layer3_outputs(7369)) and (layer3_outputs(2006));
    layer4_outputs(5709) <= not(layer3_outputs(2470));
    layer4_outputs(5710) <= layer3_outputs(4636);
    layer4_outputs(5711) <= not(layer3_outputs(6835));
    layer4_outputs(5712) <= not(layer3_outputs(6358));
    layer4_outputs(5713) <= not(layer3_outputs(3155)) or (layer3_outputs(1074));
    layer4_outputs(5714) <= layer3_outputs(3865);
    layer4_outputs(5715) <= layer3_outputs(6950);
    layer4_outputs(5716) <= not(layer3_outputs(2140)) or (layer3_outputs(7556));
    layer4_outputs(5717) <= layer3_outputs(85);
    layer4_outputs(5718) <= layer3_outputs(9279);
    layer4_outputs(5719) <= (layer3_outputs(1424)) and not (layer3_outputs(6943));
    layer4_outputs(5720) <= (layer3_outputs(7986)) xor (layer3_outputs(5269));
    layer4_outputs(5721) <= (layer3_outputs(9480)) and not (layer3_outputs(4847));
    layer4_outputs(5722) <= (layer3_outputs(6047)) and not (layer3_outputs(6666));
    layer4_outputs(5723) <= layer3_outputs(8426);
    layer4_outputs(5724) <= layer3_outputs(1572);
    layer4_outputs(5725) <= not(layer3_outputs(5258));
    layer4_outputs(5726) <= not((layer3_outputs(4179)) or (layer3_outputs(8818)));
    layer4_outputs(5727) <= (layer3_outputs(4090)) xor (layer3_outputs(815));
    layer4_outputs(5728) <= not(layer3_outputs(3079));
    layer4_outputs(5729) <= (layer3_outputs(7535)) or (layer3_outputs(9012));
    layer4_outputs(5730) <= not(layer3_outputs(4249));
    layer4_outputs(5731) <= not(layer3_outputs(7333));
    layer4_outputs(5732) <= layer3_outputs(3605);
    layer4_outputs(5733) <= not(layer3_outputs(897)) or (layer3_outputs(5455));
    layer4_outputs(5734) <= not(layer3_outputs(6131));
    layer4_outputs(5735) <= (layer3_outputs(7909)) xor (layer3_outputs(6615));
    layer4_outputs(5736) <= layer3_outputs(4915);
    layer4_outputs(5737) <= not(layer3_outputs(4130));
    layer4_outputs(5738) <= (layer3_outputs(10176)) or (layer3_outputs(4528));
    layer4_outputs(5739) <= layer3_outputs(7111);
    layer4_outputs(5740) <= layer3_outputs(2321);
    layer4_outputs(5741) <= not((layer3_outputs(675)) or (layer3_outputs(8400)));
    layer4_outputs(5742) <= (layer3_outputs(3873)) and not (layer3_outputs(1869));
    layer4_outputs(5743) <= not(layer3_outputs(132));
    layer4_outputs(5744) <= not(layer3_outputs(1465)) or (layer3_outputs(2311));
    layer4_outputs(5745) <= layer3_outputs(6369);
    layer4_outputs(5746) <= layer3_outputs(478);
    layer4_outputs(5747) <= '0';
    layer4_outputs(5748) <= not(layer3_outputs(1638));
    layer4_outputs(5749) <= not(layer3_outputs(8617));
    layer4_outputs(5750) <= not(layer3_outputs(8444));
    layer4_outputs(5751) <= layer3_outputs(7635);
    layer4_outputs(5752) <= not(layer3_outputs(1276));
    layer4_outputs(5753) <= layer3_outputs(6573);
    layer4_outputs(5754) <= not(layer3_outputs(1896));
    layer4_outputs(5755) <= not(layer3_outputs(492));
    layer4_outputs(5756) <= layer3_outputs(9429);
    layer4_outputs(5757) <= not(layer3_outputs(8964)) or (layer3_outputs(7213));
    layer4_outputs(5758) <= not((layer3_outputs(4312)) xor (layer3_outputs(6562)));
    layer4_outputs(5759) <= not(layer3_outputs(2017));
    layer4_outputs(5760) <= not(layer3_outputs(5652));
    layer4_outputs(5761) <= not(layer3_outputs(6837));
    layer4_outputs(5762) <= not(layer3_outputs(7590));
    layer4_outputs(5763) <= not(layer3_outputs(4588));
    layer4_outputs(5764) <= not(layer3_outputs(804));
    layer4_outputs(5765) <= (layer3_outputs(5941)) and not (layer3_outputs(9157));
    layer4_outputs(5766) <= (layer3_outputs(2482)) xor (layer3_outputs(2907));
    layer4_outputs(5767) <= not((layer3_outputs(4132)) or (layer3_outputs(3553)));
    layer4_outputs(5768) <= not((layer3_outputs(1402)) xor (layer3_outputs(9068)));
    layer4_outputs(5769) <= layer3_outputs(1054);
    layer4_outputs(5770) <= not(layer3_outputs(8490));
    layer4_outputs(5771) <= not((layer3_outputs(1570)) or (layer3_outputs(3967)));
    layer4_outputs(5772) <= not(layer3_outputs(7375));
    layer4_outputs(5773) <= not((layer3_outputs(3395)) xor (layer3_outputs(9697)));
    layer4_outputs(5774) <= not(layer3_outputs(2147)) or (layer3_outputs(2598));
    layer4_outputs(5775) <= not(layer3_outputs(6963));
    layer4_outputs(5776) <= (layer3_outputs(3766)) and not (layer3_outputs(9574));
    layer4_outputs(5777) <= not(layer3_outputs(9888)) or (layer3_outputs(3880));
    layer4_outputs(5778) <= layer3_outputs(9572);
    layer4_outputs(5779) <= layer3_outputs(8162);
    layer4_outputs(5780) <= not(layer3_outputs(4585));
    layer4_outputs(5781) <= not(layer3_outputs(7936));
    layer4_outputs(5782) <= not(layer3_outputs(719));
    layer4_outputs(5783) <= not(layer3_outputs(8895));
    layer4_outputs(5784) <= layer3_outputs(4342);
    layer4_outputs(5785) <= '0';
    layer4_outputs(5786) <= not((layer3_outputs(824)) xor (layer3_outputs(6367)));
    layer4_outputs(5787) <= layer3_outputs(1718);
    layer4_outputs(5788) <= not(layer3_outputs(4408));
    layer4_outputs(5789) <= not(layer3_outputs(3052));
    layer4_outputs(5790) <= not(layer3_outputs(638)) or (layer3_outputs(7833));
    layer4_outputs(5791) <= not(layer3_outputs(7836));
    layer4_outputs(5792) <= not(layer3_outputs(932));
    layer4_outputs(5793) <= not((layer3_outputs(1451)) xor (layer3_outputs(3118)));
    layer4_outputs(5794) <= layer3_outputs(226);
    layer4_outputs(5795) <= not((layer3_outputs(5186)) or (layer3_outputs(3524)));
    layer4_outputs(5796) <= not(layer3_outputs(5362));
    layer4_outputs(5797) <= not(layer3_outputs(6867));
    layer4_outputs(5798) <= (layer3_outputs(9938)) or (layer3_outputs(7776));
    layer4_outputs(5799) <= layer3_outputs(2009);
    layer4_outputs(5800) <= not((layer3_outputs(4684)) and (layer3_outputs(3478)));
    layer4_outputs(5801) <= not(layer3_outputs(3387));
    layer4_outputs(5802) <= layer3_outputs(8098);
    layer4_outputs(5803) <= layer3_outputs(1161);
    layer4_outputs(5804) <= layer3_outputs(8042);
    layer4_outputs(5805) <= (layer3_outputs(909)) and not (layer3_outputs(3176));
    layer4_outputs(5806) <= (layer3_outputs(4824)) and not (layer3_outputs(3251));
    layer4_outputs(5807) <= layer3_outputs(1605);
    layer4_outputs(5808) <= layer3_outputs(6208);
    layer4_outputs(5809) <= not((layer3_outputs(6013)) and (layer3_outputs(8590)));
    layer4_outputs(5810) <= layer3_outputs(1028);
    layer4_outputs(5811) <= not(layer3_outputs(5063));
    layer4_outputs(5812) <= not(layer3_outputs(5311));
    layer4_outputs(5813) <= not(layer3_outputs(702)) or (layer3_outputs(740));
    layer4_outputs(5814) <= layer3_outputs(4044);
    layer4_outputs(5815) <= not((layer3_outputs(7271)) and (layer3_outputs(1221)));
    layer4_outputs(5816) <= layer3_outputs(2844);
    layer4_outputs(5817) <= (layer3_outputs(10228)) and not (layer3_outputs(8423));
    layer4_outputs(5818) <= layer3_outputs(1222);
    layer4_outputs(5819) <= not((layer3_outputs(7150)) or (layer3_outputs(1653)));
    layer4_outputs(5820) <= (layer3_outputs(678)) xor (layer3_outputs(4497));
    layer4_outputs(5821) <= layer3_outputs(4031);
    layer4_outputs(5822) <= not(layer3_outputs(8883));
    layer4_outputs(5823) <= not(layer3_outputs(941));
    layer4_outputs(5824) <= (layer3_outputs(7693)) or (layer3_outputs(4545));
    layer4_outputs(5825) <= (layer3_outputs(9969)) and not (layer3_outputs(8525));
    layer4_outputs(5826) <= not(layer3_outputs(3745)) or (layer3_outputs(4151));
    layer4_outputs(5827) <= layer3_outputs(4805);
    layer4_outputs(5828) <= not((layer3_outputs(3625)) or (layer3_outputs(2934)));
    layer4_outputs(5829) <= not(layer3_outputs(218));
    layer4_outputs(5830) <= layer3_outputs(82);
    layer4_outputs(5831) <= (layer3_outputs(8871)) and not (layer3_outputs(3966));
    layer4_outputs(5832) <= layer3_outputs(2298);
    layer4_outputs(5833) <= layer3_outputs(8316);
    layer4_outputs(5834) <= (layer3_outputs(1133)) xor (layer3_outputs(5519));
    layer4_outputs(5835) <= layer3_outputs(513);
    layer4_outputs(5836) <= layer3_outputs(7304);
    layer4_outputs(5837) <= layer3_outputs(5848);
    layer4_outputs(5838) <= layer3_outputs(8362);
    layer4_outputs(5839) <= not(layer3_outputs(3582));
    layer4_outputs(5840) <= (layer3_outputs(7451)) or (layer3_outputs(3700));
    layer4_outputs(5841) <= (layer3_outputs(3437)) or (layer3_outputs(756));
    layer4_outputs(5842) <= (layer3_outputs(629)) or (layer3_outputs(10119));
    layer4_outputs(5843) <= not((layer3_outputs(1767)) and (layer3_outputs(3047)));
    layer4_outputs(5844) <= (layer3_outputs(6720)) and not (layer3_outputs(6023));
    layer4_outputs(5845) <= not(layer3_outputs(7700));
    layer4_outputs(5846) <= (layer3_outputs(8408)) and not (layer3_outputs(6945));
    layer4_outputs(5847) <= not(layer3_outputs(8402)) or (layer3_outputs(1199));
    layer4_outputs(5848) <= not(layer3_outputs(8046));
    layer4_outputs(5849) <= (layer3_outputs(5004)) or (layer3_outputs(2227));
    layer4_outputs(5850) <= (layer3_outputs(3357)) xor (layer3_outputs(823));
    layer4_outputs(5851) <= (layer3_outputs(3109)) xor (layer3_outputs(2542));
    layer4_outputs(5852) <= (layer3_outputs(3762)) xor (layer3_outputs(706));
    layer4_outputs(5853) <= layer3_outputs(6198);
    layer4_outputs(5854) <= (layer3_outputs(3911)) and not (layer3_outputs(9079));
    layer4_outputs(5855) <= (layer3_outputs(8180)) xor (layer3_outputs(1385));
    layer4_outputs(5856) <= not((layer3_outputs(2337)) and (layer3_outputs(2557)));
    layer4_outputs(5857) <= (layer3_outputs(5002)) and not (layer3_outputs(6162));
    layer4_outputs(5858) <= not((layer3_outputs(7203)) xor (layer3_outputs(6409)));
    layer4_outputs(5859) <= layer3_outputs(8185);
    layer4_outputs(5860) <= layer3_outputs(6847);
    layer4_outputs(5861) <= not(layer3_outputs(7409)) or (layer3_outputs(4822));
    layer4_outputs(5862) <= (layer3_outputs(4591)) and not (layer3_outputs(1339));
    layer4_outputs(5863) <= not((layer3_outputs(8637)) xor (layer3_outputs(7076)));
    layer4_outputs(5864) <= layer3_outputs(7786);
    layer4_outputs(5865) <= layer3_outputs(1408);
    layer4_outputs(5866) <= not((layer3_outputs(8040)) or (layer3_outputs(5215)));
    layer4_outputs(5867) <= layer3_outputs(1355);
    layer4_outputs(5868) <= layer3_outputs(7245);
    layer4_outputs(5869) <= not(layer3_outputs(9495)) or (layer3_outputs(194));
    layer4_outputs(5870) <= not(layer3_outputs(1016));
    layer4_outputs(5871) <= not(layer3_outputs(4088));
    layer4_outputs(5872) <= not(layer3_outputs(8796));
    layer4_outputs(5873) <= layer3_outputs(7910);
    layer4_outputs(5874) <= '0';
    layer4_outputs(5875) <= not(layer3_outputs(1872));
    layer4_outputs(5876) <= layer3_outputs(1504);
    layer4_outputs(5877) <= not(layer3_outputs(1112));
    layer4_outputs(5878) <= (layer3_outputs(6772)) and not (layer3_outputs(6099));
    layer4_outputs(5879) <= not(layer3_outputs(5007));
    layer4_outputs(5880) <= not(layer3_outputs(9803));
    layer4_outputs(5881) <= not(layer3_outputs(1163));
    layer4_outputs(5882) <= (layer3_outputs(6453)) and not (layer3_outputs(6253));
    layer4_outputs(5883) <= not((layer3_outputs(3559)) and (layer3_outputs(8421)));
    layer4_outputs(5884) <= not(layer3_outputs(7920));
    layer4_outputs(5885) <= layer3_outputs(1415);
    layer4_outputs(5886) <= (layer3_outputs(3979)) and (layer3_outputs(5629));
    layer4_outputs(5887) <= not(layer3_outputs(3933));
    layer4_outputs(5888) <= layer3_outputs(8150);
    layer4_outputs(5889) <= not((layer3_outputs(7211)) xor (layer3_outputs(4501)));
    layer4_outputs(5890) <= layer3_outputs(426);
    layer4_outputs(5891) <= not(layer3_outputs(7296));
    layer4_outputs(5892) <= not(layer3_outputs(6823));
    layer4_outputs(5893) <= layer3_outputs(7988);
    layer4_outputs(5894) <= not(layer3_outputs(2412));
    layer4_outputs(5895) <= not(layer3_outputs(4206));
    layer4_outputs(5896) <= layer3_outputs(261);
    layer4_outputs(5897) <= not(layer3_outputs(2676));
    layer4_outputs(5898) <= layer3_outputs(5754);
    layer4_outputs(5899) <= not(layer3_outputs(6186));
    layer4_outputs(5900) <= not(layer3_outputs(8649)) or (layer3_outputs(794));
    layer4_outputs(5901) <= not(layer3_outputs(5069));
    layer4_outputs(5902) <= (layer3_outputs(8051)) xor (layer3_outputs(708));
    layer4_outputs(5903) <= not((layer3_outputs(3048)) xor (layer3_outputs(4807)));
    layer4_outputs(5904) <= (layer3_outputs(8371)) or (layer3_outputs(156));
    layer4_outputs(5905) <= not(layer3_outputs(4645));
    layer4_outputs(5906) <= not((layer3_outputs(7038)) xor (layer3_outputs(1357)));
    layer4_outputs(5907) <= not((layer3_outputs(3786)) xor (layer3_outputs(4595)));
    layer4_outputs(5908) <= (layer3_outputs(9413)) or (layer3_outputs(5369));
    layer4_outputs(5909) <= layer3_outputs(5138);
    layer4_outputs(5910) <= (layer3_outputs(2736)) and not (layer3_outputs(4954));
    layer4_outputs(5911) <= not(layer3_outputs(4855));
    layer4_outputs(5912) <= '0';
    layer4_outputs(5913) <= not(layer3_outputs(6840)) or (layer3_outputs(1899));
    layer4_outputs(5914) <= (layer3_outputs(8198)) or (layer3_outputs(6705));
    layer4_outputs(5915) <= (layer3_outputs(7101)) xor (layer3_outputs(6880));
    layer4_outputs(5916) <= not((layer3_outputs(3249)) and (layer3_outputs(8388)));
    layer4_outputs(5917) <= (layer3_outputs(6904)) xor (layer3_outputs(5530));
    layer4_outputs(5918) <= layer3_outputs(10183);
    layer4_outputs(5919) <= (layer3_outputs(7085)) and (layer3_outputs(935));
    layer4_outputs(5920) <= (layer3_outputs(9328)) and (layer3_outputs(4239));
    layer4_outputs(5921) <= not((layer3_outputs(1414)) xor (layer3_outputs(7975)));
    layer4_outputs(5922) <= not(layer3_outputs(8604));
    layer4_outputs(5923) <= (layer3_outputs(5303)) or (layer3_outputs(3535));
    layer4_outputs(5924) <= not(layer3_outputs(4785));
    layer4_outputs(5925) <= not(layer3_outputs(8381));
    layer4_outputs(5926) <= not(layer3_outputs(1723));
    layer4_outputs(5927) <= (layer3_outputs(6737)) or (layer3_outputs(1151));
    layer4_outputs(5928) <= layer3_outputs(7273);
    layer4_outputs(5929) <= not((layer3_outputs(712)) xor (layer3_outputs(7925)));
    layer4_outputs(5930) <= not((layer3_outputs(2357)) xor (layer3_outputs(1052)));
    layer4_outputs(5931) <= layer3_outputs(3774);
    layer4_outputs(5932) <= layer3_outputs(4159);
    layer4_outputs(5933) <= not(layer3_outputs(1411));
    layer4_outputs(5934) <= layer3_outputs(5001);
    layer4_outputs(5935) <= not(layer3_outputs(2226));
    layer4_outputs(5936) <= not(layer3_outputs(5926));
    layer4_outputs(5937) <= (layer3_outputs(6750)) and (layer3_outputs(2903));
    layer4_outputs(5938) <= layer3_outputs(5687);
    layer4_outputs(5939) <= not(layer3_outputs(4477)) or (layer3_outputs(5505));
    layer4_outputs(5940) <= not((layer3_outputs(6758)) or (layer3_outputs(2947)));
    layer4_outputs(5941) <= not((layer3_outputs(1136)) or (layer3_outputs(2488)));
    layer4_outputs(5942) <= layer3_outputs(8851);
    layer4_outputs(5943) <= layer3_outputs(7404);
    layer4_outputs(5944) <= (layer3_outputs(1633)) or (layer3_outputs(4825));
    layer4_outputs(5945) <= '1';
    layer4_outputs(5946) <= (layer3_outputs(304)) and (layer3_outputs(1320));
    layer4_outputs(5947) <= (layer3_outputs(7475)) and not (layer3_outputs(9686));
    layer4_outputs(5948) <= not(layer3_outputs(6905));
    layer4_outputs(5949) <= not(layer3_outputs(482));
    layer4_outputs(5950) <= (layer3_outputs(4508)) and not (layer3_outputs(689));
    layer4_outputs(5951) <= not(layer3_outputs(6468));
    layer4_outputs(5952) <= layer3_outputs(9942);
    layer4_outputs(5953) <= layer3_outputs(3035);
    layer4_outputs(5954) <= not(layer3_outputs(7156));
    layer4_outputs(5955) <= layer3_outputs(3212);
    layer4_outputs(5956) <= not((layer3_outputs(6216)) or (layer3_outputs(6479)));
    layer4_outputs(5957) <= (layer3_outputs(5698)) and not (layer3_outputs(3663));
    layer4_outputs(5958) <= layer3_outputs(3416);
    layer4_outputs(5959) <= not((layer3_outputs(8414)) xor (layer3_outputs(3934)));
    layer4_outputs(5960) <= not(layer3_outputs(2683));
    layer4_outputs(5961) <= not((layer3_outputs(6099)) or (layer3_outputs(7412)));
    layer4_outputs(5962) <= layer3_outputs(8637);
    layer4_outputs(5963) <= layer3_outputs(8794);
    layer4_outputs(5964) <= layer3_outputs(4895);
    layer4_outputs(5965) <= layer3_outputs(9680);
    layer4_outputs(5966) <= (layer3_outputs(1836)) xor (layer3_outputs(5196));
    layer4_outputs(5967) <= layer3_outputs(6129);
    layer4_outputs(5968) <= not(layer3_outputs(9257));
    layer4_outputs(5969) <= not((layer3_outputs(8864)) xor (layer3_outputs(8624)));
    layer4_outputs(5970) <= not(layer3_outputs(2625)) or (layer3_outputs(1877));
    layer4_outputs(5971) <= not(layer3_outputs(4114));
    layer4_outputs(5972) <= not((layer3_outputs(7865)) xor (layer3_outputs(3380)));
    layer4_outputs(5973) <= (layer3_outputs(5973)) xor (layer3_outputs(2756));
    layer4_outputs(5974) <= layer3_outputs(6574);
    layer4_outputs(5975) <= (layer3_outputs(8683)) and not (layer3_outputs(646));
    layer4_outputs(5976) <= not(layer3_outputs(7234));
    layer4_outputs(5977) <= not((layer3_outputs(4291)) or (layer3_outputs(4062)));
    layer4_outputs(5978) <= (layer3_outputs(274)) and not (layer3_outputs(4929));
    layer4_outputs(5979) <= not((layer3_outputs(2549)) or (layer3_outputs(4124)));
    layer4_outputs(5980) <= not((layer3_outputs(7965)) or (layer3_outputs(3013)));
    layer4_outputs(5981) <= not(layer3_outputs(9461));
    layer4_outputs(5982) <= not((layer3_outputs(8299)) or (layer3_outputs(4461)));
    layer4_outputs(5983) <= layer3_outputs(975);
    layer4_outputs(5984) <= (layer3_outputs(7141)) xor (layer3_outputs(3933));
    layer4_outputs(5985) <= not(layer3_outputs(7443)) or (layer3_outputs(6165));
    layer4_outputs(5986) <= not(layer3_outputs(10060));
    layer4_outputs(5987) <= (layer3_outputs(9774)) xor (layer3_outputs(1453));
    layer4_outputs(5988) <= not(layer3_outputs(5107));
    layer4_outputs(5989) <= not(layer3_outputs(1041));
    layer4_outputs(5990) <= not(layer3_outputs(2623));
    layer4_outputs(5991) <= not((layer3_outputs(256)) xor (layer3_outputs(6604)));
    layer4_outputs(5992) <= not(layer3_outputs(5026));
    layer4_outputs(5993) <= not((layer3_outputs(5777)) and (layer3_outputs(7367)));
    layer4_outputs(5994) <= layer3_outputs(7922);
    layer4_outputs(5995) <= not(layer3_outputs(8450)) or (layer3_outputs(8825));
    layer4_outputs(5996) <= not(layer3_outputs(1934)) or (layer3_outputs(9792));
    layer4_outputs(5997) <= not(layer3_outputs(4681));
    layer4_outputs(5998) <= layer3_outputs(2261);
    layer4_outputs(5999) <= not(layer3_outputs(4703));
    layer4_outputs(6000) <= (layer3_outputs(6021)) xor (layer3_outputs(5678));
    layer4_outputs(6001) <= not(layer3_outputs(6519)) or (layer3_outputs(3021));
    layer4_outputs(6002) <= layer3_outputs(642);
    layer4_outputs(6003) <= not(layer3_outputs(4910));
    layer4_outputs(6004) <= not((layer3_outputs(1456)) xor (layer3_outputs(2619)));
    layer4_outputs(6005) <= (layer3_outputs(3577)) and (layer3_outputs(7013));
    layer4_outputs(6006) <= layer3_outputs(5863);
    layer4_outputs(6007) <= layer3_outputs(6105);
    layer4_outputs(6008) <= not((layer3_outputs(4688)) xor (layer3_outputs(9842)));
    layer4_outputs(6009) <= (layer3_outputs(3249)) or (layer3_outputs(7334));
    layer4_outputs(6010) <= not(layer3_outputs(5387)) or (layer3_outputs(5582));
    layer4_outputs(6011) <= not(layer3_outputs(3858));
    layer4_outputs(6012) <= not(layer3_outputs(3959));
    layer4_outputs(6013) <= layer3_outputs(29);
    layer4_outputs(6014) <= not((layer3_outputs(6872)) xor (layer3_outputs(6132)));
    layer4_outputs(6015) <= layer3_outputs(9428);
    layer4_outputs(6016) <= not((layer3_outputs(1532)) xor (layer3_outputs(10119)));
    layer4_outputs(6017) <= (layer3_outputs(1820)) and not (layer3_outputs(6614));
    layer4_outputs(6018) <= not(layer3_outputs(4778));
    layer4_outputs(6019) <= (layer3_outputs(4704)) xor (layer3_outputs(38));
    layer4_outputs(6020) <= not(layer3_outputs(5441));
    layer4_outputs(6021) <= not(layer3_outputs(4010)) or (layer3_outputs(4335));
    layer4_outputs(6022) <= (layer3_outputs(2068)) and (layer3_outputs(5180));
    layer4_outputs(6023) <= layer3_outputs(1263);
    layer4_outputs(6024) <= layer3_outputs(6333);
    layer4_outputs(6025) <= not(layer3_outputs(8223));
    layer4_outputs(6026) <= not(layer3_outputs(5975));
    layer4_outputs(6027) <= layer3_outputs(3190);
    layer4_outputs(6028) <= layer3_outputs(5327);
    layer4_outputs(6029) <= layer3_outputs(5805);
    layer4_outputs(6030) <= not(layer3_outputs(8934));
    layer4_outputs(6031) <= layer3_outputs(2338);
    layer4_outputs(6032) <= not((layer3_outputs(9049)) or (layer3_outputs(3946)));
    layer4_outputs(6033) <= not(layer3_outputs(8564));
    layer4_outputs(6034) <= layer3_outputs(10221);
    layer4_outputs(6035) <= layer3_outputs(9538);
    layer4_outputs(6036) <= not(layer3_outputs(8068));
    layer4_outputs(6037) <= not(layer3_outputs(2359));
    layer4_outputs(6038) <= not(layer3_outputs(3014)) or (layer3_outputs(4348));
    layer4_outputs(6039) <= not(layer3_outputs(5424));
    layer4_outputs(6040) <= not(layer3_outputs(8799));
    layer4_outputs(6041) <= layer3_outputs(3338);
    layer4_outputs(6042) <= not(layer3_outputs(6538));
    layer4_outputs(6043) <= (layer3_outputs(3452)) and not (layer3_outputs(8448));
    layer4_outputs(6044) <= not((layer3_outputs(6563)) xor (layer3_outputs(9996)));
    layer4_outputs(6045) <= layer3_outputs(3740);
    layer4_outputs(6046) <= (layer3_outputs(5654)) xor (layer3_outputs(267));
    layer4_outputs(6047) <= (layer3_outputs(3004)) and not (layer3_outputs(4016));
    layer4_outputs(6048) <= layer3_outputs(8888);
    layer4_outputs(6049) <= layer3_outputs(6424);
    layer4_outputs(6050) <= (layer3_outputs(3108)) xor (layer3_outputs(3578));
    layer4_outputs(6051) <= not((layer3_outputs(5223)) and (layer3_outputs(320)));
    layer4_outputs(6052) <= not(layer3_outputs(845));
    layer4_outputs(6053) <= not(layer3_outputs(821)) or (layer3_outputs(1687));
    layer4_outputs(6054) <= not(layer3_outputs(9205)) or (layer3_outputs(9167));
    layer4_outputs(6055) <= not(layer3_outputs(5927));
    layer4_outputs(6056) <= layer3_outputs(2788);
    layer4_outputs(6057) <= (layer3_outputs(4503)) xor (layer3_outputs(3494));
    layer4_outputs(6058) <= (layer3_outputs(7588)) or (layer3_outputs(5987));
    layer4_outputs(6059) <= (layer3_outputs(8695)) xor (layer3_outputs(1517));
    layer4_outputs(6060) <= not((layer3_outputs(4600)) or (layer3_outputs(3005)));
    layer4_outputs(6061) <= not(layer3_outputs(8091)) or (layer3_outputs(9283));
    layer4_outputs(6062) <= not(layer3_outputs(5823));
    layer4_outputs(6063) <= layer3_outputs(5397);
    layer4_outputs(6064) <= not(layer3_outputs(1650));
    layer4_outputs(6065) <= layer3_outputs(1259);
    layer4_outputs(6066) <= (layer3_outputs(6400)) or (layer3_outputs(10096));
    layer4_outputs(6067) <= not(layer3_outputs(1861));
    layer4_outputs(6068) <= not(layer3_outputs(9869));
    layer4_outputs(6069) <= not(layer3_outputs(561));
    layer4_outputs(6070) <= (layer3_outputs(6774)) xor (layer3_outputs(9321));
    layer4_outputs(6071) <= not(layer3_outputs(2926));
    layer4_outputs(6072) <= not(layer3_outputs(3977));
    layer4_outputs(6073) <= not((layer3_outputs(4024)) and (layer3_outputs(3611)));
    layer4_outputs(6074) <= not(layer3_outputs(8586));
    layer4_outputs(6075) <= not(layer3_outputs(3990)) or (layer3_outputs(4597));
    layer4_outputs(6076) <= not((layer3_outputs(8215)) xor (layer3_outputs(6030)));
    layer4_outputs(6077) <= not(layer3_outputs(4577));
    layer4_outputs(6078) <= layer3_outputs(5088);
    layer4_outputs(6079) <= not(layer3_outputs(7302));
    layer4_outputs(6080) <= (layer3_outputs(2459)) and not (layer3_outputs(5986));
    layer4_outputs(6081) <= (layer3_outputs(1181)) and not (layer3_outputs(2649));
    layer4_outputs(6082) <= not((layer3_outputs(4742)) and (layer3_outputs(5473)));
    layer4_outputs(6083) <= (layer3_outputs(378)) or (layer3_outputs(5457));
    layer4_outputs(6084) <= not((layer3_outputs(7314)) xor (layer3_outputs(2944)));
    layer4_outputs(6085) <= layer3_outputs(803);
    layer4_outputs(6086) <= not(layer3_outputs(3326));
    layer4_outputs(6087) <= (layer3_outputs(106)) and not (layer3_outputs(2388));
    layer4_outputs(6088) <= not(layer3_outputs(8234)) or (layer3_outputs(3723));
    layer4_outputs(6089) <= not(layer3_outputs(2394));
    layer4_outputs(6090) <= not((layer3_outputs(3005)) xor (layer3_outputs(8734)));
    layer4_outputs(6091) <= layer3_outputs(8857);
    layer4_outputs(6092) <= not(layer3_outputs(9142)) or (layer3_outputs(7029));
    layer4_outputs(6093) <= (layer3_outputs(7911)) and not (layer3_outputs(955));
    layer4_outputs(6094) <= layer3_outputs(4912);
    layer4_outputs(6095) <= (layer3_outputs(3059)) xor (layer3_outputs(936));
    layer4_outputs(6096) <= not((layer3_outputs(5521)) xor (layer3_outputs(7539)));
    layer4_outputs(6097) <= layer3_outputs(31);
    layer4_outputs(6098) <= not(layer3_outputs(260));
    layer4_outputs(6099) <= layer3_outputs(10005);
    layer4_outputs(6100) <= not(layer3_outputs(1364));
    layer4_outputs(6101) <= (layer3_outputs(6394)) and (layer3_outputs(2356));
    layer4_outputs(6102) <= not(layer3_outputs(9361));
    layer4_outputs(6103) <= layer3_outputs(7232);
    layer4_outputs(6104) <= layer3_outputs(7507);
    layer4_outputs(6105) <= (layer3_outputs(5271)) and not (layer3_outputs(4755));
    layer4_outputs(6106) <= (layer3_outputs(4131)) and not (layer3_outputs(10109));
    layer4_outputs(6107) <= (layer3_outputs(7291)) and (layer3_outputs(1915));
    layer4_outputs(6108) <= not(layer3_outputs(3982));
    layer4_outputs(6109) <= not(layer3_outputs(7108));
    layer4_outputs(6110) <= not(layer3_outputs(2216));
    layer4_outputs(6111) <= not(layer3_outputs(1364));
    layer4_outputs(6112) <= (layer3_outputs(2025)) xor (layer3_outputs(6518));
    layer4_outputs(6113) <= not(layer3_outputs(4430));
    layer4_outputs(6114) <= (layer3_outputs(637)) xor (layer3_outputs(6917));
    layer4_outputs(6115) <= (layer3_outputs(483)) and not (layer3_outputs(3493));
    layer4_outputs(6116) <= not(layer3_outputs(2030));
    layer4_outputs(6117) <= not(layer3_outputs(3235));
    layer4_outputs(6118) <= layer3_outputs(1199);
    layer4_outputs(6119) <= not(layer3_outputs(7639)) or (layer3_outputs(6995));
    layer4_outputs(6120) <= not(layer3_outputs(2492)) or (layer3_outputs(4715));
    layer4_outputs(6121) <= layer3_outputs(1408);
    layer4_outputs(6122) <= not(layer3_outputs(1235));
    layer4_outputs(6123) <= (layer3_outputs(6215)) and not (layer3_outputs(2870));
    layer4_outputs(6124) <= layer3_outputs(8196);
    layer4_outputs(6125) <= layer3_outputs(1781);
    layer4_outputs(6126) <= not(layer3_outputs(2097));
    layer4_outputs(6127) <= not(layer3_outputs(9));
    layer4_outputs(6128) <= not(layer3_outputs(3085));
    layer4_outputs(6129) <= not((layer3_outputs(7382)) or (layer3_outputs(5989)));
    layer4_outputs(6130) <= not((layer3_outputs(3687)) or (layer3_outputs(2629)));
    layer4_outputs(6131) <= layer3_outputs(7985);
    layer4_outputs(6132) <= layer3_outputs(5801);
    layer4_outputs(6133) <= (layer3_outputs(6712)) and (layer3_outputs(9111));
    layer4_outputs(6134) <= not(layer3_outputs(2110));
    layer4_outputs(6135) <= (layer3_outputs(8885)) and (layer3_outputs(10046));
    layer4_outputs(6136) <= layer3_outputs(8696);
    layer4_outputs(6137) <= '1';
    layer4_outputs(6138) <= not(layer3_outputs(3294));
    layer4_outputs(6139) <= layer3_outputs(5279);
    layer4_outputs(6140) <= layer3_outputs(9046);
    layer4_outputs(6141) <= not(layer3_outputs(7090));
    layer4_outputs(6142) <= layer3_outputs(5682);
    layer4_outputs(6143) <= layer3_outputs(950);
    layer4_outputs(6144) <= not((layer3_outputs(4588)) xor (layer3_outputs(3549)));
    layer4_outputs(6145) <= layer3_outputs(10052);
    layer4_outputs(6146) <= not(layer3_outputs(9465));
    layer4_outputs(6147) <= layer3_outputs(5974);
    layer4_outputs(6148) <= layer3_outputs(6564);
    layer4_outputs(6149) <= (layer3_outputs(6444)) and not (layer3_outputs(9016));
    layer4_outputs(6150) <= layer3_outputs(3624);
    layer4_outputs(6151) <= not((layer3_outputs(4984)) xor (layer3_outputs(8776)));
    layer4_outputs(6152) <= (layer3_outputs(1732)) xor (layer3_outputs(1545));
    layer4_outputs(6153) <= not(layer3_outputs(8817));
    layer4_outputs(6154) <= (layer3_outputs(6957)) or (layer3_outputs(9716));
    layer4_outputs(6155) <= layer3_outputs(208);
    layer4_outputs(6156) <= not(layer3_outputs(9190)) or (layer3_outputs(6783));
    layer4_outputs(6157) <= layer3_outputs(9576);
    layer4_outputs(6158) <= not((layer3_outputs(2956)) xor (layer3_outputs(2931)));
    layer4_outputs(6159) <= (layer3_outputs(9220)) xor (layer3_outputs(7565));
    layer4_outputs(6160) <= layer3_outputs(6039);
    layer4_outputs(6161) <= not(layer3_outputs(2087));
    layer4_outputs(6162) <= not((layer3_outputs(9403)) and (layer3_outputs(4791)));
    layer4_outputs(6163) <= not(layer3_outputs(5343));
    layer4_outputs(6164) <= (layer3_outputs(2397)) or (layer3_outputs(1));
    layer4_outputs(6165) <= not((layer3_outputs(9162)) xor (layer3_outputs(6958)));
    layer4_outputs(6166) <= layer3_outputs(7196);
    layer4_outputs(6167) <= not(layer3_outputs(7368));
    layer4_outputs(6168) <= (layer3_outputs(9324)) and not (layer3_outputs(4064));
    layer4_outputs(6169) <= not(layer3_outputs(8709));
    layer4_outputs(6170) <= layer3_outputs(8923);
    layer4_outputs(6171) <= not(layer3_outputs(2681));
    layer4_outputs(6172) <= not(layer3_outputs(292));
    layer4_outputs(6173) <= not(layer3_outputs(5750)) or (layer3_outputs(2595));
    layer4_outputs(6174) <= not(layer3_outputs(7065));
    layer4_outputs(6175) <= not((layer3_outputs(5178)) xor (layer3_outputs(1248)));
    layer4_outputs(6176) <= layer3_outputs(9271);
    layer4_outputs(6177) <= not(layer3_outputs(94));
    layer4_outputs(6178) <= (layer3_outputs(363)) or (layer3_outputs(7400));
    layer4_outputs(6179) <= not((layer3_outputs(1397)) xor (layer3_outputs(3131)));
    layer4_outputs(6180) <= (layer3_outputs(5629)) and not (layer3_outputs(9822));
    layer4_outputs(6181) <= not(layer3_outputs(6180));
    layer4_outputs(6182) <= not(layer3_outputs(1977));
    layer4_outputs(6183) <= not(layer3_outputs(2572));
    layer4_outputs(6184) <= layer3_outputs(6764);
    layer4_outputs(6185) <= not((layer3_outputs(4335)) and (layer3_outputs(2221)));
    layer4_outputs(6186) <= (layer3_outputs(210)) and not (layer3_outputs(8524));
    layer4_outputs(6187) <= not(layer3_outputs(6015));
    layer4_outputs(6188) <= not((layer3_outputs(4404)) or (layer3_outputs(5609)));
    layer4_outputs(6189) <= (layer3_outputs(7574)) or (layer3_outputs(1285));
    layer4_outputs(6190) <= (layer3_outputs(5453)) and (layer3_outputs(4369));
    layer4_outputs(6191) <= not(layer3_outputs(5847));
    layer4_outputs(6192) <= layer3_outputs(224);
    layer4_outputs(6193) <= not(layer3_outputs(2862)) or (layer3_outputs(3550));
    layer4_outputs(6194) <= layer3_outputs(9432);
    layer4_outputs(6195) <= not((layer3_outputs(6392)) or (layer3_outputs(9550)));
    layer4_outputs(6196) <= not(layer3_outputs(1512));
    layer4_outputs(6197) <= (layer3_outputs(9408)) xor (layer3_outputs(10025));
    layer4_outputs(6198) <= not((layer3_outputs(2685)) xor (layer3_outputs(7318)));
    layer4_outputs(6199) <= (layer3_outputs(2100)) or (layer3_outputs(5151));
    layer4_outputs(6200) <= not(layer3_outputs(5904)) or (layer3_outputs(7932));
    layer4_outputs(6201) <= (layer3_outputs(7231)) xor (layer3_outputs(8104));
    layer4_outputs(6202) <= not(layer3_outputs(5575));
    layer4_outputs(6203) <= layer3_outputs(3139);
    layer4_outputs(6204) <= not(layer3_outputs(1350));
    layer4_outputs(6205) <= (layer3_outputs(7557)) and (layer3_outputs(5167));
    layer4_outputs(6206) <= not(layer3_outputs(2975)) or (layer3_outputs(9117));
    layer4_outputs(6207) <= (layer3_outputs(9231)) and (layer3_outputs(2377));
    layer4_outputs(6208) <= not(layer3_outputs(4792));
    layer4_outputs(6209) <= not((layer3_outputs(3248)) xor (layer3_outputs(7505)));
    layer4_outputs(6210) <= not((layer3_outputs(5498)) or (layer3_outputs(1840)));
    layer4_outputs(6211) <= (layer3_outputs(1817)) or (layer3_outputs(4283));
    layer4_outputs(6212) <= layer3_outputs(3230);
    layer4_outputs(6213) <= layer3_outputs(4350);
    layer4_outputs(6214) <= layer3_outputs(8509);
    layer4_outputs(6215) <= (layer3_outputs(313)) xor (layer3_outputs(1795));
    layer4_outputs(6216) <= not(layer3_outputs(4305));
    layer4_outputs(6217) <= not(layer3_outputs(1060)) or (layer3_outputs(4319));
    layer4_outputs(6218) <= not(layer3_outputs(4325));
    layer4_outputs(6219) <= not((layer3_outputs(10239)) or (layer3_outputs(9762)));
    layer4_outputs(6220) <= not((layer3_outputs(1327)) xor (layer3_outputs(5569)));
    layer4_outputs(6221) <= not(layer3_outputs(3218));
    layer4_outputs(6222) <= (layer3_outputs(5222)) or (layer3_outputs(3356));
    layer4_outputs(6223) <= layer3_outputs(6335);
    layer4_outputs(6224) <= not(layer3_outputs(1068));
    layer4_outputs(6225) <= (layer3_outputs(5398)) and (layer3_outputs(6469));
    layer4_outputs(6226) <= not((layer3_outputs(7946)) xor (layer3_outputs(9383)));
    layer4_outputs(6227) <= layer3_outputs(8879);
    layer4_outputs(6228) <= (layer3_outputs(5345)) xor (layer3_outputs(10149));
    layer4_outputs(6229) <= layer3_outputs(5813);
    layer4_outputs(6230) <= layer3_outputs(6366);
    layer4_outputs(6231) <= (layer3_outputs(2009)) and not (layer3_outputs(8054));
    layer4_outputs(6232) <= (layer3_outputs(602)) or (layer3_outputs(1630));
    layer4_outputs(6233) <= layer3_outputs(3298);
    layer4_outputs(6234) <= not(layer3_outputs(5203)) or (layer3_outputs(10142));
    layer4_outputs(6235) <= not(layer3_outputs(5862)) or (layer3_outputs(3371));
    layer4_outputs(6236) <= not((layer3_outputs(4242)) xor (layer3_outputs(127)));
    layer4_outputs(6237) <= layer3_outputs(9200);
    layer4_outputs(6238) <= layer3_outputs(9826);
    layer4_outputs(6239) <= not((layer3_outputs(5584)) xor (layer3_outputs(2583)));
    layer4_outputs(6240) <= (layer3_outputs(9435)) and (layer3_outputs(9981));
    layer4_outputs(6241) <= not((layer3_outputs(44)) or (layer3_outputs(9562)));
    layer4_outputs(6242) <= not(layer3_outputs(145)) or (layer3_outputs(3824));
    layer4_outputs(6243) <= not(layer3_outputs(8376));
    layer4_outputs(6244) <= (layer3_outputs(448)) and not (layer3_outputs(9384));
    layer4_outputs(6245) <= layer3_outputs(4922);
    layer4_outputs(6246) <= not(layer3_outputs(1096)) or (layer3_outputs(9426));
    layer4_outputs(6247) <= layer3_outputs(5932);
    layer4_outputs(6248) <= not((layer3_outputs(7934)) xor (layer3_outputs(3478)));
    layer4_outputs(6249) <= not(layer3_outputs(4432));
    layer4_outputs(6250) <= not(layer3_outputs(448));
    layer4_outputs(6251) <= layer3_outputs(3917);
    layer4_outputs(6252) <= not(layer3_outputs(1970)) or (layer3_outputs(7181));
    layer4_outputs(6253) <= (layer3_outputs(8910)) or (layer3_outputs(3241));
    layer4_outputs(6254) <= layer3_outputs(6030);
    layer4_outputs(6255) <= layer3_outputs(909);
    layer4_outputs(6256) <= (layer3_outputs(8719)) or (layer3_outputs(9860));
    layer4_outputs(6257) <= not(layer3_outputs(3017)) or (layer3_outputs(3066));
    layer4_outputs(6258) <= layer3_outputs(1429);
    layer4_outputs(6259) <= not(layer3_outputs(3092)) or (layer3_outputs(11));
    layer4_outputs(6260) <= layer3_outputs(3431);
    layer4_outputs(6261) <= '0';
    layer4_outputs(6262) <= not(layer3_outputs(1273));
    layer4_outputs(6263) <= not(layer3_outputs(9684)) or (layer3_outputs(7787));
    layer4_outputs(6264) <= not(layer3_outputs(3453));
    layer4_outputs(6265) <= layer3_outputs(4441);
    layer4_outputs(6266) <= (layer3_outputs(3403)) xor (layer3_outputs(5921));
    layer4_outputs(6267) <= not(layer3_outputs(1664)) or (layer3_outputs(9073));
    layer4_outputs(6268) <= layer3_outputs(7114);
    layer4_outputs(6269) <= (layer3_outputs(8841)) and not (layer3_outputs(3205));
    layer4_outputs(6270) <= not((layer3_outputs(7732)) and (layer3_outputs(6905)));
    layer4_outputs(6271) <= not(layer3_outputs(6174));
    layer4_outputs(6272) <= layer3_outputs(7255);
    layer4_outputs(6273) <= (layer3_outputs(6571)) xor (layer3_outputs(2689));
    layer4_outputs(6274) <= not(layer3_outputs(4887));
    layer4_outputs(6275) <= not((layer3_outputs(6619)) and (layer3_outputs(3548)));
    layer4_outputs(6276) <= layer3_outputs(5842);
    layer4_outputs(6277) <= not((layer3_outputs(609)) xor (layer3_outputs(6002)));
    layer4_outputs(6278) <= not(layer3_outputs(8));
    layer4_outputs(6279) <= not(layer3_outputs(3513));
    layer4_outputs(6280) <= not((layer3_outputs(8985)) and (layer3_outputs(6129)));
    layer4_outputs(6281) <= layer3_outputs(3596);
    layer4_outputs(6282) <= not(layer3_outputs(5320));
    layer4_outputs(6283) <= (layer3_outputs(10082)) and not (layer3_outputs(1791));
    layer4_outputs(6284) <= layer3_outputs(6042);
    layer4_outputs(6285) <= layer3_outputs(1069);
    layer4_outputs(6286) <= not(layer3_outputs(113));
    layer4_outputs(6287) <= (layer3_outputs(5799)) or (layer3_outputs(9608));
    layer4_outputs(6288) <= layer3_outputs(7326);
    layer4_outputs(6289) <= not(layer3_outputs(800));
    layer4_outputs(6290) <= layer3_outputs(4202);
    layer4_outputs(6291) <= (layer3_outputs(6786)) and not (layer3_outputs(3098));
    layer4_outputs(6292) <= layer3_outputs(7924);
    layer4_outputs(6293) <= layer3_outputs(389);
    layer4_outputs(6294) <= layer3_outputs(5240);
    layer4_outputs(6295) <= not(layer3_outputs(2034));
    layer4_outputs(6296) <= not(layer3_outputs(6185));
    layer4_outputs(6297) <= not((layer3_outputs(9220)) xor (layer3_outputs(153)));
    layer4_outputs(6298) <= '0';
    layer4_outputs(6299) <= not(layer3_outputs(8879));
    layer4_outputs(6300) <= (layer3_outputs(386)) and not (layer3_outputs(9560));
    layer4_outputs(6301) <= not(layer3_outputs(9651));
    layer4_outputs(6302) <= not(layer3_outputs(7140)) or (layer3_outputs(5808));
    layer4_outputs(6303) <= not((layer3_outputs(2348)) and (layer3_outputs(2358)));
    layer4_outputs(6304) <= layer3_outputs(622);
    layer4_outputs(6305) <= layer3_outputs(136);
    layer4_outputs(6306) <= layer3_outputs(7059);
    layer4_outputs(6307) <= (layer3_outputs(9042)) xor (layer3_outputs(2587));
    layer4_outputs(6308) <= layer3_outputs(6609);
    layer4_outputs(6309) <= (layer3_outputs(9166)) xor (layer3_outputs(5726));
    layer4_outputs(6310) <= not(layer3_outputs(5916));
    layer4_outputs(6311) <= layer3_outputs(3386);
    layer4_outputs(6312) <= layer3_outputs(1190);
    layer4_outputs(6313) <= not((layer3_outputs(9218)) and (layer3_outputs(846)));
    layer4_outputs(6314) <= layer3_outputs(7771);
    layer4_outputs(6315) <= layer3_outputs(9587);
    layer4_outputs(6316) <= (layer3_outputs(8147)) or (layer3_outputs(10144));
    layer4_outputs(6317) <= not((layer3_outputs(5544)) xor (layer3_outputs(737)));
    layer4_outputs(6318) <= not(layer3_outputs(2851)) or (layer3_outputs(2810));
    layer4_outputs(6319) <= not(layer3_outputs(2410)) or (layer3_outputs(3153));
    layer4_outputs(6320) <= (layer3_outputs(9139)) and (layer3_outputs(2560));
    layer4_outputs(6321) <= not(layer3_outputs(8288));
    layer4_outputs(6322) <= not((layer3_outputs(5899)) or (layer3_outputs(6334)));
    layer4_outputs(6323) <= (layer3_outputs(3955)) and not (layer3_outputs(3083));
    layer4_outputs(6324) <= not((layer3_outputs(3121)) and (layer3_outputs(8887)));
    layer4_outputs(6325) <= layer3_outputs(1958);
    layer4_outputs(6326) <= not(layer3_outputs(7168)) or (layer3_outputs(10026));
    layer4_outputs(6327) <= layer3_outputs(2038);
    layer4_outputs(6328) <= layer3_outputs(4746);
    layer4_outputs(6329) <= layer3_outputs(5881);
    layer4_outputs(6330) <= layer3_outputs(9070);
    layer4_outputs(6331) <= not((layer3_outputs(9566)) or (layer3_outputs(3430)));
    layer4_outputs(6332) <= (layer3_outputs(7082)) and (layer3_outputs(3177));
    layer4_outputs(6333) <= not((layer3_outputs(2840)) xor (layer3_outputs(8934)));
    layer4_outputs(6334) <= layer3_outputs(7551);
    layer4_outputs(6335) <= not(layer3_outputs(1787)) or (layer3_outputs(3830));
    layer4_outputs(6336) <= not(layer3_outputs(3619));
    layer4_outputs(6337) <= (layer3_outputs(9436)) and (layer3_outputs(9002));
    layer4_outputs(6338) <= not((layer3_outputs(8142)) xor (layer3_outputs(7034)));
    layer4_outputs(6339) <= not(layer3_outputs(2714));
    layer4_outputs(6340) <= layer3_outputs(3501);
    layer4_outputs(6341) <= layer3_outputs(2482);
    layer4_outputs(6342) <= layer3_outputs(2639);
    layer4_outputs(6343) <= layer3_outputs(7603);
    layer4_outputs(6344) <= not((layer3_outputs(7052)) and (layer3_outputs(6120)));
    layer4_outputs(6345) <= not(layer3_outputs(6489)) or (layer3_outputs(1096));
    layer4_outputs(6346) <= layer3_outputs(8659);
    layer4_outputs(6347) <= not(layer3_outputs(6539));
    layer4_outputs(6348) <= layer3_outputs(295);
    layer4_outputs(6349) <= not(layer3_outputs(349));
    layer4_outputs(6350) <= not((layer3_outputs(4175)) xor (layer3_outputs(9040)));
    layer4_outputs(6351) <= not(layer3_outputs(5417));
    layer4_outputs(6352) <= (layer3_outputs(10197)) and not (layer3_outputs(5232));
    layer4_outputs(6353) <= (layer3_outputs(6277)) or (layer3_outputs(9485));
    layer4_outputs(6354) <= not(layer3_outputs(7977));
    layer4_outputs(6355) <= (layer3_outputs(4927)) and not (layer3_outputs(4753));
    layer4_outputs(6356) <= not(layer3_outputs(2301)) or (layer3_outputs(3430));
    layer4_outputs(6357) <= not((layer3_outputs(6447)) and (layer3_outputs(1110)));
    layer4_outputs(6358) <= not((layer3_outputs(2764)) xor (layer3_outputs(2151)));
    layer4_outputs(6359) <= not(layer3_outputs(6911));
    layer4_outputs(6360) <= not(layer3_outputs(3076));
    layer4_outputs(6361) <= (layer3_outputs(146)) and (layer3_outputs(6116));
    layer4_outputs(6362) <= layer3_outputs(5404);
    layer4_outputs(6363) <= not((layer3_outputs(7298)) xor (layer3_outputs(5514)));
    layer4_outputs(6364) <= not((layer3_outputs(10041)) and (layer3_outputs(8029)));
    layer4_outputs(6365) <= layer3_outputs(4496);
    layer4_outputs(6366) <= not(layer3_outputs(10082)) or (layer3_outputs(4441));
    layer4_outputs(6367) <= not((layer3_outputs(3704)) or (layer3_outputs(8231)));
    layer4_outputs(6368) <= not(layer3_outputs(1689));
    layer4_outputs(6369) <= not(layer3_outputs(8177));
    layer4_outputs(6370) <= not(layer3_outputs(4848));
    layer4_outputs(6371) <= not((layer3_outputs(10227)) or (layer3_outputs(4449)));
    layer4_outputs(6372) <= not(layer3_outputs(840));
    layer4_outputs(6373) <= not(layer3_outputs(9721)) or (layer3_outputs(7225));
    layer4_outputs(6374) <= not(layer3_outputs(6227));
    layer4_outputs(6375) <= layer3_outputs(4984);
    layer4_outputs(6376) <= '0';
    layer4_outputs(6377) <= layer3_outputs(10233);
    layer4_outputs(6378) <= layer3_outputs(5423);
    layer4_outputs(6379) <= not(layer3_outputs(986));
    layer4_outputs(6380) <= not(layer3_outputs(6152));
    layer4_outputs(6381) <= not(layer3_outputs(1919));
    layer4_outputs(6382) <= not((layer3_outputs(9422)) or (layer3_outputs(679)));
    layer4_outputs(6383) <= not(layer3_outputs(9567));
    layer4_outputs(6384) <= not((layer3_outputs(2583)) xor (layer3_outputs(2664)));
    layer4_outputs(6385) <= (layer3_outputs(8781)) xor (layer3_outputs(4795));
    layer4_outputs(6386) <= layer3_outputs(7018);
    layer4_outputs(6387) <= layer3_outputs(5043);
    layer4_outputs(6388) <= not((layer3_outputs(4322)) or (layer3_outputs(446)));
    layer4_outputs(6389) <= '1';
    layer4_outputs(6390) <= not(layer3_outputs(4192));
    layer4_outputs(6391) <= not(layer3_outputs(4091));
    layer4_outputs(6392) <= layer3_outputs(842);
    layer4_outputs(6393) <= (layer3_outputs(10128)) xor (layer3_outputs(3359));
    layer4_outputs(6394) <= '0';
    layer4_outputs(6395) <= layer3_outputs(7277);
    layer4_outputs(6396) <= not(layer3_outputs(170));
    layer4_outputs(6397) <= not(layer3_outputs(4491));
    layer4_outputs(6398) <= not(layer3_outputs(8031));
    layer4_outputs(6399) <= not(layer3_outputs(1528));
    layer4_outputs(6400) <= not(layer3_outputs(8849));
    layer4_outputs(6401) <= layer3_outputs(9173);
    layer4_outputs(6402) <= layer3_outputs(4539);
    layer4_outputs(6403) <= layer3_outputs(2695);
    layer4_outputs(6404) <= not((layer3_outputs(179)) xor (layer3_outputs(1825)));
    layer4_outputs(6405) <= not((layer3_outputs(8409)) or (layer3_outputs(40)));
    layer4_outputs(6406) <= layer3_outputs(4742);
    layer4_outputs(6407) <= layer3_outputs(7202);
    layer4_outputs(6408) <= (layer3_outputs(9966)) and not (layer3_outputs(1799));
    layer4_outputs(6409) <= not(layer3_outputs(4020));
    layer4_outputs(6410) <= layer3_outputs(7800);
    layer4_outputs(6411) <= not(layer3_outputs(3914));
    layer4_outputs(6412) <= not(layer3_outputs(3196));
    layer4_outputs(6413) <= layer3_outputs(906);
    layer4_outputs(6414) <= not(layer3_outputs(1196)) or (layer3_outputs(4872));
    layer4_outputs(6415) <= not(layer3_outputs(8540));
    layer4_outputs(6416) <= (layer3_outputs(4774)) xor (layer3_outputs(2780));
    layer4_outputs(6417) <= (layer3_outputs(5855)) xor (layer3_outputs(9389));
    layer4_outputs(6418) <= not((layer3_outputs(6292)) and (layer3_outputs(135)));
    layer4_outputs(6419) <= '0';
    layer4_outputs(6420) <= layer3_outputs(8677);
    layer4_outputs(6421) <= not(layer3_outputs(3913));
    layer4_outputs(6422) <= not(layer3_outputs(4007));
    layer4_outputs(6423) <= not(layer3_outputs(7503)) or (layer3_outputs(105));
    layer4_outputs(6424) <= not(layer3_outputs(9270)) or (layer3_outputs(429));
    layer4_outputs(6425) <= (layer3_outputs(4596)) and not (layer3_outputs(1303));
    layer4_outputs(6426) <= not((layer3_outputs(5588)) and (layer3_outputs(7276)));
    layer4_outputs(6427) <= not(layer3_outputs(8830));
    layer4_outputs(6428) <= layer3_outputs(4820);
    layer4_outputs(6429) <= not((layer3_outputs(10172)) xor (layer3_outputs(3663)));
    layer4_outputs(6430) <= not(layer3_outputs(6887));
    layer4_outputs(6431) <= layer3_outputs(4709);
    layer4_outputs(6432) <= (layer3_outputs(3811)) or (layer3_outputs(2237));
    layer4_outputs(6433) <= layer3_outputs(3462);
    layer4_outputs(6434) <= not(layer3_outputs(7978));
    layer4_outputs(6435) <= not(layer3_outputs(9216));
    layer4_outputs(6436) <= layer3_outputs(9795);
    layer4_outputs(6437) <= not(layer3_outputs(229));
    layer4_outputs(6438) <= layer3_outputs(3349);
    layer4_outputs(6439) <= not(layer3_outputs(2734));
    layer4_outputs(6440) <= not((layer3_outputs(4938)) xor (layer3_outputs(6126)));
    layer4_outputs(6441) <= not(layer3_outputs(3110));
    layer4_outputs(6442) <= (layer3_outputs(7069)) xor (layer3_outputs(3203));
    layer4_outputs(6443) <= not(layer3_outputs(4126));
    layer4_outputs(6444) <= layer3_outputs(7760);
    layer4_outputs(6445) <= not((layer3_outputs(608)) or (layer3_outputs(6303)));
    layer4_outputs(6446) <= not(layer3_outputs(10237));
    layer4_outputs(6447) <= not((layer3_outputs(3855)) or (layer3_outputs(7692)));
    layer4_outputs(6448) <= not((layer3_outputs(6536)) xor (layer3_outputs(2301)));
    layer4_outputs(6449) <= not((layer3_outputs(1218)) xor (layer3_outputs(21)));
    layer4_outputs(6450) <= layer3_outputs(7619);
    layer4_outputs(6451) <= (layer3_outputs(6061)) and not (layer3_outputs(5502));
    layer4_outputs(6452) <= layer3_outputs(2704);
    layer4_outputs(6453) <= not((layer3_outputs(8164)) and (layer3_outputs(1231)));
    layer4_outputs(6454) <= layer3_outputs(1188);
    layer4_outputs(6455) <= not(layer3_outputs(8672)) or (layer3_outputs(6691));
    layer4_outputs(6456) <= not((layer3_outputs(2673)) xor (layer3_outputs(7945)));
    layer4_outputs(6457) <= not(layer3_outputs(7331)) or (layer3_outputs(3450));
    layer4_outputs(6458) <= not((layer3_outputs(6224)) and (layer3_outputs(3343)));
    layer4_outputs(6459) <= layer3_outputs(499);
    layer4_outputs(6460) <= (layer3_outputs(4950)) and not (layer3_outputs(9542));
    layer4_outputs(6461) <= layer3_outputs(5280);
    layer4_outputs(6462) <= (layer3_outputs(4510)) xor (layer3_outputs(6067));
    layer4_outputs(6463) <= layer3_outputs(6585);
    layer4_outputs(6464) <= not(layer3_outputs(6328));
    layer4_outputs(6465) <= not(layer3_outputs(1714)) or (layer3_outputs(7911));
    layer4_outputs(6466) <= not((layer3_outputs(1328)) xor (layer3_outputs(1050)));
    layer4_outputs(6467) <= '0';
    layer4_outputs(6468) <= '1';
    layer4_outputs(6469) <= not(layer3_outputs(7189));
    layer4_outputs(6470) <= (layer3_outputs(9805)) xor (layer3_outputs(7746));
    layer4_outputs(6471) <= not(layer3_outputs(905));
    layer4_outputs(6472) <= (layer3_outputs(9285)) and not (layer3_outputs(4679));
    layer4_outputs(6473) <= not(layer3_outputs(2294)) or (layer3_outputs(8404));
    layer4_outputs(6474) <= not(layer3_outputs(6060)) or (layer3_outputs(5023));
    layer4_outputs(6475) <= layer3_outputs(5475);
    layer4_outputs(6476) <= (layer3_outputs(2791)) or (layer3_outputs(458));
    layer4_outputs(6477) <= not(layer3_outputs(5820));
    layer4_outputs(6478) <= layer3_outputs(1546);
    layer4_outputs(6479) <= layer3_outputs(3080);
    layer4_outputs(6480) <= not((layer3_outputs(3161)) or (layer3_outputs(5490)));
    layer4_outputs(6481) <= not(layer3_outputs(3824));
    layer4_outputs(6482) <= layer3_outputs(2878);
    layer4_outputs(6483) <= not((layer3_outputs(4720)) and (layer3_outputs(5002)));
    layer4_outputs(6484) <= (layer3_outputs(4793)) and not (layer3_outputs(1383));
    layer4_outputs(6485) <= layer3_outputs(6008);
    layer4_outputs(6486) <= layer3_outputs(8858);
    layer4_outputs(6487) <= layer3_outputs(9961);
    layer4_outputs(6488) <= not((layer3_outputs(9195)) or (layer3_outputs(116)));
    layer4_outputs(6489) <= (layer3_outputs(4947)) and (layer3_outputs(8999));
    layer4_outputs(6490) <= layer3_outputs(6870);
    layer4_outputs(6491) <= layer3_outputs(5413);
    layer4_outputs(6492) <= (layer3_outputs(4093)) or (layer3_outputs(2755));
    layer4_outputs(6493) <= (layer3_outputs(1522)) or (layer3_outputs(1658));
    layer4_outputs(6494) <= (layer3_outputs(9493)) xor (layer3_outputs(10038));
    layer4_outputs(6495) <= not(layer3_outputs(90));
    layer4_outputs(6496) <= not((layer3_outputs(9251)) xor (layer3_outputs(8173)));
    layer4_outputs(6497) <= not(layer3_outputs(6084));
    layer4_outputs(6498) <= not((layer3_outputs(2218)) xor (layer3_outputs(4869)));
    layer4_outputs(6499) <= layer3_outputs(5670);
    layer4_outputs(6500) <= (layer3_outputs(4127)) and not (layer3_outputs(6038));
    layer4_outputs(6501) <= layer3_outputs(3097);
    layer4_outputs(6502) <= not((layer3_outputs(9301)) xor (layer3_outputs(4789)));
    layer4_outputs(6503) <= (layer3_outputs(338)) and (layer3_outputs(7655));
    layer4_outputs(6504) <= not(layer3_outputs(9859));
    layer4_outputs(6505) <= not(layer3_outputs(6043)) or (layer3_outputs(372));
    layer4_outputs(6506) <= layer3_outputs(9288);
    layer4_outputs(6507) <= (layer3_outputs(10132)) xor (layer3_outputs(2389));
    layer4_outputs(6508) <= not(layer3_outputs(3684)) or (layer3_outputs(5464));
    layer4_outputs(6509) <= not(layer3_outputs(5255));
    layer4_outputs(6510) <= (layer3_outputs(5734)) xor (layer3_outputs(610));
    layer4_outputs(6511) <= (layer3_outputs(5766)) xor (layer3_outputs(7365));
    layer4_outputs(6512) <= not(layer3_outputs(8963));
    layer4_outputs(6513) <= not(layer3_outputs(5379));
    layer4_outputs(6514) <= (layer3_outputs(2835)) xor (layer3_outputs(3614));
    layer4_outputs(6515) <= not((layer3_outputs(9793)) or (layer3_outputs(5284)));
    layer4_outputs(6516) <= not(layer3_outputs(1998));
    layer4_outputs(6517) <= not((layer3_outputs(709)) and (layer3_outputs(8460)));
    layer4_outputs(6518) <= not((layer3_outputs(7964)) or (layer3_outputs(9554)));
    layer4_outputs(6519) <= layer3_outputs(4304);
    layer4_outputs(6520) <= not(layer3_outputs(669));
    layer4_outputs(6521) <= not((layer3_outputs(1104)) or (layer3_outputs(5545)));
    layer4_outputs(6522) <= layer3_outputs(10204);
    layer4_outputs(6523) <= layer3_outputs(6157);
    layer4_outputs(6524) <= not(layer3_outputs(4118)) or (layer3_outputs(6049));
    layer4_outputs(6525) <= layer3_outputs(2773);
    layer4_outputs(6526) <= not(layer3_outputs(2269));
    layer4_outputs(6527) <= (layer3_outputs(5825)) and not (layer3_outputs(5759));
    layer4_outputs(6528) <= (layer3_outputs(1708)) xor (layer3_outputs(2852));
    layer4_outputs(6529) <= not(layer3_outputs(5821));
    layer4_outputs(6530) <= not((layer3_outputs(7254)) xor (layer3_outputs(1663)));
    layer4_outputs(6531) <= not(layer3_outputs(9512)) or (layer3_outputs(8441));
    layer4_outputs(6532) <= layer3_outputs(3048);
    layer4_outputs(6533) <= layer3_outputs(2843);
    layer4_outputs(6534) <= layer3_outputs(3412);
    layer4_outputs(6535) <= not(layer3_outputs(1233));
    layer4_outputs(6536) <= not((layer3_outputs(3024)) and (layer3_outputs(2070)));
    layer4_outputs(6537) <= (layer3_outputs(1640)) and not (layer3_outputs(3174));
    layer4_outputs(6538) <= layer3_outputs(6106);
    layer4_outputs(6539) <= not(layer3_outputs(9909));
    layer4_outputs(6540) <= not((layer3_outputs(1244)) xor (layer3_outputs(8334)));
    layer4_outputs(6541) <= layer3_outputs(5496);
    layer4_outputs(6542) <= not(layer3_outputs(4893));
    layer4_outputs(6543) <= not(layer3_outputs(5417));
    layer4_outputs(6544) <= '0';
    layer4_outputs(6545) <= (layer3_outputs(1246)) and not (layer3_outputs(8132));
    layer4_outputs(6546) <= not(layer3_outputs(2032));
    layer4_outputs(6547) <= not((layer3_outputs(2970)) or (layer3_outputs(9814)));
    layer4_outputs(6548) <= not((layer3_outputs(1486)) xor (layer3_outputs(8261)));
    layer4_outputs(6549) <= not(layer3_outputs(5330)) or (layer3_outputs(5692));
    layer4_outputs(6550) <= layer3_outputs(7868);
    layer4_outputs(6551) <= not(layer3_outputs(1480));
    layer4_outputs(6552) <= not((layer3_outputs(5081)) or (layer3_outputs(2743)));
    layer4_outputs(6553) <= not(layer3_outputs(452));
    layer4_outputs(6554) <= layer3_outputs(9534);
    layer4_outputs(6555) <= not((layer3_outputs(8238)) and (layer3_outputs(4165)));
    layer4_outputs(6556) <= not((layer3_outputs(3618)) xor (layer3_outputs(4816)));
    layer4_outputs(6557) <= not(layer3_outputs(9536)) or (layer3_outputs(1734));
    layer4_outputs(6558) <= layer3_outputs(4530);
    layer4_outputs(6559) <= (layer3_outputs(8861)) and not (layer3_outputs(2767));
    layer4_outputs(6560) <= not((layer3_outputs(9715)) xor (layer3_outputs(3058)));
    layer4_outputs(6561) <= (layer3_outputs(3381)) xor (layer3_outputs(2487));
    layer4_outputs(6562) <= (layer3_outputs(9440)) or (layer3_outputs(4129));
    layer4_outputs(6563) <= not((layer3_outputs(373)) or (layer3_outputs(733)));
    layer4_outputs(6564) <= not(layer3_outputs(2069));
    layer4_outputs(6565) <= (layer3_outputs(3758)) xor (layer3_outputs(447));
    layer4_outputs(6566) <= not((layer3_outputs(2053)) and (layer3_outputs(860)));
    layer4_outputs(6567) <= layer3_outputs(7912);
    layer4_outputs(6568) <= layer3_outputs(7903);
    layer4_outputs(6569) <= (layer3_outputs(6716)) xor (layer3_outputs(1541));
    layer4_outputs(6570) <= (layer3_outputs(8229)) and not (layer3_outputs(2429));
    layer4_outputs(6571) <= not(layer3_outputs(220));
    layer4_outputs(6572) <= not(layer3_outputs(2231));
    layer4_outputs(6573) <= not(layer3_outputs(768));
    layer4_outputs(6574) <= (layer3_outputs(4140)) and (layer3_outputs(2093));
    layer4_outputs(6575) <= layer3_outputs(4149);
    layer4_outputs(6576) <= not(layer3_outputs(2138));
    layer4_outputs(6577) <= layer3_outputs(8468);
    layer4_outputs(6578) <= not((layer3_outputs(3564)) xor (layer3_outputs(4051)));
    layer4_outputs(6579) <= layer3_outputs(2352);
    layer4_outputs(6580) <= not(layer3_outputs(1085)) or (layer3_outputs(8390));
    layer4_outputs(6581) <= (layer3_outputs(7298)) xor (layer3_outputs(2573));
    layer4_outputs(6582) <= (layer3_outputs(1198)) and (layer3_outputs(3131));
    layer4_outputs(6583) <= layer3_outputs(4384);
    layer4_outputs(6584) <= not((layer3_outputs(8599)) or (layer3_outputs(2581)));
    layer4_outputs(6585) <= (layer3_outputs(7094)) xor (layer3_outputs(3234));
    layer4_outputs(6586) <= not(layer3_outputs(9170));
    layer4_outputs(6587) <= not(layer3_outputs(9275));
    layer4_outputs(6588) <= not(layer3_outputs(1689));
    layer4_outputs(6589) <= not((layer3_outputs(1302)) or (layer3_outputs(8446)));
    layer4_outputs(6590) <= (layer3_outputs(1937)) and not (layer3_outputs(5005));
    layer4_outputs(6591) <= not(layer3_outputs(4584));
    layer4_outputs(6592) <= layer3_outputs(8250);
    layer4_outputs(6593) <= (layer3_outputs(9609)) or (layer3_outputs(3790));
    layer4_outputs(6594) <= layer3_outputs(8256);
    layer4_outputs(6595) <= not(layer3_outputs(4641)) or (layer3_outputs(1806));
    layer4_outputs(6596) <= not(layer3_outputs(9320));
    layer4_outputs(6597) <= layer3_outputs(1602);
    layer4_outputs(6598) <= not((layer3_outputs(4345)) xor (layer3_outputs(6387)));
    layer4_outputs(6599) <= layer3_outputs(7500);
    layer4_outputs(6600) <= not((layer3_outputs(39)) xor (layer3_outputs(4708)));
    layer4_outputs(6601) <= (layer3_outputs(6039)) or (layer3_outputs(2486));
    layer4_outputs(6602) <= layer3_outputs(2039);
    layer4_outputs(6603) <= not(layer3_outputs(5351));
    layer4_outputs(6604) <= layer3_outputs(8749);
    layer4_outputs(6605) <= not(layer3_outputs(2613));
    layer4_outputs(6606) <= layer3_outputs(9795);
    layer4_outputs(6607) <= not(layer3_outputs(651));
    layer4_outputs(6608) <= layer3_outputs(3996);
    layer4_outputs(6609) <= not(layer3_outputs(156));
    layer4_outputs(6610) <= not(layer3_outputs(1627));
    layer4_outputs(6611) <= layer3_outputs(8853);
    layer4_outputs(6612) <= '0';
    layer4_outputs(6613) <= not((layer3_outputs(4109)) xor (layer3_outputs(2488)));
    layer4_outputs(6614) <= not(layer3_outputs(8983));
    layer4_outputs(6615) <= layer3_outputs(2240);
    layer4_outputs(6616) <= layer3_outputs(6131);
    layer4_outputs(6617) <= not(layer3_outputs(7012)) or (layer3_outputs(9490));
    layer4_outputs(6618) <= layer3_outputs(6384);
    layer4_outputs(6619) <= layer3_outputs(4527);
    layer4_outputs(6620) <= layer3_outputs(6121);
    layer4_outputs(6621) <= (layer3_outputs(1319)) and not (layer3_outputs(7484));
    layer4_outputs(6622) <= layer3_outputs(3221);
    layer4_outputs(6623) <= layer3_outputs(830);
    layer4_outputs(6624) <= layer3_outputs(6916);
    layer4_outputs(6625) <= (layer3_outputs(7542)) and not (layer3_outputs(750));
    layer4_outputs(6626) <= layer3_outputs(3864);
    layer4_outputs(6627) <= not(layer3_outputs(7318)) or (layer3_outputs(5047));
    layer4_outputs(6628) <= (layer3_outputs(9497)) or (layer3_outputs(2534));
    layer4_outputs(6629) <= not((layer3_outputs(8878)) and (layer3_outputs(5365)));
    layer4_outputs(6630) <= not((layer3_outputs(8510)) or (layer3_outputs(233)));
    layer4_outputs(6631) <= not(layer3_outputs(7010));
    layer4_outputs(6632) <= not((layer3_outputs(4153)) and (layer3_outputs(4230)));
    layer4_outputs(6633) <= not(layer3_outputs(5363));
    layer4_outputs(6634) <= layer3_outputs(7479);
    layer4_outputs(6635) <= not(layer3_outputs(7245)) or (layer3_outputs(1805));
    layer4_outputs(6636) <= not((layer3_outputs(9803)) xor (layer3_outputs(2096)));
    layer4_outputs(6637) <= '1';
    layer4_outputs(6638) <= layer3_outputs(9478);
    layer4_outputs(6639) <= not(layer3_outputs(6626));
    layer4_outputs(6640) <= not((layer3_outputs(5366)) and (layer3_outputs(7714)));
    layer4_outputs(6641) <= '1';
    layer4_outputs(6642) <= not((layer3_outputs(657)) and (layer3_outputs(6243)));
    layer4_outputs(6643) <= not((layer3_outputs(1145)) or (layer3_outputs(7299)));
    layer4_outputs(6644) <= layer3_outputs(9171);
    layer4_outputs(6645) <= (layer3_outputs(8155)) and not (layer3_outputs(9414));
    layer4_outputs(6646) <= layer3_outputs(9742);
    layer4_outputs(6647) <= not(layer3_outputs(8615));
    layer4_outputs(6648) <= layer3_outputs(8348);
    layer4_outputs(6649) <= not((layer3_outputs(9420)) xor (layer3_outputs(4013)));
    layer4_outputs(6650) <= not(layer3_outputs(6517));
    layer4_outputs(6651) <= not((layer3_outputs(896)) or (layer3_outputs(5999)));
    layer4_outputs(6652) <= not((layer3_outputs(774)) xor (layer3_outputs(8422)));
    layer4_outputs(6653) <= layer3_outputs(7521);
    layer4_outputs(6654) <= not(layer3_outputs(1362));
    layer4_outputs(6655) <= not((layer3_outputs(5515)) and (layer3_outputs(6971)));
    layer4_outputs(6656) <= layer3_outputs(5803);
    layer4_outputs(6657) <= not((layer3_outputs(5484)) and (layer3_outputs(1863)));
    layer4_outputs(6658) <= not(layer3_outputs(8235));
    layer4_outputs(6659) <= not(layer3_outputs(4042));
    layer4_outputs(6660) <= layer3_outputs(3008);
    layer4_outputs(6661) <= layer3_outputs(1087);
    layer4_outputs(6662) <= (layer3_outputs(2700)) and (layer3_outputs(10170));
    layer4_outputs(6663) <= (layer3_outputs(6611)) xor (layer3_outputs(4291));
    layer4_outputs(6664) <= (layer3_outputs(4459)) and not (layer3_outputs(7330));
    layer4_outputs(6665) <= layer3_outputs(2951);
    layer4_outputs(6666) <= layer3_outputs(894);
    layer4_outputs(6667) <= layer3_outputs(7002);
    layer4_outputs(6668) <= not((layer3_outputs(6331)) xor (layer3_outputs(6364)));
    layer4_outputs(6669) <= layer3_outputs(566);
    layer4_outputs(6670) <= layer3_outputs(5185);
    layer4_outputs(6671) <= not(layer3_outputs(9151));
    layer4_outputs(6672) <= layer3_outputs(4936);
    layer4_outputs(6673) <= layer3_outputs(8249);
    layer4_outputs(6674) <= layer3_outputs(4575);
    layer4_outputs(6675) <= not(layer3_outputs(3368));
    layer4_outputs(6676) <= not(layer3_outputs(8714));
    layer4_outputs(6677) <= not(layer3_outputs(2381));
    layer4_outputs(6678) <= not(layer3_outputs(3306));
    layer4_outputs(6679) <= (layer3_outputs(9548)) xor (layer3_outputs(7627));
    layer4_outputs(6680) <= not(layer3_outputs(9896));
    layer4_outputs(6681) <= not(layer3_outputs(4250));
    layer4_outputs(6682) <= (layer3_outputs(2360)) and (layer3_outputs(5489));
    layer4_outputs(6683) <= not((layer3_outputs(5310)) xor (layer3_outputs(6409)));
    layer4_outputs(6684) <= not(layer3_outputs(2600));
    layer4_outputs(6685) <= layer3_outputs(1423);
    layer4_outputs(6686) <= not(layer3_outputs(1052));
    layer4_outputs(6687) <= layer3_outputs(9642);
    layer4_outputs(6688) <= layer3_outputs(8251);
    layer4_outputs(6689) <= (layer3_outputs(5998)) xor (layer3_outputs(454));
    layer4_outputs(6690) <= not(layer3_outputs(2389));
    layer4_outputs(6691) <= not(layer3_outputs(402));
    layer4_outputs(6692) <= not(layer3_outputs(2586));
    layer4_outputs(6693) <= (layer3_outputs(3368)) and not (layer3_outputs(1298));
    layer4_outputs(6694) <= not(layer3_outputs(7233));
    layer4_outputs(6695) <= not((layer3_outputs(5824)) and (layer3_outputs(6544)));
    layer4_outputs(6696) <= not(layer3_outputs(5320));
    layer4_outputs(6697) <= not((layer3_outputs(9380)) or (layer3_outputs(3029)));
    layer4_outputs(6698) <= not((layer3_outputs(9876)) xor (layer3_outputs(6468)));
    layer4_outputs(6699) <= layer3_outputs(1983);
    layer4_outputs(6700) <= not(layer3_outputs(2813)) or (layer3_outputs(9058));
    layer4_outputs(6701) <= not(layer3_outputs(4568)) or (layer3_outputs(9272));
    layer4_outputs(6702) <= not(layer3_outputs(9956)) or (layer3_outputs(6306));
    layer4_outputs(6703) <= layer3_outputs(1742);
    layer4_outputs(6704) <= layer3_outputs(263);
    layer4_outputs(6705) <= not(layer3_outputs(585));
    layer4_outputs(6706) <= not(layer3_outputs(2414)) or (layer3_outputs(7139));
    layer4_outputs(6707) <= (layer3_outputs(9429)) and not (layer3_outputs(3082));
    layer4_outputs(6708) <= not((layer3_outputs(2621)) xor (layer3_outputs(2968)));
    layer4_outputs(6709) <= not((layer3_outputs(4445)) xor (layer3_outputs(3141)));
    layer4_outputs(6710) <= layer3_outputs(4097);
    layer4_outputs(6711) <= (layer3_outputs(1249)) xor (layer3_outputs(2287));
    layer4_outputs(6712) <= not((layer3_outputs(8023)) xor (layer3_outputs(4558)));
    layer4_outputs(6713) <= layer3_outputs(1399);
    layer4_outputs(6714) <= '1';
    layer4_outputs(6715) <= layer3_outputs(5671);
    layer4_outputs(6716) <= (layer3_outputs(1434)) and not (layer3_outputs(2919));
    layer4_outputs(6717) <= not(layer3_outputs(9397));
    layer4_outputs(6718) <= not((layer3_outputs(4648)) and (layer3_outputs(8455)));
    layer4_outputs(6719) <= layer3_outputs(3888);
    layer4_outputs(6720) <= not(layer3_outputs(2942));
    layer4_outputs(6721) <= (layer3_outputs(2636)) xor (layer3_outputs(1347));
    layer4_outputs(6722) <= (layer3_outputs(7037)) xor (layer3_outputs(3372));
    layer4_outputs(6723) <= not((layer3_outputs(8782)) or (layer3_outputs(465)));
    layer4_outputs(6724) <= not((layer3_outputs(10196)) and (layer3_outputs(403)));
    layer4_outputs(6725) <= not(layer3_outputs(8351));
    layer4_outputs(6726) <= not(layer3_outputs(10203));
    layer4_outputs(6727) <= not(layer3_outputs(4964));
    layer4_outputs(6728) <= layer3_outputs(8413);
    layer4_outputs(6729) <= not(layer3_outputs(776)) or (layer3_outputs(8544));
    layer4_outputs(6730) <= (layer3_outputs(9035)) or (layer3_outputs(7490));
    layer4_outputs(6731) <= (layer3_outputs(6720)) and not (layer3_outputs(4189));
    layer4_outputs(6732) <= layer3_outputs(10097);
    layer4_outputs(6733) <= layer3_outputs(762);
    layer4_outputs(6734) <= layer3_outputs(7289);
    layer4_outputs(6735) <= not(layer3_outputs(915)) or (layer3_outputs(5402));
    layer4_outputs(6736) <= not(layer3_outputs(560)) or (layer3_outputs(1405));
    layer4_outputs(6737) <= layer3_outputs(8048);
    layer4_outputs(6738) <= not((layer3_outputs(9519)) xor (layer3_outputs(9400)));
    layer4_outputs(6739) <= not(layer3_outputs(4558));
    layer4_outputs(6740) <= layer3_outputs(5915);
    layer4_outputs(6741) <= layer3_outputs(4951);
    layer4_outputs(6742) <= layer3_outputs(565);
    layer4_outputs(6743) <= not(layer3_outputs(9347));
    layer4_outputs(6744) <= (layer3_outputs(9099)) and not (layer3_outputs(8056));
    layer4_outputs(6745) <= not(layer3_outputs(7971)) or (layer3_outputs(9743));
    layer4_outputs(6746) <= (layer3_outputs(4216)) and (layer3_outputs(6068));
    layer4_outputs(6747) <= layer3_outputs(8917);
    layer4_outputs(6748) <= (layer3_outputs(7951)) xor (layer3_outputs(6417));
    layer4_outputs(6749) <= layer3_outputs(6624);
    layer4_outputs(6750) <= not(layer3_outputs(8652)) or (layer3_outputs(4642));
    layer4_outputs(6751) <= layer3_outputs(7765);
    layer4_outputs(6752) <= '0';
    layer4_outputs(6753) <= layer3_outputs(9663);
    layer4_outputs(6754) <= (layer3_outputs(9115)) or (layer3_outputs(1644));
    layer4_outputs(6755) <= (layer3_outputs(8810)) xor (layer3_outputs(6687));
    layer4_outputs(6756) <= layer3_outputs(9728);
    layer4_outputs(6757) <= not(layer3_outputs(2384)) or (layer3_outputs(5414));
    layer4_outputs(6758) <= not(layer3_outputs(3012)) or (layer3_outputs(9443));
    layer4_outputs(6759) <= not((layer3_outputs(3164)) and (layer3_outputs(4669)));
    layer4_outputs(6760) <= not(layer3_outputs(83));
    layer4_outputs(6761) <= layer3_outputs(332);
    layer4_outputs(6762) <= not(layer3_outputs(1516));
    layer4_outputs(6763) <= not((layer3_outputs(9950)) xor (layer3_outputs(3719)));
    layer4_outputs(6764) <= layer3_outputs(4985);
    layer4_outputs(6765) <= not(layer3_outputs(992));
    layer4_outputs(6766) <= (layer3_outputs(340)) xor (layer3_outputs(9986));
    layer4_outputs(6767) <= layer3_outputs(8516);
    layer4_outputs(6768) <= not(layer3_outputs(4571));
    layer4_outputs(6769) <= layer3_outputs(6831);
    layer4_outputs(6770) <= (layer3_outputs(1186)) and (layer3_outputs(8066));
    layer4_outputs(6771) <= (layer3_outputs(7851)) or (layer3_outputs(2729));
    layer4_outputs(6772) <= layer3_outputs(7363);
    layer4_outputs(6773) <= layer3_outputs(5601);
    layer4_outputs(6774) <= layer3_outputs(5405);
    layer4_outputs(6775) <= not(layer3_outputs(2225));
    layer4_outputs(6776) <= layer3_outputs(6894);
    layer4_outputs(6777) <= layer3_outputs(3695);
    layer4_outputs(6778) <= not(layer3_outputs(2027));
    layer4_outputs(6779) <= (layer3_outputs(7470)) xor (layer3_outputs(8812));
    layer4_outputs(6780) <= not(layer3_outputs(3419));
    layer4_outputs(6781) <= not(layer3_outputs(3302));
    layer4_outputs(6782) <= not(layer3_outputs(6743));
    layer4_outputs(6783) <= layer3_outputs(3604);
    layer4_outputs(6784) <= layer3_outputs(6379);
    layer4_outputs(6785) <= not((layer3_outputs(5292)) xor (layer3_outputs(9812)));
    layer4_outputs(6786) <= not((layer3_outputs(1666)) and (layer3_outputs(9284)));
    layer4_outputs(6787) <= not(layer3_outputs(3655));
    layer4_outputs(6788) <= '0';
    layer4_outputs(6789) <= not(layer3_outputs(7258));
    layer4_outputs(6790) <= not(layer3_outputs(2230)) or (layer3_outputs(1205));
    layer4_outputs(6791) <= (layer3_outputs(8535)) or (layer3_outputs(5606));
    layer4_outputs(6792) <= (layer3_outputs(431)) and not (layer3_outputs(8304));
    layer4_outputs(6793) <= (layer3_outputs(8681)) or (layer3_outputs(4303));
    layer4_outputs(6794) <= not((layer3_outputs(432)) and (layer3_outputs(4997)));
    layer4_outputs(6795) <= layer3_outputs(324);
    layer4_outputs(6796) <= layer3_outputs(7491);
    layer4_outputs(6797) <= (layer3_outputs(5737)) and (layer3_outputs(5772));
    layer4_outputs(6798) <= not(layer3_outputs(5974));
    layer4_outputs(6799) <= layer3_outputs(9250);
    layer4_outputs(6800) <= (layer3_outputs(8200)) and not (layer3_outputs(2753));
    layer4_outputs(6801) <= layer3_outputs(6464);
    layer4_outputs(6802) <= not((layer3_outputs(10222)) xor (layer3_outputs(6486)));
    layer4_outputs(6803) <= not(layer3_outputs(635));
    layer4_outputs(6804) <= (layer3_outputs(1501)) or (layer3_outputs(7693));
    layer4_outputs(6805) <= not(layer3_outputs(604));
    layer4_outputs(6806) <= (layer3_outputs(2095)) or (layer3_outputs(3104));
    layer4_outputs(6807) <= not(layer3_outputs(8986)) or (layer3_outputs(543));
    layer4_outputs(6808) <= layer3_outputs(7396);
    layer4_outputs(6809) <= (layer3_outputs(6057)) and (layer3_outputs(9064));
    layer4_outputs(6810) <= not(layer3_outputs(3508)) or (layer3_outputs(9713));
    layer4_outputs(6811) <= not(layer3_outputs(9244));
    layer4_outputs(6812) <= not((layer3_outputs(6113)) xor (layer3_outputs(8678)));
    layer4_outputs(6813) <= (layer3_outputs(8005)) and (layer3_outputs(8958));
    layer4_outputs(6814) <= not(layer3_outputs(2158));
    layer4_outputs(6815) <= (layer3_outputs(8058)) and not (layer3_outputs(3659));
    layer4_outputs(6816) <= (layer3_outputs(3856)) xor (layer3_outputs(6762));
    layer4_outputs(6817) <= not((layer3_outputs(3568)) or (layer3_outputs(1520)));
    layer4_outputs(6818) <= (layer3_outputs(4407)) and not (layer3_outputs(3816));
    layer4_outputs(6819) <= layer3_outputs(8599);
    layer4_outputs(6820) <= layer3_outputs(6866);
    layer4_outputs(6821) <= not(layer3_outputs(9315)) or (layer3_outputs(3717));
    layer4_outputs(6822) <= (layer3_outputs(4150)) and (layer3_outputs(7392));
    layer4_outputs(6823) <= (layer3_outputs(6417)) and not (layer3_outputs(753));
    layer4_outputs(6824) <= not((layer3_outputs(9702)) xor (layer3_outputs(5555)));
    layer4_outputs(6825) <= not(layer3_outputs(5056));
    layer4_outputs(6826) <= layer3_outputs(3776);
    layer4_outputs(6827) <= (layer3_outputs(9251)) and not (layer3_outputs(4596));
    layer4_outputs(6828) <= (layer3_outputs(10175)) and not (layer3_outputs(4677));
    layer4_outputs(6829) <= layer3_outputs(8275);
    layer4_outputs(6830) <= not(layer3_outputs(2172));
    layer4_outputs(6831) <= not(layer3_outputs(4429));
    layer4_outputs(6832) <= not(layer3_outputs(7529));
    layer4_outputs(6833) <= (layer3_outputs(1589)) and not (layer3_outputs(2835));
    layer4_outputs(6834) <= layer3_outputs(6664);
    layer4_outputs(6835) <= (layer3_outputs(6406)) xor (layer3_outputs(6671));
    layer4_outputs(6836) <= (layer3_outputs(9561)) xor (layer3_outputs(9509));
    layer4_outputs(6837) <= not(layer3_outputs(10021));
    layer4_outputs(6838) <= not(layer3_outputs(4919));
    layer4_outputs(6839) <= not((layer3_outputs(5717)) xor (layer3_outputs(4213)));
    layer4_outputs(6840) <= not((layer3_outputs(1014)) xor (layer3_outputs(8085)));
    layer4_outputs(6841) <= not(layer3_outputs(7325));
    layer4_outputs(6842) <= not((layer3_outputs(2079)) xor (layer3_outputs(6434)));
    layer4_outputs(6843) <= (layer3_outputs(2913)) and (layer3_outputs(5513));
    layer4_outputs(6844) <= not(layer3_outputs(4417));
    layer4_outputs(6845) <= not(layer3_outputs(7589));
    layer4_outputs(6846) <= not(layer3_outputs(5821));
    layer4_outputs(6847) <= (layer3_outputs(8093)) and (layer3_outputs(3734));
    layer4_outputs(6848) <= not(layer3_outputs(6564));
    layer4_outputs(6849) <= not(layer3_outputs(4918));
    layer4_outputs(6850) <= (layer3_outputs(538)) and (layer3_outputs(9114));
    layer4_outputs(6851) <= not((layer3_outputs(6989)) and (layer3_outputs(9535)));
    layer4_outputs(6852) <= not(layer3_outputs(3344));
    layer4_outputs(6853) <= not(layer3_outputs(6848));
    layer4_outputs(6854) <= not(layer3_outputs(1449));
    layer4_outputs(6855) <= layer3_outputs(532);
    layer4_outputs(6856) <= not(layer3_outputs(8608));
    layer4_outputs(6857) <= not((layer3_outputs(9063)) or (layer3_outputs(3780)));
    layer4_outputs(6858) <= not(layer3_outputs(1162));
    layer4_outputs(6859) <= not((layer3_outputs(8737)) xor (layer3_outputs(6465)));
    layer4_outputs(6860) <= (layer3_outputs(5602)) and not (layer3_outputs(4623));
    layer4_outputs(6861) <= layer3_outputs(3596);
    layer4_outputs(6862) <= (layer3_outputs(1091)) or (layer3_outputs(3113));
    layer4_outputs(6863) <= not(layer3_outputs(7343)) or (layer3_outputs(4104));
    layer4_outputs(6864) <= layer3_outputs(9915);
    layer4_outputs(6865) <= (layer3_outputs(2572)) or (layer3_outputs(9196));
    layer4_outputs(6866) <= not(layer3_outputs(2912)) or (layer3_outputs(4270));
    layer4_outputs(6867) <= (layer3_outputs(4983)) or (layer3_outputs(7770));
    layer4_outputs(6868) <= layer3_outputs(7995);
    layer4_outputs(6869) <= not(layer3_outputs(6599)) or (layer3_outputs(5944));
    layer4_outputs(6870) <= not(layer3_outputs(10128));
    layer4_outputs(6871) <= layer3_outputs(3763);
    layer4_outputs(6872) <= (layer3_outputs(7170)) and not (layer3_outputs(7329));
    layer4_outputs(6873) <= not((layer3_outputs(3969)) xor (layer3_outputs(5264)));
    layer4_outputs(6874) <= (layer3_outputs(2744)) xor (layer3_outputs(4299));
    layer4_outputs(6875) <= not(layer3_outputs(4732)) or (layer3_outputs(10077));
    layer4_outputs(6876) <= not(layer3_outputs(1615));
    layer4_outputs(6877) <= (layer3_outputs(9408)) and (layer3_outputs(4273));
    layer4_outputs(6878) <= not(layer3_outputs(282));
    layer4_outputs(6879) <= (layer3_outputs(9241)) and not (layer3_outputs(597));
    layer4_outputs(6880) <= not(layer3_outputs(2936));
    layer4_outputs(6881) <= (layer3_outputs(4721)) xor (layer3_outputs(8133));
    layer4_outputs(6882) <= (layer3_outputs(8790)) and not (layer3_outputs(1739));
    layer4_outputs(6883) <= not((layer3_outputs(7915)) xor (layer3_outputs(330)));
    layer4_outputs(6884) <= not(layer3_outputs(5770));
    layer4_outputs(6885) <= (layer3_outputs(973)) and (layer3_outputs(6321));
    layer4_outputs(6886) <= layer3_outputs(8707);
    layer4_outputs(6887) <= layer3_outputs(8260);
    layer4_outputs(6888) <= (layer3_outputs(7024)) and not (layer3_outputs(5161));
    layer4_outputs(6889) <= (layer3_outputs(9748)) xor (layer3_outputs(2184));
    layer4_outputs(6890) <= layer3_outputs(1232);
    layer4_outputs(6891) <= not(layer3_outputs(2650));
    layer4_outputs(6892) <= not(layer3_outputs(8312));
    layer4_outputs(6893) <= not(layer3_outputs(936));
    layer4_outputs(6894) <= layer3_outputs(2690);
    layer4_outputs(6895) <= not(layer3_outputs(2937));
    layer4_outputs(6896) <= layer3_outputs(283);
    layer4_outputs(6897) <= (layer3_outputs(2466)) and not (layer3_outputs(4976));
    layer4_outputs(6898) <= not(layer3_outputs(6794)) or (layer3_outputs(7685));
    layer4_outputs(6899) <= (layer3_outputs(109)) xor (layer3_outputs(394));
    layer4_outputs(6900) <= layer3_outputs(3111);
    layer4_outputs(6901) <= not(layer3_outputs(7129));
    layer4_outputs(6902) <= layer3_outputs(7584);
    layer4_outputs(6903) <= layer3_outputs(7923);
    layer4_outputs(6904) <= not(layer3_outputs(2179)) or (layer3_outputs(9095));
    layer4_outputs(6905) <= not(layer3_outputs(1950));
    layer4_outputs(6906) <= not(layer3_outputs(2486));
    layer4_outputs(6907) <= not(layer3_outputs(3482));
    layer4_outputs(6908) <= layer3_outputs(2933);
    layer4_outputs(6909) <= not(layer3_outputs(2836));
    layer4_outputs(6910) <= (layer3_outputs(7290)) xor (layer3_outputs(8984));
    layer4_outputs(6911) <= not(layer3_outputs(7947)) or (layer3_outputs(6083));
    layer4_outputs(6912) <= not((layer3_outputs(586)) xor (layer3_outputs(5411)));
    layer4_outputs(6913) <= not(layer3_outputs(5800));
    layer4_outputs(6914) <= (layer3_outputs(1807)) and not (layer3_outputs(5328));
    layer4_outputs(6915) <= not(layer3_outputs(4806));
    layer4_outputs(6916) <= not(layer3_outputs(7099));
    layer4_outputs(6917) <= (layer3_outputs(10219)) and not (layer3_outputs(5143));
    layer4_outputs(6918) <= layer3_outputs(4354);
    layer4_outputs(6919) <= (layer3_outputs(5831)) or (layer3_outputs(5474));
    layer4_outputs(6920) <= (layer3_outputs(6695)) xor (layer3_outputs(250));
    layer4_outputs(6921) <= layer3_outputs(2831);
    layer4_outputs(6922) <= not(layer3_outputs(5525));
    layer4_outputs(6923) <= layer3_outputs(6286);
    layer4_outputs(6924) <= not(layer3_outputs(3187));
    layer4_outputs(6925) <= not(layer3_outputs(6467));
    layer4_outputs(6926) <= not(layer3_outputs(8653));
    layer4_outputs(6927) <= layer3_outputs(2192);
    layer4_outputs(6928) <= not(layer3_outputs(1960)) or (layer3_outputs(496));
    layer4_outputs(6929) <= not(layer3_outputs(7133));
    layer4_outputs(6930) <= layer3_outputs(3709);
    layer4_outputs(6931) <= layer3_outputs(9268);
    layer4_outputs(6932) <= not((layer3_outputs(10104)) xor (layer3_outputs(203)));
    layer4_outputs(6933) <= (layer3_outputs(4702)) xor (layer3_outputs(8136));
    layer4_outputs(6934) <= layer3_outputs(5452);
    layer4_outputs(6935) <= (layer3_outputs(1458)) and not (layer3_outputs(6621));
    layer4_outputs(6936) <= not((layer3_outputs(1103)) or (layer3_outputs(5560)));
    layer4_outputs(6937) <= not(layer3_outputs(6559)) or (layer3_outputs(8284));
    layer4_outputs(6938) <= not((layer3_outputs(3408)) xor (layer3_outputs(353)));
    layer4_outputs(6939) <= (layer3_outputs(5291)) and (layer3_outputs(6364));
    layer4_outputs(6940) <= (layer3_outputs(244)) and not (layer3_outputs(1893));
    layer4_outputs(6941) <= (layer3_outputs(8997)) xor (layer3_outputs(1207));
    layer4_outputs(6942) <= not(layer3_outputs(10008)) or (layer3_outputs(9127));
    layer4_outputs(6943) <= layer3_outputs(9296);
    layer4_outputs(6944) <= not(layer3_outputs(10044));
    layer4_outputs(6945) <= not(layer3_outputs(6792)) or (layer3_outputs(5797));
    layer4_outputs(6946) <= layer3_outputs(7123);
    layer4_outputs(6947) <= layer3_outputs(6561);
    layer4_outputs(6948) <= layer3_outputs(1145);
    layer4_outputs(6949) <= not(layer3_outputs(7039));
    layer4_outputs(6950) <= (layer3_outputs(6188)) and not (layer3_outputs(8889));
    layer4_outputs(6951) <= layer3_outputs(9414);
    layer4_outputs(6952) <= not(layer3_outputs(3340));
    layer4_outputs(6953) <= not((layer3_outputs(3273)) and (layer3_outputs(129)));
    layer4_outputs(6954) <= layer3_outputs(8264);
    layer4_outputs(6955) <= (layer3_outputs(8333)) and not (layer3_outputs(1990));
    layer4_outputs(6956) <= not(layer3_outputs(3488));
    layer4_outputs(6957) <= layer3_outputs(2839);
    layer4_outputs(6958) <= not((layer3_outputs(993)) or (layer3_outputs(5116)));
    layer4_outputs(6959) <= not(layer3_outputs(2908));
    layer4_outputs(6960) <= (layer3_outputs(3304)) and (layer3_outputs(5340));
    layer4_outputs(6961) <= (layer3_outputs(8925)) xor (layer3_outputs(1308));
    layer4_outputs(6962) <= not(layer3_outputs(2164));
    layer4_outputs(6963) <= not(layer3_outputs(4701));
    layer4_outputs(6964) <= layer3_outputs(6151);
    layer4_outputs(6965) <= not((layer3_outputs(3966)) or (layer3_outputs(888)));
    layer4_outputs(6966) <= (layer3_outputs(6248)) and not (layer3_outputs(8486));
    layer4_outputs(6967) <= not(layer3_outputs(3619));
    layer4_outputs(6968) <= (layer3_outputs(5240)) or (layer3_outputs(2104));
    layer4_outputs(6969) <= not((layer3_outputs(5949)) or (layer3_outputs(5367)));
    layer4_outputs(6970) <= not(layer3_outputs(10174));
    layer4_outputs(6971) <= not(layer3_outputs(2339)) or (layer3_outputs(4966));
    layer4_outputs(6972) <= not(layer3_outputs(7393));
    layer4_outputs(6973) <= layer3_outputs(9145);
    layer4_outputs(6974) <= not(layer3_outputs(8074));
    layer4_outputs(6975) <= layer3_outputs(9386);
    layer4_outputs(6976) <= layer3_outputs(7336);
    layer4_outputs(6977) <= not(layer3_outputs(9833));
    layer4_outputs(6978) <= not(layer3_outputs(3491));
    layer4_outputs(6979) <= layer3_outputs(4368);
    layer4_outputs(6980) <= not(layer3_outputs(1069));
    layer4_outputs(6981) <= not(layer3_outputs(8844));
    layer4_outputs(6982) <= (layer3_outputs(9305)) and not (layer3_outputs(8050));
    layer4_outputs(6983) <= (layer3_outputs(74)) xor (layer3_outputs(3645));
    layer4_outputs(6984) <= (layer3_outputs(3657)) and (layer3_outputs(9730));
    layer4_outputs(6985) <= not((layer3_outputs(4207)) xor (layer3_outputs(8938)));
    layer4_outputs(6986) <= layer3_outputs(7450);
    layer4_outputs(6987) <= not(layer3_outputs(2960));
    layer4_outputs(6988) <= layer3_outputs(2960);
    layer4_outputs(6989) <= not((layer3_outputs(1290)) and (layer3_outputs(3631)));
    layer4_outputs(6990) <= (layer3_outputs(3078)) and not (layer3_outputs(5322));
    layer4_outputs(6991) <= layer3_outputs(9583);
    layer4_outputs(6992) <= (layer3_outputs(5408)) and not (layer3_outputs(8342));
    layer4_outputs(6993) <= (layer3_outputs(178)) xor (layer3_outputs(6351));
    layer4_outputs(6994) <= layer3_outputs(4371);
    layer4_outputs(6995) <= (layer3_outputs(1695)) and not (layer3_outputs(9223));
    layer4_outputs(6996) <= not(layer3_outputs(8417));
    layer4_outputs(6997) <= not((layer3_outputs(8210)) or (layer3_outputs(8311)));
    layer4_outputs(6998) <= not(layer3_outputs(707));
    layer4_outputs(6999) <= layer3_outputs(4209);
    layer4_outputs(7000) <= not((layer3_outputs(5659)) or (layer3_outputs(5897)));
    layer4_outputs(7001) <= not(layer3_outputs(4045)) or (layer3_outputs(6023));
    layer4_outputs(7002) <= layer3_outputs(5658);
    layer4_outputs(7003) <= not(layer3_outputs(9013));
    layer4_outputs(7004) <= not(layer3_outputs(3823));
    layer4_outputs(7005) <= layer3_outputs(7405);
    layer4_outputs(7006) <= layer3_outputs(59);
    layer4_outputs(7007) <= (layer3_outputs(3418)) and not (layer3_outputs(9157));
    layer4_outputs(7008) <= (layer3_outputs(2872)) and not (layer3_outputs(5750));
    layer4_outputs(7009) <= layer3_outputs(6112);
    layer4_outputs(7010) <= layer3_outputs(7080);
    layer4_outputs(7011) <= (layer3_outputs(9102)) xor (layer3_outputs(5016));
    layer4_outputs(7012) <= not(layer3_outputs(3311));
    layer4_outputs(7013) <= not(layer3_outputs(2538));
    layer4_outputs(7014) <= not(layer3_outputs(2647)) or (layer3_outputs(9818));
    layer4_outputs(7015) <= not(layer3_outputs(10111));
    layer4_outputs(7016) <= (layer3_outputs(1178)) xor (layer3_outputs(3129));
    layer4_outputs(7017) <= layer3_outputs(1968);
    layer4_outputs(7018) <= layer3_outputs(6423);
    layer4_outputs(7019) <= not(layer3_outputs(2495));
    layer4_outputs(7020) <= (layer3_outputs(725)) xor (layer3_outputs(4466));
    layer4_outputs(7021) <= not(layer3_outputs(6037));
    layer4_outputs(7022) <= not(layer3_outputs(2927));
    layer4_outputs(7023) <= not((layer3_outputs(6531)) xor (layer3_outputs(962)));
    layer4_outputs(7024) <= not(layer3_outputs(3383));
    layer4_outputs(7025) <= not(layer3_outputs(6481));
    layer4_outputs(7026) <= not(layer3_outputs(2491));
    layer4_outputs(7027) <= not((layer3_outputs(4699)) xor (layer3_outputs(9505)));
    layer4_outputs(7028) <= not((layer3_outputs(8662)) and (layer3_outputs(2102)));
    layer4_outputs(7029) <= not(layer3_outputs(9440));
    layer4_outputs(7030) <= layer3_outputs(8686);
    layer4_outputs(7031) <= (layer3_outputs(8718)) xor (layer3_outputs(3595));
    layer4_outputs(7032) <= not((layer3_outputs(2646)) or (layer3_outputs(9975)));
    layer4_outputs(7033) <= (layer3_outputs(4554)) xor (layer3_outputs(8676));
    layer4_outputs(7034) <= not(layer3_outputs(254));
    layer4_outputs(7035) <= layer3_outputs(4562);
    layer4_outputs(7036) <= layer3_outputs(8562);
    layer4_outputs(7037) <= not((layer3_outputs(4245)) xor (layer3_outputs(8785)));
    layer4_outputs(7038) <= layer3_outputs(8302);
    layer4_outputs(7039) <= not(layer3_outputs(4110));
    layer4_outputs(7040) <= not(layer3_outputs(7051)) or (layer3_outputs(9023));
    layer4_outputs(7041) <= (layer3_outputs(8704)) xor (layer3_outputs(4050));
    layer4_outputs(7042) <= layer3_outputs(2537);
    layer4_outputs(7043) <= layer3_outputs(465);
    layer4_outputs(7044) <= not((layer3_outputs(8022)) and (layer3_outputs(9516)));
    layer4_outputs(7045) <= not((layer3_outputs(2316)) and (layer3_outputs(2501)));
    layer4_outputs(7046) <= '1';
    layer4_outputs(7047) <= not(layer3_outputs(9125));
    layer4_outputs(7048) <= not(layer3_outputs(8483)) or (layer3_outputs(9053));
    layer4_outputs(7049) <= layer3_outputs(7348);
    layer4_outputs(7050) <= layer3_outputs(188);
    layer4_outputs(7051) <= not(layer3_outputs(1294));
    layer4_outputs(7052) <= not((layer3_outputs(1001)) and (layer3_outputs(438)));
    layer4_outputs(7053) <= layer3_outputs(5567);
    layer4_outputs(7054) <= layer3_outputs(2361);
    layer4_outputs(7055) <= not(layer3_outputs(3858));
    layer4_outputs(7056) <= (layer3_outputs(6627)) and not (layer3_outputs(3200));
    layer4_outputs(7057) <= (layer3_outputs(1067)) and not (layer3_outputs(3777));
    layer4_outputs(7058) <= layer3_outputs(7256);
    layer4_outputs(7059) <= not(layer3_outputs(6643)) or (layer3_outputs(3122));
    layer4_outputs(7060) <= not(layer3_outputs(1039));
    layer4_outputs(7061) <= not(layer3_outputs(6151));
    layer4_outputs(7062) <= layer3_outputs(7163);
    layer4_outputs(7063) <= not((layer3_outputs(1833)) and (layer3_outputs(8766)));
    layer4_outputs(7064) <= not(layer3_outputs(592));
    layer4_outputs(7065) <= (layer3_outputs(2137)) and not (layer3_outputs(2202));
    layer4_outputs(7066) <= '1';
    layer4_outputs(7067) <= not(layer3_outputs(1250));
    layer4_outputs(7068) <= layer3_outputs(9299);
    layer4_outputs(7069) <= not((layer3_outputs(406)) xor (layer3_outputs(7425)));
    layer4_outputs(7070) <= not((layer3_outputs(3923)) and (layer3_outputs(1476)));
    layer4_outputs(7071) <= (layer3_outputs(7639)) and not (layer3_outputs(4649));
    layer4_outputs(7072) <= not((layer3_outputs(3187)) xor (layer3_outputs(9886)));
    layer4_outputs(7073) <= not(layer3_outputs(3866));
    layer4_outputs(7074) <= not(layer3_outputs(3592));
    layer4_outputs(7075) <= (layer3_outputs(1863)) and (layer3_outputs(3398));
    layer4_outputs(7076) <= not(layer3_outputs(4143));
    layer4_outputs(7077) <= layer3_outputs(1000);
    layer4_outputs(7078) <= (layer3_outputs(6210)) xor (layer3_outputs(2054));
    layer4_outputs(7079) <= layer3_outputs(9590);
    layer4_outputs(7080) <= not(layer3_outputs(7410));
    layer4_outputs(7081) <= layer3_outputs(2927);
    layer4_outputs(7082) <= layer3_outputs(1455);
    layer4_outputs(7083) <= layer3_outputs(5679);
    layer4_outputs(7084) <= not(layer3_outputs(7474));
    layer4_outputs(7085) <= layer3_outputs(3910);
    layer4_outputs(7086) <= layer3_outputs(2170);
    layer4_outputs(7087) <= not((layer3_outputs(243)) and (layer3_outputs(2449)));
    layer4_outputs(7088) <= not((layer3_outputs(3742)) xor (layer3_outputs(677)));
    layer4_outputs(7089) <= layer3_outputs(8168);
    layer4_outputs(7090) <= (layer3_outputs(3637)) or (layer3_outputs(913));
    layer4_outputs(7091) <= '0';
    layer4_outputs(7092) <= (layer3_outputs(9217)) or (layer3_outputs(8981));
    layer4_outputs(7093) <= not(layer3_outputs(110));
    layer4_outputs(7094) <= layer3_outputs(968);
    layer4_outputs(7095) <= (layer3_outputs(8921)) or (layer3_outputs(2149));
    layer4_outputs(7096) <= not(layer3_outputs(5091));
    layer4_outputs(7097) <= not(layer3_outputs(4373));
    layer4_outputs(7098) <= not(layer3_outputs(4700));
    layer4_outputs(7099) <= layer3_outputs(863);
    layer4_outputs(7100) <= layer3_outputs(5164);
    layer4_outputs(7101) <= not((layer3_outputs(8303)) or (layer3_outputs(4541)));
    layer4_outputs(7102) <= not(layer3_outputs(8455));
    layer4_outputs(7103) <= not(layer3_outputs(5864));
    layer4_outputs(7104) <= (layer3_outputs(5086)) and not (layer3_outputs(6279));
    layer4_outputs(7105) <= not(layer3_outputs(3056));
    layer4_outputs(7106) <= not(layer3_outputs(5490)) or (layer3_outputs(8520));
    layer4_outputs(7107) <= (layer3_outputs(4540)) and (layer3_outputs(3938));
    layer4_outputs(7108) <= layer3_outputs(4083);
    layer4_outputs(7109) <= (layer3_outputs(75)) and not (layer3_outputs(3204));
    layer4_outputs(7110) <= layer3_outputs(3706);
    layer4_outputs(7111) <= layer3_outputs(7379);
    layer4_outputs(7112) <= not((layer3_outputs(8570)) xor (layer3_outputs(7921)));
    layer4_outputs(7113) <= not(layer3_outputs(6214));
    layer4_outputs(7114) <= layer3_outputs(9441);
    layer4_outputs(7115) <= not((layer3_outputs(6192)) and (layer3_outputs(2542)));
    layer4_outputs(7116) <= layer3_outputs(2421);
    layer4_outputs(7117) <= not(layer3_outputs(5314));
    layer4_outputs(7118) <= not(layer3_outputs(4440));
    layer4_outputs(7119) <= not(layer3_outputs(2849));
    layer4_outputs(7120) <= layer3_outputs(9821);
    layer4_outputs(7121) <= not(layer3_outputs(2631));
    layer4_outputs(7122) <= not(layer3_outputs(739));
    layer4_outputs(7123) <= not(layer3_outputs(1388));
    layer4_outputs(7124) <= '1';
    layer4_outputs(7125) <= not(layer3_outputs(4499));
    layer4_outputs(7126) <= (layer3_outputs(8442)) and not (layer3_outputs(8654));
    layer4_outputs(7127) <= layer3_outputs(9322);
    layer4_outputs(7128) <= (layer3_outputs(2484)) and not (layer3_outputs(9311));
    layer4_outputs(7129) <= not(layer3_outputs(2198));
    layer4_outputs(7130) <= not(layer3_outputs(4862)) or (layer3_outputs(9644));
    layer4_outputs(7131) <= not((layer3_outputs(4670)) xor (layer3_outputs(3661)));
    layer4_outputs(7132) <= not(layer3_outputs(5125)) or (layer3_outputs(5495));
    layer4_outputs(7133) <= layer3_outputs(5227);
    layer4_outputs(7134) <= not(layer3_outputs(3864));
    layer4_outputs(7135) <= (layer3_outputs(6990)) xor (layer3_outputs(2675));
    layer4_outputs(7136) <= layer3_outputs(3147);
    layer4_outputs(7137) <= (layer3_outputs(5736)) or (layer3_outputs(343));
    layer4_outputs(7138) <= (layer3_outputs(6421)) xor (layer3_outputs(7871));
    layer4_outputs(7139) <= not((layer3_outputs(8285)) xor (layer3_outputs(4629)));
    layer4_outputs(7140) <= layer3_outputs(2120);
    layer4_outputs(7141) <= layer3_outputs(9913);
    layer4_outputs(7142) <= layer3_outputs(1099);
    layer4_outputs(7143) <= not((layer3_outputs(5346)) xor (layer3_outputs(8705)));
    layer4_outputs(7144) <= layer3_outputs(3480);
    layer4_outputs(7145) <= (layer3_outputs(9132)) xor (layer3_outputs(9512));
    layer4_outputs(7146) <= not((layer3_outputs(1495)) or (layer3_outputs(5159)));
    layer4_outputs(7147) <= layer3_outputs(9223);
    layer4_outputs(7148) <= not(layer3_outputs(1748));
    layer4_outputs(7149) <= not(layer3_outputs(5759));
    layer4_outputs(7150) <= not(layer3_outputs(7347)) or (layer3_outputs(3096));
    layer4_outputs(7151) <= not(layer3_outputs(5617));
    layer4_outputs(7152) <= layer3_outputs(8265);
    layer4_outputs(7153) <= (layer3_outputs(2204)) and not (layer3_outputs(3895));
    layer4_outputs(7154) <= not(layer3_outputs(5226));
    layer4_outputs(7155) <= not(layer3_outputs(8531)) or (layer3_outputs(9830));
    layer4_outputs(7156) <= (layer3_outputs(4178)) xor (layer3_outputs(35));
    layer4_outputs(7157) <= not(layer3_outputs(2898));
    layer4_outputs(7158) <= not((layer3_outputs(5146)) or (layer3_outputs(9192)));
    layer4_outputs(7159) <= not(layer3_outputs(1555));
    layer4_outputs(7160) <= not(layer3_outputs(4446));
    layer4_outputs(7161) <= layer3_outputs(641);
    layer4_outputs(7162) <= not(layer3_outputs(8966)) or (layer3_outputs(6745));
    layer4_outputs(7163) <= not(layer3_outputs(7058));
    layer4_outputs(7164) <= not(layer3_outputs(1342));
    layer4_outputs(7165) <= layer3_outputs(6739);
    layer4_outputs(7166) <= (layer3_outputs(6624)) or (layer3_outputs(9118));
    layer4_outputs(7167) <= layer3_outputs(8556);
    layer4_outputs(7168) <= layer3_outputs(3487);
    layer4_outputs(7169) <= not((layer3_outputs(6982)) xor (layer3_outputs(8200)));
    layer4_outputs(7170) <= layer3_outputs(9977);
    layer4_outputs(7171) <= layer3_outputs(1636);
    layer4_outputs(7172) <= not(layer3_outputs(2148));
    layer4_outputs(7173) <= not(layer3_outputs(1295));
    layer4_outputs(7174) <= not(layer3_outputs(7102));
    layer4_outputs(7175) <= layer3_outputs(4610);
    layer4_outputs(7176) <= layer3_outputs(6284);
    layer4_outputs(7177) <= layer3_outputs(5069);
    layer4_outputs(7178) <= (layer3_outputs(5120)) xor (layer3_outputs(4722));
    layer4_outputs(7179) <= not(layer3_outputs(9682));
    layer4_outputs(7180) <= (layer3_outputs(6339)) xor (layer3_outputs(4982));
    layer4_outputs(7181) <= (layer3_outputs(1813)) and not (layer3_outputs(3668));
    layer4_outputs(7182) <= layer3_outputs(4572);
    layer4_outputs(7183) <= not(layer3_outputs(2351));
    layer4_outputs(7184) <= not((layer3_outputs(2821)) or (layer3_outputs(771)));
    layer4_outputs(7185) <= not(layer3_outputs(5119)) or (layer3_outputs(1023));
    layer4_outputs(7186) <= not((layer3_outputs(3359)) or (layer3_outputs(9930)));
    layer4_outputs(7187) <= not(layer3_outputs(2360));
    layer4_outputs(7188) <= not(layer3_outputs(8414)) or (layer3_outputs(9919));
    layer4_outputs(7189) <= not(layer3_outputs(7401));
    layer4_outputs(7190) <= not(layer3_outputs(534)) or (layer3_outputs(5842));
    layer4_outputs(7191) <= layer3_outputs(249);
    layer4_outputs(7192) <= layer3_outputs(3204);
    layer4_outputs(7193) <= not(layer3_outputs(8791));
    layer4_outputs(7194) <= (layer3_outputs(3100)) and (layer3_outputs(9879));
    layer4_outputs(7195) <= layer3_outputs(8325);
    layer4_outputs(7196) <= layer3_outputs(6940);
    layer4_outputs(7197) <= (layer3_outputs(7009)) xor (layer3_outputs(8812));
    layer4_outputs(7198) <= layer3_outputs(8069);
    layer4_outputs(7199) <= layer3_outputs(8475);
    layer4_outputs(7200) <= not(layer3_outputs(2511)) or (layer3_outputs(5611));
    layer4_outputs(7201) <= not(layer3_outputs(7541)) or (layer3_outputs(5391));
    layer4_outputs(7202) <= not(layer3_outputs(711));
    layer4_outputs(7203) <= not(layer3_outputs(1118)) or (layer3_outputs(5058));
    layer4_outputs(7204) <= layer3_outputs(10017);
    layer4_outputs(7205) <= not(layer3_outputs(9197));
    layer4_outputs(7206) <= (layer3_outputs(5041)) and (layer3_outputs(3648));
    layer4_outputs(7207) <= not(layer3_outputs(5531)) or (layer3_outputs(7011));
    layer4_outputs(7208) <= not(layer3_outputs(5462));
    layer4_outputs(7209) <= not(layer3_outputs(424)) or (layer3_outputs(6373));
    layer4_outputs(7210) <= (layer3_outputs(884)) xor (layer3_outputs(8386));
    layer4_outputs(7211) <= (layer3_outputs(8920)) xor (layer3_outputs(6976));
    layer4_outputs(7212) <= not(layer3_outputs(9849));
    layer4_outputs(7213) <= not(layer3_outputs(9482));
    layer4_outputs(7214) <= not((layer3_outputs(6317)) or (layer3_outputs(4575)));
    layer4_outputs(7215) <= layer3_outputs(8469);
    layer4_outputs(7216) <= layer3_outputs(272);
    layer4_outputs(7217) <= '0';
    layer4_outputs(7218) <= (layer3_outputs(7333)) and (layer3_outputs(1932));
    layer4_outputs(7219) <= not((layer3_outputs(1281)) xor (layer3_outputs(1007)));
    layer4_outputs(7220) <= not((layer3_outputs(722)) xor (layer3_outputs(242)));
    layer4_outputs(7221) <= not(layer3_outputs(9266));
    layer4_outputs(7222) <= not(layer3_outputs(3168));
    layer4_outputs(7223) <= (layer3_outputs(6283)) and not (layer3_outputs(2541));
    layer4_outputs(7224) <= (layer3_outputs(4083)) xor (layer3_outputs(2794));
    layer4_outputs(7225) <= not(layer3_outputs(2915)) or (layer3_outputs(2450));
    layer4_outputs(7226) <= not(layer3_outputs(4268));
    layer4_outputs(7227) <= (layer3_outputs(8007)) xor (layer3_outputs(3072));
    layer4_outputs(7228) <= not(layer3_outputs(1912));
    layer4_outputs(7229) <= layer3_outputs(967);
    layer4_outputs(7230) <= not(layer3_outputs(5380));
    layer4_outputs(7231) <= layer3_outputs(2475);
    layer4_outputs(7232) <= not(layer3_outputs(1577));
    layer4_outputs(7233) <= layer3_outputs(3099);
    layer4_outputs(7234) <= layer3_outputs(7565);
    layer4_outputs(7235) <= not(layer3_outputs(2558));
    layer4_outputs(7236) <= not(layer3_outputs(2319)) or (layer3_outputs(3293));
    layer4_outputs(7237) <= not(layer3_outputs(9734)) or (layer3_outputs(8149));
    layer4_outputs(7238) <= (layer3_outputs(9289)) xor (layer3_outputs(3247));
    layer4_outputs(7239) <= not(layer3_outputs(9379)) or (layer3_outputs(6257));
    layer4_outputs(7240) <= not((layer3_outputs(271)) xor (layer3_outputs(4348)));
    layer4_outputs(7241) <= layer3_outputs(4962);
    layer4_outputs(7242) <= not((layer3_outputs(5631)) xor (layer3_outputs(7511)));
    layer4_outputs(7243) <= not(layer3_outputs(4624));
    layer4_outputs(7244) <= not(layer3_outputs(2114));
    layer4_outputs(7245) <= not((layer3_outputs(307)) xor (layer3_outputs(8305)));
    layer4_outputs(7246) <= not(layer3_outputs(865)) or (layer3_outputs(926));
    layer4_outputs(7247) <= (layer3_outputs(3844)) and not (layer3_outputs(9691));
    layer4_outputs(7248) <= not((layer3_outputs(3320)) xor (layer3_outputs(7589)));
    layer4_outputs(7249) <= (layer3_outputs(2316)) or (layer3_outputs(2407));
    layer4_outputs(7250) <= not((layer3_outputs(476)) xor (layer3_outputs(2088)));
    layer4_outputs(7251) <= layer3_outputs(8585);
    layer4_outputs(7252) <= layer3_outputs(542);
    layer4_outputs(7253) <= (layer3_outputs(7657)) xor (layer3_outputs(4030));
    layer4_outputs(7254) <= not(layer3_outputs(8458));
    layer4_outputs(7255) <= not(layer3_outputs(395)) or (layer3_outputs(9653));
    layer4_outputs(7256) <= not(layer3_outputs(478));
    layer4_outputs(7257) <= layer3_outputs(6181);
    layer4_outputs(7258) <= not((layer3_outputs(9187)) and (layer3_outputs(8613)));
    layer4_outputs(7259) <= not((layer3_outputs(567)) xor (layer3_outputs(7463)));
    layer4_outputs(7260) <= layer3_outputs(2894);
    layer4_outputs(7261) <= layer3_outputs(7862);
    layer4_outputs(7262) <= not(layer3_outputs(1519)) or (layer3_outputs(6569));
    layer4_outputs(7263) <= not(layer3_outputs(4613));
    layer4_outputs(7264) <= (layer3_outputs(7078)) and not (layer3_outputs(8087));
    layer4_outputs(7265) <= '0';
    layer4_outputs(7266) <= layer3_outputs(1214);
    layer4_outputs(7267) <= (layer3_outputs(2964)) and (layer3_outputs(2905));
    layer4_outputs(7268) <= not(layer3_outputs(9140));
    layer4_outputs(7269) <= not(layer3_outputs(6940));
    layer4_outputs(7270) <= not((layer3_outputs(3007)) xor (layer3_outputs(1559)));
    layer4_outputs(7271) <= not(layer3_outputs(755));
    layer4_outputs(7272) <= not((layer3_outputs(5856)) and (layer3_outputs(3608)));
    layer4_outputs(7273) <= not(layer3_outputs(4861));
    layer4_outputs(7274) <= (layer3_outputs(3969)) and (layer3_outputs(4863));
    layer4_outputs(7275) <= (layer3_outputs(871)) xor (layer3_outputs(4420));
    layer4_outputs(7276) <= (layer3_outputs(2317)) and (layer3_outputs(7718));
    layer4_outputs(7277) <= layer3_outputs(4332);
    layer4_outputs(7278) <= (layer3_outputs(6801)) xor (layer3_outputs(6142));
    layer4_outputs(7279) <= not(layer3_outputs(5378)) or (layer3_outputs(1152));
    layer4_outputs(7280) <= not(layer3_outputs(6845));
    layer4_outputs(7281) <= not((layer3_outputs(8706)) xor (layer3_outputs(9968)));
    layer4_outputs(7282) <= layer3_outputs(3662);
    layer4_outputs(7283) <= not(layer3_outputs(9985));
    layer4_outputs(7284) <= layer3_outputs(1180);
    layer4_outputs(7285) <= not(layer3_outputs(590)) or (layer3_outputs(3853));
    layer4_outputs(7286) <= layer3_outputs(4235);
    layer4_outputs(7287) <= '1';
    layer4_outputs(7288) <= (layer3_outputs(1163)) xor (layer3_outputs(8343));
    layer4_outputs(7289) <= not(layer3_outputs(5889));
    layer4_outputs(7290) <= not(layer3_outputs(1789));
    layer4_outputs(7291) <= layer3_outputs(2013);
    layer4_outputs(7292) <= layer3_outputs(3501);
    layer4_outputs(7293) <= not(layer3_outputs(9433)) or (layer3_outputs(7661));
    layer4_outputs(7294) <= layer3_outputs(9436);
    layer4_outputs(7295) <= not(layer3_outputs(1636));
    layer4_outputs(7296) <= layer3_outputs(8612);
    layer4_outputs(7297) <= layer3_outputs(3538);
    layer4_outputs(7298) <= not(layer3_outputs(1105));
    layer4_outputs(7299) <= not((layer3_outputs(3930)) xor (layer3_outputs(9606)));
    layer4_outputs(7300) <= layer3_outputs(1904);
    layer4_outputs(7301) <= not(layer3_outputs(8642));
    layer4_outputs(7302) <= not((layer3_outputs(9456)) and (layer3_outputs(440)));
    layer4_outputs(7303) <= not(layer3_outputs(8817)) or (layer3_outputs(6993));
    layer4_outputs(7304) <= not(layer3_outputs(3573));
    layer4_outputs(7305) <= layer3_outputs(1377);
    layer4_outputs(7306) <= not(layer3_outputs(2059));
    layer4_outputs(7307) <= (layer3_outputs(4511)) and not (layer3_outputs(5416));
    layer4_outputs(7308) <= layer3_outputs(5260);
    layer4_outputs(7309) <= layer3_outputs(1344);
    layer4_outputs(7310) <= layer3_outputs(414);
    layer4_outputs(7311) <= layer3_outputs(7731);
    layer4_outputs(7312) <= (layer3_outputs(3949)) and not (layer3_outputs(9733));
    layer4_outputs(7313) <= not((layer3_outputs(5071)) or (layer3_outputs(2230)));
    layer4_outputs(7314) <= (layer3_outputs(2187)) or (layer3_outputs(8138));
    layer4_outputs(7315) <= not(layer3_outputs(8513));
    layer4_outputs(7316) <= layer3_outputs(2800);
    layer4_outputs(7317) <= not(layer3_outputs(2880));
    layer4_outputs(7318) <= not(layer3_outputs(1515)) or (layer3_outputs(3903));
    layer4_outputs(7319) <= layer3_outputs(1588);
    layer4_outputs(7320) <= layer3_outputs(6441);
    layer4_outputs(7321) <= layer3_outputs(1847);
    layer4_outputs(7322) <= layer3_outputs(8033);
    layer4_outputs(7323) <= (layer3_outputs(2314)) xor (layer3_outputs(8399));
    layer4_outputs(7324) <= layer3_outputs(4113);
    layer4_outputs(7325) <= layer3_outputs(5570);
    layer4_outputs(7326) <= layer3_outputs(9846);
    layer4_outputs(7327) <= not((layer3_outputs(2375)) or (layer3_outputs(4717)));
    layer4_outputs(7328) <= (layer3_outputs(8914)) xor (layer3_outputs(3975));
    layer4_outputs(7329) <= not(layer3_outputs(3987));
    layer4_outputs(7330) <= (layer3_outputs(2413)) and not (layer3_outputs(1154));
    layer4_outputs(7331) <= not((layer3_outputs(1288)) xor (layer3_outputs(3765)));
    layer4_outputs(7332) <= (layer3_outputs(4032)) xor (layer3_outputs(8799));
    layer4_outputs(7333) <= not(layer3_outputs(5270));
    layer4_outputs(7334) <= not(layer3_outputs(1301));
    layer4_outputs(7335) <= not(layer3_outputs(5432));
    layer4_outputs(7336) <= not((layer3_outputs(3459)) and (layer3_outputs(5165)));
    layer4_outputs(7337) <= layer3_outputs(7842);
    layer4_outputs(7338) <= layer3_outputs(165);
    layer4_outputs(7339) <= not(layer3_outputs(4963));
    layer4_outputs(7340) <= (layer3_outputs(7204)) and not (layer3_outputs(4315));
    layer4_outputs(7341) <= not((layer3_outputs(1966)) xor (layer3_outputs(8424)));
    layer4_outputs(7342) <= (layer3_outputs(6525)) xor (layer3_outputs(7600));
    layer4_outputs(7343) <= not(layer3_outputs(777)) or (layer3_outputs(4035));
    layer4_outputs(7344) <= not(layer3_outputs(6889));
    layer4_outputs(7345) <= not(layer3_outputs(7248));
    layer4_outputs(7346) <= layer3_outputs(6787);
    layer4_outputs(7347) <= (layer3_outputs(984)) xor (layer3_outputs(3558));
    layer4_outputs(7348) <= not(layer3_outputs(3332));
    layer4_outputs(7349) <= layer3_outputs(8243);
    layer4_outputs(7350) <= not((layer3_outputs(8481)) xor (layer3_outputs(8152)));
    layer4_outputs(7351) <= (layer3_outputs(8150)) and not (layer3_outputs(2588));
    layer4_outputs(7352) <= not(layer3_outputs(5102)) or (layer3_outputs(1332));
    layer4_outputs(7353) <= not((layer3_outputs(7117)) xor (layer3_outputs(7449)));
    layer4_outputs(7354) <= not(layer3_outputs(3803)) or (layer3_outputs(434));
    layer4_outputs(7355) <= layer3_outputs(6807);
    layer4_outputs(7356) <= layer3_outputs(2614);
    layer4_outputs(7357) <= not(layer3_outputs(4514));
    layer4_outputs(7358) <= layer3_outputs(5771);
    layer4_outputs(7359) <= not((layer3_outputs(1131)) and (layer3_outputs(2334)));
    layer4_outputs(7360) <= not(layer3_outputs(1363));
    layer4_outputs(7361) <= not(layer3_outputs(2702));
    layer4_outputs(7362) <= (layer3_outputs(9360)) or (layer3_outputs(6340));
    layer4_outputs(7363) <= layer3_outputs(9918);
    layer4_outputs(7364) <= not(layer3_outputs(5142));
    layer4_outputs(7365) <= layer3_outputs(2932);
    layer4_outputs(7366) <= layer3_outputs(5828);
    layer4_outputs(7367) <= layer3_outputs(6127);
    layer4_outputs(7368) <= not((layer3_outputs(323)) and (layer3_outputs(6275)));
    layer4_outputs(7369) <= (layer3_outputs(3065)) and not (layer3_outputs(2313));
    layer4_outputs(7370) <= layer3_outputs(8113);
    layer4_outputs(7371) <= (layer3_outputs(435)) and not (layer3_outputs(7247));
    layer4_outputs(7372) <= not((layer3_outputs(6118)) xor (layer3_outputs(1345)));
    layer4_outputs(7373) <= not(layer3_outputs(5241));
    layer4_outputs(7374) <= not(layer3_outputs(4187));
    layer4_outputs(7375) <= (layer3_outputs(1321)) and not (layer3_outputs(4706));
    layer4_outputs(7376) <= layer3_outputs(8932);
    layer4_outputs(7377) <= (layer3_outputs(6395)) or (layer3_outputs(3279));
    layer4_outputs(7378) <= (layer3_outputs(1511)) xor (layer3_outputs(7317));
    layer4_outputs(7379) <= (layer3_outputs(9889)) xor (layer3_outputs(3742));
    layer4_outputs(7380) <= not(layer3_outputs(7795));
    layer4_outputs(7381) <= layer3_outputs(882);
    layer4_outputs(7382) <= (layer3_outputs(7466)) xor (layer3_outputs(7443));
    layer4_outputs(7383) <= (layer3_outputs(422)) and not (layer3_outputs(9460));
    layer4_outputs(7384) <= not(layer3_outputs(1522));
    layer4_outputs(7385) <= layer3_outputs(2025);
    layer4_outputs(7386) <= (layer3_outputs(4354)) xor (layer3_outputs(8596));
    layer4_outputs(7387) <= not((layer3_outputs(4301)) xor (layer3_outputs(3536)));
    layer4_outputs(7388) <= (layer3_outputs(2387)) and (layer3_outputs(3819));
    layer4_outputs(7389) <= layer3_outputs(5760);
    layer4_outputs(7390) <= not(layer3_outputs(3134));
    layer4_outputs(7391) <= not(layer3_outputs(1030));
    layer4_outputs(7392) <= (layer3_outputs(1331)) or (layer3_outputs(8545));
    layer4_outputs(7393) <= not((layer3_outputs(6947)) xor (layer3_outputs(8686)));
    layer4_outputs(7394) <= not(layer3_outputs(418));
    layer4_outputs(7395) <= layer3_outputs(1042);
    layer4_outputs(7396) <= not(layer3_outputs(806));
    layer4_outputs(7397) <= layer3_outputs(4529);
    layer4_outputs(7398) <= layer3_outputs(3627);
    layer4_outputs(7399) <= layer3_outputs(3291);
    layer4_outputs(7400) <= layer3_outputs(3046);
    layer4_outputs(7401) <= not(layer3_outputs(3040)) or (layer3_outputs(571));
    layer4_outputs(7402) <= not((layer3_outputs(6732)) xor (layer3_outputs(4021)));
    layer4_outputs(7403) <= layer3_outputs(5840);
    layer4_outputs(7404) <= not(layer3_outputs(2213));
    layer4_outputs(7405) <= not((layer3_outputs(9891)) xor (layer3_outputs(1366)));
    layer4_outputs(7406) <= not(layer3_outputs(8347));
    layer4_outputs(7407) <= not(layer3_outputs(9771));
    layer4_outputs(7408) <= (layer3_outputs(8923)) or (layer3_outputs(9225));
    layer4_outputs(7409) <= (layer3_outputs(2663)) xor (layer3_outputs(4654));
    layer4_outputs(7410) <= not(layer3_outputs(9626));
    layer4_outputs(7411) <= not(layer3_outputs(9610));
    layer4_outputs(7412) <= layer3_outputs(8744);
    layer4_outputs(7413) <= not(layer3_outputs(2362));
    layer4_outputs(7414) <= (layer3_outputs(4289)) and not (layer3_outputs(7991));
    layer4_outputs(7415) <= not(layer3_outputs(9263));
    layer4_outputs(7416) <= not((layer3_outputs(3874)) and (layer3_outputs(3030)));
    layer4_outputs(7417) <= (layer3_outputs(4455)) and not (layer3_outputs(3355));
    layer4_outputs(7418) <= (layer3_outputs(5461)) xor (layer3_outputs(5938));
    layer4_outputs(7419) <= (layer3_outputs(2469)) xor (layer3_outputs(8332));
    layer4_outputs(7420) <= layer3_outputs(7075);
    layer4_outputs(7421) <= layer3_outputs(6067);
    layer4_outputs(7422) <= layer3_outputs(3406);
    layer4_outputs(7423) <= layer3_outputs(9165);
    layer4_outputs(7424) <= not(layer3_outputs(9047));
    layer4_outputs(7425) <= not(layer3_outputs(6348));
    layer4_outputs(7426) <= layer3_outputs(9528);
    layer4_outputs(7427) <= not(layer3_outputs(3254));
    layer4_outputs(7428) <= (layer3_outputs(981)) and not (layer3_outputs(7121));
    layer4_outputs(7429) <= not(layer3_outputs(2106));
    layer4_outputs(7430) <= not(layer3_outputs(923));
    layer4_outputs(7431) <= not(layer3_outputs(2966));
    layer4_outputs(7432) <= not((layer3_outputs(7870)) xor (layer3_outputs(3974)));
    layer4_outputs(7433) <= (layer3_outputs(8975)) and (layer3_outputs(901));
    layer4_outputs(7434) <= layer3_outputs(8802);
    layer4_outputs(7435) <= not(layer3_outputs(9445));
    layer4_outputs(7436) <= layer3_outputs(1560);
    layer4_outputs(7437) <= layer3_outputs(816);
    layer4_outputs(7438) <= (layer3_outputs(7476)) xor (layer3_outputs(7350));
    layer4_outputs(7439) <= layer3_outputs(6336);
    layer4_outputs(7440) <= layer3_outputs(9732);
    layer4_outputs(7441) <= '0';
    layer4_outputs(7442) <= not(layer3_outputs(8958));
    layer4_outputs(7443) <= not((layer3_outputs(2587)) or (layer3_outputs(34)));
    layer4_outputs(7444) <= not(layer3_outputs(6398)) or (layer3_outputs(5952));
    layer4_outputs(7445) <= (layer3_outputs(6380)) and (layer3_outputs(5460));
    layer4_outputs(7446) <= (layer3_outputs(8742)) and not (layer3_outputs(6785));
    layer4_outputs(7447) <= layer3_outputs(7074);
    layer4_outputs(7448) <= not(layer3_outputs(252));
    layer4_outputs(7449) <= not((layer3_outputs(9193)) xor (layer3_outputs(6617)));
    layer4_outputs(7450) <= (layer3_outputs(10137)) and not (layer3_outputs(1332));
    layer4_outputs(7451) <= (layer3_outputs(4516)) and not (layer3_outputs(9777));
    layer4_outputs(7452) <= layer3_outputs(8869);
    layer4_outputs(7453) <= not((layer3_outputs(8919)) xor (layer3_outputs(4392)));
    layer4_outputs(7454) <= layer3_outputs(9980);
    layer4_outputs(7455) <= not(layer3_outputs(732));
    layer4_outputs(7456) <= layer3_outputs(15);
    layer4_outputs(7457) <= not(layer3_outputs(9594));
    layer4_outputs(7458) <= layer3_outputs(355);
    layer4_outputs(7459) <= (layer3_outputs(6524)) and not (layer3_outputs(3226));
    layer4_outputs(7460) <= not((layer3_outputs(8211)) or (layer3_outputs(7457)));
    layer4_outputs(7461) <= not((layer3_outputs(4916)) or (layer3_outputs(3598)));
    layer4_outputs(7462) <= (layer3_outputs(1691)) and not (layer3_outputs(5104));
    layer4_outputs(7463) <= not(layer3_outputs(6451));
    layer4_outputs(7464) <= not(layer3_outputs(6718));
    layer4_outputs(7465) <= layer3_outputs(1390);
    layer4_outputs(7466) <= (layer3_outputs(971)) and not (layer3_outputs(455));
    layer4_outputs(7467) <= not((layer3_outputs(616)) xor (layer3_outputs(6141)));
    layer4_outputs(7468) <= not((layer3_outputs(5214)) and (layer3_outputs(8350)));
    layer4_outputs(7469) <= not(layer3_outputs(1672));
    layer4_outputs(7470) <= not(layer3_outputs(8052)) or (layer3_outputs(1809));
    layer4_outputs(7471) <= (layer3_outputs(695)) xor (layer3_outputs(2374));
    layer4_outputs(7472) <= not((layer3_outputs(4729)) xor (layer3_outputs(7104)));
    layer4_outputs(7473) <= layer3_outputs(8565);
    layer4_outputs(7474) <= layer3_outputs(545);
    layer4_outputs(7475) <= not(layer3_outputs(8193)) or (layer3_outputs(9743));
    layer4_outputs(7476) <= not(layer3_outputs(8186));
    layer4_outputs(7477) <= not(layer3_outputs(6837));
    layer4_outputs(7478) <= not((layer3_outputs(2976)) or (layer3_outputs(9623)));
    layer4_outputs(7479) <= not(layer3_outputs(7019));
    layer4_outputs(7480) <= not(layer3_outputs(3261)) or (layer3_outputs(201));
    layer4_outputs(7481) <= not(layer3_outputs(1870));
    layer4_outputs(7482) <= not(layer3_outputs(3760));
    layer4_outputs(7483) <= layer3_outputs(10200);
    layer4_outputs(7484) <= (layer3_outputs(4671)) xor (layer3_outputs(1059));
    layer4_outputs(7485) <= not(layer3_outputs(5013));
    layer4_outputs(7486) <= (layer3_outputs(7828)) or (layer3_outputs(8094));
    layer4_outputs(7487) <= not((layer3_outputs(5583)) xor (layer3_outputs(9710)));
    layer4_outputs(7488) <= layer3_outputs(9637);
    layer4_outputs(7489) <= not((layer3_outputs(6704)) xor (layer3_outputs(3018)));
    layer4_outputs(7490) <= not(layer3_outputs(8045));
    layer4_outputs(7491) <= layer3_outputs(3183);
    layer4_outputs(7492) <= not(layer3_outputs(5133)) or (layer3_outputs(5412));
    layer4_outputs(7493) <= not((layer3_outputs(5051)) xor (layer3_outputs(8296)));
    layer4_outputs(7494) <= not(layer3_outputs(841));
    layer4_outputs(7495) <= not(layer3_outputs(650));
    layer4_outputs(7496) <= layer3_outputs(1915);
    layer4_outputs(7497) <= layer3_outputs(8055);
    layer4_outputs(7498) <= not((layer3_outputs(9200)) or (layer3_outputs(7915)));
    layer4_outputs(7499) <= layer3_outputs(8583);
    layer4_outputs(7500) <= not(layer3_outputs(5449));
    layer4_outputs(7501) <= (layer3_outputs(8635)) and not (layer3_outputs(4125));
    layer4_outputs(7502) <= not(layer3_outputs(2782));
    layer4_outputs(7503) <= layer3_outputs(3616);
    layer4_outputs(7504) <= not(layer3_outputs(7461));
    layer4_outputs(7505) <= layer3_outputs(9189);
    layer4_outputs(7506) <= (layer3_outputs(1744)) and not (layer3_outputs(1195));
    layer4_outputs(7507) <= not(layer3_outputs(2699));
    layer4_outputs(7508) <= layer3_outputs(1712);
    layer4_outputs(7509) <= (layer3_outputs(2060)) and (layer3_outputs(1941));
    layer4_outputs(7510) <= not(layer3_outputs(6977));
    layer4_outputs(7511) <= not(layer3_outputs(3423)) or (layer3_outputs(4193));
    layer4_outputs(7512) <= not(layer3_outputs(105)) or (layer3_outputs(1271));
    layer4_outputs(7513) <= layer3_outputs(8557);
    layer4_outputs(7514) <= layer3_outputs(6045);
    layer4_outputs(7515) <= not(layer3_outputs(5336));
    layer4_outputs(7516) <= not(layer3_outputs(5832));
    layer4_outputs(7517) <= not(layer3_outputs(524)) or (layer3_outputs(3599));
    layer4_outputs(7518) <= layer3_outputs(1531);
    layer4_outputs(7519) <= layer3_outputs(1691);
    layer4_outputs(7520) <= not(layer3_outputs(133));
    layer4_outputs(7521) <= layer3_outputs(6935);
    layer4_outputs(7522) <= not((layer3_outputs(1431)) xor (layer3_outputs(1394)));
    layer4_outputs(7523) <= not(layer3_outputs(1707));
    layer4_outputs(7524) <= (layer3_outputs(8398)) xor (layer3_outputs(9069));
    layer4_outputs(7525) <= not((layer3_outputs(3460)) xor (layer3_outputs(7996)));
    layer4_outputs(7526) <= not((layer3_outputs(9541)) and (layer3_outputs(2569)));
    layer4_outputs(7527) <= not((layer3_outputs(5089)) xor (layer3_outputs(4197)));
    layer4_outputs(7528) <= not(layer3_outputs(4750));
    layer4_outputs(7529) <= layer3_outputs(282);
    layer4_outputs(7530) <= not((layer3_outputs(3025)) xor (layer3_outputs(2074)));
    layer4_outputs(7531) <= not((layer3_outputs(7625)) xor (layer3_outputs(9169)));
    layer4_outputs(7532) <= layer3_outputs(7267);
    layer4_outputs(7533) <= layer3_outputs(5883);
    layer4_outputs(7534) <= not((layer3_outputs(7208)) and (layer3_outputs(8232)));
    layer4_outputs(7535) <= not((layer3_outputs(8089)) xor (layer3_outputs(4154)));
    layer4_outputs(7536) <= '1';
    layer4_outputs(7537) <= layer3_outputs(6226);
    layer4_outputs(7538) <= not(layer3_outputs(2306));
    layer4_outputs(7539) <= layer3_outputs(4163);
    layer4_outputs(7540) <= not((layer3_outputs(7621)) or (layer3_outputs(3891)));
    layer4_outputs(7541) <= not(layer3_outputs(1901)) or (layer3_outputs(2092));
    layer4_outputs(7542) <= not((layer3_outputs(1427)) xor (layer3_outputs(3644)));
    layer4_outputs(7543) <= not(layer3_outputs(6143));
    layer4_outputs(7544) <= not(layer3_outputs(5467));
    layer4_outputs(7545) <= (layer3_outputs(7908)) and not (layer3_outputs(479));
    layer4_outputs(7546) <= (layer3_outputs(7088)) and not (layer3_outputs(5152));
    layer4_outputs(7547) <= not(layer3_outputs(2661));
    layer4_outputs(7548) <= not((layer3_outputs(648)) xor (layer3_outputs(724)));
    layer4_outputs(7549) <= (layer3_outputs(9920)) and not (layer3_outputs(47));
    layer4_outputs(7550) <= layer3_outputs(9315);
    layer4_outputs(7551) <= not(layer3_outputs(3206)) or (layer3_outputs(4507));
    layer4_outputs(7552) <= not((layer3_outputs(9194)) and (layer3_outputs(3737)));
    layer4_outputs(7553) <= layer3_outputs(2145);
    layer4_outputs(7554) <= not((layer3_outputs(592)) and (layer3_outputs(5595)));
    layer4_outputs(7555) <= not(layer3_outputs(4617));
    layer4_outputs(7556) <= (layer3_outputs(8096)) xor (layer3_outputs(4803));
    layer4_outputs(7557) <= (layer3_outputs(3885)) and not (layer3_outputs(481));
    layer4_outputs(7558) <= not(layer3_outputs(7765));
    layer4_outputs(7559) <= layer3_outputs(2424);
    layer4_outputs(7560) <= not(layer3_outputs(1581));
    layer4_outputs(7561) <= (layer3_outputs(5025)) and not (layer3_outputs(217));
    layer4_outputs(7562) <= not((layer3_outputs(3105)) xor (layer3_outputs(1988)));
    layer4_outputs(7563) <= layer3_outputs(6403);
    layer4_outputs(7564) <= not(layer3_outputs(5884));
    layer4_outputs(7565) <= not(layer3_outputs(9615));
    layer4_outputs(7566) <= (layer3_outputs(6339)) xor (layer3_outputs(6001));
    layer4_outputs(7567) <= layer3_outputs(617);
    layer4_outputs(7568) <= (layer3_outputs(4008)) xor (layer3_outputs(6965));
    layer4_outputs(7569) <= not(layer3_outputs(73));
    layer4_outputs(7570) <= not(layer3_outputs(1221));
    layer4_outputs(7571) <= '1';
    layer4_outputs(7572) <= (layer3_outputs(1651)) xor (layer3_outputs(9948));
    layer4_outputs(7573) <= (layer3_outputs(1610)) or (layer3_outputs(1693));
    layer4_outputs(7574) <= (layer3_outputs(2148)) xor (layer3_outputs(10145));
    layer4_outputs(7575) <= not((layer3_outputs(6202)) and (layer3_outputs(4723)));
    layer4_outputs(7576) <= layer3_outputs(9608);
    layer4_outputs(7577) <= (layer3_outputs(4386)) and not (layer3_outputs(171));
    layer4_outputs(7578) <= (layer3_outputs(9451)) xor (layer3_outputs(3565));
    layer4_outputs(7579) <= (layer3_outputs(6240)) or (layer3_outputs(2589));
    layer4_outputs(7580) <= layer3_outputs(9105);
    layer4_outputs(7581) <= not(layer3_outputs(419));
    layer4_outputs(7582) <= not((layer3_outputs(9335)) or (layer3_outputs(4805)));
    layer4_outputs(7583) <= not(layer3_outputs(8497)) or (layer3_outputs(9731));
    layer4_outputs(7584) <= not((layer3_outputs(7803)) xor (layer3_outputs(7958)));
    layer4_outputs(7585) <= layer3_outputs(6199);
    layer4_outputs(7586) <= not(layer3_outputs(2809));
    layer4_outputs(7587) <= not((layer3_outputs(8308)) or (layer3_outputs(201)));
    layer4_outputs(7588) <= not((layer3_outputs(8916)) xor (layer3_outputs(9648)));
    layer4_outputs(7589) <= not((layer3_outputs(4330)) or (layer3_outputs(3649)));
    layer4_outputs(7590) <= (layer3_outputs(3856)) and not (layer3_outputs(5911));
    layer4_outputs(7591) <= not((layer3_outputs(6217)) xor (layer3_outputs(210)));
    layer4_outputs(7592) <= not(layer3_outputs(4320));
    layer4_outputs(7593) <= not(layer3_outputs(7611));
    layer4_outputs(7594) <= not(layer3_outputs(5510)) or (layer3_outputs(3691));
    layer4_outputs(7595) <= (layer3_outputs(1124)) and not (layer3_outputs(8295));
    layer4_outputs(7596) <= layer3_outputs(7675);
    layer4_outputs(7597) <= (layer3_outputs(4938)) xor (layer3_outputs(5708));
    layer4_outputs(7598) <= not(layer3_outputs(9403));
    layer4_outputs(7599) <= not((layer3_outputs(1450)) xor (layer3_outputs(1299)));
    layer4_outputs(7600) <= not((layer3_outputs(1186)) and (layer3_outputs(7936)));
    layer4_outputs(7601) <= layer3_outputs(4234);
    layer4_outputs(7602) <= not((layer3_outputs(1901)) xor (layer3_outputs(4612)));
    layer4_outputs(7603) <= (layer3_outputs(3151)) and not (layer3_outputs(6860));
    layer4_outputs(7604) <= layer3_outputs(1502);
    layer4_outputs(7605) <= not(layer3_outputs(8877));
    layer4_outputs(7606) <= not(layer3_outputs(5539));
    layer4_outputs(7607) <= layer3_outputs(3641);
    layer4_outputs(7608) <= layer3_outputs(700);
    layer4_outputs(7609) <= not(layer3_outputs(6441));
    layer4_outputs(7610) <= not(layer3_outputs(5204));
    layer4_outputs(7611) <= (layer3_outputs(9772)) or (layer3_outputs(8127));
    layer4_outputs(7612) <= not((layer3_outputs(3893)) or (layer3_outputs(3739)));
    layer4_outputs(7613) <= layer3_outputs(4993);
    layer4_outputs(7614) <= layer3_outputs(6670);
    layer4_outputs(7615) <= not((layer3_outputs(4023)) xor (layer3_outputs(8807)));
    layer4_outputs(7616) <= (layer3_outputs(6836)) or (layer3_outputs(3274));
    layer4_outputs(7617) <= '0';
    layer4_outputs(7618) <= (layer3_outputs(8793)) xor (layer3_outputs(8071));
    layer4_outputs(7619) <= (layer3_outputs(6013)) xor (layer3_outputs(1628));
    layer4_outputs(7620) <= not(layer3_outputs(2682));
    layer4_outputs(7621) <= layer3_outputs(5485);
    layer4_outputs(7622) <= not(layer3_outputs(9908));
    layer4_outputs(7623) <= not(layer3_outputs(8831));
    layer4_outputs(7624) <= not(layer3_outputs(9726));
    layer4_outputs(7625) <= not((layer3_outputs(7307)) or (layer3_outputs(2015)));
    layer4_outputs(7626) <= layer3_outputs(9596);
    layer4_outputs(7627) <= layer3_outputs(7579);
    layer4_outputs(7628) <= '0';
    layer4_outputs(7629) <= not(layer3_outputs(2745));
    layer4_outputs(7630) <= not((layer3_outputs(3126)) or (layer3_outputs(1167)));
    layer4_outputs(7631) <= layer3_outputs(2178);
    layer4_outputs(7632) <= not(layer3_outputs(8027));
    layer4_outputs(7633) <= not((layer3_outputs(7768)) xor (layer3_outputs(2764)));
    layer4_outputs(7634) <= layer3_outputs(7697);
    layer4_outputs(7635) <= layer3_outputs(7963);
    layer4_outputs(7636) <= layer3_outputs(437);
    layer4_outputs(7637) <= not(layer3_outputs(3688));
    layer4_outputs(7638) <= not(layer3_outputs(6010));
    layer4_outputs(7639) <= layer3_outputs(1510);
    layer4_outputs(7640) <= not((layer3_outputs(8475)) xor (layer3_outputs(7746)));
    layer4_outputs(7641) <= layer3_outputs(1389);
    layer4_outputs(7642) <= (layer3_outputs(5837)) and not (layer3_outputs(487));
    layer4_outputs(7643) <= not(layer3_outputs(4716));
    layer4_outputs(7644) <= not((layer3_outputs(4095)) or (layer3_outputs(7837)));
    layer4_outputs(7645) <= not(layer3_outputs(53));
    layer4_outputs(7646) <= (layer3_outputs(6986)) or (layer3_outputs(6128));
    layer4_outputs(7647) <= not(layer3_outputs(6804));
    layer4_outputs(7648) <= not(layer3_outputs(2474)) or (layer3_outputs(9227));
    layer4_outputs(7649) <= layer3_outputs(7552);
    layer4_outputs(7650) <= (layer3_outputs(10138)) and (layer3_outputs(10038));
    layer4_outputs(7651) <= (layer3_outputs(3717)) xor (layer3_outputs(7110));
    layer4_outputs(7652) <= not(layer3_outputs(9128)) or (layer3_outputs(5229));
    layer4_outputs(7653) <= (layer3_outputs(4343)) xor (layer3_outputs(6581));
    layer4_outputs(7654) <= (layer3_outputs(7001)) or (layer3_outputs(7384));
    layer4_outputs(7655) <= layer3_outputs(4650);
    layer4_outputs(7656) <= not(layer3_outputs(5256));
    layer4_outputs(7657) <= not(layer3_outputs(7413));
    layer4_outputs(7658) <= not((layer3_outputs(9021)) xor (layer3_outputs(7136)));
    layer4_outputs(7659) <= (layer3_outputs(4100)) xor (layer3_outputs(321));
    layer4_outputs(7660) <= not((layer3_outputs(9491)) and (layer3_outputs(4331)));
    layer4_outputs(7661) <= (layer3_outputs(1466)) and (layer3_outputs(2594));
    layer4_outputs(7662) <= (layer3_outputs(167)) or (layer3_outputs(2472));
    layer4_outputs(7663) <= layer3_outputs(5696);
    layer4_outputs(7664) <= not(layer3_outputs(3807));
    layer4_outputs(7665) <= not((layer3_outputs(3837)) xor (layer3_outputs(10123)));
    layer4_outputs(7666) <= (layer3_outputs(958)) and not (layer3_outputs(7699));
    layer4_outputs(7667) <= not((layer3_outputs(9034)) xor (layer3_outputs(6802)));
    layer4_outputs(7668) <= layer3_outputs(4114);
    layer4_outputs(7669) <= not(layer3_outputs(2541));
    layer4_outputs(7670) <= (layer3_outputs(5176)) xor (layer3_outputs(7006));
    layer4_outputs(7671) <= not((layer3_outputs(7642)) xor (layer3_outputs(9877)));
    layer4_outputs(7672) <= layer3_outputs(7457);
    layer4_outputs(7673) <= not((layer3_outputs(1674)) or (layer3_outputs(3382)));
    layer4_outputs(7674) <= layer3_outputs(4654);
    layer4_outputs(7675) <= not(layer3_outputs(500));
    layer4_outputs(7676) <= not(layer3_outputs(9978));
    layer4_outputs(7677) <= (layer3_outputs(8062)) xor (layer3_outputs(8638));
    layer4_outputs(7678) <= layer3_outputs(12);
    layer4_outputs(7679) <= layer3_outputs(245);
    layer4_outputs(7680) <= not(layer3_outputs(5094));
    layer4_outputs(7681) <= layer3_outputs(4550);
    layer4_outputs(7682) <= not(layer3_outputs(2972));
    layer4_outputs(7683) <= (layer3_outputs(9557)) and not (layer3_outputs(3363));
    layer4_outputs(7684) <= layer3_outputs(9362);
    layer4_outputs(7685) <= not((layer3_outputs(9384)) or (layer3_outputs(6834)));
    layer4_outputs(7686) <= not((layer3_outputs(9249)) xor (layer3_outputs(1505)));
    layer4_outputs(7687) <= (layer3_outputs(5304)) and (layer3_outputs(5549));
    layer4_outputs(7688) <= not(layer3_outputs(9411));
    layer4_outputs(7689) <= layer3_outputs(3787);
    layer4_outputs(7690) <= layer3_outputs(3638);
    layer4_outputs(7691) <= not((layer3_outputs(1524)) xor (layer3_outputs(443)));
    layer4_outputs(7692) <= layer3_outputs(4809);
    layer4_outputs(7693) <= layer3_outputs(9654);
    layer4_outputs(7694) <= not((layer3_outputs(7253)) xor (layer3_outputs(9361)));
    layer4_outputs(7695) <= not(layer3_outputs(3346));
    layer4_outputs(7696) <= not(layer3_outputs(2503));
    layer4_outputs(7697) <= not((layer3_outputs(8192)) xor (layer3_outputs(1341)));
    layer4_outputs(7698) <= not((layer3_outputs(7344)) xor (layer3_outputs(2568)));
    layer4_outputs(7699) <= layer3_outputs(4203);
    layer4_outputs(7700) <= (layer3_outputs(3991)) or (layer3_outputs(8692));
    layer4_outputs(7701) <= not(layer3_outputs(1706)) or (layer3_outputs(5161));
    layer4_outputs(7702) <= not(layer3_outputs(6595));
    layer4_outputs(7703) <= (layer3_outputs(9725)) and (layer3_outputs(5065));
    layer4_outputs(7704) <= (layer3_outputs(6191)) xor (layer3_outputs(3772));
    layer4_outputs(7705) <= (layer3_outputs(3695)) and not (layer3_outputs(3152));
    layer4_outputs(7706) <= layer3_outputs(4965);
    layer4_outputs(7707) <= (layer3_outputs(8866)) and (layer3_outputs(9342));
    layer4_outputs(7708) <= not(layer3_outputs(6961));
    layer4_outputs(7709) <= layer3_outputs(2719);
    layer4_outputs(7710) <= not(layer3_outputs(5720));
    layer4_outputs(7711) <= layer3_outputs(1454);
    layer4_outputs(7712) <= not((layer3_outputs(104)) and (layer3_outputs(4601)));
    layer4_outputs(7713) <= not((layer3_outputs(8214)) xor (layer3_outputs(5943)));
    layer4_outputs(7714) <= (layer3_outputs(2501)) xor (layer3_outputs(8885));
    layer4_outputs(7715) <= (layer3_outputs(3459)) or (layer3_outputs(5675));
    layer4_outputs(7716) <= layer3_outputs(7829);
    layer4_outputs(7717) <= not(layer3_outputs(1985));
    layer4_outputs(7718) <= (layer3_outputs(6014)) and not (layer3_outputs(7749));
    layer4_outputs(7719) <= (layer3_outputs(4981)) and not (layer3_outputs(2948));
    layer4_outputs(7720) <= not((layer3_outputs(7673)) xor (layer3_outputs(6521)));
    layer4_outputs(7721) <= not(layer3_outputs(2638)) or (layer3_outputs(7794));
    layer4_outputs(7722) <= layer3_outputs(10059);
    layer4_outputs(7723) <= not(layer3_outputs(9011));
    layer4_outputs(7724) <= not(layer3_outputs(3557));
    layer4_outputs(7725) <= layer3_outputs(5191);
    layer4_outputs(7726) <= not((layer3_outputs(127)) xor (layer3_outputs(8251)));
    layer4_outputs(7727) <= not((layer3_outputs(800)) or (layer3_outputs(9564)));
    layer4_outputs(7728) <= not((layer3_outputs(2238)) and (layer3_outputs(241)));
    layer4_outputs(7729) <= not((layer3_outputs(2929)) and (layer3_outputs(8641)));
    layer4_outputs(7730) <= not((layer3_outputs(9783)) or (layer3_outputs(3149)));
    layer4_outputs(7731) <= not(layer3_outputs(7129));
    layer4_outputs(7732) <= not(layer3_outputs(3860)) or (layer3_outputs(591));
    layer4_outputs(7733) <= layer3_outputs(7056);
    layer4_outputs(7734) <= (layer3_outputs(10079)) xor (layer3_outputs(8886));
    layer4_outputs(7735) <= not(layer3_outputs(9999));
    layer4_outputs(7736) <= (layer3_outputs(2328)) and not (layer3_outputs(3384));
    layer4_outputs(7737) <= layer3_outputs(8831);
    layer4_outputs(7738) <= (layer3_outputs(6088)) or (layer3_outputs(8360));
    layer4_outputs(7739) <= not(layer3_outputs(1999));
    layer4_outputs(7740) <= layer3_outputs(4517);
    layer4_outputs(7741) <= not((layer3_outputs(4482)) xor (layer3_outputs(3667)));
    layer4_outputs(7742) <= not((layer3_outputs(5430)) xor (layer3_outputs(4549)));
    layer4_outputs(7743) <= layer3_outputs(7338);
    layer4_outputs(7744) <= not(layer3_outputs(1295));
    layer4_outputs(7745) <= not(layer3_outputs(9487));
    layer4_outputs(7746) <= not(layer3_outputs(1679));
    layer4_outputs(7747) <= not((layer3_outputs(1381)) and (layer3_outputs(8968)));
    layer4_outputs(7748) <= not(layer3_outputs(4252));
    layer4_outputs(7749) <= not(layer3_outputs(634));
    layer4_outputs(7750) <= layer3_outputs(8276);
    layer4_outputs(7751) <= not((layer3_outputs(9286)) xor (layer3_outputs(2346)));
    layer4_outputs(7752) <= not((layer3_outputs(7672)) or (layer3_outputs(5115)));
    layer4_outputs(7753) <= layer3_outputs(982);
    layer4_outputs(7754) <= not(layer3_outputs(5400));
    layer4_outputs(7755) <= layer3_outputs(5270);
    layer4_outputs(7756) <= (layer3_outputs(9863)) and not (layer3_outputs(5598));
    layer4_outputs(7757) <= (layer3_outputs(3570)) and not (layer3_outputs(7613));
    layer4_outputs(7758) <= (layer3_outputs(8004)) or (layer3_outputs(8281));
    layer4_outputs(7759) <= not(layer3_outputs(5423));
    layer4_outputs(7760) <= (layer3_outputs(1433)) xor (layer3_outputs(2552));
    layer4_outputs(7761) <= not(layer3_outputs(9860)) or (layer3_outputs(9744));
    layer4_outputs(7762) <= not((layer3_outputs(7319)) and (layer3_outputs(488)));
    layer4_outputs(7763) <= layer3_outputs(809);
    layer4_outputs(7764) <= not((layer3_outputs(6999)) xor (layer3_outputs(6156)));
    layer4_outputs(7765) <= (layer3_outputs(2772)) xor (layer3_outputs(5818));
    layer4_outputs(7766) <= (layer3_outputs(6290)) and not (layer3_outputs(558));
    layer4_outputs(7767) <= (layer3_outputs(7729)) and not (layer3_outputs(3165));
    layer4_outputs(7768) <= not((layer3_outputs(5469)) xor (layer3_outputs(3585)));
    layer4_outputs(7769) <= layer3_outputs(6919);
    layer4_outputs(7770) <= (layer3_outputs(4413)) or (layer3_outputs(1567));
    layer4_outputs(7771) <= layer3_outputs(810);
    layer4_outputs(7772) <= layer3_outputs(7153);
    layer4_outputs(7773) <= not(layer3_outputs(5785));
    layer4_outputs(7774) <= not(layer3_outputs(6411)) or (layer3_outputs(6911));
    layer4_outputs(7775) <= (layer3_outputs(5441)) xor (layer3_outputs(10060));
    layer4_outputs(7776) <= (layer3_outputs(9089)) xor (layer3_outputs(7519));
    layer4_outputs(7777) <= not(layer3_outputs(407));
    layer4_outputs(7778) <= (layer3_outputs(5210)) or (layer3_outputs(8546));
    layer4_outputs(7779) <= (layer3_outputs(2250)) xor (layer3_outputs(6519));
    layer4_outputs(7780) <= layer3_outputs(9410);
    layer4_outputs(7781) <= layer3_outputs(8184);
    layer4_outputs(7782) <= (layer3_outputs(6155)) and not (layer3_outputs(6692));
    layer4_outputs(7783) <= layer3_outputs(9603);
    layer4_outputs(7784) <= layer3_outputs(1181);
    layer4_outputs(7785) <= (layer3_outputs(1754)) and not (layer3_outputs(736));
    layer4_outputs(7786) <= not(layer3_outputs(2859));
    layer4_outputs(7787) <= not((layer3_outputs(3779)) xor (layer3_outputs(6516)));
    layer4_outputs(7788) <= (layer3_outputs(7173)) and not (layer3_outputs(5869));
    layer4_outputs(7789) <= (layer3_outputs(8525)) and (layer3_outputs(9432));
    layer4_outputs(7790) <= layer3_outputs(2020);
    layer4_outputs(7791) <= layer3_outputs(415);
    layer4_outputs(7792) <= layer3_outputs(9075);
    layer4_outputs(7793) <= (layer3_outputs(5120)) and not (layer3_outputs(3626));
    layer4_outputs(7794) <= not(layer3_outputs(7594)) or (layer3_outputs(9951));
    layer4_outputs(7795) <= layer3_outputs(255);
    layer4_outputs(7796) <= not(layer3_outputs(4647));
    layer4_outputs(7797) <= not((layer3_outputs(5257)) xor (layer3_outputs(3101)));
    layer4_outputs(7798) <= not(layer3_outputs(8521));
    layer4_outputs(7799) <= not(layer3_outputs(6694));
    layer4_outputs(7800) <= (layer3_outputs(3339)) xor (layer3_outputs(9909));
    layer4_outputs(7801) <= layer3_outputs(5710);
    layer4_outputs(7802) <= not(layer3_outputs(10156));
    layer4_outputs(7803) <= layer3_outputs(30);
    layer4_outputs(7804) <= layer3_outputs(7628);
    layer4_outputs(7805) <= not(layer3_outputs(7536));
    layer4_outputs(7806) <= layer3_outputs(8593);
    layer4_outputs(7807) <= not(layer3_outputs(7763));
    layer4_outputs(7808) <= (layer3_outputs(5942)) xor (layer3_outputs(7818));
    layer4_outputs(7809) <= layer3_outputs(8890);
    layer4_outputs(7810) <= (layer3_outputs(3410)) and (layer3_outputs(7720));
    layer4_outputs(7811) <= (layer3_outputs(436)) and not (layer3_outputs(5390));
    layer4_outputs(7812) <= '1';
    layer4_outputs(7813) <= layer3_outputs(945);
    layer4_outputs(7814) <= (layer3_outputs(9785)) and (layer3_outputs(6833));
    layer4_outputs(7815) <= not(layer3_outputs(1439));
    layer4_outputs(7816) <= layer3_outputs(1428);
    layer4_outputs(7817) <= layer3_outputs(594);
    layer4_outputs(7818) <= (layer3_outputs(2715)) or (layer3_outputs(1479));
    layer4_outputs(7819) <= layer3_outputs(9983);
    layer4_outputs(7820) <= not(layer3_outputs(9197));
    layer4_outputs(7821) <= layer3_outputs(3879);
    layer4_outputs(7822) <= not(layer3_outputs(8988)) or (layer3_outputs(4061));
    layer4_outputs(7823) <= layer3_outputs(8590);
    layer4_outputs(7824) <= not(layer3_outputs(6004));
    layer4_outputs(7825) <= not(layer3_outputs(4188));
    layer4_outputs(7826) <= not(layer3_outputs(4545));
    layer4_outputs(7827) <= '0';
    layer4_outputs(7828) <= layer3_outputs(6390);
    layer4_outputs(7829) <= layer3_outputs(3321);
    layer4_outputs(7830) <= not(layer3_outputs(2712));
    layer4_outputs(7831) <= not(layer3_outputs(7537));
    layer4_outputs(7832) <= not(layer3_outputs(9267));
    layer4_outputs(7833) <= (layer3_outputs(1934)) xor (layer3_outputs(4079));
    layer4_outputs(7834) <= not((layer3_outputs(876)) and (layer3_outputs(3732)));
    layer4_outputs(7835) <= not(layer3_outputs(289)) or (layer3_outputs(1234));
    layer4_outputs(7836) <= not(layer3_outputs(9784));
    layer4_outputs(7837) <= not(layer3_outputs(1578));
    layer4_outputs(7838) <= not(layer3_outputs(6045));
    layer4_outputs(7839) <= not(layer3_outputs(4342)) or (layer3_outputs(4307));
    layer4_outputs(7840) <= not(layer3_outputs(3150));
    layer4_outputs(7841) <= not(layer3_outputs(3228)) or (layer3_outputs(7444));
    layer4_outputs(7842) <= layer3_outputs(60);
    layer4_outputs(7843) <= not(layer3_outputs(7816));
    layer4_outputs(7844) <= layer3_outputs(3834);
    layer4_outputs(7845) <= not(layer3_outputs(7821)) or (layer3_outputs(4658));
    layer4_outputs(7846) <= (layer3_outputs(7968)) xor (layer3_outputs(3945));
    layer4_outputs(7847) <= not(layer3_outputs(2291));
    layer4_outputs(7848) <= (layer3_outputs(8560)) or (layer3_outputs(1849));
    layer4_outputs(7849) <= (layer3_outputs(3820)) and (layer3_outputs(4900));
    layer4_outputs(7850) <= layer3_outputs(6211);
    layer4_outputs(7851) <= not(layer3_outputs(3728));
    layer4_outputs(7852) <= not((layer3_outputs(4671)) or (layer3_outputs(2322)));
    layer4_outputs(7853) <= layer3_outputs(6586);
    layer4_outputs(7854) <= layer3_outputs(5290);
    layer4_outputs(7855) <= layer3_outputs(2686);
    layer4_outputs(7856) <= layer3_outputs(4518);
    layer4_outputs(7857) <= (layer3_outputs(3434)) and not (layer3_outputs(5817));
    layer4_outputs(7858) <= (layer3_outputs(1563)) and not (layer3_outputs(486));
    layer4_outputs(7859) <= not(layer3_outputs(9825));
    layer4_outputs(7860) <= not(layer3_outputs(9363)) or (layer3_outputs(3139));
    layer4_outputs(7861) <= not(layer3_outputs(7547));
    layer4_outputs(7862) <= layer3_outputs(4);
    layer4_outputs(7863) <= not((layer3_outputs(3747)) xor (layer3_outputs(9590)));
    layer4_outputs(7864) <= (layer3_outputs(6378)) xor (layer3_outputs(2480));
    layer4_outputs(7865) <= layer3_outputs(1211);
    layer4_outputs(7866) <= layer3_outputs(3215);
    layer4_outputs(7867) <= not(layer3_outputs(3467));
    layer4_outputs(7868) <= (layer3_outputs(6520)) or (layer3_outputs(4590));
    layer4_outputs(7869) <= layer3_outputs(5301);
    layer4_outputs(7870) <= (layer3_outputs(3248)) xor (layer3_outputs(3023));
    layer4_outputs(7871) <= (layer3_outputs(3404)) and (layer3_outputs(954));
    layer4_outputs(7872) <= not(layer3_outputs(166));
    layer4_outputs(7873) <= layer3_outputs(21);
    layer4_outputs(7874) <= not((layer3_outputs(7438)) or (layer3_outputs(4577)));
    layer4_outputs(7875) <= not((layer3_outputs(5292)) xor (layer3_outputs(8888)));
    layer4_outputs(7876) <= not(layer3_outputs(5914));
    layer4_outputs(7877) <= not((layer3_outputs(7161)) xor (layer3_outputs(8099)));
    layer4_outputs(7878) <= (layer3_outputs(4269)) and not (layer3_outputs(2376));
    layer4_outputs(7879) <= (layer3_outputs(8756)) and not (layer3_outputs(1850));
    layer4_outputs(7880) <= layer3_outputs(5329);
    layer4_outputs(7881) <= (layer3_outputs(1773)) xor (layer3_outputs(6972));
    layer4_outputs(7882) <= (layer3_outputs(3944)) xor (layer3_outputs(8800));
    layer4_outputs(7883) <= layer3_outputs(5099);
    layer4_outputs(7884) <= layer3_outputs(67);
    layer4_outputs(7885) <= not((layer3_outputs(8362)) or (layer3_outputs(7836)));
    layer4_outputs(7886) <= layer3_outputs(5333);
    layer4_outputs(7887) <= layer3_outputs(190);
    layer4_outputs(7888) <= not((layer3_outputs(8423)) xor (layer3_outputs(5344)));
    layer4_outputs(7889) <= not((layer3_outputs(7500)) xor (layer3_outputs(9545)));
    layer4_outputs(7890) <= (layer3_outputs(3727)) and not (layer3_outputs(4499));
    layer4_outputs(7891) <= layer3_outputs(6950);
    layer4_outputs(7892) <= (layer3_outputs(6395)) or (layer3_outputs(1027));
    layer4_outputs(7893) <= not((layer3_outputs(7764)) and (layer3_outputs(4047)));
    layer4_outputs(7894) <= not(layer3_outputs(2515));
    layer4_outputs(7895) <= not((layer3_outputs(7098)) xor (layer3_outputs(5589)));
    layer4_outputs(7896) <= (layer3_outputs(8559)) or (layer3_outputs(5347));
    layer4_outputs(7897) <= (layer3_outputs(297)) and not (layer3_outputs(3750));
    layer4_outputs(7898) <= layer3_outputs(3001);
    layer4_outputs(7899) <= (layer3_outputs(8790)) and not (layer3_outputs(2824));
    layer4_outputs(7900) <= not((layer3_outputs(8158)) and (layer3_outputs(2705)));
    layer4_outputs(7901) <= not(layer3_outputs(9254));
    layer4_outputs(7902) <= (layer3_outputs(5508)) and (layer3_outputs(8142));
    layer4_outputs(7903) <= not((layer3_outputs(1095)) and (layer3_outputs(7944)));
    layer4_outputs(7904) <= not(layer3_outputs(8767));
    layer4_outputs(7905) <= layer3_outputs(8019);
    layer4_outputs(7906) <= not(layer3_outputs(5209));
    layer4_outputs(7907) <= not(layer3_outputs(6075)) or (layer3_outputs(8896));
    layer4_outputs(7908) <= not((layer3_outputs(4463)) or (layer3_outputs(3891)));
    layer4_outputs(7909) <= layer3_outputs(1920);
    layer4_outputs(7910) <= not(layer3_outputs(5879)) or (layer3_outputs(4298));
    layer4_outputs(7911) <= not(layer3_outputs(7739));
    layer4_outputs(7912) <= layer3_outputs(2463);
    layer4_outputs(7913) <= (layer3_outputs(304)) xor (layer3_outputs(8054));
    layer4_outputs(7914) <= (layer3_outputs(7322)) and not (layer3_outputs(4510));
    layer4_outputs(7915) <= not((layer3_outputs(3373)) or (layer3_outputs(9046)));
    layer4_outputs(7916) <= layer3_outputs(8379);
    layer4_outputs(7917) <= (layer3_outputs(8682)) and not (layer3_outputs(4722));
    layer4_outputs(7918) <= layer3_outputs(3498);
    layer4_outputs(7919) <= not(layer3_outputs(487));
    layer4_outputs(7920) <= not((layer3_outputs(3444)) xor (layer3_outputs(2150)));
    layer4_outputs(7921) <= layer3_outputs(973);
    layer4_outputs(7922) <= not((layer3_outputs(3876)) xor (layer3_outputs(9577)));
    layer4_outputs(7923) <= not(layer3_outputs(5516)) or (layer3_outputs(3771));
    layer4_outputs(7924) <= not((layer3_outputs(6788)) xor (layer3_outputs(150)));
    layer4_outputs(7925) <= not((layer3_outputs(3184)) or (layer3_outputs(5662)));
    layer4_outputs(7926) <= not(layer3_outputs(7983));
    layer4_outputs(7927) <= not((layer3_outputs(2717)) xor (layer3_outputs(6767)));
    layer4_outputs(7928) <= layer3_outputs(8924);
    layer4_outputs(7929) <= layer3_outputs(6920);
    layer4_outputs(7930) <= not((layer3_outputs(9939)) and (layer3_outputs(8445)));
    layer4_outputs(7931) <= not(layer3_outputs(6354));
    layer4_outputs(7932) <= layer3_outputs(1869);
    layer4_outputs(7933) <= layer3_outputs(8896);
    layer4_outputs(7934) <= not(layer3_outputs(10032));
    layer4_outputs(7935) <= (layer3_outputs(2111)) xor (layer3_outputs(9211));
    layer4_outputs(7936) <= (layer3_outputs(4103)) xor (layer3_outputs(2467));
    layer4_outputs(7937) <= layer3_outputs(6026);
    layer4_outputs(7938) <= not((layer3_outputs(7527)) xor (layer3_outputs(6069)));
    layer4_outputs(7939) <= (layer3_outputs(8057)) xor (layer3_outputs(1657));
    layer4_outputs(7940) <= (layer3_outputs(498)) and (layer3_outputs(2020));
    layer4_outputs(7941) <= not(layer3_outputs(1540));
    layer4_outputs(7942) <= not(layer3_outputs(8426));
    layer4_outputs(7943) <= not(layer3_outputs(2017));
    layer4_outputs(7944) <= not(layer3_outputs(3722));
    layer4_outputs(7945) <= (layer3_outputs(3309)) and not (layer3_outputs(7402));
    layer4_outputs(7946) <= not(layer3_outputs(2167)) or (layer3_outputs(3043));
    layer4_outputs(7947) <= (layer3_outputs(5787)) and (layer3_outputs(9928));
    layer4_outputs(7948) <= layer3_outputs(306);
    layer4_outputs(7949) <= layer3_outputs(4096);
    layer4_outputs(7950) <= not((layer3_outputs(3896)) xor (layer3_outputs(2436)));
    layer4_outputs(7951) <= layer3_outputs(5603);
    layer4_outputs(7952) <= (layer3_outputs(231)) and not (layer3_outputs(5338));
    layer4_outputs(7953) <= not((layer3_outputs(2129)) and (layer3_outputs(10015)));
    layer4_outputs(7954) <= not(layer3_outputs(3612));
    layer4_outputs(7955) <= layer3_outputs(5827);
    layer4_outputs(7956) <= not((layer3_outputs(10218)) or (layer3_outputs(8705)));
    layer4_outputs(7957) <= layer3_outputs(4244);
    layer4_outputs(7958) <= not(layer3_outputs(1957));
    layer4_outputs(7959) <= not(layer3_outputs(3840));
    layer4_outputs(7960) <= (layer3_outputs(5350)) and not (layer3_outputs(6183));
    layer4_outputs(7961) <= (layer3_outputs(4609)) or (layer3_outputs(5782));
    layer4_outputs(7962) <= layer3_outputs(7230);
    layer4_outputs(7963) <= layer3_outputs(9513);
    layer4_outputs(7964) <= not(layer3_outputs(4851));
    layer4_outputs(7965) <= not(layer3_outputs(9466)) or (layer3_outputs(9533));
    layer4_outputs(7966) <= layer3_outputs(309);
    layer4_outputs(7967) <= not(layer3_outputs(2988));
    layer4_outputs(7968) <= not((layer3_outputs(9815)) and (layer3_outputs(10102)));
    layer4_outputs(7969) <= (layer3_outputs(9334)) xor (layer3_outputs(1577));
    layer4_outputs(7970) <= not(layer3_outputs(2545));
    layer4_outputs(7971) <= '1';
    layer4_outputs(7972) <= not(layer3_outputs(92));
    layer4_outputs(7973) <= not(layer3_outputs(9176));
    layer4_outputs(7974) <= not(layer3_outputs(5894));
    layer4_outputs(7975) <= not(layer3_outputs(9133));
    layer4_outputs(7976) <= '1';
    layer4_outputs(7977) <= not(layer3_outputs(5421));
    layer4_outputs(7978) <= not(layer3_outputs(1644));
    layer4_outputs(7979) <= not((layer3_outputs(2457)) xor (layer3_outputs(7949)));
    layer4_outputs(7980) <= (layer3_outputs(1029)) xor (layer3_outputs(7148));
    layer4_outputs(7981) <= (layer3_outputs(6244)) and not (layer3_outputs(6022));
    layer4_outputs(7982) <= layer3_outputs(8193);
    layer4_outputs(7983) <= not(layer3_outputs(8212));
    layer4_outputs(7984) <= layer3_outputs(4208);
    layer4_outputs(7985) <= not((layer3_outputs(6107)) or (layer3_outputs(8571)));
    layer4_outputs(7986) <= not(layer3_outputs(3611));
    layer4_outputs(7987) <= not(layer3_outputs(3749)) or (layer3_outputs(7236));
    layer4_outputs(7988) <= not(layer3_outputs(3045));
    layer4_outputs(7989) <= (layer3_outputs(7293)) and not (layer3_outputs(8335));
    layer4_outputs(7990) <= layer3_outputs(6450);
    layer4_outputs(7991) <= not(layer3_outputs(5476));
    layer4_outputs(7992) <= '0';
    layer4_outputs(7993) <= layer3_outputs(7240);
    layer4_outputs(7994) <= not((layer3_outputs(8029)) or (layer3_outputs(4274)));
    layer4_outputs(7995) <= layer3_outputs(7645);
    layer4_outputs(7996) <= layer3_outputs(7090);
    layer4_outputs(7997) <= layer3_outputs(2971);
    layer4_outputs(7998) <= not(layer3_outputs(8688));
    layer4_outputs(7999) <= not(layer3_outputs(9884));
    layer4_outputs(8000) <= not(layer3_outputs(1338));
    layer4_outputs(8001) <= '0';
    layer4_outputs(8002) <= (layer3_outputs(3265)) xor (layer3_outputs(8630));
    layer4_outputs(8003) <= layer3_outputs(7573);
    layer4_outputs(8004) <= not(layer3_outputs(531));
    layer4_outputs(8005) <= not(layer3_outputs(7263));
    layer4_outputs(8006) <= (layer3_outputs(545)) xor (layer3_outputs(9176));
    layer4_outputs(8007) <= layer3_outputs(1159);
    layer4_outputs(8008) <= layer3_outputs(686);
    layer4_outputs(8009) <= not((layer3_outputs(2259)) and (layer3_outputs(6798)));
    layer4_outputs(8010) <= not(layer3_outputs(5003));
    layer4_outputs(8011) <= (layer3_outputs(4328)) xor (layer3_outputs(6345));
    layer4_outputs(8012) <= layer3_outputs(2447);
    layer4_outputs(8013) <= (layer3_outputs(904)) and not (layer3_outputs(6638));
    layer4_outputs(8014) <= (layer3_outputs(2110)) and not (layer3_outputs(2008));
    layer4_outputs(8015) <= not(layer3_outputs(8575));
    layer4_outputs(8016) <= layer3_outputs(10191);
    layer4_outputs(8017) <= not(layer3_outputs(1682));
    layer4_outputs(8018) <= layer3_outputs(785);
    layer4_outputs(8019) <= not((layer3_outputs(726)) and (layer3_outputs(2866)));
    layer4_outputs(8020) <= (layer3_outputs(8508)) xor (layer3_outputs(360));
    layer4_outputs(8021) <= not((layer3_outputs(9942)) and (layer3_outputs(4999)));
    layer4_outputs(8022) <= (layer3_outputs(2141)) or (layer3_outputs(7480));
    layer4_outputs(8023) <= not(layer3_outputs(3143));
    layer4_outputs(8024) <= not(layer3_outputs(9262));
    layer4_outputs(8025) <= not(layer3_outputs(463));
    layer4_outputs(8026) <= layer3_outputs(1980);
    layer4_outputs(8027) <= not(layer3_outputs(3519)) or (layer3_outputs(228));
    layer4_outputs(8028) <= (layer3_outputs(5917)) xor (layer3_outputs(5619));
    layer4_outputs(8029) <= not(layer3_outputs(6276));
    layer4_outputs(8030) <= layer3_outputs(6587);
    layer4_outputs(8031) <= layer3_outputs(7207);
    layer4_outputs(8032) <= not(layer3_outputs(4959));
    layer4_outputs(8033) <= layer3_outputs(4581);
    layer4_outputs(8034) <= not(layer3_outputs(1324));
    layer4_outputs(8035) <= (layer3_outputs(263)) and not (layer3_outputs(3862));
    layer4_outputs(8036) <= layer3_outputs(9649);
    layer4_outputs(8037) <= not((layer3_outputs(4594)) or (layer3_outputs(4260)));
    layer4_outputs(8038) <= not(layer3_outputs(2332));
    layer4_outputs(8039) <= not(layer3_outputs(2391));
    layer4_outputs(8040) <= not(layer3_outputs(3797));
    layer4_outputs(8041) <= layer3_outputs(28);
    layer4_outputs(8042) <= not((layer3_outputs(4056)) xor (layer3_outputs(2877)));
    layer4_outputs(8043) <= not(layer3_outputs(8660));
    layer4_outputs(8044) <= not(layer3_outputs(6353));
    layer4_outputs(8045) <= layer3_outputs(7731);
    layer4_outputs(8046) <= not((layer3_outputs(4184)) and (layer3_outputs(2938)));
    layer4_outputs(8047) <= not(layer3_outputs(8112));
    layer4_outputs(8048) <= (layer3_outputs(3530)) and not (layer3_outputs(7418));
    layer4_outputs(8049) <= (layer3_outputs(9809)) xor (layer3_outputs(1473));
    layer4_outputs(8050) <= not(layer3_outputs(4442));
    layer4_outputs(8051) <= layer3_outputs(8125);
    layer4_outputs(8052) <= not(layer3_outputs(6650)) or (layer3_outputs(3630));
    layer4_outputs(8053) <= not((layer3_outputs(5433)) xor (layer3_outputs(7956)));
    layer4_outputs(8054) <= (layer3_outputs(8647)) and not (layer3_outputs(8707));
    layer4_outputs(8055) <= not(layer3_outputs(8366));
    layer4_outputs(8056) <= not(layer3_outputs(4362));
    layer4_outputs(8057) <= (layer3_outputs(4431)) xor (layer3_outputs(9705));
    layer4_outputs(8058) <= layer3_outputs(2216);
    layer4_outputs(8059) <= (layer3_outputs(921)) and not (layer3_outputs(2981));
    layer4_outputs(8060) <= not(layer3_outputs(6362)) or (layer3_outputs(9198));
    layer4_outputs(8061) <= not(layer3_outputs(1230));
    layer4_outputs(8062) <= not(layer3_outputs(6893)) or (layer3_outputs(875));
    layer4_outputs(8063) <= not(layer3_outputs(34));
    layer4_outputs(8064) <= not(layer3_outputs(6700)) or (layer3_outputs(4633));
    layer4_outputs(8065) <= layer3_outputs(1659);
    layer4_outputs(8066) <= not(layer3_outputs(1515));
    layer4_outputs(8067) <= not((layer3_outputs(7165)) and (layer3_outputs(3142)));
    layer4_outputs(8068) <= layer3_outputs(9011);
    layer4_outputs(8069) <= layer3_outputs(7029);
    layer4_outputs(8070) <= (layer3_outputs(5136)) or (layer3_outputs(3197));
    layer4_outputs(8071) <= (layer3_outputs(1531)) and not (layer3_outputs(1288));
    layer4_outputs(8072) <= not(layer3_outputs(1514));
    layer4_outputs(8073) <= not(layer3_outputs(4604));
    layer4_outputs(8074) <= layer3_outputs(7422);
    layer4_outputs(8075) <= (layer3_outputs(1940)) and not (layer3_outputs(9084));
    layer4_outputs(8076) <= not((layer3_outputs(5987)) xor (layer3_outputs(71)));
    layer4_outputs(8077) <= not(layer3_outputs(3781));
    layer4_outputs(8078) <= not(layer3_outputs(2691));
    layer4_outputs(8079) <= not((layer3_outputs(3387)) xor (layer3_outputs(9971)));
    layer4_outputs(8080) <= not(layer3_outputs(7575));
    layer4_outputs(8081) <= not(layer3_outputs(8204));
    layer4_outputs(8082) <= layer3_outputs(405);
    layer4_outputs(8083) <= not(layer3_outputs(9499)) or (layer3_outputs(9688));
    layer4_outputs(8084) <= layer3_outputs(3017);
    layer4_outputs(8085) <= not(layer3_outputs(3787));
    layer4_outputs(8086) <= not((layer3_outputs(5938)) xor (layer3_outputs(2048)));
    layer4_outputs(8087) <= (layer3_outputs(55)) and not (layer3_outputs(3142));
    layer4_outputs(8088) <= not((layer3_outputs(472)) xor (layer3_outputs(4680)));
    layer4_outputs(8089) <= (layer3_outputs(5205)) xor (layer3_outputs(1459));
    layer4_outputs(8090) <= not((layer3_outputs(5641)) xor (layer3_outputs(8907)));
    layer4_outputs(8091) <= (layer3_outputs(1746)) xor (layer3_outputs(9550));
    layer4_outputs(8092) <= layer3_outputs(7428);
    layer4_outputs(8093) <= layer3_outputs(1946);
    layer4_outputs(8094) <= not(layer3_outputs(10008));
    layer4_outputs(8095) <= not(layer3_outputs(3421));
    layer4_outputs(8096) <= not(layer3_outputs(5439));
    layer4_outputs(8097) <= layer3_outputs(5532);
    layer4_outputs(8098) <= not(layer3_outputs(9845));
    layer4_outputs(8099) <= (layer3_outputs(7041)) and not (layer3_outputs(3441));
    layer4_outputs(8100) <= (layer3_outputs(1430)) or (layer3_outputs(391));
    layer4_outputs(8101) <= not((layer3_outputs(3231)) and (layer3_outputs(7366)));
    layer4_outputs(8102) <= not(layer3_outputs(172)) or (layer3_outputs(4487));
    layer4_outputs(8103) <= layer3_outputs(10042);
    layer4_outputs(8104) <= not((layer3_outputs(7560)) xor (layer3_outputs(5796)));
    layer4_outputs(8105) <= (layer3_outputs(2857)) and not (layer3_outputs(4410));
    layer4_outputs(8106) <= '1';
    layer4_outputs(8107) <= not(layer3_outputs(1841));
    layer4_outputs(8108) <= layer3_outputs(1022);
    layer4_outputs(8109) <= layer3_outputs(3153);
    layer4_outputs(8110) <= layer3_outputs(4201);
    layer4_outputs(8111) <= layer3_outputs(5233);
    layer4_outputs(8112) <= (layer3_outputs(5704)) and not (layer3_outputs(4375));
    layer4_outputs(8113) <= (layer3_outputs(9632)) and not (layer3_outputs(2722));
    layer4_outputs(8114) <= layer3_outputs(7447);
    layer4_outputs(8115) <= not(layer3_outputs(5566)) or (layer3_outputs(1455));
    layer4_outputs(8116) <= layer3_outputs(8598);
    layer4_outputs(8117) <= not((layer3_outputs(5451)) xor (layer3_outputs(9337)));
    layer4_outputs(8118) <= layer3_outputs(5627);
    layer4_outputs(8119) <= not((layer3_outputs(2564)) or (layer3_outputs(4579)));
    layer4_outputs(8120) <= layer3_outputs(3167);
    layer4_outputs(8121) <= layer3_outputs(1002);
    layer4_outputs(8122) <= layer3_outputs(8074);
    layer4_outputs(8123) <= not((layer3_outputs(1611)) xor (layer3_outputs(3126)));
    layer4_outputs(8124) <= not(layer3_outputs(2386));
    layer4_outputs(8125) <= not(layer3_outputs(6964));
    layer4_outputs(8126) <= not(layer3_outputs(1609));
    layer4_outputs(8127) <= (layer3_outputs(1687)) and not (layer3_outputs(1478));
    layer4_outputs(8128) <= layer3_outputs(4856);
    layer4_outputs(8129) <= not((layer3_outputs(7335)) or (layer3_outputs(4476)));
    layer4_outputs(8130) <= not(layer3_outputs(8359));
    layer4_outputs(8131) <= not(layer3_outputs(3287));
    layer4_outputs(8132) <= (layer3_outputs(1017)) xor (layer3_outputs(2829));
    layer4_outputs(8133) <= not(layer3_outputs(9185));
    layer4_outputs(8134) <= not(layer3_outputs(6428));
    layer4_outputs(8135) <= not((layer3_outputs(4817)) xor (layer3_outputs(6630)));
    layer4_outputs(8136) <= not((layer3_outputs(6923)) xor (layer3_outputs(9130)));
    layer4_outputs(8137) <= layer3_outputs(7607);
    layer4_outputs(8138) <= not(layer3_outputs(8678)) or (layer3_outputs(8043));
    layer4_outputs(8139) <= layer3_outputs(9422);
    layer4_outputs(8140) <= not((layer3_outputs(3258)) or (layer3_outputs(205)));
    layer4_outputs(8141) <= not(layer3_outputs(6858)) or (layer3_outputs(5556));
    layer4_outputs(8142) <= not((layer3_outputs(5914)) xor (layer3_outputs(148)));
    layer4_outputs(8143) <= layer3_outputs(7937);
    layer4_outputs(8144) <= layer3_outputs(5836);
    layer4_outputs(8145) <= not(layer3_outputs(10073));
    layer4_outputs(8146) <= not((layer3_outputs(3921)) and (layer3_outputs(5636)));
    layer4_outputs(8147) <= layer3_outputs(3556);
    layer4_outputs(8148) <= not(layer3_outputs(4340));
    layer4_outputs(8149) <= (layer3_outputs(8842)) and not (layer3_outputs(3191));
    layer4_outputs(8150) <= not(layer3_outputs(5352));
    layer4_outputs(8151) <= not(layer3_outputs(1472));
    layer4_outputs(8152) <= (layer3_outputs(3544)) xor (layer3_outputs(6910));
    layer4_outputs(8153) <= layer3_outputs(4700);
    layer4_outputs(8154) <= not(layer3_outputs(5738));
    layer4_outputs(8155) <= layer3_outputs(7118);
    layer4_outputs(8156) <= layer3_outputs(3865);
    layer4_outputs(8157) <= layer3_outputs(5912);
    layer4_outputs(8158) <= not(layer3_outputs(7357)) or (layer3_outputs(4316));
    layer4_outputs(8159) <= layer3_outputs(8887);
    layer4_outputs(8160) <= '1';
    layer4_outputs(8161) <= not(layer3_outputs(6605));
    layer4_outputs(8162) <= not(layer3_outputs(3587));
    layer4_outputs(8163) <= not(layer3_outputs(968));
    layer4_outputs(8164) <= not((layer3_outputs(8806)) and (layer3_outputs(3266)));
    layer4_outputs(8165) <= not((layer3_outputs(1424)) xor (layer3_outputs(132)));
    layer4_outputs(8166) <= layer3_outputs(8795);
    layer4_outputs(8167) <= not(layer3_outputs(6955));
    layer4_outputs(8168) <= layer3_outputs(5482);
    layer4_outputs(8169) <= layer3_outputs(2124);
    layer4_outputs(8170) <= not((layer3_outputs(7032)) xor (layer3_outputs(7897)));
    layer4_outputs(8171) <= not((layer3_outputs(2914)) xor (layer3_outputs(9659)));
    layer4_outputs(8172) <= layer3_outputs(8046);
    layer4_outputs(8173) <= (layer3_outputs(7680)) and (layer3_outputs(6443));
    layer4_outputs(8174) <= layer3_outputs(730);
    layer4_outputs(8175) <= (layer3_outputs(153)) and not (layer3_outputs(5757));
    layer4_outputs(8176) <= layer3_outputs(4978);
    layer4_outputs(8177) <= layer3_outputs(4175);
    layer4_outputs(8178) <= layer3_outputs(8247);
    layer4_outputs(8179) <= not((layer3_outputs(9750)) or (layer3_outputs(7320)));
    layer4_outputs(8180) <= (layer3_outputs(2635)) xor (layer3_outputs(4659));
    layer4_outputs(8181) <= not(layer3_outputs(3952));
    layer4_outputs(8182) <= not(layer3_outputs(4208));
    layer4_outputs(8183) <= layer3_outputs(1139);
    layer4_outputs(8184) <= (layer3_outputs(5551)) and not (layer3_outputs(6233));
    layer4_outputs(8185) <= not((layer3_outputs(6607)) and (layer3_outputs(7177)));
    layer4_outputs(8186) <= not(layer3_outputs(3286)) or (layer3_outputs(4171));
    layer4_outputs(8187) <= not(layer3_outputs(9391));
    layer4_outputs(8188) <= (layer3_outputs(8080)) or (layer3_outputs(10091));
    layer4_outputs(8189) <= (layer3_outputs(6694)) or (layer3_outputs(2246));
    layer4_outputs(8190) <= not(layer3_outputs(8876));
    layer4_outputs(8191) <= (layer3_outputs(2574)) and not (layer3_outputs(4735));
    layer4_outputs(8192) <= not(layer3_outputs(3337));
    layer4_outputs(8193) <= layer3_outputs(622);
    layer4_outputs(8194) <= layer3_outputs(10057);
    layer4_outputs(8195) <= layer3_outputs(1984);
    layer4_outputs(8196) <= layer3_outputs(10171);
    layer4_outputs(8197) <= not(layer3_outputs(5044));
    layer4_outputs(8198) <= layer3_outputs(6606);
    layer4_outputs(8199) <= (layer3_outputs(9330)) xor (layer3_outputs(1963));
    layer4_outputs(8200) <= (layer3_outputs(7354)) xor (layer3_outputs(7524));
    layer4_outputs(8201) <= not((layer3_outputs(2093)) xor (layer3_outputs(7899)));
    layer4_outputs(8202) <= not(layer3_outputs(7086));
    layer4_outputs(8203) <= layer3_outputs(3144);
    layer4_outputs(8204) <= not((layer3_outputs(2418)) and (layer3_outputs(9208)));
    layer4_outputs(8205) <= not(layer3_outputs(4026)) or (layer3_outputs(5924));
    layer4_outputs(8206) <= not(layer3_outputs(1991));
    layer4_outputs(8207) <= (layer3_outputs(2183)) and not (layer3_outputs(1722));
    layer4_outputs(8208) <= layer3_outputs(4033);
    layer4_outputs(8209) <= layer3_outputs(1539);
    layer4_outputs(8210) <= (layer3_outputs(10188)) or (layer3_outputs(2066));
    layer4_outputs(8211) <= not(layer3_outputs(7813));
    layer4_outputs(8212) <= not(layer3_outputs(4564)) or (layer3_outputs(1492));
    layer4_outputs(8213) <= not(layer3_outputs(182));
    layer4_outputs(8214) <= (layer3_outputs(7399)) and (layer3_outputs(9756));
    layer4_outputs(8215) <= (layer3_outputs(1286)) and not (layer3_outputs(4106));
    layer4_outputs(8216) <= (layer3_outputs(9168)) and not (layer3_outputs(3681));
    layer4_outputs(8217) <= not(layer3_outputs(1371));
    layer4_outputs(8218) <= (layer3_outputs(3729)) or (layer3_outputs(6319));
    layer4_outputs(8219) <= not(layer3_outputs(7901)) or (layer3_outputs(3214));
    layer4_outputs(8220) <= not(layer3_outputs(7799));
    layer4_outputs(8221) <= layer3_outputs(2697);
    layer4_outputs(8222) <= not((layer3_outputs(5097)) xor (layer3_outputs(9916)));
    layer4_outputs(8223) <= (layer3_outputs(2031)) and (layer3_outputs(8310));
    layer4_outputs(8224) <= not(layer3_outputs(8676));
    layer4_outputs(8225) <= (layer3_outputs(3417)) xor (layer3_outputs(7984));
    layer4_outputs(8226) <= (layer3_outputs(9328)) xor (layer3_outputs(8132));
    layer4_outputs(8227) <= not(layer3_outputs(3432));
    layer4_outputs(8228) <= layer3_outputs(2955);
    layer4_outputs(8229) <= not(layer3_outputs(1694));
    layer4_outputs(8230) <= layer3_outputs(8250);
    layer4_outputs(8231) <= layer3_outputs(9823);
    layer4_outputs(8232) <= (layer3_outputs(3648)) and not (layer3_outputs(5564));
    layer4_outputs(8233) <= not(layer3_outputs(9453));
    layer4_outputs(8234) <= not((layer3_outputs(331)) xor (layer3_outputs(730)));
    layer4_outputs(8235) <= not(layer3_outputs(33)) or (layer3_outputs(6604));
    layer4_outputs(8236) <= (layer3_outputs(9829)) and (layer3_outputs(311));
    layer4_outputs(8237) <= not(layer3_outputs(6106));
    layer4_outputs(8238) <= not(layer3_outputs(5818));
    layer4_outputs(8239) <= layer3_outputs(1360);
    layer4_outputs(8240) <= not(layer3_outputs(79));
    layer4_outputs(8241) <= layer3_outputs(7890);
    layer4_outputs(8242) <= (layer3_outputs(6292)) or (layer3_outputs(3038));
    layer4_outputs(8243) <= layer3_outputs(9949);
    layer4_outputs(8244) <= not(layer3_outputs(9275));
    layer4_outputs(8245) <= layer3_outputs(5074);
    layer4_outputs(8246) <= not(layer3_outputs(858));
    layer4_outputs(8247) <= layer3_outputs(5075);
    layer4_outputs(8248) <= not(layer3_outputs(8474));
    layer4_outputs(8249) <= (layer3_outputs(5869)) xor (layer3_outputs(3558));
    layer4_outputs(8250) <= not(layer3_outputs(2962));
    layer4_outputs(8251) <= (layer3_outputs(3953)) and not (layer3_outputs(10037));
    layer4_outputs(8252) <= not(layer3_outputs(8548));
    layer4_outputs(8253) <= not(layer3_outputs(6291));
    layer4_outputs(8254) <= layer3_outputs(9700);
    layer4_outputs(8255) <= not(layer3_outputs(6934)) or (layer3_outputs(2985));
    layer4_outputs(8256) <= layer3_outputs(1279);
    layer4_outputs(8257) <= not(layer3_outputs(205));
    layer4_outputs(8258) <= not(layer3_outputs(8722));
    layer4_outputs(8259) <= not(layer3_outputs(5632));
    layer4_outputs(8260) <= not((layer3_outputs(3458)) and (layer3_outputs(5576)));
    layer4_outputs(8261) <= not(layer3_outputs(3720));
    layer4_outputs(8262) <= not(layer3_outputs(7751)) or (layer3_outputs(9020));
    layer4_outputs(8263) <= layer3_outputs(8076);
    layer4_outputs(8264) <= (layer3_outputs(4593)) or (layer3_outputs(5681));
    layer4_outputs(8265) <= layer3_outputs(280);
    layer4_outputs(8266) <= (layer3_outputs(7640)) xor (layer3_outputs(6480));
    layer4_outputs(8267) <= not(layer3_outputs(7815));
    layer4_outputs(8268) <= layer3_outputs(8134);
    layer4_outputs(8269) <= not(layer3_outputs(9973));
    layer4_outputs(8270) <= (layer3_outputs(2967)) xor (layer3_outputs(251));
    layer4_outputs(8271) <= (layer3_outputs(775)) xor (layer3_outputs(303));
    layer4_outputs(8272) <= '1';
    layer4_outputs(8273) <= layer3_outputs(5997);
    layer4_outputs(8274) <= layer3_outputs(1569);
    layer4_outputs(8275) <= (layer3_outputs(202)) xor (layer3_outputs(3342));
    layer4_outputs(8276) <= layer3_outputs(7266);
    layer4_outputs(8277) <= (layer3_outputs(9925)) and not (layer3_outputs(3178));
    layer4_outputs(8278) <= (layer3_outputs(7316)) xor (layer3_outputs(1635));
    layer4_outputs(8279) <= (layer3_outputs(5018)) and not (layer3_outputs(3524));
    layer4_outputs(8280) <= layer3_outputs(4280);
    layer4_outputs(8281) <= not((layer3_outputs(9248)) or (layer3_outputs(8502)));
    layer4_outputs(8282) <= not(layer3_outputs(4776));
    layer4_outputs(8283) <= not(layer3_outputs(235));
    layer4_outputs(8284) <= layer3_outputs(6855);
    layer4_outputs(8285) <= (layer3_outputs(5803)) and not (layer3_outputs(4579));
    layer4_outputs(8286) <= not(layer3_outputs(6886)) or (layer3_outputs(6425));
    layer4_outputs(8287) <= not(layer3_outputs(4232));
    layer4_outputs(8288) <= layer3_outputs(4416);
    layer4_outputs(8289) <= '0';
    layer4_outputs(8290) <= not((layer3_outputs(175)) xor (layer3_outputs(6847)));
    layer4_outputs(8291) <= not(layer3_outputs(2974));
    layer4_outputs(8292) <= layer3_outputs(7201);
    layer4_outputs(8293) <= (layer3_outputs(3773)) and not (layer3_outputs(5197));
    layer4_outputs(8294) <= not(layer3_outputs(7380));
    layer4_outputs(8295) <= layer3_outputs(1767);
    layer4_outputs(8296) <= not((layer3_outputs(2977)) and (layer3_outputs(7221)));
    layer4_outputs(8297) <= (layer3_outputs(2210)) xor (layer3_outputs(6480));
    layer4_outputs(8298) <= not(layer3_outputs(9888));
    layer4_outputs(8299) <= not((layer3_outputs(455)) xor (layer3_outputs(7056)));
    layer4_outputs(8300) <= not(layer3_outputs(6160));
    layer4_outputs(8301) <= not(layer3_outputs(6048));
    layer4_outputs(8302) <= layer3_outputs(1770);
    layer4_outputs(8303) <= layer3_outputs(8342);
    layer4_outputs(8304) <= not(layer3_outputs(2643));
    layer4_outputs(8305) <= (layer3_outputs(4873)) xor (layer3_outputs(4401));
    layer4_outputs(8306) <= (layer3_outputs(8064)) or (layer3_outputs(5127));
    layer4_outputs(8307) <= not(layer3_outputs(2411));
    layer4_outputs(8308) <= not((layer3_outputs(280)) and (layer3_outputs(8839)));
    layer4_outputs(8309) <= layer3_outputs(9424);
    layer4_outputs(8310) <= layer3_outputs(2408);
    layer4_outputs(8311) <= not((layer3_outputs(2967)) and (layer3_outputs(8963)));
    layer4_outputs(8312) <= not((layer3_outputs(4397)) xor (layer3_outputs(4359)));
    layer4_outputs(8313) <= not((layer3_outputs(9745)) xor (layer3_outputs(4243)));
    layer4_outputs(8314) <= not(layer3_outputs(4062));
    layer4_outputs(8315) <= not(layer3_outputs(8568));
    layer4_outputs(8316) <= not(layer3_outputs(2373));
    layer4_outputs(8317) <= '0';
    layer4_outputs(8318) <= not(layer3_outputs(4128));
    layer4_outputs(8319) <= not(layer3_outputs(694));
    layer4_outputs(8320) <= layer3_outputs(4423);
    layer4_outputs(8321) <= (layer3_outputs(10018)) xor (layer3_outputs(9588));
    layer4_outputs(8322) <= not((layer3_outputs(2326)) xor (layer3_outputs(3384)));
    layer4_outputs(8323) <= not(layer3_outputs(9129)) or (layer3_outputs(6095));
    layer4_outputs(8324) <= layer3_outputs(7016);
    layer4_outputs(8325) <= (layer3_outputs(8850)) and not (layer3_outputs(4108));
    layer4_outputs(8326) <= layer3_outputs(7790);
    layer4_outputs(8327) <= layer3_outputs(9186);
    layer4_outputs(8328) <= layer3_outputs(9137);
    layer4_outputs(8329) <= (layer3_outputs(5507)) xor (layer3_outputs(944));
    layer4_outputs(8330) <= not(layer3_outputs(488));
    layer4_outputs(8331) <= layer3_outputs(5123);
    layer4_outputs(8332) <= not(layer3_outputs(477)) or (layer3_outputs(2580));
    layer4_outputs(8333) <= not(layer3_outputs(5689));
    layer4_outputs(8334) <= not(layer3_outputs(553)) or (layer3_outputs(2452));
    layer4_outputs(8335) <= not(layer3_outputs(9840)) or (layer3_outputs(5950));
    layer4_outputs(8336) <= (layer3_outputs(8596)) and not (layer3_outputs(24));
    layer4_outputs(8337) <= not(layer3_outputs(9522));
    layer4_outputs(8338) <= not(layer3_outputs(7319));
    layer4_outputs(8339) <= layer3_outputs(858);
    layer4_outputs(8340) <= not(layer3_outputs(2021));
    layer4_outputs(8341) <= not(layer3_outputs(3464)) or (layer3_outputs(4740));
    layer4_outputs(8342) <= layer3_outputs(7278);
    layer4_outputs(8343) <= (layer3_outputs(615)) and (layer3_outputs(1613));
    layer4_outputs(8344) <= not(layer3_outputs(9344));
    layer4_outputs(8345) <= not(layer3_outputs(9553));
    layer4_outputs(8346) <= not(layer3_outputs(4674));
    layer4_outputs(8347) <= (layer3_outputs(2067)) or (layer3_outputs(4675));
    layer4_outputs(8348) <= not(layer3_outputs(947));
    layer4_outputs(8349) <= layer3_outputs(4810);
    layer4_outputs(8350) <= '0';
    layer4_outputs(8351) <= not(layer3_outputs(988));
    layer4_outputs(8352) <= not(layer3_outputs(801));
    layer4_outputs(8353) <= not(layer3_outputs(7946));
    layer4_outputs(8354) <= not((layer3_outputs(7441)) or (layer3_outputs(2440)));
    layer4_outputs(8355) <= not((layer3_outputs(1018)) or (layer3_outputs(1031)));
    layer4_outputs(8356) <= not(layer3_outputs(576)) or (layer3_outputs(7967));
    layer4_outputs(8357) <= layer3_outputs(6210);
    layer4_outputs(8358) <= layer3_outputs(6591);
    layer4_outputs(8359) <= not(layer3_outputs(6093)) or (layer3_outputs(2082));
    layer4_outputs(8360) <= not(layer3_outputs(5166));
    layer4_outputs(8361) <= not(layer3_outputs(8499));
    layer4_outputs(8362) <= (layer3_outputs(3096)) xor (layer3_outputs(9679));
    layer4_outputs(8363) <= (layer3_outputs(6283)) or (layer3_outputs(6042));
    layer4_outputs(8364) <= not(layer3_outputs(5807));
    layer4_outputs(8365) <= layer3_outputs(7486);
    layer4_outputs(8366) <= layer3_outputs(9252);
    layer4_outputs(8367) <= not(layer3_outputs(7118));
    layer4_outputs(8368) <= (layer3_outputs(4898)) and not (layer3_outputs(9424));
    layer4_outputs(8369) <= layer3_outputs(6709);
    layer4_outputs(8370) <= layer3_outputs(2117);
    layer4_outputs(8371) <= (layer3_outputs(95)) xor (layer3_outputs(6603));
    layer4_outputs(8372) <= layer3_outputs(4630);
    layer4_outputs(8373) <= not(layer3_outputs(7158));
    layer4_outputs(8374) <= layer3_outputs(5976);
    layer4_outputs(8375) <= not(layer3_outputs(6805));
    layer4_outputs(8376) <= layer3_outputs(7458);
    layer4_outputs(8377) <= not(layer3_outputs(3958));
    layer4_outputs(8378) <= not(layer3_outputs(1626));
    layer4_outputs(8379) <= not(layer3_outputs(1098));
    layer4_outputs(8380) <= not((layer3_outputs(9714)) or (layer3_outputs(6338)));
    layer4_outputs(8381) <= not((layer3_outputs(8453)) xor (layer3_outputs(6427)));
    layer4_outputs(8382) <= layer3_outputs(5977);
    layer4_outputs(8383) <= layer3_outputs(8884);
    layer4_outputs(8384) <= not(layer3_outputs(9088));
    layer4_outputs(8385) <= (layer3_outputs(3860)) and not (layer3_outputs(6379));
    layer4_outputs(8386) <= not(layer3_outputs(7800));
    layer4_outputs(8387) <= layer3_outputs(8800);
    layer4_outputs(8388) <= layer3_outputs(4606);
    layer4_outputs(8389) <= layer3_outputs(335);
    layer4_outputs(8390) <= not(layer3_outputs(4969)) or (layer3_outputs(2656));
    layer4_outputs(8391) <= layer3_outputs(5945);
    layer4_outputs(8392) <= not(layer3_outputs(7327));
    layer4_outputs(8393) <= not(layer3_outputs(8106));
    layer4_outputs(8394) <= layer3_outputs(4110);
    layer4_outputs(8395) <= (layer3_outputs(10047)) and not (layer3_outputs(9341));
    layer4_outputs(8396) <= layer3_outputs(2783);
    layer4_outputs(8397) <= layer3_outputs(5333);
    layer4_outputs(8398) <= not(layer3_outputs(4032));
    layer4_outputs(8399) <= layer3_outputs(5449);
    layer4_outputs(8400) <= not(layer3_outputs(2650));
    layer4_outputs(8401) <= not((layer3_outputs(4627)) xor (layer3_outputs(3404)));
    layer4_outputs(8402) <= not((layer3_outputs(1526)) and (layer3_outputs(1996)));
    layer4_outputs(8403) <= not(layer3_outputs(3390));
    layer4_outputs(8404) <= (layer3_outputs(211)) and (layer3_outputs(1790));
    layer4_outputs(8405) <= not(layer3_outputs(7817));
    layer4_outputs(8406) <= not(layer3_outputs(758)) or (layer3_outputs(8063));
    layer4_outputs(8407) <= (layer3_outputs(7807)) and not (layer3_outputs(3420));
    layer4_outputs(8408) <= not(layer3_outputs(191));
    layer4_outputs(8409) <= not(layer3_outputs(5522));
    layer4_outputs(8410) <= not((layer3_outputs(2976)) and (layer3_outputs(792)));
    layer4_outputs(8411) <= not((layer3_outputs(3186)) or (layer3_outputs(5635)));
    layer4_outputs(8412) <= layer3_outputs(2021);
    layer4_outputs(8413) <= not(layer3_outputs(4379));
    layer4_outputs(8414) <= layer3_outputs(2698);
    layer4_outputs(8415) <= not(layer3_outputs(3303)) or (layer3_outputs(1808));
    layer4_outputs(8416) <= not((layer3_outputs(4783)) xor (layer3_outputs(7883)));
    layer4_outputs(8417) <= not((layer3_outputs(6765)) xor (layer3_outputs(9642)));
    layer4_outputs(8418) <= layer3_outputs(7783);
    layer4_outputs(8419) <= not(layer3_outputs(4398));
    layer4_outputs(8420) <= not(layer3_outputs(3715));
    layer4_outputs(8421) <= layer3_outputs(7501);
    layer4_outputs(8422) <= layer3_outputs(10088);
    layer4_outputs(8423) <= not(layer3_outputs(4176));
    layer4_outputs(8424) <= (layer3_outputs(8047)) or (layer3_outputs(1414));
    layer4_outputs(8425) <= layer3_outputs(5826);
    layer4_outputs(8426) <= not(layer3_outputs(1090));
    layer4_outputs(8427) <= not((layer3_outputs(7421)) and (layer3_outputs(4962)));
    layer4_outputs(8428) <= layer3_outputs(3185);
    layer4_outputs(8429) <= not(layer3_outputs(4134));
    layer4_outputs(8430) <= not(layer3_outputs(8177));
    layer4_outputs(8431) <= not((layer3_outputs(9135)) xor (layer3_outputs(9102)));
    layer4_outputs(8432) <= (layer3_outputs(4730)) and (layer3_outputs(8037));
    layer4_outputs(8433) <= (layer3_outputs(4697)) or (layer3_outputs(2076));
    layer4_outputs(8434) <= not((layer3_outputs(895)) xor (layer3_outputs(10211)));
    layer4_outputs(8435) <= layer3_outputs(5824);
    layer4_outputs(8436) <= not((layer3_outputs(633)) or (layer3_outputs(1763)));
    layer4_outputs(8437) <= (layer3_outputs(2953)) or (layer3_outputs(1469));
    layer4_outputs(8438) <= layer3_outputs(8898);
    layer4_outputs(8439) <= layer3_outputs(1294);
    layer4_outputs(8440) <= not(layer3_outputs(7918));
    layer4_outputs(8441) <= (layer3_outputs(3244)) xor (layer3_outputs(672));
    layer4_outputs(8442) <= (layer3_outputs(9451)) xor (layer3_outputs(57));
    layer4_outputs(8443) <= not((layer3_outputs(7621)) or (layer3_outputs(6863)));
    layer4_outputs(8444) <= not(layer3_outputs(3467));
    layer4_outputs(8445) <= (layer3_outputs(10139)) xor (layer3_outputs(9272));
    layer4_outputs(8446) <= not((layer3_outputs(9800)) xor (layer3_outputs(4436)));
    layer4_outputs(8447) <= not(layer3_outputs(4188));
    layer4_outputs(8448) <= (layer3_outputs(4546)) xor (layer3_outputs(944));
    layer4_outputs(8449) <= layer3_outputs(666);
    layer4_outputs(8450) <= not(layer3_outputs(6309));
    layer4_outputs(8451) <= not(layer3_outputs(9578));
    layer4_outputs(8452) <= layer3_outputs(6820);
    layer4_outputs(8453) <= (layer3_outputs(847)) xor (layer3_outputs(4966));
    layer4_outputs(8454) <= (layer3_outputs(2080)) and not (layer3_outputs(5249));
    layer4_outputs(8455) <= not(layer3_outputs(4440));
    layer4_outputs(8456) <= not(layer3_outputs(1406));
    layer4_outputs(8457) <= not(layer3_outputs(2808));
    layer4_outputs(8458) <= layer3_outputs(5248);
    layer4_outputs(8459) <= (layer3_outputs(3740)) and not (layer3_outputs(4662));
    layer4_outputs(8460) <= not(layer3_outputs(1215)) or (layer3_outputs(8456));
    layer4_outputs(8461) <= layer3_outputs(8498);
    layer4_outputs(8462) <= (layer3_outputs(1006)) xor (layer3_outputs(9640));
    layer4_outputs(8463) <= not(layer3_outputs(4917)) or (layer3_outputs(7080));
    layer4_outputs(8464) <= (layer3_outputs(9785)) and not (layer3_outputs(4215));
    layer4_outputs(8465) <= not((layer3_outputs(8257)) and (layer3_outputs(4229)));
    layer4_outputs(8466) <= (layer3_outputs(1930)) and not (layer3_outputs(5647));
    layer4_outputs(8467) <= layer3_outputs(4528);
    layer4_outputs(8468) <= not((layer3_outputs(2654)) xor (layer3_outputs(212)));
    layer4_outputs(8469) <= not(layer3_outputs(9144));
    layer4_outputs(8470) <= (layer3_outputs(10130)) and not (layer3_outputs(1810));
    layer4_outputs(8471) <= layer3_outputs(3267);
    layer4_outputs(8472) <= not(layer3_outputs(3318));
    layer4_outputs(8473) <= layer3_outputs(1816);
    layer4_outputs(8474) <= layer3_outputs(4704);
    layer4_outputs(8475) <= not(layer3_outputs(1719));
    layer4_outputs(8476) <= not((layer3_outputs(1341)) and (layer3_outputs(8573)));
    layer4_outputs(8477) <= not(layer3_outputs(6451));
    layer4_outputs(8478) <= not((layer3_outputs(6149)) and (layer3_outputs(5839)));
    layer4_outputs(8479) <= layer3_outputs(2106);
    layer4_outputs(8480) <= (layer3_outputs(8491)) xor (layer3_outputs(199));
    layer4_outputs(8481) <= layer3_outputs(2788);
    layer4_outputs(8482) <= layer3_outputs(1193);
    layer4_outputs(8483) <= not((layer3_outputs(4649)) xor (layer3_outputs(7756)));
    layer4_outputs(8484) <= (layer3_outputs(967)) or (layer3_outputs(6686));
    layer4_outputs(8485) <= layer3_outputs(6625);
    layer4_outputs(8486) <= not(layer3_outputs(7458));
    layer4_outputs(8487) <= (layer3_outputs(2595)) or (layer3_outputs(9295));
    layer4_outputs(8488) <= not((layer3_outputs(2186)) or (layer3_outputs(9475)));
    layer4_outputs(8489) <= (layer3_outputs(2416)) xor (layer3_outputs(4416));
    layer4_outputs(8490) <= layer3_outputs(4030);
    layer4_outputs(8491) <= (layer3_outputs(7273)) xor (layer3_outputs(636));
    layer4_outputs(8492) <= (layer3_outputs(9373)) or (layer3_outputs(5648));
    layer4_outputs(8493) <= not((layer3_outputs(5953)) xor (layer3_outputs(8763)));
    layer4_outputs(8494) <= not((layer3_outputs(4469)) xor (layer3_outputs(3697)));
    layer4_outputs(8495) <= '1';
    layer4_outputs(8496) <= not(layer3_outputs(411));
    layer4_outputs(8497) <= (layer3_outputs(7255)) and not (layer3_outputs(265));
    layer4_outputs(8498) <= layer3_outputs(5031);
    layer4_outputs(8499) <= (layer3_outputs(2)) and (layer3_outputs(7553));
    layer4_outputs(8500) <= not((layer3_outputs(5460)) and (layer3_outputs(1497)));
    layer4_outputs(8501) <= not((layer3_outputs(8780)) xor (layer3_outputs(3495)));
    layer4_outputs(8502) <= '1';
    layer4_outputs(8503) <= (layer3_outputs(6070)) and not (layer3_outputs(6873));
    layer4_outputs(8504) <= not((layer3_outputs(3696)) and (layer3_outputs(5052)));
    layer4_outputs(8505) <= not(layer3_outputs(5685));
    layer4_outputs(8506) <= not(layer3_outputs(422));
    layer4_outputs(8507) <= not(layer3_outputs(1322));
    layer4_outputs(8508) <= not(layer3_outputs(8401)) or (layer3_outputs(5406));
    layer4_outputs(8509) <= (layer3_outputs(7014)) or (layer3_outputs(875));
    layer4_outputs(8510) <= (layer3_outputs(7598)) or (layer3_outputs(5208));
    layer4_outputs(8511) <= not((layer3_outputs(8553)) and (layer3_outputs(9302)));
    layer4_outputs(8512) <= not((layer3_outputs(7807)) or (layer3_outputs(2428)));
    layer4_outputs(8513) <= layer3_outputs(7811);
    layer4_outputs(8514) <= not(layer3_outputs(2605));
    layer4_outputs(8515) <= layer3_outputs(3376);
    layer4_outputs(8516) <= not(layer3_outputs(370)) or (layer3_outputs(7643));
    layer4_outputs(8517) <= layer3_outputs(633);
    layer4_outputs(8518) <= not(layer3_outputs(6884)) or (layer3_outputs(2995));
    layer4_outputs(8519) <= (layer3_outputs(8699)) and not (layer3_outputs(8319));
    layer4_outputs(8520) <= (layer3_outputs(4117)) xor (layer3_outputs(9485));
    layer4_outputs(8521) <= not(layer3_outputs(9073));
    layer4_outputs(8522) <= not(layer3_outputs(3795));
    layer4_outputs(8523) <= not((layer3_outputs(1939)) xor (layer3_outputs(5635)));
    layer4_outputs(8524) <= not(layer3_outputs(7262));
    layer4_outputs(8525) <= layer3_outputs(8381);
    layer4_outputs(8526) <= layer3_outputs(4011);
    layer4_outputs(8527) <= layer3_outputs(8070);
    layer4_outputs(8528) <= not(layer3_outputs(7939));
    layer4_outputs(8529) <= not((layer3_outputs(2111)) and (layer3_outputs(3940)));
    layer4_outputs(8530) <= (layer3_outputs(9224)) and not (layer3_outputs(3203));
    layer4_outputs(8531) <= not((layer3_outputs(1326)) xor (layer3_outputs(3534)));
    layer4_outputs(8532) <= layer3_outputs(6561);
    layer4_outputs(8533) <= not(layer3_outputs(1066)) or (layer3_outputs(1500));
    layer4_outputs(8534) <= '0';
    layer4_outputs(8535) <= not(layer3_outputs(8063));
    layer4_outputs(8536) <= layer3_outputs(9800);
    layer4_outputs(8537) <= not(layer3_outputs(5693));
    layer4_outputs(8538) <= not(layer3_outputs(497));
    layer4_outputs(8539) <= not(layer3_outputs(4226));
    layer4_outputs(8540) <= (layer3_outputs(3826)) xor (layer3_outputs(4025));
    layer4_outputs(8541) <= layer3_outputs(5622);
    layer4_outputs(8542) <= layer3_outputs(5285);
    layer4_outputs(8543) <= not(layer3_outputs(9115));
    layer4_outputs(8544) <= not(layer3_outputs(9578));
    layer4_outputs(8545) <= not(layer3_outputs(7711));
    layer4_outputs(8546) <= not(layer3_outputs(5393)) or (layer3_outputs(1793));
    layer4_outputs(8547) <= not((layer3_outputs(5593)) and (layer3_outputs(2081)));
    layer4_outputs(8548) <= (layer3_outputs(8769)) and not (layer3_outputs(9031));
    layer4_outputs(8549) <= not(layer3_outputs(8485)) or (layer3_outputs(7847));
    layer4_outputs(8550) <= layer3_outputs(1956);
    layer4_outputs(8551) <= not(layer3_outputs(7433));
    layer4_outputs(8552) <= (layer3_outputs(1037)) or (layer3_outputs(4565));
    layer4_outputs(8553) <= not(layer3_outputs(2477));
    layer4_outputs(8554) <= (layer3_outputs(1835)) xor (layer3_outputs(1596));
    layer4_outputs(8555) <= not((layer3_outputs(3573)) xor (layer3_outputs(9506)));
    layer4_outputs(8556) <= not((layer3_outputs(8086)) xor (layer3_outputs(8439)));
    layer4_outputs(8557) <= not(layer3_outputs(4752)) or (layer3_outputs(6102));
    layer4_outputs(8558) <= '0';
    layer4_outputs(8559) <= not((layer3_outputs(10072)) or (layer3_outputs(539)));
    layer4_outputs(8560) <= not(layer3_outputs(7625));
    layer4_outputs(8561) <= (layer3_outputs(9850)) xor (layer3_outputs(7542));
    layer4_outputs(8562) <= layer3_outputs(7007);
    layer4_outputs(8563) <= not((layer3_outputs(8082)) and (layer3_outputs(7434)));
    layer4_outputs(8564) <= not((layer3_outputs(4074)) or (layer3_outputs(6757)));
    layer4_outputs(8565) <= not(layer3_outputs(5746));
    layer4_outputs(8566) <= layer3_outputs(7419);
    layer4_outputs(8567) <= '0';
    layer4_outputs(8568) <= not(layer3_outputs(2435));
    layer4_outputs(8569) <= layer3_outputs(3010);
    layer4_outputs(8570) <= not((layer3_outputs(4928)) xor (layer3_outputs(3192)));
    layer4_outputs(8571) <= not((layer3_outputs(1950)) and (layer3_outputs(1393)));
    layer4_outputs(8572) <= layer3_outputs(75);
    layer4_outputs(8573) <= not((layer3_outputs(10201)) xor (layer3_outputs(9017)));
    layer4_outputs(8574) <= not(layer3_outputs(4668)) or (layer3_outputs(2288));
    layer4_outputs(8575) <= not(layer3_outputs(7831));
    layer4_outputs(8576) <= not(layer3_outputs(2929));
    layer4_outputs(8577) <= layer3_outputs(8026);
    layer4_outputs(8578) <= not(layer3_outputs(8218)) or (layer3_outputs(7699));
    layer4_outputs(8579) <= not(layer3_outputs(6994));
    layer4_outputs(8580) <= not((layer3_outputs(9928)) or (layer3_outputs(585)));
    layer4_outputs(8581) <= layer3_outputs(8770);
    layer4_outputs(8582) <= (layer3_outputs(172)) and not (layer3_outputs(2352));
    layer4_outputs(8583) <= not(layer3_outputs(5616));
    layer4_outputs(8584) <= (layer3_outputs(6226)) xor (layer3_outputs(9709));
    layer4_outputs(8585) <= not(layer3_outputs(4672));
    layer4_outputs(8586) <= layer3_outputs(2054);
    layer4_outputs(8587) <= layer3_outputs(9240);
    layer4_outputs(8588) <= not((layer3_outputs(6385)) xor (layer3_outputs(2099)));
    layer4_outputs(8589) <= not(layer3_outputs(7322));
    layer4_outputs(8590) <= not(layer3_outputs(7919));
    layer4_outputs(8591) <= (layer3_outputs(4637)) and not (layer3_outputs(5716));
    layer4_outputs(8592) <= (layer3_outputs(9449)) or (layer3_outputs(9343));
    layer4_outputs(8593) <= not((layer3_outputs(9412)) xor (layer3_outputs(8899)));
    layer4_outputs(8594) <= (layer3_outputs(7846)) xor (layer3_outputs(3366));
    layer4_outputs(8595) <= layer3_outputs(7213);
    layer4_outputs(8596) <= layer3_outputs(10224);
    layer4_outputs(8597) <= (layer3_outputs(8635)) xor (layer3_outputs(5957));
    layer4_outputs(8598) <= '0';
    layer4_outputs(8599) <= (layer3_outputs(6998)) xor (layer3_outputs(1768));
    layer4_outputs(8600) <= not(layer3_outputs(4586)) or (layer3_outputs(4214));
    layer4_outputs(8601) <= not(layer3_outputs(1569));
    layer4_outputs(8602) <= not(layer3_outputs(3593));
    layer4_outputs(8603) <= not(layer3_outputs(9225));
    layer4_outputs(8604) <= layer3_outputs(357);
    layer4_outputs(8605) <= layer3_outputs(4947);
    layer4_outputs(8606) <= layer3_outputs(7517);
    layer4_outputs(8607) <= (layer3_outputs(6428)) xor (layer3_outputs(7591));
    layer4_outputs(8608) <= not(layer3_outputs(5612));
    layer4_outputs(8609) <= layer3_outputs(392);
    layer4_outputs(8610) <= (layer3_outputs(7341)) xor (layer3_outputs(9856));
    layer4_outputs(8611) <= not(layer3_outputs(1066));
    layer4_outputs(8612) <= not(layer3_outputs(4346));
    layer4_outputs(8613) <= '0';
    layer4_outputs(8614) <= layer3_outputs(9298);
    layer4_outputs(8615) <= layer3_outputs(9498);
    layer4_outputs(8616) <= not(layer3_outputs(1685));
    layer4_outputs(8617) <= (layer3_outputs(9602)) and (layer3_outputs(6556));
    layer4_outputs(8618) <= layer3_outputs(387);
    layer4_outputs(8619) <= not(layer3_outputs(7812)) or (layer3_outputs(2113));
    layer4_outputs(8620) <= layer3_outputs(6551);
    layer4_outputs(8621) <= layer3_outputs(8176);
    layer4_outputs(8622) <= not(layer3_outputs(177));
    layer4_outputs(8623) <= '0';
    layer4_outputs(8624) <= not(layer3_outputs(544));
    layer4_outputs(8625) <= not(layer3_outputs(2959)) or (layer3_outputs(9892));
    layer4_outputs(8626) <= not(layer3_outputs(9681));
    layer4_outputs(8627) <= layer3_outputs(248);
    layer4_outputs(8628) <= not(layer3_outputs(5305)) or (layer3_outputs(1783));
    layer4_outputs(8629) <= (layer3_outputs(7268)) and (layer3_outputs(7775));
    layer4_outputs(8630) <= (layer3_outputs(840)) xor (layer3_outputs(8452));
    layer4_outputs(8631) <= not(layer3_outputs(6901));
    layer4_outputs(8632) <= layer3_outputs(5141);
    layer4_outputs(8633) <= (layer3_outputs(7402)) and not (layer3_outputs(5331));
    layer4_outputs(8634) <= not(layer3_outputs(6625));
    layer4_outputs(8635) <= not(layer3_outputs(7943)) or (layer3_outputs(2510));
    layer4_outputs(8636) <= layer3_outputs(8289);
    layer4_outputs(8637) <= layer3_outputs(5557);
    layer4_outputs(8638) <= not(layer3_outputs(5990));
    layer4_outputs(8639) <= (layer3_outputs(6789)) and (layer3_outputs(4880));
    layer4_outputs(8640) <= not(layer3_outputs(5368));
    layer4_outputs(8641) <= not(layer3_outputs(3835));
    layer4_outputs(8642) <= not(layer3_outputs(9660));
    layer4_outputs(8643) <= not(layer3_outputs(981));
    layer4_outputs(8644) <= not(layer3_outputs(3366));
    layer4_outputs(8645) <= layer3_outputs(2231);
    layer4_outputs(8646) <= not(layer3_outputs(1158));
    layer4_outputs(8647) <= not(layer3_outputs(4237));
    layer4_outputs(8648) <= not(layer3_outputs(4682));
    layer4_outputs(8649) <= not(layer3_outputs(6242));
    layer4_outputs(8650) <= layer3_outputs(7284);
    layer4_outputs(8651) <= not(layer3_outputs(2575));
    layer4_outputs(8652) <= not(layer3_outputs(1717));
    layer4_outputs(8653) <= not(layer3_outputs(7702)) or (layer3_outputs(5740));
    layer4_outputs(8654) <= layer3_outputs(3708);
    layer4_outputs(8655) <= not(layer3_outputs(2922));
    layer4_outputs(8656) <= not(layer3_outputs(377));
    layer4_outputs(8657) <= layer3_outputs(10174);
    layer4_outputs(8658) <= (layer3_outputs(9107)) or (layer3_outputs(8369));
    layer4_outputs(8659) <= not((layer3_outputs(3776)) and (layer3_outputs(7155)));
    layer4_outputs(8660) <= layer3_outputs(9749);
    layer4_outputs(8661) <= not(layer3_outputs(4444)) or (layer3_outputs(7981));
    layer4_outputs(8662) <= layer3_outputs(188);
    layer4_outputs(8663) <= not((layer3_outputs(8692)) xor (layer3_outputs(4809)));
    layer4_outputs(8664) <= not(layer3_outputs(4359));
    layer4_outputs(8665) <= not((layer3_outputs(8276)) xor (layer3_outputs(5237)));
    layer4_outputs(8666) <= not(layer3_outputs(4643)) or (layer3_outputs(495));
    layer4_outputs(8667) <= not(layer3_outputs(8356)) or (layer3_outputs(6850));
    layer4_outputs(8668) <= not(layer3_outputs(10163));
    layer4_outputs(8669) <= not((layer3_outputs(5104)) xor (layer3_outputs(2264)));
    layer4_outputs(8670) <= not((layer3_outputs(4169)) and (layer3_outputs(4770)));
    layer4_outputs(8671) <= not(layer3_outputs(4711));
    layer4_outputs(8672) <= not(layer3_outputs(5236));
    layer4_outputs(8673) <= layer3_outputs(949);
    layer4_outputs(8674) <= layer3_outputs(8571);
    layer4_outputs(8675) <= not(layer3_outputs(2819)) or (layer3_outputs(7626));
    layer4_outputs(8676) <= not(layer3_outputs(7270));
    layer4_outputs(8677) <= not(layer3_outputs(1182));
    layer4_outputs(8678) <= (layer3_outputs(7295)) or (layer3_outputs(1177));
    layer4_outputs(8679) <= layer3_outputs(7905);
    layer4_outputs(8680) <= not(layer3_outputs(5246));
    layer4_outputs(8681) <= (layer3_outputs(489)) and (layer3_outputs(9665));
    layer4_outputs(8682) <= not(layer3_outputs(1661));
    layer4_outputs(8683) <= (layer3_outputs(7884)) xor (layer3_outputs(5491));
    layer4_outputs(8684) <= layer3_outputs(511);
    layer4_outputs(8685) <= layer3_outputs(7266);
    layer4_outputs(8686) <= not(layer3_outputs(6146));
    layer4_outputs(8687) <= (layer3_outputs(5669)) and (layer3_outputs(4167));
    layer4_outputs(8688) <= (layer3_outputs(6770)) and not (layer3_outputs(5783));
    layer4_outputs(8689) <= (layer3_outputs(9075)) and not (layer3_outputs(6368));
    layer4_outputs(8690) <= not((layer3_outputs(314)) and (layer3_outputs(4053)));
    layer4_outputs(8691) <= layer3_outputs(8996);
    layer4_outputs(8692) <= not((layer3_outputs(8137)) and (layer3_outputs(5991)));
    layer4_outputs(8693) <= layer3_outputs(7403);
    layer4_outputs(8694) <= (layer3_outputs(7647)) and (layer3_outputs(9488));
    layer4_outputs(8695) <= (layer3_outputs(8123)) and not (layer3_outputs(8921));
    layer4_outputs(8696) <= not(layer3_outputs(7813));
    layer4_outputs(8697) <= layer3_outputs(9111);
    layer4_outputs(8698) <= not((layer3_outputs(3435)) or (layer3_outputs(6897)));
    layer4_outputs(8699) <= layer3_outputs(6104);
    layer4_outputs(8700) <= not(layer3_outputs(9738)) or (layer3_outputs(9080));
    layer4_outputs(8701) <= not(layer3_outputs(2620)) or (layer3_outputs(8805));
    layer4_outputs(8702) <= not(layer3_outputs(7180));
    layer4_outputs(8703) <= not(layer3_outputs(9395));
    layer4_outputs(8704) <= not(layer3_outputs(141));
    layer4_outputs(8705) <= (layer3_outputs(7663)) xor (layer3_outputs(6448));
    layer4_outputs(8706) <= not(layer3_outputs(4228));
    layer4_outputs(8707) <= layer3_outputs(5150);
    layer4_outputs(8708) <= not((layer3_outputs(1872)) xor (layer3_outputs(7555)));
    layer4_outputs(8709) <= not(layer3_outputs(3200));
    layer4_outputs(8710) <= not(layer3_outputs(3999));
    layer4_outputs(8711) <= layer3_outputs(3977);
    layer4_outputs(8712) <= not(layer3_outputs(1844));
    layer4_outputs(8713) <= not((layer3_outputs(7572)) or (layer3_outputs(1187)));
    layer4_outputs(8714) <= layer3_outputs(7075);
    layer4_outputs(8715) <= layer3_outputs(961);
    layer4_outputs(8716) <= (layer3_outputs(8492)) xor (layer3_outputs(4839));
    layer4_outputs(8717) <= layer3_outputs(3266);
    layer4_outputs(8718) <= not(layer3_outputs(8440));
    layer4_outputs(8719) <= not(layer3_outputs(7031));
    layer4_outputs(8720) <= layer3_outputs(9735);
    layer4_outputs(8721) <= layer3_outputs(4858);
    layer4_outputs(8722) <= (layer3_outputs(1140)) and (layer3_outputs(3301));
    layer4_outputs(8723) <= (layer3_outputs(4306)) and not (layer3_outputs(7781));
    layer4_outputs(8724) <= not((layer3_outputs(1599)) xor (layer3_outputs(4402)));
    layer4_outputs(8725) <= not(layer3_outputs(7190));
    layer4_outputs(8726) <= not(layer3_outputs(3497));
    layer4_outputs(8727) <= not(layer3_outputs(1610));
    layer4_outputs(8728) <= layer3_outputs(7079);
    layer4_outputs(8729) <= (layer3_outputs(8167)) and (layer3_outputs(539));
    layer4_outputs(8730) <= layer3_outputs(2513);
    layer4_outputs(8731) <= not(layer3_outputs(5871));
    layer4_outputs(8732) <= (layer3_outputs(2408)) xor (layer3_outputs(5705));
    layer4_outputs(8733) <= layer3_outputs(5379);
    layer4_outputs(8734) <= not((layer3_outputs(9375)) xor (layer3_outputs(4414)));
    layer4_outputs(8735) <= not(layer3_outputs(2233));
    layer4_outputs(8736) <= (layer3_outputs(7431)) xor (layer3_outputs(2403));
    layer4_outputs(8737) <= not((layer3_outputs(9383)) xor (layer3_outputs(9156)));
    layer4_outputs(8738) <= (layer3_outputs(933)) and not (layer3_outputs(1002));
    layer4_outputs(8739) <= not(layer3_outputs(1826)) or (layer3_outputs(8406));
    layer4_outputs(8740) <= (layer3_outputs(4420)) xor (layer3_outputs(4122));
    layer4_outputs(8741) <= not(layer3_outputs(1130));
    layer4_outputs(8742) <= not(layer3_outputs(675));
    layer4_outputs(8743) <= not(layer3_outputs(7749));
    layer4_outputs(8744) <= (layer3_outputs(8039)) xor (layer3_outputs(4707));
    layer4_outputs(8745) <= not(layer3_outputs(6026)) or (layer3_outputs(5348));
    layer4_outputs(8746) <= (layer3_outputs(9081)) and not (layer3_outputs(7391));
    layer4_outputs(8747) <= not(layer3_outputs(2990));
    layer4_outputs(8748) <= not(layer3_outputs(9303));
    layer4_outputs(8749) <= not(layer3_outputs(1766)) or (layer3_outputs(5853));
    layer4_outputs(8750) <= not(layer3_outputs(600)) or (layer3_outputs(5185));
    layer4_outputs(8751) <= layer3_outputs(3286);
    layer4_outputs(8752) <= (layer3_outputs(4086)) and (layer3_outputs(292));
    layer4_outputs(8753) <= layer3_outputs(2561);
    layer4_outputs(8754) <= not(layer3_outputs(5550));
    layer4_outputs(8755) <= layer3_outputs(1457);
    layer4_outputs(8756) <= (layer3_outputs(9875)) or (layer3_outputs(2952));
    layer4_outputs(8757) <= not((layer3_outputs(4206)) xor (layer3_outputs(8833)));
    layer4_outputs(8758) <= layer3_outputs(9369);
    layer4_outputs(8759) <= not(layer3_outputs(3842));
    layer4_outputs(8760) <= layer3_outputs(5753);
    layer4_outputs(8761) <= layer3_outputs(9500);
    layer4_outputs(8762) <= layer3_outputs(2867);
    layer4_outputs(8763) <= (layer3_outputs(548)) and not (layer3_outputs(655));
    layer4_outputs(8764) <= not(layer3_outputs(869)) or (layer3_outputs(30));
    layer4_outputs(8765) <= not(layer3_outputs(8720)) or (layer3_outputs(6335));
    layer4_outputs(8766) <= (layer3_outputs(760)) and not (layer3_outputs(7371));
    layer4_outputs(8767) <= not(layer3_outputs(9457));
    layer4_outputs(8768) <= layer3_outputs(4979);
    layer4_outputs(8769) <= not(layer3_outputs(1911));
    layer4_outputs(8770) <= not(layer3_outputs(3347));
    layer4_outputs(8771) <= not(layer3_outputs(10029));
    layer4_outputs(8772) <= layer3_outputs(2901);
    layer4_outputs(8773) <= (layer3_outputs(410)) and not (layer3_outputs(4573));
    layer4_outputs(8774) <= not(layer3_outputs(5386));
    layer4_outputs(8775) <= layer3_outputs(5705);
    layer4_outputs(8776) <= layer3_outputs(6341);
    layer4_outputs(8777) <= not(layer3_outputs(3956));
    layer4_outputs(8778) <= layer3_outputs(6193);
    layer4_outputs(8779) <= layer3_outputs(6360);
    layer4_outputs(8780) <= layer3_outputs(9932);
    layer4_outputs(8781) <= layer3_outputs(7365);
    layer4_outputs(8782) <= not(layer3_outputs(485));
    layer4_outputs(8783) <= not(layer3_outputs(4490));
    layer4_outputs(8784) <= not(layer3_outputs(960));
    layer4_outputs(8785) <= (layer3_outputs(6381)) and (layer3_outputs(3132));
    layer4_outputs(8786) <= layer3_outputs(1810);
    layer4_outputs(8787) <= layer3_outputs(5764);
    layer4_outputs(8788) <= layer3_outputs(2046);
    layer4_outputs(8789) <= not(layer3_outputs(246));
    layer4_outputs(8790) <= not((layer3_outputs(8725)) or (layer3_outputs(1325)));
    layer4_outputs(8791) <= layer3_outputs(8100);
    layer4_outputs(8792) <= layer3_outputs(8339);
    layer4_outputs(8793) <= (layer3_outputs(5650)) and not (layer3_outputs(3872));
    layer4_outputs(8794) <= not((layer3_outputs(8493)) or (layer3_outputs(8864)));
    layer4_outputs(8795) <= (layer3_outputs(5349)) xor (layer3_outputs(5829));
    layer4_outputs(8796) <= not((layer3_outputs(4386)) xor (layer3_outputs(5239)));
    layer4_outputs(8797) <= (layer3_outputs(2212)) and (layer3_outputs(8667));
    layer4_outputs(8798) <= not(layer3_outputs(5988)) or (layer3_outputs(4523));
    layer4_outputs(8799) <= (layer3_outputs(4046)) xor (layer3_outputs(5356));
    layer4_outputs(8800) <= layer3_outputs(5634);
    layer4_outputs(8801) <= layer3_outputs(5335);
    layer4_outputs(8802) <= not(layer3_outputs(3012));
    layer4_outputs(8803) <= (layer3_outputs(9372)) xor (layer3_outputs(7006));
    layer4_outputs(8804) <= not(layer3_outputs(9205));
    layer4_outputs(8805) <= not((layer3_outputs(6563)) and (layer3_outputs(6272)));
    layer4_outputs(8806) <= not((layer3_outputs(2768)) and (layer3_outputs(4425)));
    layer4_outputs(8807) <= layer3_outputs(6271);
    layer4_outputs(8808) <= layer3_outputs(9134);
    layer4_outputs(8809) <= not(layer3_outputs(8995));
    layer4_outputs(8810) <= (layer3_outputs(1120)) xor (layer3_outputs(7179));
    layer4_outputs(8811) <= (layer3_outputs(7828)) and (layer3_outputs(9724));
    layer4_outputs(8812) <= not((layer3_outputs(4682)) and (layer3_outputs(6310)));
    layer4_outputs(8813) <= not((layer3_outputs(2749)) and (layer3_outputs(8684)));
    layer4_outputs(8814) <= layer3_outputs(1172);
    layer4_outputs(8815) <= not(layer3_outputs(3567));
    layer4_outputs(8816) <= (layer3_outputs(7083)) and not (layer3_outputs(836));
    layer4_outputs(8817) <= not(layer3_outputs(8396));
    layer4_outputs(8818) <= (layer3_outputs(4874)) and (layer3_outputs(5549));
    layer4_outputs(8819) <= layer3_outputs(806);
    layer4_outputs(8820) <= (layer3_outputs(8461)) and not (layer3_outputs(342));
    layer4_outputs(8821) <= layer3_outputs(2186);
    layer4_outputs(8822) <= layer3_outputs(5742);
    layer4_outputs(8823) <= not(layer3_outputs(7916));
    layer4_outputs(8824) <= not(layer3_outputs(9874));
    layer4_outputs(8825) <= not((layer3_outputs(84)) or (layer3_outputs(4689)));
    layer4_outputs(8826) <= layer3_outputs(2426);
    layer4_outputs(8827) <= not(layer3_outputs(1170)) or (layer3_outputs(1894));
    layer4_outputs(8828) <= layer3_outputs(6235);
    layer4_outputs(8829) <= (layer3_outputs(3036)) xor (layer3_outputs(10110));
    layer4_outputs(8830) <= not(layer3_outputs(5348));
    layer4_outputs(8831) <= not(layer3_outputs(8267));
    layer4_outputs(8832) <= (layer3_outputs(765)) and not (layer3_outputs(7445));
    layer4_outputs(8833) <= not((layer3_outputs(7361)) xor (layer3_outputs(387)));
    layer4_outputs(8834) <= (layer3_outputs(409)) and not (layer3_outputs(7721));
    layer4_outputs(8835) <= not(layer3_outputs(2143));
    layer4_outputs(8836) <= not((layer3_outputs(6280)) or (layer3_outputs(3907)));
    layer4_outputs(8837) <= not(layer3_outputs(5474)) or (layer3_outputs(9762));
    layer4_outputs(8838) <= not(layer3_outputs(2665)) or (layer3_outputs(618));
    layer4_outputs(8839) <= not(layer3_outputs(397));
    layer4_outputs(8840) <= (layer3_outputs(9496)) and not (layer3_outputs(5649));
    layer4_outputs(8841) <= not(layer3_outputs(6376));
    layer4_outputs(8842) <= layer3_outputs(5048);
    layer4_outputs(8843) <= layer3_outputs(1528);
    layer4_outputs(8844) <= (layer3_outputs(6293)) xor (layer3_outputs(7285));
    layer4_outputs(8845) <= layer3_outputs(1468);
    layer4_outputs(8846) <= not(layer3_outputs(5983)) or (layer3_outputs(1401));
    layer4_outputs(8847) <= (layer3_outputs(317)) xor (layer3_outputs(2423));
    layer4_outputs(8848) <= not((layer3_outputs(999)) xor (layer3_outputs(4748)));
    layer4_outputs(8849) <= not(layer3_outputs(1578));
    layer4_outputs(8850) <= layer3_outputs(6218);
    layer4_outputs(8851) <= not(layer3_outputs(2089));
    layer4_outputs(8852) <= layer3_outputs(9233);
    layer4_outputs(8853) <= (layer3_outputs(4316)) and not (layer3_outputs(6065));
    layer4_outputs(8854) <= layer3_outputs(9934);
    layer4_outputs(8855) <= not(layer3_outputs(4380));
    layer4_outputs(8856) <= (layer3_outputs(3665)) xor (layer3_outputs(6414));
    layer4_outputs(8857) <= (layer3_outputs(3562)) or (layer3_outputs(8443));
    layer4_outputs(8858) <= not((layer3_outputs(5935)) or (layer3_outputs(8368)));
    layer4_outputs(8859) <= (layer3_outputs(5212)) and not (layer3_outputs(2048));
    layer4_outputs(8860) <= not(layer3_outputs(6123));
    layer4_outputs(8861) <= not((layer3_outputs(5553)) xor (layer3_outputs(4339)));
    layer4_outputs(8862) <= layer3_outputs(1203);
    layer4_outputs(8863) <= not(layer3_outputs(8065));
    layer4_outputs(8864) <= not(layer3_outputs(214));
    layer4_outputs(8865) <= layer3_outputs(4554);
    layer4_outputs(8866) <= not((layer3_outputs(1305)) and (layer3_outputs(6036)));
    layer4_outputs(8867) <= (layer3_outputs(2579)) and not (layer3_outputs(9871));
    layer4_outputs(8868) <= not((layer3_outputs(8792)) xor (layer3_outputs(3010)));
    layer4_outputs(8869) <= not(layer3_outputs(7144));
    layer4_outputs(8870) <= not(layer3_outputs(1277));
    layer4_outputs(8871) <= layer3_outputs(4421);
    layer4_outputs(8872) <= (layer3_outputs(9872)) xor (layer3_outputs(3330));
    layer4_outputs(8873) <= '0';
    layer4_outputs(8874) <= not((layer3_outputs(6136)) or (layer3_outputs(9378)));
    layer4_outputs(8875) <= layer3_outputs(5395);
    layer4_outputs(8876) <= layer3_outputs(3936);
    layer4_outputs(8877) <= (layer3_outputs(4886)) and not (layer3_outputs(3552));
    layer4_outputs(8878) <= (layer3_outputs(7028)) and not (layer3_outputs(2220));
    layer4_outputs(8879) <= not((layer3_outputs(1396)) and (layer3_outputs(1061)));
    layer4_outputs(8880) <= layer3_outputs(2341);
    layer4_outputs(8881) <= layer3_outputs(3389);
    layer4_outputs(8882) <= not(layer3_outputs(9465));
    layer4_outputs(8883) <= not(layer3_outputs(832));
    layer4_outputs(8884) <= not((layer3_outputs(5054)) xor (layer3_outputs(8371)));
    layer4_outputs(8885) <= (layer3_outputs(8351)) and not (layer3_outputs(3984));
    layer4_outputs(8886) <= (layer3_outputs(7733)) xor (layer3_outputs(1275));
    layer4_outputs(8887) <= (layer3_outputs(7835)) xor (layer3_outputs(5010));
    layer4_outputs(8888) <= (layer3_outputs(7030)) or (layer3_outputs(884));
    layer4_outputs(8889) <= (layer3_outputs(8576)) and (layer3_outputs(2430));
    layer4_outputs(8890) <= layer3_outputs(1975);
    layer4_outputs(8891) <= not(layer3_outputs(9168));
    layer4_outputs(8892) <= not(layer3_outputs(1543));
    layer4_outputs(8893) <= '1';
    layer4_outputs(8894) <= (layer3_outputs(2055)) and (layer3_outputs(6585));
    layer4_outputs(8895) <= not(layer3_outputs(7224));
    layer4_outputs(8896) <= not(layer3_outputs(3218)) or (layer3_outputs(9385));
    layer4_outputs(8897) <= (layer3_outputs(4578)) and not (layer3_outputs(5030));
    layer4_outputs(8898) <= (layer3_outputs(8016)) and (layer3_outputs(6352));
    layer4_outputs(8899) <= layer3_outputs(6319);
    layer4_outputs(8900) <= not(layer3_outputs(7546));
    layer4_outputs(8901) <= not(layer3_outputs(2321)) or (layer3_outputs(1333));
    layer4_outputs(8902) <= '0';
    layer4_outputs(8903) <= not(layer3_outputs(920));
    layer4_outputs(8904) <= not(layer3_outputs(4203));
    layer4_outputs(8905) <= not(layer3_outputs(9839));
    layer4_outputs(8906) <= layer3_outputs(6495);
    layer4_outputs(8907) <= layer3_outputs(1229);
    layer4_outputs(8908) <= not(layer3_outputs(2027)) or (layer3_outputs(9984));
    layer4_outputs(8909) <= (layer3_outputs(1792)) or (layer3_outputs(5354));
    layer4_outputs(8910) <= layer3_outputs(2732);
    layer4_outputs(8911) <= not(layer3_outputs(1973));
    layer4_outputs(8912) <= not(layer3_outputs(3160));
    layer4_outputs(8913) <= layer3_outputs(5500);
    layer4_outputs(8914) <= not(layer3_outputs(9276)) or (layer3_outputs(886));
    layer4_outputs(8915) <= (layer3_outputs(4564)) xor (layer3_outputs(9755));
    layer4_outputs(8916) <= layer3_outputs(6329);
    layer4_outputs(8917) <= layer3_outputs(6848);
    layer4_outputs(8918) <= (layer3_outputs(7144)) or (layer3_outputs(149));
    layer4_outputs(8919) <= (layer3_outputs(9103)) xor (layer3_outputs(57));
    layer4_outputs(8920) <= layer3_outputs(4540);
    layer4_outputs(8921) <= (layer3_outputs(4173)) or (layer3_outputs(4771));
    layer4_outputs(8922) <= layer3_outputs(2286);
    layer4_outputs(8923) <= not(layer3_outputs(1788));
    layer4_outputs(8924) <= not(layer3_outputs(4663));
    layer4_outputs(8925) <= (layer3_outputs(2981)) or (layer3_outputs(8964));
    layer4_outputs(8926) <= layer3_outputs(6305);
    layer4_outputs(8927) <= not(layer3_outputs(429));
    layer4_outputs(8928) <= (layer3_outputs(2790)) and not (layer3_outputs(347));
    layer4_outputs(8929) <= not(layer3_outputs(7943)) or (layer3_outputs(9060));
    layer4_outputs(8930) <= layer3_outputs(9348);
    layer4_outputs(8931) <= not(layer3_outputs(7109));
    layer4_outputs(8932) <= layer3_outputs(6957);
    layer4_outputs(8933) <= (layer3_outputs(8111)) and not (layer3_outputs(4807));
    layer4_outputs(8934) <= layer3_outputs(8856);
    layer4_outputs(8935) <= not(layer3_outputs(2141));
    layer4_outputs(8936) <= (layer3_outputs(6359)) xor (layer3_outputs(5845));
    layer4_outputs(8937) <= not(layer3_outputs(5481)) or (layer3_outputs(5598));
    layer4_outputs(8938) <= not(layer3_outputs(1098));
    layer4_outputs(8939) <= not(layer3_outputs(6333));
    layer4_outputs(8940) <= layer3_outputs(9301);
    layer4_outputs(8941) <= not((layer3_outputs(1715)) xor (layer3_outputs(767)));
    layer4_outputs(8942) <= (layer3_outputs(7308)) and not (layer3_outputs(7115));
    layer4_outputs(8943) <= not((layer3_outputs(7214)) xor (layer3_outputs(9325)));
    layer4_outputs(8944) <= (layer3_outputs(8089)) or (layer3_outputs(2304));
    layer4_outputs(8945) <= not(layer3_outputs(7113)) or (layer3_outputs(341));
    layer4_outputs(8946) <= (layer3_outputs(6632)) xor (layer3_outputs(7539));
    layer4_outputs(8947) <= not(layer3_outputs(4837));
    layer4_outputs(8948) <= not(layer3_outputs(2073));
    layer4_outputs(8949) <= (layer3_outputs(639)) and not (layer3_outputs(508));
    layer4_outputs(8950) <= not(layer3_outputs(3848));
    layer4_outputs(8951) <= not(layer3_outputs(4102));
    layer4_outputs(8952) <= '1';
    layer4_outputs(8953) <= not(layer3_outputs(10117));
    layer4_outputs(8954) <= (layer3_outputs(441)) and not (layer3_outputs(9482));
    layer4_outputs(8955) <= not(layer3_outputs(4936));
    layer4_outputs(8956) <= layer3_outputs(9774);
    layer4_outputs(8957) <= not(layer3_outputs(6222)) or (layer3_outputs(6115));
    layer4_outputs(8958) <= not((layer3_outputs(4380)) xor (layer3_outputs(4561)));
    layer4_outputs(8959) <= not(layer3_outputs(1404)) or (layer3_outputs(5930));
    layer4_outputs(8960) <= layer3_outputs(1583);
    layer4_outputs(8961) <= not(layer3_outputs(6530));
    layer4_outputs(8962) <= layer3_outputs(789);
    layer4_outputs(8963) <= not(layer3_outputs(8624)) or (layer3_outputs(3850));
    layer4_outputs(8964) <= layer3_outputs(4660);
    layer4_outputs(8965) <= layer3_outputs(5122);
    layer4_outputs(8966) <= not((layer3_outputs(9701)) xor (layer3_outputs(7826)));
    layer4_outputs(8967) <= not(layer3_outputs(1217));
    layer4_outputs(8968) <= not(layer3_outputs(1618)) or (layer3_outputs(1799));
    layer4_outputs(8969) <= layer3_outputs(6003);
    layer4_outputs(8970) <= not((layer3_outputs(8380)) xor (layer3_outputs(3881)));
    layer4_outputs(8971) <= not(layer3_outputs(9255));
    layer4_outputs(8972) <= (layer3_outputs(2608)) and not (layer3_outputs(1206));
    layer4_outputs(8973) <= not(layer3_outputs(656));
    layer4_outputs(8974) <= not((layer3_outputs(7125)) and (layer3_outputs(732)));
    layer4_outputs(8975) <= (layer3_outputs(5966)) and not (layer3_outputs(4639));
    layer4_outputs(8976) <= (layer3_outputs(8775)) or (layer3_outputs(3583));
    layer4_outputs(8977) <= not(layer3_outputs(9239));
    layer4_outputs(8978) <= not(layer3_outputs(9989));
    layer4_outputs(8979) <= not(layer3_outputs(7265)) or (layer3_outputs(6490));
    layer4_outputs(8980) <= not(layer3_outputs(8035));
    layer4_outputs(8981) <= not(layer3_outputs(7279)) or (layer3_outputs(5794));
    layer4_outputs(8982) <= (layer3_outputs(6597)) or (layer3_outputs(728));
    layer4_outputs(8983) <= not(layer3_outputs(7462));
    layer4_outputs(8984) <= not((layer3_outputs(9455)) xor (layer3_outputs(8086)));
    layer4_outputs(8985) <= not((layer3_outputs(5697)) and (layer3_outputs(6822)));
    layer4_outputs(8986) <= layer3_outputs(6028);
    layer4_outputs(8987) <= (layer3_outputs(10208)) and not (layer3_outputs(7209));
    layer4_outputs(8988) <= not(layer3_outputs(5848)) or (layer3_outputs(7358));
    layer4_outputs(8989) <= layer3_outputs(3749);
    layer4_outputs(8990) <= (layer3_outputs(542)) xor (layer3_outputs(5233));
    layer4_outputs(8991) <= (layer3_outputs(7599)) and not (layer3_outputs(5939));
    layer4_outputs(8992) <= not(layer3_outputs(8819));
    layer4_outputs(8993) <= not((layer3_outputs(6303)) xor (layer3_outputs(1239)));
    layer4_outputs(8994) <= not(layer3_outputs(6478));
    layer4_outputs(8995) <= (layer3_outputs(718)) or (layer3_outputs(6483));
    layer4_outputs(8996) <= not(layer3_outputs(7637)) or (layer3_outputs(2140));
    layer4_outputs(8997) <= (layer3_outputs(1867)) xor (layer3_outputs(9676));
    layer4_outputs(8998) <= not(layer3_outputs(7374));
    layer4_outputs(8999) <= not(layer3_outputs(2078));
    layer4_outputs(9000) <= layer3_outputs(1923);
    layer4_outputs(9001) <= (layer3_outputs(9392)) and not (layer3_outputs(4415));
    layer4_outputs(9002) <= (layer3_outputs(721)) and not (layer3_outputs(2735));
    layer4_outputs(9003) <= not(layer3_outputs(6826));
    layer4_outputs(9004) <= not((layer3_outputs(531)) and (layer3_outputs(7506)));
    layer4_outputs(9005) <= '1';
    layer4_outputs(9006) <= not(layer3_outputs(1811));
    layer4_outputs(9007) <= (layer3_outputs(5049)) or (layer3_outputs(1521));
    layer4_outputs(9008) <= (layer3_outputs(9857)) and not (layer3_outputs(9935));
    layer4_outputs(9009) <= not(layer3_outputs(914));
    layer4_outputs(9010) <= not(layer3_outputs(8439));
    layer4_outputs(9011) <= (layer3_outputs(7336)) or (layer3_outputs(3561));
    layer4_outputs(9012) <= not(layer3_outputs(5497)) or (layer3_outputs(5972));
    layer4_outputs(9013) <= not(layer3_outputs(9823));
    layer4_outputs(9014) <= not(layer3_outputs(2108)) or (layer3_outputs(8840));
    layer4_outputs(9015) <= (layer3_outputs(9997)) and (layer3_outputs(5122));
    layer4_outputs(9016) <= not(layer3_outputs(5028));
    layer4_outputs(9017) <= layer3_outputs(6916);
    layer4_outputs(9018) <= not((layer3_outputs(1176)) xor (layer3_outputs(4423)));
    layer4_outputs(9019) <= not(layer3_outputs(6759));
    layer4_outputs(9020) <= layer3_outputs(5164);
    layer4_outputs(9021) <= layer3_outputs(7235);
    layer4_outputs(9022) <= (layer3_outputs(718)) xor (layer3_outputs(6111));
    layer4_outputs(9023) <= not((layer3_outputs(5876)) xor (layer3_outputs(10209)));
    layer4_outputs(9024) <= layer3_outputs(7242);
    layer4_outputs(9025) <= not(layer3_outputs(5192)) or (layer3_outputs(576));
    layer4_outputs(9026) <= not((layer3_outputs(5868)) or (layer3_outputs(5712)));
    layer4_outputs(9027) <= not(layer3_outputs(565)) or (layer3_outputs(4041));
    layer4_outputs(9028) <= (layer3_outputs(166)) xor (layer3_outputs(2151));
    layer4_outputs(9029) <= not((layer3_outputs(8388)) and (layer3_outputs(5654)));
    layer4_outputs(9030) <= (layer3_outputs(1564)) or (layer3_outputs(3542));
    layer4_outputs(9031) <= layer3_outputs(4616);
    layer4_outputs(9032) <= (layer3_outputs(5965)) and (layer3_outputs(7906));
    layer4_outputs(9033) <= (layer3_outputs(5630)) and (layer3_outputs(6356));
    layer4_outputs(9034) <= layer3_outputs(8621);
    layer4_outputs(9035) <= not(layer3_outputs(3069)) or (layer3_outputs(3664));
    layer4_outputs(9036) <= layer3_outputs(386);
    layer4_outputs(9037) <= layer3_outputs(124);
    layer4_outputs(9038) <= not(layer3_outputs(284));
    layer4_outputs(9039) <= not(layer3_outputs(5042));
    layer4_outputs(9040) <= not(layer3_outputs(84)) or (layer3_outputs(5489));
    layer4_outputs(9041) <= (layer3_outputs(9283)) xor (layer3_outputs(2747));
    layer4_outputs(9042) <= layer3_outputs(3957);
    layer4_outputs(9043) <= layer3_outputs(266);
    layer4_outputs(9044) <= layer3_outputs(8237);
    layer4_outputs(9045) <= (layer3_outputs(8438)) xor (layer3_outputs(7364));
    layer4_outputs(9046) <= (layer3_outputs(5512)) or (layer3_outputs(5134));
    layer4_outputs(9047) <= (layer3_outputs(1772)) xor (layer3_outputs(3063));
    layer4_outputs(9048) <= not(layer3_outputs(83));
    layer4_outputs(9049) <= layer3_outputs(9861);
    layer4_outputs(9050) <= not((layer3_outputs(2949)) and (layer3_outputs(2427)));
    layer4_outputs(9051) <= layer3_outputs(8420);
    layer4_outputs(9052) <= not(layer3_outputs(6542));
    layer4_outputs(9053) <= (layer3_outputs(1269)) and not (layer3_outputs(7670));
    layer4_outputs(9054) <= not(layer3_outputs(6442));
    layer4_outputs(9055) <= not(layer3_outputs(820));
    layer4_outputs(9056) <= not(layer3_outputs(2899));
    layer4_outputs(9057) <= not(layer3_outputs(3496));
    layer4_outputs(9058) <= not(layer3_outputs(2242)) or (layer3_outputs(3760));
    layer4_outputs(9059) <= not(layer3_outputs(9210));
    layer4_outputs(9060) <= not(layer3_outputs(3634)) or (layer3_outputs(4694));
    layer4_outputs(9061) <= not((layer3_outputs(6142)) and (layer3_outputs(5811)));
    layer4_outputs(9062) <= not(layer3_outputs(6799));
    layer4_outputs(9063) <= not((layer3_outputs(9531)) xor (layer3_outputs(5394)));
    layer4_outputs(9064) <= layer3_outputs(2799);
    layer4_outputs(9065) <= not(layer3_outputs(1978));
    layer4_outputs(9066) <= not((layer3_outputs(1019)) or (layer3_outputs(5287)));
    layer4_outputs(9067) <= not(layer3_outputs(9260));
    layer4_outputs(9068) <= not(layer3_outputs(6806)) or (layer3_outputs(2058));
    layer4_outputs(9069) <= not((layer3_outputs(9877)) and (layer3_outputs(7317)));
    layer4_outputs(9070) <= layer3_outputs(1598);
    layer4_outputs(9071) <= layer3_outputs(3994);
    layer4_outputs(9072) <= layer3_outputs(7620);
    layer4_outputs(9073) <= not(layer3_outputs(9054));
    layer4_outputs(9074) <= not(layer3_outputs(3287));
    layer4_outputs(9075) <= layer3_outputs(4688);
    layer4_outputs(9076) <= not(layer3_outputs(4812));
    layer4_outputs(9077) <= layer3_outputs(7888);
    layer4_outputs(9078) <= layer3_outputs(9044);
    layer4_outputs(9079) <= (layer3_outputs(6568)) and not (layer3_outputs(1959));
    layer4_outputs(9080) <= layer3_outputs(2848);
    layer4_outputs(9081) <= not((layer3_outputs(8528)) and (layer3_outputs(2119)));
    layer4_outputs(9082) <= (layer3_outputs(9398)) xor (layer3_outputs(543));
    layer4_outputs(9083) <= '0';
    layer4_outputs(9084) <= not(layer3_outputs(2169));
    layer4_outputs(9085) <= not(layer3_outputs(6736));
    layer4_outputs(9086) <= layer3_outputs(3149);
    layer4_outputs(9087) <= not(layer3_outputs(5505));
    layer4_outputs(9088) <= not(layer3_outputs(700));
    layer4_outputs(9089) <= not(layer3_outputs(8384));
    layer4_outputs(9090) <= not(layer3_outputs(682));
    layer4_outputs(9091) <= not((layer3_outputs(1265)) and (layer3_outputs(4067)));
    layer4_outputs(9092) <= (layer3_outputs(5293)) xor (layer3_outputs(940));
    layer4_outputs(9093) <= (layer3_outputs(4884)) and not (layer3_outputs(460));
    layer4_outputs(9094) <= not(layer3_outputs(10037)) or (layer3_outputs(5868));
    layer4_outputs(9095) <= not(layer3_outputs(8623)) or (layer3_outputs(8526));
    layer4_outputs(9096) <= not((layer3_outputs(3906)) xor (layer3_outputs(1025)));
    layer4_outputs(9097) <= layer3_outputs(567);
    layer4_outputs(9098) <= layer3_outputs(8234);
    layer4_outputs(9099) <= (layer3_outputs(6945)) and (layer3_outputs(8307));
    layer4_outputs(9100) <= layer3_outputs(3746);
    layer4_outputs(9101) <= not(layer3_outputs(3310)) or (layer3_outputs(4054));
    layer4_outputs(9102) <= (layer3_outputs(8536)) and (layer3_outputs(1612));
    layer4_outputs(9103) <= not(layer3_outputs(5160)) or (layer3_outputs(5889));
    layer4_outputs(9104) <= layer3_outputs(8166);
    layer4_outputs(9105) <= (layer3_outputs(4455)) and not (layer3_outputs(3469));
    layer4_outputs(9106) <= not(layer3_outputs(9214)) or (layer3_outputs(3721));
    layer4_outputs(9107) <= (layer3_outputs(4637)) xor (layer3_outputs(4851));
    layer4_outputs(9108) <= not((layer3_outputs(6661)) or (layer3_outputs(6699)));
    layer4_outputs(9109) <= (layer3_outputs(427)) and (layer3_outputs(7082));
    layer4_outputs(9110) <= not(layer3_outputs(2347)) or (layer3_outputs(7658));
    layer4_outputs(9111) <= (layer3_outputs(6466)) and not (layer3_outputs(2028));
    layer4_outputs(9112) <= layer3_outputs(6457);
    layer4_outputs(9113) <= not((layer3_outputs(4222)) and (layer3_outputs(3275)));
    layer4_outputs(9114) <= not((layer3_outputs(1231)) xor (layer3_outputs(8329)));
    layer4_outputs(9115) <= layer3_outputs(8322);
    layer4_outputs(9116) <= not(layer3_outputs(6816));
    layer4_outputs(9117) <= layer3_outputs(8917);
    layer4_outputs(9118) <= not((layer3_outputs(4325)) or (layer3_outputs(2753)));
    layer4_outputs(9119) <= layer3_outputs(2905);
    layer4_outputs(9120) <= not((layer3_outputs(9646)) or (layer3_outputs(7770)));
    layer4_outputs(9121) <= not(layer3_outputs(9579));
    layer4_outputs(9122) <= layer3_outputs(2782);
    layer4_outputs(9123) <= not(layer3_outputs(704));
    layer4_outputs(9124) <= (layer3_outputs(1492)) xor (layer3_outputs(9333));
    layer4_outputs(9125) <= not(layer3_outputs(4908));
    layer4_outputs(9126) <= layer3_outputs(9782);
    layer4_outputs(9127) <= layer3_outputs(4070);
    layer4_outputs(9128) <= not(layer3_outputs(2359)) or (layer3_outputs(4871));
    layer4_outputs(9129) <= layer3_outputs(6296);
    layer4_outputs(9130) <= not((layer3_outputs(4614)) or (layer3_outputs(1669)));
    layer4_outputs(9131) <= (layer3_outputs(4042)) and not (layer3_outputs(736));
    layer4_outputs(9132) <= layer3_outputs(5146);
    layer4_outputs(9133) <= not(layer3_outputs(6086));
    layer4_outputs(9134) <= not(layer3_outputs(9456));
    layer4_outputs(9135) <= layer3_outputs(7945);
    layer4_outputs(9136) <= (layer3_outputs(4621)) and not (layer3_outputs(2760));
    layer4_outputs(9137) <= not((layer3_outputs(2553)) and (layer3_outputs(6036)));
    layer4_outputs(9138) <= not(layer3_outputs(965));
    layer4_outputs(9139) <= layer3_outputs(2660);
    layer4_outputs(9140) <= (layer3_outputs(8274)) and not (layer3_outputs(6515));
    layer4_outputs(9141) <= layer3_outputs(3794);
    layer4_outputs(9142) <= not(layer3_outputs(5312)) or (layer3_outputs(938));
    layer4_outputs(9143) <= layer3_outputs(8797);
    layer4_outputs(9144) <= layer3_outputs(927);
    layer4_outputs(9145) <= (layer3_outputs(7879)) xor (layer3_outputs(6985));
    layer4_outputs(9146) <= layer3_outputs(7627);
    layer4_outputs(9147) <= not((layer3_outputs(163)) xor (layer3_outputs(3455)));
    layer4_outputs(9148) <= not(layer3_outputs(5219));
    layer4_outputs(9149) <= (layer3_outputs(1400)) or (layer3_outputs(1189));
    layer4_outputs(9150) <= (layer3_outputs(7861)) and not (layer3_outputs(3926));
    layer4_outputs(9151) <= layer3_outputs(7994);
    layer4_outputs(9152) <= not(layer3_outputs(319));
    layer4_outputs(9153) <= not(layer3_outputs(7276));
    layer4_outputs(9154) <= not(layer3_outputs(9245));
    layer4_outputs(9155) <= (layer3_outputs(5852)) and not (layer3_outputs(871));
    layer4_outputs(9156) <= (layer3_outputs(1886)) and (layer3_outputs(4382));
    layer4_outputs(9157) <= not(layer3_outputs(4813));
    layer4_outputs(9158) <= (layer3_outputs(1617)) and (layer3_outputs(5111));
    layer4_outputs(9159) <= not(layer3_outputs(6134));
    layer4_outputs(9160) <= layer3_outputs(3509);
    layer4_outputs(9161) <= not(layer3_outputs(6403));
    layer4_outputs(9162) <= layer3_outputs(8211);
    layer4_outputs(9163) <= layer3_outputs(3622);
    layer4_outputs(9164) <= not(layer3_outputs(7321));
    layer4_outputs(9165) <= layer3_outputs(2876);
    layer4_outputs(9166) <= not(layer3_outputs(420));
    layer4_outputs(9167) <= layer3_outputs(9558);
    layer4_outputs(9168) <= not(layer3_outputs(10098)) or (layer3_outputs(823));
    layer4_outputs(9169) <= (layer3_outputs(9958)) and not (layer3_outputs(5247));
    layer4_outputs(9170) <= (layer3_outputs(9340)) and (layer3_outputs(1779));
    layer4_outputs(9171) <= (layer3_outputs(774)) xor (layer3_outputs(2122));
    layer4_outputs(9172) <= not(layer3_outputs(8311));
    layer4_outputs(9173) <= not(layer3_outputs(6654));
    layer4_outputs(9174) <= (layer3_outputs(141)) xor (layer3_outputs(7804));
    layer4_outputs(9175) <= layer3_outputs(10169);
    layer4_outputs(9176) <= not((layer3_outputs(6749)) xor (layer3_outputs(1078)));
    layer4_outputs(9177) <= layer3_outputs(3942);
    layer4_outputs(9178) <= not(layer3_outputs(7572));
    layer4_outputs(9179) <= (layer3_outputs(6463)) and not (layer3_outputs(2606));
    layer4_outputs(9180) <= not(layer3_outputs(7993)) or (layer3_outputs(6598));
    layer4_outputs(9181) <= not(layer3_outputs(1351));
    layer4_outputs(9182) <= not(layer3_outputs(5745));
    layer4_outputs(9183) <= not(layer3_outputs(1229));
    layer4_outputs(9184) <= layer3_outputs(2499);
    layer4_outputs(9185) <= not(layer3_outputs(6897));
    layer4_outputs(9186) <= layer3_outputs(6912);
    layer4_outputs(9187) <= not((layer3_outputs(3039)) and (layer3_outputs(1362)));
    layer4_outputs(9188) <= not(layer3_outputs(8356)) or (layer3_outputs(1092));
    layer4_outputs(9189) <= layer3_outputs(8822);
    layer4_outputs(9190) <= layer3_outputs(5334);
    layer4_outputs(9191) <= not((layer3_outputs(491)) or (layer3_outputs(5696)));
    layer4_outputs(9192) <= not(layer3_outputs(7198));
    layer4_outputs(9193) <= not(layer3_outputs(10216));
    layer4_outputs(9194) <= layer3_outputs(3159);
    layer4_outputs(9195) <= not(layer3_outputs(8587)) or (layer3_outputs(4373));
    layer4_outputs(9196) <= not(layer3_outputs(3923));
    layer4_outputs(9197) <= not(layer3_outputs(2336));
    layer4_outputs(9198) <= layer3_outputs(1179);
    layer4_outputs(9199) <= layer3_outputs(4861);
    layer4_outputs(9200) <= not((layer3_outputs(3914)) and (layer3_outputs(1715)));
    layer4_outputs(9201) <= (layer3_outputs(6969)) and not (layer3_outputs(8482));
    layer4_outputs(9202) <= layer3_outputs(8249);
    layer4_outputs(9203) <= layer3_outputs(4556);
    layer4_outputs(9204) <= not((layer3_outputs(1743)) xor (layer3_outputs(6349)));
    layer4_outputs(9205) <= layer3_outputs(1215);
    layer4_outputs(9206) <= (layer3_outputs(2056)) or (layer3_outputs(4723));
    layer4_outputs(9207) <= not((layer3_outputs(9012)) and (layer3_outputs(7695)));
    layer4_outputs(9208) <= not(layer3_outputs(2228)) or (layer3_outputs(4063));
    layer4_outputs(9209) <= (layer3_outputs(1853)) and (layer3_outputs(5063));
    layer4_outputs(9210) <= layer3_outputs(9155);
    layer4_outputs(9211) <= not((layer3_outputs(4634)) xor (layer3_outputs(6762)));
    layer4_outputs(9212) <= (layer3_outputs(120)) xor (layer3_outputs(2850));
    layer4_outputs(9213) <= layer3_outputs(4383);
    layer4_outputs(9214) <= (layer3_outputs(4443)) and (layer3_outputs(7558));
    layer4_outputs(9215) <= not(layer3_outputs(6438)) or (layer3_outputs(8948));
    layer4_outputs(9216) <= (layer3_outputs(2784)) and (layer3_outputs(5991));
    layer4_outputs(9217) <= not((layer3_outputs(2001)) and (layer3_outputs(2431)));
    layer4_outputs(9218) <= layer3_outputs(6648);
    layer4_outputs(9219) <= layer3_outputs(4075);
    layer4_outputs(9220) <= not(layer3_outputs(5049));
    layer4_outputs(9221) <= layer3_outputs(8892);
    layer4_outputs(9222) <= not((layer3_outputs(2546)) xor (layer3_outputs(9761)));
    layer4_outputs(9223) <= layer3_outputs(9834);
    layer4_outputs(9224) <= (layer3_outputs(914)) and not (layer3_outputs(2232));
    layer4_outputs(9225) <= not(layer3_outputs(9014));
    layer4_outputs(9226) <= layer3_outputs(9869);
    layer4_outputs(9227) <= layer3_outputs(6011);
    layer4_outputs(9228) <= not(layer3_outputs(6832));
    layer4_outputs(9229) <= layer3_outputs(9297);
    layer4_outputs(9230) <= layer3_outputs(10055);
    layer4_outputs(9231) <= layer3_outputs(2571);
    layer4_outputs(9232) <= not(layer3_outputs(7130));
    layer4_outputs(9233) <= not(layer3_outputs(7015));
    layer4_outputs(9234) <= layer3_outputs(7258);
    layer4_outputs(9235) <= not((layer3_outputs(4350)) xor (layer3_outputs(8427)));
    layer4_outputs(9236) <= layer3_outputs(5663);
    layer4_outputs(9237) <= layer3_outputs(9033);
    layer4_outputs(9238) <= not(layer3_outputs(1101)) or (layer3_outputs(5369));
    layer4_outputs(9239) <= (layer3_outputs(9113)) or (layer3_outputs(5419));
    layer4_outputs(9240) <= layer3_outputs(6488);
    layer4_outputs(9241) <= (layer3_outputs(10220)) and (layer3_outputs(9852));
    layer4_outputs(9242) <= not(layer3_outputs(5969));
    layer4_outputs(9243) <= not(layer3_outputs(2705));
    layer4_outputs(9244) <= layer3_outputs(7426);
    layer4_outputs(9245) <= not(layer3_outputs(1902));
    layer4_outputs(9246) <= layer3_outputs(3117);
    layer4_outputs(9247) <= (layer3_outputs(1307)) xor (layer3_outputs(6096));
    layer4_outputs(9248) <= not(layer3_outputs(5388));
    layer4_outputs(9249) <= layer3_outputs(7575);
    layer4_outputs(9250) <= (layer3_outputs(8609)) or (layer3_outputs(3645));
    layer4_outputs(9251) <= (layer3_outputs(9496)) xor (layer3_outputs(9651));
    layer4_outputs(9252) <= layer3_outputs(2880);
    layer4_outputs(9253) <= layer3_outputs(8561);
    layer4_outputs(9254) <= not(layer3_outputs(4915)) or (layer3_outputs(1315));
    layer4_outputs(9255) <= (layer3_outputs(9108)) xor (layer3_outputs(2671));
    layer4_outputs(9256) <= layer3_outputs(9267);
    layer4_outputs(9257) <= (layer3_outputs(2956)) xor (layer3_outputs(8352));
    layer4_outputs(9258) <= (layer3_outputs(9508)) or (layer3_outputs(4583));
    layer4_outputs(9259) <= layer3_outputs(4759);
    layer4_outputs(9260) <= not(layer3_outputs(4763)) or (layer3_outputs(2907));
    layer4_outputs(9261) <= not(layer3_outputs(6973));
    layer4_outputs(9262) <= not((layer3_outputs(685)) xor (layer3_outputs(212)));
    layer4_outputs(9263) <= layer3_outputs(1699);
    layer4_outputs(9264) <= layer3_outputs(6500);
    layer4_outputs(9265) <= (layer3_outputs(7609)) xor (layer3_outputs(2899));
    layer4_outputs(9266) <= (layer3_outputs(3474)) and (layer3_outputs(4224));
    layer4_outputs(9267) <= layer3_outputs(2973);
    layer4_outputs(9268) <= not((layer3_outputs(8494)) xor (layer3_outputs(8786)));
    layer4_outputs(9269) <= not(layer3_outputs(123));
    layer4_outputs(9270) <= not(layer3_outputs(9336));
    layer4_outputs(9271) <= not(layer3_outputs(9601));
    layer4_outputs(9272) <= not(layer3_outputs(2505)) or (layer3_outputs(7493));
    layer4_outputs(9273) <= layer3_outputs(9406);
    layer4_outputs(9274) <= not((layer3_outputs(2847)) and (layer3_outputs(9313)));
    layer4_outputs(9275) <= (layer3_outputs(234)) and not (layer3_outputs(1534));
    layer4_outputs(9276) <= (layer3_outputs(5931)) and not (layer3_outputs(3315));
    layer4_outputs(9277) <= layer3_outputs(928);
    layer4_outputs(9278) <= (layer3_outputs(6176)) or (layer3_outputs(1953));
    layer4_outputs(9279) <= layer3_outputs(2475);
    layer4_outputs(9280) <= layer3_outputs(5399);
    layer4_outputs(9281) <= layer3_outputs(9817);
    layer4_outputs(9282) <= not((layer3_outputs(2884)) xor (layer3_outputs(8528)));
    layer4_outputs(9283) <= not(layer3_outputs(599));
    layer4_outputs(9284) <= layer3_outputs(8503);
    layer4_outputs(9285) <= layer3_outputs(8049);
    layer4_outputs(9286) <= layer3_outputs(1083);
    layer4_outputs(9287) <= not((layer3_outputs(5128)) xor (layer3_outputs(2016)));
    layer4_outputs(9288) <= not(layer3_outputs(893)) or (layer3_outputs(4944));
    layer4_outputs(9289) <= layer3_outputs(6457);
    layer4_outputs(9290) <= not(layer3_outputs(6930));
    layer4_outputs(9291) <= not(layer3_outputs(3905)) or (layer3_outputs(7187));
    layer4_outputs(9292) <= not(layer3_outputs(8020));
    layer4_outputs(9293) <= not((layer3_outputs(6476)) and (layer3_outputs(7628)));
    layer4_outputs(9294) <= layer3_outputs(9268);
    layer4_outputs(9295) <= layer3_outputs(6526);
    layer4_outputs(9296) <= not(layer3_outputs(9098)) or (layer3_outputs(4265));
    layer4_outputs(9297) <= layer3_outputs(6290);
    layer4_outputs(9298) <= not(layer3_outputs(8916));
    layer4_outputs(9299) <= not(layer3_outputs(6189));
    layer4_outputs(9300) <= (layer3_outputs(6016)) and (layer3_outputs(5427));
    layer4_outputs(9301) <= not(layer3_outputs(8882)) or (layer3_outputs(1858));
    layer4_outputs(9302) <= (layer3_outputs(5533)) xor (layer3_outputs(5442));
    layer4_outputs(9303) <= (layer3_outputs(5103)) and (layer3_outputs(2917));
    layer4_outputs(9304) <= layer3_outputs(9010);
    layer4_outputs(9305) <= layer3_outputs(6394);
    layer4_outputs(9306) <= not(layer3_outputs(7345));
    layer4_outputs(9307) <= (layer3_outputs(7871)) xor (layer3_outputs(3230));
    layer4_outputs(9308) <= (layer3_outputs(6949)) or (layer3_outputs(3832));
    layer4_outputs(9309) <= (layer3_outputs(6032)) xor (layer3_outputs(7904));
    layer4_outputs(9310) <= not((layer3_outputs(9507)) xor (layer3_outputs(2648)));
    layer4_outputs(9311) <= layer3_outputs(7420);
    layer4_outputs(9312) <= not(layer3_outputs(7564));
    layer4_outputs(9313) <= layer3_outputs(8527);
    layer4_outputs(9314) <= (layer3_outputs(5466)) and not (layer3_outputs(1027));
    layer4_outputs(9315) <= (layer3_outputs(6295)) and not (layer3_outputs(2152));
    layer4_outputs(9316) <= layer3_outputs(7354);
    layer4_outputs(9317) <= layer3_outputs(6256);
    layer4_outputs(9318) <= (layer3_outputs(4999)) and not (layer3_outputs(3964));
    layer4_outputs(9319) <= not(layer3_outputs(6103));
    layer4_outputs(9320) <= (layer3_outputs(6566)) xor (layer3_outputs(7392));
    layer4_outputs(9321) <= not(layer3_outputs(8398));
    layer4_outputs(9322) <= not((layer3_outputs(4845)) or (layer3_outputs(7939)));
    layer4_outputs(9323) <= not(layer3_outputs(4248));
    layer4_outputs(9324) <= not((layer3_outputs(4977)) xor (layer3_outputs(1292)));
    layer4_outputs(9325) <= not(layer3_outputs(3397));
    layer4_outputs(9326) <= (layer3_outputs(3728)) xor (layer3_outputs(6641));
    layer4_outputs(9327) <= (layer3_outputs(9000)) and not (layer3_outputs(5261));
    layer4_outputs(9328) <= (layer3_outputs(6469)) or (layer3_outputs(7864));
    layer4_outputs(9329) <= not(layer3_outputs(1576));
    layer4_outputs(9330) <= not(layer3_outputs(1075));
    layer4_outputs(9331) <= layer3_outputs(2669);
    layer4_outputs(9332) <= layer3_outputs(741);
    layer4_outputs(9333) <= not((layer3_outputs(9003)) xor (layer3_outputs(6231)));
    layer4_outputs(9334) <= layer3_outputs(5920);
    layer4_outputs(9335) <= (layer3_outputs(3162)) xor (layer3_outputs(8363));
    layer4_outputs(9336) <= not(layer3_outputs(934));
    layer4_outputs(9337) <= (layer3_outputs(551)) and not (layer3_outputs(7396));
    layer4_outputs(9338) <= (layer3_outputs(5440)) or (layer3_outputs(1240));
    layer4_outputs(9339) <= layer3_outputs(5893);
    layer4_outputs(9340) <= not(layer3_outputs(889));
    layer4_outputs(9341) <= layer3_outputs(10006);
    layer4_outputs(9342) <= not((layer3_outputs(8582)) or (layer3_outputs(5674)));
    layer4_outputs(9343) <= not(layer3_outputs(684));
    layer4_outputs(9344) <= layer3_outputs(3576);
    layer4_outputs(9345) <= layer3_outputs(324);
    layer4_outputs(9346) <= not(layer3_outputs(4607));
    layer4_outputs(9347) <= not(layer3_outputs(1057));
    layer4_outputs(9348) <= not(layer3_outputs(1692)) or (layer3_outputs(5036));
    layer4_outputs(9349) <= not(layer3_outputs(8470));
    layer4_outputs(9350) <= (layer3_outputs(6518)) and (layer3_outputs(6922));
    layer4_outputs(9351) <= (layer3_outputs(7446)) and not (layer3_outputs(4360));
    layer4_outputs(9352) <= not(layer3_outputs(3983));
    layer4_outputs(9353) <= layer3_outputs(5919);
    layer4_outputs(9354) <= (layer3_outputs(8522)) and not (layer3_outputs(4664));
    layer4_outputs(9355) <= layer3_outputs(3652);
    layer4_outputs(9356) <= not(layer3_outputs(37)) or (layer3_outputs(8973));
    layer4_outputs(9357) <= not(layer3_outputs(1986));
    layer4_outputs(9358) <= (layer3_outputs(8325)) and not (layer3_outputs(1406));
    layer4_outputs(9359) <= (layer3_outputs(7710)) xor (layer3_outputs(8823));
    layer4_outputs(9360) <= layer3_outputs(3535);
    layer4_outputs(9361) <= (layer3_outputs(4428)) and not (layer3_outputs(5232));
    layer4_outputs(9362) <= layer3_outputs(8419);
    layer4_outputs(9363) <= layer3_outputs(4432);
    layer4_outputs(9364) <= (layer3_outputs(4282)) and not (layer3_outputs(1198));
    layer4_outputs(9365) <= not(layer3_outputs(4563));
    layer4_outputs(9366) <= (layer3_outputs(6062)) or (layer3_outputs(6114));
    layer4_outputs(9367) <= (layer3_outputs(6505)) and not (layer3_outputs(1013));
    layer4_outputs(9368) <= layer3_outputs(2540);
    layer4_outputs(9369) <= (layer3_outputs(1512)) xor (layer3_outputs(2007));
    layer4_outputs(9370) <= layer3_outputs(1151);
    layer4_outputs(9371) <= not((layer3_outputs(1931)) or (layer3_outputs(8803)));
    layer4_outputs(9372) <= (layer3_outputs(9374)) and not (layer3_outputs(7287));
    layer4_outputs(9373) <= not((layer3_outputs(339)) xor (layer3_outputs(1879)));
    layer4_outputs(9374) <= (layer3_outputs(1654)) and not (layer3_outputs(893));
    layer4_outputs(9375) <= '0';
    layer4_outputs(9376) <= not((layer3_outputs(3894)) xor (layer3_outputs(7633)));
    layer4_outputs(9377) <= (layer3_outputs(6347)) xor (layer3_outputs(8766));
    layer4_outputs(9378) <= layer3_outputs(9502);
    layer4_outputs(9379) <= not(layer3_outputs(8491)) or (layer3_outputs(4909));
    layer4_outputs(9380) <= not(layer3_outputs(5873));
    layer4_outputs(9381) <= (layer3_outputs(6337)) and not (layer3_outputs(7948));
    layer4_outputs(9382) <= not(layer3_outputs(345));
    layer4_outputs(9383) <= (layer3_outputs(3107)) or (layer3_outputs(1301));
    layer4_outputs(9384) <= layer3_outputs(7585);
    layer4_outputs(9385) <= (layer3_outputs(2696)) xor (layer3_outputs(3550));
    layer4_outputs(9386) <= not((layer3_outputs(9048)) xor (layer3_outputs(8128)));
    layer4_outputs(9387) <= not(layer3_outputs(9488)) or (layer3_outputs(6705));
    layer4_outputs(9388) <= not(layer3_outputs(5724));
    layer4_outputs(9389) <= not((layer3_outputs(5160)) or (layer3_outputs(123)));
    layer4_outputs(9390) <= not(layer3_outputs(10030));
    layer4_outputs(9391) <= layer3_outputs(7559);
    layer4_outputs(9392) <= not(layer3_outputs(8510)) or (layer3_outputs(9243));
    layer4_outputs(9393) <= not((layer3_outputs(4610)) xor (layer3_outputs(2309)));
    layer4_outputs(9394) <= (layer3_outputs(1678)) or (layer3_outputs(8820));
    layer4_outputs(9395) <= (layer3_outputs(8998)) xor (layer3_outputs(5694));
    layer4_outputs(9396) <= (layer3_outputs(6162)) and not (layer3_outputs(2874));
    layer4_outputs(9397) <= layer3_outputs(2968);
    layer4_outputs(9398) <= layer3_outputs(289);
    layer4_outputs(9399) <= (layer3_outputs(5677)) or (layer3_outputs(5843));
    layer4_outputs(9400) <= layer3_outputs(8658);
    layer4_outputs(9401) <= not(layer3_outputs(2155));
    layer4_outputs(9402) <= not(layer3_outputs(7739));
    layer4_outputs(9403) <= (layer3_outputs(6555)) xor (layer3_outputs(5075));
    layer4_outputs(9404) <= layer3_outputs(3056);
    layer4_outputs(9405) <= layer3_outputs(7747);
    layer4_outputs(9406) <= layer3_outputs(1888);
    layer4_outputs(9407) <= layer3_outputs(9427);
    layer4_outputs(9408) <= (layer3_outputs(1757)) and not (layer3_outputs(6199));
    layer4_outputs(9409) <= (layer3_outputs(9434)) xor (layer3_outputs(2604));
    layer4_outputs(9410) <= (layer3_outputs(1716)) or (layer3_outputs(7987));
    layer4_outputs(9411) <= not(layer3_outputs(2988));
    layer4_outputs(9412) <= not(layer3_outputs(1240));
    layer4_outputs(9413) <= not(layer3_outputs(6659));
    layer4_outputs(9414) <= not(layer3_outputs(8552));
    layer4_outputs(9415) <= layer3_outputs(4168);
    layer4_outputs(9416) <= (layer3_outputs(7528)) xor (layer3_outputs(4537));
    layer4_outputs(9417) <= layer3_outputs(525);
    layer4_outputs(9418) <= not(layer3_outputs(3332));
    layer4_outputs(9419) <= '1';
    layer4_outputs(9420) <= layer3_outputs(1614);
    layer4_outputs(9421) <= not((layer3_outputs(3636)) xor (layer3_outputs(2096)));
    layer4_outputs(9422) <= layer3_outputs(7153);
    layer4_outputs(9423) <= (layer3_outputs(4765)) and (layer3_outputs(2922));
    layer4_outputs(9424) <= not(layer3_outputs(1777));
    layer4_outputs(9425) <= not(layer3_outputs(4154));
    layer4_outputs(9426) <= (layer3_outputs(3223)) or (layer3_outputs(1733));
    layer4_outputs(9427) <= not(layer3_outputs(8835)) or (layer3_outputs(5288));
    layer4_outputs(9428) <= not((layer3_outputs(8661)) or (layer3_outputs(6731)));
    layer4_outputs(9429) <= layer3_outputs(972);
    layer4_outputs(9430) <= layer3_outputs(9821);
    layer4_outputs(9431) <= not(layer3_outputs(1303));
    layer4_outputs(9432) <= not(layer3_outputs(505));
    layer4_outputs(9433) <= layer3_outputs(5494);
    layer4_outputs(9434) <= not(layer3_outputs(8385));
    layer4_outputs(9435) <= not(layer3_outputs(1189));
    layer4_outputs(9436) <= layer3_outputs(6609);
    layer4_outputs(9437) <= layer3_outputs(962);
    layer4_outputs(9438) <= not(layer3_outputs(1270));
    layer4_outputs(9439) <= layer3_outputs(1074);
    layer4_outputs(9440) <= layer3_outputs(9595);
    layer4_outputs(9441) <= not(layer3_outputs(9083));
    layer4_outputs(9442) <= (layer3_outputs(10197)) or (layer3_outputs(5766));
    layer4_outputs(9443) <= (layer3_outputs(340)) xor (layer3_outputs(8338));
    layer4_outputs(9444) <= layer3_outputs(9089);
    layer4_outputs(9445) <= (layer3_outputs(10223)) and (layer3_outputs(4462));
    layer4_outputs(9446) <= not(layer3_outputs(9228)) or (layer3_outputs(4266));
    layer4_outputs(9447) <= layer3_outputs(606);
    layer4_outputs(9448) <= not(layer3_outputs(1261));
    layer4_outputs(9449) <= layer3_outputs(389);
    layer4_outputs(9450) <= (layer3_outputs(8871)) xor (layer3_outputs(2234));
    layer4_outputs(9451) <= not((layer3_outputs(175)) and (layer3_outputs(5297)));
    layer4_outputs(9452) <= (layer3_outputs(900)) xor (layer3_outputs(1933));
    layer4_outputs(9453) <= (layer3_outputs(3333)) or (layer3_outputs(5643));
    layer4_outputs(9454) <= not(layer3_outputs(8045));
    layer4_outputs(9455) <= layer3_outputs(6931);
    layer4_outputs(9456) <= not(layer3_outputs(7937));
    layer4_outputs(9457) <= layer3_outputs(8187);
    layer4_outputs(9458) <= not(layer3_outputs(9893));
    layer4_outputs(9459) <= (layer3_outputs(3128)) xor (layer3_outputs(999));
    layer4_outputs(9460) <= not((layer3_outputs(6819)) or (layer3_outputs(4875)));
    layer4_outputs(9461) <= not(layer3_outputs(7303));
    layer4_outputs(9462) <= layer3_outputs(1556);
    layer4_outputs(9463) <= not(layer3_outputs(8427));
    layer4_outputs(9464) <= (layer3_outputs(3324)) xor (layer3_outputs(6803));
    layer4_outputs(9465) <= layer3_outputs(748);
    layer4_outputs(9466) <= not((layer3_outputs(2882)) or (layer3_outputs(6839)));
    layer4_outputs(9467) <= not(layer3_outputs(2528));
    layer4_outputs(9468) <= (layer3_outputs(555)) xor (layer3_outputs(5159));
    layer4_outputs(9469) <= (layer3_outputs(2249)) and not (layer3_outputs(8242));
    layer4_outputs(9470) <= (layer3_outputs(2706)) and not (layer3_outputs(7304));
    layer4_outputs(9471) <= not(layer3_outputs(10230));
    layer4_outputs(9472) <= not(layer3_outputs(5297));
    layer4_outputs(9473) <= not((layer3_outputs(7534)) xor (layer3_outputs(5245)));
    layer4_outputs(9474) <= not((layer3_outputs(4672)) or (layer3_outputs(4038)));
    layer4_outputs(9475) <= (layer3_outputs(2943)) and (layer3_outputs(7903));
    layer4_outputs(9476) <= '0';
    layer4_outputs(9477) <= (layer3_outputs(5136)) xor (layer3_outputs(7887));
    layer4_outputs(9478) <= layer3_outputs(1454);
    layer4_outputs(9479) <= (layer3_outputs(2829)) and not (layer3_outputs(7907));
    layer4_outputs(9480) <= not(layer3_outputs(9409));
    layer4_outputs(9481) <= layer3_outputs(3456);
    layer4_outputs(9482) <= '0';
    layer4_outputs(9483) <= not(layer3_outputs(5339));
    layer4_outputs(9484) <= not(layer3_outputs(1736)) or (layer3_outputs(595));
    layer4_outputs(9485) <= not(layer3_outputs(7970));
    layer4_outputs(9486) <= not(layer3_outputs(5068));
    layer4_outputs(9487) <= layer3_outputs(8496);
    layer4_outputs(9488) <= '0';
    layer4_outputs(9489) <= layer3_outputs(4066);
    layer4_outputs(9490) <= layer3_outputs(4363);
    layer4_outputs(9491) <= not(layer3_outputs(2716));
    layer4_outputs(9492) <= not(layer3_outputs(6040));
    layer4_outputs(9493) <= (layer3_outputs(7596)) and not (layer3_outputs(7654));
    layer4_outputs(9494) <= layer3_outputs(790);
    layer4_outputs(9495) <= not(layer3_outputs(899));
    layer4_outputs(9496) <= layer3_outputs(6859);
    layer4_outputs(9497) <= layer3_outputs(7997);
    layer4_outputs(9498) <= layer3_outputs(761);
    layer4_outputs(9499) <= not((layer3_outputs(10103)) or (layer3_outputs(8001)));
    layer4_outputs(9500) <= not((layer3_outputs(2385)) xor (layer3_outputs(7346)));
    layer4_outputs(9501) <= not((layer3_outputs(8298)) and (layer3_outputs(4675)));
    layer4_outputs(9502) <= not((layer3_outputs(1748)) and (layer3_outputs(8159)));
    layer4_outputs(9503) <= not((layer3_outputs(3839)) xor (layer3_outputs(4197)));
    layer4_outputs(9504) <= layer3_outputs(3158);
    layer4_outputs(9505) <= not(layer3_outputs(7466));
    layer4_outputs(9506) <= layer3_outputs(6836);
    layer4_outputs(9507) <= not(layer3_outputs(3484)) or (layer3_outputs(9846));
    layer4_outputs(9508) <= not((layer3_outputs(2799)) and (layer3_outputs(1948)));
    layer4_outputs(9509) <= layer3_outputs(2558);
    layer4_outputs(9510) <= not((layer3_outputs(3570)) xor (layer3_outputs(7756)));
    layer4_outputs(9511) <= not(layer3_outputs(1815)) or (layer3_outputs(6161));
    layer4_outputs(9512) <= (layer3_outputs(337)) and not (layer3_outputs(4310));
    layer4_outputs(9513) <= (layer3_outputs(2222)) and not (layer3_outputs(4239));
    layer4_outputs(9514) <= not(layer3_outputs(6355));
    layer4_outputs(9515) <= layer3_outputs(3205);
    layer4_outputs(9516) <= layer3_outputs(1452);
    layer4_outputs(9517) <= (layer3_outputs(6644)) and (layer3_outputs(2924));
    layer4_outputs(9518) <= layer3_outputs(238);
    layer4_outputs(9519) <= not(layer3_outputs(7136));
    layer4_outputs(9520) <= not(layer3_outputs(729));
    layer4_outputs(9521) <= not(layer3_outputs(670)) or (layer3_outputs(9415));
    layer4_outputs(9522) <= (layer3_outputs(8822)) and not (layer3_outputs(7652));
    layer4_outputs(9523) <= not(layer3_outputs(5952));
    layer4_outputs(9524) <= not(layer3_outputs(9763));
    layer4_outputs(9525) <= layer3_outputs(2762);
    layer4_outputs(9526) <= (layer3_outputs(5017)) xor (layer3_outputs(3029));
    layer4_outputs(9527) <= not((layer3_outputs(4355)) xor (layer3_outputs(10195)));
    layer4_outputs(9528) <= (layer3_outputs(3788)) and not (layer3_outputs(5555));
    layer4_outputs(9529) <= not((layer3_outputs(77)) xor (layer3_outputs(5169)));
    layer4_outputs(9530) <= (layer3_outputs(5151)) xor (layer3_outputs(6788));
    layer4_outputs(9531) <= not(layer3_outputs(4132)) or (layer3_outputs(1093));
    layer4_outputs(9532) <= not(layer3_outputs(8673));
    layer4_outputs(9533) <= (layer3_outputs(10062)) xor (layer3_outputs(2604));
    layer4_outputs(9534) <= (layer3_outputs(227)) xor (layer3_outputs(6071));
    layer4_outputs(9535) <= (layer3_outputs(6727)) and not (layer3_outputs(8751));
    layer4_outputs(9536) <= not(layer3_outputs(6446));
    layer4_outputs(9537) <= not(layer3_outputs(3660));
    layer4_outputs(9538) <= not(layer3_outputs(4617));
    layer4_outputs(9539) <= not(layer3_outputs(1018)) or (layer3_outputs(7061));
    layer4_outputs(9540) <= not(layer3_outputs(9393));
    layer4_outputs(9541) <= not(layer3_outputs(9134));
    layer4_outputs(9542) <= '1';
    layer4_outputs(9543) <= not((layer3_outputs(7985)) xor (layer3_outputs(7368)));
    layer4_outputs(9544) <= (layer3_outputs(1460)) and not (layer3_outputs(1053));
    layer4_outputs(9545) <= (layer3_outputs(10069)) and not (layer3_outputs(308));
    layer4_outputs(9546) <= not(layer3_outputs(295));
    layer4_outputs(9547) <= not((layer3_outputs(8094)) xor (layer3_outputs(1594)));
    layer4_outputs(9548) <= layer3_outputs(1033);
    layer4_outputs(9549) <= not(layer3_outputs(10054));
    layer4_outputs(9550) <= layer3_outputs(6325);
    layer4_outputs(9551) <= not(layer3_outputs(5875));
    layer4_outputs(9552) <= not((layer3_outputs(6342)) or (layer3_outputs(8912)));
    layer4_outputs(9553) <= (layer3_outputs(6327)) and not (layer3_outputs(2727));
    layer4_outputs(9554) <= layer3_outputs(380);
    layer4_outputs(9555) <= not(layer3_outputs(4194));
    layer4_outputs(9556) <= not(layer3_outputs(8016));
    layer4_outputs(9557) <= layer3_outputs(7002);
    layer4_outputs(9558) <= not((layer3_outputs(433)) or (layer3_outputs(6701)));
    layer4_outputs(9559) <= (layer3_outputs(6454)) or (layer3_outputs(8024));
    layer4_outputs(9560) <= not(layer3_outputs(7981)) or (layer3_outputs(572));
    layer4_outputs(9561) <= not((layer3_outputs(3465)) or (layer3_outputs(9366)));
    layer4_outputs(9562) <= not((layer3_outputs(4657)) or (layer3_outputs(7066)));
    layer4_outputs(9563) <= not((layer3_outputs(5751)) and (layer3_outputs(8999)));
    layer4_outputs(9564) <= layer3_outputs(9094);
    layer4_outputs(9565) <= not(layer3_outputs(5711));
    layer4_outputs(9566) <= layer3_outputs(882);
    layer4_outputs(9567) <= layer3_outputs(6952);
    layer4_outputs(9568) <= layer3_outputs(7225);
    layer4_outputs(9569) <= not(layer3_outputs(5506)) or (layer3_outputs(4332));
    layer4_outputs(9570) <= layer3_outputs(7488);
    layer4_outputs(9571) <= (layer3_outputs(2758)) and not (layer3_outputs(3369));
    layer4_outputs(9572) <= not(layer3_outputs(1750));
    layer4_outputs(9573) <= layer3_outputs(8542);
    layer4_outputs(9574) <= (layer3_outputs(2618)) xor (layer3_outputs(7342));
    layer4_outputs(9575) <= not((layer3_outputs(7695)) xor (layer3_outputs(9284)));
    layer4_outputs(9576) <= layer3_outputs(10080);
    layer4_outputs(9577) <= not(layer3_outputs(5));
    layer4_outputs(9578) <= not((layer3_outputs(2626)) xor (layer3_outputs(7512)));
    layer4_outputs(9579) <= (layer3_outputs(3328)) xor (layer3_outputs(4248));
    layer4_outputs(9580) <= (layer3_outputs(837)) or (layer3_outputs(8446));
    layer4_outputs(9581) <= (layer3_outputs(3164)) xor (layer3_outputs(9120));
    layer4_outputs(9582) <= layer3_outputs(4130);
    layer4_outputs(9583) <= layer3_outputs(7474);
    layer4_outputs(9584) <= layer3_outputs(3228);
    layer4_outputs(9585) <= not(layer3_outputs(5816)) or (layer3_outputs(2817));
    layer4_outputs(9586) <= not(layer3_outputs(1024));
    layer4_outputs(9587) <= not(layer3_outputs(5173));
    layer4_outputs(9588) <= not(layer3_outputs(7808));
    layer4_outputs(9589) <= not(layer3_outputs(1500));
    layer4_outputs(9590) <= (layer3_outputs(5732)) and (layer3_outputs(9636));
    layer4_outputs(9591) <= layer3_outputs(8665);
    layer4_outputs(9592) <= not((layer3_outputs(7003)) and (layer3_outputs(7962)));
    layer4_outputs(9593) <= (layer3_outputs(9781)) and (layer3_outputs(7089));
    layer4_outputs(9594) <= not(layer3_outputs(7880)) or (layer3_outputs(6724));
    layer4_outputs(9595) <= not(layer3_outputs(3537));
    layer4_outputs(9596) <= layer3_outputs(1964);
    layer4_outputs(9597) <= layer3_outputs(2160);
    layer4_outputs(9598) <= layer3_outputs(3898);
    layer4_outputs(9599) <= layer3_outputs(3093);
    layer4_outputs(9600) <= layer3_outputs(10072);
    layer4_outputs(9601) <= (layer3_outputs(1269)) and (layer3_outputs(1988));
    layer4_outputs(9602) <= not((layer3_outputs(19)) or (layer3_outputs(2396)));
    layer4_outputs(9603) <= (layer3_outputs(9862)) or (layer3_outputs(9790));
    layer4_outputs(9604) <= not(layer3_outputs(8454));
    layer4_outputs(9605) <= not((layer3_outputs(2494)) and (layer3_outputs(8346)));
    layer4_outputs(9606) <= not(layer3_outputs(4939)) or (layer3_outputs(10069));
    layer4_outputs(9607) <= not(layer3_outputs(724)) or (layer3_outputs(6996));
    layer4_outputs(9608) <= not(layer3_outputs(10066));
    layer4_outputs(9609) <= '0';
    layer4_outputs(9610) <= layer3_outputs(4768);
    layer4_outputs(9611) <= not(layer3_outputs(9793));
    layer4_outputs(9612) <= not(layer3_outputs(8898));
    layer4_outputs(9613) <= layer3_outputs(9734);
    layer4_outputs(9614) <= not((layer3_outputs(9070)) xor (layer3_outputs(8982)));
    layer4_outputs(9615) <= layer3_outputs(4785);
    layer4_outputs(9616) <= layer3_outputs(2367);
    layer4_outputs(9617) <= not(layer3_outputs(7578)) or (layer3_outputs(6859));
    layer4_outputs(9618) <= not(layer3_outputs(3201));
    layer4_outputs(9619) <= not(layer3_outputs(8993));
    layer4_outputs(9620) <= not((layer3_outputs(2246)) and (layer3_outputs(8609)));
    layer4_outputs(9621) <= (layer3_outputs(204)) xor (layer3_outputs(8262));
    layer4_outputs(9622) <= not(layer3_outputs(1062));
    layer4_outputs(9623) <= layer3_outputs(797);
    layer4_outputs(9624) <= not(layer3_outputs(5059));
    layer4_outputs(9625) <= not(layer3_outputs(708)) or (layer3_outputs(9166));
    layer4_outputs(9626) <= (layer3_outputs(272)) xor (layer3_outputs(5908));
    layer4_outputs(9627) <= layer3_outputs(3877);
    layer4_outputs(9628) <= not(layer3_outputs(3202));
    layer4_outputs(9629) <= not((layer3_outputs(1507)) xor (layer3_outputs(5021)));
    layer4_outputs(9630) <= not(layer3_outputs(1952));
    layer4_outputs(9631) <= not(layer3_outputs(4555));
    layer4_outputs(9632) <= not(layer3_outputs(9199)) or (layer3_outputs(6202));
    layer4_outputs(9633) <= not((layer3_outputs(4198)) xor (layer3_outputs(8463)));
    layer4_outputs(9634) <= not(layer3_outputs(3623));
    layer4_outputs(9635) <= not((layer3_outputs(8878)) or (layer3_outputs(6874)));
    layer4_outputs(9636) <= layer3_outputs(9665);
    layer4_outputs(9637) <= layer3_outputs(8915);
    layer4_outputs(9638) <= (layer3_outputs(9835)) and not (layer3_outputs(4427));
    layer4_outputs(9639) <= layer3_outputs(1241);
    layer4_outputs(9640) <= layer3_outputs(5593);
    layer4_outputs(9641) <= (layer3_outputs(5728)) and not (layer3_outputs(3782));
    layer4_outputs(9642) <= not((layer3_outputs(3339)) xor (layer3_outputs(9977)));
    layer4_outputs(9643) <= not(layer3_outputs(2674));
    layer4_outputs(9644) <= (layer3_outputs(9695)) xor (layer3_outputs(6582));
    layer4_outputs(9645) <= '0';
    layer4_outputs(9646) <= layer3_outputs(4092);
    layer4_outputs(9647) <= not((layer3_outputs(2069)) and (layer3_outputs(5188)));
    layer4_outputs(9648) <= not((layer3_outputs(3794)) and (layer3_outputs(4437)));
    layer4_outputs(9649) <= not(layer3_outputs(5039));
    layer4_outputs(9650) <= not((layer3_outputs(9265)) xor (layer3_outputs(6212)));
    layer4_outputs(9651) <= not(layer3_outputs(6717));
    layer4_outputs(9652) <= layer3_outputs(1047);
    layer4_outputs(9653) <= (layer3_outputs(2271)) xor (layer3_outputs(3712));
    layer4_outputs(9654) <= not(layer3_outputs(9960));
    layer4_outputs(9655) <= not((layer3_outputs(3955)) xor (layer3_outputs(9015)));
    layer4_outputs(9656) <= not(layer3_outputs(4447));
    layer4_outputs(9657) <= (layer3_outputs(861)) xor (layer3_outputs(6818));
    layer4_outputs(9658) <= layer3_outputs(6000);
    layer4_outputs(9659) <= layer3_outputs(673);
    layer4_outputs(9660) <= not((layer3_outputs(8287)) and (layer3_outputs(1226)));
    layer4_outputs(9661) <= layer3_outputs(6090);
    layer4_outputs(9662) <= not(layer3_outputs(784));
    layer4_outputs(9663) <= (layer3_outputs(4749)) xor (layer3_outputs(3884));
    layer4_outputs(9664) <= not(layer3_outputs(8622));
    layer4_outputs(9665) <= layer3_outputs(5894);
    layer4_outputs(9666) <= not(layer3_outputs(2725));
    layer4_outputs(9667) <= not((layer3_outputs(8521)) and (layer3_outputs(3325)));
    layer4_outputs(9668) <= not((layer3_outputs(3338)) and (layer3_outputs(3320)));
    layer4_outputs(9669) <= not(layer3_outputs(7913));
    layer4_outputs(9670) <= (layer3_outputs(1444)) xor (layer3_outputs(2526));
    layer4_outputs(9671) <= layer3_outputs(6714);
    layer4_outputs(9672) <= layer3_outputs(3584);
    layer4_outputs(9673) <= layer3_outputs(6094);
    layer4_outputs(9674) <= layer3_outputs(4656);
    layer4_outputs(9675) <= (layer3_outputs(457)) xor (layer3_outputs(5752));
    layer4_outputs(9676) <= not((layer3_outputs(10065)) and (layer3_outputs(2730)));
    layer4_outputs(9677) <= not(layer3_outputs(5600)) or (layer3_outputs(10058));
    layer4_outputs(9678) <= (layer3_outputs(8221)) xor (layer3_outputs(7459));
    layer4_outputs(9679) <= layer3_outputs(2044);
    layer4_outputs(9680) <= not((layer3_outputs(5943)) or (layer3_outputs(9407)));
    layer4_outputs(9681) <= layer3_outputs(6813);
    layer4_outputs(9682) <= not(layer3_outputs(6983)) or (layer3_outputs(9468));
    layer4_outputs(9683) <= not(layer3_outputs(5779));
    layer4_outputs(9684) <= (layer3_outputs(1005)) xor (layer3_outputs(6060));
    layer4_outputs(9685) <= (layer3_outputs(72)) and not (layer3_outputs(7514));
    layer4_outputs(9686) <= layer3_outputs(6322);
    layer4_outputs(9687) <= '1';
    layer4_outputs(9688) <= not(layer3_outputs(7464));
    layer4_outputs(9689) <= not(layer3_outputs(754));
    layer4_outputs(9690) <= (layer3_outputs(6726)) xor (layer3_outputs(3076));
    layer4_outputs(9691) <= (layer3_outputs(10155)) xor (layer3_outputs(2273));
    layer4_outputs(9692) <= (layer3_outputs(4236)) xor (layer3_outputs(6388));
    layer4_outputs(9693) <= layer3_outputs(7649);
    layer4_outputs(9694) <= (layer3_outputs(1283)) and not (layer3_outputs(5090));
    layer4_outputs(9695) <= layer3_outputs(9377);
    layer4_outputs(9696) <= (layer3_outputs(7345)) xor (layer3_outputs(625));
    layer4_outputs(9697) <= (layer3_outputs(1778)) and (layer3_outputs(5601));
    layer4_outputs(9698) <= not(layer3_outputs(1461));
    layer4_outputs(9699) <= not((layer3_outputs(329)) and (layer3_outputs(3493)));
    layer4_outputs(9700) <= not(layer3_outputs(5582));
    layer4_outputs(9701) <= layer3_outputs(112);
    layer4_outputs(9702) <= (layer3_outputs(8253)) and (layer3_outputs(7516));
    layer4_outputs(9703) <= (layer3_outputs(523)) and not (layer3_outputs(5813));
    layer4_outputs(9704) <= (layer3_outputs(6482)) xor (layer3_outputs(7268));
    layer4_outputs(9705) <= not((layer3_outputs(4713)) xor (layer3_outputs(2697)));
    layer4_outputs(9706) <= not(layer3_outputs(1925));
    layer4_outputs(9707) <= not(layer3_outputs(9306)) or (layer3_outputs(6051));
    layer4_outputs(9708) <= (layer3_outputs(366)) or (layer3_outputs(2175));
    layer4_outputs(9709) <= not(layer3_outputs(4744));
    layer4_outputs(9710) <= not(layer3_outputs(9898));
    layer4_outputs(9711) <= not((layer3_outputs(10040)) xor (layer3_outputs(3426)));
    layer4_outputs(9712) <= not((layer3_outputs(8863)) and (layer3_outputs(3694)));
    layer4_outputs(9713) <= (layer3_outputs(533)) and not (layer3_outputs(1242));
    layer4_outputs(9714) <= not((layer3_outputs(7895)) xor (layer3_outputs(8194)));
    layer4_outputs(9715) <= (layer3_outputs(4519)) or (layer3_outputs(7737));
    layer4_outputs(9716) <= not(layer3_outputs(9842));
    layer4_outputs(9717) <= layer3_outputs(7478);
    layer4_outputs(9718) <= layer3_outputs(5562);
    layer4_outputs(9719) <= not(layer3_outputs(1323));
    layer4_outputs(9720) <= not((layer3_outputs(4658)) xor (layer3_outputs(1800)));
    layer4_outputs(9721) <= (layer3_outputs(385)) and not (layer3_outputs(3843));
    layer4_outputs(9722) <= (layer3_outputs(5440)) xor (layer3_outputs(3027));
    layer4_outputs(9723) <= layer3_outputs(7048);
    layer4_outputs(9724) <= not((layer3_outputs(249)) or (layer3_outputs(1141)));
    layer4_outputs(9725) <= (layer3_outputs(4268)) and (layer3_outputs(8804));
    layer4_outputs(9726) <= layer3_outputs(658);
    layer4_outputs(9727) <= not(layer3_outputs(8809));
    layer4_outputs(9728) <= layer3_outputs(1313);
    layer4_outputs(9729) <= layer3_outputs(4471);
    layer4_outputs(9730) <= not(layer3_outputs(649));
    layer4_outputs(9731) <= layer3_outputs(1234);
    layer4_outputs(9732) <= not(layer3_outputs(6690));
    layer4_outputs(9733) <= not((layer3_outputs(7926)) xor (layer3_outputs(7618)));
    layer4_outputs(9734) <= not((layer3_outputs(8301)) xor (layer3_outputs(5156)));
    layer4_outputs(9735) <= layer3_outputs(8084);
    layer4_outputs(9736) <= layer3_outputs(2600);
    layer4_outputs(9737) <= layer3_outputs(8811);
    layer4_outputs(9738) <= not(layer3_outputs(8927));
    layer4_outputs(9739) <= not((layer3_outputs(9975)) or (layer3_outputs(4761)));
    layer4_outputs(9740) <= layer3_outputs(1461);
    layer4_outputs(9741) <= not(layer3_outputs(6741));
    layer4_outputs(9742) <= (layer3_outputs(5817)) and not (layer3_outputs(91));
    layer4_outputs(9743) <= not(layer3_outputs(6034));
    layer4_outputs(9744) <= (layer3_outputs(10157)) and (layer3_outputs(3396));
    layer4_outputs(9745) <= layer3_outputs(530);
    layer4_outputs(9746) <= (layer3_outputs(924)) xor (layer3_outputs(7669));
    layer4_outputs(9747) <= not(layer3_outputs(3212));
    layer4_outputs(9748) <= layer3_outputs(8378);
    layer4_outputs(9749) <= not(layer3_outputs(8309)) or (layer3_outputs(4419));
    layer4_outputs(9750) <= not(layer3_outputs(5202));
    layer4_outputs(9751) <= (layer3_outputs(7219)) or (layer3_outputs(5509));
    layer4_outputs(9752) <= not(layer3_outputs(4889));
    layer4_outputs(9753) <= not(layer3_outputs(6190)) or (layer3_outputs(10136));
    layer4_outputs(9754) <= (layer3_outputs(6232)) and not (layer3_outputs(9346));
    layer4_outputs(9755) <= not((layer3_outputs(1954)) xor (layer3_outputs(6796)));
    layer4_outputs(9756) <= layer3_outputs(5523);
    layer4_outputs(9757) <= layer3_outputs(6766);
    layer4_outputs(9758) <= not((layer3_outputs(4293)) or (layer3_outputs(9037)));
    layer4_outputs(9759) <= (layer3_outputs(4460)) xor (layer3_outputs(10031));
    layer4_outputs(9760) <= not(layer3_outputs(4930));
    layer4_outputs(9761) <= layer3_outputs(1560);
    layer4_outputs(9762) <= (layer3_outputs(1235)) xor (layer3_outputs(7222));
    layer4_outputs(9763) <= layer3_outputs(7281);
    layer4_outputs(9764) <= (layer3_outputs(4888)) xor (layer3_outputs(2489));
    layer4_outputs(9765) <= (layer3_outputs(4959)) and not (layer3_outputs(4542));
    layer4_outputs(9766) <= layer3_outputs(1102);
    layer4_outputs(9767) <= not(layer3_outputs(8839));
    layer4_outputs(9768) <= layer3_outputs(2255);
    layer4_outputs(9769) <= (layer3_outputs(5028)) xor (layer3_outputs(2327));
    layer4_outputs(9770) <= not(layer3_outputs(1594));
    layer4_outputs(9771) <= (layer3_outputs(867)) and (layer3_outputs(984));
    layer4_outputs(9772) <= '0';
    layer4_outputs(9773) <= not((layer3_outputs(8569)) xor (layer3_outputs(6025)));
    layer4_outputs(9774) <= layer3_outputs(6010);
    layer4_outputs(9775) <= (layer3_outputs(9000)) xor (layer3_outputs(5230));
    layer4_outputs(9776) <= not(layer3_outputs(6713));
    layer4_outputs(9777) <= layer3_outputs(7688);
    layer4_outputs(9778) <= not(layer3_outputs(7203)) or (layer3_outputs(9100));
    layer4_outputs(9779) <= not((layer3_outputs(9417)) xor (layer3_outputs(7841)));
    layer4_outputs(9780) <= (layer3_outputs(10105)) and not (layer3_outputs(7780));
    layer4_outputs(9781) <= layer3_outputs(3392);
    layer4_outputs(9782) <= not(layer3_outputs(9828));
    layer4_outputs(9783) <= not((layer3_outputs(8905)) xor (layer3_outputs(43)));
    layer4_outputs(9784) <= layer3_outputs(9321);
    layer4_outputs(9785) <= layer3_outputs(6260);
    layer4_outputs(9786) <= layer3_outputs(5923);
    layer4_outputs(9787) <= not(layer3_outputs(5995));
    layer4_outputs(9788) <= layer3_outputs(1365);
    layer4_outputs(9789) <= not(layer3_outputs(5909));
    layer4_outputs(9790) <= not(layer3_outputs(7390)) or (layer3_outputs(9810));
    layer4_outputs(9791) <= not(layer3_outputs(1549)) or (layer3_outputs(1371));
    layer4_outputs(9792) <= not((layer3_outputs(9694)) or (layer3_outputs(6906)));
    layer4_outputs(9793) <= (layer3_outputs(4483)) and (layer3_outputs(1791));
    layer4_outputs(9794) <= layer3_outputs(3841);
    layer4_outputs(9795) <= layer3_outputs(1827);
    layer4_outputs(9796) <= layer3_outputs(8216);
    layer4_outputs(9797) <= not(layer3_outputs(121)) or (layer3_outputs(1421));
    layer4_outputs(9798) <= layer3_outputs(10122);
    layer4_outputs(9799) <= layer3_outputs(9599);
    layer4_outputs(9800) <= layer3_outputs(3568);
    layer4_outputs(9801) <= (layer3_outputs(6201)) xor (layer3_outputs(6330));
    layer4_outputs(9802) <= (layer3_outputs(4872)) and (layer3_outputs(7414));
    layer4_outputs(9803) <= layer3_outputs(5636);
    layer4_outputs(9804) <= layer3_outputs(9553);
    layer4_outputs(9805) <= not(layer3_outputs(9662));
    layer4_outputs(9806) <= layer3_outputs(3968);
    layer4_outputs(9807) <= layer3_outputs(2118);
    layer4_outputs(9808) <= not((layer3_outputs(8030)) or (layer3_outputs(5544)));
    layer4_outputs(9809) <= (layer3_outputs(8375)) and not (layer3_outputs(8061));
    layer4_outputs(9810) <= layer3_outputs(155);
    layer4_outputs(9811) <= layer3_outputs(990);
    layer4_outputs(9812) <= not((layer3_outputs(5000)) or (layer3_outputs(4304)));
    layer4_outputs(9813) <= layer3_outputs(8468);
    layer4_outputs(9814) <= layer3_outputs(3219);
    layer4_outputs(9815) <= not(layer3_outputs(7772));
    layer4_outputs(9816) <= layer3_outputs(1407);
    layer4_outputs(9817) <= not((layer3_outputs(7167)) xor (layer3_outputs(8991)));
    layer4_outputs(9818) <= not(layer3_outputs(6753));
    layer4_outputs(9819) <= layer3_outputs(5589);
    layer4_outputs(9820) <= not(layer3_outputs(4931));
    layer4_outputs(9821) <= (layer3_outputs(9175)) or (layer3_outputs(8370));
    layer4_outputs(9822) <= layer3_outputs(7805);
    layer4_outputs(9823) <= not((layer3_outputs(8504)) xor (layer3_outputs(4566)));
    layer4_outputs(9824) <= (layer3_outputs(1735)) xor (layer3_outputs(8317));
    layer4_outputs(9825) <= layer3_outputs(8457);
    layer4_outputs(9826) <= not((layer3_outputs(7893)) xor (layer3_outputs(4839)));
    layer4_outputs(9827) <= not(layer3_outputs(5543));
    layer4_outputs(9828) <= not(layer3_outputs(503)) or (layer3_outputs(4389));
    layer4_outputs(9829) <= not(layer3_outputs(7570));
    layer4_outputs(9830) <= not(layer3_outputs(4765));
    layer4_outputs(9831) <= (layer3_outputs(8953)) xor (layer3_outputs(5234));
    layer4_outputs(9832) <= not((layer3_outputs(6280)) and (layer3_outputs(3088)));
    layer4_outputs(9833) <= not(layer3_outputs(7734));
    layer4_outputs(9834) <= (layer3_outputs(7562)) xor (layer3_outputs(2696));
    layer4_outputs(9835) <= (layer3_outputs(5436)) and not (layer3_outputs(8929));
    layer4_outputs(9836) <= not(layer3_outputs(3263)) or (layer3_outputs(3689));
    layer4_outputs(9837) <= not(layer3_outputs(10022)) or (layer3_outputs(4906));
    layer4_outputs(9838) <= (layer3_outputs(8183)) and not (layer3_outputs(4308));
    layer4_outputs(9839) <= not(layer3_outputs(7551));
    layer4_outputs(9840) <= layer3_outputs(5883);
    layer4_outputs(9841) <= layer3_outputs(6307);
    layer4_outputs(9842) <= layer3_outputs(2759);
    layer4_outputs(9843) <= layer3_outputs(8636);
    layer4_outputs(9844) <= not(layer3_outputs(1557));
    layer4_outputs(9845) <= not(layer3_outputs(1728));
    layer4_outputs(9846) <= not(layer3_outputs(1480));
    layer4_outputs(9847) <= layer3_outputs(4773);
    layer4_outputs(9848) <= not(layer3_outputs(2570));
    layer4_outputs(9849) <= (layer3_outputs(2276)) and not (layer3_outputs(9430));
    layer4_outputs(9850) <= not(layer3_outputs(4087));
    layer4_outputs(9851) <= not(layer3_outputs(5496));
    layer4_outputs(9852) <= layer3_outputs(4683);
    layer4_outputs(9853) <= not(layer3_outputs(498));
    layer4_outputs(9854) <= layer3_outputs(1822);
    layer4_outputs(9855) <= not((layer3_outputs(1044)) and (layer3_outputs(7196)));
    layer4_outputs(9856) <= not(layer3_outputs(167));
    layer4_outputs(9857) <= layer3_outputs(1989);
    layer4_outputs(9858) <= layer3_outputs(6040);
    layer4_outputs(9859) <= not(layer3_outputs(8579));
    layer4_outputs(9860) <= layer3_outputs(2297);
    layer4_outputs(9861) <= layer3_outputs(3330);
    layer4_outputs(9862) <= (layer3_outputs(8502)) and (layer3_outputs(4754));
    layer4_outputs(9863) <= layer3_outputs(4484);
    layer4_outputs(9864) <= not((layer3_outputs(1268)) xor (layer3_outputs(6002)));
    layer4_outputs(9865) <= not((layer3_outputs(4447)) or (layer3_outputs(4592)));
    layer4_outputs(9866) <= not(layer3_outputs(3989)) or (layer3_outputs(7727));
    layer4_outputs(9867) <= not(layer3_outputs(8901));
    layer4_outputs(9868) <= layer3_outputs(7089);
    layer4_outputs(9869) <= not((layer3_outputs(5428)) xor (layer3_outputs(3479)));
    layer4_outputs(9870) <= (layer3_outputs(2198)) xor (layer3_outputs(7923));
    layer4_outputs(9871) <= not(layer3_outputs(1400));
    layer4_outputs(9872) <= layer3_outputs(7874);
    layer4_outputs(9873) <= not(layer3_outputs(3469));
    layer4_outputs(9874) <= not((layer3_outputs(1616)) xor (layer3_outputs(3409)));
    layer4_outputs(9875) <= (layer3_outputs(8190)) and not (layer3_outputs(8319));
    layer4_outputs(9876) <= not(layer3_outputs(4232));
    layer4_outputs(9877) <= layer3_outputs(5870);
    layer4_outputs(9878) <= not(layer3_outputs(597)) or (layer3_outputs(787));
    layer4_outputs(9879) <= not(layer3_outputs(4060));
    layer4_outputs(9880) <= layer3_outputs(10007);
    layer4_outputs(9881) <= (layer3_outputs(3342)) and not (layer3_outputs(6081));
    layer4_outputs(9882) <= layer3_outputs(7869);
    layer4_outputs(9883) <= layer3_outputs(291);
    layer4_outputs(9884) <= not((layer3_outputs(6576)) xor (layer3_outputs(693)));
    layer4_outputs(9885) <= (layer3_outputs(4744)) xor (layer3_outputs(2656));
    layer4_outputs(9886) <= not((layer3_outputs(1680)) or (layer3_outputs(1926)));
    layer4_outputs(9887) <= not((layer3_outputs(1614)) or (layer3_outputs(376)));
    layer4_outputs(9888) <= not((layer3_outputs(9035)) or (layer3_outputs(874)));
    layer4_outputs(9889) <= not(layer3_outputs(2168)) or (layer3_outputs(2306));
    layer4_outputs(9890) <= not(layer3_outputs(8267));
    layer4_outputs(9891) <= not(layer3_outputs(4607));
    layer4_outputs(9892) <= not(layer3_outputs(5012)) or (layer3_outputs(2101));
    layer4_outputs(9893) <= layer3_outputs(6782);
    layer4_outputs(9894) <= not((layer3_outputs(8846)) or (layer3_outputs(9072)));
    layer4_outputs(9895) <= not(layer3_outputs(7013));
    layer4_outputs(9896) <= not((layer3_outputs(2989)) xor (layer3_outputs(3317)));
    layer4_outputs(9897) <= not(layer3_outputs(5184));
    layer4_outputs(9898) <= not((layer3_outputs(1910)) xor (layer3_outputs(5786)));
    layer4_outputs(9899) <= not(layer3_outputs(5162));
    layer4_outputs(9900) <= layer3_outputs(10218);
    layer4_outputs(9901) <= not(layer3_outputs(10164));
    layer4_outputs(9902) <= layer3_outputs(6560);
    layer4_outputs(9903) <= layer3_outputs(2713);
    layer4_outputs(9904) <= not((layer3_outputs(5124)) xor (layer3_outputs(4458)));
    layer4_outputs(9905) <= (layer3_outputs(7393)) or (layer3_outputs(5536));
    layer4_outputs(9906) <= '0';
    layer4_outputs(9907) <= layer3_outputs(348);
    layer4_outputs(9908) <= (layer3_outputs(3609)) and not (layer3_outputs(7152));
    layer4_outputs(9909) <= not(layer3_outputs(8148));
    layer4_outputs(9910) <= not(layer3_outputs(4960));
    layer4_outputs(9911) <= not((layer3_outputs(2593)) and (layer3_outputs(7388)));
    layer4_outputs(9912) <= layer3_outputs(3783);
    layer4_outputs(9913) <= not(layer3_outputs(6608));
    layer4_outputs(9914) <= layer3_outputs(3723);
    layer4_outputs(9915) <= (layer3_outputs(9825)) and (layer3_outputs(3922));
    layer4_outputs(9916) <= not(layer3_outputs(8044));
    layer4_outputs(9917) <= (layer3_outputs(5926)) xor (layer3_outputs(9545));
    layer4_outputs(9918) <= layer3_outputs(8636);
    layer4_outputs(9919) <= layer3_outputs(9779);
    layer4_outputs(9920) <= not(layer3_outputs(604));
    layer4_outputs(9921) <= layer3_outputs(8610);
    layer4_outputs(9922) <= layer3_outputs(2311);
    layer4_outputs(9923) <= layer3_outputs(5305);
    layer4_outputs(9924) <= not((layer3_outputs(4361)) xor (layer3_outputs(3734)));
    layer4_outputs(9925) <= (layer3_outputs(4645)) xor (layer3_outputs(6715));
    layer4_outputs(9926) <= not(layer3_outputs(9963));
    layer4_outputs(9927) <= not(layer3_outputs(10034));
    layer4_outputs(9928) <= not(layer3_outputs(93));
    layer4_outputs(9929) <= (layer3_outputs(9019)) xor (layer3_outputs(146));
    layer4_outputs(9930) <= layer3_outputs(1035);
    layer4_outputs(9931) <= not((layer3_outputs(5540)) or (layer3_outputs(3132)));
    layer4_outputs(9932) <= not(layer3_outputs(8880));
    layer4_outputs(9933) <= layer3_outputs(8959);
    layer4_outputs(9934) <= layer3_outputs(2312);
    layer4_outputs(9935) <= not(layer3_outputs(5580));
    layer4_outputs(9936) <= (layer3_outputs(1763)) xor (layer3_outputs(2028));
    layer4_outputs(9937) <= (layer3_outputs(5149)) xor (layer3_outputs(1698));
    layer4_outputs(9938) <= not(layer3_outputs(8503));
    layer4_outputs(9939) <= not(layer3_outputs(5569));
    layer4_outputs(9940) <= not((layer3_outputs(1363)) xor (layer3_outputs(1725)));
    layer4_outputs(9941) <= layer3_outputs(4651);
    layer4_outputs(9942) <= not(layer3_outputs(8447));
    layer4_outputs(9943) <= not((layer3_outputs(1505)) xor (layer3_outputs(1028)));
    layer4_outputs(9944) <= not(layer3_outputs(2853)) or (layer3_outputs(5519));
    layer4_outputs(9945) <= not((layer3_outputs(9858)) xor (layer3_outputs(5531)));
    layer4_outputs(9946) <= '0';
    layer4_outputs(9947) <= layer3_outputs(5278);
    layer4_outputs(9948) <= not(layer3_outputs(4842));
    layer4_outputs(9949) <= (layer3_outputs(5407)) xor (layer3_outputs(9696));
    layer4_outputs(9950) <= layer3_outputs(4968);
    layer4_outputs(9951) <= not(layer3_outputs(6781)) or (layer3_outputs(6101));
    layer4_outputs(9952) <= not((layer3_outputs(8900)) xor (layer3_outputs(6311)));
    layer4_outputs(9953) <= not(layer3_outputs(4017));
    layer4_outputs(9954) <= not(layer3_outputs(3081));
    layer4_outputs(9955) <= not((layer3_outputs(6461)) and (layer3_outputs(7477)));
    layer4_outputs(9956) <= not(layer3_outputs(3666)) or (layer3_outputs(6927));
    layer4_outputs(9957) <= layer3_outputs(7366);
    layer4_outputs(9958) <= not(layer3_outputs(1731)) or (layer3_outputs(2531));
    layer4_outputs(9959) <= (layer3_outputs(5137)) xor (layer3_outputs(4896));
    layer4_outputs(9960) <= layer3_outputs(9358);
    layer4_outputs(9961) <= not((layer3_outputs(8983)) or (layer3_outputs(1778)));
    layer4_outputs(9962) <= (layer3_outputs(2875)) and not (layer3_outputs(5131));
    layer4_outputs(9963) <= not((layer3_outputs(757)) or (layer3_outputs(5546)));
    layer4_outputs(9964) <= layer3_outputs(3732);
    layer4_outputs(9965) <= (layer3_outputs(6987)) or (layer3_outputs(7356));
    layer4_outputs(9966) <= not(layer3_outputs(300)) or (layer3_outputs(948));
    layer4_outputs(9967) <= not((layer3_outputs(10135)) and (layer3_outputs(2470)));
    layer4_outputs(9968) <= (layer3_outputs(5316)) or (layer3_outputs(8013));
    layer4_outputs(9969) <= (layer3_outputs(1941)) xor (layer3_outputs(1260));
    layer4_outputs(9970) <= '0';
    layer4_outputs(9971) <= layer3_outputs(4453);
    layer4_outputs(9972) <= not(layer3_outputs(5753));
    layer4_outputs(9973) <= not(layer3_outputs(10076));
    layer4_outputs(9974) <= layer3_outputs(8305);
    layer4_outputs(9975) <= not(layer3_outputs(8651));
    layer4_outputs(9976) <= not(layer3_outputs(3026)) or (layer3_outputs(104));
    layer4_outputs(9977) <= layer3_outputs(5576);
    layer4_outputs(9978) <= not(layer3_outputs(2928));
    layer4_outputs(9979) <= not(layer3_outputs(5152));
    layer4_outputs(9980) <= not((layer3_outputs(3043)) and (layer3_outputs(8295)));
    layer4_outputs(9981) <= layer3_outputs(5257);
    layer4_outputs(9982) <= not(layer3_outputs(2941));
    layer4_outputs(9983) <= not(layer3_outputs(3400));
    layer4_outputs(9984) <= (layer3_outputs(8485)) and not (layer3_outputs(4238));
    layer4_outputs(9985) <= (layer3_outputs(8567)) xor (layer3_outputs(9628));
    layer4_outputs(9986) <= not(layer3_outputs(6944));
    layer4_outputs(9987) <= not((layer3_outputs(2223)) xor (layer3_outputs(7735)));
    layer4_outputs(9988) <= (layer3_outputs(7113)) and not (layer3_outputs(3691));
    layer4_outputs(9989) <= layer3_outputs(2830);
    layer4_outputs(9990) <= layer3_outputs(8746);
    layer4_outputs(9991) <= not(layer3_outputs(7518));
    layer4_outputs(9992) <= not((layer3_outputs(4547)) and (layer3_outputs(2051)));
    layer4_outputs(9993) <= not((layer3_outputs(5003)) or (layer3_outputs(7417)));
    layer4_outputs(9994) <= (layer3_outputs(8238)) or (layer3_outputs(3070));
    layer4_outputs(9995) <= not(layer3_outputs(4233));
    layer4_outputs(9996) <= layer3_outputs(8203);
    layer4_outputs(9997) <= not(layer3_outputs(3034));
    layer4_outputs(9998) <= layer3_outputs(4088);
    layer4_outputs(9999) <= layer3_outputs(4145);
    layer4_outputs(10000) <= (layer3_outputs(9995)) and not (layer3_outputs(7463));
    layer4_outputs(10001) <= layer3_outputs(8285);
    layer4_outputs(10002) <= not((layer3_outputs(1741)) xor (layer3_outputs(9333)));
    layer4_outputs(10003) <= not(layer3_outputs(4302));
    layer4_outputs(10004) <= not(layer3_outputs(4111));
    layer4_outputs(10005) <= layer3_outputs(1441);
    layer4_outputs(10006) <= not(layer3_outputs(848)) or (layer3_outputs(7608));
    layer4_outputs(10007) <= layer3_outputs(7115);
    layer4_outputs(10008) <= not(layer3_outputs(8677));
    layer4_outputs(10009) <= layer3_outputs(1212);
    layer4_outputs(10010) <= not(layer3_outputs(10011)) or (layer3_outputs(9043));
    layer4_outputs(10011) <= not(layer3_outputs(2338));
    layer4_outputs(10012) <= (layer3_outputs(4532)) and not (layer3_outputs(9412));
    layer4_outputs(10013) <= layer3_outputs(6149);
    layer4_outputs(10014) <= layer3_outputs(5986);
    layer4_outputs(10015) <= not((layer3_outputs(9013)) xor (layer3_outputs(5432)));
    layer4_outputs(10016) <= layer3_outputs(1257);
    layer4_outputs(10017) <= not(layer3_outputs(933));
    layer4_outputs(10018) <= not((layer3_outputs(953)) xor (layer3_outputs(2182)));
    layer4_outputs(10019) <= not(layer3_outputs(7085)) or (layer3_outputs(959));
    layer4_outputs(10020) <= not((layer3_outputs(7353)) and (layer3_outputs(7197)));
    layer4_outputs(10021) <= layer3_outputs(868);
    layer4_outputs(10022) <= '1';
    layer4_outputs(10023) <= layer3_outputs(3300);
    layer4_outputs(10024) <= (layer3_outputs(6473)) xor (layer3_outputs(3253));
    layer4_outputs(10025) <= not(layer3_outputs(7467));
    layer4_outputs(10026) <= not(layer3_outputs(5656));
    layer4_outputs(10027) <= (layer3_outputs(111)) and not (layer3_outputs(5101));
    layer4_outputs(10028) <= not(layer3_outputs(169));
    layer4_outputs(10029) <= layer3_outputs(142);
    layer4_outputs(10030) <= not(layer3_outputs(6632)) or (layer3_outputs(6286));
    layer4_outputs(10031) <= not(layer3_outputs(569));
    layer4_outputs(10032) <= layer3_outputs(3970);
    layer4_outputs(10033) <= (layer3_outputs(4479)) xor (layer3_outputs(496));
    layer4_outputs(10034) <= layer3_outputs(6622);
    layer4_outputs(10035) <= layer3_outputs(2123);
    layer4_outputs(10036) <= not(layer3_outputs(63));
    layer4_outputs(10037) <= not(layer3_outputs(7399)) or (layer3_outputs(755));
    layer4_outputs(10038) <= (layer3_outputs(8726)) xor (layer3_outputs(4762));
    layer4_outputs(10039) <= (layer3_outputs(3112)) and not (layer3_outputs(305));
    layer4_outputs(10040) <= not(layer3_outputs(6092)) or (layer3_outputs(669));
    layer4_outputs(10041) <= not(layer3_outputs(8603));
    layer4_outputs(10042) <= layer3_outputs(517);
    layer4_outputs(10043) <= not(layer3_outputs(7442));
    layer4_outputs(10044) <= layer3_outputs(5875);
    layer4_outputs(10045) <= not(layer3_outputs(9708));
    layer4_outputs(10046) <= layer3_outputs(8005);
    layer4_outputs(10047) <= layer3_outputs(5250);
    layer4_outputs(10048) <= layer3_outputs(5071);
    layer4_outputs(10049) <= (layer3_outputs(1562)) and (layer3_outputs(9158));
    layer4_outputs(10050) <= not(layer3_outputs(8567)) or (layer3_outputs(1331));
    layer4_outputs(10051) <= layer3_outputs(4287);
    layer4_outputs(10052) <= not((layer3_outputs(5945)) xor (layer3_outputs(3940)));
    layer4_outputs(10053) <= not(layer3_outputs(8357));
    layer4_outputs(10054) <= (layer3_outputs(8421)) xor (layer3_outputs(4000));
    layer4_outputs(10055) <= not(layer3_outputs(9778)) or (layer3_outputs(8207));
    layer4_outputs(10056) <= (layer3_outputs(1979)) and not (layer3_outputs(8020));
    layer4_outputs(10057) <= (layer3_outputs(2155)) or (layer3_outputs(2292));
    layer4_outputs(10058) <= layer3_outputs(10135);
    layer4_outputs(10059) <= not(layer3_outputs(9172));
    layer4_outputs(10060) <= not(layer3_outputs(620)) or (layer3_outputs(8862));
    layer4_outputs(10061) <= not(layer3_outputs(5846));
    layer4_outputs(10062) <= not(layer3_outputs(4981));
    layer4_outputs(10063) <= not(layer3_outputs(9667));
    layer4_outputs(10064) <= layer3_outputs(939);
    layer4_outputs(10065) <= not((layer3_outputs(6326)) and (layer3_outputs(8835)));
    layer4_outputs(10066) <= not(layer3_outputs(8512));
    layer4_outputs(10067) <= not((layer3_outputs(4703)) xor (layer3_outputs(7791)));
    layer4_outputs(10068) <= (layer3_outputs(3242)) and not (layer3_outputs(5722));
    layer4_outputs(10069) <= not(layer3_outputs(4259));
    layer4_outputs(10070) <= layer3_outputs(3264);
    layer4_outputs(10071) <= layer3_outputs(1600);
    layer4_outputs(10072) <= (layer3_outputs(4049)) and not (layer3_outputs(8577));
    layer4_outputs(10073) <= layer3_outputs(2657);
    layer4_outputs(10074) <= not((layer3_outputs(9614)) xor (layer3_outputs(6868)));
    layer4_outputs(10075) <= layer3_outputs(7533);
    layer4_outputs(10076) <= layer3_outputs(5444);
    layer4_outputs(10077) <= layer3_outputs(6782);
    layer4_outputs(10078) <= not((layer3_outputs(9995)) xor (layer3_outputs(601)));
    layer4_outputs(10079) <= layer3_outputs(4860);
    layer4_outputs(10080) <= (layer3_outputs(8116)) or (layer3_outputs(8130));
    layer4_outputs(10081) <= not(layer3_outputs(2396));
    layer4_outputs(10082) <= layer3_outputs(5055);
    layer4_outputs(10083) <= layer3_outputs(9770);
    layer4_outputs(10084) <= layer3_outputs(9522);
    layer4_outputs(10085) <= not((layer3_outputs(7601)) or (layer3_outputs(3675)));
    layer4_outputs(10086) <= not((layer3_outputs(3399)) xor (layer3_outputs(7124)));
    layer4_outputs(10087) <= layer3_outputs(2740);
    layer4_outputs(10088) <= not(layer3_outputs(1122)) or (layer3_outputs(7472));
    layer4_outputs(10089) <= not((layer3_outputs(1237)) xor (layer3_outputs(10170)));
    layer4_outputs(10090) <= not(layer3_outputs(8613));
    layer4_outputs(10091) <= not(layer3_outputs(9741));
    layer4_outputs(10092) <= not((layer3_outputs(5167)) or (layer3_outputs(4565)));
    layer4_outputs(10093) <= not((layer3_outputs(1219)) and (layer3_outputs(3421)));
    layer4_outputs(10094) <= (layer3_outputs(5368)) xor (layer3_outputs(7237));
    layer4_outputs(10095) <= (layer3_outputs(2712)) xor (layer3_outputs(4954));
    layer4_outputs(10096) <= not(layer3_outputs(7473));
    layer4_outputs(10097) <= not(layer3_outputs(3685));
    layer4_outputs(10098) <= layer3_outputs(1257);
    layer4_outputs(10099) <= (layer3_outputs(6728)) xor (layer3_outputs(2643));
    layer4_outputs(10100) <= not(layer3_outputs(4502));
    layer4_outputs(10101) <= layer3_outputs(8644);
    layer4_outputs(10102) <= not(layer3_outputs(9899));
    layer4_outputs(10103) <= not(layer3_outputs(9691));
    layer4_outputs(10104) <= not((layer3_outputs(916)) or (layer3_outputs(1091)));
    layer4_outputs(10105) <= (layer3_outputs(8003)) and not (layer3_outputs(4405));
    layer4_outputs(10106) <= (layer3_outputs(9700)) or (layer3_outputs(7626));
    layer4_outputs(10107) <= '1';
    layer4_outputs(10108) <= not(layer3_outputs(8710));
    layer4_outputs(10109) <= layer3_outputs(1309);
    layer4_outputs(10110) <= layer3_outputs(3710);
    layer4_outputs(10111) <= (layer3_outputs(6931)) and (layer3_outputs(5326));
    layer4_outputs(10112) <= not(layer3_outputs(9372));
    layer4_outputs(10113) <= layer3_outputs(5774);
    layer4_outputs(10114) <= layer3_outputs(7262);
    layer4_outputs(10115) <= layer3_outputs(1548);
    layer4_outputs(10116) <= layer3_outputs(1201);
    layer4_outputs(10117) <= '0';
    layer4_outputs(10118) <= not(layer3_outputs(9030)) or (layer3_outputs(7307));
    layer4_outputs(10119) <= layer3_outputs(6740);
    layer4_outputs(10120) <= layer3_outputs(8985);
    layer4_outputs(10121) <= layer3_outputs(2123);
    layer4_outputs(10122) <= not(layer3_outputs(3388));
    layer4_outputs(10123) <= (layer3_outputs(6878)) or (layer3_outputs(8529));
    layer4_outputs(10124) <= (layer3_outputs(9863)) and not (layer3_outputs(6747));
    layer4_outputs(10125) <= not(layer3_outputs(4081));
    layer4_outputs(10126) <= layer3_outputs(2468);
    layer4_outputs(10127) <= not(layer3_outputs(6533));
    layer4_outputs(10128) <= layer3_outputs(6626);
    layer4_outputs(10129) <= (layer3_outputs(1256)) and not (layer3_outputs(2910));
    layer4_outputs(10130) <= not((layer3_outputs(704)) xor (layer3_outputs(8443)));
    layer4_outputs(10131) <= layer3_outputs(5084);
    layer4_outputs(10132) <= '0';
    layer4_outputs(10133) <= (layer3_outputs(9474)) xor (layer3_outputs(6296));
    layer4_outputs(10134) <= not(layer3_outputs(7218)) or (layer3_outputs(986));
    layer4_outputs(10135) <= not((layer3_outputs(78)) xor (layer3_outputs(4252)));
    layer4_outputs(10136) <= layer3_outputs(8833);
    layer4_outputs(10137) <= (layer3_outputs(417)) xor (layer3_outputs(5064));
    layer4_outputs(10138) <= layer3_outputs(8172);
    layer4_outputs(10139) <= layer3_outputs(6920);
    layer4_outputs(10140) <= (layer3_outputs(371)) and (layer3_outputs(6415));
    layer4_outputs(10141) <= layer3_outputs(3308);
    layer4_outputs(10142) <= layer3_outputs(8908);
    layer4_outputs(10143) <= not(layer3_outputs(8832)) or (layer3_outputs(9174));
    layer4_outputs(10144) <= not((layer3_outputs(2295)) xor (layer3_outputs(4472)));
    layer4_outputs(10145) <= (layer3_outputs(7223)) or (layer3_outputs(1663));
    layer4_outputs(10146) <= not(layer3_outputs(6008));
    layer4_outputs(10147) <= '0';
    layer4_outputs(10148) <= not(layer3_outputs(3751));
    layer4_outputs(10149) <= not((layer3_outputs(9617)) or (layer3_outputs(4059)));
    layer4_outputs(10150) <= not(layer3_outputs(4726)) or (layer3_outputs(8780));
    layer4_outputs(10151) <= not(layer3_outputs(3819));
    layer4_outputs(10152) <= layer3_outputs(8495);
    layer4_outputs(10153) <= layer3_outputs(8178);
    layer4_outputs(10154) <= layer3_outputs(7449);
    layer4_outputs(10155) <= not(layer3_outputs(9375));
    layer4_outputs(10156) <= not(layer3_outputs(2084));
    layer4_outputs(10157) <= not(layer3_outputs(1381));
    layer4_outputs(10158) <= not(layer3_outputs(7689));
    layer4_outputs(10159) <= (layer3_outputs(8326)) and not (layer3_outputs(5313));
    layer4_outputs(10160) <= not(layer3_outputs(7032));
    layer4_outputs(10161) <= not((layer3_outputs(6866)) xor (layer3_outputs(963)));
    layer4_outputs(10162) <= not(layer3_outputs(4605));
    layer4_outputs(10163) <= not(layer3_outputs(5668));
    layer4_outputs(10164) <= not(layer3_outputs(10130));
    layer4_outputs(10165) <= (layer3_outputs(6760)) xor (layer3_outputs(8247));
    layer4_outputs(10166) <= layer3_outputs(2022);
    layer4_outputs(10167) <= (layer3_outputs(8403)) and not (layer3_outputs(6245));
    layer4_outputs(10168) <= layer3_outputs(8197);
    layer4_outputs(10169) <= not(layer3_outputs(9961));
    layer4_outputs(10170) <= '0';
    layer4_outputs(10171) <= not(layer3_outputs(9672));
    layer4_outputs(10172) <= not(layer3_outputs(1868));
    layer4_outputs(10173) <= layer3_outputs(5276);
    layer4_outputs(10174) <= not(layer3_outputs(6196));
    layer4_outputs(10175) <= not(layer3_outputs(2942));
    layer4_outputs(10176) <= layer3_outputs(6881);
    layer4_outputs(10177) <= not((layer3_outputs(9591)) xor (layer3_outputs(3811)));
    layer4_outputs(10178) <= layer3_outputs(6263);
    layer4_outputs(10179) <= (layer3_outputs(1704)) and (layer3_outputs(6618));
    layer4_outputs(10180) <= (layer3_outputs(3670)) xor (layer3_outputs(10194));
    layer4_outputs(10181) <= not(layer3_outputs(758));
    layer4_outputs(10182) <= (layer3_outputs(8014)) or (layer3_outputs(477));
    layer4_outputs(10183) <= layer3_outputs(9976);
    layer4_outputs(10184) <= not((layer3_outputs(5554)) or (layer3_outputs(7929)));
    layer4_outputs(10185) <= not(layer3_outputs(3447));
    layer4_outputs(10186) <= not(layer3_outputs(5501));
    layer4_outputs(10187) <= (layer3_outputs(8618)) xor (layer3_outputs(8589));
    layer4_outputs(10188) <= not(layer3_outputs(3136));
    layer4_outputs(10189) <= layer3_outputs(2593);
    layer4_outputs(10190) <= not(layer3_outputs(698));
    layer4_outputs(10191) <= (layer3_outputs(8777)) xor (layer3_outputs(1629));
    layer4_outputs(10192) <= not(layer3_outputs(1827));
    layer4_outputs(10193) <= not(layer3_outputs(10067)) or (layer3_outputs(7164));
    layer4_outputs(10194) <= (layer3_outputs(8131)) and not (layer3_outputs(7045));
    layer4_outputs(10195) <= (layer3_outputs(974)) xor (layer3_outputs(770));
    layer4_outputs(10196) <= not((layer3_outputs(9669)) or (layer3_outputs(5748)));
    layer4_outputs(10197) <= not((layer3_outputs(7755)) or (layer3_outputs(10173)));
    layer4_outputs(10198) <= not(layer3_outputs(6776)) or (layer3_outputs(6413));
    layer4_outputs(10199) <= not(layer3_outputs(9964));
    layer4_outputs(10200) <= layer3_outputs(3227);
    layer4_outputs(10201) <= layer3_outputs(5250);
    layer4_outputs(10202) <= layer3_outputs(9552);
    layer4_outputs(10203) <= layer3_outputs(9887);
    layer4_outputs(10204) <= (layer3_outputs(7638)) xor (layer3_outputs(2793));
    layer4_outputs(10205) <= (layer3_outputs(9678)) and (layer3_outputs(764));
    layer4_outputs(10206) <= not(layer3_outputs(8415)) or (layer3_outputs(290));
    layer4_outputs(10207) <= not(layer3_outputs(7185));
    layer4_outputs(10208) <= (layer3_outputs(5509)) and not (layer3_outputs(814));
    layer4_outputs(10209) <= not(layer3_outputs(1802));
    layer4_outputs(10210) <= layer3_outputs(780);
    layer4_outputs(10211) <= not((layer3_outputs(9719)) xor (layer3_outputs(4864)));
    layer4_outputs(10212) <= not(layer3_outputs(8222));
    layer4_outputs(10213) <= not(layer3_outputs(243));
    layer4_outputs(10214) <= not(layer3_outputs(2866));
    layer4_outputs(10215) <= layer3_outputs(1123);
    layer4_outputs(10216) <= layer3_outputs(1685);
    layer4_outputs(10217) <= (layer3_outputs(9240)) and (layer3_outputs(1090));
    layer4_outputs(10218) <= not(layer3_outputs(956));
    layer4_outputs(10219) <= layer3_outputs(1307);
    layer4_outputs(10220) <= layer3_outputs(8487);
    layer4_outputs(10221) <= layer3_outputs(1343);
    layer4_outputs(10222) <= not(layer3_outputs(8239));
    layer4_outputs(10223) <= not(layer3_outputs(8244));
    layer4_outputs(10224) <= not(layer3_outputs(6730));
    layer4_outputs(10225) <= not((layer3_outputs(3169)) xor (layer3_outputs(9498)));
    layer4_outputs(10226) <= not(layer3_outputs(8107));
    layer4_outputs(10227) <= not(layer3_outputs(4181));
    layer4_outputs(10228) <= layer3_outputs(6358);
    layer4_outputs(10229) <= (layer3_outputs(1529)) and not (layer3_outputs(4970));
    layer4_outputs(10230) <= layer3_outputs(3225);
    layer4_outputs(10231) <= layer3_outputs(3687);
    layer4_outputs(10232) <= not(layer3_outputs(9835)) or (layer3_outputs(1571));
    layer4_outputs(10233) <= not(layer3_outputs(5289)) or (layer3_outputs(1410));
    layer4_outputs(10234) <= not(layer3_outputs(6550));
    layer4_outputs(10235) <= layer3_outputs(10014);
    layer4_outputs(10236) <= layer3_outputs(5867);
    layer4_outputs(10237) <= layer3_outputs(8860);
    layer4_outputs(10238) <= layer3_outputs(1305);
    layer4_outputs(10239) <= not(layer3_outputs(3290));
    outputs(0) <= layer4_outputs(2425);
    outputs(1) <= layer4_outputs(4804);
    outputs(2) <= (layer4_outputs(9896)) xor (layer4_outputs(4676));
    outputs(3) <= not(layer4_outputs(8498));
    outputs(4) <= layer4_outputs(1416);
    outputs(5) <= layer4_outputs(4222);
    outputs(6) <= not(layer4_outputs(2649));
    outputs(7) <= layer4_outputs(10183);
    outputs(8) <= not(layer4_outputs(2126));
    outputs(9) <= layer4_outputs(140);
    outputs(10) <= layer4_outputs(3000);
    outputs(11) <= layer4_outputs(9659);
    outputs(12) <= not(layer4_outputs(9949)) or (layer4_outputs(7089));
    outputs(13) <= not((layer4_outputs(9206)) xor (layer4_outputs(5535)));
    outputs(14) <= layer4_outputs(4987);
    outputs(15) <= layer4_outputs(895);
    outputs(16) <= (layer4_outputs(4861)) xor (layer4_outputs(7484));
    outputs(17) <= not((layer4_outputs(7819)) and (layer4_outputs(8583)));
    outputs(18) <= (layer4_outputs(9563)) xor (layer4_outputs(8465));
    outputs(19) <= layer4_outputs(10100);
    outputs(20) <= (layer4_outputs(8484)) xor (layer4_outputs(1452));
    outputs(21) <= layer4_outputs(8632);
    outputs(22) <= not(layer4_outputs(1931));
    outputs(23) <= layer4_outputs(6571);
    outputs(24) <= (layer4_outputs(7231)) xor (layer4_outputs(3861));
    outputs(25) <= not(layer4_outputs(7552)) or (layer4_outputs(9812));
    outputs(26) <= layer4_outputs(7953);
    outputs(27) <= layer4_outputs(2871);
    outputs(28) <= not((layer4_outputs(3176)) xor (layer4_outputs(5194)));
    outputs(29) <= not((layer4_outputs(6065)) or (layer4_outputs(6405)));
    outputs(30) <= not(layer4_outputs(8394));
    outputs(31) <= layer4_outputs(7524);
    outputs(32) <= (layer4_outputs(204)) or (layer4_outputs(3117));
    outputs(33) <= layer4_outputs(481);
    outputs(34) <= not(layer4_outputs(9828)) or (layer4_outputs(7395));
    outputs(35) <= not(layer4_outputs(3914));
    outputs(36) <= layer4_outputs(138);
    outputs(37) <= not(layer4_outputs(7750));
    outputs(38) <= not(layer4_outputs(227));
    outputs(39) <= not(layer4_outputs(2387));
    outputs(40) <= layer4_outputs(1818);
    outputs(41) <= not(layer4_outputs(8673));
    outputs(42) <= layer4_outputs(7961);
    outputs(43) <= layer4_outputs(2259);
    outputs(44) <= (layer4_outputs(6388)) xor (layer4_outputs(2493));
    outputs(45) <= (layer4_outputs(4452)) xor (layer4_outputs(4527));
    outputs(46) <= layer4_outputs(8735);
    outputs(47) <= (layer4_outputs(4746)) xor (layer4_outputs(7736));
    outputs(48) <= (layer4_outputs(2271)) xor (layer4_outputs(10234));
    outputs(49) <= not(layer4_outputs(9192));
    outputs(50) <= not(layer4_outputs(453));
    outputs(51) <= not(layer4_outputs(3153)) or (layer4_outputs(7857));
    outputs(52) <= not((layer4_outputs(3451)) xor (layer4_outputs(9453)));
    outputs(53) <= not(layer4_outputs(2974));
    outputs(54) <= layer4_outputs(1380);
    outputs(55) <= not((layer4_outputs(4386)) xor (layer4_outputs(1809)));
    outputs(56) <= not(layer4_outputs(6594));
    outputs(57) <= layer4_outputs(5404);
    outputs(58) <= not((layer4_outputs(5320)) or (layer4_outputs(9119)));
    outputs(59) <= not(layer4_outputs(7086));
    outputs(60) <= not(layer4_outputs(3871)) or (layer4_outputs(5391));
    outputs(61) <= not((layer4_outputs(8966)) and (layer4_outputs(6023)));
    outputs(62) <= (layer4_outputs(8633)) xor (layer4_outputs(7442));
    outputs(63) <= (layer4_outputs(1494)) and (layer4_outputs(8068));
    outputs(64) <= not(layer4_outputs(8022));
    outputs(65) <= not(layer4_outputs(6297));
    outputs(66) <= layer4_outputs(2976);
    outputs(67) <= not(layer4_outputs(3980));
    outputs(68) <= layer4_outputs(3684);
    outputs(69) <= layer4_outputs(10036);
    outputs(70) <= (layer4_outputs(5771)) xor (layer4_outputs(707));
    outputs(71) <= not(layer4_outputs(9601));
    outputs(72) <= not((layer4_outputs(715)) xor (layer4_outputs(9030)));
    outputs(73) <= (layer4_outputs(3860)) or (layer4_outputs(9993));
    outputs(74) <= layer4_outputs(5948);
    outputs(75) <= layer4_outputs(7928);
    outputs(76) <= not(layer4_outputs(5830));
    outputs(77) <= not(layer4_outputs(6572)) or (layer4_outputs(1475));
    outputs(78) <= layer4_outputs(1896);
    outputs(79) <= layer4_outputs(1467);
    outputs(80) <= not(layer4_outputs(6080));
    outputs(81) <= not((layer4_outputs(872)) xor (layer4_outputs(8424)));
    outputs(82) <= not(layer4_outputs(9911));
    outputs(83) <= layer4_outputs(9311);
    outputs(84) <= not((layer4_outputs(9148)) xor (layer4_outputs(7958)));
    outputs(85) <= layer4_outputs(1829);
    outputs(86) <= not(layer4_outputs(6893)) or (layer4_outputs(3628));
    outputs(87) <= layer4_outputs(2844);
    outputs(88) <= layer4_outputs(5177);
    outputs(89) <= layer4_outputs(8016);
    outputs(90) <= (layer4_outputs(2002)) and (layer4_outputs(8691));
    outputs(91) <= not(layer4_outputs(9875));
    outputs(92) <= not(layer4_outputs(6638));
    outputs(93) <= layer4_outputs(2665);
    outputs(94) <= not(layer4_outputs(9667));
    outputs(95) <= layer4_outputs(1226);
    outputs(96) <= not(layer4_outputs(408));
    outputs(97) <= (layer4_outputs(7073)) and not (layer4_outputs(4610));
    outputs(98) <= not((layer4_outputs(6949)) or (layer4_outputs(8482)));
    outputs(99) <= not((layer4_outputs(1785)) xor (layer4_outputs(7476)));
    outputs(100) <= not(layer4_outputs(8619));
    outputs(101) <= not(layer4_outputs(1296));
    outputs(102) <= (layer4_outputs(1906)) xor (layer4_outputs(2623));
    outputs(103) <= not(layer4_outputs(96));
    outputs(104) <= layer4_outputs(6071);
    outputs(105) <= layer4_outputs(4097);
    outputs(106) <= not(layer4_outputs(8308));
    outputs(107) <= not(layer4_outputs(6293));
    outputs(108) <= layer4_outputs(9690);
    outputs(109) <= not(layer4_outputs(6447));
    outputs(110) <= (layer4_outputs(2723)) or (layer4_outputs(9728));
    outputs(111) <= not((layer4_outputs(961)) or (layer4_outputs(9619)));
    outputs(112) <= not(layer4_outputs(7009));
    outputs(113) <= not(layer4_outputs(1686));
    outputs(114) <= not(layer4_outputs(3314));
    outputs(115) <= layer4_outputs(5253);
    outputs(116) <= not(layer4_outputs(9875));
    outputs(117) <= (layer4_outputs(7057)) or (layer4_outputs(7264));
    outputs(118) <= (layer4_outputs(3725)) and not (layer4_outputs(9876));
    outputs(119) <= not(layer4_outputs(3823));
    outputs(120) <= not(layer4_outputs(7353));
    outputs(121) <= not((layer4_outputs(8057)) xor (layer4_outputs(9186)));
    outputs(122) <= layer4_outputs(5736);
    outputs(123) <= layer4_outputs(3935);
    outputs(124) <= layer4_outputs(3197);
    outputs(125) <= layer4_outputs(8929);
    outputs(126) <= not(layer4_outputs(2168));
    outputs(127) <= not((layer4_outputs(4953)) xor (layer4_outputs(560)));
    outputs(128) <= layer4_outputs(5241);
    outputs(129) <= layer4_outputs(6849);
    outputs(130) <= not(layer4_outputs(3844)) or (layer4_outputs(8313));
    outputs(131) <= layer4_outputs(5237);
    outputs(132) <= not(layer4_outputs(8308));
    outputs(133) <= not(layer4_outputs(5060));
    outputs(134) <= layer4_outputs(6774);
    outputs(135) <= (layer4_outputs(4609)) xor (layer4_outputs(3487));
    outputs(136) <= not((layer4_outputs(5992)) xor (layer4_outputs(2933)));
    outputs(137) <= layer4_outputs(4550);
    outputs(138) <= layer4_outputs(9639);
    outputs(139) <= not(layer4_outputs(6461));
    outputs(140) <= not(layer4_outputs(2473));
    outputs(141) <= not(layer4_outputs(3042));
    outputs(142) <= not(layer4_outputs(3672));
    outputs(143) <= layer4_outputs(7280);
    outputs(144) <= not(layer4_outputs(1927));
    outputs(145) <= layer4_outputs(5044);
    outputs(146) <= layer4_outputs(2532);
    outputs(147) <= layer4_outputs(4439);
    outputs(148) <= not(layer4_outputs(9425));
    outputs(149) <= not((layer4_outputs(3867)) xor (layer4_outputs(7779)));
    outputs(150) <= (layer4_outputs(4334)) and not (layer4_outputs(456));
    outputs(151) <= (layer4_outputs(5700)) and not (layer4_outputs(6843));
    outputs(152) <= (layer4_outputs(9886)) xor (layer4_outputs(5388));
    outputs(153) <= not(layer4_outputs(8538));
    outputs(154) <= layer4_outputs(9281);
    outputs(155) <= (layer4_outputs(9484)) xor (layer4_outputs(783));
    outputs(156) <= layer4_outputs(8948);
    outputs(157) <= not((layer4_outputs(4075)) and (layer4_outputs(7485)));
    outputs(158) <= (layer4_outputs(393)) and (layer4_outputs(10218));
    outputs(159) <= not(layer4_outputs(5899));
    outputs(160) <= not(layer4_outputs(681));
    outputs(161) <= not(layer4_outputs(7157));
    outputs(162) <= not(layer4_outputs(4183));
    outputs(163) <= not(layer4_outputs(2704));
    outputs(164) <= not(layer4_outputs(8092));
    outputs(165) <= layer4_outputs(7962);
    outputs(166) <= not(layer4_outputs(9670));
    outputs(167) <= (layer4_outputs(6582)) or (layer4_outputs(6618));
    outputs(168) <= not(layer4_outputs(6474));
    outputs(169) <= layer4_outputs(1845);
    outputs(170) <= not(layer4_outputs(8263));
    outputs(171) <= layer4_outputs(1538);
    outputs(172) <= '0';
    outputs(173) <= layer4_outputs(8750);
    outputs(174) <= layer4_outputs(1100);
    outputs(175) <= (layer4_outputs(1559)) or (layer4_outputs(9358));
    outputs(176) <= not(layer4_outputs(4853));
    outputs(177) <= layer4_outputs(2357);
    outputs(178) <= layer4_outputs(10167);
    outputs(179) <= (layer4_outputs(6403)) or (layer4_outputs(9515));
    outputs(180) <= not(layer4_outputs(172));
    outputs(181) <= layer4_outputs(5339);
    outputs(182) <= (layer4_outputs(3069)) and (layer4_outputs(9524));
    outputs(183) <= layer4_outputs(8443);
    outputs(184) <= layer4_outputs(8153);
    outputs(185) <= not(layer4_outputs(1572));
    outputs(186) <= (layer4_outputs(4958)) or (layer4_outputs(6589));
    outputs(187) <= not(layer4_outputs(6934));
    outputs(188) <= layer4_outputs(6776);
    outputs(189) <= not((layer4_outputs(3175)) xor (layer4_outputs(4055)));
    outputs(190) <= not((layer4_outputs(2862)) xor (layer4_outputs(2781)));
    outputs(191) <= layer4_outputs(650);
    outputs(192) <= (layer4_outputs(9703)) xor (layer4_outputs(5160));
    outputs(193) <= layer4_outputs(8668);
    outputs(194) <= layer4_outputs(4658);
    outputs(195) <= layer4_outputs(1562);
    outputs(196) <= not((layer4_outputs(9618)) xor (layer4_outputs(4100)));
    outputs(197) <= not((layer4_outputs(2601)) xor (layer4_outputs(5693)));
    outputs(198) <= not((layer4_outputs(3809)) xor (layer4_outputs(5027)));
    outputs(199) <= layer4_outputs(1419);
    outputs(200) <= not(layer4_outputs(5738));
    outputs(201) <= not((layer4_outputs(2921)) xor (layer4_outputs(3434)));
    outputs(202) <= layer4_outputs(4263);
    outputs(203) <= not(layer4_outputs(1174));
    outputs(204) <= layer4_outputs(6378);
    outputs(205) <= not(layer4_outputs(2352));
    outputs(206) <= not(layer4_outputs(5710));
    outputs(207) <= layer4_outputs(770);
    outputs(208) <= layer4_outputs(6578);
    outputs(209) <= not(layer4_outputs(6336));
    outputs(210) <= layer4_outputs(8286);
    outputs(211) <= layer4_outputs(1848);
    outputs(212) <= layer4_outputs(9846);
    outputs(213) <= layer4_outputs(8566);
    outputs(214) <= not(layer4_outputs(5873));
    outputs(215) <= (layer4_outputs(8009)) xor (layer4_outputs(1686));
    outputs(216) <= not((layer4_outputs(6520)) and (layer4_outputs(4538)));
    outputs(217) <= not(layer4_outputs(6971)) or (layer4_outputs(9164));
    outputs(218) <= layer4_outputs(5021);
    outputs(219) <= not(layer4_outputs(2439));
    outputs(220) <= not((layer4_outputs(5158)) xor (layer4_outputs(9700)));
    outputs(221) <= not(layer4_outputs(3397));
    outputs(222) <= not((layer4_outputs(9612)) xor (layer4_outputs(1252)));
    outputs(223) <= layer4_outputs(5569);
    outputs(224) <= layer4_outputs(3403);
    outputs(225) <= layer4_outputs(6570);
    outputs(226) <= layer4_outputs(6671);
    outputs(227) <= not(layer4_outputs(686));
    outputs(228) <= (layer4_outputs(6616)) xor (layer4_outputs(9549));
    outputs(229) <= not(layer4_outputs(2970));
    outputs(230) <= not(layer4_outputs(9850));
    outputs(231) <= layer4_outputs(4785);
    outputs(232) <= layer4_outputs(8237);
    outputs(233) <= (layer4_outputs(10142)) xor (layer4_outputs(4160));
    outputs(234) <= not(layer4_outputs(2190));
    outputs(235) <= not(layer4_outputs(1976));
    outputs(236) <= not(layer4_outputs(7914)) or (layer4_outputs(8877));
    outputs(237) <= not((layer4_outputs(7768)) xor (layer4_outputs(9810)));
    outputs(238) <= layer4_outputs(6497);
    outputs(239) <= not(layer4_outputs(1381));
    outputs(240) <= not((layer4_outputs(2044)) xor (layer4_outputs(2073)));
    outputs(241) <= (layer4_outputs(2055)) and not (layer4_outputs(1765));
    outputs(242) <= not(layer4_outputs(7732));
    outputs(243) <= not(layer4_outputs(4627));
    outputs(244) <= layer4_outputs(5381);
    outputs(245) <= not(layer4_outputs(1679));
    outputs(246) <= layer4_outputs(4490);
    outputs(247) <= not(layer4_outputs(8533));
    outputs(248) <= not(layer4_outputs(4443)) or (layer4_outputs(8133));
    outputs(249) <= (layer4_outputs(9136)) and not (layer4_outputs(8297));
    outputs(250) <= not(layer4_outputs(4268));
    outputs(251) <= layer4_outputs(5568);
    outputs(252) <= (layer4_outputs(6549)) and not (layer4_outputs(10017));
    outputs(253) <= not(layer4_outputs(3599));
    outputs(254) <= layer4_outputs(5400);
    outputs(255) <= not(layer4_outputs(2152));
    outputs(256) <= not(layer4_outputs(3592));
    outputs(257) <= not(layer4_outputs(5512));
    outputs(258) <= (layer4_outputs(4405)) xor (layer4_outputs(7605));
    outputs(259) <= not(layer4_outputs(4556));
    outputs(260) <= not(layer4_outputs(2692));
    outputs(261) <= not(layer4_outputs(1437));
    outputs(262) <= not(layer4_outputs(2394));
    outputs(263) <= (layer4_outputs(76)) and (layer4_outputs(8377));
    outputs(264) <= layer4_outputs(6295);
    outputs(265) <= layer4_outputs(2611);
    outputs(266) <= layer4_outputs(7743);
    outputs(267) <= not(layer4_outputs(6718));
    outputs(268) <= not(layer4_outputs(2852));
    outputs(269) <= not(layer4_outputs(6506));
    outputs(270) <= (layer4_outputs(4615)) xor (layer4_outputs(6416));
    outputs(271) <= not(layer4_outputs(4947));
    outputs(272) <= not(layer4_outputs(7238));
    outputs(273) <= not(layer4_outputs(5098));
    outputs(274) <= layer4_outputs(5030);
    outputs(275) <= (layer4_outputs(10201)) xor (layer4_outputs(3280));
    outputs(276) <= not((layer4_outputs(9963)) xor (layer4_outputs(3358)));
    outputs(277) <= not(layer4_outputs(4674));
    outputs(278) <= layer4_outputs(7462);
    outputs(279) <= not((layer4_outputs(624)) and (layer4_outputs(4922)));
    outputs(280) <= layer4_outputs(3742);
    outputs(281) <= layer4_outputs(78);
    outputs(282) <= layer4_outputs(6806);
    outputs(283) <= (layer4_outputs(6344)) and not (layer4_outputs(1106));
    outputs(284) <= not(layer4_outputs(3177));
    outputs(285) <= not(layer4_outputs(7067));
    outputs(286) <= layer4_outputs(5751);
    outputs(287) <= (layer4_outputs(5813)) xor (layer4_outputs(6126));
    outputs(288) <= not(layer4_outputs(9036));
    outputs(289) <= layer4_outputs(2667);
    outputs(290) <= not(layer4_outputs(4959));
    outputs(291) <= not(layer4_outputs(1137));
    outputs(292) <= layer4_outputs(1636);
    outputs(293) <= layer4_outputs(3946);
    outputs(294) <= (layer4_outputs(1968)) and (layer4_outputs(8939));
    outputs(295) <= not(layer4_outputs(2705));
    outputs(296) <= (layer4_outputs(5411)) and not (layer4_outputs(4786));
    outputs(297) <= not(layer4_outputs(9856));
    outputs(298) <= layer4_outputs(6713);
    outputs(299) <= not(layer4_outputs(6893));
    outputs(300) <= (layer4_outputs(1135)) xor (layer4_outputs(7642));
    outputs(301) <= layer4_outputs(6876);
    outputs(302) <= layer4_outputs(9212);
    outputs(303) <= layer4_outputs(4494);
    outputs(304) <= (layer4_outputs(7243)) and (layer4_outputs(9873));
    outputs(305) <= not((layer4_outputs(10064)) xor (layer4_outputs(5137)));
    outputs(306) <= (layer4_outputs(4159)) xor (layer4_outputs(9910));
    outputs(307) <= '0';
    outputs(308) <= layer4_outputs(3546);
    outputs(309) <= (layer4_outputs(7570)) xor (layer4_outputs(7647));
    outputs(310) <= not((layer4_outputs(6999)) xor (layer4_outputs(4341)));
    outputs(311) <= not(layer4_outputs(7387));
    outputs(312) <= layer4_outputs(2690);
    outputs(313) <= not(layer4_outputs(779));
    outputs(314) <= not((layer4_outputs(7631)) or (layer4_outputs(8175)));
    outputs(315) <= not((layer4_outputs(7266)) or (layer4_outputs(4685)));
    outputs(316) <= layer4_outputs(5751);
    outputs(317) <= (layer4_outputs(5584)) xor (layer4_outputs(7349));
    outputs(318) <= not(layer4_outputs(2214)) or (layer4_outputs(6855));
    outputs(319) <= layer4_outputs(4507);
    outputs(320) <= layer4_outputs(5971);
    outputs(321) <= layer4_outputs(9993);
    outputs(322) <= (layer4_outputs(3821)) xor (layer4_outputs(2413));
    outputs(323) <= not(layer4_outputs(9945));
    outputs(324) <= (layer4_outputs(3925)) xor (layer4_outputs(8552));
    outputs(325) <= not(layer4_outputs(8619));
    outputs(326) <= layer4_outputs(1779);
    outputs(327) <= not((layer4_outputs(6060)) xor (layer4_outputs(8075)));
    outputs(328) <= not(layer4_outputs(446));
    outputs(329) <= layer4_outputs(3676);
    outputs(330) <= not(layer4_outputs(6304));
    outputs(331) <= (layer4_outputs(9050)) and (layer4_outputs(8010));
    outputs(332) <= (layer4_outputs(4181)) or (layer4_outputs(8290));
    outputs(333) <= not(layer4_outputs(6979));
    outputs(334) <= not((layer4_outputs(9046)) xor (layer4_outputs(2192)));
    outputs(335) <= not(layer4_outputs(1274));
    outputs(336) <= layer4_outputs(4274);
    outputs(337) <= layer4_outputs(5496);
    outputs(338) <= not(layer4_outputs(3694));
    outputs(339) <= not((layer4_outputs(514)) and (layer4_outputs(2155)));
    outputs(340) <= (layer4_outputs(6026)) and (layer4_outputs(3199));
    outputs(341) <= not(layer4_outputs(9470));
    outputs(342) <= not(layer4_outputs(976));
    outputs(343) <= not(layer4_outputs(10083)) or (layer4_outputs(2808));
    outputs(344) <= (layer4_outputs(3705)) or (layer4_outputs(1566));
    outputs(345) <= not(layer4_outputs(249));
    outputs(346) <= layer4_outputs(3105);
    outputs(347) <= not(layer4_outputs(1630));
    outputs(348) <= layer4_outputs(596);
    outputs(349) <= not(layer4_outputs(8770));
    outputs(350) <= not(layer4_outputs(5989)) or (layer4_outputs(4305));
    outputs(351) <= not(layer4_outputs(6873));
    outputs(352) <= layer4_outputs(500);
    outputs(353) <= (layer4_outputs(7138)) xor (layer4_outputs(4525));
    outputs(354) <= layer4_outputs(7164);
    outputs(355) <= not(layer4_outputs(4522));
    outputs(356) <= not((layer4_outputs(7869)) xor (layer4_outputs(7045)));
    outputs(357) <= not((layer4_outputs(3904)) xor (layer4_outputs(5893)));
    outputs(358) <= not(layer4_outputs(4483));
    outputs(359) <= layer4_outputs(826);
    outputs(360) <= layer4_outputs(1644);
    outputs(361) <= (layer4_outputs(1947)) and (layer4_outputs(3256));
    outputs(362) <= layer4_outputs(1235);
    outputs(363) <= layer4_outputs(318);
    outputs(364) <= not(layer4_outputs(7619));
    outputs(365) <= (layer4_outputs(1119)) xor (layer4_outputs(9043));
    outputs(366) <= not((layer4_outputs(4969)) and (layer4_outputs(5328)));
    outputs(367) <= not((layer4_outputs(5002)) or (layer4_outputs(169)));
    outputs(368) <= layer4_outputs(7268);
    outputs(369) <= layer4_outputs(3012);
    outputs(370) <= not(layer4_outputs(6863));
    outputs(371) <= layer4_outputs(2081);
    outputs(372) <= not((layer4_outputs(2833)) or (layer4_outputs(8854)));
    outputs(373) <= not(layer4_outputs(8776));
    outputs(374) <= (layer4_outputs(8202)) xor (layer4_outputs(7289));
    outputs(375) <= layer4_outputs(881);
    outputs(376) <= layer4_outputs(868);
    outputs(377) <= not(layer4_outputs(10215));
    outputs(378) <= layer4_outputs(729);
    outputs(379) <= layer4_outputs(6670);
    outputs(380) <= (layer4_outputs(4539)) xor (layer4_outputs(5679));
    outputs(381) <= (layer4_outputs(1392)) and not (layer4_outputs(3474));
    outputs(382) <= layer4_outputs(4721);
    outputs(383) <= not(layer4_outputs(8075));
    outputs(384) <= not((layer4_outputs(4584)) xor (layer4_outputs(2960)));
    outputs(385) <= not(layer4_outputs(2335));
    outputs(386) <= not(layer4_outputs(272));
    outputs(387) <= layer4_outputs(9821);
    outputs(388) <= not((layer4_outputs(8900)) xor (layer4_outputs(1831)));
    outputs(389) <= layer4_outputs(714);
    outputs(390) <= not(layer4_outputs(4108));
    outputs(391) <= not(layer4_outputs(6994));
    outputs(392) <= not(layer4_outputs(7735));
    outputs(393) <= layer4_outputs(4957);
    outputs(394) <= not(layer4_outputs(5710));
    outputs(395) <= not((layer4_outputs(7959)) xor (layer4_outputs(6433)));
    outputs(396) <= layer4_outputs(9241);
    outputs(397) <= not(layer4_outputs(3965));
    outputs(398) <= not(layer4_outputs(9522));
    outputs(399) <= not((layer4_outputs(5981)) xor (layer4_outputs(7086)));
    outputs(400) <= not(layer4_outputs(6956));
    outputs(401) <= layer4_outputs(1516);
    outputs(402) <= not(layer4_outputs(319));
    outputs(403) <= not(layer4_outputs(7405));
    outputs(404) <= not(layer4_outputs(930));
    outputs(405) <= not(layer4_outputs(2435)) or (layer4_outputs(3427));
    outputs(406) <= (layer4_outputs(8613)) xor (layer4_outputs(8199));
    outputs(407) <= not(layer4_outputs(8000));
    outputs(408) <= (layer4_outputs(6348)) and (layer4_outputs(4611));
    outputs(409) <= not(layer4_outputs(8505));
    outputs(410) <= (layer4_outputs(3294)) xor (layer4_outputs(5117));
    outputs(411) <= not(layer4_outputs(5800));
    outputs(412) <= layer4_outputs(931);
    outputs(413) <= layer4_outputs(369);
    outputs(414) <= not((layer4_outputs(5028)) xor (layer4_outputs(6073)));
    outputs(415) <= not(layer4_outputs(1742));
    outputs(416) <= not(layer4_outputs(5485)) or (layer4_outputs(2625));
    outputs(417) <= not((layer4_outputs(9256)) xor (layer4_outputs(4611)));
    outputs(418) <= (layer4_outputs(2331)) xor (layer4_outputs(3590));
    outputs(419) <= (layer4_outputs(7194)) and not (layer4_outputs(6891));
    outputs(420) <= not(layer4_outputs(2475));
    outputs(421) <= not(layer4_outputs(10094));
    outputs(422) <= not(layer4_outputs(10015));
    outputs(423) <= not(layer4_outputs(10154));
    outputs(424) <= not((layer4_outputs(1487)) or (layer4_outputs(7723)));
    outputs(425) <= not(layer4_outputs(10185));
    outputs(426) <= layer4_outputs(2533);
    outputs(427) <= (layer4_outputs(6361)) xor (layer4_outputs(4601));
    outputs(428) <= not(layer4_outputs(1300));
    outputs(429) <= not(layer4_outputs(6538));
    outputs(430) <= layer4_outputs(9263);
    outputs(431) <= not(layer4_outputs(2780));
    outputs(432) <= not(layer4_outputs(2702));
    outputs(433) <= not(layer4_outputs(4085));
    outputs(434) <= layer4_outputs(1164);
    outputs(435) <= layer4_outputs(3022);
    outputs(436) <= (layer4_outputs(5269)) xor (layer4_outputs(1325));
    outputs(437) <= layer4_outputs(3744);
    outputs(438) <= layer4_outputs(1237);
    outputs(439) <= layer4_outputs(1656);
    outputs(440) <= not(layer4_outputs(4083));
    outputs(441) <= layer4_outputs(3760);
    outputs(442) <= (layer4_outputs(2299)) and not (layer4_outputs(4143));
    outputs(443) <= not(layer4_outputs(1382));
    outputs(444) <= not(layer4_outputs(997));
    outputs(445) <= (layer4_outputs(7569)) and (layer4_outputs(9620));
    outputs(446) <= not(layer4_outputs(2382));
    outputs(447) <= not(layer4_outputs(9425)) or (layer4_outputs(3735));
    outputs(448) <= not(layer4_outputs(611));
    outputs(449) <= (layer4_outputs(8876)) or (layer4_outputs(3338));
    outputs(450) <= (layer4_outputs(5582)) or (layer4_outputs(5159));
    outputs(451) <= not((layer4_outputs(1513)) and (layer4_outputs(2517)));
    outputs(452) <= not((layer4_outputs(293)) xor (layer4_outputs(5224)));
    outputs(453) <= (layer4_outputs(7998)) xor (layer4_outputs(1944));
    outputs(454) <= layer4_outputs(7681);
    outputs(455) <= layer4_outputs(1573);
    outputs(456) <= layer4_outputs(4823);
    outputs(457) <= not((layer4_outputs(4995)) xor (layer4_outputs(6439)));
    outputs(458) <= not((layer4_outputs(4999)) and (layer4_outputs(4890)));
    outputs(459) <= not(layer4_outputs(4185));
    outputs(460) <= not((layer4_outputs(276)) xor (layer4_outputs(9194)));
    outputs(461) <= layer4_outputs(6997);
    outputs(462) <= not(layer4_outputs(5595));
    outputs(463) <= (layer4_outputs(254)) or (layer4_outputs(8349));
    outputs(464) <= not(layer4_outputs(4328));
    outputs(465) <= layer4_outputs(5318);
    outputs(466) <= not((layer4_outputs(6464)) and (layer4_outputs(4095)));
    outputs(467) <= (layer4_outputs(602)) and not (layer4_outputs(6312));
    outputs(468) <= not((layer4_outputs(3246)) and (layer4_outputs(5486)));
    outputs(469) <= layer4_outputs(2092);
    outputs(470) <= not(layer4_outputs(4260));
    outputs(471) <= not(layer4_outputs(5873));
    outputs(472) <= (layer4_outputs(2291)) or (layer4_outputs(5387));
    outputs(473) <= not(layer4_outputs(1632));
    outputs(474) <= not(layer4_outputs(7142));
    outputs(475) <= layer4_outputs(4420);
    outputs(476) <= layer4_outputs(5827);
    outputs(477) <= layer4_outputs(8512);
    outputs(478) <= not(layer4_outputs(3606));
    outputs(479) <= layer4_outputs(6382);
    outputs(480) <= (layer4_outputs(2160)) xor (layer4_outputs(5380));
    outputs(481) <= layer4_outputs(5742);
    outputs(482) <= not(layer4_outputs(7852));
    outputs(483) <= layer4_outputs(2830);
    outputs(484) <= layer4_outputs(7985);
    outputs(485) <= not((layer4_outputs(7179)) xor (layer4_outputs(2545)));
    outputs(486) <= not(layer4_outputs(7897));
    outputs(487) <= not(layer4_outputs(4369));
    outputs(488) <= (layer4_outputs(2509)) and not (layer4_outputs(6322));
    outputs(489) <= (layer4_outputs(7376)) and (layer4_outputs(3661));
    outputs(490) <= layer4_outputs(8276);
    outputs(491) <= (layer4_outputs(4127)) and not (layer4_outputs(5912));
    outputs(492) <= not(layer4_outputs(3185));
    outputs(493) <= layer4_outputs(8559);
    outputs(494) <= layer4_outputs(5310);
    outputs(495) <= layer4_outputs(4817);
    outputs(496) <= not((layer4_outputs(9840)) xor (layer4_outputs(9876)));
    outputs(497) <= not(layer4_outputs(5032));
    outputs(498) <= not(layer4_outputs(4214));
    outputs(499) <= not(layer4_outputs(2469));
    outputs(500) <= (layer4_outputs(2525)) xor (layer4_outputs(2340));
    outputs(501) <= not(layer4_outputs(9787));
    outputs(502) <= (layer4_outputs(4007)) or (layer4_outputs(2869));
    outputs(503) <= not(layer4_outputs(4952));
    outputs(504) <= layer4_outputs(9537);
    outputs(505) <= layer4_outputs(4174);
    outputs(506) <= layer4_outputs(8865);
    outputs(507) <= not(layer4_outputs(1032));
    outputs(508) <= not(layer4_outputs(6464));
    outputs(509) <= not((layer4_outputs(8611)) xor (layer4_outputs(5376)));
    outputs(510) <= layer4_outputs(2140);
    outputs(511) <= not(layer4_outputs(9368));
    outputs(512) <= layer4_outputs(7524);
    outputs(513) <= layer4_outputs(9100);
    outputs(514) <= (layer4_outputs(2541)) xor (layer4_outputs(9185));
    outputs(515) <= not(layer4_outputs(5309));
    outputs(516) <= (layer4_outputs(9238)) xor (layer4_outputs(8781));
    outputs(517) <= not(layer4_outputs(5402)) or (layer4_outputs(2292));
    outputs(518) <= (layer4_outputs(4147)) xor (layer4_outputs(9296));
    outputs(519) <= layer4_outputs(424);
    outputs(520) <= not((layer4_outputs(3042)) xor (layer4_outputs(2121)));
    outputs(521) <= (layer4_outputs(7938)) xor (layer4_outputs(775));
    outputs(522) <= not(layer4_outputs(4850));
    outputs(523) <= layer4_outputs(3143);
    outputs(524) <= not((layer4_outputs(4354)) xor (layer4_outputs(9947)));
    outputs(525) <= (layer4_outputs(4375)) and (layer4_outputs(7164));
    outputs(526) <= not(layer4_outputs(3335));
    outputs(527) <= not(layer4_outputs(1182));
    outputs(528) <= not(layer4_outputs(9979));
    outputs(529) <= not(layer4_outputs(7567));
    outputs(530) <= not(layer4_outputs(3150));
    outputs(531) <= not(layer4_outputs(1012)) or (layer4_outputs(5069));
    outputs(532) <= layer4_outputs(1301);
    outputs(533) <= not((layer4_outputs(6012)) xor (layer4_outputs(9994)));
    outputs(534) <= not(layer4_outputs(9202)) or (layer4_outputs(4741));
    outputs(535) <= layer4_outputs(5771);
    outputs(536) <= layer4_outputs(1520);
    outputs(537) <= not(layer4_outputs(5007));
    outputs(538) <= not(layer4_outputs(3549));
    outputs(539) <= not(layer4_outputs(6448));
    outputs(540) <= layer4_outputs(9462);
    outputs(541) <= layer4_outputs(6491);
    outputs(542) <= layer4_outputs(2863);
    outputs(543) <= (layer4_outputs(1568)) xor (layer4_outputs(168));
    outputs(544) <= layer4_outputs(7158);
    outputs(545) <= not((layer4_outputs(7194)) xor (layer4_outputs(9606)));
    outputs(546) <= not((layer4_outputs(9943)) and (layer4_outputs(4149)));
    outputs(547) <= not(layer4_outputs(8334));
    outputs(548) <= not(layer4_outputs(2556));
    outputs(549) <= not(layer4_outputs(4934));
    outputs(550) <= (layer4_outputs(2965)) xor (layer4_outputs(8641));
    outputs(551) <= layer4_outputs(2065);
    outputs(552) <= not(layer4_outputs(9284));
    outputs(553) <= layer4_outputs(7036);
    outputs(554) <= not(layer4_outputs(2255));
    outputs(555) <= layer4_outputs(271);
    outputs(556) <= not(layer4_outputs(7523));
    outputs(557) <= layer4_outputs(3681);
    outputs(558) <= not((layer4_outputs(3001)) and (layer4_outputs(5860)));
    outputs(559) <= not(layer4_outputs(6661));
    outputs(560) <= layer4_outputs(6613);
    outputs(561) <= not((layer4_outputs(4109)) xor (layer4_outputs(7597)));
    outputs(562) <= layer4_outputs(7180);
    outputs(563) <= not((layer4_outputs(5068)) or (layer4_outputs(285)));
    outputs(564) <= not(layer4_outputs(5941));
    outputs(565) <= not(layer4_outputs(9973)) or (layer4_outputs(3193));
    outputs(566) <= not(layer4_outputs(4251));
    outputs(567) <= not(layer4_outputs(7146));
    outputs(568) <= layer4_outputs(3926);
    outputs(569) <= not(layer4_outputs(9323));
    outputs(570) <= not(layer4_outputs(250));
    outputs(571) <= (layer4_outputs(9124)) xor (layer4_outputs(5132));
    outputs(572) <= not(layer4_outputs(98)) or (layer4_outputs(5956));
    outputs(573) <= (layer4_outputs(2785)) xor (layer4_outputs(2310));
    outputs(574) <= not((layer4_outputs(7121)) xor (layer4_outputs(7776)));
    outputs(575) <= (layer4_outputs(989)) xor (layer4_outputs(1393));
    outputs(576) <= layer4_outputs(6734);
    outputs(577) <= layer4_outputs(7439);
    outputs(578) <= not((layer4_outputs(4161)) xor (layer4_outputs(8869)));
    outputs(579) <= layer4_outputs(5284);
    outputs(580) <= layer4_outputs(9745);
    outputs(581) <= layer4_outputs(9962);
    outputs(582) <= layer4_outputs(264);
    outputs(583) <= layer4_outputs(9398);
    outputs(584) <= layer4_outputs(671);
    outputs(585) <= not(layer4_outputs(7785));
    outputs(586) <= layer4_outputs(1915);
    outputs(587) <= layer4_outputs(542);
    outputs(588) <= layer4_outputs(20);
    outputs(589) <= not(layer4_outputs(726)) or (layer4_outputs(2955));
    outputs(590) <= not(layer4_outputs(2816));
    outputs(591) <= layer4_outputs(3792);
    outputs(592) <= (layer4_outputs(6952)) and (layer4_outputs(5510));
    outputs(593) <= not(layer4_outputs(359)) or (layer4_outputs(5712));
    outputs(594) <= not(layer4_outputs(6802));
    outputs(595) <= (layer4_outputs(1413)) and (layer4_outputs(9540));
    outputs(596) <= not(layer4_outputs(8804));
    outputs(597) <= layer4_outputs(3826);
    outputs(598) <= layer4_outputs(2410);
    outputs(599) <= not(layer4_outputs(9814));
    outputs(600) <= not(layer4_outputs(3708)) or (layer4_outputs(8456));
    outputs(601) <= layer4_outputs(7806);
    outputs(602) <= layer4_outputs(1234);
    outputs(603) <= layer4_outputs(4139);
    outputs(604) <= not(layer4_outputs(1105));
    outputs(605) <= not(layer4_outputs(5034)) or (layer4_outputs(952));
    outputs(606) <= not(layer4_outputs(1843));
    outputs(607) <= layer4_outputs(6703);
    outputs(608) <= not(layer4_outputs(4084));
    outputs(609) <= not((layer4_outputs(7351)) xor (layer4_outputs(8436)));
    outputs(610) <= not(layer4_outputs(4478));
    outputs(611) <= (layer4_outputs(9594)) xor (layer4_outputs(3807));
    outputs(612) <= layer4_outputs(156);
    outputs(613) <= layer4_outputs(5104);
    outputs(614) <= not(layer4_outputs(8658));
    outputs(615) <= (layer4_outputs(8890)) or (layer4_outputs(1283));
    outputs(616) <= not((layer4_outputs(7256)) xor (layer4_outputs(316)));
    outputs(617) <= layer4_outputs(3296);
    outputs(618) <= layer4_outputs(239);
    outputs(619) <= not((layer4_outputs(6014)) xor (layer4_outputs(6243)));
    outputs(620) <= not(layer4_outputs(3041));
    outputs(621) <= (layer4_outputs(2432)) xor (layer4_outputs(4493));
    outputs(622) <= layer4_outputs(3169);
    outputs(623) <= not(layer4_outputs(9418));
    outputs(624) <= (layer4_outputs(6820)) or (layer4_outputs(6900));
    outputs(625) <= layer4_outputs(7346);
    outputs(626) <= not(layer4_outputs(8968)) or (layer4_outputs(8878));
    outputs(627) <= not(layer4_outputs(973));
    outputs(628) <= layer4_outputs(3275);
    outputs(629) <= layer4_outputs(2233);
    outputs(630) <= not(layer4_outputs(5821));
    outputs(631) <= (layer4_outputs(2535)) xor (layer4_outputs(6753));
    outputs(632) <= layer4_outputs(8606);
    outputs(633) <= layer4_outputs(8430);
    outputs(634) <= layer4_outputs(6696);
    outputs(635) <= not(layer4_outputs(6974));
    outputs(636) <= layer4_outputs(2929);
    outputs(637) <= (layer4_outputs(1806)) xor (layer4_outputs(5528));
    outputs(638) <= layer4_outputs(9485);
    outputs(639) <= not((layer4_outputs(6249)) and (layer4_outputs(9743)));
    outputs(640) <= not(layer4_outputs(1423));
    outputs(641) <= (layer4_outputs(213)) xor (layer4_outputs(3079));
    outputs(642) <= not(layer4_outputs(5628));
    outputs(643) <= not(layer4_outputs(9818));
    outputs(644) <= (layer4_outputs(4566)) or (layer4_outputs(4089));
    outputs(645) <= (layer4_outputs(5457)) xor (layer4_outputs(7541));
    outputs(646) <= not((layer4_outputs(1166)) xor (layer4_outputs(544)));
    outputs(647) <= not(layer4_outputs(3993));
    outputs(648) <= layer4_outputs(9121);
    outputs(649) <= not(layer4_outputs(9725));
    outputs(650) <= layer4_outputs(4180);
    outputs(651) <= (layer4_outputs(8956)) or (layer4_outputs(1396));
    outputs(652) <= not(layer4_outputs(4329));
    outputs(653) <= not(layer4_outputs(9595));
    outputs(654) <= (layer4_outputs(1781)) or (layer4_outputs(1039));
    outputs(655) <= not((layer4_outputs(5767)) xor (layer4_outputs(8022)));
    outputs(656) <= layer4_outputs(6198);
    outputs(657) <= layer4_outputs(9136);
    outputs(658) <= layer4_outputs(7295);
    outputs(659) <= not(layer4_outputs(6580)) or (layer4_outputs(4699));
    outputs(660) <= not(layer4_outputs(6745));
    outputs(661) <= layer4_outputs(10205);
    outputs(662) <= not((layer4_outputs(8612)) or (layer4_outputs(1835)));
    outputs(663) <= layer4_outputs(3478);
    outputs(664) <= not(layer4_outputs(5059));
    outputs(665) <= (layer4_outputs(4993)) or (layer4_outputs(7187));
    outputs(666) <= (layer4_outputs(860)) or (layer4_outputs(7183));
    outputs(667) <= not(layer4_outputs(1704)) or (layer4_outputs(3593));
    outputs(668) <= not((layer4_outputs(1618)) xor (layer4_outputs(2413)));
    outputs(669) <= layer4_outputs(4569);
    outputs(670) <= layer4_outputs(7864);
    outputs(671) <= (layer4_outputs(8002)) and not (layer4_outputs(2019));
    outputs(672) <= (layer4_outputs(4707)) and not (layer4_outputs(4838));
    outputs(673) <= not(layer4_outputs(3340));
    outputs(674) <= not(layer4_outputs(4454)) or (layer4_outputs(4224));
    outputs(675) <= layer4_outputs(2729);
    outputs(676) <= (layer4_outputs(9128)) and (layer4_outputs(3880));
    outputs(677) <= layer4_outputs(53);
    outputs(678) <= layer4_outputs(1464);
    outputs(679) <= not((layer4_outputs(2936)) xor (layer4_outputs(1060)));
    outputs(680) <= not(layer4_outputs(5786));
    outputs(681) <= not(layer4_outputs(5635));
    outputs(682) <= not(layer4_outputs(1344)) or (layer4_outputs(724));
    outputs(683) <= not(layer4_outputs(3602)) or (layer4_outputs(2218));
    outputs(684) <= not(layer4_outputs(2982));
    outputs(685) <= layer4_outputs(9990);
    outputs(686) <= layer4_outputs(6961);
    outputs(687) <= layer4_outputs(5939);
    outputs(688) <= (layer4_outputs(538)) xor (layer4_outputs(3418));
    outputs(689) <= not(layer4_outputs(421));
    outputs(690) <= layer4_outputs(2311);
    outputs(691) <= not(layer4_outputs(3515)) or (layer4_outputs(786));
    outputs(692) <= layer4_outputs(5556);
    outputs(693) <= layer4_outputs(6820);
    outputs(694) <= not(layer4_outputs(1087));
    outputs(695) <= (layer4_outputs(9360)) xor (layer4_outputs(1501));
    outputs(696) <= not((layer4_outputs(7213)) or (layer4_outputs(8400)));
    outputs(697) <= not(layer4_outputs(1043));
    outputs(698) <= layer4_outputs(943);
    outputs(699) <= (layer4_outputs(2358)) and (layer4_outputs(6367));
    outputs(700) <= not(layer4_outputs(9187));
    outputs(701) <= not(layer4_outputs(6247));
    outputs(702) <= layer4_outputs(6604);
    outputs(703) <= (layer4_outputs(9956)) xor (layer4_outputs(7734));
    outputs(704) <= layer4_outputs(2311);
    outputs(705) <= layer4_outputs(3081);
    outputs(706) <= (layer4_outputs(3521)) xor (layer4_outputs(8622));
    outputs(707) <= not((layer4_outputs(5011)) xor (layer4_outputs(5791)));
    outputs(708) <= layer4_outputs(3273);
    outputs(709) <= layer4_outputs(5752);
    outputs(710) <= not(layer4_outputs(5271));
    outputs(711) <= not(layer4_outputs(2620));
    outputs(712) <= (layer4_outputs(2599)) and not (layer4_outputs(7624));
    outputs(713) <= not(layer4_outputs(987));
    outputs(714) <= layer4_outputs(3395);
    outputs(715) <= layer4_outputs(6094);
    outputs(716) <= not(layer4_outputs(975));
    outputs(717) <= (layer4_outputs(10039)) xor (layer4_outputs(6606));
    outputs(718) <= layer4_outputs(93);
    outputs(719) <= not((layer4_outputs(6484)) xor (layer4_outputs(1758)));
    outputs(720) <= not(layer4_outputs(4680));
    outputs(721) <= not(layer4_outputs(9332)) or (layer4_outputs(4467));
    outputs(722) <= not(layer4_outputs(2562));
    outputs(723) <= layer4_outputs(8696);
    outputs(724) <= (layer4_outputs(3123)) and not (layer4_outputs(5251));
    outputs(725) <= (layer4_outputs(200)) or (layer4_outputs(1734));
    outputs(726) <= layer4_outputs(6373);
    outputs(727) <= not(layer4_outputs(1778));
    outputs(728) <= not(layer4_outputs(3775));
    outputs(729) <= not(layer4_outputs(5753));
    outputs(730) <= not(layer4_outputs(4072));
    outputs(731) <= not(layer4_outputs(7579));
    outputs(732) <= not((layer4_outputs(2036)) xor (layer4_outputs(7478)));
    outputs(733) <= layer4_outputs(4408);
    outputs(734) <= layer4_outputs(5006);
    outputs(735) <= not(layer4_outputs(6247));
    outputs(736) <= not(layer4_outputs(3175));
    outputs(737) <= not((layer4_outputs(5437)) xor (layer4_outputs(10170)));
    outputs(738) <= not(layer4_outputs(9600));
    outputs(739) <= not(layer4_outputs(1770));
    outputs(740) <= layer4_outputs(4046);
    outputs(741) <= not((layer4_outputs(7583)) and (layer4_outputs(6340)));
    outputs(742) <= not(layer4_outputs(5761)) or (layer4_outputs(3674));
    outputs(743) <= not((layer4_outputs(8037)) xor (layer4_outputs(4499)));
    outputs(744) <= not(layer4_outputs(8324)) or (layer4_outputs(2762));
    outputs(745) <= not((layer4_outputs(9560)) xor (layer4_outputs(5011)));
    outputs(746) <= (layer4_outputs(7170)) or (layer4_outputs(3023));
    outputs(747) <= layer4_outputs(7148);
    outputs(748) <= not(layer4_outputs(8169));
    outputs(749) <= not((layer4_outputs(2013)) xor (layer4_outputs(8664)));
    outputs(750) <= not((layer4_outputs(6291)) xor (layer4_outputs(3610)));
    outputs(751) <= not(layer4_outputs(7205));
    outputs(752) <= not(layer4_outputs(7942));
    outputs(753) <= not(layer4_outputs(3633));
    outputs(754) <= layer4_outputs(2369);
    outputs(755) <= '1';
    outputs(756) <= (layer4_outputs(1136)) and (layer4_outputs(8477));
    outputs(757) <= (layer4_outputs(4092)) or (layer4_outputs(5500));
    outputs(758) <= not((layer4_outputs(603)) or (layer4_outputs(4328)));
    outputs(759) <= not(layer4_outputs(5514));
    outputs(760) <= not(layer4_outputs(9340));
    outputs(761) <= not(layer4_outputs(2040));
    outputs(762) <= layer4_outputs(7196);
    outputs(763) <= not(layer4_outputs(5525));
    outputs(764) <= (layer4_outputs(8295)) and (layer4_outputs(7662));
    outputs(765) <= (layer4_outputs(317)) or (layer4_outputs(632));
    outputs(766) <= not((layer4_outputs(7494)) and (layer4_outputs(3950)));
    outputs(767) <= '0';
    outputs(768) <= (layer4_outputs(10113)) and not (layer4_outputs(1942));
    outputs(769) <= not(layer4_outputs(4128));
    outputs(770) <= (layer4_outputs(10135)) and not (layer4_outputs(5741));
    outputs(771) <= layer4_outputs(8782);
    outputs(772) <= not(layer4_outputs(8636));
    outputs(773) <= layer4_outputs(2922);
    outputs(774) <= not(layer4_outputs(13));
    outputs(775) <= (layer4_outputs(7314)) and (layer4_outputs(7408));
    outputs(776) <= not((layer4_outputs(1415)) xor (layer4_outputs(2143)));
    outputs(777) <= not((layer4_outputs(5844)) or (layer4_outputs(1102)));
    outputs(778) <= not(layer4_outputs(5667));
    outputs(779) <= not(layer4_outputs(1206));
    outputs(780) <= layer4_outputs(1293);
    outputs(781) <= not((layer4_outputs(3103)) xor (layer4_outputs(66)));
    outputs(782) <= not(layer4_outputs(8527));
    outputs(783) <= layer4_outputs(2922);
    outputs(784) <= (layer4_outputs(2084)) xor (layer4_outputs(5789));
    outputs(785) <= layer4_outputs(7653);
    outputs(786) <= layer4_outputs(10002);
    outputs(787) <= not(layer4_outputs(4048));
    outputs(788) <= not((layer4_outputs(7129)) xor (layer4_outputs(382)));
    outputs(789) <= (layer4_outputs(915)) and (layer4_outputs(345));
    outputs(790) <= layer4_outputs(10129);
    outputs(791) <= layer4_outputs(4038);
    outputs(792) <= layer4_outputs(5213);
    outputs(793) <= not(layer4_outputs(7282));
    outputs(794) <= layer4_outputs(9199);
    outputs(795) <= layer4_outputs(5335);
    outputs(796) <= not(layer4_outputs(8816));
    outputs(797) <= not((layer4_outputs(764)) xor (layer4_outputs(3981)));
    outputs(798) <= not(layer4_outputs(2168));
    outputs(799) <= not(layer4_outputs(639));
    outputs(800) <= '0';
    outputs(801) <= layer4_outputs(8850);
    outputs(802) <= layer4_outputs(5302);
    outputs(803) <= not(layer4_outputs(5484));
    outputs(804) <= layer4_outputs(1958);
    outputs(805) <= layer4_outputs(8061);
    outputs(806) <= not(layer4_outputs(7171));
    outputs(807) <= not(layer4_outputs(8310));
    outputs(808) <= layer4_outputs(7563);
    outputs(809) <= layer4_outputs(4249);
    outputs(810) <= not(layer4_outputs(6804));
    outputs(811) <= layer4_outputs(1314);
    outputs(812) <= layer4_outputs(7111);
    outputs(813) <= not((layer4_outputs(17)) xor (layer4_outputs(5590)));
    outputs(814) <= not(layer4_outputs(3993));
    outputs(815) <= not(layer4_outputs(10096));
    outputs(816) <= not(layer4_outputs(7023));
    outputs(817) <= not(layer4_outputs(1953));
    outputs(818) <= layer4_outputs(424);
    outputs(819) <= layer4_outputs(8050);
    outputs(820) <= not(layer4_outputs(4013));
    outputs(821) <= not((layer4_outputs(8712)) xor (layer4_outputs(9293)));
    outputs(822) <= (layer4_outputs(5982)) xor (layer4_outputs(9666));
    outputs(823) <= not(layer4_outputs(7004));
    outputs(824) <= not(layer4_outputs(7287)) or (layer4_outputs(2860));
    outputs(825) <= layer4_outputs(8974);
    outputs(826) <= layer4_outputs(3829);
    outputs(827) <= (layer4_outputs(2866)) and not (layer4_outputs(7878));
    outputs(828) <= not(layer4_outputs(8831));
    outputs(829) <= not(layer4_outputs(7078));
    outputs(830) <= not(layer4_outputs(1026));
    outputs(831) <= not(layer4_outputs(10180)) or (layer4_outputs(6736));
    outputs(832) <= not(layer4_outputs(7537));
    outputs(833) <= layer4_outputs(621);
    outputs(834) <= layer4_outputs(3261);
    outputs(835) <= layer4_outputs(7221);
    outputs(836) <= not(layer4_outputs(2536));
    outputs(837) <= layer4_outputs(1086);
    outputs(838) <= layer4_outputs(7226);
    outputs(839) <= (layer4_outputs(3703)) xor (layer4_outputs(2177));
    outputs(840) <= not((layer4_outputs(5508)) xor (layer4_outputs(5105)));
    outputs(841) <= layer4_outputs(9084);
    outputs(842) <= not(layer4_outputs(184));
    outputs(843) <= (layer4_outputs(5867)) xor (layer4_outputs(3757));
    outputs(844) <= not((layer4_outputs(5954)) and (layer4_outputs(9771)));
    outputs(845) <= (layer4_outputs(1214)) or (layer4_outputs(7111));
    outputs(846) <= layer4_outputs(4875);
    outputs(847) <= not(layer4_outputs(7972));
    outputs(848) <= not(layer4_outputs(27));
    outputs(849) <= not(layer4_outputs(4506));
    outputs(850) <= layer4_outputs(5638);
    outputs(851) <= layer4_outputs(1190);
    outputs(852) <= layer4_outputs(6808);
    outputs(853) <= layer4_outputs(1479);
    outputs(854) <= layer4_outputs(9153);
    outputs(855) <= not(layer4_outputs(2489));
    outputs(856) <= layer4_outputs(7361);
    outputs(857) <= layer4_outputs(2799);
    outputs(858) <= (layer4_outputs(6488)) xor (layer4_outputs(3997));
    outputs(859) <= not((layer4_outputs(1916)) xor (layer4_outputs(6395)));
    outputs(860) <= layer4_outputs(234);
    outputs(861) <= layer4_outputs(5510);
    outputs(862) <= layer4_outputs(9634);
    outputs(863) <= not(layer4_outputs(8189)) or (layer4_outputs(1213));
    outputs(864) <= not((layer4_outputs(5470)) and (layer4_outputs(3474)));
    outputs(865) <= not(layer4_outputs(5100));
    outputs(866) <= layer4_outputs(3181);
    outputs(867) <= not(layer4_outputs(5766));
    outputs(868) <= (layer4_outputs(4429)) xor (layer4_outputs(9559));
    outputs(869) <= layer4_outputs(1042);
    outputs(870) <= (layer4_outputs(9206)) and (layer4_outputs(3961));
    outputs(871) <= not(layer4_outputs(182));
    outputs(872) <= not(layer4_outputs(8594));
    outputs(873) <= layer4_outputs(6885);
    outputs(874) <= not(layer4_outputs(8110));
    outputs(875) <= not((layer4_outputs(4206)) and (layer4_outputs(5155)));
    outputs(876) <= not(layer4_outputs(6738));
    outputs(877) <= not(layer4_outputs(2557));
    outputs(878) <= (layer4_outputs(8980)) and not (layer4_outputs(4242));
    outputs(879) <= not(layer4_outputs(1509));
    outputs(880) <= not(layer4_outputs(2280));
    outputs(881) <= not(layer4_outputs(3927)) or (layer4_outputs(5943));
    outputs(882) <= not(layer4_outputs(3804));
    outputs(883) <= not(layer4_outputs(1299));
    outputs(884) <= layer4_outputs(4375);
    outputs(885) <= layer4_outputs(3635);
    outputs(886) <= layer4_outputs(2746);
    outputs(887) <= not(layer4_outputs(1730));
    outputs(888) <= not(layer4_outputs(1477)) or (layer4_outputs(2680));
    outputs(889) <= not(layer4_outputs(2501));
    outputs(890) <= not((layer4_outputs(4728)) xor (layer4_outputs(4626)));
    outputs(891) <= (layer4_outputs(569)) xor (layer4_outputs(1367));
    outputs(892) <= (layer4_outputs(6150)) xor (layer4_outputs(9215));
    outputs(893) <= layer4_outputs(9897);
    outputs(894) <= layer4_outputs(7662);
    outputs(895) <= layer4_outputs(9708);
    outputs(896) <= (layer4_outputs(7308)) xor (layer4_outputs(1800));
    outputs(897) <= not(layer4_outputs(10171));
    outputs(898) <= layer4_outputs(3483);
    outputs(899) <= not(layer4_outputs(5701));
    outputs(900) <= layer4_outputs(7948);
    outputs(901) <= not(layer4_outputs(6141));
    outputs(902) <= not(layer4_outputs(1210));
    outputs(903) <= not(layer4_outputs(5258));
    outputs(904) <= not((layer4_outputs(6678)) xor (layer4_outputs(2418)));
    outputs(905) <= not(layer4_outputs(4664));
    outputs(906) <= layer4_outputs(10160);
    outputs(907) <= layer4_outputs(9321);
    outputs(908) <= (layer4_outputs(3794)) xor (layer4_outputs(4964));
    outputs(909) <= not(layer4_outputs(6756));
    outputs(910) <= not(layer4_outputs(8824));
    outputs(911) <= layer4_outputs(2583);
    outputs(912) <= layer4_outputs(4377);
    outputs(913) <= layer4_outputs(5130);
    outputs(914) <= not(layer4_outputs(4702)) or (layer4_outputs(8590));
    outputs(915) <= not(layer4_outputs(7848)) or (layer4_outputs(8564));
    outputs(916) <= layer4_outputs(1246);
    outputs(917) <= not((layer4_outputs(4869)) xor (layer4_outputs(9627)));
    outputs(918) <= layer4_outputs(8513);
    outputs(919) <= not((layer4_outputs(7607)) xor (layer4_outputs(3423)));
    outputs(920) <= layer4_outputs(2824);
    outputs(921) <= not(layer4_outputs(10045));
    outputs(922) <= layer4_outputs(9338);
    outputs(923) <= not(layer4_outputs(1679));
    outputs(924) <= layer4_outputs(8711);
    outputs(925) <= (layer4_outputs(6962)) xor (layer4_outputs(864));
    outputs(926) <= (layer4_outputs(8641)) xor (layer4_outputs(9113));
    outputs(927) <= layer4_outputs(833);
    outputs(928) <= (layer4_outputs(2029)) and not (layer4_outputs(3072));
    outputs(929) <= layer4_outputs(7159);
    outputs(930) <= layer4_outputs(4127);
    outputs(931) <= not(layer4_outputs(7703));
    outputs(932) <= not(layer4_outputs(6724)) or (layer4_outputs(8073));
    outputs(933) <= layer4_outputs(10063);
    outputs(934) <= not(layer4_outputs(7445));
    outputs(935) <= layer4_outputs(587);
    outputs(936) <= layer4_outputs(1634);
    outputs(937) <= layer4_outputs(4476);
    outputs(938) <= layer4_outputs(364);
    outputs(939) <= layer4_outputs(7403);
    outputs(940) <= not(layer4_outputs(3366));
    outputs(941) <= not((layer4_outputs(385)) xor (layer4_outputs(3853)));
    outputs(942) <= (layer4_outputs(7562)) xor (layer4_outputs(2388));
    outputs(943) <= layer4_outputs(3278);
    outputs(944) <= not(layer4_outputs(761));
    outputs(945) <= layer4_outputs(4027);
    outputs(946) <= (layer4_outputs(8615)) xor (layer4_outputs(6770));
    outputs(947) <= (layer4_outputs(3401)) and (layer4_outputs(3838));
    outputs(948) <= not(layer4_outputs(4163));
    outputs(949) <= layer4_outputs(4420);
    outputs(950) <= not(layer4_outputs(1497));
    outputs(951) <= layer4_outputs(4366);
    outputs(952) <= not(layer4_outputs(122));
    outputs(953) <= not(layer4_outputs(3235));
    outputs(954) <= not(layer4_outputs(3556));
    outputs(955) <= not(layer4_outputs(7390));
    outputs(956) <= not(layer4_outputs(9703));
    outputs(957) <= not(layer4_outputs(8655));
    outputs(958) <= layer4_outputs(1373);
    outputs(959) <= not(layer4_outputs(2879));
    outputs(960) <= layer4_outputs(8067);
    outputs(961) <= layer4_outputs(7841);
    outputs(962) <= not((layer4_outputs(5869)) and (layer4_outputs(6592)));
    outputs(963) <= layer4_outputs(3944);
    outputs(964) <= layer4_outputs(5033);
    outputs(965) <= not(layer4_outputs(7514));
    outputs(966) <= (layer4_outputs(6720)) and not (layer4_outputs(7767));
    outputs(967) <= not(layer4_outputs(3468));
    outputs(968) <= not(layer4_outputs(7789));
    outputs(969) <= layer4_outputs(7147);
    outputs(970) <= not(layer4_outputs(7657));
    outputs(971) <= layer4_outputs(4806);
    outputs(972) <= layer4_outputs(4722);
    outputs(973) <= not(layer4_outputs(8587));
    outputs(974) <= layer4_outputs(4679);
    outputs(975) <= not(layer4_outputs(3452));
    outputs(976) <= not(layer4_outputs(9939));
    outputs(977) <= not((layer4_outputs(6978)) xor (layer4_outputs(2591)));
    outputs(978) <= (layer4_outputs(6371)) xor (layer4_outputs(5409));
    outputs(979) <= not(layer4_outputs(8409)) or (layer4_outputs(9460));
    outputs(980) <= layer4_outputs(6513);
    outputs(981) <= not(layer4_outputs(681));
    outputs(982) <= layer4_outputs(4441);
    outputs(983) <= not(layer4_outputs(5118));
    outputs(984) <= (layer4_outputs(8573)) xor (layer4_outputs(8135));
    outputs(985) <= not(layer4_outputs(7233));
    outputs(986) <= not((layer4_outputs(7796)) xor (layer4_outputs(9053)));
    outputs(987) <= not(layer4_outputs(2686));
    outputs(988) <= (layer4_outputs(9635)) or (layer4_outputs(5041));
    outputs(989) <= not((layer4_outputs(10013)) xor (layer4_outputs(8634)));
    outputs(990) <= not(layer4_outputs(7748));
    outputs(991) <= not(layer4_outputs(4504));
    outputs(992) <= not(layer4_outputs(3112));
    outputs(993) <= not(layer4_outputs(368));
    outputs(994) <= layer4_outputs(9480);
    outputs(995) <= not(layer4_outputs(7034));
    outputs(996) <= not(layer4_outputs(2313)) or (layer4_outputs(7199));
    outputs(997) <= (layer4_outputs(3130)) xor (layer4_outputs(3467));
    outputs(998) <= layer4_outputs(5111);
    outputs(999) <= not(layer4_outputs(3279));
    outputs(1000) <= not(layer4_outputs(5817));
    outputs(1001) <= not((layer4_outputs(3146)) and (layer4_outputs(3283)));
    outputs(1002) <= not((layer4_outputs(10225)) xor (layer4_outputs(6013)));
    outputs(1003) <= not(layer4_outputs(1697));
    outputs(1004) <= layer4_outputs(8514);
    outputs(1005) <= not(layer4_outputs(5844));
    outputs(1006) <= not(layer4_outputs(4231));
    outputs(1007) <= layer4_outputs(2798);
    outputs(1008) <= layer4_outputs(3392);
    outputs(1009) <= not(layer4_outputs(9017));
    outputs(1010) <= (layer4_outputs(6435)) and not (layer4_outputs(829));
    outputs(1011) <= (layer4_outputs(2034)) and not (layer4_outputs(3053));
    outputs(1012) <= not((layer4_outputs(2963)) xor (layer4_outputs(2304)));
    outputs(1013) <= not(layer4_outputs(2873));
    outputs(1014) <= not(layer4_outputs(1465));
    outputs(1015) <= layer4_outputs(5031);
    outputs(1016) <= layer4_outputs(932);
    outputs(1017) <= (layer4_outputs(3985)) or (layer4_outputs(9115));
    outputs(1018) <= not(layer4_outputs(2836));
    outputs(1019) <= not(layer4_outputs(3262)) or (layer4_outputs(691));
    outputs(1020) <= not(layer4_outputs(3802));
    outputs(1021) <= not((layer4_outputs(2064)) xor (layer4_outputs(1319)));
    outputs(1022) <= not(layer4_outputs(9556));
    outputs(1023) <= not((layer4_outputs(9923)) xor (layer4_outputs(1045)));
    outputs(1024) <= not(layer4_outputs(7300));
    outputs(1025) <= not(layer4_outputs(3749));
    outputs(1026) <= not(layer4_outputs(6931));
    outputs(1027) <= not(layer4_outputs(2094));
    outputs(1028) <= layer4_outputs(8568);
    outputs(1029) <= not((layer4_outputs(5890)) xor (layer4_outputs(6545)));
    outputs(1030) <= not(layer4_outputs(8762));
    outputs(1031) <= not(layer4_outputs(4613));
    outputs(1032) <= (layer4_outputs(446)) and (layer4_outputs(607));
    outputs(1033) <= not(layer4_outputs(8406));
    outputs(1034) <= layer4_outputs(1040);
    outputs(1035) <= not(layer4_outputs(402)) or (layer4_outputs(1510));
    outputs(1036) <= (layer4_outputs(50)) or (layer4_outputs(2306));
    outputs(1037) <= not(layer4_outputs(309));
    outputs(1038) <= layer4_outputs(8012);
    outputs(1039) <= layer4_outputs(5064);
    outputs(1040) <= layer4_outputs(685);
    outputs(1041) <= not((layer4_outputs(3830)) xor (layer4_outputs(9772)));
    outputs(1042) <= (layer4_outputs(1085)) and not (layer4_outputs(3106));
    outputs(1043) <= layer4_outputs(7223);
    outputs(1044) <= not(layer4_outputs(9506));
    outputs(1045) <= layer4_outputs(2091);
    outputs(1046) <= layer4_outputs(4487);
    outputs(1047) <= (layer4_outputs(7440)) xor (layer4_outputs(9454));
    outputs(1048) <= not(layer4_outputs(7817));
    outputs(1049) <= not((layer4_outputs(10221)) xor (layer4_outputs(4696)));
    outputs(1050) <= not((layer4_outputs(10120)) or (layer4_outputs(4479)));
    outputs(1051) <= (layer4_outputs(1344)) xor (layer4_outputs(5987));
    outputs(1052) <= layer4_outputs(1868);
    outputs(1053) <= not(layer4_outputs(9539));
    outputs(1054) <= '0';
    outputs(1055) <= not(layer4_outputs(6036)) or (layer4_outputs(2142));
    outputs(1056) <= not(layer4_outputs(5675));
    outputs(1057) <= not(layer4_outputs(6923));
    outputs(1058) <= not(layer4_outputs(10128));
    outputs(1059) <= layer4_outputs(4287);
    outputs(1060) <= layer4_outputs(1564);
    outputs(1061) <= not(layer4_outputs(9634));
    outputs(1062) <= layer4_outputs(8812);
    outputs(1063) <= layer4_outputs(4454);
    outputs(1064) <= (layer4_outputs(4403)) and not (layer4_outputs(4227));
    outputs(1065) <= not((layer4_outputs(4734)) xor (layer4_outputs(4882)));
    outputs(1066) <= not(layer4_outputs(1603));
    outputs(1067) <= (layer4_outputs(8150)) and not (layer4_outputs(3168));
    outputs(1068) <= not(layer4_outputs(2452)) or (layer4_outputs(3135));
    outputs(1069) <= not((layer4_outputs(9996)) or (layer4_outputs(5810)));
    outputs(1070) <= not(layer4_outputs(904));
    outputs(1071) <= layer4_outputs(5271);
    outputs(1072) <= layer4_outputs(5300);
    outputs(1073) <= layer4_outputs(10207);
    outputs(1074) <= layer4_outputs(3180);
    outputs(1075) <= not(layer4_outputs(2756));
    outputs(1076) <= (layer4_outputs(2475)) and (layer4_outputs(5615));
    outputs(1077) <= not((layer4_outputs(391)) xor (layer4_outputs(3242)));
    outputs(1078) <= not(layer4_outputs(9938));
    outputs(1079) <= not(layer4_outputs(1762));
    outputs(1080) <= (layer4_outputs(4338)) xor (layer4_outputs(6058));
    outputs(1081) <= layer4_outputs(2449);
    outputs(1082) <= layer4_outputs(4083);
    outputs(1083) <= not(layer4_outputs(4015)) or (layer4_outputs(7901));
    outputs(1084) <= (layer4_outputs(3388)) xor (layer4_outputs(7216));
    outputs(1085) <= (layer4_outputs(8130)) and not (layer4_outputs(9513));
    outputs(1086) <= (layer4_outputs(7082)) xor (layer4_outputs(4476));
    outputs(1087) <= layer4_outputs(6124);
    outputs(1088) <= not(layer4_outputs(202));
    outputs(1089) <= not(layer4_outputs(1853));
    outputs(1090) <= not(layer4_outputs(5709));
    outputs(1091) <= not((layer4_outputs(4625)) or (layer4_outputs(3738)));
    outputs(1092) <= layer4_outputs(5036);
    outputs(1093) <= not((layer4_outputs(3109)) xor (layer4_outputs(3491)));
    outputs(1094) <= (layer4_outputs(5587)) xor (layer4_outputs(6077));
    outputs(1095) <= layer4_outputs(106);
    outputs(1096) <= (layer4_outputs(2582)) and not (layer4_outputs(7977));
    outputs(1097) <= not(layer4_outputs(1435));
    outputs(1098) <= not(layer4_outputs(7726));
    outputs(1099) <= not(layer4_outputs(4293));
    outputs(1100) <= (layer4_outputs(2161)) and not (layer4_outputs(4197));
    outputs(1101) <= (layer4_outputs(7228)) and not (layer4_outputs(6421));
    outputs(1102) <= not((layer4_outputs(8874)) or (layer4_outputs(8717)));
    outputs(1103) <= not(layer4_outputs(7260));
    outputs(1104) <= not(layer4_outputs(4728));
    outputs(1105) <= (layer4_outputs(3884)) xor (layer4_outputs(662));
    outputs(1106) <= (layer4_outputs(464)) xor (layer4_outputs(8307));
    outputs(1107) <= (layer4_outputs(828)) xor (layer4_outputs(7036));
    outputs(1108) <= not(layer4_outputs(5262));
    outputs(1109) <= not((layer4_outputs(7377)) or (layer4_outputs(9510)));
    outputs(1110) <= (layer4_outputs(9715)) xor (layer4_outputs(1080));
    outputs(1111) <= layer4_outputs(4436);
    outputs(1112) <= not(layer4_outputs(2978));
    outputs(1113) <= (layer4_outputs(4787)) xor (layer4_outputs(5230));
    outputs(1114) <= (layer4_outputs(8618)) and not (layer4_outputs(2639));
    outputs(1115) <= (layer4_outputs(9508)) and not (layer4_outputs(960));
    outputs(1116) <= (layer4_outputs(6920)) and not (layer4_outputs(6107));
    outputs(1117) <= layer4_outputs(4207);
    outputs(1118) <= not(layer4_outputs(167));
    outputs(1119) <= layer4_outputs(303);
    outputs(1120) <= (layer4_outputs(6634)) and not (layer4_outputs(2134));
    outputs(1121) <= (layer4_outputs(2689)) and (layer4_outputs(8731));
    outputs(1122) <= not(layer4_outputs(5228));
    outputs(1123) <= not(layer4_outputs(9125));
    outputs(1124) <= (layer4_outputs(7835)) and not (layer4_outputs(6758));
    outputs(1125) <= not(layer4_outputs(6964));
    outputs(1126) <= (layer4_outputs(2482)) and (layer4_outputs(5818));
    outputs(1127) <= (layer4_outputs(4043)) and not (layer4_outputs(6204));
    outputs(1128) <= (layer4_outputs(1436)) and not (layer4_outputs(9313));
    outputs(1129) <= not((layer4_outputs(10046)) xor (layer4_outputs(5704)));
    outputs(1130) <= not(layer4_outputs(3541));
    outputs(1131) <= not(layer4_outputs(2877));
    outputs(1132) <= not(layer4_outputs(141));
    outputs(1133) <= not(layer4_outputs(7475));
    outputs(1134) <= not(layer4_outputs(6631));
    outputs(1135) <= layer4_outputs(9131);
    outputs(1136) <= not(layer4_outputs(6704));
    outputs(1137) <= not(layer4_outputs(5372));
    outputs(1138) <= layer4_outputs(3323);
    outputs(1139) <= layer4_outputs(9894);
    outputs(1140) <= layer4_outputs(4747);
    outputs(1141) <= (layer4_outputs(8109)) xor (layer4_outputs(4270));
    outputs(1142) <= not(layer4_outputs(2235));
    outputs(1143) <= layer4_outputs(8924);
    outputs(1144) <= (layer4_outputs(9837)) xor (layer4_outputs(317));
    outputs(1145) <= (layer4_outputs(8024)) and not (layer4_outputs(4681));
    outputs(1146) <= (layer4_outputs(2550)) xor (layer4_outputs(1154));
    outputs(1147) <= (layer4_outputs(4010)) and not (layer4_outputs(7253));
    outputs(1148) <= (layer4_outputs(7191)) and not (layer4_outputs(1616));
    outputs(1149) <= layer4_outputs(6811);
    outputs(1150) <= not(layer4_outputs(5504));
    outputs(1151) <= not((layer4_outputs(7422)) xor (layer4_outputs(4259)));
    outputs(1152) <= layer4_outputs(1757);
    outputs(1153) <= layer4_outputs(4332);
    outputs(1154) <= (layer4_outputs(7272)) xor (layer4_outputs(6913));
    outputs(1155) <= layer4_outputs(9602);
    outputs(1156) <= layer4_outputs(1457);
    outputs(1157) <= not(layer4_outputs(6075));
    outputs(1158) <= not(layer4_outputs(9106)) or (layer4_outputs(7656));
    outputs(1159) <= not((layer4_outputs(8064)) xor (layer4_outputs(4753)));
    outputs(1160) <= not(layer4_outputs(3925));
    outputs(1161) <= (layer4_outputs(9045)) and (layer4_outputs(6062));
    outputs(1162) <= layer4_outputs(2556);
    outputs(1163) <= not(layer4_outputs(1009));
    outputs(1164) <= (layer4_outputs(8521)) and not (layer4_outputs(6172));
    outputs(1165) <= not(layer4_outputs(5025));
    outputs(1166) <= not(layer4_outputs(4034));
    outputs(1167) <= layer4_outputs(1775);
    outputs(1168) <= not(layer4_outputs(5736));
    outputs(1169) <= (layer4_outputs(8508)) xor (layer4_outputs(7635));
    outputs(1170) <= not(layer4_outputs(4246));
    outputs(1171) <= layer4_outputs(844);
    outputs(1172) <= layer4_outputs(3677);
    outputs(1173) <= (layer4_outputs(1137)) xor (layer4_outputs(3686));
    outputs(1174) <= (layer4_outputs(9333)) xor (layer4_outputs(7762));
    outputs(1175) <= (layer4_outputs(4917)) xor (layer4_outputs(6043));
    outputs(1176) <= layer4_outputs(8056);
    outputs(1177) <= not(layer4_outputs(2406));
    outputs(1178) <= layer4_outputs(5624);
    outputs(1179) <= not(layer4_outputs(9847));
    outputs(1180) <= (layer4_outputs(4573)) and not (layer4_outputs(4863));
    outputs(1181) <= (layer4_outputs(545)) xor (layer4_outputs(4463));
    outputs(1182) <= layer4_outputs(1081);
    outputs(1183) <= not(layer4_outputs(4240));
    outputs(1184) <= (layer4_outputs(8854)) xor (layer4_outputs(9203));
    outputs(1185) <= not(layer4_outputs(10227));
    outputs(1186) <= (layer4_outputs(7924)) xor (layer4_outputs(5198));
    outputs(1187) <= layer4_outputs(1455);
    outputs(1188) <= not(layer4_outputs(380));
    outputs(1189) <= '1';
    outputs(1190) <= (layer4_outputs(5759)) and (layer4_outputs(1021));
    outputs(1191) <= (layer4_outputs(3860)) and not (layer4_outputs(10093));
    outputs(1192) <= not(layer4_outputs(6375));
    outputs(1193) <= (layer4_outputs(8677)) xor (layer4_outputs(2784));
    outputs(1194) <= not((layer4_outputs(531)) or (layer4_outputs(5298)));
    outputs(1195) <= layer4_outputs(2348);
    outputs(1196) <= (layer4_outputs(1858)) and not (layer4_outputs(6493));
    outputs(1197) <= '0';
    outputs(1198) <= (layer4_outputs(7509)) and (layer4_outputs(7389));
    outputs(1199) <= not(layer4_outputs(32));
    outputs(1200) <= layer4_outputs(8998);
    outputs(1201) <= layer4_outputs(8123);
    outputs(1202) <= (layer4_outputs(7013)) xor (layer4_outputs(718));
    outputs(1203) <= not(layer4_outputs(7321)) or (layer4_outputs(1358));
    outputs(1204) <= (layer4_outputs(1881)) and not (layer4_outputs(2154));
    outputs(1205) <= layer4_outputs(6478);
    outputs(1206) <= (layer4_outputs(4837)) and (layer4_outputs(5760));
    outputs(1207) <= not(layer4_outputs(406));
    outputs(1208) <= not(layer4_outputs(5863));
    outputs(1209) <= layer4_outputs(1707);
    outputs(1210) <= not(layer4_outputs(2298));
    outputs(1211) <= not((layer4_outputs(4014)) or (layer4_outputs(8416)));
    outputs(1212) <= (layer4_outputs(4656)) xor (layer4_outputs(7105));
    outputs(1213) <= not(layer4_outputs(7907));
    outputs(1214) <= layer4_outputs(2017);
    outputs(1215) <= not(layer4_outputs(7318));
    outputs(1216) <= not(layer4_outputs(7248));
    outputs(1217) <= not(layer4_outputs(8710));
    outputs(1218) <= not(layer4_outputs(226));
    outputs(1219) <= layer4_outputs(651);
    outputs(1220) <= not(layer4_outputs(481));
    outputs(1221) <= not((layer4_outputs(7886)) xor (layer4_outputs(9546)));
    outputs(1222) <= layer4_outputs(1614);
    outputs(1223) <= not((layer4_outputs(2094)) or (layer4_outputs(6368)));
    outputs(1224) <= (layer4_outputs(112)) and not (layer4_outputs(6001));
    outputs(1225) <= not((layer4_outputs(2572)) or (layer4_outputs(3104)));
    outputs(1226) <= layer4_outputs(10149);
    outputs(1227) <= (layer4_outputs(1886)) and not (layer4_outputs(88));
    outputs(1228) <= (layer4_outputs(3099)) or (layer4_outputs(3569));
    outputs(1229) <= layer4_outputs(3985);
    outputs(1230) <= layer4_outputs(9679);
    outputs(1231) <= (layer4_outputs(3181)) xor (layer4_outputs(3717));
    outputs(1232) <= layer4_outputs(2626);
    outputs(1233) <= not(layer4_outputs(1857));
    outputs(1234) <= not(layer4_outputs(2078));
    outputs(1235) <= not((layer4_outputs(1262)) or (layer4_outputs(1903)));
    outputs(1236) <= (layer4_outputs(4229)) xor (layer4_outputs(873));
    outputs(1237) <= not((layer4_outputs(510)) xor (layer4_outputs(7011)));
    outputs(1238) <= (layer4_outputs(6489)) xor (layer4_outputs(9465));
    outputs(1239) <= layer4_outputs(4168);
    outputs(1240) <= not((layer4_outputs(3484)) xor (layer4_outputs(1491)));
    outputs(1241) <= not(layer4_outputs(9909));
    outputs(1242) <= '0';
    outputs(1243) <= (layer4_outputs(2690)) xor (layer4_outputs(2874));
    outputs(1244) <= not(layer4_outputs(1220));
    outputs(1245) <= layer4_outputs(6382);
    outputs(1246) <= (layer4_outputs(5639)) xor (layer4_outputs(9138));
    outputs(1247) <= not(layer4_outputs(9996));
    outputs(1248) <= layer4_outputs(5553);
    outputs(1249) <= (layer4_outputs(529)) xor (layer4_outputs(3266));
    outputs(1250) <= layer4_outputs(7993);
    outputs(1251) <= layer4_outputs(3886);
    outputs(1252) <= (layer4_outputs(8658)) xor (layer4_outputs(3221));
    outputs(1253) <= (layer4_outputs(5596)) xor (layer4_outputs(2179));
    outputs(1254) <= (layer4_outputs(4113)) and not (layer4_outputs(5364));
    outputs(1255) <= (layer4_outputs(9933)) or (layer4_outputs(3250));
    outputs(1256) <= not((layer4_outputs(82)) xor (layer4_outputs(5305)));
    outputs(1257) <= not((layer4_outputs(5579)) or (layer4_outputs(4822)));
    outputs(1258) <= '0';
    outputs(1259) <= (layer4_outputs(1450)) and (layer4_outputs(2163));
    outputs(1260) <= (layer4_outputs(9019)) and (layer4_outputs(10076));
    outputs(1261) <= layer4_outputs(1174);
    outputs(1262) <= (layer4_outputs(7645)) and (layer4_outputs(5240));
    outputs(1263) <= not(layer4_outputs(9489));
    outputs(1264) <= (layer4_outputs(7283)) xor (layer4_outputs(8567));
    outputs(1265) <= not(layer4_outputs(2857));
    outputs(1266) <= not((layer4_outputs(8238)) xor (layer4_outputs(114)));
    outputs(1267) <= layer4_outputs(5955);
    outputs(1268) <= layer4_outputs(9144);
    outputs(1269) <= (layer4_outputs(9152)) xor (layer4_outputs(6869));
    outputs(1270) <= not(layer4_outputs(7071));
    outputs(1271) <= (layer4_outputs(4459)) and not (layer4_outputs(4461));
    outputs(1272) <= layer4_outputs(2153);
    outputs(1273) <= not((layer4_outputs(7807)) or (layer4_outputs(1637)));
    outputs(1274) <= (layer4_outputs(3748)) xor (layer4_outputs(7163));
    outputs(1275) <= not(layer4_outputs(8750));
    outputs(1276) <= not((layer4_outputs(8915)) xor (layer4_outputs(10218)));
    outputs(1277) <= (layer4_outputs(4623)) xor (layer4_outputs(117));
    outputs(1278) <= not(layer4_outputs(8479));
    outputs(1279) <= not((layer4_outputs(3149)) xor (layer4_outputs(2905)));
    outputs(1280) <= (layer4_outputs(2732)) xor (layer4_outputs(4645));
    outputs(1281) <= (layer4_outputs(4368)) xor (layer4_outputs(2792));
    outputs(1282) <= not(layer4_outputs(1192));
    outputs(1283) <= (layer4_outputs(2837)) and not (layer4_outputs(6897));
    outputs(1284) <= not(layer4_outputs(696));
    outputs(1285) <= (layer4_outputs(9574)) and not (layer4_outputs(855));
    outputs(1286) <= not(layer4_outputs(1811));
    outputs(1287) <= not(layer4_outputs(6778));
    outputs(1288) <= not(layer4_outputs(301));
    outputs(1289) <= layer4_outputs(4737);
    outputs(1290) <= (layer4_outputs(209)) and not (layer4_outputs(9571));
    outputs(1291) <= not(layer4_outputs(534));
    outputs(1292) <= not((layer4_outputs(5910)) or (layer4_outputs(8040)));
    outputs(1293) <= layer4_outputs(284);
    outputs(1294) <= layer4_outputs(9611);
    outputs(1295) <= (layer4_outputs(8275)) xor (layer4_outputs(8175));
    outputs(1296) <= not((layer4_outputs(9943)) xor (layer4_outputs(2112)));
    outputs(1297) <= (layer4_outputs(7826)) xor (layer4_outputs(3693));
    outputs(1298) <= (layer4_outputs(6065)) xor (layer4_outputs(145));
    outputs(1299) <= layer4_outputs(8792);
    outputs(1300) <= not(layer4_outputs(210));
    outputs(1301) <= (layer4_outputs(5987)) and not (layer4_outputs(5218));
    outputs(1302) <= (layer4_outputs(2088)) xor (layer4_outputs(488));
    outputs(1303) <= layer4_outputs(1511);
    outputs(1304) <= (layer4_outputs(1064)) xor (layer4_outputs(7357));
    outputs(1305) <= not(layer4_outputs(1293));
    outputs(1306) <= not((layer4_outputs(7045)) xor (layer4_outputs(6106)));
    outputs(1307) <= not((layer4_outputs(1261)) xor (layer4_outputs(8572)));
    outputs(1308) <= not(layer4_outputs(9149));
    outputs(1309) <= not(layer4_outputs(9832));
    outputs(1310) <= not(layer4_outputs(2929));
    outputs(1311) <= layer4_outputs(3333);
    outputs(1312) <= not(layer4_outputs(8810));
    outputs(1313) <= (layer4_outputs(4)) xor (layer4_outputs(3503));
    outputs(1314) <= not((layer4_outputs(6871)) or (layer4_outputs(7555)));
    outputs(1315) <= (layer4_outputs(3346)) and (layer4_outputs(6292));
    outputs(1316) <= (layer4_outputs(7592)) and not (layer4_outputs(3947));
    outputs(1317) <= not(layer4_outputs(327));
    outputs(1318) <= layer4_outputs(9517);
    outputs(1319) <= layer4_outputs(7205);
    outputs(1320) <= (layer4_outputs(6444)) or (layer4_outputs(6129));
    outputs(1321) <= (layer4_outputs(4939)) and not (layer4_outputs(8789));
    outputs(1322) <= layer4_outputs(7795);
    outputs(1323) <= (layer4_outputs(6391)) xor (layer4_outputs(9313));
    outputs(1324) <= not((layer4_outputs(8368)) xor (layer4_outputs(8229)));
    outputs(1325) <= not(layer4_outputs(362));
    outputs(1326) <= (layer4_outputs(3247)) xor (layer4_outputs(9438));
    outputs(1327) <= (layer4_outputs(8388)) and (layer4_outputs(8210));
    outputs(1328) <= layer4_outputs(601);
    outputs(1329) <= layer4_outputs(9369);
    outputs(1330) <= (layer4_outputs(8045)) xor (layer4_outputs(6639));
    outputs(1331) <= not(layer4_outputs(1589));
    outputs(1332) <= layer4_outputs(680);
    outputs(1333) <= layer4_outputs(9751);
    outputs(1334) <= (layer4_outputs(6332)) or (layer4_outputs(1278));
    outputs(1335) <= not(layer4_outputs(7754));
    outputs(1336) <= (layer4_outputs(5737)) and not (layer4_outputs(610));
    outputs(1337) <= (layer4_outputs(6136)) and not (layer4_outputs(7254));
    outputs(1338) <= (layer4_outputs(3495)) and (layer4_outputs(326));
    outputs(1339) <= not((layer4_outputs(2530)) xor (layer4_outputs(8826)));
    outputs(1340) <= not((layer4_outputs(1112)) xor (layer4_outputs(3790)));
    outputs(1341) <= layer4_outputs(5005);
    outputs(1342) <= layer4_outputs(5246);
    outputs(1343) <= (layer4_outputs(5537)) xor (layer4_outputs(8670));
    outputs(1344) <= (layer4_outputs(9891)) and not (layer4_outputs(6218));
    outputs(1345) <= layer4_outputs(7931);
    outputs(1346) <= not((layer4_outputs(2768)) xor (layer4_outputs(7586)));
    outputs(1347) <= (layer4_outputs(8526)) xor (layer4_outputs(8347));
    outputs(1348) <= not(layer4_outputs(4973));
    outputs(1349) <= (layer4_outputs(9995)) and not (layer4_outputs(5612));
    outputs(1350) <= (layer4_outputs(7922)) xor (layer4_outputs(9803));
    outputs(1351) <= not(layer4_outputs(4682));
    outputs(1352) <= layer4_outputs(9003);
    outputs(1353) <= '0';
    outputs(1354) <= not(layer4_outputs(4909));
    outputs(1355) <= layer4_outputs(8551);
    outputs(1356) <= (layer4_outputs(4579)) and (layer4_outputs(7685));
    outputs(1357) <= (layer4_outputs(5401)) xor (layer4_outputs(2193));
    outputs(1358) <= not((layer4_outputs(814)) xor (layer4_outputs(5231)));
    outputs(1359) <= layer4_outputs(6797);
    outputs(1360) <= not((layer4_outputs(10027)) or (layer4_outputs(5509)));
    outputs(1361) <= not((layer4_outputs(6653)) or (layer4_outputs(8534)));
    outputs(1362) <= not(layer4_outputs(4718));
    outputs(1363) <= (layer4_outputs(4278)) and not (layer4_outputs(2615));
    outputs(1364) <= layer4_outputs(8904);
    outputs(1365) <= not((layer4_outputs(7652)) or (layer4_outputs(1530)));
    outputs(1366) <= not(layer4_outputs(8576));
    outputs(1367) <= not(layer4_outputs(5589));
    outputs(1368) <= (layer4_outputs(313)) and (layer4_outputs(5438));
    outputs(1369) <= not(layer4_outputs(1172));
    outputs(1370) <= layer4_outputs(150);
    outputs(1371) <= (layer4_outputs(6476)) and not (layer4_outputs(6879));
    outputs(1372) <= not(layer4_outputs(4795));
    outputs(1373) <= not((layer4_outputs(4441)) xor (layer4_outputs(4986)));
    outputs(1374) <= not(layer4_outputs(1034));
    outputs(1375) <= (layer4_outputs(3303)) and not (layer4_outputs(683));
    outputs(1376) <= (layer4_outputs(1970)) and not (layer4_outputs(794));
    outputs(1377) <= not((layer4_outputs(2554)) xor (layer4_outputs(7535)));
    outputs(1378) <= not(layer4_outputs(8084));
    outputs(1379) <= (layer4_outputs(121)) xor (layer4_outputs(8898));
    outputs(1380) <= (layer4_outputs(738)) and not (layer4_outputs(4340));
    outputs(1381) <= layer4_outputs(2277);
    outputs(1382) <= not(layer4_outputs(10066));
    outputs(1383) <= layer4_outputs(4736);
    outputs(1384) <= layer4_outputs(7978);
    outputs(1385) <= not(layer4_outputs(5817));
    outputs(1386) <= not(layer4_outputs(10181));
    outputs(1387) <= not(layer4_outputs(3996));
    outputs(1388) <= not(layer4_outputs(8481));
    outputs(1389) <= not((layer4_outputs(2159)) xor (layer4_outputs(515)));
    outputs(1390) <= layer4_outputs(9827);
    outputs(1391) <= (layer4_outputs(1722)) and not (layer4_outputs(5779));
    outputs(1392) <= not(layer4_outputs(7608));
    outputs(1393) <= not(layer4_outputs(7755));
    outputs(1394) <= not(layer4_outputs(9366));
    outputs(1395) <= layer4_outputs(4193);
    outputs(1396) <= not(layer4_outputs(2569));
    outputs(1397) <= (layer4_outputs(7434)) xor (layer4_outputs(336));
    outputs(1398) <= not(layer4_outputs(6003));
    outputs(1399) <= not(layer4_outputs(9967)) or (layer4_outputs(6323));
    outputs(1400) <= layer4_outputs(2430);
    outputs(1401) <= not(layer4_outputs(2815));
    outputs(1402) <= '0';
    outputs(1403) <= (layer4_outputs(8250)) and not (layer4_outputs(2696));
    outputs(1404) <= (layer4_outputs(2553)) xor (layer4_outputs(3570));
    outputs(1405) <= not((layer4_outputs(6449)) or (layer4_outputs(4617)));
    outputs(1406) <= not(layer4_outputs(3979));
    outputs(1407) <= not(layer4_outputs(4881));
    outputs(1408) <= (layer4_outputs(2861)) xor (layer4_outputs(8694));
    outputs(1409) <= layer4_outputs(6455);
    outputs(1410) <= not((layer4_outputs(5449)) or (layer4_outputs(493)));
    outputs(1411) <= not(layer4_outputs(4066)) or (layer4_outputs(950));
    outputs(1412) <= layer4_outputs(564);
    outputs(1413) <= layer4_outputs(9556);
    outputs(1414) <= (layer4_outputs(5774)) and not (layer4_outputs(7711));
    outputs(1415) <= layer4_outputs(8942);
    outputs(1416) <= layer4_outputs(1340);
    outputs(1417) <= not((layer4_outputs(4435)) or (layer4_outputs(486)));
    outputs(1418) <= not((layer4_outputs(7729)) or (layer4_outputs(8113)));
    outputs(1419) <= not(layer4_outputs(223));
    outputs(1420) <= (layer4_outputs(3747)) and not (layer4_outputs(5272));
    outputs(1421) <= not((layer4_outputs(7097)) or (layer4_outputs(8933)));
    outputs(1422) <= not(layer4_outputs(8195));
    outputs(1423) <= not((layer4_outputs(9590)) xor (layer4_outputs(1231)));
    outputs(1424) <= '0';
    outputs(1425) <= not((layer4_outputs(1268)) xor (layer4_outputs(5352)));
    outputs(1426) <= not((layer4_outputs(6869)) xor (layer4_outputs(4644)));
    outputs(1427) <= layer4_outputs(2711);
    outputs(1428) <= layer4_outputs(3835);
    outputs(1429) <= not(layer4_outputs(2315));
    outputs(1430) <= (layer4_outputs(1453)) and (layer4_outputs(5628));
    outputs(1431) <= layer4_outputs(4607);
    outputs(1432) <= not((layer4_outputs(2284)) or (layer4_outputs(5918)));
    outputs(1433) <= (layer4_outputs(9157)) and (layer4_outputs(5238));
    outputs(1434) <= (layer4_outputs(4579)) xor (layer4_outputs(4012));
    outputs(1435) <= layer4_outputs(8856);
    outputs(1436) <= layer4_outputs(4589);
    outputs(1437) <= not(layer4_outputs(4189));
    outputs(1438) <= not(layer4_outputs(10227)) or (layer4_outputs(8594));
    outputs(1439) <= not((layer4_outputs(2314)) xor (layer4_outputs(1149)));
    outputs(1440) <= not(layer4_outputs(8740));
    outputs(1441) <= not((layer4_outputs(7385)) xor (layer4_outputs(7761)));
    outputs(1442) <= layer4_outputs(3681);
    outputs(1443) <= layer4_outputs(5931);
    outputs(1444) <= not(layer4_outputs(5201));
    outputs(1445) <= not(layer4_outputs(8142));
    outputs(1446) <= layer4_outputs(6451);
    outputs(1447) <= not((layer4_outputs(981)) xor (layer4_outputs(4594)));
    outputs(1448) <= layer4_outputs(761);
    outputs(1449) <= not(layer4_outputs(9502));
    outputs(1450) <= not(layer4_outputs(8416));
    outputs(1451) <= layer4_outputs(6200);
    outputs(1452) <= not((layer4_outputs(2083)) xor (layer4_outputs(7894)));
    outputs(1453) <= not((layer4_outputs(6033)) xor (layer4_outputs(7070)));
    outputs(1454) <= (layer4_outputs(3735)) xor (layer4_outputs(682));
    outputs(1455) <= (layer4_outputs(5816)) xor (layer4_outputs(7005));
    outputs(1456) <= (layer4_outputs(7576)) and (layer4_outputs(2803));
    outputs(1457) <= layer4_outputs(5681);
    outputs(1458) <= (layer4_outputs(6656)) xor (layer4_outputs(9807));
    outputs(1459) <= (layer4_outputs(5764)) xor (layer4_outputs(5696));
    outputs(1460) <= layer4_outputs(8722);
    outputs(1461) <= not(layer4_outputs(9762));
    outputs(1462) <= not((layer4_outputs(8623)) or (layer4_outputs(4119)));
    outputs(1463) <= not(layer4_outputs(3801));
    outputs(1464) <= (layer4_outputs(8279)) and not (layer4_outputs(8293));
    outputs(1465) <= (layer4_outputs(5038)) xor (layer4_outputs(9794));
    outputs(1466) <= layer4_outputs(3436);
    outputs(1467) <= (layer4_outputs(9157)) and not (layer4_outputs(2703));
    outputs(1468) <= not(layer4_outputs(7331));
    outputs(1469) <= not(layer4_outputs(4090));
    outputs(1470) <= (layer4_outputs(197)) and (layer4_outputs(3155));
    outputs(1471) <= layer4_outputs(7881);
    outputs(1472) <= not(layer4_outputs(4156));
    outputs(1473) <= not(layer4_outputs(782));
    outputs(1474) <= (layer4_outputs(8086)) and not (layer4_outputs(1339));
    outputs(1475) <= not((layer4_outputs(367)) xor (layer4_outputs(2098)));
    outputs(1476) <= not(layer4_outputs(4575));
    outputs(1477) <= not(layer4_outputs(8330));
    outputs(1478) <= not(layer4_outputs(6345));
    outputs(1479) <= not(layer4_outputs(3544));
    outputs(1480) <= layer4_outputs(7450);
    outputs(1481) <= not((layer4_outputs(9795)) or (layer4_outputs(3663)));
    outputs(1482) <= not((layer4_outputs(5962)) xor (layer4_outputs(1524)));
    outputs(1483) <= not(layer4_outputs(7432));
    outputs(1484) <= (layer4_outputs(1511)) and not (layer4_outputs(923));
    outputs(1485) <= layer4_outputs(4372);
    outputs(1486) <= not(layer4_outputs(2885));
    outputs(1487) <= (layer4_outputs(1007)) and not (layer4_outputs(9680));
    outputs(1488) <= not(layer4_outputs(7695));
    outputs(1489) <= not(layer4_outputs(8079));
    outputs(1490) <= layer4_outputs(8540);
    outputs(1491) <= (layer4_outputs(6381)) and not (layer4_outputs(9930));
    outputs(1492) <= not(layer4_outputs(3306));
    outputs(1493) <= (layer4_outputs(1994)) xor (layer4_outputs(1397));
    outputs(1494) <= (layer4_outputs(7344)) and not (layer4_outputs(2369));
    outputs(1495) <= not(layer4_outputs(696));
    outputs(1496) <= layer4_outputs(2244);
    outputs(1497) <= not(layer4_outputs(6757));
    outputs(1498) <= layer4_outputs(7576);
    outputs(1499) <= layer4_outputs(10052);
    outputs(1500) <= (layer4_outputs(6678)) and not (layer4_outputs(2825));
    outputs(1501) <= (layer4_outputs(7742)) and not (layer4_outputs(6422));
    outputs(1502) <= not(layer4_outputs(3001));
    outputs(1503) <= (layer4_outputs(10006)) and (layer4_outputs(3413));
    outputs(1504) <= layer4_outputs(105);
    outputs(1505) <= not(layer4_outputs(3841));
    outputs(1506) <= (layer4_outputs(9890)) and not (layer4_outputs(8421));
    outputs(1507) <= not(layer4_outputs(8115));
    outputs(1508) <= layer4_outputs(8631);
    outputs(1509) <= (layer4_outputs(4547)) xor (layer4_outputs(4845));
    outputs(1510) <= (layer4_outputs(5719)) and not (layer4_outputs(1675));
    outputs(1511) <= not(layer4_outputs(692)) or (layer4_outputs(4063));
    outputs(1512) <= not(layer4_outputs(4494));
    outputs(1513) <= not(layer4_outputs(4874));
    outputs(1514) <= layer4_outputs(4429);
    outputs(1515) <= layer4_outputs(1442);
    outputs(1516) <= (layer4_outputs(9698)) and (layer4_outputs(9929));
    outputs(1517) <= (layer4_outputs(10163)) and not (layer4_outputs(2421));
    outputs(1518) <= (layer4_outputs(5362)) and not (layer4_outputs(3229));
    outputs(1519) <= not(layer4_outputs(7207));
    outputs(1520) <= not(layer4_outputs(5837));
    outputs(1521) <= layer4_outputs(4582);
    outputs(1522) <= (layer4_outputs(8593)) and not (layer4_outputs(2713));
    outputs(1523) <= not(layer4_outputs(6875));
    outputs(1524) <= not(layer4_outputs(3591));
    outputs(1525) <= (layer4_outputs(2432)) xor (layer4_outputs(8376));
    outputs(1526) <= layer4_outputs(5620);
    outputs(1527) <= not(layer4_outputs(5939));
    outputs(1528) <= not((layer4_outputs(6426)) xor (layer4_outputs(4416)));
    outputs(1529) <= layer4_outputs(7206);
    outputs(1530) <= (layer4_outputs(3198)) and not (layer4_outputs(4989));
    outputs(1531) <= not(layer4_outputs(3439));
    outputs(1532) <= layer4_outputs(2776);
    outputs(1533) <= (layer4_outputs(6527)) and not (layer4_outputs(5876));
    outputs(1534) <= (layer4_outputs(5043)) xor (layer4_outputs(194));
    outputs(1535) <= not((layer4_outputs(9734)) or (layer4_outputs(99)));
    outputs(1536) <= not((layer4_outputs(9386)) or (layer4_outputs(10187)));
    outputs(1537) <= (layer4_outputs(7680)) or (layer4_outputs(5861));
    outputs(1538) <= layer4_outputs(3856);
    outputs(1539) <= not(layer4_outputs(3360));
    outputs(1540) <= not(layer4_outputs(8205));
    outputs(1541) <= not((layer4_outputs(10075)) or (layer4_outputs(3038)));
    outputs(1542) <= layer4_outputs(6914);
    outputs(1543) <= layer4_outputs(6151);
    outputs(1544) <= (layer4_outputs(1713)) xor (layer4_outputs(3431));
    outputs(1545) <= not(layer4_outputs(2621));
    outputs(1546) <= not(layer4_outputs(5370));
    outputs(1547) <= not(layer4_outputs(2392)) or (layer4_outputs(699));
    outputs(1548) <= not(layer4_outputs(7055));
    outputs(1549) <= (layer4_outputs(9138)) xor (layer4_outputs(6915));
    outputs(1550) <= not((layer4_outputs(7731)) xor (layer4_outputs(6742)));
    outputs(1551) <= not(layer4_outputs(2954));
    outputs(1552) <= (layer4_outputs(3782)) and not (layer4_outputs(451));
    outputs(1553) <= not((layer4_outputs(8904)) xor (layer4_outputs(4703)));
    outputs(1554) <= not(layer4_outputs(183));
    outputs(1555) <= layer4_outputs(6609);
    outputs(1556) <= (layer4_outputs(61)) and not (layer4_outputs(10237));
    outputs(1557) <= not(layer4_outputs(5365));
    outputs(1558) <= layer4_outputs(4149);
    outputs(1559) <= not((layer4_outputs(6089)) or (layer4_outputs(417)));
    outputs(1560) <= not((layer4_outputs(3251)) xor (layer4_outputs(6015)));
    outputs(1561) <= (layer4_outputs(1671)) xor (layer4_outputs(4250));
    outputs(1562) <= not(layer4_outputs(5885));
    outputs(1563) <= not(layer4_outputs(5807));
    outputs(1564) <= layer4_outputs(5963);
    outputs(1565) <= not(layer4_outputs(994));
    outputs(1566) <= layer4_outputs(2294);
    outputs(1567) <= not((layer4_outputs(1286)) xor (layer4_outputs(1764)));
    outputs(1568) <= (layer4_outputs(3128)) xor (layer4_outputs(6174));
    outputs(1569) <= not(layer4_outputs(3541));
    outputs(1570) <= not(layer4_outputs(2199));
    outputs(1571) <= not(layer4_outputs(5801));
    outputs(1572) <= not(layer4_outputs(618));
    outputs(1573) <= not((layer4_outputs(7809)) xor (layer4_outputs(5416)));
    outputs(1574) <= (layer4_outputs(290)) xor (layer4_outputs(3192));
    outputs(1575) <= not(layer4_outputs(891));
    outputs(1576) <= (layer4_outputs(2962)) xor (layer4_outputs(6160));
    outputs(1577) <= not(layer4_outputs(2151));
    outputs(1578) <= not(layer4_outputs(5529));
    outputs(1579) <= not(layer4_outputs(3892));
    outputs(1580) <= not(layer4_outputs(8680));
    outputs(1581) <= (layer4_outputs(1083)) and (layer4_outputs(6968));
    outputs(1582) <= not((layer4_outputs(7029)) xor (layer4_outputs(506)));
    outputs(1583) <= (layer4_outputs(8637)) xor (layer4_outputs(3162));
    outputs(1584) <= (layer4_outputs(6814)) and not (layer4_outputs(9098));
    outputs(1585) <= not(layer4_outputs(2831));
    outputs(1586) <= (layer4_outputs(5348)) and (layer4_outputs(6601));
    outputs(1587) <= (layer4_outputs(9839)) xor (layer4_outputs(8105));
    outputs(1588) <= not((layer4_outputs(1451)) xor (layer4_outputs(3678)));
    outputs(1589) <= not(layer4_outputs(2133));
    outputs(1590) <= not(layer4_outputs(6274));
    outputs(1591) <= not(layer4_outputs(9538));
    outputs(1592) <= not(layer4_outputs(3568));
    outputs(1593) <= (layer4_outputs(4421)) and not (layer4_outputs(6178));
    outputs(1594) <= not((layer4_outputs(2819)) or (layer4_outputs(897)));
    outputs(1595) <= layer4_outputs(8517);
    outputs(1596) <= (layer4_outputs(7040)) and not (layer4_outputs(4504));
    outputs(1597) <= layer4_outputs(5034);
    outputs(1598) <= not((layer4_outputs(2189)) or (layer4_outputs(9678)));
    outputs(1599) <= layer4_outputs(3097);
    outputs(1600) <= layer4_outputs(2058);
    outputs(1601) <= (layer4_outputs(945)) xor (layer4_outputs(4098));
    outputs(1602) <= layer4_outputs(980);
    outputs(1603) <= not((layer4_outputs(507)) or (layer4_outputs(3021)));
    outputs(1604) <= layer4_outputs(2484);
    outputs(1605) <= (layer4_outputs(970)) and not (layer4_outputs(491));
    outputs(1606) <= not((layer4_outputs(4936)) or (layer4_outputs(2087)));
    outputs(1607) <= (layer4_outputs(82)) and not (layer4_outputs(8009));
    outputs(1608) <= (layer4_outputs(6868)) and not (layer4_outputs(2654));
    outputs(1609) <= (layer4_outputs(1934)) xor (layer4_outputs(9383));
    outputs(1610) <= not(layer4_outputs(3200));
    outputs(1611) <= not(layer4_outputs(4930));
    outputs(1612) <= (layer4_outputs(9262)) xor (layer4_outputs(1051));
    outputs(1613) <= (layer4_outputs(7842)) and (layer4_outputs(1847));
    outputs(1614) <= not(layer4_outputs(4171));
    outputs(1615) <= not(layer4_outputs(6121));
    outputs(1616) <= layer4_outputs(5408);
    outputs(1617) <= not(layer4_outputs(6412));
    outputs(1618) <= not(layer4_outputs(2569));
    outputs(1619) <= not(layer4_outputs(7618));
    outputs(1620) <= layer4_outputs(3703);
    outputs(1621) <= (layer4_outputs(8655)) and not (layer4_outputs(4515));
    outputs(1622) <= not(layer4_outputs(1335));
    outputs(1623) <= not(layer4_outputs(5661));
    outputs(1624) <= not(layer4_outputs(4727));
    outputs(1625) <= layer4_outputs(5601);
    outputs(1626) <= layer4_outputs(3436);
    outputs(1627) <= layer4_outputs(3603);
    outputs(1628) <= (layer4_outputs(6263)) and not (layer4_outputs(2625));
    outputs(1629) <= (layer4_outputs(1977)) and (layer4_outputs(9315));
    outputs(1630) <= (layer4_outputs(9279)) and not (layer4_outputs(2548));
    outputs(1631) <= layer4_outputs(9765);
    outputs(1632) <= layer4_outputs(8776);
    outputs(1633) <= layer4_outputs(2307);
    outputs(1634) <= not((layer4_outputs(7853)) xor (layer4_outputs(1547)));
    outputs(1635) <= layer4_outputs(5354);
    outputs(1636) <= not(layer4_outputs(2380));
    outputs(1637) <= not(layer4_outputs(5258));
    outputs(1638) <= layer4_outputs(9371);
    outputs(1639) <= layer4_outputs(8773);
    outputs(1640) <= not((layer4_outputs(814)) xor (layer4_outputs(7664)));
    outputs(1641) <= layer4_outputs(7637);
    outputs(1642) <= (layer4_outputs(2370)) xor (layer4_outputs(7454));
    outputs(1643) <= (layer4_outputs(1015)) xor (layer4_outputs(587));
    outputs(1644) <= layer4_outputs(2879);
    outputs(1645) <= (layer4_outputs(3241)) and not (layer4_outputs(5368));
    outputs(1646) <= (layer4_outputs(9006)) xor (layer4_outputs(2390));
    outputs(1647) <= layer4_outputs(8307);
    outputs(1648) <= layer4_outputs(1296);
    outputs(1649) <= not((layer4_outputs(1627)) xor (layer4_outputs(836)));
    outputs(1650) <= not(layer4_outputs(5223));
    outputs(1651) <= not((layer4_outputs(693)) xor (layer4_outputs(8703)));
    outputs(1652) <= not((layer4_outputs(4913)) xor (layer4_outputs(309)));
    outputs(1653) <= layer4_outputs(2035);
    outputs(1654) <= not(layer4_outputs(3700));
    outputs(1655) <= (layer4_outputs(6735)) and not (layer4_outputs(952));
    outputs(1656) <= not(layer4_outputs(4053)) or (layer4_outputs(9784));
    outputs(1657) <= not(layer4_outputs(8822));
    outputs(1658) <= not(layer4_outputs(83));
    outputs(1659) <= layer4_outputs(601);
    outputs(1660) <= layer4_outputs(3601);
    outputs(1661) <= layer4_outputs(3310);
    outputs(1662) <= (layer4_outputs(1838)) and (layer4_outputs(3561));
    outputs(1663) <= (layer4_outputs(3584)) and not (layer4_outputs(7501));
    outputs(1664) <= (layer4_outputs(7472)) and not (layer4_outputs(148));
    outputs(1665) <= layer4_outputs(7590);
    outputs(1666) <= (layer4_outputs(4964)) xor (layer4_outputs(5990));
    outputs(1667) <= not(layer4_outputs(7226));
    outputs(1668) <= (layer4_outputs(2801)) and not (layer4_outputs(1282));
    outputs(1669) <= not(layer4_outputs(3563));
    outputs(1670) <= layer4_outputs(4394);
    outputs(1671) <= layer4_outputs(4023);
    outputs(1672) <= not(layer4_outputs(1454));
    outputs(1673) <= layer4_outputs(4612);
    outputs(1674) <= layer4_outputs(7673);
    outputs(1675) <= not(layer4_outputs(5025));
    outputs(1676) <= (layer4_outputs(8712)) xor (layer4_outputs(9084));
    outputs(1677) <= not(layer4_outputs(4171));
    outputs(1678) <= (layer4_outputs(797)) and not (layer4_outputs(70));
    outputs(1679) <= (layer4_outputs(6728)) and (layer4_outputs(9647));
    outputs(1680) <= not(layer4_outputs(6189));
    outputs(1681) <= (layer4_outputs(5035)) and (layer4_outputs(6656));
    outputs(1682) <= not(layer4_outputs(6754));
    outputs(1683) <= (layer4_outputs(5090)) and not (layer4_outputs(2355));
    outputs(1684) <= (layer4_outputs(2095)) and not (layer4_outputs(2399));
    outputs(1685) <= (layer4_outputs(3640)) and not (layer4_outputs(4971));
    outputs(1686) <= '0';
    outputs(1687) <= not(layer4_outputs(7729));
    outputs(1688) <= not(layer4_outputs(5412));
    outputs(1689) <= (layer4_outputs(2283)) and not (layer4_outputs(5370));
    outputs(1690) <= layer4_outputs(9062);
    outputs(1691) <= (layer4_outputs(7883)) and not (layer4_outputs(9695));
    outputs(1692) <= layer4_outputs(3476);
    outputs(1693) <= not(layer4_outputs(9487));
    outputs(1694) <= not(layer4_outputs(5367));
    outputs(1695) <= not(layer4_outputs(265)) or (layer4_outputs(2319));
    outputs(1696) <= layer4_outputs(9915);
    outputs(1697) <= (layer4_outputs(3724)) and (layer4_outputs(10004));
    outputs(1698) <= layer4_outputs(7908);
    outputs(1699) <= (layer4_outputs(9167)) or (layer4_outputs(8357));
    outputs(1700) <= (layer4_outputs(2870)) xor (layer4_outputs(4817));
    outputs(1701) <= not(layer4_outputs(361));
    outputs(1702) <= not(layer4_outputs(412));
    outputs(1703) <= not(layer4_outputs(4762));
    outputs(1704) <= not(layer4_outputs(7235));
    outputs(1705) <= not(layer4_outputs(5504));
    outputs(1706) <= layer4_outputs(1081);
    outputs(1707) <= not(layer4_outputs(7433));
    outputs(1708) <= layer4_outputs(5016);
    outputs(1709) <= not(layer4_outputs(946));
    outputs(1710) <= (layer4_outputs(6914)) and not (layer4_outputs(110));
    outputs(1711) <= not(layer4_outputs(1888));
    outputs(1712) <= (layer4_outputs(5646)) and not (layer4_outputs(6744));
    outputs(1713) <= not((layer4_outputs(7676)) and (layer4_outputs(816)));
    outputs(1714) <= not((layer4_outputs(1515)) xor (layer4_outputs(2434)));
    outputs(1715) <= not((layer4_outputs(8888)) xor (layer4_outputs(1447)));
    outputs(1716) <= not(layer4_outputs(2241));
    outputs(1717) <= layer4_outputs(1916);
    outputs(1718) <= layer4_outputs(3863);
    outputs(1719) <= (layer4_outputs(4319)) and not (layer4_outputs(5096));
    outputs(1720) <= not((layer4_outputs(3934)) or (layer4_outputs(1566)));
    outputs(1721) <= layer4_outputs(9570);
    outputs(1722) <= not((layer4_outputs(9169)) xor (layer4_outputs(9201)));
    outputs(1723) <= not((layer4_outputs(5217)) xor (layer4_outputs(2619)));
    outputs(1724) <= layer4_outputs(6072);
    outputs(1725) <= not(layer4_outputs(175));
    outputs(1726) <= not(layer4_outputs(7427));
    outputs(1727) <= (layer4_outputs(7478)) and (layer4_outputs(6771));
    outputs(1728) <= (layer4_outputs(7545)) and not (layer4_outputs(8598));
    outputs(1729) <= (layer4_outputs(8722)) and (layer4_outputs(2287));
    outputs(1730) <= not((layer4_outputs(4353)) or (layer4_outputs(5280)));
    outputs(1731) <= not(layer4_outputs(3264));
    outputs(1732) <= layer4_outputs(4586);
    outputs(1733) <= layer4_outputs(9421);
    outputs(1734) <= (layer4_outputs(75)) and not (layer4_outputs(9950));
    outputs(1735) <= (layer4_outputs(7846)) and (layer4_outputs(8837));
    outputs(1736) <= not(layer4_outputs(5630));
    outputs(1737) <= (layer4_outputs(8392)) and not (layer4_outputs(2996));
    outputs(1738) <= layer4_outputs(4393);
    outputs(1739) <= (layer4_outputs(4259)) and (layer4_outputs(3407));
    outputs(1740) <= not(layer4_outputs(3184));
    outputs(1741) <= layer4_outputs(1090);
    outputs(1742) <= not(layer4_outputs(2584));
    outputs(1743) <= not(layer4_outputs(2316));
    outputs(1744) <= not((layer4_outputs(10168)) or (layer4_outputs(9921)));
    outputs(1745) <= (layer4_outputs(4040)) and (layer4_outputs(786));
    outputs(1746) <= not(layer4_outputs(8286));
    outputs(1747) <= (layer4_outputs(4319)) and not (layer4_outputs(4560));
    outputs(1748) <= (layer4_outputs(2069)) and not (layer4_outputs(2736));
    outputs(1749) <= (layer4_outputs(4887)) and (layer4_outputs(7064));
    outputs(1750) <= (layer4_outputs(2459)) and (layer4_outputs(2549));
    outputs(1751) <= not(layer4_outputs(6141));
    outputs(1752) <= layer4_outputs(5935);
    outputs(1753) <= layer4_outputs(2359);
    outputs(1754) <= not(layer4_outputs(6600));
    outputs(1755) <= not((layer4_outputs(5391)) xor (layer4_outputs(539)));
    outputs(1756) <= layer4_outputs(953);
    outputs(1757) <= layer4_outputs(3618);
    outputs(1758) <= layer4_outputs(5377);
    outputs(1759) <= not(layer4_outputs(5396));
    outputs(1760) <= not((layer4_outputs(9156)) xor (layer4_outputs(5146)));
    outputs(1761) <= not(layer4_outputs(9310));
    outputs(1762) <= layer4_outputs(742);
    outputs(1763) <= not((layer4_outputs(6985)) xor (layer4_outputs(3441)));
    outputs(1764) <= layer4_outputs(6682);
    outputs(1765) <= (layer4_outputs(3010)) xor (layer4_outputs(6803));
    outputs(1766) <= not(layer4_outputs(10025));
    outputs(1767) <= not(layer4_outputs(8578));
    outputs(1768) <= not(layer4_outputs(9244));
    outputs(1769) <= (layer4_outputs(5103)) xor (layer4_outputs(421));
    outputs(1770) <= not(layer4_outputs(3183));
    outputs(1771) <= not(layer4_outputs(7230));
    outputs(1772) <= (layer4_outputs(5750)) and not (layer4_outputs(3255));
    outputs(1773) <= layer4_outputs(7099);
    outputs(1774) <= not(layer4_outputs(65));
    outputs(1775) <= (layer4_outputs(2697)) and not (layer4_outputs(9061));
    outputs(1776) <= not(layer4_outputs(6924));
    outputs(1777) <= (layer4_outputs(4052)) xor (layer4_outputs(4148));
    outputs(1778) <= (layer4_outputs(4726)) and not (layer4_outputs(7336));
    outputs(1779) <= not(layer4_outputs(8249));
    outputs(1780) <= not(layer4_outputs(7285));
    outputs(1781) <= not(layer4_outputs(9241));
    outputs(1782) <= (layer4_outputs(4006)) xor (layer4_outputs(2942));
    outputs(1783) <= not(layer4_outputs(8301));
    outputs(1784) <= not(layer4_outputs(8146));
    outputs(1785) <= '0';
    outputs(1786) <= (layer4_outputs(4435)) xor (layer4_outputs(2662));
    outputs(1787) <= not(layer4_outputs(3332));
    outputs(1788) <= (layer4_outputs(700)) and not (layer4_outputs(1532));
    outputs(1789) <= layer4_outputs(6959);
    outputs(1790) <= (layer4_outputs(7993)) and not (layer4_outputs(9776));
    outputs(1791) <= not(layer4_outputs(2488));
    outputs(1792) <= (layer4_outputs(2923)) xor (layer4_outputs(992));
    outputs(1793) <= not(layer4_outputs(263));
    outputs(1794) <= not(layer4_outputs(785));
    outputs(1795) <= (layer4_outputs(6529)) xor (layer4_outputs(511));
    outputs(1796) <= not(layer4_outputs(10146));
    outputs(1797) <= layer4_outputs(7863);
    outputs(1798) <= layer4_outputs(1580);
    outputs(1799) <= (layer4_outputs(7829)) and not (layer4_outputs(8177));
    outputs(1800) <= not((layer4_outputs(8531)) xor (layer4_outputs(9759)));
    outputs(1801) <= layer4_outputs(8336);
    outputs(1802) <= layer4_outputs(546);
    outputs(1803) <= not(layer4_outputs(767));
    outputs(1804) <= not(layer4_outputs(6075));
    outputs(1805) <= not(layer4_outputs(4452));
    outputs(1806) <= layer4_outputs(8933);
    outputs(1807) <= layer4_outputs(1193);
    outputs(1808) <= layer4_outputs(1433);
    outputs(1809) <= not(layer4_outputs(8311));
    outputs(1810) <= (layer4_outputs(7119)) xor (layer4_outputs(793));
    outputs(1811) <= layer4_outputs(3724);
    outputs(1812) <= layer4_outputs(2046);
    outputs(1813) <= not((layer4_outputs(4287)) or (layer4_outputs(9531)));
    outputs(1814) <= (layer4_outputs(1259)) and not (layer4_outputs(8041));
    outputs(1815) <= (layer4_outputs(3360)) and not (layer4_outputs(1530));
    outputs(1816) <= (layer4_outputs(3870)) and (layer4_outputs(7952));
    outputs(1817) <= not(layer4_outputs(6345)) or (layer4_outputs(3144));
    outputs(1818) <= not(layer4_outputs(6687));
    outputs(1819) <= (layer4_outputs(3679)) xor (layer4_outputs(3542));
    outputs(1820) <= not(layer4_outputs(7413));
    outputs(1821) <= layer4_outputs(4415);
    outputs(1822) <= not(layer4_outputs(9538));
    outputs(1823) <= not((layer4_outputs(9473)) or (layer4_outputs(1609)));
    outputs(1824) <= (layer4_outputs(4405)) and (layer4_outputs(8059));
    outputs(1825) <= not((layer4_outputs(2824)) xor (layer4_outputs(5663)));
    outputs(1826) <= layer4_outputs(7117);
    outputs(1827) <= not(layer4_outputs(5971));
    outputs(1828) <= layer4_outputs(608);
    outputs(1829) <= (layer4_outputs(4082)) and not (layer4_outputs(2438));
    outputs(1830) <= not(layer4_outputs(7839));
    outputs(1831) <= layer4_outputs(1885);
    outputs(1832) <= not((layer4_outputs(1304)) xor (layer4_outputs(6748)));
    outputs(1833) <= not(layer4_outputs(1236));
    outputs(1834) <= not(layer4_outputs(6199));
    outputs(1835) <= not(layer4_outputs(9451));
    outputs(1836) <= layer4_outputs(4163);
    outputs(1837) <= not(layer4_outputs(97));
    outputs(1838) <= '0';
    outputs(1839) <= not((layer4_outputs(2100)) or (layer4_outputs(3130)));
    outputs(1840) <= (layer4_outputs(4460)) xor (layer4_outputs(9472));
    outputs(1841) <= layer4_outputs(9407);
    outputs(1842) <= (layer4_outputs(2906)) xor (layer4_outputs(499));
    outputs(1843) <= layer4_outputs(818);
    outputs(1844) <= layer4_outputs(3770);
    outputs(1845) <= not(layer4_outputs(801));
    outputs(1846) <= (layer4_outputs(2439)) and not (layer4_outputs(7093));
    outputs(1847) <= not(layer4_outputs(428));
    outputs(1848) <= not(layer4_outputs(7838));
    outputs(1849) <= not(layer4_outputs(9652));
    outputs(1850) <= layer4_outputs(7797);
    outputs(1851) <= layer4_outputs(3440);
    outputs(1852) <= (layer4_outputs(9293)) and not (layer4_outputs(8120));
    outputs(1853) <= not(layer4_outputs(1062));
    outputs(1854) <= not((layer4_outputs(1124)) or (layer4_outputs(4822)));
    outputs(1855) <= not(layer4_outputs(2890));
    outputs(1856) <= (layer4_outputs(2652)) and not (layer4_outputs(3756));
    outputs(1857) <= (layer4_outputs(8166)) and not (layer4_outputs(7733));
    outputs(1858) <= (layer4_outputs(9751)) and (layer4_outputs(3777));
    outputs(1859) <= layer4_outputs(8456);
    outputs(1860) <= (layer4_outputs(2342)) or (layer4_outputs(2188));
    outputs(1861) <= not((layer4_outputs(7367)) xor (layer4_outputs(1225)));
    outputs(1862) <= layer4_outputs(8240);
    outputs(1863) <= layer4_outputs(1960);
    outputs(1864) <= layer4_outputs(295);
    outputs(1865) <= (layer4_outputs(5896)) and (layer4_outputs(9550));
    outputs(1866) <= (layer4_outputs(9820)) and (layer4_outputs(1250));
    outputs(1867) <= (layer4_outputs(4460)) and not (layer4_outputs(5309));
    outputs(1868) <= (layer4_outputs(4199)) xor (layer4_outputs(10044));
    outputs(1869) <= (layer4_outputs(1801)) xor (layer4_outputs(6939));
    outputs(1870) <= layer4_outputs(8582);
    outputs(1871) <= not(layer4_outputs(7331));
    outputs(1872) <= not(layer4_outputs(5418));
    outputs(1873) <= layer4_outputs(965);
    outputs(1874) <= (layer4_outputs(1268)) and (layer4_outputs(4602));
    outputs(1875) <= layer4_outputs(2120);
    outputs(1876) <= not(layer4_outputs(3273));
    outputs(1877) <= layer4_outputs(8702);
    outputs(1878) <= layer4_outputs(9688);
    outputs(1879) <= (layer4_outputs(4390)) xor (layer4_outputs(5304));
    outputs(1880) <= (layer4_outputs(2183)) and (layer4_outputs(10162));
    outputs(1881) <= layer4_outputs(9968);
    outputs(1882) <= not(layer4_outputs(5098));
    outputs(1883) <= (layer4_outputs(267)) xor (layer4_outputs(2999));
    outputs(1884) <= not(layer4_outputs(9551));
    outputs(1885) <= not(layer4_outputs(6729));
    outputs(1886) <= (layer4_outputs(5105)) and not (layer4_outputs(8807));
    outputs(1887) <= not(layer4_outputs(8522));
    outputs(1888) <= layer4_outputs(6480);
    outputs(1889) <= layer4_outputs(578);
    outputs(1890) <= (layer4_outputs(7350)) and not (layer4_outputs(4608));
    outputs(1891) <= not(layer4_outputs(78)) or (layer4_outputs(6850));
    outputs(1892) <= layer4_outputs(3285);
    outputs(1893) <= layer4_outputs(1059);
    outputs(1894) <= (layer4_outputs(3119)) and not (layer4_outputs(375));
    outputs(1895) <= not(layer4_outputs(6252));
    outputs(1896) <= not((layer4_outputs(9559)) xor (layer4_outputs(9088)));
    outputs(1897) <= layer4_outputs(4002);
    outputs(1898) <= not(layer4_outputs(8176));
    outputs(1899) <= not(layer4_outputs(7300));
    outputs(1900) <= (layer4_outputs(10148)) and not (layer4_outputs(660));
    outputs(1901) <= layer4_outputs(1536);
    outputs(1902) <= not((layer4_outputs(8857)) xor (layer4_outputs(6450)));
    outputs(1903) <= not(layer4_outputs(6181));
    outputs(1904) <= not((layer4_outputs(1691)) or (layer4_outputs(785)));
    outputs(1905) <= not((layer4_outputs(1962)) xor (layer4_outputs(4562)));
    outputs(1906) <= (layer4_outputs(6331)) and (layer4_outputs(1178));
    outputs(1907) <= (layer4_outputs(8539)) or (layer4_outputs(9243));
    outputs(1908) <= (layer4_outputs(6870)) xor (layer4_outputs(905));
    outputs(1909) <= layer4_outputs(6890);
    outputs(1910) <= layer4_outputs(3820);
    outputs(1911) <= not((layer4_outputs(8467)) xor (layer4_outputs(6358)));
    outputs(1912) <= not(layer4_outputs(4550));
    outputs(1913) <= layer4_outputs(3898);
    outputs(1914) <= (layer4_outputs(5825)) and (layer4_outputs(754));
    outputs(1915) <= not(layer4_outputs(6110)) or (layer4_outputs(2983));
    outputs(1916) <= not(layer4_outputs(2915));
    outputs(1917) <= not((layer4_outputs(6836)) xor (layer4_outputs(8738)));
    outputs(1918) <= layer4_outputs(5163);
    outputs(1919) <= not((layer4_outputs(6070)) xor (layer4_outputs(8842)));
    outputs(1920) <= not(layer4_outputs(6949));
    outputs(1921) <= (layer4_outputs(8615)) xor (layer4_outputs(435));
    outputs(1922) <= not(layer4_outputs(64));
    outputs(1923) <= layer4_outputs(5947);
    outputs(1924) <= layer4_outputs(6739);
    outputs(1925) <= layer4_outputs(8796);
    outputs(1926) <= layer4_outputs(9475);
    outputs(1927) <= not((layer4_outputs(7473)) or (layer4_outputs(9590)));
    outputs(1928) <= not(layer4_outputs(4020));
    outputs(1929) <= not(layer4_outputs(1666));
    outputs(1930) <= (layer4_outputs(4495)) and not (layer4_outputs(7235));
    outputs(1931) <= not(layer4_outputs(8589));
    outputs(1932) <= not((layer4_outputs(2526)) or (layer4_outputs(3521)));
    outputs(1933) <= not((layer4_outputs(2390)) xor (layer4_outputs(5051)));
    outputs(1934) <= not(layer4_outputs(5373));
    outputs(1935) <= not((layer4_outputs(8177)) or (layer4_outputs(3212)));
    outputs(1936) <= not(layer4_outputs(3421));
    outputs(1937) <= layer4_outputs(2045);
    outputs(1938) <= layer4_outputs(4207);
    outputs(1939) <= (layer4_outputs(2038)) and (layer4_outputs(2595));
    outputs(1940) <= (layer4_outputs(2223)) and not (layer4_outputs(3390));
    outputs(1941) <= not(layer4_outputs(7655));
    outputs(1942) <= (layer4_outputs(3662)) xor (layer4_outputs(5030));
    outputs(1943) <= (layer4_outputs(6963)) xor (layer4_outputs(9602));
    outputs(1944) <= (layer4_outputs(3163)) xor (layer4_outputs(3688));
    outputs(1945) <= layer4_outputs(6506);
    outputs(1946) <= not(layer4_outputs(9323));
    outputs(1947) <= layer4_outputs(137);
    outputs(1948) <= layer4_outputs(2682);
    outputs(1949) <= not((layer4_outputs(9191)) xor (layer4_outputs(3797)));
    outputs(1950) <= not(layer4_outputs(10151));
    outputs(1951) <= layer4_outputs(6988);
    outputs(1952) <= not((layer4_outputs(7905)) xor (layer4_outputs(2613)));
    outputs(1953) <= not(layer4_outputs(315));
    outputs(1954) <= layer4_outputs(5040);
    outputs(1955) <= not(layer4_outputs(9746));
    outputs(1956) <= not((layer4_outputs(9705)) xor (layer4_outputs(4898)));
    outputs(1957) <= not(layer4_outputs(10023));
    outputs(1958) <= not(layer4_outputs(5152)) or (layer4_outputs(449));
    outputs(1959) <= not((layer4_outputs(59)) or (layer4_outputs(4877)));
    outputs(1960) <= not((layer4_outputs(3999)) or (layer4_outputs(1852)));
    outputs(1961) <= not(layer4_outputs(3024));
    outputs(1962) <= layer4_outputs(6746);
    outputs(1963) <= not(layer4_outputs(57));
    outputs(1964) <= not((layer4_outputs(4003)) xor (layer4_outputs(1719)));
    outputs(1965) <= not((layer4_outputs(8221)) xor (layer4_outputs(10233)));
    outputs(1966) <= not((layer4_outputs(5488)) or (layer4_outputs(6001)));
    outputs(1967) <= layer4_outputs(6093);
    outputs(1968) <= layer4_outputs(7626);
    outputs(1969) <= layer4_outputs(2281);
    outputs(1970) <= layer4_outputs(2114);
    outputs(1971) <= not(layer4_outputs(7726));
    outputs(1972) <= not(layer4_outputs(7021));
    outputs(1973) <= (layer4_outputs(9109)) and not (layer4_outputs(9474));
    outputs(1974) <= not((layer4_outputs(2180)) and (layer4_outputs(8195)));
    outputs(1975) <= (layer4_outputs(916)) and not (layer4_outputs(1507));
    outputs(1976) <= (layer4_outputs(4524)) xor (layer4_outputs(397));
    outputs(1977) <= (layer4_outputs(1203)) xor (layer4_outputs(2594));
    outputs(1978) <= not(layer4_outputs(1264));
    outputs(1979) <= layer4_outputs(9952);
    outputs(1980) <= (layer4_outputs(1095)) and (layer4_outputs(570));
    outputs(1981) <= not(layer4_outputs(311));
    outputs(1982) <= not(layer4_outputs(8795));
    outputs(1983) <= (layer4_outputs(9045)) and not (layer4_outputs(3722));
    outputs(1984) <= not(layer4_outputs(396));
    outputs(1985) <= layer4_outputs(9055);
    outputs(1986) <= not(layer4_outputs(4016));
    outputs(1987) <= not(layer4_outputs(6413));
    outputs(1988) <= (layer4_outputs(1337)) xor (layer4_outputs(3710));
    outputs(1989) <= not(layer4_outputs(4387)) or (layer4_outputs(2191));
    outputs(1990) <= layer4_outputs(2780);
    outputs(1991) <= not(layer4_outputs(3666));
    outputs(1992) <= not((layer4_outputs(8715)) xor (layer4_outputs(3104)));
    outputs(1993) <= not(layer4_outputs(9128));
    outputs(1994) <= not((layer4_outputs(2430)) xor (layer4_outputs(7406)));
    outputs(1995) <= not(layer4_outputs(1399));
    outputs(1996) <= layer4_outputs(1219);
    outputs(1997) <= (layer4_outputs(9092)) and (layer4_outputs(1263));
    outputs(1998) <= layer4_outputs(6027);
    outputs(1999) <= (layer4_outputs(3545)) and not (layer4_outputs(7258));
    outputs(2000) <= not(layer4_outputs(9442));
    outputs(2001) <= not(layer4_outputs(5373));
    outputs(2002) <= layer4_outputs(2433);
    outputs(2003) <= not(layer4_outputs(3050));
    outputs(2004) <= layer4_outputs(7127);
    outputs(2005) <= not(layer4_outputs(6904));
    outputs(2006) <= (layer4_outputs(4234)) and not (layer4_outputs(8882));
    outputs(2007) <= not(layer4_outputs(2924));
    outputs(2008) <= not((layer4_outputs(6026)) or (layer4_outputs(4925)));
    outputs(2009) <= layer4_outputs(4627);
    outputs(2010) <= layer4_outputs(2586);
    outputs(2011) <= not(layer4_outputs(5757));
    outputs(2012) <= (layer4_outputs(8865)) xor (layer4_outputs(3064));
    outputs(2013) <= (layer4_outputs(6353)) and (layer4_outputs(6347));
    outputs(2014) <= layer4_outputs(4086);
    outputs(2015) <= not(layer4_outputs(7006));
    outputs(2016) <= layer4_outputs(5604);
    outputs(2017) <= not(layer4_outputs(8917));
    outputs(2018) <= not((layer4_outputs(7975)) xor (layer4_outputs(7700)));
    outputs(2019) <= layer4_outputs(6562);
    outputs(2020) <= (layer4_outputs(2363)) and (layer4_outputs(7516));
    outputs(2021) <= layer4_outputs(9304);
    outputs(2022) <= layer4_outputs(2542);
    outputs(2023) <= not(layer4_outputs(9343));
    outputs(2024) <= not(layer4_outputs(9951));
    outputs(2025) <= not((layer4_outputs(5338)) xor (layer4_outputs(6512)));
    outputs(2026) <= not(layer4_outputs(5139));
    outputs(2027) <= not(layer4_outputs(2710));
    outputs(2028) <= (layer4_outputs(7697)) xor (layer4_outputs(7879));
    outputs(2029) <= layer4_outputs(351);
    outputs(2030) <= not(layer4_outputs(10128));
    outputs(2031) <= not(layer4_outputs(6185)) or (layer4_outputs(2017));
    outputs(2032) <= layer4_outputs(4697);
    outputs(2033) <= (layer4_outputs(8781)) and not (layer4_outputs(8332));
    outputs(2034) <= (layer4_outputs(8006)) and not (layer4_outputs(6793));
    outputs(2035) <= layer4_outputs(5009);
    outputs(2036) <= (layer4_outputs(1750)) xor (layer4_outputs(7460));
    outputs(2037) <= layer4_outputs(1915);
    outputs(2038) <= layer4_outputs(6462);
    outputs(2039) <= not(layer4_outputs(2187)) or (layer4_outputs(792));
    outputs(2040) <= (layer4_outputs(3972)) xor (layer4_outputs(8691));
    outputs(2041) <= layer4_outputs(3548);
    outputs(2042) <= not((layer4_outputs(8061)) or (layer4_outputs(8970)));
    outputs(2043) <= layer4_outputs(6444);
    outputs(2044) <= layer4_outputs(404);
    outputs(2045) <= not((layer4_outputs(5308)) xor (layer4_outputs(8131)));
    outputs(2046) <= not(layer4_outputs(25));
    outputs(2047) <= layer4_outputs(3304);
    outputs(2048) <= layer4_outputs(7600);
    outputs(2049) <= not((layer4_outputs(4663)) xor (layer4_outputs(688)));
    outputs(2050) <= not((layer4_outputs(5261)) xor (layer4_outputs(5570)));
    outputs(2051) <= not(layer4_outputs(2145));
    outputs(2052) <= not((layer4_outputs(8263)) xor (layer4_outputs(2577)));
    outputs(2053) <= layer4_outputs(3531);
    outputs(2054) <= (layer4_outputs(4508)) xor (layer4_outputs(8829));
    outputs(2055) <= not((layer4_outputs(9985)) xor (layer4_outputs(777)));
    outputs(2056) <= not((layer4_outputs(3836)) and (layer4_outputs(3854)));
    outputs(2057) <= not(layer4_outputs(3620));
    outputs(2058) <= layer4_outputs(5472);
    outputs(2059) <= layer4_outputs(8439);
    outputs(2060) <= not((layer4_outputs(7766)) xor (layer4_outputs(9275)));
    outputs(2061) <= not(layer4_outputs(6162));
    outputs(2062) <= layer4_outputs(1807);
    outputs(2063) <= (layer4_outputs(5215)) xor (layer4_outputs(371));
    outputs(2064) <= not(layer4_outputs(2851));
    outputs(2065) <= layer4_outputs(4802);
    outputs(2066) <= not(layer4_outputs(3513));
    outputs(2067) <= not(layer4_outputs(1872));
    outputs(2068) <= (layer4_outputs(4312)) xor (layer4_outputs(2829));
    outputs(2069) <= (layer4_outputs(10108)) xor (layer4_outputs(7254));
    outputs(2070) <= (layer4_outputs(6585)) and not (layer4_outputs(6844));
    outputs(2071) <= (layer4_outputs(811)) xor (layer4_outputs(9071));
    outputs(2072) <= (layer4_outputs(4284)) xor (layer4_outputs(10194));
    outputs(2073) <= not(layer4_outputs(4132));
    outputs(2074) <= not((layer4_outputs(9504)) xor (layer4_outputs(6730)));
    outputs(2075) <= not(layer4_outputs(953));
    outputs(2076) <= (layer4_outputs(3346)) and not (layer4_outputs(2830));
    outputs(2077) <= layer4_outputs(7232);
    outputs(2078) <= not((layer4_outputs(6558)) and (layer4_outputs(3344)));
    outputs(2079) <= not(layer4_outputs(9670));
    outputs(2080) <= (layer4_outputs(5858)) and not (layer4_outputs(6355));
    outputs(2081) <= not(layer4_outputs(425));
    outputs(2082) <= not(layer4_outputs(6471));
    outputs(2083) <= layer4_outputs(9944);
    outputs(2084) <= layer4_outputs(4140);
    outputs(2085) <= layer4_outputs(6611);
    outputs(2086) <= not(layer4_outputs(3134));
    outputs(2087) <= not(layer4_outputs(7041));
    outputs(2088) <= not(layer4_outputs(3312));
    outputs(2089) <= not(layer4_outputs(6231));
    outputs(2090) <= not(layer4_outputs(7957));
    outputs(2091) <= not((layer4_outputs(2542)) and (layer4_outputs(8731)));
    outputs(2092) <= not(layer4_outputs(4434));
    outputs(2093) <= (layer4_outputs(9205)) and not (layer4_outputs(4444));
    outputs(2094) <= not(layer4_outputs(8438));
    outputs(2095) <= not(layer4_outputs(3612));
    outputs(2096) <= not(layer4_outputs(2572));
    outputs(2097) <= not(layer4_outputs(6292));
    outputs(2098) <= '1';
    outputs(2099) <= layer4_outputs(8326);
    outputs(2100) <= layer4_outputs(7004);
    outputs(2101) <= not(layer4_outputs(5240));
    outputs(2102) <= not(layer4_outputs(1760));
    outputs(2103) <= not(layer4_outputs(4675)) or (layer4_outputs(635));
    outputs(2104) <= (layer4_outputs(1291)) and (layer4_outputs(8104));
    outputs(2105) <= not((layer4_outputs(1905)) and (layer4_outputs(2994)));
    outputs(2106) <= not(layer4_outputs(8239));
    outputs(2107) <= (layer4_outputs(4765)) xor (layer4_outputs(10091));
    outputs(2108) <= not(layer4_outputs(4596));
    outputs(2109) <= not(layer4_outputs(9728));
    outputs(2110) <= layer4_outputs(4354);
    outputs(2111) <= not(layer4_outputs(10179));
    outputs(2112) <= not(layer4_outputs(1351));
    outputs(2113) <= not(layer4_outputs(3712));
    outputs(2114) <= (layer4_outputs(8991)) xor (layer4_outputs(6264));
    outputs(2115) <= not(layer4_outputs(918));
    outputs(2116) <= layer4_outputs(7640);
    outputs(2117) <= not(layer4_outputs(9180)) or (layer4_outputs(991));
    outputs(2118) <= (layer4_outputs(1730)) or (layer4_outputs(949));
    outputs(2119) <= layer4_outputs(1153);
    outputs(2120) <= not((layer4_outputs(2810)) and (layer4_outputs(3358)));
    outputs(2121) <= not(layer4_outputs(3182));
    outputs(2122) <= not(layer4_outputs(2560)) or (layer4_outputs(5656));
    outputs(2123) <= layer4_outputs(6554);
    outputs(2124) <= not(layer4_outputs(9802)) or (layer4_outputs(6311));
    outputs(2125) <= layer4_outputs(3799);
    outputs(2126) <= (layer4_outputs(1002)) xor (layer4_outputs(337));
    outputs(2127) <= not(layer4_outputs(9816));
    outputs(2128) <= not(layer4_outputs(886));
    outputs(2129) <= not((layer4_outputs(8032)) or (layer4_outputs(5619)));
    outputs(2130) <= not((layer4_outputs(951)) xor (layer4_outputs(2791)));
    outputs(2131) <= not(layer4_outputs(6201));
    outputs(2132) <= not(layer4_outputs(2437));
    outputs(2133) <= layer4_outputs(2796);
    outputs(2134) <= not(layer4_outputs(9920));
    outputs(2135) <= not((layer4_outputs(716)) xor (layer4_outputs(3060)));
    outputs(2136) <= not(layer4_outputs(6462));
    outputs(2137) <= not(layer4_outputs(3879));
    outputs(2138) <= (layer4_outputs(1323)) or (layer4_outputs(567));
    outputs(2139) <= not(layer4_outputs(1244));
    outputs(2140) <= not(layer4_outputs(8772));
    outputs(2141) <= layer4_outputs(7510);
    outputs(2142) <= (layer4_outputs(4308)) xor (layer4_outputs(4645));
    outputs(2143) <= layer4_outputs(10062);
    outputs(2144) <= (layer4_outputs(2773)) xor (layer4_outputs(4272));
    outputs(2145) <= layer4_outputs(5583);
    outputs(2146) <= not(layer4_outputs(9347));
    outputs(2147) <= not(layer4_outputs(3843));
    outputs(2148) <= layer4_outputs(7364);
    outputs(2149) <= layer4_outputs(4415);
    outputs(2150) <= (layer4_outputs(8663)) and (layer4_outputs(8311));
    outputs(2151) <= not(layer4_outputs(7967));
    outputs(2152) <= layer4_outputs(5097);
    outputs(2153) <= not(layer4_outputs(3769));
    outputs(2154) <= not((layer4_outputs(4367)) xor (layer4_outputs(6281)));
    outputs(2155) <= (layer4_outputs(7648)) xor (layer4_outputs(839));
    outputs(2156) <= not(layer4_outputs(3658));
    outputs(2157) <= not((layer4_outputs(7219)) xor (layer4_outputs(1109)));
    outputs(2158) <= layer4_outputs(9196);
    outputs(2159) <= not(layer4_outputs(1274));
    outputs(2160) <= layer4_outputs(4552);
    outputs(2161) <= not(layer4_outputs(132));
    outputs(2162) <= layer4_outputs(4744);
    outputs(2163) <= not((layer4_outputs(986)) xor (layer4_outputs(1139)));
    outputs(2164) <= not(layer4_outputs(7900));
    outputs(2165) <= not(layer4_outputs(7221)) or (layer4_outputs(6188));
    outputs(2166) <= not(layer4_outputs(2676));
    outputs(2167) <= not((layer4_outputs(653)) xor (layer4_outputs(7898)));
    outputs(2168) <= layer4_outputs(8069);
    outputs(2169) <= not(layer4_outputs(6872));
    outputs(2170) <= not(layer4_outputs(5876));
    outputs(2171) <= not(layer4_outputs(5942));
    outputs(2172) <= layer4_outputs(2071);
    outputs(2173) <= layer4_outputs(930);
    outputs(2174) <= not(layer4_outputs(8883));
    outputs(2175) <= not((layer4_outputs(7648)) xor (layer4_outputs(9747)));
    outputs(2176) <= not(layer4_outputs(4086));
    outputs(2177) <= layer4_outputs(3736);
    outputs(2178) <= not((layer4_outputs(7337)) xor (layer4_outputs(9689)));
    outputs(2179) <= not(layer4_outputs(648)) or (layer4_outputs(6856));
    outputs(2180) <= not((layer4_outputs(6220)) or (layer4_outputs(2167)));
    outputs(2181) <= layer4_outputs(3477);
    outputs(2182) <= not(layer4_outputs(10047));
    outputs(2183) <= layer4_outputs(6633);
    outputs(2184) <= not(layer4_outputs(9661));
    outputs(2185) <= not(layer4_outputs(4481));
    outputs(2186) <= not(layer4_outputs(5706)) or (layer4_outputs(5242));
    outputs(2187) <= (layer4_outputs(5060)) xor (layer4_outputs(1155));
    outputs(2188) <= layer4_outputs(10220);
    outputs(2189) <= not(layer4_outputs(9135));
    outputs(2190) <= not(layer4_outputs(4509));
    outputs(2191) <= layer4_outputs(4468);
    outputs(2192) <= not(layer4_outputs(4105));
    outputs(2193) <= not(layer4_outputs(5605));
    outputs(2194) <= layer4_outputs(7880);
    outputs(2195) <= not(layer4_outputs(599));
    outputs(2196) <= not((layer4_outputs(147)) xor (layer4_outputs(2315)));
    outputs(2197) <= not(layer4_outputs(2120));
    outputs(2198) <= not(layer4_outputs(8118)) or (layer4_outputs(2730));
    outputs(2199) <= (layer4_outputs(8511)) xor (layer4_outputs(5922));
    outputs(2200) <= (layer4_outputs(3579)) xor (layer4_outputs(5583));
    outputs(2201) <= (layer4_outputs(3015)) and not (layer4_outputs(5648));
    outputs(2202) <= not((layer4_outputs(9351)) or (layer4_outputs(6363)));
    outputs(2203) <= layer4_outputs(342);
    outputs(2204) <= layer4_outputs(6299);
    outputs(2205) <= not(layer4_outputs(7479));
    outputs(2206) <= not((layer4_outputs(492)) or (layer4_outputs(6535)));
    outputs(2207) <= layer4_outputs(1635);
    outputs(2208) <= layer4_outputs(9257);
    outputs(2209) <= not(layer4_outputs(725)) or (layer4_outputs(563));
    outputs(2210) <= (layer4_outputs(3102)) xor (layer4_outputs(3321));
    outputs(2211) <= not(layer4_outputs(5685)) or (layer4_outputs(9503));
    outputs(2212) <= layer4_outputs(4847);
    outputs(2213) <= layer4_outputs(9825);
    outputs(2214) <= layer4_outputs(7275);
    outputs(2215) <= not(layer4_outputs(6078));
    outputs(2216) <= not(layer4_outputs(1140));
    outputs(2217) <= not(layer4_outputs(2056));
    outputs(2218) <= not(layer4_outputs(5446));
    outputs(2219) <= (layer4_outputs(7409)) and not (layer4_outputs(4546));
    outputs(2220) <= not((layer4_outputs(1252)) xor (layer4_outputs(929)));
    outputs(2221) <= not(layer4_outputs(4764));
    outputs(2222) <= not(layer4_outputs(2739));
    outputs(2223) <= not(layer4_outputs(9580)) or (layer4_outputs(9141));
    outputs(2224) <= not(layer4_outputs(9260));
    outputs(2225) <= not(layer4_outputs(6654));
    outputs(2226) <= layer4_outputs(2865);
    outputs(2227) <= layer4_outputs(8017);
    outputs(2228) <= layer4_outputs(5651);
    outputs(2229) <= not((layer4_outputs(1634)) xor (layer4_outputs(5163)));
    outputs(2230) <= layer4_outputs(325);
    outputs(2231) <= not(layer4_outputs(9114));
    outputs(2232) <= not((layer4_outputs(2019)) and (layer4_outputs(7198)));
    outputs(2233) <= not(layer4_outputs(8528));
    outputs(2234) <= not(layer4_outputs(3877)) or (layer4_outputs(1172));
    outputs(2235) <= layer4_outputs(8224);
    outputs(2236) <= not(layer4_outputs(4104));
    outputs(2237) <= not(layer4_outputs(9260));
    outputs(2238) <= layer4_outputs(3532);
    outputs(2239) <= not((layer4_outputs(9721)) xor (layer4_outputs(7489)));
    outputs(2240) <= not((layer4_outputs(5831)) xor (layer4_outputs(2132)));
    outputs(2241) <= not((layer4_outputs(1520)) xor (layer4_outputs(10152)));
    outputs(2242) <= layer4_outputs(8510);
    outputs(2243) <= not(layer4_outputs(3790));
    outputs(2244) <= (layer4_outputs(5758)) xor (layer4_outputs(2130));
    outputs(2245) <= not(layer4_outputs(782));
    outputs(2246) <= not(layer4_outputs(7025));
    outputs(2247) <= layer4_outputs(1505);
    outputs(2248) <= not(layer4_outputs(5177));
    outputs(2249) <= not(layer4_outputs(4035)) or (layer4_outputs(4963));
    outputs(2250) <= not(layer4_outputs(5748));
    outputs(2251) <= layer4_outputs(8953);
    outputs(2252) <= layer4_outputs(2418);
    outputs(2253) <= layer4_outputs(1545);
    outputs(2254) <= not((layer4_outputs(763)) xor (layer4_outputs(228)));
    outputs(2255) <= not((layer4_outputs(5726)) xor (layer4_outputs(9614)));
    outputs(2256) <= layer4_outputs(1347);
    outputs(2257) <= layer4_outputs(6953);
    outputs(2258) <= not(layer4_outputs(2133));
    outputs(2259) <= '0';
    outputs(2260) <= not(layer4_outputs(1560)) or (layer4_outputs(9422));
    outputs(2261) <= (layer4_outputs(6966)) or (layer4_outputs(4242));
    outputs(2262) <= not((layer4_outputs(6702)) or (layer4_outputs(2826)));
    outputs(2263) <= not(layer4_outputs(9417)) or (layer4_outputs(8870));
    outputs(2264) <= not(layer4_outputs(4101));
    outputs(2265) <= not((layer4_outputs(955)) xor (layer4_outputs(2131)));
    outputs(2266) <= layer4_outputs(4203);
    outputs(2267) <= layer4_outputs(2388);
    outputs(2268) <= layer4_outputs(1211);
    outputs(2269) <= (layer4_outputs(2865)) and (layer4_outputs(8959));
    outputs(2270) <= layer4_outputs(3113);
    outputs(2271) <= (layer4_outputs(5246)) or (layer4_outputs(2350));
    outputs(2272) <= (layer4_outputs(2215)) xor (layer4_outputs(2197));
    outputs(2273) <= not(layer4_outputs(396));
    outputs(2274) <= layer4_outputs(1374);
    outputs(2275) <= layer4_outputs(8050);
    outputs(2276) <= layer4_outputs(9764);
    outputs(2277) <= not(layer4_outputs(7574));
    outputs(2278) <= not(layer4_outputs(2988));
    outputs(2279) <= not(layer4_outputs(9291));
    outputs(2280) <= not((layer4_outputs(1860)) xor (layer4_outputs(1983)));
    outputs(2281) <= layer4_outputs(8706);
    outputs(2282) <= not(layer4_outputs(3017)) or (layer4_outputs(321));
    outputs(2283) <= layer4_outputs(1440);
    outputs(2284) <= not((layer4_outputs(6268)) xor (layer4_outputs(890)));
    outputs(2285) <= layer4_outputs(4914);
    outputs(2286) <= not(layer4_outputs(8909));
    outputs(2287) <= layer4_outputs(9829);
    outputs(2288) <= not(layer4_outputs(9114));
    outputs(2289) <= not((layer4_outputs(8699)) or (layer4_outputs(5308)));
    outputs(2290) <= (layer4_outputs(6846)) xor (layer4_outputs(4555));
    outputs(2291) <= not(layer4_outputs(6493));
    outputs(2292) <= layer4_outputs(4553);
    outputs(2293) <= layer4_outputs(1189);
    outputs(2294) <= not((layer4_outputs(5116)) or (layer4_outputs(9150)));
    outputs(2295) <= layer4_outputs(7873);
    outputs(2296) <= not((layer4_outputs(2593)) or (layer4_outputs(2610)));
    outputs(2297) <= layer4_outputs(7426);
    outputs(2298) <= not(layer4_outputs(8105));
    outputs(2299) <= not(layer4_outputs(5423));
    outputs(2300) <= layer4_outputs(1472);
    outputs(2301) <= (layer4_outputs(9341)) xor (layer4_outputs(6669));
    outputs(2302) <= not(layer4_outputs(5837));
    outputs(2303) <= not(layer4_outputs(9248));
    outputs(2304) <= not((layer4_outputs(10215)) xor (layer4_outputs(2900)));
    outputs(2305) <= layer4_outputs(8868);
    outputs(2306) <= not((layer4_outputs(1208)) xor (layer4_outputs(2678)));
    outputs(2307) <= (layer4_outputs(6925)) xor (layer4_outputs(6924));
    outputs(2308) <= layer4_outputs(1983);
    outputs(2309) <= (layer4_outputs(5858)) xor (layer4_outputs(7008));
    outputs(2310) <= layer4_outputs(3995);
    outputs(2311) <= layer4_outputs(9521);
    outputs(2312) <= (layer4_outputs(4216)) xor (layer4_outputs(1284));
    outputs(2313) <= not(layer4_outputs(11));
    outputs(2314) <= not((layer4_outputs(9977)) xor (layer4_outputs(4996)));
    outputs(2315) <= not((layer4_outputs(5581)) and (layer4_outputs(7865)));
    outputs(2316) <= layer4_outputs(24);
    outputs(2317) <= not((layer4_outputs(8395)) xor (layer4_outputs(6886)));
    outputs(2318) <= not((layer4_outputs(5745)) or (layer4_outputs(7307)));
    outputs(2319) <= layer4_outputs(5530);
    outputs(2320) <= (layer4_outputs(791)) xor (layer4_outputs(7795));
    outputs(2321) <= (layer4_outputs(479)) and (layer4_outputs(6541));
    outputs(2322) <= not(layer4_outputs(6672));
    outputs(2323) <= layer4_outputs(3555);
    outputs(2324) <= layer4_outputs(7118);
    outputs(2325) <= (layer4_outputs(2360)) xor (layer4_outputs(3542));
    outputs(2326) <= not(layer4_outputs(6818));
    outputs(2327) <= not(layer4_outputs(6511));
    outputs(2328) <= (layer4_outputs(3208)) xor (layer4_outputs(6135));
    outputs(2329) <= not(layer4_outputs(5468));
    outputs(2330) <= (layer4_outputs(5466)) and not (layer4_outputs(3372));
    outputs(2331) <= layer4_outputs(6597);
    outputs(2332) <= layer4_outputs(6655);
    outputs(2333) <= not(layer4_outputs(838));
    outputs(2334) <= layer4_outputs(2263);
    outputs(2335) <= layer4_outputs(956);
    outputs(2336) <= layer4_outputs(9165);
    outputs(2337) <= layer4_outputs(4969);
    outputs(2338) <= (layer4_outputs(6094)) xor (layer4_outputs(3062));
    outputs(2339) <= not((layer4_outputs(9766)) and (layer4_outputs(6649)));
    outputs(2340) <= not(layer4_outputs(7783));
    outputs(2341) <= layer4_outputs(4712);
    outputs(2342) <= (layer4_outputs(8402)) xor (layer4_outputs(9604));
    outputs(2343) <= not(layer4_outputs(5796));
    outputs(2344) <= not((layer4_outputs(189)) and (layer4_outputs(7343)));
    outputs(2345) <= not((layer4_outputs(9283)) xor (layer4_outputs(4136)));
    outputs(2346) <= not(layer4_outputs(7005));
    outputs(2347) <= layer4_outputs(2472);
    outputs(2348) <= layer4_outputs(169);
    outputs(2349) <= (layer4_outputs(3810)) or (layer4_outputs(4992));
    outputs(2350) <= layer4_outputs(8579);
    outputs(2351) <= not(layer4_outputs(3697));
    outputs(2352) <= layer4_outputs(5292);
    outputs(2353) <= layer4_outputs(1230);
    outputs(2354) <= not(layer4_outputs(2665));
    outputs(2355) <= not((layer4_outputs(8280)) and (layer4_outputs(922)));
    outputs(2356) <= not((layer4_outputs(3950)) xor (layer4_outputs(8586)));
    outputs(2357) <= layer4_outputs(3873);
    outputs(2358) <= '1';
    outputs(2359) <= layer4_outputs(7173);
    outputs(2360) <= layer4_outputs(5226);
    outputs(2361) <= not((layer4_outputs(1812)) xor (layer4_outputs(7664)));
    outputs(2362) <= not(layer4_outputs(3930));
    outputs(2363) <= layer4_outputs(3460);
    outputs(2364) <= (layer4_outputs(3811)) xor (layer4_outputs(8261));
    outputs(2365) <= (layer4_outputs(1204)) or (layer4_outputs(5001));
    outputs(2366) <= not(layer4_outputs(2238));
    outputs(2367) <= (layer4_outputs(2686)) xor (layer4_outputs(2729));
    outputs(2368) <= not((layer4_outputs(8562)) and (layer4_outputs(7492)));
    outputs(2369) <= (layer4_outputs(4708)) and not (layer4_outputs(10141));
    outputs(2370) <= not(layer4_outputs(387));
    outputs(2371) <= layer4_outputs(6852);
    outputs(2372) <= layer4_outputs(3316);
    outputs(2373) <= layer4_outputs(978);
    outputs(2374) <= not(layer4_outputs(7458));
    outputs(2375) <= not(layer4_outputs(9536));
    outputs(2376) <= (layer4_outputs(4609)) xor (layer4_outputs(3984));
    outputs(2377) <= not((layer4_outputs(7149)) xor (layer4_outputs(6342)));
    outputs(2378) <= layer4_outputs(2099);
    outputs(2379) <= layer4_outputs(902);
    outputs(2380) <= layer4_outputs(9760);
    outputs(2381) <= not((layer4_outputs(4955)) xor (layer4_outputs(6602)));
    outputs(2382) <= not((layer4_outputs(5748)) xor (layer4_outputs(6207)));
    outputs(2383) <= not(layer4_outputs(3511));
    outputs(2384) <= (layer4_outputs(9687)) and not (layer4_outputs(9224));
    outputs(2385) <= not(layer4_outputs(4786));
    outputs(2386) <= not(layer4_outputs(3579));
    outputs(2387) <= layer4_outputs(6347);
    outputs(2388) <= not(layer4_outputs(3664)) or (layer4_outputs(7838));
    outputs(2389) <= (layer4_outputs(2219)) xor (layer4_outputs(353));
    outputs(2390) <= not((layer4_outputs(8449)) or (layer4_outputs(6612)));
    outputs(2391) <= not(layer4_outputs(10203));
    outputs(2392) <= not((layer4_outputs(4290)) xor (layer4_outputs(5316)));
    outputs(2393) <= (layer4_outputs(9775)) xor (layer4_outputs(9416));
    outputs(2394) <= not(layer4_outputs(4051));
    outputs(2395) <= not((layer4_outputs(6646)) and (layer4_outputs(2314)));
    outputs(2396) <= layer4_outputs(1285);
    outputs(2397) <= (layer4_outputs(5612)) or (layer4_outputs(4380));
    outputs(2398) <= (layer4_outputs(10012)) and (layer4_outputs(8213));
    outputs(2399) <= not(layer4_outputs(6148));
    outputs(2400) <= layer4_outputs(7644);
    outputs(2401) <= not((layer4_outputs(4361)) xor (layer4_outputs(4011)));
    outputs(2402) <= layer4_outputs(354);
    outputs(2403) <= (layer4_outputs(10239)) xor (layer4_outputs(4814));
    outputs(2404) <= (layer4_outputs(2814)) and not (layer4_outputs(1755));
    outputs(2405) <= not(layer4_outputs(6999));
    outputs(2406) <= layer4_outputs(1297);
    outputs(2407) <= (layer4_outputs(4820)) xor (layer4_outputs(7168));
    outputs(2408) <= not((layer4_outputs(9868)) xor (layer4_outputs(3425)));
    outputs(2409) <= not((layer4_outputs(2563)) xor (layer4_outputs(2713)));
    outputs(2410) <= layer4_outputs(7944);
    outputs(2411) <= layer4_outputs(539);
    outputs(2412) <= layer4_outputs(1683);
    outputs(2413) <= not(layer4_outputs(7784));
    outputs(2414) <= layer4_outputs(9771);
    outputs(2415) <= not(layer4_outputs(8154));
    outputs(2416) <= layer4_outputs(6325);
    outputs(2417) <= layer4_outputs(4580);
    outputs(2418) <= layer4_outputs(7690);
    outputs(2419) <= not(layer4_outputs(965));
    outputs(2420) <= layer4_outputs(7813);
    outputs(2421) <= (layer4_outputs(1074)) and not (layer4_outputs(10208));
    outputs(2422) <= not(layer4_outputs(538));
    outputs(2423) <= (layer4_outputs(6990)) xor (layer4_outputs(4106));
    outputs(2424) <= layer4_outputs(878);
    outputs(2425) <= not((layer4_outputs(3488)) and (layer4_outputs(4363)));
    outputs(2426) <= layer4_outputs(6413);
    outputs(2427) <= not(layer4_outputs(8569));
    outputs(2428) <= layer4_outputs(4267);
    outputs(2429) <= not((layer4_outputs(8214)) xor (layer4_outputs(4982)));
    outputs(2430) <= layer4_outputs(2419);
    outputs(2431) <= not((layer4_outputs(5905)) and (layer4_outputs(9382)));
    outputs(2432) <= not((layer4_outputs(2992)) xor (layer4_outputs(2269)));
    outputs(2433) <= not(layer4_outputs(8425));
    outputs(2434) <= not(layer4_outputs(9796));
    outputs(2435) <= layer4_outputs(6946);
    outputs(2436) <= layer4_outputs(6113);
    outputs(2437) <= (layer4_outputs(2079)) and not (layer4_outputs(8949));
    outputs(2438) <= not(layer4_outputs(8370));
    outputs(2439) <= not(layer4_outputs(3416));
    outputs(2440) <= not(layer4_outputs(8367)) or (layer4_outputs(7568));
    outputs(2441) <= layer4_outputs(4490);
    outputs(2442) <= (layer4_outputs(9430)) xor (layer4_outputs(9113));
    outputs(2443) <= '0';
    outputs(2444) <= layer4_outputs(3911);
    outputs(2445) <= (layer4_outputs(9000)) xor (layer4_outputs(9140));
    outputs(2446) <= layer4_outputs(8251);
    outputs(2447) <= layer4_outputs(6962);
    outputs(2448) <= layer4_outputs(5956);
    outputs(2449) <= not((layer4_outputs(161)) or (layer4_outputs(882)));
    outputs(2450) <= layer4_outputs(6460);
    outputs(2451) <= layer4_outputs(3183);
    outputs(2452) <= not(layer4_outputs(3567));
    outputs(2453) <= (layer4_outputs(6741)) xor (layer4_outputs(5017));
    outputs(2454) <= not(layer4_outputs(2454));
    outputs(2455) <= layer4_outputs(8961);
    outputs(2456) <= not(layer4_outputs(3933));
    outputs(2457) <= layer4_outputs(1557);
    outputs(2458) <= not(layer4_outputs(3213));
    outputs(2459) <= layer4_outputs(8839);
    outputs(2460) <= not((layer4_outputs(3955)) xor (layer4_outputs(6905)));
    outputs(2461) <= not((layer4_outputs(7294)) xor (layer4_outputs(9577)));
    outputs(2462) <= not(layer4_outputs(9717)) or (layer4_outputs(87));
    outputs(2463) <= not((layer4_outputs(1111)) and (layer4_outputs(9682)));
    outputs(2464) <= not(layer4_outputs(7469));
    outputs(2465) <= layer4_outputs(10226);
    outputs(2466) <= not((layer4_outputs(9947)) and (layer4_outputs(3633)));
    outputs(2467) <= (layer4_outputs(6092)) and not (layer4_outputs(9057));
    outputs(2468) <= not(layer4_outputs(7134));
    outputs(2469) <= not((layer4_outputs(7845)) xor (layer4_outputs(1153)));
    outputs(2470) <= not(layer4_outputs(2820));
    outputs(2471) <= not(layer4_outputs(2873));
    outputs(2472) <= (layer4_outputs(9250)) xor (layer4_outputs(1623));
    outputs(2473) <= (layer4_outputs(9982)) or (layer4_outputs(1228));
    outputs(2474) <= layer4_outputs(461);
    outputs(2475) <= layer4_outputs(5500);
    outputs(2476) <= not(layer4_outputs(10079));
    outputs(2477) <= layer4_outputs(6727);
    outputs(2478) <= not(layer4_outputs(6041));
    outputs(2479) <= not(layer4_outputs(3759)) or (layer4_outputs(5012));
    outputs(2480) <= not(layer4_outputs(5155)) or (layer4_outputs(4411));
    outputs(2481) <= layer4_outputs(6280);
    outputs(2482) <= layer4_outputs(6079);
    outputs(2483) <= (layer4_outputs(6995)) xor (layer4_outputs(10226));
    outputs(2484) <= not((layer4_outputs(468)) xor (layer4_outputs(6326)));
    outputs(2485) <= layer4_outputs(5088);
    outputs(2486) <= not(layer4_outputs(8331));
    outputs(2487) <= (layer4_outputs(2629)) xor (layer4_outputs(1255));
    outputs(2488) <= not(layer4_outputs(8741));
    outputs(2489) <= not(layer4_outputs(4564));
    outputs(2490) <= (layer4_outputs(3915)) xor (layer4_outputs(6470));
    outputs(2491) <= (layer4_outputs(1594)) xor (layer4_outputs(8986));
    outputs(2492) <= not(layer4_outputs(2279)) or (layer4_outputs(3814));
    outputs(2493) <= not((layer4_outputs(6114)) or (layer4_outputs(4570)));
    outputs(2494) <= not(layer4_outputs(7012));
    outputs(2495) <= layer4_outputs(10230);
    outputs(2496) <= not(layer4_outputs(9663));
    outputs(2497) <= (layer4_outputs(3206)) xor (layer4_outputs(9381));
    outputs(2498) <= not(layer4_outputs(152));
    outputs(2499) <= not((layer4_outputs(248)) xor (layer4_outputs(5814)));
    outputs(2500) <= layer4_outputs(1549);
    outputs(2501) <= (layer4_outputs(9847)) xor (layer4_outputs(2229));
    outputs(2502) <= layer4_outputs(8);
    outputs(2503) <= (layer4_outputs(111)) xor (layer4_outputs(3829));
    outputs(2504) <= layer4_outputs(3920);
    outputs(2505) <= (layer4_outputs(3404)) xor (layer4_outputs(5201));
    outputs(2506) <= layer4_outputs(8989);
    outputs(2507) <= (layer4_outputs(7868)) xor (layer4_outputs(5121));
    outputs(2508) <= not((layer4_outputs(9236)) xor (layer4_outputs(8046)));
    outputs(2509) <= (layer4_outputs(884)) or (layer4_outputs(7015));
    outputs(2510) <= not((layer4_outputs(8228)) xor (layer4_outputs(3325)));
    outputs(2511) <= not((layer4_outputs(7906)) xor (layer4_outputs(7898)));
    outputs(2512) <= not((layer4_outputs(572)) or (layer4_outputs(713)));
    outputs(2513) <= layer4_outputs(4977);
    outputs(2514) <= not((layer4_outputs(3927)) xor (layer4_outputs(2228)));
    outputs(2515) <= layer4_outputs(7137);
    outputs(2516) <= layer4_outputs(7172);
    outputs(2517) <= layer4_outputs(1880);
    outputs(2518) <= not(layer4_outputs(4283));
    outputs(2519) <= (layer4_outputs(3809)) xor (layer4_outputs(6811));
    outputs(2520) <= layer4_outputs(5973);
    outputs(2521) <= layer4_outputs(9718);
    outputs(2522) <= not(layer4_outputs(1437));
    outputs(2523) <= not((layer4_outputs(5503)) and (layer4_outputs(275)));
    outputs(2524) <= (layer4_outputs(7152)) xor (layer4_outputs(8995));
    outputs(2525) <= not(layer4_outputs(1961));
    outputs(2526) <= layer4_outputs(8803);
    outputs(2527) <= (layer4_outputs(2747)) xor (layer4_outputs(6352));
    outputs(2528) <= not((layer4_outputs(3973)) or (layer4_outputs(7960)));
    outputs(2529) <= not((layer4_outputs(7062)) xor (layer4_outputs(5422)));
    outputs(2530) <= not(layer4_outputs(9665)) or (layer4_outputs(5750));
    outputs(2531) <= not(layer4_outputs(422));
    outputs(2532) <= not(layer4_outputs(6596));
    outputs(2533) <= not(layer4_outputs(6233));
    outputs(2534) <= not((layer4_outputs(8875)) xor (layer4_outputs(8471)));
    outputs(2535) <= layer4_outputs(2519);
    outputs(2536) <= not(layer4_outputs(5650));
    outputs(2537) <= not((layer4_outputs(9058)) and (layer4_outputs(6600)));
    outputs(2538) <= not(layer4_outputs(9322));
    outputs(2539) <= not(layer4_outputs(2710));
    outputs(2540) <= not((layer4_outputs(1313)) xor (layer4_outputs(6788)));
    outputs(2541) <= (layer4_outputs(8372)) xor (layer4_outputs(489));
    outputs(2542) <= not(layer4_outputs(2373));
    outputs(2543) <= layer4_outputs(7887);
    outputs(2544) <= layer4_outputs(3519);
    outputs(2545) <= not(layer4_outputs(5572));
    outputs(2546) <= not((layer4_outputs(3444)) xor (layer4_outputs(6660)));
    outputs(2547) <= layer4_outputs(1647);
    outputs(2548) <= not(layer4_outputs(7362)) or (layer4_outputs(5549));
    outputs(2549) <= not(layer4_outputs(7195));
    outputs(2550) <= not(layer4_outputs(7083));
    outputs(2551) <= not((layer4_outputs(7017)) xor (layer4_outputs(1542)));
    outputs(2552) <= not(layer4_outputs(4637));
    outputs(2553) <= layer4_outputs(120);
    outputs(2554) <= (layer4_outputs(1701)) xor (layer4_outputs(3963));
    outputs(2555) <= not(layer4_outputs(4960));
    outputs(2556) <= not((layer4_outputs(2187)) xor (layer4_outputs(1600)));
    outputs(2557) <= (layer4_outputs(8418)) and not (layer4_outputs(4206));
    outputs(2558) <= not(layer4_outputs(10031)) or (layer4_outputs(10000));
    outputs(2559) <= not((layer4_outputs(8821)) and (layer4_outputs(435)));
    outputs(2560) <= layer4_outputs(2374);
    outputs(2561) <= not(layer4_outputs(2198)) or (layer4_outputs(9833));
    outputs(2562) <= layer4_outputs(3054);
    outputs(2563) <= not(layer4_outputs(6710));
    outputs(2564) <= layer4_outputs(6157);
    outputs(2565) <= layer4_outputs(2845);
    outputs(2566) <= layer4_outputs(9669);
    outputs(2567) <= layer4_outputs(3503);
    outputs(2568) <= not(layer4_outputs(4480));
    outputs(2569) <= not(layer4_outputs(2817));
    outputs(2570) <= layer4_outputs(661);
    outputs(2571) <= not(layer4_outputs(741));
    outputs(2572) <= not(layer4_outputs(4831));
    outputs(2573) <= (layer4_outputs(2868)) and (layer4_outputs(7191));
    outputs(2574) <= not((layer4_outputs(8508)) and (layer4_outputs(5560)));
    outputs(2575) <= layer4_outputs(2558);
    outputs(2576) <= (layer4_outputs(3840)) xor (layer4_outputs(3298));
    outputs(2577) <= not(layer4_outputs(7295));
    outputs(2578) <= not((layer4_outputs(9373)) xor (layer4_outputs(3384)));
    outputs(2579) <= not(layer4_outputs(6346));
    outputs(2580) <= not(layer4_outputs(8630));
    outputs(2581) <= layer4_outputs(42);
    outputs(2582) <= not(layer4_outputs(8672));
    outputs(2583) <= layer4_outputs(5673);
    outputs(2584) <= not(layer4_outputs(1581));
    outputs(2585) <= layer4_outputs(1803);
    outputs(2586) <= not(layer4_outputs(10131));
    outputs(2587) <= not(layer4_outputs(8159)) or (layer4_outputs(4738));
    outputs(2588) <= not(layer4_outputs(957));
    outputs(2589) <= layer4_outputs(1493);
    outputs(2590) <= layer4_outputs(7252);
    outputs(2591) <= (layer4_outputs(2236)) or (layer4_outputs(5669));
    outputs(2592) <= not(layer4_outputs(9028));
    outputs(2593) <= (layer4_outputs(2)) xor (layer4_outputs(3338));
    outputs(2594) <= not((layer4_outputs(6666)) xor (layer4_outputs(2342)));
    outputs(2595) <= not(layer4_outputs(647));
    outputs(2596) <= (layer4_outputs(2284)) and not (layer4_outputs(5437));
    outputs(2597) <= not((layer4_outputs(3652)) xor (layer4_outputs(6149)));
    outputs(2598) <= layer4_outputs(1253);
    outputs(2599) <= (layer4_outputs(305)) xor (layer4_outputs(1796));
    outputs(2600) <= layer4_outputs(3959);
    outputs(2601) <= layer4_outputs(7127);
    outputs(2602) <= (layer4_outputs(2226)) xor (layer4_outputs(2260));
    outputs(2603) <= (layer4_outputs(1741)) xor (layer4_outputs(935));
    outputs(2604) <= layer4_outputs(8544);
    outputs(2605) <= layer4_outputs(2712);
    outputs(2606) <= not((layer4_outputs(4910)) xor (layer4_outputs(5522)));
    outputs(2607) <= (layer4_outputs(8320)) and (layer4_outputs(8051));
    outputs(2608) <= not(layer4_outputs(1162)) or (layer4_outputs(1658));
    outputs(2609) <= not(layer4_outputs(338));
    outputs(2610) <= layer4_outputs(4530);
    outputs(2611) <= layer4_outputs(7996);
    outputs(2612) <= (layer4_outputs(5464)) and not (layer4_outputs(214));
    outputs(2613) <= not(layer4_outputs(6116));
    outputs(2614) <= not(layer4_outputs(1156));
    outputs(2615) <= not((layer4_outputs(8825)) or (layer4_outputs(7712)));
    outputs(2616) <= not(layer4_outputs(6027));
    outputs(2617) <= not((layer4_outputs(7483)) xor (layer4_outputs(7786)));
    outputs(2618) <= layer4_outputs(5233);
    outputs(2619) <= (layer4_outputs(306)) and not (layer4_outputs(2913));
    outputs(2620) <= (layer4_outputs(612)) and not (layer4_outputs(8368));
    outputs(2621) <= not(layer4_outputs(6880));
    outputs(2622) <= not(layer4_outputs(6043));
    outputs(2623) <= (layer4_outputs(6846)) xor (layer4_outputs(1984));
    outputs(2624) <= layer4_outputs(898);
    outputs(2625) <= not(layer4_outputs(10165));
    outputs(2626) <= not((layer4_outputs(7411)) xor (layer4_outputs(3954)));
    outputs(2627) <= not(layer4_outputs(5846));
    outputs(2628) <= not(layer4_outputs(9700));
    outputs(2629) <= not(layer4_outputs(8243));
    outputs(2630) <= not(layer4_outputs(3492));
    outputs(2631) <= not((layer4_outputs(7428)) xor (layer4_outputs(1521)));
    outputs(2632) <= (layer4_outputs(1119)) xor (layer4_outputs(6514));
    outputs(2633) <= layer4_outputs(1186);
    outputs(2634) <= not((layer4_outputs(3806)) and (layer4_outputs(1064)));
    outputs(2635) <= layer4_outputs(7039);
    outputs(2636) <= (layer4_outputs(1981)) or (layer4_outputs(2431));
    outputs(2637) <= (layer4_outputs(1529)) xor (layer4_outputs(9837));
    outputs(2638) <= (layer4_outputs(4385)) xor (layer4_outputs(4882));
    outputs(2639) <= (layer4_outputs(9097)) xor (layer4_outputs(3598));
    outputs(2640) <= layer4_outputs(7773);
    outputs(2641) <= (layer4_outputs(3865)) xor (layer4_outputs(8662));
    outputs(2642) <= (layer4_outputs(1720)) xor (layer4_outputs(2673));
    outputs(2643) <= not(layer4_outputs(7319));
    outputs(2644) <= layer4_outputs(10085);
    outputs(2645) <= not(layer4_outputs(6899));
    outputs(2646) <= layer4_outputs(3669);
    outputs(2647) <= not((layer4_outputs(8783)) and (layer4_outputs(8220)));
    outputs(2648) <= not(layer4_outputs(4956));
    outputs(2649) <= not(layer4_outputs(390)) or (layer4_outputs(8534));
    outputs(2650) <= not((layer4_outputs(3781)) and (layer4_outputs(6273)));
    outputs(2651) <= not(layer4_outputs(5458));
    outputs(2652) <= layer4_outputs(1508);
    outputs(2653) <= '0';
    outputs(2654) <= not((layer4_outputs(3307)) xor (layer4_outputs(3409)));
    outputs(2655) <= layer4_outputs(4512);
    outputs(2656) <= layer4_outputs(735);
    outputs(2657) <= not(layer4_outputs(4210));
    outputs(2658) <= layer4_outputs(4243);
    outputs(2659) <= layer4_outputs(4223);
    outputs(2660) <= (layer4_outputs(3824)) and not (layer4_outputs(6394));
    outputs(2661) <= not(layer4_outputs(3353));
    outputs(2662) <= layer4_outputs(6563);
    outputs(2663) <= layer4_outputs(8721);
    outputs(2664) <= not((layer4_outputs(173)) or (layer4_outputs(2268)));
    outputs(2665) <= not(layer4_outputs(3972));
    outputs(2666) <= not(layer4_outputs(7420)) or (layer4_outputs(3682));
    outputs(2667) <= not(layer4_outputs(9253));
    outputs(2668) <= layer4_outputs(8832);
    outputs(2669) <= layer4_outputs(3642);
    outputs(2670) <= layer4_outputs(4078);
    outputs(2671) <= not(layer4_outputs(2301));
    outputs(2672) <= not((layer4_outputs(5875)) xor (layer4_outputs(9199)));
    outputs(2673) <= not(layer4_outputs(5495));
    outputs(2674) <= (layer4_outputs(6916)) xor (layer4_outputs(4187));
    outputs(2675) <= (layer4_outputs(3844)) xor (layer4_outputs(7186));
    outputs(2676) <= not((layer4_outputs(4110)) xor (layer4_outputs(8660)));
    outputs(2677) <= layer4_outputs(280);
    outputs(2678) <= layer4_outputs(1106);
    outputs(2679) <= (layer4_outputs(2026)) xor (layer4_outputs(1382));
    outputs(2680) <= (layer4_outputs(7933)) xor (layer4_outputs(7673));
    outputs(2681) <= not((layer4_outputs(6547)) xor (layer4_outputs(1478)));
    outputs(2682) <= not((layer4_outputs(9542)) xor (layer4_outputs(2280)));
    outputs(2683) <= not(layer4_outputs(846));
    outputs(2684) <= not(layer4_outputs(8089));
    outputs(2685) <= not(layer4_outputs(5273));
    outputs(2686) <= not(layer4_outputs(7691));
    outputs(2687) <= not((layer4_outputs(3659)) xor (layer4_outputs(1322)));
    outputs(2688) <= (layer4_outputs(1036)) and not (layer4_outputs(4322));
    outputs(2689) <= not((layer4_outputs(2262)) xor (layer4_outputs(2401)));
    outputs(2690) <= not(layer4_outputs(8630));
    outputs(2691) <= not(layer4_outputs(1037));
    outputs(2692) <= not((layer4_outputs(9371)) xor (layer4_outputs(5037)));
    outputs(2693) <= (layer4_outputs(9888)) and not (layer4_outputs(3847));
    outputs(2694) <= not(layer4_outputs(7654));
    outputs(2695) <= not(layer4_outputs(7592));
    outputs(2696) <= (layer4_outputs(2872)) xor (layer4_outputs(3025));
    outputs(2697) <= layer4_outputs(9268);
    outputs(2698) <= (layer4_outputs(5544)) xor (layer4_outputs(1735));
    outputs(2699) <= layer4_outputs(3048);
    outputs(2700) <= not((layer4_outputs(8610)) xor (layer4_outputs(6111)));
    outputs(2701) <= (layer4_outputs(8843)) xor (layer4_outputs(8440));
    outputs(2702) <= not((layer4_outputs(4184)) xor (layer4_outputs(4564)));
    outputs(2703) <= layer4_outputs(1937);
    outputs(2704) <= not(layer4_outputs(3746));
    outputs(2705) <= not(layer4_outputs(8928));
    outputs(2706) <= not((layer4_outputs(2265)) xor (layer4_outputs(4898)));
    outputs(2707) <= (layer4_outputs(3000)) and (layer4_outputs(6284));
    outputs(2708) <= not((layer4_outputs(2258)) xor (layer4_outputs(10008)));
    outputs(2709) <= (layer4_outputs(1735)) xor (layer4_outputs(3373));
    outputs(2710) <= (layer4_outputs(4032)) or (layer4_outputs(9110));
    outputs(2711) <= not(layer4_outputs(4717));
    outputs(2712) <= not(layer4_outputs(384));
    outputs(2713) <= not(layer4_outputs(1776));
    outputs(2714) <= (layer4_outputs(870)) and not (layer4_outputs(5931));
    outputs(2715) <= not(layer4_outputs(10093));
    outputs(2716) <= layer4_outputs(7744);
    outputs(2717) <= (layer4_outputs(9177)) and not (layer4_outputs(1946));
    outputs(2718) <= (layer4_outputs(998)) xor (layer4_outputs(1001));
    outputs(2719) <= not(layer4_outputs(5281));
    outputs(2720) <= not((layer4_outputs(7934)) xor (layer4_outputs(6398)));
    outputs(2721) <= layer4_outputs(9287);
    outputs(2722) <= (layer4_outputs(6620)) xor (layer4_outputs(7210));
    outputs(2723) <= layer4_outputs(6508);
    outputs(2724) <= layer4_outputs(8152);
    outputs(2725) <= not(layer4_outputs(6952)) or (layer4_outputs(4921));
    outputs(2726) <= (layer4_outputs(7773)) xor (layer4_outputs(5588));
    outputs(2727) <= not(layer4_outputs(693));
    outputs(2728) <= layer4_outputs(277);
    outputs(2729) <= (layer4_outputs(8371)) xor (layer4_outputs(9903));
    outputs(2730) <= not(layer4_outputs(4359));
    outputs(2731) <= (layer4_outputs(3222)) xor (layer4_outputs(6550));
    outputs(2732) <= (layer4_outputs(5398)) xor (layer4_outputs(4299));
    outputs(2733) <= '1';
    outputs(2734) <= not(layer4_outputs(6576));
    outputs(2735) <= not(layer4_outputs(8403));
    outputs(2736) <= not((layer4_outputs(245)) xor (layer4_outputs(8215)));
    outputs(2737) <= layer4_outputs(9131);
    outputs(2738) <= (layer4_outputs(7347)) and (layer4_outputs(3002));
    outputs(2739) <= layer4_outputs(157);
    outputs(2740) <= not(layer4_outputs(5984));
    outputs(2741) <= (layer4_outputs(7037)) or (layer4_outputs(5483));
    outputs(2742) <= (layer4_outputs(8017)) xor (layer4_outputs(8353));
    outputs(2743) <= not((layer4_outputs(6699)) xor (layer4_outputs(314)));
    outputs(2744) <= layer4_outputs(5142);
    outputs(2745) <= layer4_outputs(5687);
    outputs(2746) <= layer4_outputs(4281);
    outputs(2747) <= layer4_outputs(3008);
    outputs(2748) <= (layer4_outputs(4510)) or (layer4_outputs(4950));
    outputs(2749) <= layer4_outputs(3805);
    outputs(2750) <= not(layer4_outputs(2759)) or (layer4_outputs(5731));
    outputs(2751) <= not(layer4_outputs(1207));
    outputs(2752) <= layer4_outputs(8822);
    outputs(2753) <= layer4_outputs(3594);
    outputs(2754) <= not((layer4_outputs(7831)) or (layer4_outputs(5257)));
    outputs(2755) <= not(layer4_outputs(6346));
    outputs(2756) <= layer4_outputs(8028);
    outputs(2757) <= not(layer4_outputs(4404));
    outputs(2758) <= layer4_outputs(800);
    outputs(2759) <= (layer4_outputs(465)) and (layer4_outputs(6779));
    outputs(2760) <= not(layer4_outputs(3160));
    outputs(2761) <= not((layer4_outputs(7119)) xor (layer4_outputs(2516)));
    outputs(2762) <= not(layer4_outputs(8389));
    outputs(2763) <= layer4_outputs(5091);
    outputs(2764) <= not(layer4_outputs(6041)) or (layer4_outputs(1031));
    outputs(2765) <= not(layer4_outputs(9246));
    outputs(2766) <= layer4_outputs(2620);
    outputs(2767) <= not((layer4_outputs(9583)) xor (layer4_outputs(1832)));
    outputs(2768) <= not((layer4_outputs(5918)) xor (layer4_outputs(3512)));
    outputs(2769) <= layer4_outputs(8085);
    outputs(2770) <= layer4_outputs(6570);
    outputs(2771) <= layer4_outputs(6825);
    outputs(2772) <= not(layer4_outputs(6497));
    outputs(2773) <= layer4_outputs(2153);
    outputs(2774) <= layer4_outputs(8734);
    outputs(2775) <= not(layer4_outputs(8184)) or (layer4_outputs(9801));
    outputs(2776) <= not((layer4_outputs(2805)) xor (layer4_outputs(8940)));
    outputs(2777) <= layer4_outputs(3871);
    outputs(2778) <= layer4_outputs(5006);
    outputs(2779) <= not(layer4_outputs(4403));
    outputs(2780) <= not(layer4_outputs(1145));
    outputs(2781) <= not((layer4_outputs(3990)) xor (layer4_outputs(8242)));
    outputs(2782) <= (layer4_outputs(1177)) xor (layer4_outputs(3614));
    outputs(2783) <= not(layer4_outputs(4732));
    outputs(2784) <= layer4_outputs(7297);
    outputs(2785) <= layer4_outputs(7203);
    outputs(2786) <= layer4_outputs(8348);
    outputs(2787) <= layer4_outputs(7211);
    outputs(2788) <= not((layer4_outputs(8749)) xor (layer4_outputs(6186)));
    outputs(2789) <= not((layer4_outputs(5239)) xor (layer4_outputs(8272)));
    outputs(2790) <= layer4_outputs(3608);
    outputs(2791) <= not(layer4_outputs(6146));
    outputs(2792) <= layer4_outputs(4344);
    outputs(2793) <= not(layer4_outputs(5520)) or (layer4_outputs(1063));
    outputs(2794) <= not(layer4_outputs(10005));
    outputs(2795) <= (layer4_outputs(7740)) xor (layer4_outputs(7738));
    outputs(2796) <= (layer4_outputs(8026)) or (layer4_outputs(4867));
    outputs(2797) <= not(layer4_outputs(1473));
    outputs(2798) <= not(layer4_outputs(6135));
    outputs(2799) <= not((layer4_outputs(744)) xor (layer4_outputs(9492)));
    outputs(2800) <= layer4_outputs(7446);
    outputs(2801) <= layer4_outputs(5811);
    outputs(2802) <= not(layer4_outputs(3983));
    outputs(2803) <= layer4_outputs(464);
    outputs(2804) <= not((layer4_outputs(10116)) xor (layer4_outputs(6450)));
    outputs(2805) <= layer4_outputs(9569);
    outputs(2806) <= not((layer4_outputs(4397)) xor (layer4_outputs(6407)));
    outputs(2807) <= (layer4_outputs(6984)) xor (layer4_outputs(467));
    outputs(2808) <= layer4_outputs(1190);
    outputs(2809) <= not(layer4_outputs(9575));
    outputs(2810) <= layer4_outputs(2566);
    outputs(2811) <= not(layer4_outputs(4758)) or (layer4_outputs(8639));
    outputs(2812) <= layer4_outputs(4867);
    outputs(2813) <= layer4_outputs(6280);
    outputs(2814) <= (layer4_outputs(7393)) and not (layer4_outputs(2128));
    outputs(2815) <= not(layer4_outputs(928));
    outputs(2816) <= not((layer4_outputs(8788)) xor (layer4_outputs(6064)));
    outputs(2817) <= not(layer4_outputs(1576)) or (layer4_outputs(8429));
    outputs(2818) <= (layer4_outputs(8317)) xor (layer4_outputs(9505));
    outputs(2819) <= not(layer4_outputs(9723));
    outputs(2820) <= layer4_outputs(4704);
    outputs(2821) <= not((layer4_outputs(8789)) or (layer4_outputs(6599)));
    outputs(2822) <= not(layer4_outputs(8791));
    outputs(2823) <= layer4_outputs(1823);
    outputs(2824) <= not(layer4_outputs(8647));
    outputs(2825) <= not((layer4_outputs(7465)) xor (layer4_outputs(7871)));
    outputs(2826) <= not(layer4_outputs(3483));
    outputs(2827) <= layer4_outputs(2199);
    outputs(2828) <= layer4_outputs(3110);
    outputs(2829) <= layer4_outputs(10123);
    outputs(2830) <= not(layer4_outputs(8675));
    outputs(2831) <= (layer4_outputs(5841)) and not (layer4_outputs(9368));
    outputs(2832) <= not((layer4_outputs(1482)) xor (layer4_outputs(5080)));
    outputs(2833) <= not(layer4_outputs(395));
    outputs(2834) <= not(layer4_outputs(9297));
    outputs(2835) <= layer4_outputs(9969);
    outputs(2836) <= not((layer4_outputs(4279)) and (layer4_outputs(6429)));
    outputs(2837) <= not((layer4_outputs(6316)) and (layer4_outputs(6202)));
    outputs(2838) <= layer4_outputs(8029);
    outputs(2839) <= layer4_outputs(5052);
    outputs(2840) <= not(layer4_outputs(1266));
    outputs(2841) <= not(layer4_outputs(4681));
    outputs(2842) <= not(layer4_outputs(6));
    outputs(2843) <= not(layer4_outputs(5134));
    outputs(2844) <= not(layer4_outputs(4320));
    outputs(2845) <= not((layer4_outputs(5329)) and (layer4_outputs(3695)));
    outputs(2846) <= not(layer4_outputs(1802)) or (layer4_outputs(3258));
    outputs(2847) <= not(layer4_outputs(3908));
    outputs(2848) <= not(layer4_outputs(9889));
    outputs(2849) <= layer4_outputs(4309);
    outputs(2850) <= not(layer4_outputs(8335));
    outputs(2851) <= layer4_outputs(2443);
    outputs(2852) <= layer4_outputs(6289);
    outputs(2853) <= layer4_outputs(2838);
    outputs(2854) <= not(layer4_outputs(8836));
    outputs(2855) <= not(layer4_outputs(4051));
    outputs(2856) <= not(layer4_outputs(6510));
    outputs(2857) <= not((layer4_outputs(9856)) or (layer4_outputs(6608)));
    outputs(2858) <= (layer4_outputs(9038)) xor (layer4_outputs(8860));
    outputs(2859) <= (layer4_outputs(1684)) xor (layer4_outputs(7984));
    outputs(2860) <= layer4_outputs(8212);
    outputs(2861) <= layer4_outputs(1866);
    outputs(2862) <= (layer4_outputs(6157)) and not (layer4_outputs(8928));
    outputs(2863) <= not(layer4_outputs(5089)) or (layer4_outputs(5529));
    outputs(2864) <= not(layer4_outputs(440));
    outputs(2865) <= not(layer4_outputs(3377));
    outputs(2866) <= not(layer4_outputs(7433));
    outputs(2867) <= layer4_outputs(1684);
    outputs(2868) <= layer4_outputs(9432);
    outputs(2869) <= not(layer4_outputs(6375));
    outputs(2870) <= not(layer4_outputs(9209));
    outputs(2871) <= (layer4_outputs(2886)) xor (layer4_outputs(720));
    outputs(2872) <= (layer4_outputs(4209)) or (layer4_outputs(859));
    outputs(2873) <= not((layer4_outputs(9093)) xor (layer4_outputs(1744)));
    outputs(2874) <= not((layer4_outputs(2422)) xor (layer4_outputs(1478)));
    outputs(2875) <= '1';
    outputs(2876) <= not((layer4_outputs(3819)) xor (layer4_outputs(2576)));
    outputs(2877) <= layer4_outputs(6446);
    outputs(2878) <= not((layer4_outputs(9878)) xor (layer4_outputs(5778)));
    outputs(2879) <= not((layer4_outputs(2097)) xor (layer4_outputs(3327)));
    outputs(2880) <= (layer4_outputs(1568)) xor (layer4_outputs(8711));
    outputs(2881) <= layer4_outputs(6848);
    outputs(2882) <= not((layer4_outputs(6340)) and (layer4_outputs(2662)));
    outputs(2883) <= layer4_outputs(1434);
    outputs(2884) <= layer4_outputs(8065);
    outputs(2885) <= not(layer4_outputs(8364));
    outputs(2886) <= layer4_outputs(6366);
    outputs(2887) <= layer4_outputs(443);
    outputs(2888) <= not(layer4_outputs(3006)) or (layer4_outputs(3009));
    outputs(2889) <= not(layer4_outputs(3930));
    outputs(2890) <= (layer4_outputs(7683)) or (layer4_outputs(8911));
    outputs(2891) <= not(layer4_outputs(29));
    outputs(2892) <= layer4_outputs(285);
    outputs(2893) <= not(layer4_outputs(5597));
    outputs(2894) <= layer4_outputs(7089);
    outputs(2895) <= layer4_outputs(710);
    outputs(2896) <= not(layer4_outputs(6672));
    outputs(2897) <= not(layer4_outputs(7532));
    outputs(2898) <= layer4_outputs(6035);
    outputs(2899) <= layer4_outputs(7038);
    outputs(2900) <= (layer4_outputs(711)) xor (layer4_outputs(2211));
    outputs(2901) <= (layer4_outputs(5472)) and not (layer4_outputs(4180));
    outputs(2902) <= not((layer4_outputs(7491)) xor (layer4_outputs(5237)));
    outputs(2903) <= layer4_outputs(9933);
    outputs(2904) <= not((layer4_outputs(10109)) xor (layer4_outputs(8614)));
    outputs(2905) <= (layer4_outputs(9976)) and not (layer4_outputs(6894));
    outputs(2906) <= not((layer4_outputs(5639)) xor (layer4_outputs(9653)));
    outputs(2907) <= layer4_outputs(4292);
    outputs(2908) <= not(layer4_outputs(3702)) or (layer4_outputs(7980));
    outputs(2909) <= layer4_outputs(2493);
    outputs(2910) <= not(layer4_outputs(824));
    outputs(2911) <= layer4_outputs(875);
    outputs(2912) <= not(layer4_outputs(5065));
    outputs(2913) <= layer4_outputs(1016);
    outputs(2914) <= layer4_outputs(808);
    outputs(2915) <= not((layer4_outputs(7589)) and (layer4_outputs(9081)));
    outputs(2916) <= layer4_outputs(2681);
    outputs(2917) <= layer4_outputs(2613);
    outputs(2918) <= not((layer4_outputs(6437)) or (layer4_outputs(7097)));
    outputs(2919) <= layer4_outputs(10035);
    outputs(2920) <= not(layer4_outputs(3232));
    outputs(2921) <= layer4_outputs(1077);
    outputs(2922) <= (layer4_outputs(1747)) xor (layer4_outputs(7468));
    outputs(2923) <= (layer4_outputs(5589)) and not (layer4_outputs(4225));
    outputs(2924) <= not(layer4_outputs(2685));
    outputs(2925) <= (layer4_outputs(12)) xor (layer4_outputs(3141));
    outputs(2926) <= (layer4_outputs(10026)) or (layer4_outputs(2213));
    outputs(2927) <= not(layer4_outputs(3692));
    outputs(2928) <= not(layer4_outputs(3448));
    outputs(2929) <= not(layer4_outputs(5563)) or (layer4_outputs(4445));
    outputs(2930) <= not(layer4_outputs(9516)) or (layer4_outputs(8703));
    outputs(2931) <= not(layer4_outputs(4225));
    outputs(2932) <= layer4_outputs(5890);
    outputs(2933) <= (layer4_outputs(1643)) xor (layer4_outputs(7301));
    outputs(2934) <= not(layer4_outputs(6288)) or (layer4_outputs(10061));
    outputs(2935) <= layer4_outputs(266);
    outputs(2936) <= layer4_outputs(1602);
    outputs(2937) <= not(layer4_outputs(8005));
    outputs(2938) <= not(layer4_outputs(4145));
    outputs(2939) <= (layer4_outputs(4640)) and not (layer4_outputs(5903));
    outputs(2940) <= not((layer4_outputs(8278)) xor (layer4_outputs(5103)));
    outputs(2941) <= layer4_outputs(7372);
    outputs(2942) <= not(layer4_outputs(8916));
    outputs(2943) <= layer4_outputs(7522);
    outputs(2944) <= not(layer4_outputs(8496));
    outputs(2945) <= layer4_outputs(5026);
    outputs(2946) <= (layer4_outputs(462)) and not (layer4_outputs(10192));
    outputs(2947) <= (layer4_outputs(1074)) and not (layer4_outputs(5802));
    outputs(2948) <= not(layer4_outputs(8518));
    outputs(2949) <= layer4_outputs(284);
    outputs(2950) <= (layer4_outputs(5870)) xor (layer4_outputs(3952));
    outputs(2951) <= not(layer4_outputs(8099));
    outputs(2952) <= (layer4_outputs(10069)) or (layer4_outputs(4485));
    outputs(2953) <= not((layer4_outputs(8391)) xor (layer4_outputs(5606)));
    outputs(2954) <= not(layer4_outputs(6762));
    outputs(2955) <= not((layer4_outputs(1322)) and (layer4_outputs(8458)));
    outputs(2956) <= not((layer4_outputs(3522)) xor (layer4_outputs(1264)));
    outputs(2957) <= layer4_outputs(8971);
    outputs(2958) <= layer4_outputs(8094);
    outputs(2959) <= layer4_outputs(9006);
    outputs(2960) <= layer4_outputs(7393);
    outputs(2961) <= not(layer4_outputs(8115)) or (layer4_outputs(3317));
    outputs(2962) <= not((layer4_outputs(2157)) xor (layer4_outputs(1816)));
    outputs(2963) <= (layer4_outputs(177)) xor (layer4_outputs(3991));
    outputs(2964) <= layer4_outputs(3276);
    outputs(2965) <= not(layer4_outputs(2782));
    outputs(2966) <= not(layer4_outputs(2854));
    outputs(2967) <= (layer4_outputs(9133)) and not (layer4_outputs(2175));
    outputs(2968) <= layer4_outputs(3817);
    outputs(2969) <= (layer4_outputs(3400)) xor (layer4_outputs(5342));
    outputs(2970) <= not((layer4_outputs(951)) and (layer4_outputs(629)));
    outputs(2971) <= not(layer4_outputs(1715));
    outputs(2972) <= not((layer4_outputs(8921)) xor (layer4_outputs(1495)));
    outputs(2973) <= (layer4_outputs(1471)) xor (layer4_outputs(5660));
    outputs(2974) <= not(layer4_outputs(8305));
    outputs(2975) <= (layer4_outputs(10054)) xor (layer4_outputs(3455));
    outputs(2976) <= not(layer4_outputs(8605));
    outputs(2977) <= not(layer4_outputs(7946));
    outputs(2978) <= layer4_outputs(6760);
    outputs(2979) <= not(layer4_outputs(8381));
    outputs(2980) <= layer4_outputs(5556);
    outputs(2981) <= layer4_outputs(6903);
    outputs(2982) <= not(layer4_outputs(311));
    outputs(2983) <= layer4_outputs(3148);
    outputs(2984) <= not(layer4_outputs(5802));
    outputs(2985) <= layer4_outputs(8650);
    outputs(2986) <= layer4_outputs(2362);
    outputs(2987) <= layer4_outputs(7751);
    outputs(2988) <= not(layer4_outputs(6828));
    outputs(2989) <= not(layer4_outputs(7292));
    outputs(2990) <= not(layer4_outputs(4827));
    outputs(2991) <= not((layer4_outputs(607)) and (layer4_outputs(1839)));
    outputs(2992) <= layer4_outputs(3352);
    outputs(2993) <= not((layer4_outputs(1447)) xor (layer4_outputs(1118)));
    outputs(2994) <= not((layer4_outputs(9851)) xor (layer4_outputs(1295)));
    outputs(2995) <= layer4_outputs(10003);
    outputs(2996) <= layer4_outputs(6147);
    outputs(2997) <= not(layer4_outputs(2907));
    outputs(2998) <= layer4_outputs(3336);
    outputs(2999) <= not(layer4_outputs(7306));
    outputs(3000) <= (layer4_outputs(8947)) xor (layer4_outputs(7750));
    outputs(3001) <= not(layer4_outputs(2499));
    outputs(3002) <= not((layer4_outputs(2386)) xor (layer4_outputs(2307)));
    outputs(3003) <= not(layer4_outputs(3241));
    outputs(3004) <= layer4_outputs(2253);
    outputs(3005) <= not(layer4_outputs(6557));
    outputs(3006) <= layer4_outputs(8036);
    outputs(3007) <= layer4_outputs(153);
    outputs(3008) <= layer4_outputs(6937);
    outputs(3009) <= layer4_outputs(4974);
    outputs(3010) <= not((layer4_outputs(6517)) and (layer4_outputs(5092)));
    outputs(3011) <= (layer4_outputs(9160)) and (layer4_outputs(4929));
    outputs(3012) <= not(layer4_outputs(6380));
    outputs(3013) <= (layer4_outputs(4275)) xor (layer4_outputs(8909));
    outputs(3014) <= layer4_outputs(4201);
    outputs(3015) <= (layer4_outputs(9294)) xor (layer4_outputs(2007));
    outputs(3016) <= (layer4_outputs(6308)) xor (layer4_outputs(5828));
    outputs(3017) <= layer4_outputs(6024);
    outputs(3018) <= not((layer4_outputs(4905)) or (layer4_outputs(9170)));
    outputs(3019) <= not((layer4_outputs(7482)) xor (layer4_outputs(5355)));
    outputs(3020) <= not(layer4_outputs(7798));
    outputs(3021) <= (layer4_outputs(1535)) xor (layer4_outputs(3193));
    outputs(3022) <= not(layer4_outputs(2422)) or (layer4_outputs(9711));
    outputs(3023) <= not((layer4_outputs(3782)) xor (layer4_outputs(7156)));
    outputs(3024) <= layer4_outputs(3090);
    outputs(3025) <= not(layer4_outputs(6195));
    outputs(3026) <= (layer4_outputs(5247)) xor (layer4_outputs(1029));
    outputs(3027) <= layer4_outputs(8844);
    outputs(3028) <= not((layer4_outputs(9934)) xor (layer4_outputs(4807)));
    outputs(3029) <= layer4_outputs(2698);
    outputs(3030) <= (layer4_outputs(1601)) xor (layer4_outputs(157));
    outputs(3031) <= not(layer4_outputs(2995));
    outputs(3032) <= not(layer4_outputs(1562));
    outputs(3033) <= layer4_outputs(7030);
    outputs(3034) <= (layer4_outputs(5429)) xor (layer4_outputs(6815));
    outputs(3035) <= '0';
    outputs(3036) <= layer4_outputs(8871);
    outputs(3037) <= (layer4_outputs(5229)) xor (layer4_outputs(3426));
    outputs(3038) <= not(layer4_outputs(2459));
    outputs(3039) <= not((layer4_outputs(9097)) xor (layer4_outputs(906)));
    outputs(3040) <= not(layer4_outputs(8565));
    outputs(3041) <= not(layer4_outputs(780)) or (layer4_outputs(638));
    outputs(3042) <= not(layer4_outputs(6751)) or (layer4_outputs(6625));
    outputs(3043) <= layer4_outputs(516);
    outputs(3044) <= not(layer4_outputs(1783));
    outputs(3045) <= not(layer4_outputs(6542));
    outputs(3046) <= (layer4_outputs(1485)) xor (layer4_outputs(4385));
    outputs(3047) <= layer4_outputs(9655);
    outputs(3048) <= layer4_outputs(1885);
    outputs(3049) <= layer4_outputs(4326);
    outputs(3050) <= not((layer4_outputs(1452)) xor (layer4_outputs(3698)));
    outputs(3051) <= layer4_outputs(10045);
    outputs(3052) <= not(layer4_outputs(5980)) or (layer4_outputs(6799));
    outputs(3053) <= not((layer4_outputs(4844)) xor (layer4_outputs(537)));
    outputs(3054) <= (layer4_outputs(7738)) and (layer4_outputs(7155));
    outputs(3055) <= not(layer4_outputs(10194));
    outputs(3056) <= not((layer4_outputs(9039)) and (layer4_outputs(5150)));
    outputs(3057) <= layer4_outputs(3547);
    outputs(3058) <= layer4_outputs(431);
    outputs(3059) <= layer4_outputs(4512);
    outputs(3060) <= layer4_outputs(6222);
    outputs(3061) <= not((layer4_outputs(2210)) xor (layer4_outputs(9812)));
    outputs(3062) <= (layer4_outputs(2706)) xor (layer4_outputs(4578));
    outputs(3063) <= not(layer4_outputs(3355));
    outputs(3064) <= layer4_outputs(8756);
    outputs(3065) <= layer4_outputs(2911);
    outputs(3066) <= layer4_outputs(7473);
    outputs(3067) <= not(layer4_outputs(1847));
    outputs(3068) <= not((layer4_outputs(7766)) xor (layer4_outputs(9441)));
    outputs(3069) <= layer4_outputs(2384);
    outputs(3070) <= layer4_outputs(1341);
    outputs(3071) <= not(layer4_outputs(734)) or (layer4_outputs(6622));
    outputs(3072) <= not(layer4_outputs(3769));
    outputs(3073) <= not((layer4_outputs(6480)) xor (layer4_outputs(2327)));
    outputs(3074) <= layer4_outputs(379);
    outputs(3075) <= layer4_outputs(8737);
    outputs(3076) <= not(layer4_outputs(8431));
    outputs(3077) <= not(layer4_outputs(9032));
    outputs(3078) <= not(layer4_outputs(4646));
    outputs(3079) <= layer4_outputs(6182);
    outputs(3080) <= layer4_outputs(9763);
    outputs(3081) <= not((layer4_outputs(9867)) xor (layer4_outputs(118)));
    outputs(3082) <= layer4_outputs(9757);
    outputs(3083) <= not(layer4_outputs(3549));
    outputs(3084) <= not((layer4_outputs(320)) xor (layer4_outputs(9166)));
    outputs(3085) <= not(layer4_outputs(186));
    outputs(3086) <= layer4_outputs(7021);
    outputs(3087) <= not((layer4_outputs(49)) and (layer4_outputs(3224)));
    outputs(3088) <= (layer4_outputs(8935)) and (layer4_outputs(8700));
    outputs(3089) <= not((layer4_outputs(2991)) and (layer4_outputs(1896)));
    outputs(3090) <= layer4_outputs(3789);
    outputs(3091) <= not(layer4_outputs(5440));
    outputs(3092) <= layer4_outputs(8451);
    outputs(3093) <= layer4_outputs(4291);
    outputs(3094) <= not(layer4_outputs(4841));
    outputs(3095) <= not(layer4_outputs(9901));
    outputs(3096) <= layer4_outputs(9041);
    outputs(3097) <= not((layer4_outputs(9558)) and (layer4_outputs(6826)));
    outputs(3098) <= layer4_outputs(7853);
    outputs(3099) <= (layer4_outputs(7982)) xor (layer4_outputs(5449));
    outputs(3100) <= (layer4_outputs(2695)) xor (layer4_outputs(4983));
    outputs(3101) <= not(layer4_outputs(3646));
    outputs(3102) <= not(layer4_outputs(259));
    outputs(3103) <= not((layer4_outputs(4823)) xor (layer4_outputs(1200)));
    outputs(3104) <= not(layer4_outputs(4911));
    outputs(3105) <= layer4_outputs(4481);
    outputs(3106) <= not(layer4_outputs(2416));
    outputs(3107) <= not(layer4_outputs(10053));
    outputs(3108) <= layer4_outputs(473);
    outputs(3109) <= layer4_outputs(3813);
    outputs(3110) <= (layer4_outputs(9561)) xor (layer4_outputs(8332));
    outputs(3111) <= not((layer4_outputs(6337)) xor (layer4_outputs(5436)));
    outputs(3112) <= not((layer4_outputs(796)) and (layer4_outputs(6639)));
    outputs(3113) <= not(layer4_outputs(8417));
    outputs(3114) <= layer4_outputs(7230);
    outputs(3115) <= not(layer4_outputs(6004));
    outputs(3116) <= not((layer4_outputs(1180)) or (layer4_outputs(3498)));
    outputs(3117) <= not(layer4_outputs(6381)) or (layer4_outputs(5495));
    outputs(3118) <= not(layer4_outputs(3654));
    outputs(3119) <= (layer4_outputs(2039)) or (layer4_outputs(3890));
    outputs(3120) <= not(layer4_outputs(7622));
    outputs(3121) <= layer4_outputs(5390);
    outputs(3122) <= layer4_outputs(2884);
    outputs(3123) <= not(layer4_outputs(2144));
    outputs(3124) <= layer4_outputs(9228);
    outputs(3125) <= (layer4_outputs(5397)) xor (layer4_outputs(1102));
    outputs(3126) <= not(layer4_outputs(4971));
    outputs(3127) <= layer4_outputs(9134);
    outputs(3128) <= (layer4_outputs(8312)) xor (layer4_outputs(1412));
    outputs(3129) <= not((layer4_outputs(803)) xor (layer4_outputs(6837)));
    outputs(3130) <= layer4_outputs(7985);
    outputs(3131) <= not(layer4_outputs(6782));
    outputs(3132) <= (layer4_outputs(3233)) xor (layer4_outputs(2062));
    outputs(3133) <= (layer4_outputs(2692)) and not (layer4_outputs(1442));
    outputs(3134) <= layer4_outputs(4507);
    outputs(3135) <= layer4_outputs(5676);
    outputs(3136) <= layer4_outputs(3792);
    outputs(3137) <= layer4_outputs(9233);
    outputs(3138) <= not((layer4_outputs(4937)) xor (layer4_outputs(2135)));
    outputs(3139) <= (layer4_outputs(5747)) or (layer4_outputs(6766));
    outputs(3140) <= layer4_outputs(3509);
    outputs(3141) <= layer4_outputs(8890);
    outputs(3142) <= layer4_outputs(8994);
    outputs(3143) <= layer4_outputs(4724);
    outputs(3144) <= not(layer4_outputs(8763));
    outputs(3145) <= not((layer4_outputs(8555)) xor (layer4_outputs(3668)));
    outputs(3146) <= not((layer4_outputs(9455)) and (layer4_outputs(5627)));
    outputs(3147) <= not(layer4_outputs(6429));
    outputs(3148) <= (layer4_outputs(3698)) and (layer4_outputs(8441));
    outputs(3149) <= not((layer4_outputs(3739)) xor (layer4_outputs(10174)));
    outputs(3150) <= layer4_outputs(7161);
    outputs(3151) <= (layer4_outputs(9121)) xor (layer4_outputs(3902));
    outputs(3152) <= (layer4_outputs(7374)) and not (layer4_outputs(5577));
    outputs(3153) <= (layer4_outputs(4936)) and not (layer4_outputs(2664));
    outputs(3154) <= not(layer4_outputs(333));
    outputs(3155) <= layer4_outputs(9878);
    outputs(3156) <= not(layer4_outputs(3600));
    outputs(3157) <= layer4_outputs(9842);
    outputs(3158) <= layer4_outputs(2618);
    outputs(3159) <= not(layer4_outputs(6780));
    outputs(3160) <= layer4_outputs(8178);
    outputs(3161) <= layer4_outputs(3843);
    outputs(3162) <= (layer4_outputs(7608)) and not (layer4_outputs(7342));
    outputs(3163) <= (layer4_outputs(3910)) xor (layer4_outputs(2276));
    outputs(3164) <= (layer4_outputs(7616)) and not (layer4_outputs(6650));
    outputs(3165) <= layer4_outputs(3401);
    outputs(3166) <= layer4_outputs(9445);
    outputs(3167) <= not(layer4_outputs(1222)) or (layer4_outputs(8550));
    outputs(3168) <= not(layer4_outputs(9261));
    outputs(3169) <= not((layer4_outputs(1217)) or (layer4_outputs(8992)));
    outputs(3170) <= (layer4_outputs(2186)) and not (layer4_outputs(1167));
    outputs(3171) <= layer4_outputs(205);
    outputs(3172) <= not(layer4_outputs(278));
    outputs(3173) <= not(layer4_outputs(3064));
    outputs(3174) <= layer4_outputs(7892);
    outputs(3175) <= not(layer4_outputs(200));
    outputs(3176) <= not((layer4_outputs(8545)) xor (layer4_outputs(7396)));
    outputs(3177) <= (layer4_outputs(9626)) and not (layer4_outputs(3093));
    outputs(3178) <= not(layer4_outputs(5601));
    outputs(3179) <= layer4_outputs(2676);
    outputs(3180) <= layer4_outputs(1163);
    outputs(3181) <= not(layer4_outputs(7520));
    outputs(3182) <= layer4_outputs(8315);
    outputs(3183) <= not(layer4_outputs(8530)) or (layer4_outputs(1370));
    outputs(3184) <= not((layer4_outputs(2797)) and (layer4_outputs(7130)));
    outputs(3185) <= layer4_outputs(2088);
    outputs(3186) <= (layer4_outputs(4816)) xor (layer4_outputs(9242));
    outputs(3187) <= not(layer4_outputs(4010));
    outputs(3188) <= (layer4_outputs(6260)) and (layer4_outputs(2015));
    outputs(3189) <= not((layer4_outputs(705)) and (layer4_outputs(7778)));
    outputs(3190) <= not(layer4_outputs(7732));
    outputs(3191) <= layer4_outputs(1563);
    outputs(3192) <= layer4_outputs(3418);
    outputs(3193) <= not((layer4_outputs(2119)) xor (layer4_outputs(3665)));
    outputs(3194) <= (layer4_outputs(7229)) or (layer4_outputs(4430));
    outputs(3195) <= not((layer4_outputs(3991)) xor (layer4_outputs(4825)));
    outputs(3196) <= (layer4_outputs(2081)) xor (layer4_outputs(8256));
    outputs(3197) <= (layer4_outputs(576)) xor (layer4_outputs(9655));
    outputs(3198) <= not(layer4_outputs(5463));
    outputs(3199) <= not((layer4_outputs(3469)) xor (layer4_outputs(4336)));
    outputs(3200) <= (layer4_outputs(10125)) and not (layer4_outputs(4654));
    outputs(3201) <= layer4_outputs(986);
    outputs(3202) <= not(layer4_outputs(9263)) or (layer4_outputs(7663));
    outputs(3203) <= (layer4_outputs(1890)) xor (layer4_outputs(3845));
    outputs(3204) <= layer4_outputs(2909);
    outputs(3205) <= not(layer4_outputs(7498));
    outputs(3206) <= not((layer4_outputs(5585)) xor (layer4_outputs(6750)));
    outputs(3207) <= layer4_outputs(7035);
    outputs(3208) <= not((layer4_outputs(3632)) or (layer4_outputs(2464)));
    outputs(3209) <= not((layer4_outputs(9666)) xor (layer4_outputs(3588)));
    outputs(3210) <= not((layer4_outputs(1724)) or (layer4_outputs(6927)));
    outputs(3211) <= not(layer4_outputs(1599));
    outputs(3212) <= not((layer4_outputs(7718)) xor (layer4_outputs(9739)));
    outputs(3213) <= (layer4_outputs(9825)) xor (layer4_outputs(42));
    outputs(3214) <= not(layer4_outputs(1923));
    outputs(3215) <= not(layer4_outputs(7809));
    outputs(3216) <= layer4_outputs(1414);
    outputs(3217) <= layer4_outputs(837);
    outputs(3218) <= layer4_outputs(5624);
    outputs(3219) <= not(layer4_outputs(5662));
    outputs(3220) <= (layer4_outputs(8735)) xor (layer4_outputs(5892));
    outputs(3221) <= not(layer4_outputs(2920));
    outputs(3222) <= not(layer4_outputs(5598));
    outputs(3223) <= not(layer4_outputs(8649));
    outputs(3224) <= layer4_outputs(7495);
    outputs(3225) <= layer4_outputs(8230);
    outputs(3226) <= (layer4_outputs(9367)) xor (layer4_outputs(7216));
    outputs(3227) <= layer4_outputs(1495);
    outputs(3228) <= not(layer4_outputs(6362));
    outputs(3229) <= not(layer4_outputs(2760)) or (layer4_outputs(2897));
    outputs(3230) <= not((layer4_outputs(5927)) and (layer4_outputs(2473)));
    outputs(3231) <= (layer4_outputs(1748)) xor (layer4_outputs(6863));
    outputs(3232) <= (layer4_outputs(6661)) and not (layer4_outputs(9266));
    outputs(3233) <= not(layer4_outputs(376));
    outputs(3234) <= not((layer4_outputs(10086)) xor (layer4_outputs(3386)));
    outputs(3235) <= layer4_outputs(10144);
    outputs(3236) <= layer4_outputs(2771);
    outputs(3237) <= not(layer4_outputs(9219));
    outputs(3238) <= layer4_outputs(4432);
    outputs(3239) <= not(layer4_outputs(7824));
    outputs(3240) <= not(layer4_outputs(1312)) or (layer4_outputs(5772));
    outputs(3241) <= not(layer4_outputs(872));
    outputs(3242) <= layer4_outputs(236);
    outputs(3243) <= not((layer4_outputs(6241)) xor (layer4_outputs(9350)));
    outputs(3244) <= not(layer4_outputs(6782));
    outputs(3245) <= not((layer4_outputs(820)) xor (layer4_outputs(790)));
    outputs(3246) <= not(layer4_outputs(7607));
    outputs(3247) <= not(layer4_outputs(6569));
    outputs(3248) <= not(layer4_outputs(5142));
    outputs(3249) <= not(layer4_outputs(8766)) or (layer4_outputs(1716));
    outputs(3250) <= layer4_outputs(9733);
    outputs(3251) <= not(layer4_outputs(3462));
    outputs(3252) <= not(layer4_outputs(6282)) or (layer4_outputs(1877));
    outputs(3253) <= layer4_outputs(1541);
    outputs(3254) <= not(layer4_outputs(859));
    outputs(3255) <= not(layer4_outputs(878));
    outputs(3256) <= not(layer4_outputs(7968));
    outputs(3257) <= not((layer4_outputs(1620)) and (layer4_outputs(2204)));
    outputs(3258) <= not(layer4_outputs(9072));
    outputs(3259) <= not(layer4_outputs(3429));
    outputs(3260) <= (layer4_outputs(10176)) xor (layer4_outputs(2555));
    outputs(3261) <= not((layer4_outputs(2047)) xor (layer4_outputs(4251)));
    outputs(3262) <= (layer4_outputs(9433)) and (layer4_outputs(23));
    outputs(3263) <= not(layer4_outputs(1029));
    outputs(3264) <= layer4_outputs(3644);
    outputs(3265) <= not((layer4_outputs(9828)) xor (layer4_outputs(1283)));
    outputs(3266) <= (layer4_outputs(8688)) xor (layer4_outputs(7383));
    outputs(3267) <= not((layer4_outputs(7394)) xor (layer4_outputs(2288)));
    outputs(3268) <= layer4_outputs(5964);
    outputs(3269) <= not(layer4_outputs(6864));
    outputs(3270) <= layer4_outputs(5824);
    outputs(3271) <= not(layer4_outputs(10202)) or (layer4_outputs(7273));
    outputs(3272) <= layer4_outputs(1056);
    outputs(3273) <= layer4_outputs(2967);
    outputs(3274) <= not((layer4_outputs(1051)) or (layer4_outputs(1824)));
    outputs(3275) <= layer4_outputs(1787);
    outputs(3276) <= not(layer4_outputs(8172));
    outputs(3277) <= not(layer4_outputs(1050));
    outputs(3278) <= not(layer4_outputs(6212));
    outputs(3279) <= not((layer4_outputs(5714)) or (layer4_outputs(9111)));
    outputs(3280) <= not(layer4_outputs(2193));
    outputs(3281) <= not(layer4_outputs(6538));
    outputs(3282) <= not(layer4_outputs(619)) or (layer4_outputs(3734));
    outputs(3283) <= not((layer4_outputs(7991)) or (layer4_outputs(8745)));
    outputs(3284) <= not(layer4_outputs(2923));
    outputs(3285) <= not(layer4_outputs(2991));
    outputs(3286) <= not(layer4_outputs(9292));
    outputs(3287) <= not(layer4_outputs(9471));
    outputs(3288) <= not(layer4_outputs(3379));
    outputs(3289) <= not(layer4_outputs(1484));
    outputs(3290) <= not(layer4_outputs(4651));
    outputs(3291) <= not((layer4_outputs(5756)) xor (layer4_outputs(7333)));
    outputs(3292) <= layer4_outputs(1564);
    outputs(3293) <= layer4_outputs(4668);
    outputs(3294) <= layer4_outputs(8393);
    outputs(3295) <= (layer4_outputs(8761)) and not (layer4_outputs(6889));
    outputs(3296) <= layer4_outputs(7829);
    outputs(3297) <= (layer4_outputs(1327)) xor (layer4_outputs(750));
    outputs(3298) <= not((layer4_outputs(9579)) xor (layer4_outputs(9737)));
    outputs(3299) <= not(layer4_outputs(2236));
    outputs(3300) <= (layer4_outputs(3756)) and not (layer4_outputs(9819));
    outputs(3301) <= not(layer4_outputs(7360)) or (layer4_outputs(3686));
    outputs(3302) <= not((layer4_outputs(5044)) xor (layer4_outputs(4042)));
    outputs(3303) <= (layer4_outputs(6860)) or (layer4_outputs(2784));
    outputs(3304) <= layer4_outputs(2325);
    outputs(3305) <= (layer4_outputs(3253)) xor (layer4_outputs(6056));
    outputs(3306) <= not(layer4_outputs(1272));
    outputs(3307) <= layer4_outputs(7762);
    outputs(3308) <= not((layer4_outputs(6245)) xor (layer4_outputs(2121)));
    outputs(3309) <= layer4_outputs(9733);
    outputs(3310) <= not(layer4_outputs(4736));
    outputs(3311) <= (layer4_outputs(1026)) and (layer4_outputs(7848));
    outputs(3312) <= not(layer4_outputs(5647));
    outputs(3313) <= not(layer4_outputs(3191));
    outputs(3314) <= layer4_outputs(6537);
    outputs(3315) <= layer4_outputs(7911);
    outputs(3316) <= layer4_outputs(5659);
    outputs(3317) <= layer4_outputs(280);
    outputs(3318) <= not(layer4_outputs(1945));
    outputs(3319) <= not(layer4_outputs(6427));
    outputs(3320) <= not(layer4_outputs(4621));
    outputs(3321) <= not((layer4_outputs(5358)) or (layer4_outputs(8048)));
    outputs(3322) <= not(layer4_outputs(8450));
    outputs(3323) <= (layer4_outputs(3006)) and (layer4_outputs(7024));
    outputs(3324) <= (layer4_outputs(1310)) xor (layer4_outputs(9894));
    outputs(3325) <= layer4_outputs(5512);
    outputs(3326) <= not(layer4_outputs(1124));
    outputs(3327) <= not(layer4_outputs(5505));
    outputs(3328) <= layer4_outputs(4752);
    outputs(3329) <= not(layer4_outputs(2057));
    outputs(3330) <= layer4_outputs(362);
    outputs(3331) <= (layer4_outputs(5259)) xor (layer4_outputs(1767));
    outputs(3332) <= layer4_outputs(8114);
    outputs(3333) <= not((layer4_outputs(3036)) xor (layer4_outputs(3823)));
    outputs(3334) <= (layer4_outputs(5948)) xor (layer4_outputs(9440));
    outputs(3335) <= not(layer4_outputs(7560));
    outputs(3336) <= (layer4_outputs(4057)) xor (layer4_outputs(8965));
    outputs(3337) <= layer4_outputs(6583);
    outputs(3338) <= layer4_outputs(220);
    outputs(3339) <= not(layer4_outputs(8491));
    outputs(3340) <= not(layer4_outputs(8077));
    outputs(3341) <= layer4_outputs(4175);
    outputs(3342) <= not(layer4_outputs(331));
    outputs(3343) <= not(layer4_outputs(8180));
    outputs(3344) <= layer4_outputs(7850);
    outputs(3345) <= not(layer4_outputs(7352));
    outputs(3346) <= not(layer4_outputs(4135));
    outputs(3347) <= (layer4_outputs(2581)) or (layer4_outputs(982));
    outputs(3348) <= not(layer4_outputs(4863));
    outputs(3349) <= (layer4_outputs(3721)) xor (layer4_outputs(8396));
    outputs(3350) <= not((layer4_outputs(2477)) xor (layer4_outputs(1000)));
    outputs(3351) <= layer4_outputs(9431);
    outputs(3352) <= not(layer4_outputs(8082));
    outputs(3353) <= not(layer4_outputs(411));
    outputs(3354) <= layer4_outputs(9563);
    outputs(3355) <= not(layer4_outputs(2105));
    outputs(3356) <= not((layer4_outputs(6167)) xor (layer4_outputs(9049)));
    outputs(3357) <= not((layer4_outputs(5090)) xor (layer4_outputs(2726)));
    outputs(3358) <= not(layer4_outputs(9308)) or (layer4_outputs(4548));
    outputs(3359) <= (layer4_outputs(5697)) and not (layer4_outputs(2137));
    outputs(3360) <= not(layer4_outputs(6266));
    outputs(3361) <= (layer4_outputs(3538)) or (layer4_outputs(2052));
    outputs(3362) <= not((layer4_outputs(3128)) xor (layer4_outputs(924)));
    outputs(3363) <= layer4_outputs(354);
    outputs(3364) <= not((layer4_outputs(7507)) and (layer4_outputs(4574)));
    outputs(3365) <= (layer4_outputs(6793)) and not (layer4_outputs(1196));
    outputs(3366) <= (layer4_outputs(5242)) xor (layer4_outputs(4012));
    outputs(3367) <= not(layer4_outputs(5558));
    outputs(3368) <= layer4_outputs(769);
    outputs(3369) <= not(layer4_outputs(2321)) or (layer4_outputs(109));
    outputs(3370) <= not((layer4_outputs(9583)) xor (layer4_outputs(3349)));
    outputs(3371) <= not((layer4_outputs(5695)) xor (layer4_outputs(3114)));
    outputs(3372) <= (layer4_outputs(6235)) and not (layer4_outputs(1585));
    outputs(3373) <= layer4_outputs(2527);
    outputs(3374) <= not(layer4_outputs(90));
    outputs(3375) <= layer4_outputs(2889);
    outputs(3376) <= layer4_outputs(3673);
    outputs(3377) <= layer4_outputs(8254);
    outputs(3378) <= layer4_outputs(789);
    outputs(3379) <= '1';
    outputs(3380) <= not((layer4_outputs(1939)) xor (layer4_outputs(7559)));
    outputs(3381) <= not((layer4_outputs(5664)) xor (layer4_outputs(8)));
    outputs(3382) <= (layer4_outputs(5897)) xor (layer4_outputs(2529));
    outputs(3383) <= (layer4_outputs(5741)) xor (layer4_outputs(6130));
    outputs(3384) <= layer4_outputs(6317);
    outputs(3385) <= (layer4_outputs(190)) xor (layer4_outputs(3858));
    outputs(3386) <= not(layer4_outputs(3831));
    outputs(3387) <= layer4_outputs(6471);
    outputs(3388) <= not(layer4_outputs(5875));
    outputs(3389) <= layer4_outputs(222);
    outputs(3390) <= not(layer4_outputs(8190)) or (layer4_outputs(809));
    outputs(3391) <= layer4_outputs(1759);
    outputs(3392) <= (layer4_outputs(6260)) xor (layer4_outputs(4238));
    outputs(3393) <= not(layer4_outputs(2041));
    outputs(3394) <= layer4_outputs(6487);
    outputs(3395) <= layer4_outputs(9228);
    outputs(3396) <= not(layer4_outputs(8866));
    outputs(3397) <= not((layer4_outputs(4007)) xor (layer4_outputs(6294)));
    outputs(3398) <= layer4_outputs(8517);
    outputs(3399) <= layer4_outputs(579);
    outputs(3400) <= not((layer4_outputs(5670)) xor (layer4_outputs(8058)));
    outputs(3401) <= layer4_outputs(8333);
    outputs(3402) <= layer4_outputs(1780);
    outputs(3403) <= not(layer4_outputs(307));
    outputs(3404) <= (layer4_outputs(3257)) xor (layer4_outputs(9062));
    outputs(3405) <= layer4_outputs(8349);
    outputs(3406) <= layer4_outputs(5307);
    outputs(3407) <= not((layer4_outputs(9448)) or (layer4_outputs(6568)));
    outputs(3408) <= not(layer4_outputs(6150));
    outputs(3409) <= not((layer4_outputs(4649)) xor (layer4_outputs(8276)));
    outputs(3410) <= (layer4_outputs(1875)) and not (layer4_outputs(4854));
    outputs(3411) <= not(layer4_outputs(6948));
    outputs(3412) <= (layer4_outputs(1161)) and not (layer4_outputs(3254));
    outputs(3413) <= layer4_outputs(283);
    outputs(3414) <= not(layer4_outputs(1372));
    outputs(3415) <= (layer4_outputs(8830)) xor (layer4_outputs(2220));
    outputs(3416) <= not(layer4_outputs(5283));
    outputs(3417) <= (layer4_outputs(6038)) xor (layer4_outputs(1351));
    outputs(3418) <= layer4_outputs(6537);
    outputs(3419) <= not((layer4_outputs(1633)) xor (layer4_outputs(3126)));
    outputs(3420) <= not(layer4_outputs(4448));
    outputs(3421) <= layer4_outputs(4264);
    outputs(3422) <= not(layer4_outputs(3427));
    outputs(3423) <= not(layer4_outputs(1845));
    outputs(3424) <= not(layer4_outputs(815));
    outputs(3425) <= (layer4_outputs(908)) and not (layer4_outputs(7899));
    outputs(3426) <= not(layer4_outputs(9664));
    outputs(3427) <= layer4_outputs(7663);
    outputs(3428) <= layer4_outputs(9295);
    outputs(3429) <= not((layer4_outputs(403)) xor (layer4_outputs(7679)));
    outputs(3430) <= not(layer4_outputs(3689));
    outputs(3431) <= (layer4_outputs(1569)) xor (layer4_outputs(9027));
    outputs(3432) <= layer4_outputs(6628);
    outputs(3433) <= not(layer4_outputs(5720));
    outputs(3434) <= (layer4_outputs(8258)) or (layer4_outputs(1691));
    outputs(3435) <= layer4_outputs(7759);
    outputs(3436) <= not(layer4_outputs(1556));
    outputs(3437) <= layer4_outputs(849);
    outputs(3438) <= (layer4_outputs(1610)) and (layer4_outputs(9056));
    outputs(3439) <= not((layer4_outputs(9033)) or (layer4_outputs(9805)));
    outputs(3440) <= not(layer4_outputs(7573)) or (layer4_outputs(780));
    outputs(3441) <= not(layer4_outputs(9900));
    outputs(3442) <= layer4_outputs(7027);
    outputs(3443) <= not(layer4_outputs(6618));
    outputs(3444) <= layer4_outputs(3978);
    outputs(3445) <= not(layer4_outputs(8811));
    outputs(3446) <= not(layer4_outputs(474));
    outputs(3447) <= (layer4_outputs(2487)) xor (layer4_outputs(8543));
    outputs(3448) <= not(layer4_outputs(6363));
    outputs(3449) <= not(layer4_outputs(9210));
    outputs(3450) <= not(layer4_outputs(8588));
    outputs(3451) <= layer4_outputs(10121);
    outputs(3452) <= layer4_outputs(1581);
    outputs(3453) <= not(layer4_outputs(238));
    outputs(3454) <= not((layer4_outputs(7727)) xor (layer4_outputs(5913)));
    outputs(3455) <= not(layer4_outputs(9277));
    outputs(3456) <= (layer4_outputs(5829)) and (layer4_outputs(7911));
    outputs(3457) <= (layer4_outputs(4653)) xor (layer4_outputs(3313));
    outputs(3458) <= (layer4_outputs(5191)) and (layer4_outputs(8403));
    outputs(3459) <= not((layer4_outputs(2487)) or (layer4_outputs(6710)));
    outputs(3460) <= layer4_outputs(2621);
    outputs(3461) <= not(layer4_outputs(1523));
    outputs(3462) <= not(layer4_outputs(5204));
    outputs(3463) <= layer4_outputs(516);
    outputs(3464) <= not(layer4_outputs(1654)) or (layer4_outputs(513));
    outputs(3465) <= not(layer4_outputs(3926));
    outputs(3466) <= layer4_outputs(8551);
    outputs(3467) <= not((layer4_outputs(8362)) xor (layer4_outputs(7046)));
    outputs(3468) <= layer4_outputs(5010);
    outputs(3469) <= layer4_outputs(6236);
    outputs(3470) <= not(layer4_outputs(4118));
    outputs(3471) <= '1';
    outputs(3472) <= not(layer4_outputs(1013));
    outputs(3473) <= not(layer4_outputs(7138));
    outputs(3474) <= not((layer4_outputs(8483)) and (layer4_outputs(1951)));
    outputs(3475) <= not(layer4_outputs(2395));
    outputs(3476) <= layer4_outputs(5866);
    outputs(3477) <= not(layer4_outputs(6737));
    outputs(3478) <= layer4_outputs(2631);
    outputs(3479) <= layer4_outputs(9333);
    outputs(3480) <= not(layer4_outputs(3004));
    outputs(3481) <= '1';
    outputs(3482) <= not(layer4_outputs(3604));
    outputs(3483) <= (layer4_outputs(7115)) xor (layer4_outputs(2619));
    outputs(3484) <= not(layer4_outputs(4367));
    outputs(3485) <= not(layer4_outputs(2628));
    outputs(3486) <= layer4_outputs(6268);
    outputs(3487) <= layer4_outputs(6020);
    outputs(3488) <= not((layer4_outputs(4827)) xor (layer4_outputs(848)));
    outputs(3489) <= not(layer4_outputs(6693));
    outputs(3490) <= not(layer4_outputs(5401));
    outputs(3491) <= not(layer4_outputs(5315));
    outputs(3492) <= (layer4_outputs(6681)) xor (layer4_outputs(7804));
    outputs(3493) <= (layer4_outputs(413)) xor (layer4_outputs(10031));
    outputs(3494) <= (layer4_outputs(3028)) xor (layer4_outputs(5603));
    outputs(3495) <= layer4_outputs(500);
    outputs(3496) <= not((layer4_outputs(3498)) xor (layer4_outputs(5475)));
    outputs(3497) <= layer4_outputs(1649);
    outputs(3498) <= layer4_outputs(8969);
    outputs(3499) <= not(layer4_outputs(6823));
    outputs(3500) <= (layer4_outputs(2646)) xor (layer4_outputs(4845));
    outputs(3501) <= layer4_outputs(1034);
    outputs(3502) <= (layer4_outputs(4419)) and not (layer4_outputs(3426));
    outputs(3503) <= (layer4_outputs(1126)) xor (layer4_outputs(8181));
    outputs(3504) <= not(layer4_outputs(6104));
    outputs(3505) <= (layer4_outputs(3636)) xor (layer4_outputs(4300));
    outputs(3506) <= not((layer4_outputs(4161)) xor (layer4_outputs(812)));
    outputs(3507) <= not((layer4_outputs(821)) xor (layer4_outputs(3442)));
    outputs(3508) <= not((layer4_outputs(3326)) xor (layer4_outputs(2290)));
    outputs(3509) <= layer4_outputs(4756);
    outputs(3510) <= layer4_outputs(7193);
    outputs(3511) <= (layer4_outputs(4702)) and (layer4_outputs(6909));
    outputs(3512) <= layer4_outputs(2734);
    outputs(3513) <= not((layer4_outputs(1708)) or (layer4_outputs(977)));
    outputs(3514) <= layer4_outputs(5755);
    outputs(3515) <= (layer4_outputs(595)) or (layer4_outputs(8480));
    outputs(3516) <= not((layer4_outputs(6946)) xor (layer4_outputs(5292)));
    outputs(3517) <= not(layer4_outputs(5008));
    outputs(3518) <= not(layer4_outputs(4428));
    outputs(3519) <= layer4_outputs(8603);
    outputs(3520) <= (layer4_outputs(5395)) and (layer4_outputs(3210));
    outputs(3521) <= (layer4_outputs(4146)) xor (layer4_outputs(9443));
    outputs(3522) <= layer4_outputs(2368);
    outputs(3523) <= not(layer4_outputs(5765));
    outputs(3524) <= layer4_outputs(3134);
    outputs(3525) <= layer4_outputs(9486);
    outputs(3526) <= layer4_outputs(10094);
    outputs(3527) <= layer4_outputs(1669);
    outputs(3528) <= not((layer4_outputs(3308)) xor (layer4_outputs(4317)));
    outputs(3529) <= (layer4_outputs(1477)) xor (layer4_outputs(4371));
    outputs(3530) <= not(layer4_outputs(4439));
    outputs(3531) <= (layer4_outputs(8394)) and not (layer4_outputs(5005));
    outputs(3532) <= not(layer4_outputs(4160)) or (layer4_outputs(7016));
    outputs(3533) <= (layer4_outputs(8774)) or (layer4_outputs(927));
    outputs(3534) <= not(layer4_outputs(5123));
    outputs(3535) <= layer4_outputs(1894);
    outputs(3536) <= layer4_outputs(3392);
    outputs(3537) <= layer4_outputs(5702);
    outputs(3538) <= layer4_outputs(2257);
    outputs(3539) <= layer4_outputs(4868);
    outputs(3540) <= not(layer4_outputs(3359));
    outputs(3541) <= not(layer4_outputs(475));
    outputs(3542) <= not((layer4_outputs(3668)) and (layer4_outputs(1397)));
    outputs(3543) <= not(layer4_outputs(8383));
    outputs(3544) <= layer4_outputs(5249);
    outputs(3545) <= (layer4_outputs(1698)) xor (layer4_outputs(8725));
    outputs(3546) <= layer4_outputs(4115);
    outputs(3547) <= (layer4_outputs(9282)) and not (layer4_outputs(3689));
    outputs(3548) <= layer4_outputs(6711);
    outputs(3549) <= not(layer4_outputs(5732));
    outputs(3550) <= not(layer4_outputs(2181)) or (layer4_outputs(7554));
    outputs(3551) <= (layer4_outputs(9566)) or (layer4_outputs(1202));
    outputs(3552) <= not(layer4_outputs(2826));
    outputs(3553) <= layer4_outputs(220);
    outputs(3554) <= (layer4_outputs(6619)) xor (layer4_outputs(2456));
    outputs(3555) <= not(layer4_outputs(3479));
    outputs(3556) <= not((layer4_outputs(2276)) or (layer4_outputs(3184)));
    outputs(3557) <= not(layer4_outputs(9605));
    outputs(3558) <= layer4_outputs(3362);
    outputs(3559) <= layer4_outputs(4355);
    outputs(3560) <= layer4_outputs(5359);
    outputs(3561) <= not(layer4_outputs(4526));
    outputs(3562) <= not(layer4_outputs(8931));
    outputs(3563) <= not(layer4_outputs(8103));
    outputs(3564) <= not(layer4_outputs(4042));
    outputs(3565) <= layer4_outputs(7850);
    outputs(3566) <= not((layer4_outputs(1525)) and (layer4_outputs(8260)));
    outputs(3567) <= not((layer4_outputs(4918)) xor (layer4_outputs(6821)));
    outputs(3568) <= not(layer4_outputs(6692));
    outputs(3569) <= not(layer4_outputs(600));
    outputs(3570) <= not(layer4_outputs(10198)) or (layer4_outputs(8840));
    outputs(3571) <= (layer4_outputs(4324)) xor (layer4_outputs(8029));
    outputs(3572) <= layer4_outputs(4496);
    outputs(3573) <= not(layer4_outputs(4648));
    outputs(3574) <= layer4_outputs(5270);
    outputs(3575) <= not((layer4_outputs(2154)) xor (layer4_outputs(2972)));
    outputs(3576) <= not(layer4_outputs(10030));
    outputs(3577) <= layer4_outputs(7940);
    outputs(3578) <= not(layer4_outputs(7303));
    outputs(3579) <= layer4_outputs(2457);
    outputs(3580) <= layer4_outputs(7398);
    outputs(3581) <= layer4_outputs(9614);
    outputs(3582) <= layer4_outputs(9863);
    outputs(3583) <= not(layer4_outputs(6198));
    outputs(3584) <= (layer4_outputs(2717)) xor (layer4_outputs(8362));
    outputs(3585) <= (layer4_outputs(4848)) and not (layer4_outputs(717));
    outputs(3586) <= not(layer4_outputs(7658));
    outputs(3587) <= layer4_outputs(8451);
    outputs(3588) <= (layer4_outputs(5979)) and not (layer4_outputs(7919));
    outputs(3589) <= layer4_outputs(931);
    outputs(3590) <= layer4_outputs(433);
    outputs(3591) <= layer4_outputs(3961);
    outputs(3592) <= not((layer4_outputs(6655)) xor (layer4_outputs(3631)));
    outputs(3593) <= (layer4_outputs(2668)) and not (layer4_outputs(9595));
    outputs(3594) <= not(layer4_outputs(7071));
    outputs(3595) <= layer4_outputs(1385);
    outputs(3596) <= (layer4_outputs(9447)) xor (layer4_outputs(6770));
    outputs(3597) <= layer4_outputs(4932);
    outputs(3598) <= layer4_outputs(8547);
    outputs(3599) <= layer4_outputs(2950);
    outputs(3600) <= not(layer4_outputs(6571));
    outputs(3601) <= layer4_outputs(3937);
    outputs(3602) <= not(layer4_outputs(4424));
    outputs(3603) <= layer4_outputs(6010);
    outputs(3604) <= (layer4_outputs(2839)) and (layer4_outputs(4347));
    outputs(3605) <= not(layer4_outputs(8187)) or (layer4_outputs(7131));
    outputs(3606) <= (layer4_outputs(921)) xor (layer4_outputs(8147));
    outputs(3607) <= not((layer4_outputs(9139)) xor (layer4_outputs(3564)));
    outputs(3608) <= (layer4_outputs(8143)) or (layer4_outputs(2460));
    outputs(3609) <= not(layer4_outputs(9285));
    outputs(3610) <= (layer4_outputs(5602)) xor (layer4_outputs(8800));
    outputs(3611) <= not(layer4_outputs(3180)) or (layer4_outputs(651));
    outputs(3612) <= not(layer4_outputs(3556)) or (layer4_outputs(1859));
    outputs(3613) <= not(layer4_outputs(8968));
    outputs(3614) <= not(layer4_outputs(9137));
    outputs(3615) <= layer4_outputs(5679);
    outputs(3616) <= layer4_outputs(5677);
    outputs(3617) <= not(layer4_outputs(1291));
    outputs(3618) <= layer4_outputs(8499);
    outputs(3619) <= (layer4_outputs(5898)) and (layer4_outputs(6016));
    outputs(3620) <= not((layer4_outputs(8944)) xor (layer4_outputs(9410)));
    outputs(3621) <= (layer4_outputs(9101)) and not (layer4_outputs(2472));
    outputs(3622) <= not((layer4_outputs(5974)) and (layer4_outputs(1260)));
    outputs(3623) <= not(layer4_outputs(8351));
    outputs(3624) <= not(layer4_outputs(7162));
    outputs(3625) <= (layer4_outputs(5695)) xor (layer4_outputs(2892));
    outputs(3626) <= not((layer4_outputs(3732)) and (layer4_outputs(1366)));
    outputs(3627) <= layer4_outputs(7751);
    outputs(3628) <= not(layer4_outputs(6995));
    outputs(3629) <= layer4_outputs(3578);
    outputs(3630) <= (layer4_outputs(4922)) and not (layer4_outputs(923));
    outputs(3631) <= layer4_outputs(1908);
    outputs(3632) <= not(layer4_outputs(4874));
    outputs(3633) <= (layer4_outputs(6131)) xor (layer4_outputs(2653));
    outputs(3634) <= not(layer4_outputs(7090));
    outputs(3635) <= not(layer4_outputs(3447));
    outputs(3636) <= (layer4_outputs(5264)) xor (layer4_outputs(2303));
    outputs(3637) <= (layer4_outputs(9506)) xor (layer4_outputs(7391));
    outputs(3638) <= not(layer4_outputs(6945));
    outputs(3639) <= layer4_outputs(6191);
    outputs(3640) <= layer4_outputs(9181);
    outputs(3641) <= not(layer4_outputs(988));
    outputs(3642) <= layer4_outputs(10035);
    outputs(3643) <= not(layer4_outputs(8602));
    outputs(3644) <= not(layer4_outputs(4204));
    outputs(3645) <= not(layer4_outputs(5193));
    outputs(3646) <= (layer4_outputs(615)) xor (layer4_outputs(6398));
    outputs(3647) <= not(layer4_outputs(1066));
    outputs(3648) <= (layer4_outputs(659)) xor (layer4_outputs(9193));
    outputs(3649) <= layer4_outputs(189);
    outputs(3650) <= not(layer4_outputs(8845));
    outputs(3651) <= (layer4_outputs(5232)) and not (layer4_outputs(1651));
    outputs(3652) <= layer4_outputs(1010);
    outputs(3653) <= layer4_outputs(1584);
    outputs(3654) <= not(layer4_outputs(5897));
    outputs(3655) <= not((layer4_outputs(7425)) xor (layer4_outputs(7444)));
    outputs(3656) <= not((layer4_outputs(1981)) xor (layer4_outputs(894)));
    outputs(3657) <= not(layer4_outputs(2529)) or (layer4_outputs(566));
    outputs(3658) <= layer4_outputs(10085);
    outputs(3659) <= layer4_outputs(3268);
    outputs(3660) <= not(layer4_outputs(7195));
    outputs(3661) <= not(layer4_outputs(5842)) or (layer4_outputs(6989));
    outputs(3662) <= layer4_outputs(470);
    outputs(3663) <= layer4_outputs(4123);
    outputs(3664) <= not(layer4_outputs(8565)) or (layer4_outputs(9528));
    outputs(3665) <= not(layer4_outputs(8963)) or (layer4_outputs(2831));
    outputs(3666) <= (layer4_outputs(9007)) and not (layer4_outputs(5480));
    outputs(3667) <= not(layer4_outputs(9117));
    outputs(3668) <= not(layer4_outputs(4987));
    outputs(3669) <= not((layer4_outputs(608)) and (layer4_outputs(5241)));
    outputs(3670) <= not(layer4_outputs(9708));
    outputs(3671) <= (layer4_outputs(440)) or (layer4_outputs(9042));
    outputs(3672) <= layer4_outputs(2915);
    outputs(3673) <= not(layer4_outputs(9200)) or (layer4_outputs(2412));
    outputs(3674) <= not(layer4_outputs(9821));
    outputs(3675) <= not((layer4_outputs(3422)) and (layer4_outputs(7440)));
    outputs(3676) <= not(layer4_outputs(472));
    outputs(3677) <= not(layer4_outputs(612));
    outputs(3678) <= (layer4_outputs(8191)) xor (layer4_outputs(9553));
    outputs(3679) <= (layer4_outputs(7392)) and not (layer4_outputs(134));
    outputs(3680) <= (layer4_outputs(9399)) xor (layer4_outputs(4720));
    outputs(3681) <= layer4_outputs(2607);
    outputs(3682) <= not(layer4_outputs(458));
    outputs(3683) <= not(layer4_outputs(7192));
    outputs(3684) <= not(layer4_outputs(9116));
    outputs(3685) <= layer4_outputs(6232);
    outputs(3686) <= not((layer4_outputs(1200)) xor (layer4_outputs(4465)));
    outputs(3687) <= (layer4_outputs(9599)) xor (layer4_outputs(3815));
    outputs(3688) <= not((layer4_outputs(9592)) xor (layer4_outputs(9127)));
    outputs(3689) <= (layer4_outputs(5993)) and not (layer4_outputs(7459));
    outputs(3690) <= not(layer4_outputs(466));
    outputs(3691) <= not(layer4_outputs(1779));
    outputs(3692) <= (layer4_outputs(5426)) xor (layer4_outputs(2119));
    outputs(3693) <= not(layer4_outputs(7962));
    outputs(3694) <= not((layer4_outputs(2534)) or (layer4_outputs(5331)));
    outputs(3695) <= not(layer4_outputs(10003));
    outputs(3696) <= not(layer4_outputs(850));
    outputs(3697) <= (layer4_outputs(2338)) and not (layer4_outputs(7634));
    outputs(3698) <= not((layer4_outputs(550)) xor (layer4_outputs(126)));
    outputs(3699) <= layer4_outputs(8501);
    outputs(3700) <= not(layer4_outputs(330));
    outputs(3701) <= (layer4_outputs(561)) and not (layer4_outputs(5357));
    outputs(3702) <= layer4_outputs(6288);
    outputs(3703) <= not((layer4_outputs(3868)) xor (layer4_outputs(652)));
    outputs(3704) <= not((layer4_outputs(6067)) xor (layer4_outputs(54)));
    outputs(3705) <= not(layer4_outputs(511));
    outputs(3706) <= not(layer4_outputs(8094));
    outputs(3707) <= layer4_outputs(3178);
    outputs(3708) <= not(layer4_outputs(9740));
    outputs(3709) <= (layer4_outputs(5332)) and not (layer4_outputs(1710));
    outputs(3710) <= not((layer4_outputs(3268)) or (layer4_outputs(7528)));
    outputs(3711) <= not(layer4_outputs(8482));
    outputs(3712) <= not(layer4_outputs(5878));
    outputs(3713) <= not(layer4_outputs(720)) or (layer4_outputs(7862));
    outputs(3714) <= layer4_outputs(8682);
    outputs(3715) <= (layer4_outputs(4221)) or (layer4_outputs(447));
    outputs(3716) <= '0';
    outputs(3717) <= (layer4_outputs(89)) xor (layer4_outputs(1666));
    outputs(3718) <= not(layer4_outputs(6313)) or (layer4_outputs(967));
    outputs(3719) <= layer4_outputs(6010);
    outputs(3720) <= layer4_outputs(6845);
    outputs(3721) <= not(layer4_outputs(9060)) or (layer4_outputs(9158));
    outputs(3722) <= not(layer4_outputs(1997));
    outputs(3723) <= layer4_outputs(4570);
    outputs(3724) <= not(layer4_outputs(39));
    outputs(3725) <= layer4_outputs(4458);
    outputs(3726) <= layer4_outputs(3149);
    outputs(3727) <= not((layer4_outputs(5565)) xor (layer4_outputs(7591)));
    outputs(3728) <= layer4_outputs(917);
    outputs(3729) <= not(layer4_outputs(9815));
    outputs(3730) <= not((layer4_outputs(5076)) and (layer4_outputs(2261)));
    outputs(3731) <= not(layer4_outputs(1777)) or (layer4_outputs(2677));
    outputs(3732) <= not((layer4_outputs(10177)) xor (layer4_outputs(6838)));
    outputs(3733) <= (layer4_outputs(3957)) and not (layer4_outputs(967));
    outputs(3734) <= layer4_outputs(10178);
    outputs(3735) <= not((layer4_outputs(1002)) xor (layer4_outputs(193)));
    outputs(3736) <= not(layer4_outputs(9547));
    outputs(3737) <= layer4_outputs(10188);
    outputs(3738) <= not(layer4_outputs(6364)) or (layer4_outputs(7050));
    outputs(3739) <= layer4_outputs(1016);
    outputs(3740) <= not(layer4_outputs(1773));
    outputs(3741) <= layer4_outputs(7020);
    outputs(3742) <= layer4_outputs(1271);
    outputs(3743) <= layer4_outputs(7212);
    outputs(3744) <= not((layer4_outputs(8699)) xor (layer4_outputs(7165)));
    outputs(3745) <= layer4_outputs(2129);
    outputs(3746) <= layer4_outputs(624);
    outputs(3747) <= not(layer4_outputs(6207));
    outputs(3748) <= (layer4_outputs(7360)) or (layer4_outputs(5473));
    outputs(3749) <= (layer4_outputs(2059)) or (layer4_outputs(4159));
    outputs(3750) <= layer4_outputs(7558);
    outputs(3751) <= not(layer4_outputs(9456));
    outputs(3752) <= (layer4_outputs(2445)) xor (layer4_outputs(146));
    outputs(3753) <= not(layer4_outputs(7918));
    outputs(3754) <= not(layer4_outputs(4768)) or (layer4_outputs(5995));
    outputs(3755) <= (layer4_outputs(5744)) and not (layer4_outputs(7776));
    outputs(3756) <= not((layer4_outputs(9898)) or (layer4_outputs(6603)));
    outputs(3757) <= not(layer4_outputs(3370));
    outputs(3758) <= layer4_outputs(4859);
    outputs(3759) <= not((layer4_outputs(6825)) or (layer4_outputs(2585)));
    outputs(3760) <= not(layer4_outputs(9674)) or (layer4_outputs(2502));
    outputs(3761) <= not(layer4_outputs(2498));
    outputs(3762) <= layer4_outputs(1702);
    outputs(3763) <= not(layer4_outputs(9355));
    outputs(3764) <= not(layer4_outputs(9373));
    outputs(3765) <= not(layer4_outputs(5938));
    outputs(3766) <= (layer4_outputs(9650)) xor (layer4_outputs(7399));
    outputs(3767) <= layer4_outputs(5803);
    outputs(3768) <= layer4_outputs(9857);
    outputs(3769) <= (layer4_outputs(6341)) xor (layer4_outputs(7293));
    outputs(3770) <= not((layer4_outputs(4352)) xor (layer4_outputs(9432)));
    outputs(3771) <= layer4_outputs(9105);
    outputs(3772) <= not((layer4_outputs(326)) xor (layer4_outputs(4907)));
    outputs(3773) <= not(layer4_outputs(3310));
    outputs(3774) <= not((layer4_outputs(3217)) xor (layer4_outputs(9428)));
    outputs(3775) <= not(layer4_outputs(1024));
    outputs(3776) <= not((layer4_outputs(4730)) xor (layer4_outputs(4714)));
    outputs(3777) <= layer4_outputs(3821);
    outputs(3778) <= not(layer4_outputs(2428));
    outputs(3779) <= layer4_outputs(3733);
    outputs(3780) <= layer4_outputs(8352);
    outputs(3781) <= layer4_outputs(1009);
    outputs(3782) <= (layer4_outputs(3866)) xor (layer4_outputs(8312));
    outputs(3783) <= not((layer4_outputs(6328)) xor (layer4_outputs(1130)));
    outputs(3784) <= not(layer4_outputs(14));
    outputs(3785) <= not(layer4_outputs(1133));
    outputs(3786) <= layer4_outputs(4942);
    outputs(3787) <= (layer4_outputs(4)) xor (layer4_outputs(5324));
    outputs(3788) <= not(layer4_outputs(8829));
    outputs(3789) <= layer4_outputs(4074);
    outputs(3790) <= (layer4_outputs(5838)) and not (layer4_outputs(2326));
    outputs(3791) <= layer4_outputs(1143);
    outputs(3792) <= not((layer4_outputs(1144)) xor (layer4_outputs(2560)));
    outputs(3793) <= not(layer4_outputs(9009)) or (layer4_outputs(1281));
    outputs(3794) <= not(layer4_outputs(7214)) or (layer4_outputs(8462));
    outputs(3795) <= not((layer4_outputs(8116)) or (layer4_outputs(7709)));
    outputs(3796) <= not(layer4_outputs(6990));
    outputs(3797) <= layer4_outputs(9413);
    outputs(3798) <= layer4_outputs(6854);
    outputs(3799) <= layer4_outputs(110);
    outputs(3800) <= not(layer4_outputs(7280)) or (layer4_outputs(9854));
    outputs(3801) <= not(layer4_outputs(9067));
    outputs(3802) <= layer4_outputs(1518);
    outputs(3803) <= not(layer4_outputs(7074));
    outputs(3804) <= not((layer4_outputs(5703)) or (layer4_outputs(5912)));
    outputs(3805) <= not(layer4_outputs(3949));
    outputs(3806) <= (layer4_outputs(4203)) xor (layer4_outputs(1481));
    outputs(3807) <= not(layer4_outputs(2028));
    outputs(3808) <= layer4_outputs(6584);
    outputs(3809) <= layer4_outputs(1285);
    outputs(3810) <= not(layer4_outputs(4840));
    outputs(3811) <= layer4_outputs(9175);
    outputs(3812) <= layer4_outputs(7003);
    outputs(3813) <= not(layer4_outputs(3610));
    outputs(3814) <= not(layer4_outputs(2033));
    outputs(3815) <= not((layer4_outputs(519)) xor (layer4_outputs(7312)));
    outputs(3816) <= layer4_outputs(3910);
    outputs(3817) <= layer4_outputs(6877);
    outputs(3818) <= layer4_outputs(356);
    outputs(3819) <= (layer4_outputs(4008)) xor (layer4_outputs(2247));
    outputs(3820) <= not((layer4_outputs(3729)) xor (layer4_outputs(6111)));
    outputs(3821) <= layer4_outputs(9435);
    outputs(3822) <= (layer4_outputs(6573)) xor (layer4_outputs(6794));
    outputs(3823) <= layer4_outputs(7076);
    outputs(3824) <= not((layer4_outputs(1609)) or (layer4_outputs(9858)));
    outputs(3825) <= not((layer4_outputs(2769)) xor (layer4_outputs(4873)));
    outputs(3826) <= (layer4_outputs(3340)) and not (layer4_outputs(1201));
    outputs(3827) <= (layer4_outputs(6840)) xor (layer4_outputs(5799));
    outputs(3828) <= layer4_outputs(1505);
    outputs(3829) <= not(layer4_outputs(5787));
    outputs(3830) <= layer4_outputs(1937);
    outputs(3831) <= (layer4_outputs(3025)) and not (layer4_outputs(8430));
    outputs(3832) <= layer4_outputs(3186);
    outputs(3833) <= (layer4_outputs(3612)) or (layer4_outputs(6740));
    outputs(3834) <= (layer4_outputs(6892)) xor (layer4_outputs(148));
    outputs(3835) <= not(layer4_outputs(6341));
    outputs(3836) <= not(layer4_outputs(9035));
    outputs(3837) <= not(layer4_outputs(962));
    outputs(3838) <= layer4_outputs(9980);
    outputs(3839) <= (layer4_outputs(5833)) xor (layer4_outputs(8112));
    outputs(3840) <= (layer4_outputs(1489)) xor (layer4_outputs(5367));
    outputs(3841) <= (layer4_outputs(3195)) xor (layer4_outputs(4128));
    outputs(3842) <= layer4_outputs(6812);
    outputs(3843) <= layer4_outputs(4285);
    outputs(3844) <= layer4_outputs(7690);
    outputs(3845) <= layer4_outputs(2926);
    outputs(3846) <= not((layer4_outputs(501)) xor (layer4_outputs(7265)));
    outputs(3847) <= not(layer4_outputs(8137));
    outputs(3848) <= layer4_outputs(8958);
    outputs(3849) <= not(layer4_outputs(7456));
    outputs(3850) <= (layer4_outputs(2399)) xor (layer4_outputs(5424));
    outputs(3851) <= not(layer4_outputs(6475));
    outputs(3852) <= layer4_outputs(9509);
    outputs(3853) <= layer4_outputs(5783);
    outputs(3854) <= not(layer4_outputs(3173));
    outputs(3855) <= (layer4_outputs(2177)) and not (layer4_outputs(8620));
    outputs(3856) <= not((layer4_outputs(9835)) xor (layer4_outputs(2151)));
    outputs(3857) <= layer4_outputs(1544);
    outputs(3858) <= not(layer4_outputs(10198));
    outputs(3859) <= not(layer4_outputs(9465));
    outputs(3860) <= (layer4_outputs(7141)) xor (layer4_outputs(1771));
    outputs(3861) <= not((layer4_outputs(1317)) xor (layer4_outputs(1865)));
    outputs(3862) <= not((layer4_outputs(9617)) xor (layer4_outputs(7876)));
    outputs(3863) <= not((layer4_outputs(9486)) xor (layer4_outputs(310)));
    outputs(3864) <= layer4_outputs(7596);
    outputs(3865) <= not((layer4_outputs(1326)) xor (layer4_outputs(8336)));
    outputs(3866) <= not(layer4_outputs(902));
    outputs(3867) <= layer4_outputs(8334);
    outputs(3868) <= (layer4_outputs(8376)) xor (layer4_outputs(8795));
    outputs(3869) <= not(layer4_outputs(1653));
    outputs(3870) <= not(layer4_outputs(4545));
    outputs(3871) <= not((layer4_outputs(3694)) xor (layer4_outputs(4050)));
    outputs(3872) <= not(layer4_outputs(9551));
    outputs(3873) <= layer4_outputs(8953);
    outputs(3874) <= not(layer4_outputs(9232));
    outputs(3875) <= layer4_outputs(4607);
    outputs(3876) <= layer4_outputs(5509);
    outputs(3877) <= layer4_outputs(4089);
    outputs(3878) <= not(layer4_outputs(8862));
    outputs(3879) <= (layer4_outputs(2194)) or (layer4_outputs(8564));
    outputs(3880) <= (layer4_outputs(4710)) xor (layer4_outputs(894));
    outputs(3881) <= not((layer4_outputs(8152)) and (layer4_outputs(3140)));
    outputs(3882) <= not(layer4_outputs(2256));
    outputs(3883) <= not(layer4_outputs(7426));
    outputs(3884) <= layer4_outputs(9178);
    outputs(3885) <= layer4_outputs(1788);
    outputs(3886) <= not(layer4_outputs(2035));
    outputs(3887) <= (layer4_outputs(10188)) and (layer4_outputs(1492));
    outputs(3888) <= (layer4_outputs(5547)) xor (layer4_outputs(184));
    outputs(3889) <= (layer4_outputs(4028)) xor (layer4_outputs(1105));
    outputs(3890) <= not(layer4_outputs(6379));
    outputs(3891) <= not((layer4_outputs(5954)) xor (layer4_outputs(5797)));
    outputs(3892) <= not(layer4_outputs(8916));
    outputs(3893) <= not(layer4_outputs(8817));
    outputs(3894) <= layer4_outputs(7790);
    outputs(3895) <= layer4_outputs(15);
    outputs(3896) <= (layer4_outputs(8653)) and (layer4_outputs(10080));
    outputs(3897) <= layer4_outputs(8595);
    outputs(3898) <= layer4_outputs(7669);
    outputs(3899) <= layer4_outputs(4705);
    outputs(3900) <= (layer4_outputs(4085)) and not (layer4_outputs(4418));
    outputs(3901) <= not((layer4_outputs(8144)) or (layer4_outputs(3872)));
    outputs(3902) <= not(layer4_outputs(8605));
    outputs(3903) <= layer4_outputs(2967);
    outputs(3904) <= layer4_outputs(5001);
    outputs(3905) <= layer4_outputs(1318);
    outputs(3906) <= (layer4_outputs(2344)) xor (layer4_outputs(4249));
    outputs(3907) <= not(layer4_outputs(1762));
    outputs(3908) <= not(layer4_outputs(1665));
    outputs(3909) <= (layer4_outputs(10219)) xor (layer4_outputs(38));
    outputs(3910) <= (layer4_outputs(5870)) xor (layer4_outputs(5669));
    outputs(3911) <= (layer4_outputs(7339)) or (layer4_outputs(6461));
    outputs(3912) <= (layer4_outputs(7176)) xor (layer4_outputs(1936));
    outputs(3913) <= not(layer4_outputs(6194));
    outputs(3914) <= layer4_outputs(1603);
    outputs(3915) <= layer4_outputs(4237);
    outputs(3916) <= (layer4_outputs(9668)) or (layer4_outputs(1431));
    outputs(3917) <= layer4_outputs(3875);
    outputs(3918) <= not(layer4_outputs(6169));
    outputs(3919) <= (layer4_outputs(7001)) xor (layer4_outputs(7025));
    outputs(3920) <= layer4_outputs(2410);
    outputs(3921) <= (layer4_outputs(4298)) or (layer4_outputs(7571));
    outputs(3922) <= not((layer4_outputs(7782)) xor (layer4_outputs(2731)));
    outputs(3923) <= not(layer4_outputs(4661));
    outputs(3924) <= layer4_outputs(5088);
    outputs(3925) <= layer4_outputs(6651);
    outputs(3926) <= not(layer4_outputs(1887));
    outputs(3927) <= not(layer4_outputs(7609));
    outputs(3928) <= not(layer4_outputs(4566));
    outputs(3929) <= layer4_outputs(3344);
    outputs(3930) <= layer4_outputs(8996);
    outputs(3931) <= layer4_outputs(4524);
    outputs(3932) <= layer4_outputs(974);
    outputs(3933) <= not((layer4_outputs(7671)) xor (layer4_outputs(1012)));
    outputs(3934) <= layer4_outputs(1796);
    outputs(3935) <= not(layer4_outputs(2225));
    outputs(3936) <= layer4_outputs(450);
    outputs(3937) <= layer4_outputs(6877);
    outputs(3938) <= layer4_outputs(891);
    outputs(3939) <= layer4_outputs(10040);
    outputs(3940) <= (layer4_outputs(1805)) xor (layer4_outputs(9144));
    outputs(3941) <= not(layer4_outputs(5765));
    outputs(3942) <= not((layer4_outputs(3190)) xor (layer4_outputs(7188)));
    outputs(3943) <= not(layer4_outputs(6515));
    outputs(3944) <= not((layer4_outputs(6936)) xor (layer4_outputs(9176)));
    outputs(3945) <= layer4_outputs(9786);
    outputs(3946) <= not(layer4_outputs(10112));
    outputs(3947) <= not(layer4_outputs(10076));
    outputs(3948) <= layer4_outputs(8808);
    outputs(3949) <= layer4_outputs(2293);
    outputs(3950) <= not(layer4_outputs(9619));
    outputs(3951) <= not(layer4_outputs(4070));
    outputs(3952) <= not(layer4_outputs(3635));
    outputs(3953) <= (layer4_outputs(3350)) xor (layer4_outputs(8270));
    outputs(3954) <= not(layer4_outputs(9671)) or (layer4_outputs(6115));
    outputs(3955) <= layer4_outputs(2031);
    outputs(3956) <= (layer4_outputs(7908)) and not (layer4_outputs(8894));
    outputs(3957) <= (layer4_outputs(7083)) xor (layer4_outputs(352));
    outputs(3958) <= layer4_outputs(2054);
    outputs(3959) <= layer4_outputs(2590);
    outputs(3960) <= not(layer4_outputs(7548));
    outputs(3961) <= not((layer4_outputs(3975)) xor (layer4_outputs(9702)));
    outputs(3962) <= (layer4_outputs(4732)) xor (layer4_outputs(7782));
    outputs(3963) <= (layer4_outputs(1080)) and (layer4_outputs(4053));
    outputs(3964) <= not(layer4_outputs(8167));
    outputs(3965) <= layer4_outputs(5316);
    outputs(3966) <= not(layer4_outputs(1652));
    outputs(3967) <= (layer4_outputs(2984)) and not (layer4_outputs(7638));
    outputs(3968) <= layer4_outputs(8282);
    outputs(3969) <= layer4_outputs(4340);
    outputs(3970) <= layer4_outputs(8304);
    outputs(3971) <= layer4_outputs(9049);
    outputs(3972) <= not(layer4_outputs(7704));
    outputs(3973) <= layer4_outputs(1705);
    outputs(3974) <= not(layer4_outputs(6374)) or (layer4_outputs(3403));
    outputs(3975) <= layer4_outputs(8440);
    outputs(3976) <= (layer4_outputs(2090)) and (layer4_outputs(10010));
    outputs(3977) <= not(layer4_outputs(8461)) or (layer4_outputs(26));
    outputs(3978) <= not(layer4_outputs(1191));
    outputs(3979) <= (layer4_outputs(5959)) and not (layer4_outputs(9704));
    outputs(3980) <= layer4_outputs(3083);
    outputs(3981) <= not(layer4_outputs(7716));
    outputs(3982) <= (layer4_outputs(4811)) xor (layer4_outputs(816));
    outputs(3983) <= layer4_outputs(6795);
    outputs(3984) <= (layer4_outputs(4663)) xor (layer4_outputs(8077));
    outputs(3985) <= not(layer4_outputs(9444));
    outputs(3986) <= not(layer4_outputs(8733));
    outputs(3987) <= (layer4_outputs(5784)) and not (layer4_outputs(6379));
    outputs(3988) <= (layer4_outputs(9834)) xor (layer4_outputs(2157));
    outputs(3989) <= not((layer4_outputs(5994)) xor (layer4_outputs(8986)));
    outputs(3990) <= layer4_outputs(5184);
    outputs(3991) <= layer4_outputs(4671);
    outputs(3992) <= (layer4_outputs(1008)) xor (layer4_outputs(5904));
    outputs(3993) <= (layer4_outputs(5618)) xor (layer4_outputs(6690));
    outputs(3994) <= not(layer4_outputs(10102));
    outputs(3995) <= not((layer4_outputs(2723)) or (layer4_outputs(5616)));
    outputs(3996) <= not(layer4_outputs(2946)) or (layer4_outputs(1528));
    outputs(3997) <= not((layer4_outputs(6851)) xor (layer4_outputs(3841)));
    outputs(3998) <= not(layer4_outputs(2285));
    outputs(3999) <= not(layer4_outputs(9983));
    outputs(4000) <= layer4_outputs(9041);
    outputs(4001) <= layer4_outputs(2115);
    outputs(4002) <= not((layer4_outputs(638)) xor (layer4_outputs(5208)));
    outputs(4003) <= not(layer4_outputs(6887)) or (layer4_outputs(995));
    outputs(4004) <= '1';
    outputs(4005) <= layer4_outputs(4472);
    outputs(4006) <= not(layer4_outputs(7725)) or (layer4_outputs(7649));
    outputs(4007) <= not((layer4_outputs(3022)) xor (layer4_outputs(8182)));
    outputs(4008) <= (layer4_outputs(5281)) or (layer4_outputs(6772));
    outputs(4009) <= not(layer4_outputs(7746)) or (layer4_outputs(1411));
    outputs(4010) <= (layer4_outputs(7866)) xor (layer4_outputs(6284));
    outputs(4011) <= (layer4_outputs(229)) xor (layer4_outputs(4224));
    outputs(4012) <= not(layer4_outputs(8593));
    outputs(4013) <= not((layer4_outputs(7822)) xor (layer4_outputs(4192)));
    outputs(4014) <= (layer4_outputs(6019)) xor (layer4_outputs(4760));
    outputs(4015) <= layer4_outputs(2346);
    outputs(4016) <= not(layer4_outputs(7739));
    outputs(4017) <= layer4_outputs(4501);
    outputs(4018) <= layer4_outputs(4462);
    outputs(4019) <= layer4_outputs(6161);
    outputs(4020) <= (layer4_outputs(3376)) xor (layer4_outputs(4336));
    outputs(4021) <= (layer4_outputs(8193)) xor (layer4_outputs(4993));
    outputs(4022) <= layer4_outputs(7779);
    outputs(4023) <= layer4_outputs(7596);
    outputs(4024) <= (layer4_outputs(3753)) xor (layer4_outputs(2296));
    outputs(4025) <= (layer4_outputs(7402)) xor (layer4_outputs(8095));
    outputs(4026) <= layer4_outputs(5066);
    outputs(4027) <= layer4_outputs(65);
    outputs(4028) <= not((layer4_outputs(4213)) and (layer4_outputs(1613)));
    outputs(4029) <= layer4_outputs(2384);
    outputs(4030) <= (layer4_outputs(5976)) xor (layer4_outputs(9418));
    outputs(4031) <= layer4_outputs(4175);
    outputs(4032) <= (layer4_outputs(8342)) and (layer4_outputs(3499));
    outputs(4033) <= layer4_outputs(1500);
    outputs(4034) <= (layer4_outputs(3718)) and (layer4_outputs(5431));
    outputs(4035) <= layer4_outputs(9533);
    outputs(4036) <= not(layer4_outputs(6210));
    outputs(4037) <= layer4_outputs(8936);
    outputs(4038) <= layer4_outputs(5877);
    outputs(4039) <= layer4_outputs(703);
    outputs(4040) <= not(layer4_outputs(9631));
    outputs(4041) <= (layer4_outputs(8121)) and (layer4_outputs(6790));
    outputs(4042) <= not(layer4_outputs(7384));
    outputs(4043) <= not(layer4_outputs(8520)) or (layer4_outputs(485));
    outputs(4044) <= (layer4_outputs(5085)) xor (layer4_outputs(7368));
    outputs(4045) <= not(layer4_outputs(7921));
    outputs(4046) <= not(layer4_outputs(1664)) or (layer4_outputs(4254));
    outputs(4047) <= layer4_outputs(5206);
    outputs(4048) <= not(layer4_outputs(3153));
    outputs(4049) <= layer4_outputs(2011);
    outputs(4050) <= not((layer4_outputs(6801)) xor (layer4_outputs(2289)));
    outputs(4051) <= (layer4_outputs(4016)) and not (layer4_outputs(4041));
    outputs(4052) <= layer4_outputs(9531);
    outputs(4053) <= layer4_outputs(7677);
    outputs(4054) <= '0';
    outputs(4055) <= layer4_outputs(5072);
    outputs(4056) <= (layer4_outputs(459)) xor (layer4_outputs(5450));
    outputs(4057) <= not(layer4_outputs(7709));
    outputs(4058) <= layer4_outputs(3295);
    outputs(4059) <= not(layer4_outputs(176));
    outputs(4060) <= (layer4_outputs(6285)) and not (layer4_outputs(6858));
    outputs(4061) <= (layer4_outputs(4099)) and not (layer4_outputs(1579));
    outputs(4062) <= not(layer4_outputs(10185));
    outputs(4063) <= (layer4_outputs(7543)) xor (layer4_outputs(297));
    outputs(4064) <= layer4_outputs(9001);
    outputs(4065) <= layer4_outputs(211);
    outputs(4066) <= layer4_outputs(5236);
    outputs(4067) <= layer4_outputs(1633);
    outputs(4068) <= not(layer4_outputs(3660));
    outputs(4069) <= not(layer4_outputs(5048));
    outputs(4070) <= (layer4_outputs(4307)) xor (layer4_outputs(6244));
    outputs(4071) <= layer4_outputs(8225);
    outputs(4072) <= layer4_outputs(885);
    outputs(4073) <= (layer4_outputs(8548)) or (layer4_outputs(6574));
    outputs(4074) <= not(layer4_outputs(7797));
    outputs(4075) <= layer4_outputs(2682);
    outputs(4076) <= not(layer4_outputs(3929));
    outputs(4077) <= (layer4_outputs(4360)) and not (layer4_outputs(6251));
    outputs(4078) <= not((layer4_outputs(2238)) xor (layer4_outputs(6483)));
    outputs(4079) <= layer4_outputs(7831);
    outputs(4080) <= (layer4_outputs(8838)) xor (layer4_outputs(6679));
    outputs(4081) <= layer4_outputs(9786);
    outputs(4082) <= not(layer4_outputs(2243));
    outputs(4083) <= not(layer4_outputs(6167)) or (layer4_outputs(5032));
    outputs(4084) <= layer4_outputs(9684);
    outputs(4085) <= not(layer4_outputs(9086));
    outputs(4086) <= not((layer4_outputs(6900)) or (layer4_outputs(639)));
    outputs(4087) <= not(layer4_outputs(1129));
    outputs(4088) <= not(layer4_outputs(2482));
    outputs(4089) <= not(layer4_outputs(6266));
    outputs(4090) <= layer4_outputs(4130);
    outputs(4091) <= not(layer4_outputs(2573));
    outputs(4092) <= (layer4_outputs(4410)) xor (layer4_outputs(6067));
    outputs(4093) <= layer4_outputs(9548);
    outputs(4094) <= not(layer4_outputs(1128));
    outputs(4095) <= not((layer4_outputs(165)) xor (layer4_outputs(7236)));
    outputs(4096) <= layer4_outputs(1082);
    outputs(4097) <= (layer4_outputs(3949)) xor (layer4_outputs(1628));
    outputs(4098) <= not(layer4_outputs(8274));
    outputs(4099) <= layer4_outputs(3513);
    outputs(4100) <= layer4_outputs(3039);
    outputs(4101) <= not(layer4_outputs(5902));
    outputs(4102) <= not(layer4_outputs(2106));
    outputs(4103) <= (layer4_outputs(452)) and not (layer4_outputs(1844));
    outputs(4104) <= not(layer4_outputs(5534));
    outputs(4105) <= layer4_outputs(6472);
    outputs(4106) <= not(layer4_outputs(920));
    outputs(4107) <= not(layer4_outputs(5456));
    outputs(4108) <= not((layer4_outputs(4563)) xor (layer4_outputs(10137)));
    outputs(4109) <= (layer4_outputs(188)) xor (layer4_outputs(8066));
    outputs(4110) <= (layer4_outputs(9030)) and not (layer4_outputs(9112));
    outputs(4111) <= (layer4_outputs(387)) and not (layer4_outputs(3573));
    outputs(4112) <= not((layer4_outputs(8218)) and (layer4_outputs(4332)));
    outputs(4113) <= (layer4_outputs(3562)) xor (layer4_outputs(5626));
    outputs(4114) <= layer4_outputs(1395);
    outputs(4115) <= not((layer4_outputs(1048)) xor (layer4_outputs(5864)));
    outputs(4116) <= not(layer4_outputs(3508));
    outputs(4117) <= not(layer4_outputs(8810));
    outputs(4118) <= not(layer4_outputs(3776));
    outputs(4119) <= layer4_outputs(4396);
    outputs(4120) <= (layer4_outputs(2993)) and (layer4_outputs(2674));
    outputs(4121) <= not(layer4_outputs(5804));
    outputs(4122) <= not(layer4_outputs(8361));
    outputs(4123) <= not(layer4_outputs(8476));
    outputs(4124) <= layer4_outputs(5089);
    outputs(4125) <= layer4_outputs(3442);
    outputs(4126) <= (layer4_outputs(9195)) xor (layer4_outputs(3708));
    outputs(4127) <= layer4_outputs(6085);
    outputs(4128) <= layer4_outputs(6895);
    outputs(4129) <= not((layer4_outputs(9040)) xor (layer4_outputs(6291)));
    outputs(4130) <= (layer4_outputs(8979)) xor (layer4_outputs(299));
    outputs(4131) <= layer4_outputs(2136);
    outputs(4132) <= (layer4_outputs(7533)) and not (layer4_outputs(436));
    outputs(4133) <= layer4_outputs(5238);
    outputs(4134) <= not((layer4_outputs(3643)) xor (layer4_outputs(2377)));
    outputs(4135) <= not(layer4_outputs(853));
    outputs(4136) <= layer4_outputs(4707);
    outputs(4137) <= layer4_outputs(5567);
    outputs(4138) <= not(layer4_outputs(3449));
    outputs(4139) <= not(layer4_outputs(2599));
    outputs(4140) <= not(layer4_outputs(4781));
    outputs(4141) <= (layer4_outputs(9853)) or (layer4_outputs(7506));
    outputs(4142) <= (layer4_outputs(8671)) xor (layer4_outputs(1271));
    outputs(4143) <= (layer4_outputs(1279)) xor (layer4_outputs(913));
    outputs(4144) <= not(layer4_outputs(679));
    outputs(4145) <= (layer4_outputs(627)) xor (layer4_outputs(2942));
    outputs(4146) <= not(layer4_outputs(8353));
    outputs(4147) <= (layer4_outputs(1114)) xor (layer4_outputs(8158));
    outputs(4148) <= not(layer4_outputs(5419));
    outputs(4149) <= layer4_outputs(8618);
    outputs(4150) <= not((layer4_outputs(552)) xor (layer4_outputs(9072)));
    outputs(4151) <= layer4_outputs(5349);
    outputs(4152) <= (layer4_outputs(1963)) xor (layer4_outputs(5933));
    outputs(4153) <= layer4_outputs(9095);
    outputs(4154) <= not(layer4_outputs(7775));
    outputs(4155) <= not(layer4_outputs(574)) or (layer4_outputs(4886));
    outputs(4156) <= not(layer4_outputs(3072));
    outputs(4157) <= not(layer4_outputs(1590));
    outputs(4158) <= not(layer4_outputs(520));
    outputs(4159) <= not(layer4_outputs(8862));
    outputs(4160) <= not((layer4_outputs(8125)) xor (layer4_outputs(7602)));
    outputs(4161) <= not(layer4_outputs(3766));
    outputs(4162) <= layer4_outputs(131);
    outputs(4163) <= not(layer4_outputs(8684));
    outputs(4164) <= not((layer4_outputs(9457)) xor (layer4_outputs(9162)));
    outputs(4165) <= not(layer4_outputs(7660));
    outputs(4166) <= not(layer4_outputs(8923));
    outputs(4167) <= layer4_outputs(5886);
    outputs(4168) <= (layer4_outputs(6674)) xor (layer4_outputs(8661));
    outputs(4169) <= (layer4_outputs(4807)) or (layer4_outputs(5020));
    outputs(4170) <= not((layer4_outputs(2597)) xor (layer4_outputs(9699)));
    outputs(4171) <= not(layer4_outputs(9286));
    outputs(4172) <= layer4_outputs(7183);
    outputs(4173) <= layer4_outputs(3996);
    outputs(4174) <= (layer4_outputs(714)) xor (layer4_outputs(9340));
    outputs(4175) <= not(layer4_outputs(332));
    outputs(4176) <= layer4_outputs(7064);
    outputs(4177) <= (layer4_outputs(2945)) xor (layer4_outputs(3372));
    outputs(4178) <= not(layer4_outputs(3186));
    outputs(4179) <= not(layer4_outputs(7408));
    outputs(4180) <= not(layer4_outputs(5905));
    outputs(4181) <= not(layer4_outputs(9404));
    outputs(4182) <= layer4_outputs(3099);
    outputs(4183) <= layer4_outputs(8287);
    outputs(4184) <= not((layer4_outputs(5791)) xor (layer4_outputs(631)));
    outputs(4185) <= not((layer4_outputs(7101)) xor (layer4_outputs(1638)));
    outputs(4186) <= (layer4_outputs(2470)) xor (layer4_outputs(6322));
    outputs(4187) <= not(layer4_outputs(9278));
    outputs(4188) <= layer4_outputs(2856);
    outputs(4189) <= not(layer4_outputs(3060));
    outputs(4190) <= not((layer4_outputs(2684)) and (layer4_outputs(4932)));
    outputs(4191) <= (layer4_outputs(1040)) and not (layer4_outputs(8757));
    outputs(4192) <= (layer4_outputs(756)) xor (layer4_outputs(5047));
    outputs(4193) <= not((layer4_outputs(9467)) and (layer4_outputs(4902)));
    outputs(4194) <= not(layer4_outputs(2124));
    outputs(4195) <= (layer4_outputs(4239)) and (layer4_outputs(4141));
    outputs(4196) <= (layer4_outputs(4667)) xor (layer4_outputs(1006));
    outputs(4197) <= not(layer4_outputs(3226));
    outputs(4198) <= not((layer4_outputs(4614)) xor (layer4_outputs(7101)));
    outputs(4199) <= (layer4_outputs(7072)) xor (layer4_outputs(2458));
    outputs(4200) <= (layer4_outputs(2700)) and not (layer4_outputs(4944));
    outputs(4201) <= layer4_outputs(1943);
    outputs(4202) <= layer4_outputs(5153);
    outputs(4203) <= not(layer4_outputs(5494));
    outputs(4204) <= layer4_outputs(5724);
    outputs(4205) <= not(layer4_outputs(1059));
    outputs(4206) <= layer4_outputs(9747);
    outputs(4207) <= not(layer4_outputs(5960));
    outputs(4208) <= layer4_outputs(3032);
    outputs(4209) <= layer4_outputs(6079);
    outputs(4210) <= layer4_outputs(4158);
    outputs(4211) <= layer4_outputs(8777);
    outputs(4212) <= (layer4_outputs(2905)) or (layer4_outputs(9455));
    outputs(4213) <= layer4_outputs(4976);
    outputs(4214) <= '1';
    outputs(4215) <= not((layer4_outputs(4754)) or (layer4_outputs(4471)));
    outputs(4216) <= layer4_outputs(1974);
    outputs(4217) <= not(layer4_outputs(7665));
    outputs(4218) <= (layer4_outputs(2899)) and not (layer4_outputs(3098));
    outputs(4219) <= layer4_outputs(8978);
    outputs(4220) <= layer4_outputs(3221);
    outputs(4221) <= not(layer4_outputs(739));
    outputs(4222) <= layer4_outputs(2285);
    outputs(4223) <= not(layer4_outputs(3693));
    outputs(4224) <= layer4_outputs(1057);
    outputs(4225) <= layer4_outputs(3759);
    outputs(4226) <= not((layer4_outputs(4005)) xor (layer4_outputs(3691)));
    outputs(4227) <= layer4_outputs(6898);
    outputs(4228) <= not(layer4_outputs(4520));
    outputs(4229) <= not((layer4_outputs(1393)) xor (layer4_outputs(6240)));
    outputs(4230) <= layer4_outputs(357);
    outputs(4231) <= not(layer4_outputs(1604));
    outputs(4232) <= not(layer4_outputs(6795));
    outputs(4233) <= (layer4_outputs(5428)) and not (layer4_outputs(4430));
    outputs(4234) <= not((layer4_outputs(1515)) xor (layer4_outputs(8405)));
    outputs(4235) <= not((layer4_outputs(7747)) xor (layer4_outputs(2125)));
    outputs(4236) <= not((layer4_outputs(837)) xor (layer4_outputs(2494)));
    outputs(4237) <= not(layer4_outputs(4951));
    outputs(4238) <= (layer4_outputs(811)) and (layer4_outputs(2786));
    outputs(4239) <= (layer4_outputs(2231)) xor (layer4_outputs(7301));
    outputs(4240) <= not(layer4_outputs(8937));
    outputs(4241) <= layer4_outputs(2562);
    outputs(4242) <= (layer4_outputs(2328)) and not (layer4_outputs(3339));
    outputs(4243) <= layer4_outputs(9167);
    outputs(4244) <= not(layer4_outputs(3219)) or (layer4_outputs(8537));
    outputs(4245) <= not(layer4_outputs(6494));
    outputs(4246) <= layer4_outputs(2740);
    outputs(4247) <= not((layer4_outputs(8355)) xor (layer4_outputs(4090)));
    outputs(4248) <= not(layer4_outputs(6980));
    outputs(4249) <= not(layer4_outputs(8390));
    outputs(4250) <= not(layer4_outputs(7902));
    outputs(4251) <= (layer4_outputs(9674)) and not (layer4_outputs(2540));
    outputs(4252) <= layer4_outputs(6221);
    outputs(4253) <= layer4_outputs(9200);
    outputs(4254) <= not(layer4_outputs(3014));
    outputs(4255) <= not(layer4_outputs(2904));
    outputs(4256) <= (layer4_outputs(7968)) xor (layer4_outputs(3683));
    outputs(4257) <= layer4_outputs(3921);
    outputs(4258) <= not(layer4_outputs(6068));
    outputs(4259) <= not((layer4_outputs(8028)) xor (layer4_outputs(272)));
    outputs(4260) <= layer4_outputs(9576);
    outputs(4261) <= not(layer4_outputs(3230));
    outputs(4262) <= layer4_outputs(3559);
    outputs(4263) <= not((layer4_outputs(2414)) xor (layer4_outputs(8378)));
    outputs(4264) <= (layer4_outputs(7558)) xor (layer4_outputs(7201));
    outputs(4265) <= not(layer4_outputs(5157));
    outputs(4266) <= layer4_outputs(4921);
    outputs(4267) <= not(layer4_outputs(8649));
    outputs(4268) <= layer4_outputs(223);
    outputs(4269) <= not((layer4_outputs(699)) or (layer4_outputs(3419)));
    outputs(4270) <= not((layer4_outputs(7927)) xor (layer4_outputs(8804)));
    outputs(4271) <= not((layer4_outputs(6170)) xor (layer4_outputs(3143)));
    outputs(4272) <= layer4_outputs(7388);
    outputs(4273) <= layer4_outputs(8942);
    outputs(4274) <= (layer4_outputs(8458)) xor (layer4_outputs(4834));
    outputs(4275) <= layer4_outputs(9205);
    outputs(4276) <= layer4_outputs(9914);
    outputs(4277) <= not(layer4_outputs(9334));
    outputs(4278) <= (layer4_outputs(5484)) and not (layer4_outputs(6958));
    outputs(4279) <= not(layer4_outputs(1199));
    outputs(4280) <= layer4_outputs(2183);
    outputs(4281) <= (layer4_outputs(7880)) and not (layer4_outputs(5287));
    outputs(4282) <= not(layer4_outputs(2283));
    outputs(4283) <= not((layer4_outputs(7233)) xor (layer4_outputs(3486)));
    outputs(4284) <= not(layer4_outputs(5108));
    outputs(4285) <= (layer4_outputs(5805)) xor (layer4_outputs(4861));
    outputs(4286) <= not(layer4_outputs(2042)) or (layer4_outputs(7899));
    outputs(4287) <= not(layer4_outputs(2598));
    outputs(4288) <= layer4_outputs(3622);
    outputs(4289) <= not(layer4_outputs(5069));
    outputs(4290) <= not((layer4_outputs(1198)) or (layer4_outputs(2850)));
    outputs(4291) <= layer4_outputs(2070);
    outputs(4292) <= layer4_outputs(8248);
    outputs(4293) <= (layer4_outputs(3469)) or (layer4_outputs(5324));
    outputs(4294) <= layer4_outputs(6411);
    outputs(4295) <= not(layer4_outputs(1846));
    outputs(4296) <= not(layer4_outputs(2160)) or (layer4_outputs(2669));
    outputs(4297) <= not(layer4_outputs(9296)) or (layer4_outputs(9754));
    outputs(4298) <= layer4_outputs(4059);
    outputs(4299) <= not((layer4_outputs(7059)) xor (layer4_outputs(7407)));
    outputs(4300) <= not((layer4_outputs(6689)) and (layer4_outputs(8396)));
    outputs(4301) <= not(layer4_outputs(8901));
    outputs(4302) <= layer4_outputs(4594);
    outputs(4303) <= layer4_outputs(8907);
    outputs(4304) <= layer4_outputs(9365);
    outputs(4305) <= not((layer4_outputs(3510)) xor (layer4_outputs(8366)));
    outputs(4306) <= layer4_outputs(1673);
    outputs(4307) <= not(layer4_outputs(5482));
    outputs(4308) <= layer4_outputs(7570);
    outputs(4309) <= (layer4_outputs(3141)) and not (layer4_outputs(7920));
    outputs(4310) <= (layer4_outputs(8527)) xor (layer4_outputs(2916));
    outputs(4311) <= not(layer4_outputs(7818));
    outputs(4312) <= layer4_outputs(6944);
    outputs(4313) <= not(layer4_outputs(1772));
    outputs(4314) <= (layer4_outputs(5754)) xor (layer4_outputs(46));
    outputs(4315) <= not(layer4_outputs(7218));
    outputs(4316) <= not(layer4_outputs(8399));
    outputs(4317) <= (layer4_outputs(1464)) and not (layer4_outputs(10014));
    outputs(4318) <= not(layer4_outputs(8266));
    outputs(4319) <= not(layer4_outputs(9673));
    outputs(4320) <= (layer4_outputs(8217)) and not (layer4_outputs(8302));
    outputs(4321) <= not((layer4_outputs(3710)) xor (layer4_outputs(1423)));
    outputs(4322) <= layer4_outputs(8820);
    outputs(4323) <= not((layer4_outputs(712)) xor (layer4_outputs(2273)));
    outputs(4324) <= not(layer4_outputs(2813));
    outputs(4325) <= layer4_outputs(3283);
    outputs(4326) <= layer4_outputs(7825);
    outputs(4327) <= (layer4_outputs(254)) and not (layer4_outputs(2927));
    outputs(4328) <= layer4_outputs(9749);
    outputs(4329) <= (layer4_outputs(3727)) and not (layer4_outputs(7720));
    outputs(4330) <= not(layer4_outputs(4212));
    outputs(4331) <= not((layer4_outputs(5883)) xor (layer4_outputs(4678)));
    outputs(4332) <= layer4_outputs(7404);
    outputs(4333) <= (layer4_outputs(279)) and not (layer4_outputs(2603));
    outputs(4334) <= not(layer4_outputs(7325));
    outputs(4335) <= layer4_outputs(5363);
    outputs(4336) <= not(layer4_outputs(6401));
    outputs(4337) <= not(layer4_outputs(491));
    outputs(4338) <= not(layer4_outputs(3009));
    outputs(4339) <= not(layer4_outputs(8293));
    outputs(4340) <= not(layer4_outputs(6601));
    outputs(4341) <= not((layer4_outputs(9705)) xor (layer4_outputs(697)));
    outputs(4342) <= not(layer4_outputs(3896));
    outputs(4343) <= (layer4_outputs(6389)) and (layer4_outputs(8572));
    outputs(4344) <= not(layer4_outputs(3308));
    outputs(4345) <= (layer4_outputs(4503)) xor (layer4_outputs(4190));
    outputs(4346) <= layer4_outputs(8346);
    outputs(4347) <= not((layer4_outputs(6964)) or (layer4_outputs(1444)));
    outputs(4348) <= layer4_outputs(565);
    outputs(4349) <= layer4_outputs(1320);
    outputs(4350) <= not(layer4_outputs(457));
    outputs(4351) <= layer4_outputs(2596);
    outputs(4352) <= not(layer4_outputs(8153));
    outputs(4353) <= (layer4_outputs(5713)) and not (layer4_outputs(207));
    outputs(4354) <= not(layer4_outputs(3580));
    outputs(4355) <= not((layer4_outputs(3916)) xor (layer4_outputs(10123)));
    outputs(4356) <= (layer4_outputs(2787)) xor (layer4_outputs(8246));
    outputs(4357) <= layer4_outputs(8940);
    outputs(4358) <= not((layer4_outputs(3276)) xor (layer4_outputs(7170)));
    outputs(4359) <= layer4_outputs(4794);
    outputs(4360) <= not(layer4_outputs(2937));
    outputs(4361) <= layer4_outputs(4660);
    outputs(4362) <= not((layer4_outputs(8470)) or (layer4_outputs(8341)));
    outputs(4363) <= not(layer4_outputs(5390));
    outputs(4364) <= (layer4_outputs(10209)) and not (layer4_outputs(6935));
    outputs(4365) <= not((layer4_outputs(9413)) xor (layer4_outputs(3187)));
    outputs(4366) <= not(layer4_outputs(8043));
    outputs(4367) <= layer4_outputs(9010);
    outputs(4368) <= layer4_outputs(9589);
    outputs(4369) <= (layer4_outputs(6319)) and (layer4_outputs(1621));
    outputs(4370) <= not(layer4_outputs(3091));
    outputs(4371) <= not((layer4_outputs(1824)) xor (layer4_outputs(1213)));
    outputs(4372) <= not((layer4_outputs(9730)) or (layer4_outputs(4549)));
    outputs(4373) <= not((layer4_outputs(5776)) and (layer4_outputs(4753)));
    outputs(4374) <= not((layer4_outputs(9485)) xor (layer4_outputs(974)));
    outputs(4375) <= not(layer4_outputs(6416));
    outputs(4376) <= layer4_outputs(7855);
    outputs(4377) <= (layer4_outputs(968)) and not (layer4_outputs(3194));
    outputs(4378) <= not(layer4_outputs(2528)) or (layer4_outputs(1892));
    outputs(4379) <= not(layer4_outputs(9412));
    outputs(4380) <= not(layer4_outputs(4740));
    outputs(4381) <= (layer4_outputs(3971)) xor (layer4_outputs(1736));
    outputs(4382) <= layer4_outputs(1356);
    outputs(4383) <= layer4_outputs(4666);
    outputs(4384) <= layer4_outputs(6849);
    outputs(4385) <= not(layer4_outputs(1221));
    outputs(4386) <= not(layer4_outputs(308));
    outputs(4387) <= not((layer4_outputs(1275)) xor (layer4_outputs(2026)));
    outputs(4388) <= not((layer4_outputs(6359)) or (layer4_outputs(2534)));
    outputs(4389) <= not((layer4_outputs(7007)) xor (layer4_outputs(795)));
    outputs(4390) <= (layer4_outputs(1830)) or (layer4_outputs(2353));
    outputs(4391) <= layer4_outputs(2181);
    outputs(4392) <= (layer4_outputs(7994)) xor (layer4_outputs(1098));
    outputs(4393) <= layer4_outputs(9752);
    outputs(4394) <= (layer4_outputs(1987)) and (layer4_outputs(3413));
    outputs(4395) <= layer4_outputs(7010);
    outputs(4396) <= not(layer4_outputs(8070));
    outputs(4397) <= not(layer4_outputs(6529));
    outputs(4398) <= layer4_outputs(406);
    outputs(4399) <= (layer4_outputs(6701)) and not (layer4_outputs(3955));
    outputs(4400) <= not((layer4_outputs(2434)) xor (layer4_outputs(9488)));
    outputs(4401) <= (layer4_outputs(2603)) xor (layer4_outputs(9653));
    outputs(4402) <= not((layer4_outputs(3220)) xor (layer4_outputs(3165)));
    outputs(4403) <= not((layer4_outputs(2132)) xor (layer4_outputs(250)));
    outputs(4404) <= layer4_outputs(1104);
    outputs(4405) <= '1';
    outputs(4406) <= not(layer4_outputs(6246));
    outputs(4407) <= layer4_outputs(8951);
    outputs(4408) <= '0';
    outputs(4409) <= not((layer4_outputs(2461)) xor (layer4_outputs(7865)));
    outputs(4410) <= not(layer4_outputs(4541));
    outputs(4411) <= (layer4_outputs(8570)) and (layer4_outputs(8187));
    outputs(4412) <= layer4_outputs(3696);
    outputs(4413) <= layer4_outputs(434);
    outputs(4414) <= not((layer4_outputs(5742)) or (layer4_outputs(2270)));
    outputs(4415) <= layer4_outputs(249);
    outputs(4416) <= not((layer4_outputs(7239)) xor (layer4_outputs(8768)));
    outputs(4417) <= not(layer4_outputs(7154));
    outputs(4418) <= (layer4_outputs(9222)) and not (layer4_outputs(5877));
    outputs(4419) <= not(layer4_outputs(3818));
    outputs(4420) <= layer4_outputs(427);
    outputs(4421) <= not(layer4_outputs(569));
    outputs(4422) <= not(layer4_outputs(2341));
    outputs(4423) <= layer4_outputs(9357);
    outputs(4424) <= not(layer4_outputs(1394)) or (layer4_outputs(240));
    outputs(4425) <= not(layer4_outputs(1902));
    outputs(4426) <= not(layer4_outputs(5534)) or (layer4_outputs(2945));
    outputs(4427) <= not((layer4_outputs(1358)) or (layer4_outputs(9361)));
    outputs(4428) <= (layer4_outputs(9638)) and not (layer4_outputs(8423));
    outputs(4429) <= not(layer4_outputs(9342));
    outputs(4430) <= not(layer4_outputs(1538));
    outputs(4431) <= layer4_outputs(9923);
    outputs(4432) <= (layer4_outputs(4530)) and (layer4_outputs(3526));
    outputs(4433) <= not(layer4_outputs(4980));
    outputs(4434) <= not(layer4_outputs(7974));
    outputs(4435) <= not(layer4_outputs(2312)) or (layer4_outputs(2635));
    outputs(4436) <= not(layer4_outputs(4765));
    outputs(4437) <= not(layer4_outputs(9951));
    outputs(4438) <= not((layer4_outputs(3245)) xor (layer4_outputs(8423)));
    outputs(4439) <= not(layer4_outputs(1556));
    outputs(4440) <= not((layer4_outputs(9142)) xor (layer4_outputs(841)));
    outputs(4441) <= layer4_outputs(331);
    outputs(4442) <= not(layer4_outputs(5140));
    outputs(4443) <= layer4_outputs(7241);
    outputs(4444) <= (layer4_outputs(1964)) xor (layer4_outputs(5506));
    outputs(4445) <= layer4_outputs(5262);
    outputs(4446) <= not(layer4_outputs(5830));
    outputs(4447) <= not((layer4_outputs(3737)) or (layer4_outputs(1602)));
    outputs(4448) <= (layer4_outputs(7448)) xor (layer4_outputs(1243));
    outputs(4449) <= layer4_outputs(4948);
    outputs(4450) <= not(layer4_outputs(1640));
    outputs(4451) <= not((layer4_outputs(7599)) or (layer4_outputs(2623)));
    outputs(4452) <= layer4_outputs(4041);
    outputs(4453) <= not((layer4_outputs(4569)) xor (layer4_outputs(2602)));
    outputs(4454) <= layer4_outputs(749);
    outputs(4455) <= not(layer4_outputs(9288));
    outputs(4456) <= not(layer4_outputs(8487));
    outputs(4457) <= not((layer4_outputs(2248)) xor (layer4_outputs(6786)));
    outputs(4458) <= (layer4_outputs(1713)) xor (layer4_outputs(9897));
    outputs(4459) <= (layer4_outputs(9217)) and (layer4_outputs(4231));
    outputs(4460) <= not(layer4_outputs(10219));
    outputs(4461) <= (layer4_outputs(4347)) xor (layer4_outputs(571));
    outputs(4462) <= not((layer4_outputs(2334)) xor (layer4_outputs(4061)));
    outputs(4463) <= (layer4_outputs(8267)) and not (layer4_outputs(8800));
    outputs(4464) <= layer4_outputs(1567);
    outputs(4465) <= (layer4_outputs(9874)) and not (layer4_outputs(113));
    outputs(4466) <= layer4_outputs(544);
    outputs(4467) <= not((layer4_outputs(1547)) xor (layer4_outputs(9913)));
    outputs(4468) <= not((layer4_outputs(441)) and (layer4_outputs(2440)));
    outputs(4469) <= not((layer4_outputs(1289)) xor (layer4_outputs(6532)));
    outputs(4470) <= layer4_outputs(1339);
    outputs(4471) <= layer4_outputs(1786);
    outputs(4472) <= layer4_outputs(8775);
    outputs(4473) <= not(layer4_outputs(6536));
    outputs(4474) <= not(layer4_outputs(8646));
    outputs(4475) <= not((layer4_outputs(336)) and (layer4_outputs(7201)));
    outputs(4476) <= layer4_outputs(3093);
    outputs(4477) <= layer4_outputs(3801);
    outputs(4478) <= layer4_outputs(8718);
    outputs(4479) <= (layer4_outputs(4104)) xor (layer4_outputs(7049));
    outputs(4480) <= layer4_outputs(3655);
    outputs(4481) <= (layer4_outputs(3539)) xor (layer4_outputs(3798));
    outputs(4482) <= not((layer4_outputs(3524)) or (layer4_outputs(2275)));
    outputs(4483) <= '0';
    outputs(4484) <= '0';
    outputs(4485) <= layer4_outputs(6624);
    outputs(4486) <= layer4_outputs(5740);
    outputs(4487) <= (layer4_outputs(116)) and not (layer4_outputs(9560));
    outputs(4488) <= not(layer4_outputs(3201));
    outputs(4489) <= not(layer4_outputs(7893));
    outputs(4490) <= not(layer4_outputs(979));
    outputs(4491) <= not(layer4_outputs(6095));
    outputs(4492) <= not(layer4_outputs(2495));
    outputs(4493) <= (layer4_outputs(3532)) and not (layer4_outputs(10087));
    outputs(4494) <= layer4_outputs(10102);
    outputs(4495) <= not(layer4_outputs(320));
    outputs(4496) <= not(layer4_outputs(8373));
    outputs(4497) <= (layer4_outputs(6873)) xor (layer4_outputs(669));
    outputs(4498) <= not(layer4_outputs(7169));
    outputs(4499) <= layer4_outputs(6297);
    outputs(4500) <= not(layer4_outputs(3839)) or (layer4_outputs(3191));
    outputs(4501) <= (layer4_outputs(8335)) and not (layer4_outputs(5447));
    outputs(4502) <= not(layer4_outputs(6492));
    outputs(4503) <= layer4_outputs(3306);
    outputs(4504) <= (layer4_outputs(8290)) xor (layer4_outputs(8198));
    outputs(4505) <= not((layer4_outputs(5253)) and (layer4_outputs(8410)));
    outputs(4506) <= not(layer4_outputs(7068));
    outputs(4507) <= not(layer4_outputs(6104));
    outputs(4508) <= layer4_outputs(2021);
    outputs(4509) <= not((layer4_outputs(9988)) xor (layer4_outputs(7269)));
    outputs(4510) <= not(layer4_outputs(8935));
    outputs(4511) <= not((layer4_outputs(7836)) xor (layer4_outputs(4901)));
    outputs(4512) <= layer4_outputs(2436);
    outputs(4513) <= not((layer4_outputs(6436)) and (layer4_outputs(533)));
    outputs(4514) <= not(layer4_outputs(3630));
    outputs(4515) <= not(layer4_outputs(2932));
    outputs(4516) <= not(layer4_outputs(3196));
    outputs(4517) <= not(layer4_outputs(5552));
    outputs(4518) <= (layer4_outputs(6594)) xor (layer4_outputs(1155));
    outputs(4519) <= layer4_outputs(6555);
    outputs(4520) <= not(layer4_outputs(1132));
    outputs(4521) <= (layer4_outputs(9402)) xor (layer4_outputs(9735));
    outputs(4522) <= (layer4_outputs(6217)) and (layer4_outputs(4556));
    outputs(4523) <= layer4_outputs(6327);
    outputs(4524) <= (layer4_outputs(1833)) and (layer4_outputs(6414));
    outputs(4525) <= not((layer4_outputs(606)) xor (layer4_outputs(8827)));
    outputs(4526) <= layer4_outputs(3913);
    outputs(4527) <= not((layer4_outputs(5097)) xor (layer4_outputs(2305)));
    outputs(4528) <= layer4_outputs(2198);
    outputs(4529) <= not((layer4_outputs(2457)) or (layer4_outputs(1253)));
    outputs(4530) <= layer4_outputs(6098);
    outputs(4531) <= layer4_outputs(5122);
    outputs(4532) <= layer4_outputs(1792);
    outputs(4533) <= not((layer4_outputs(4943)) xor (layer4_outputs(6298)));
    outputs(4534) <= layer4_outputs(4183);
    outputs(4535) <= not((layer4_outputs(1527)) or (layer4_outputs(7650)));
    outputs(4536) <= layer4_outputs(5646);
    outputs(4537) <= layer4_outputs(3389);
    outputs(4538) <= not(layer4_outputs(2016));
    outputs(4539) <= not(layer4_outputs(3154));
    outputs(4540) <= (layer4_outputs(1929)) and (layer4_outputs(8538));
    outputs(4541) <= not(layer4_outputs(8302));
    outputs(4542) <= not((layer4_outputs(7715)) xor (layer4_outputs(7395)));
    outputs(4543) <= layer4_outputs(898);
    outputs(4544) <= layer4_outputs(6761);
    outputs(4545) <= not(layer4_outputs(9035));
    outputs(4546) <= (layer4_outputs(9235)) and not (layer4_outputs(2956));
    outputs(4547) <= (layer4_outputs(3970)) and not (layer4_outputs(3388));
    outputs(4548) <= layer4_outputs(6703);
    outputs(4549) <= layer4_outputs(181);
    outputs(4550) <= layer4_outputs(1545);
    outputs(4551) <= (layer4_outputs(9965)) and not (layer4_outputs(524));
    outputs(4552) <= not(layer4_outputs(5070)) or (layer4_outputs(2161));
    outputs(4553) <= not((layer4_outputs(5395)) or (layer4_outputs(6333)));
    outputs(4554) <= not((layer4_outputs(4301)) or (layer4_outputs(9311)));
    outputs(4555) <= not(layer4_outputs(5558));
    outputs(4556) <= not(layer4_outputs(5063)) or (layer4_outputs(5290));
    outputs(4557) <= layer4_outputs(889);
    outputs(4558) <= not(layer4_outputs(6693));
    outputs(4559) <= not(layer4_outputs(5160));
    outputs(4560) <= not(layer4_outputs(9741));
    outputs(4561) <= not((layer4_outputs(3873)) and (layer4_outputs(5392)));
    outputs(4562) <= not(layer4_outputs(5634));
    outputs(4563) <= layer4_outputs(7595);
    outputs(4564) <= (layer4_outputs(566)) xor (layer4_outputs(8184));
    outputs(4565) <= (layer4_outputs(5455)) xor (layer4_outputs(6376));
    outputs(4566) <= not(layer4_outputs(5274));
    outputs(4567) <= (layer4_outputs(3667)) or (layer4_outputs(1974));
    outputs(4568) <= layer4_outputs(5518);
    outputs(4569) <= (layer4_outputs(3840)) xor (layer4_outputs(9797));
    outputs(4570) <= not(layer4_outputs(6695));
    outputs(4571) <= not((layer4_outputs(6931)) and (layer4_outputs(1659)));
    outputs(4572) <= not(layer4_outputs(3709));
    outputs(4573) <= layer4_outputs(4315);
    outputs(4574) <= not((layer4_outputs(9643)) or (layer4_outputs(6817)));
    outputs(4575) <= not(layer4_outputs(401));
    outputs(4576) <= layer4_outputs(6810);
    outputs(4577) <= not(layer4_outputs(5985));
    outputs(4578) <= not((layer4_outputs(2028)) xor (layer4_outputs(1326)));
    outputs(4579) <= layer4_outputs(5843);
    outputs(4580) <= (layer4_outputs(476)) xor (layer4_outputs(1089));
    outputs(4581) <= not(layer4_outputs(7166));
    outputs(4582) <= (layer4_outputs(6912)) xor (layer4_outputs(8941));
    outputs(4583) <= layer4_outputs(246);
    outputs(4584) <= not((layer4_outputs(9936)) or (layer4_outputs(4700)));
    outputs(4585) <= layer4_outputs(1020);
    outputs(4586) <= (layer4_outputs(8363)) xor (layer4_outputs(140));
    outputs(4587) <= not((layer4_outputs(1235)) or (layer4_outputs(6994)));
    outputs(4588) <= not(layer4_outputs(4810));
    outputs(4589) <= not(layer4_outputs(431));
    outputs(4590) <= (layer4_outputs(5348)) xor (layer4_outputs(3783));
    outputs(4591) <= layer4_outputs(1398);
    outputs(4592) <= not(layer4_outputs(5209));
    outputs(4593) <= layer4_outputs(8139);
    outputs(4594) <= layer4_outputs(3865);
    outputs(4595) <= (layer4_outputs(3536)) xor (layer4_outputs(1909));
    outputs(4596) <= not((layer4_outputs(996)) xor (layer4_outputs(6149)));
    outputs(4597) <= not(layer4_outputs(6214));
    outputs(4598) <= not(layer4_outputs(4487));
    outputs(4599) <= not((layer4_outputs(1702)) or (layer4_outputs(6330)));
    outputs(4600) <= (layer4_outputs(8950)) and (layer4_outputs(9638));
    outputs(4601) <= (layer4_outputs(551)) and not (layer4_outputs(554));
    outputs(4602) <= not(layer4_outputs(7203));
    outputs(4603) <= (layer4_outputs(5580)) and (layer4_outputs(6063));
    outputs(4604) <= (layer4_outputs(7324)) xor (layer4_outputs(3323));
    outputs(4605) <= not((layer4_outputs(3112)) xor (layer4_outputs(583)));
    outputs(4606) <= not((layer4_outputs(6726)) xor (layer4_outputs(3548)));
    outputs(4607) <= not(layer4_outputs(4300));
    outputs(4608) <= (layer4_outputs(4236)) xor (layer4_outputs(4581));
    outputs(4609) <= not(layer4_outputs(530));
    outputs(4610) <= layer4_outputs(9546);
    outputs(4611) <= not((layer4_outputs(7255)) xor (layer4_outputs(7972)));
    outputs(4612) <= layer4_outputs(2452);
    outputs(4613) <= (layer4_outputs(5291)) xor (layer4_outputs(9542));
    outputs(4614) <= not(layer4_outputs(5532));
    outputs(4615) <= not(layer4_outputs(5705));
    outputs(4616) <= layer4_outputs(3869);
    outputs(4617) <= not(layer4_outputs(3578));
    outputs(4618) <= not(layer4_outputs(3533));
    outputs(4619) <= (layer4_outputs(5621)) xor (layer4_outputs(3901));
    outputs(4620) <= (layer4_outputs(9754)) or (layer4_outputs(980));
    outputs(4621) <= not(layer4_outputs(10122));
    outputs(4622) <= not(layer4_outputs(754));
    outputs(4623) <= layer4_outputs(5523);
    outputs(4624) <= layer4_outputs(5216);
    outputs(4625) <= layer4_outputs(9512);
    outputs(4626) <= not((layer4_outputs(4304)) xor (layer4_outputs(2688)));
    outputs(4627) <= layer4_outputs(7840);
    outputs(4628) <= not((layer4_outputs(8548)) xor (layer4_outputs(8236)));
    outputs(4629) <= not(layer4_outputs(5576));
    outputs(4630) <= layer4_outputs(9280);
    outputs(4631) <= (layer4_outputs(6309)) xor (layer4_outputs(6859));
    outputs(4632) <= not((layer4_outputs(8499)) or (layer4_outputs(2708)));
    outputs(4633) <= layer4_outputs(2875);
    outputs(4634) <= (layer4_outputs(1488)) xor (layer4_outputs(4941));
    outputs(4635) <= (layer4_outputs(1187)) xor (layer4_outputs(9537));
    outputs(4636) <= not(layer4_outputs(8179)) or (layer4_outputs(1171));
    outputs(4637) <= layer4_outputs(7128);
    outputs(4638) <= layer4_outputs(7328);
    outputs(4639) <= not(layer4_outputs(6302)) or (layer4_outputs(7546));
    outputs(4640) <= layer4_outputs(5617);
    outputs(4641) <= (layer4_outputs(5480)) and not (layer4_outputs(5122));
    outputs(4642) <= not(layer4_outputs(209));
    outputs(4643) <= (layer4_outputs(6069)) and (layer4_outputs(1596));
    outputs(4644) <= (layer4_outputs(8329)) xor (layer4_outputs(6482));
    outputs(4645) <= not(layer4_outputs(8388));
    outputs(4646) <= not(layer4_outputs(8973));
    outputs(4647) <= not(layer4_outputs(3490));
    outputs(4648) <= (layer4_outputs(1468)) xor (layer4_outputs(1343));
    outputs(4649) <= not(layer4_outputs(5519));
    outputs(4650) <= layer4_outputs(5792);
    outputs(4651) <= not(layer4_outputs(3289));
    outputs(4652) <= not(layer4_outputs(7867));
    outputs(4653) <= layer4_outputs(4480);
    outputs(4654) <= not(layer4_outputs(5144));
    outputs(4655) <= layer4_outputs(2836);
    outputs(4656) <= (layer4_outputs(10059)) xor (layer4_outputs(3787));
    outputs(4657) <= not(layer4_outputs(1164));
    outputs(4658) <= not(layer4_outputs(3757));
    outputs(4659) <= not(layer4_outputs(4364));
    outputs(4660) <= (layer4_outputs(7263)) and (layer4_outputs(1784));
    outputs(4661) <= layer4_outputs(9510);
    outputs(4662) <= layer4_outputs(8033);
    outputs(4663) <= layer4_outputs(1794);
    outputs(4664) <= not(layer4_outputs(5794));
    outputs(4665) <= layer4_outputs(9261);
    outputs(4666) <= not(layer4_outputs(4683));
    outputs(4667) <= (layer4_outputs(8990)) and not (layer4_outputs(798));
    outputs(4668) <= (layer4_outputs(7274)) xor (layer4_outputs(4496));
    outputs(4669) <= (layer4_outputs(1111)) xor (layer4_outputs(25));
    outputs(4670) <= (layer4_outputs(9367)) xor (layer4_outputs(1453));
    outputs(4671) <= not(layer4_outputs(5056));
    outputs(4672) <= layer4_outputs(1615);
    outputs(4673) <= (layer4_outputs(1901)) and not (layer4_outputs(9755));
    outputs(4674) <= layer4_outputs(4191);
    outputs(4675) <= not(layer4_outputs(1120));
    outputs(4676) <= layer4_outputs(4988);
    outputs(4677) <= (layer4_outputs(7192)) or (layer4_outputs(6569));
    outputs(4678) <= layer4_outputs(1065);
    outputs(4679) <= layer4_outputs(9789);
    outputs(4680) <= layer4_outputs(2289);
    outputs(4681) <= not((layer4_outputs(528)) xor (layer4_outputs(7910)));
    outputs(4682) <= (layer4_outputs(6479)) xor (layer4_outputs(9860));
    outputs(4683) <= (layer4_outputs(1187)) xor (layer4_outputs(507));
    outputs(4684) <= layer4_outputs(1359);
    outputs(4685) <= layer4_outputs(3389);
    outputs(4686) <= layer4_outputs(2056);
    outputs(4687) <= (layer4_outputs(2200)) and (layer4_outputs(10204));
    outputs(4688) <= not((layer4_outputs(9962)) xor (layer4_outputs(9273)));
    outputs(4689) <= layer4_outputs(1621);
    outputs(4690) <= (layer4_outputs(5969)) xor (layer4_outputs(3760));
    outputs(4691) <= not((layer4_outputs(2317)) and (layer4_outputs(2250)));
    outputs(4692) <= not((layer4_outputs(7425)) xor (layer4_outputs(5434)));
    outputs(4693) <= not(layer4_outputs(7860));
    outputs(4694) <= (layer4_outputs(8728)) and not (layer4_outputs(3471));
    outputs(4695) <= layer4_outputs(3835);
    outputs(4696) <= layer4_outputs(7915);
    outputs(4697) <= not(layer4_outputs(5507));
    outputs(4698) <= not(layer4_outputs(236));
    outputs(4699) <= (layer4_outputs(8815)) xor (layer4_outputs(3593));
    outputs(4700) <= not((layer4_outputs(9770)) xor (layer4_outputs(8171)));
    outputs(4701) <= not(layer4_outputs(4979));
    outputs(4702) <= not(layer4_outputs(8161));
    outputs(4703) <= (layer4_outputs(641)) xor (layer4_outputs(3337));
    outputs(4704) <= layer4_outputs(3380);
    outputs(4705) <= not((layer4_outputs(7772)) or (layer4_outputs(5426)));
    outputs(4706) <= not((layer4_outputs(6662)) xor (layer4_outputs(10044)));
    outputs(4707) <= layer4_outputs(2539);
    outputs(4708) <= not(layer4_outputs(9336));
    outputs(4709) <= layer4_outputs(2833);
    outputs(4710) <= layer4_outputs(7932);
    outputs(4711) <= layer4_outputs(700);
    outputs(4712) <= (layer4_outputs(9497)) and not (layer4_outputs(7625));
    outputs(4713) <= layer4_outputs(3152);
    outputs(4714) <= not(layer4_outputs(7077));
    outputs(4715) <= (layer4_outputs(1079)) and not (layer4_outputs(2400));
    outputs(4716) <= not(layer4_outputs(9034));
    outputs(4717) <= not(layer4_outputs(3766));
    outputs(4718) <= (layer4_outputs(5485)) and (layer4_outputs(628));
    outputs(4719) <= layer4_outputs(722);
    outputs(4720) <= not((layer4_outputs(7042)) xor (layer4_outputs(6034)));
    outputs(4721) <= not(layer4_outputs(9091));
    outputs(4722) <= not((layer4_outputs(6053)) xor (layer4_outputs(9414)));
    outputs(4723) <= layer4_outputs(9850);
    outputs(4724) <= not((layer4_outputs(6608)) and (layer4_outputs(2141)));
    outputs(4725) <= not(layer4_outputs(7722));
    outputs(4726) <= not((layer4_outputs(7668)) and (layer4_outputs(6102)));
    outputs(4727) <= not(layer4_outputs(666));
    outputs(4728) <= layer4_outputs(2745);
    outputs(4729) <= not((layer4_outputs(8126)) xor (layer4_outputs(5515)));
    outputs(4730) <= not(layer4_outputs(6628));
    outputs(4731) <= (layer4_outputs(8217)) xor (layer4_outputs(8233));
    outputs(4732) <= layer4_outputs(2981);
    outputs(4733) <= not((layer4_outputs(4568)) xor (layer4_outputs(7871)));
    outputs(4734) <= layer4_outputs(3089);
    outputs(4735) <= not(layer4_outputs(4392));
    outputs(4736) <= (layer4_outputs(10107)) xor (layer4_outputs(8872));
    outputs(4737) <= (layer4_outputs(1878)) or (layer4_outputs(2794));
    outputs(4738) <= not(layer4_outputs(4060));
    outputs(4739) <= (layer4_outputs(8947)) and not (layer4_outputs(7369));
    outputs(4740) <= layer4_outputs(8570);
    outputs(4741) <= (layer4_outputs(2158)) xor (layer4_outputs(6127));
    outputs(4742) <= not(layer4_outputs(7326));
    outputs(4743) <= not(layer4_outputs(5616));
    outputs(4744) <= not(layer4_outputs(4776));
    outputs(4745) <= not(layer4_outputs(8298));
    outputs(4746) <= layer4_outputs(5403);
    outputs(4747) <= layer4_outputs(5965);
    outputs(4748) <= not(layer4_outputs(2607));
    outputs(4749) <= not(layer4_outputs(873));
    outputs(4750) <= layer4_outputs(8777);
    outputs(4751) <= layer4_outputs(9292);
    outputs(4752) <= not(layer4_outputs(6478));
    outputs(4753) <= not(layer4_outputs(194));
    outputs(4754) <= not(layer4_outputs(1912)) or (layer4_outputs(265));
    outputs(4755) <= not((layer4_outputs(5275)) xor (layer4_outputs(6791)));
    outputs(4756) <= not((layer4_outputs(4549)) and (layer4_outputs(7092)));
    outputs(4757) <= not(layer4_outputs(8614));
    outputs(4758) <= layer4_outputs(5486);
    outputs(4759) <= (layer4_outputs(1871)) and (layer4_outputs(4857));
    outputs(4760) <= not(layer4_outputs(3605));
    outputs(4761) <= layer4_outputs(9488);
    outputs(4762) <= (layer4_outputs(6325)) and (layer4_outputs(8571));
    outputs(4763) <= (layer4_outputs(2763)) xor (layer4_outputs(3227));
    outputs(4764) <= layer4_outputs(4948);
    outputs(4765) <= layer4_outputs(9423);
    outputs(4766) <= layer4_outputs(1313);
    outputs(4767) <= not(layer4_outputs(2814));
    outputs(4768) <= not(layer4_outputs(4866));
    outputs(4769) <= layer4_outputs(3317);
    outputs(4770) <= not((layer4_outputs(8900)) or (layer4_outputs(8525)));
    outputs(4771) <= layer4_outputs(4502);
    outputs(4772) <= layer4_outputs(1802);
    outputs(4773) <= not((layer4_outputs(5351)) xor (layer4_outputs(4124)));
    outputs(4774) <= not((layer4_outputs(3581)) xor (layer4_outputs(2150)));
    outputs(4775) <= not(layer4_outputs(2080));
    outputs(4776) <= layer4_outputs(5769);
    outputs(4777) <= not(layer4_outputs(4802));
    outputs(4778) <= layer4_outputs(9470);
    outputs(4779) <= (layer4_outputs(2940)) xor (layer4_outputs(1957));
    outputs(4780) <= layer4_outputs(1887);
    outputs(4781) <= not(layer4_outputs(465));
    outputs(4782) <= not((layer4_outputs(6310)) xor (layer4_outputs(6201)));
    outputs(4783) <= (layer4_outputs(5190)) xor (layer4_outputs(1820));
    outputs(4784) <= layer4_outputs(760);
    outputs(4785) <= layer4_outputs(1455);
    outputs(4786) <= not(layer4_outputs(441));
    outputs(4787) <= not(layer4_outputs(593));
    outputs(4788) <= not(layer4_outputs(4116));
    outputs(4789) <= not(layer4_outputs(9076));
    outputs(4790) <= (layer4_outputs(2321)) and not (layer4_outputs(6254));
    outputs(4791) <= layer4_outputs(8727);
    outputs(4792) <= (layer4_outputs(4916)) xor (layer4_outputs(4649));
    outputs(4793) <= not(layer4_outputs(7903));
    outputs(4794) <= (layer4_outputs(2237)) and not (layer4_outputs(8785));
    outputs(4795) <= layer4_outputs(10199);
    outputs(4796) <= (layer4_outputs(6747)) and not (layer4_outputs(6377));
    outputs(4797) <= layer4_outputs(3168);
    outputs(4798) <= not((layer4_outputs(5919)) or (layer4_outputs(2622)));
    outputs(4799) <= layer4_outputs(7291);
    outputs(4800) <= layer4_outputs(672);
    outputs(4801) <= layer4_outputs(9649);
    outputs(4802) <= not(layer4_outputs(2063));
    outputs(4803) <= not(layer4_outputs(2641)) or (layer4_outputs(7885));
    outputs(4804) <= layer4_outputs(1758);
    outputs(4805) <= (layer4_outputs(2822)) xor (layer4_outputs(6109));
    outputs(4806) <= not(layer4_outputs(2640));
    outputs(4807) <= (layer4_outputs(8506)) xor (layer4_outputs(378));
    outputs(4808) <= (layer4_outputs(6175)) and not (layer4_outputs(6499));
    outputs(4809) <= not(layer4_outputs(3422)) or (layer4_outputs(1739));
    outputs(4810) <= not((layer4_outputs(8303)) or (layer4_outputs(869)));
    outputs(4811) <= layer4_outputs(9639);
    outputs(4812) <= not(layer4_outputs(7134));
    outputs(4813) <= not(layer4_outputs(6980));
    outputs(4814) <= (layer4_outputs(3240)) xor (layer4_outputs(1615));
    outputs(4815) <= not(layer4_outputs(2020));
    outputs(4816) <= (layer4_outputs(6549)) and (layer4_outputs(678));
    outputs(4817) <= layer4_outputs(10114);
    outputs(4818) <= not(layer4_outputs(5590));
    outputs(4819) <= not(layer4_outputs(2790));
    outputs(4820) <= (layer4_outputs(2448)) and (layer4_outputs(10050));
    outputs(4821) <= not(layer4_outputs(99));
    outputs(4822) <= layer4_outputs(5492);
    outputs(4823) <= layer4_outputs(8354);
    outputs(4824) <= (layer4_outputs(3794)) and not (layer4_outputs(6020));
    outputs(4825) <= not(layer4_outputs(7066));
    outputs(4826) <= not(layer4_outputs(5541));
    outputs(4827) <= not((layer4_outputs(5798)) xor (layer4_outputs(9908)));
    outputs(4828) <= not(layer4_outputs(3508));
    outputs(4829) <= not(layer4_outputs(8062));
    outputs(4830) <= not((layer4_outputs(3621)) xor (layer4_outputs(3932)));
    outputs(4831) <= layer4_outputs(1553);
    outputs(4832) <= not(layer4_outputs(7929));
    outputs(4833) <= layer4_outputs(7793);
    outputs(4834) <= (layer4_outputs(7131)) xor (layer4_outputs(4202));
    outputs(4835) <= layer4_outputs(3804);
    outputs(4836) <= layer4_outputs(3946);
    outputs(4837) <= layer4_outputs(7141);
    outputs(4838) <= (layer4_outputs(2408)) and (layer4_outputs(9328));
    outputs(4839) <= (layer4_outputs(9773)) and (layer4_outputs(9521));
    outputs(4840) <= (layer4_outputs(9665)) and not (layer4_outputs(9094));
    outputs(4841) <= (layer4_outputs(6037)) and not (layer4_outputs(1971));
    outputs(4842) <= (layer4_outputs(1343)) and not (layer4_outputs(10011));
    outputs(4843) <= (layer4_outputs(6965)) xor (layer4_outputs(4134));
    outputs(4844) <= not(layer4_outputs(6018));
    outputs(4845) <= (layer4_outputs(3914)) and not (layer4_outputs(2065));
    outputs(4846) <= layer4_outputs(3598);
    outputs(4847) <= not((layer4_outputs(9080)) xor (layer4_outputs(321)));
    outputs(4848) <= (layer4_outputs(9482)) or (layer4_outputs(7389));
    outputs(4849) <= not((layer4_outputs(9832)) xor (layer4_outputs(2354)));
    outputs(4850) <= not((layer4_outputs(7076)) or (layer4_outputs(4897)));
    outputs(4851) <= not(layer4_outputs(4916));
    outputs(4852) <= (layer4_outputs(5305)) and not (layer4_outputs(933));
    outputs(4853) <= layer4_outputs(9827);
    outputs(4854) <= (layer4_outputs(7643)) xor (layer4_outputs(8736));
    outputs(4855) <= not(layer4_outputs(7930)) or (layer4_outputs(6383));
    outputs(4856) <= layer4_outputs(9126);
    outputs(4857) <= (layer4_outputs(7912)) and not (layer4_outputs(356));
    outputs(4858) <= (layer4_outputs(4150)) and not (layer4_outputs(3551));
    outputs(4859) <= not(layer4_outputs(29));
    outputs(4860) <= layer4_outputs(1346);
    outputs(4861) <= not((layer4_outputs(7075)) or (layer4_outputs(5592)));
    outputs(4862) <= not(layer4_outputs(8067));
    outputs(4863) <= not((layer4_outputs(8162)) and (layer4_outputs(383)));
    outputs(4864) <= (layer4_outputs(7519)) xor (layer4_outputs(10111));
    outputs(4865) <= not((layer4_outputs(8086)) xor (layer4_outputs(8107)));
    outputs(4866) <= not((layer4_outputs(4891)) or (layer4_outputs(9803)));
    outputs(4867) <= not(layer4_outputs(6943));
    outputs(4868) <= not(layer4_outputs(7167));
    outputs(4869) <= not(layer4_outputs(7761));
    outputs(4870) <= (layer4_outputs(6367)) xor (layer4_outputs(3893));
    outputs(4871) <= not(layer4_outputs(3282));
    outputs(4872) <= not(layer4_outputs(2563));
    outputs(4873) <= layer4_outputs(7706);
    outputs(4874) <= not(layer4_outputs(2614));
    outputs(4875) <= not((layer4_outputs(9289)) or (layer4_outputs(7031)));
    outputs(4876) <= (layer4_outputs(6426)) and not (layer4_outputs(8054));
    outputs(4877) <= layer4_outputs(3092);
    outputs(4878) <= not(layer4_outputs(9791));
    outputs(4879) <= not(layer4_outputs(2711));
    outputs(4880) <= not(layer4_outputs(4774));
    outputs(4881) <= not((layer4_outputs(2014)) xor (layer4_outputs(7403)));
    outputs(4882) <= layer4_outputs(3936);
    outputs(4883) <= (layer4_outputs(4528)) and not (layer4_outputs(3721));
    outputs(4884) <= not(layer4_outputs(2725));
    outputs(4885) <= layer4_outputs(6667);
    outputs(4886) <= layer4_outputs(4998);
    outputs(4887) <= layer4_outputs(1049);
    outputs(4888) <= not((layer4_outputs(9247)) xor (layer4_outputs(7051)));
    outputs(4889) <= layer4_outputs(3101);
    outputs(4890) <= (layer4_outputs(5113)) and not (layer4_outputs(8058));
    outputs(4891) <= not(layer4_outputs(2605));
    outputs(4892) <= not(layer4_outputs(3005));
    outputs(4893) <= not(layer4_outputs(2588));
    outputs(4894) <= not(layer4_outputs(4979));
    outputs(4895) <= (layer4_outputs(8203)) or (layer4_outputs(9838));
    outputs(4896) <= not(layer4_outputs(5859));
    outputs(4897) <= not(layer4_outputs(7834));
    outputs(4898) <= not(layer4_outputs(3167));
    outputs(4899) <= (layer4_outputs(2578)) and (layer4_outputs(4219));
    outputs(4900) <= not(layer4_outputs(2519));
    outputs(4901) <= (layer4_outputs(6660)) xor (layer4_outputs(219));
    outputs(4902) <= not((layer4_outputs(2513)) xor (layer4_outputs(776)));
    outputs(4903) <= (layer4_outputs(1438)) and not (layer4_outputs(4773));
    outputs(4904) <= not(layer4_outputs(9436));
    outputs(4905) <= layer4_outputs(7963);
    outputs(4906) <= (layer4_outputs(302)) xor (layer4_outputs(6698));
    outputs(4907) <= not((layer4_outputs(3070)) xor (layer4_outputs(7794)));
    outputs(4908) <= (layer4_outputs(1793)) and (layer4_outputs(7387));
    outputs(4909) <= not((layer4_outputs(4098)) and (layer4_outputs(7594)));
    outputs(4910) <= layer4_outputs(721);
    outputs(4911) <= not((layer4_outputs(2243)) and (layer4_outputs(4892)));
    outputs(4912) <= not(layer4_outputs(10039));
    outputs(4913) <= not(layer4_outputs(8341));
    outputs(4914) <= not(layer4_outputs(705));
    outputs(4915) <= not(layer4_outputs(4662));
    outputs(4916) <= layer4_outputs(2835);
    outputs(4917) <= not((layer4_outputs(8411)) xor (layer4_outputs(7906)));
    outputs(4918) <= not(layer4_outputs(7769));
    outputs(4919) <= layer4_outputs(3903);
    outputs(4920) <= (layer4_outputs(2835)) and not (layer4_outputs(4748));
    outputs(4921) <= not(layer4_outputs(9596)) or (layer4_outputs(8837));
    outputs(4922) <= not(layer4_outputs(1154));
    outputs(4923) <= (layer4_outputs(3158)) and not (layer4_outputs(10122));
    outputs(4924) <= not(layer4_outputs(3460));
    outputs(4925) <= layer4_outputs(3864);
    outputs(4926) <= (layer4_outputs(521)) and not (layer4_outputs(4235));
    outputs(4927) <= not((layer4_outputs(8500)) xor (layer4_outputs(6923)));
    outputs(4928) <= layer4_outputs(3337);
    outputs(4929) <= layer4_outputs(5002);
    outputs(4930) <= (layer4_outputs(10051)) xor (layer4_outputs(575));
    outputs(4931) <= not(layer4_outputs(6631));
    outputs(4932) <= not((layer4_outputs(2260)) xor (layer4_outputs(9270)));
    outputs(4933) <= not(layer4_outputs(10060));
    outputs(4934) <= not(layer4_outputs(8373));
    outputs(4935) <= not(layer4_outputs(8191));
    outputs(4936) <= layer4_outputs(6321);
    outputs(4937) <= not(layer4_outputs(1479)) or (layer4_outputs(2663));
    outputs(4938) <= (layer4_outputs(5306)) and (layer4_outputs(9989));
    outputs(4939) <= not(layer4_outputs(7841));
    outputs(4940) <= layer4_outputs(2485);
    outputs(4941) <= not(layer4_outputs(6838));
    outputs(4942) <= (layer4_outputs(5545)) xor (layer4_outputs(1497));
    outputs(4943) <= layer4_outputs(6366);
    outputs(4944) <= not((layer4_outputs(3249)) xor (layer4_outputs(1114)));
    outputs(4945) <= not(layer4_outputs(1828));
    outputs(4946) <= (layer4_outputs(5676)) or (layer4_outputs(2483));
    outputs(4947) <= not(layer4_outputs(8831));
    outputs(4948) <= not(layer4_outputs(3682));
    outputs(4949) <= not(layer4_outputs(2097));
    outputs(4950) <= (layer4_outputs(1195)) xor (layer4_outputs(1659));
    outputs(4951) <= layer4_outputs(3470);
    outputs(4952) <= not((layer4_outputs(3786)) xor (layer4_outputs(4876)));
    outputs(4953) <= layer4_outputs(768);
    outputs(4954) <= not((layer4_outputs(9361)) xor (layer4_outputs(1911)));
    outputs(4955) <= not(layer4_outputs(9883));
    outputs(4956) <= not(layer4_outputs(4601));
    outputs(4957) <= layer4_outputs(5606);
    outputs(4958) <= (layer4_outputs(8425)) and (layer4_outputs(1032));
    outputs(4959) <= not(layer4_outputs(7820));
    outputs(4960) <= layer4_outputs(6153);
    outputs(4961) <= layer4_outputs(4558);
    outputs(4962) <= not(layer4_outputs(1751));
    outputs(4963) <= layer4_outputs(3453);
    outputs(4964) <= not(layer4_outputs(6290));
    outputs(4965) <= not(layer4_outputs(4229));
    outputs(4966) <= (layer4_outputs(7376)) xor (layer4_outputs(6867));
    outputs(4967) <= not((layer4_outputs(7229)) xor (layer4_outputs(166)));
    outputs(4968) <= (layer4_outputs(9991)) and (layer4_outputs(7294));
    outputs(4969) <= layer4_outputs(7368);
    outputs(4970) <= not((layer4_outputs(4576)) xor (layer4_outputs(3466)));
    outputs(4971) <= not(layer4_outputs(5654));
    outputs(4972) <= layer4_outputs(6967);
    outputs(4973) <= not((layer4_outputs(195)) or (layer4_outputs(7922)));
    outputs(4974) <= layer4_outputs(3302);
    outputs(4975) <= (layer4_outputs(1551)) xor (layer4_outputs(6663));
    outputs(4976) <= (layer4_outputs(5087)) xor (layer4_outputs(4945));
    outputs(4977) <= not(layer4_outputs(8814)) or (layer4_outputs(9057));
    outputs(4978) <= not(layer4_outputs(2600));
    outputs(4979) <= not(layer4_outputs(1799));
    outputs(4980) <= not((layer4_outputs(6828)) xor (layer4_outputs(8771)));
    outputs(4981) <= not(layer4_outputs(5966));
    outputs(4982) <= not(layer4_outputs(5013));
    outputs(4983) <= layer4_outputs(1384);
    outputs(4984) <= (layer4_outputs(3888)) and not (layer4_outputs(3169));
    outputs(4985) <= (layer4_outputs(733)) and not (layer4_outputs(7593));
    outputs(4986) <= not(layer4_outputs(5333));
    outputs(4987) <= layer4_outputs(4255);
    outputs(4988) <= not((layer4_outputs(3785)) xor (layer4_outputs(7365)));
    outputs(4989) <= not((layer4_outputs(6612)) xor (layer4_outputs(444)));
    outputs(4990) <= (layer4_outputs(559)) xor (layer4_outputs(6610));
    outputs(4991) <= not(layer4_outputs(8833));
    outputs(4992) <= not(layer4_outputs(7321));
    outputs(4993) <= not(layer4_outputs(5576));
    outputs(4994) <= not((layer4_outputs(4393)) xor (layer4_outputs(10137)));
    outputs(4995) <= layer4_outputs(10105);
    outputs(4996) <= not(layer4_outputs(5420)) or (layer4_outputs(5570));
    outputs(4997) <= not(layer4_outputs(1693));
    outputs(4998) <= layer4_outputs(3958);
    outputs(4999) <= not((layer4_outputs(10013)) xor (layer4_outputs(8360)));
    outputs(5000) <= not((layer4_outputs(2861)) xor (layer4_outputs(6809)));
    outputs(5001) <= (layer4_outputs(214)) xor (layer4_outputs(4177));
    outputs(5002) <= not(layer4_outputs(6142));
    outputs(5003) <= not(layer4_outputs(9958));
    outputs(5004) <= layer4_outputs(3754);
    outputs(5005) <= not(layer4_outputs(1364));
    outputs(5006) <= (layer4_outputs(3387)) and (layer4_outputs(2009));
    outputs(5007) <= layer4_outputs(4316);
    outputs(5008) <= layer4_outputs(5851);
    outputs(5009) <= layer4_outputs(2564);
    outputs(5010) <= '1';
    outputs(5011) <= not(layer4_outputs(7930));
    outputs(5012) <= layer4_outputs(7534);
    outputs(5013) <= not(layer4_outputs(8427));
    outputs(5014) <= (layer4_outputs(8463)) and not (layer4_outputs(1569));
    outputs(5015) <= not(layer4_outputs(510));
    outputs(5016) <= not(layer4_outputs(10063));
    outputs(5017) <= not(layer4_outputs(7019));
    outputs(5018) <= not(layer4_outputs(4222));
    outputs(5019) <= layer4_outputs(7572);
    outputs(5020) <= (layer4_outputs(5575)) and not (layer4_outputs(6966));
    outputs(5021) <= not(layer4_outputs(815));
    outputs(5022) <= layer4_outputs(1726);
    outputs(5023) <= not(layer4_outputs(3571));
    outputs(5024) <= (layer4_outputs(3489)) and not (layer4_outputs(7315));
    outputs(5025) <= not(layer4_outputs(10007));
    outputs(5026) <= not(layer4_outputs(708));
    outputs(5027) <= layer4_outputs(9249);
    outputs(5028) <= layer4_outputs(2027);
    outputs(5029) <= layer4_outputs(5467);
    outputs(5030) <= not((layer4_outputs(2992)) xor (layer4_outputs(8117)));
    outputs(5031) <= not((layer4_outputs(8214)) xor (layer4_outputs(45)));
    outputs(5032) <= layer4_outputs(7801);
    outputs(5033) <= layer4_outputs(7756);
    outputs(5034) <= (layer4_outputs(3864)) or (layer4_outputs(8232));
    outputs(5035) <= not(layer4_outputs(3265));
    outputs(5036) <= (layer4_outputs(6287)) xor (layer4_outputs(8686));
    outputs(5037) <= not(layer4_outputs(2938));
    outputs(5038) <= not(layer4_outputs(1301));
    outputs(5039) <= (layer4_outputs(8767)) xor (layer4_outputs(9568));
    outputs(5040) <= not(layer4_outputs(9339));
    outputs(5041) <= (layer4_outputs(1149)) xor (layer4_outputs(6593));
    outputs(5042) <= (layer4_outputs(7621)) xor (layer4_outputs(7177));
    outputs(5043) <= layer4_outputs(8071);
    outputs(5044) <= (layer4_outputs(4656)) and (layer4_outputs(2048));
    outputs(5045) <= layer4_outputs(7540);
    outputs(5046) <= not((layer4_outputs(5058)) xor (layer4_outputs(1070)));
    outputs(5047) <= layer4_outputs(9022);
    outputs(5048) <= not((layer4_outputs(11)) xor (layer4_outputs(8035)));
    outputs(5049) <= layer4_outputs(3032);
    outputs(5050) <= (layer4_outputs(8453)) and (layer4_outputs(2172));
    outputs(5051) <= layer4_outputs(3780);
    outputs(5052) <= not(layer4_outputs(1825));
    outputs(5053) <= layer4_outputs(5334);
    outputs(5054) <= layer4_outputs(8816);
    outputs(5055) <= not(layer4_outputs(5062));
    outputs(5056) <= (layer4_outputs(4265)) and not (layer4_outputs(97));
    outputs(5057) <= layer4_outputs(8283);
    outputs(5058) <= layer4_outputs(5235);
    outputs(5059) <= not(layer4_outputs(10043));
    outputs(5060) <= (layer4_outputs(104)) xor (layer4_outputs(9935));
    outputs(5061) <= not(layer4_outputs(594));
    outputs(5062) <= layer4_outputs(840);
    outputs(5063) <= not(layer4_outputs(8464));
    outputs(5064) <= not((layer4_outputs(295)) or (layer4_outputs(2486)));
    outputs(5065) <= layer4_outputs(8166);
    outputs(5066) <= layer4_outputs(8680);
    outputs(5067) <= layer4_outputs(1131);
    outputs(5068) <= (layer4_outputs(6430)) xor (layer4_outputs(9881));
    outputs(5069) <= not(layer4_outputs(4002));
    outputs(5070) <= layer4_outputs(9853);
    outputs(5071) <= not(layer4_outputs(4236));
    outputs(5072) <= not(layer4_outputs(9467));
    outputs(5073) <= not(layer4_outputs(1277));
    outputs(5074) <= (layer4_outputs(2770)) xor (layer4_outputs(3379));
    outputs(5075) <= layer4_outputs(4273);
    outputs(5076) <= not((layer4_outputs(339)) xor (layer4_outputs(9690)));
    outputs(5077) <= not(layer4_outputs(5209));
    outputs(5078) <= (layer4_outputs(3015)) and not (layer4_outputs(2033));
    outputs(5079) <= not((layer4_outputs(4843)) xor (layer4_outputs(867)));
    outputs(5080) <= (layer4_outputs(1769)) and (layer4_outputs(922));
    outputs(5081) <= not(layer4_outputs(755));
    outputs(5082) <= not(layer4_outputs(4835));
    outputs(5083) <= not((layer4_outputs(3810)) xor (layer4_outputs(2821)));
    outputs(5084) <= layer4_outputs(6265);
    outputs(5085) <= (layer4_outputs(2732)) and (layer4_outputs(5148));
    outputs(5086) <= not(layer4_outputs(8806));
    outputs(5087) <= not(layer4_outputs(9321));
    outputs(5088) <= not(layer4_outputs(10007));
    outputs(5089) <= (layer4_outputs(8563)) xor (layer4_outputs(2349));
    outputs(5090) <= layer4_outputs(8300);
    outputs(5091) <= layer4_outputs(8066);
    outputs(5092) <= not(layer4_outputs(348));
    outputs(5093) <= layer4_outputs(1571);
    outputs(5094) <= layer4_outputs(3319);
    outputs(5095) <= not(layer4_outputs(7988)) or (layer4_outputs(5413));
    outputs(5096) <= not(layer4_outputs(9765));
    outputs(5097) <= layer4_outputs(39);
    outputs(5098) <= (layer4_outputs(1601)) xor (layer4_outputs(1208));
    outputs(5099) <= (layer4_outputs(2656)) xor (layer4_outputs(5461));
    outputs(5100) <= not(layer4_outputs(6466));
    outputs(5101) <= not((layer4_outputs(7095)) xor (layer4_outputs(3450)));
    outputs(5102) <= not(layer4_outputs(8266));
    outputs(5103) <= not(layer4_outputs(8584));
    outputs(5104) <= '1';
    outputs(5105) <= not((layer4_outputs(2258)) xor (layer4_outputs(9256)));
    outputs(5106) <= not(layer4_outputs(3073));
    outputs(5107) <= (layer4_outputs(3505)) and not (layer4_outputs(4365));
    outputs(5108) <= (layer4_outputs(643)) and not (layer4_outputs(4741));
    outputs(5109) <= not(layer4_outputs(5705));
    outputs(5110) <= (layer4_outputs(3314)) xor (layer4_outputs(7913));
    outputs(5111) <= layer4_outputs(7753);
    outputs(5112) <= not(layer4_outputs(5244));
    outputs(5113) <= (layer4_outputs(1411)) xor (layer4_outputs(8819));
    outputs(5114) <= not(layer4_outputs(903));
    outputs(5115) <= (layer4_outputs(7689)) and not (layer4_outputs(4883));
    outputs(5116) <= not((layer4_outputs(9134)) xor (layer4_outputs(3363)));
    outputs(5117) <= layer4_outputs(8340);
    outputs(5118) <= not(layer4_outputs(5028));
    outputs(5119) <= (layer4_outputs(6179)) and not (layer4_outputs(6433));
    outputs(5120) <= not(layer4_outputs(9279));
    outputs(5121) <= (layer4_outputs(686)) and (layer4_outputs(5440));
    outputs(5122) <= not(layer4_outputs(1931));
    outputs(5123) <= (layer4_outputs(1693)) xor (layer4_outputs(3349));
    outputs(5124) <= not(layer4_outputs(7106));
    outputs(5125) <= not((layer4_outputs(4813)) or (layer4_outputs(626)));
    outputs(5126) <= not(layer4_outputs(9527)) or (layer4_outputs(3228));
    outputs(5127) <= layer4_outputs(6008);
    outputs(5128) <= (layer4_outputs(2252)) xor (layer4_outputs(4388));
    outputs(5129) <= layer4_outputs(3139);
    outputs(5130) <= not(layer4_outputs(7220));
    outputs(5131) <= not(layer4_outputs(982));
    outputs(5132) <= not((layer4_outputs(4782)) xor (layer4_outputs(6842)));
    outputs(5133) <= layer4_outputs(2592);
    outputs(5134) <= layer4_outputs(3768);
    outputs(5135) <= not((layer4_outputs(9535)) xor (layer4_outputs(5497)));
    outputs(5136) <= not((layer4_outputs(10196)) xor (layer4_outputs(4797)));
    outputs(5137) <= layer4_outputs(7504);
    outputs(5138) <= layer4_outputs(899);
    outputs(5139) <= (layer4_outputs(6724)) xor (layer4_outputs(7575));
    outputs(5140) <= not((layer4_outputs(8995)) xor (layer4_outputs(7214)));
    outputs(5141) <= (layer4_outputs(4511)) and (layer4_outputs(4975));
    outputs(5142) <= not(layer4_outputs(7001));
    outputs(5143) <= not(layer4_outputs(4350));
    outputs(5144) <= layer4_outputs(9037);
    outputs(5145) <= (layer4_outputs(3861)) xor (layer4_outputs(7410));
    outputs(5146) <= layer4_outputs(6401);
    outputs(5147) <= not((layer4_outputs(2224)) xor (layer4_outputs(4783)));
    outputs(5148) <= not(layer4_outputs(5986));
    outputs(5149) <= not((layer4_outputs(3540)) xor (layer4_outputs(8632)));
    outputs(5150) <= layer4_outputs(1941);
    outputs(5151) <= layer4_outputs(4082);
    outputs(5152) <= not((layer4_outputs(8321)) xor (layer4_outputs(6637)));
    outputs(5153) <= not((layer4_outputs(5196)) xor (layer4_outputs(8433)));
    outputs(5154) <= (layer4_outputs(3227)) xor (layer4_outputs(9777));
    outputs(5155) <= (layer4_outputs(1181)) xor (layer4_outputs(9252));
    outputs(5156) <= layer4_outputs(7753);
    outputs(5157) <= not(layer4_outputs(1784));
    outputs(5158) <= layer4_outputs(273);
    outputs(5159) <= not(layer4_outputs(10211));
    outputs(5160) <= (layer4_outputs(7842)) xor (layer4_outputs(7272));
    outputs(5161) <= not((layer4_outputs(9011)) xor (layer4_outputs(3309)));
    outputs(5162) <= not(layer4_outputs(5850));
    outputs(5163) <= layer4_outputs(2446);
    outputs(5164) <= layer4_outputs(1903);
    outputs(5165) <= layer4_outputs(8489);
    outputs(5166) <= (layer4_outputs(2609)) xor (layer4_outputs(508));
    outputs(5167) <= (layer4_outputs(865)) xor (layer4_outputs(8652));
    outputs(5168) <= not((layer4_outputs(9975)) xor (layer4_outputs(8240)));
    outputs(5169) <= not(layer4_outputs(9806));
    outputs(5170) <= not(layer4_outputs(7714));
    outputs(5171) <= (layer4_outputs(9023)) xor (layer4_outputs(6057));
    outputs(5172) <= layer4_outputs(4486);
    outputs(5173) <= layer4_outputs(3471);
    outputs(5174) <= layer4_outputs(4370);
    outputs(5175) <= not((layer4_outputs(2517)) xor (layer4_outputs(3059)));
    outputs(5176) <= not((layer4_outputs(5694)) xor (layer4_outputs(4599)));
    outputs(5177) <= (layer4_outputs(3742)) xor (layer4_outputs(5545));
    outputs(5178) <= (layer4_outputs(706)) xor (layer4_outputs(2393));
    outputs(5179) <= not(layer4_outputs(742));
    outputs(5180) <= layer4_outputs(8227);
    outputs(5181) <= not(layer4_outputs(8522));
    outputs(5182) <= not(layer4_outputs(5107));
    outputs(5183) <= not((layer4_outputs(4017)) xor (layer4_outputs(8802)));
    outputs(5184) <= layer4_outputs(5487);
    outputs(5185) <= not((layer4_outputs(7339)) xor (layer4_outputs(171)));
    outputs(5186) <= (layer4_outputs(5753)) xor (layer4_outputs(1315));
    outputs(5187) <= (layer4_outputs(1812)) xor (layer4_outputs(3179));
    outputs(5188) <= (layer4_outputs(7309)) and not (layer4_outputs(3761));
    outputs(5189) <= layer4_outputs(6635);
    outputs(5190) <= layer4_outputs(6868);
    outputs(5191) <= layer4_outputs(9077);
    outputs(5192) <= not((layer4_outputs(8797)) xor (layer4_outputs(2971)));
    outputs(5193) <= layer4_outputs(6412);
    outputs(5194) <= (layer4_outputs(6486)) and not (layer4_outputs(4788));
    outputs(5195) <= (layer4_outputs(2633)) xor (layer4_outputs(4457));
    outputs(5196) <= not(layer4_outputs(1300));
    outputs(5197) <= not(layer4_outputs(216));
    outputs(5198) <= not(layer4_outputs(4775));
    outputs(5199) <= not(layer4_outputs(4519));
    outputs(5200) <= (layer4_outputs(1678)) xor (layer4_outputs(9179));
    outputs(5201) <= (layer4_outputs(5499)) xor (layer4_outputs(3252));
    outputs(5202) <= not((layer4_outputs(9692)) xor (layer4_outputs(7248)));
    outputs(5203) <= not(layer4_outputs(5786));
    outputs(5204) <= layer4_outputs(6140);
    outputs(5205) <= not((layer4_outputs(8656)) xor (layer4_outputs(4857)));
    outputs(5206) <= (layer4_outputs(10106)) xor (layer4_outputs(4716));
    outputs(5207) <= not(layer4_outputs(5892));
    outputs(5208) <= layer4_outputs(10161);
    outputs(5209) <= (layer4_outputs(1851)) xor (layer4_outputs(9009));
    outputs(5210) <= not(layer4_outputs(2567)) or (layer4_outputs(6888));
    outputs(5211) <= layer4_outputs(1015);
    outputs(5212) <= layer4_outputs(7042);
    outputs(5213) <= not((layer4_outputs(3936)) xor (layer4_outputs(7257)));
    outputs(5214) <= not(layer4_outputs(3746));
    outputs(5215) <= not(layer4_outputs(8477));
    outputs(5216) <= layer4_outputs(6296);
    outputs(5217) <= (layer4_outputs(2266)) and (layer4_outputs(10138));
    outputs(5218) <= layer4_outputs(7532);
    outputs(5219) <= not(layer4_outputs(6163));
    outputs(5220) <= layer4_outputs(9648);
    outputs(5221) <= layer4_outputs(2998);
    outputs(5222) <= not(layer4_outputs(5378));
    outputs(5223) <= not(layer4_outputs(8938));
    outputs(5224) <= (layer4_outputs(3755)) and not (layer4_outputs(6485));
    outputs(5225) <= layer4_outputs(5346);
    outputs(5226) <= not(layer4_outputs(7859));
    outputs(5227) <= not((layer4_outputs(5252)) xor (layer4_outputs(3628)));
    outputs(5228) <= layer4_outputs(3706);
    outputs(5229) <= not((layer4_outputs(1789)) xor (layer4_outputs(10046)));
    outputs(5230) <= (layer4_outputs(9686)) xor (layer4_outputs(4900));
    outputs(5231) <= layer4_outputs(4830);
    outputs(5232) <= not((layer4_outputs(139)) xor (layer4_outputs(8809)));
    outputs(5233) <= not((layer4_outputs(6048)) xor (layer4_outputs(6468)));
    outputs(5234) <= not(layer4_outputs(3497));
    outputs(5235) <= layer4_outputs(9384);
    outputs(5236) <= layer4_outputs(5521);
    outputs(5237) <= not(layer4_outputs(3772)) or (layer4_outputs(2774));
    outputs(5238) <= layer4_outputs(3108);
    outputs(5239) <= not(layer4_outputs(6853));
    outputs(5240) <= not((layer4_outputs(5823)) xor (layer4_outputs(4792)));
    outputs(5241) <= layer4_outputs(6099);
    outputs(5242) <= (layer4_outputs(7868)) xor (layer4_outputs(8018));
    outputs(5243) <= not(layer4_outputs(2574));
    outputs(5244) <= not(layer4_outputs(6012));
    outputs(5245) <= layer4_outputs(4665);
    outputs(5246) <= not(layer4_outputs(5341));
    outputs(5247) <= not(layer4_outputs(10067));
    outputs(5248) <= not(layer4_outputs(4533));
    outputs(5249) <= (layer4_outputs(4726)) and not (layer4_outputs(3623));
    outputs(5250) <= not(layer4_outputs(7135));
    outputs(5251) <= layer4_outputs(7487);
    outputs(5252) <= layer4_outputs(95);
    outputs(5253) <= not(layer4_outputs(7038)) or (layer4_outputs(8513));
    outputs(5254) <= not((layer4_outputs(1775)) or (layer4_outputs(1552)));
    outputs(5255) <= not((layer4_outputs(6360)) and (layer4_outputs(3438)));
    outputs(5256) <= (layer4_outputs(2263)) xor (layer4_outputs(10156));
    outputs(5257) <= layer4_outputs(1991);
    outputs(5258) <= (layer4_outputs(1385)) and not (layer4_outputs(9960));
    outputs(5259) <= not((layer4_outputs(2793)) xor (layer4_outputs(3563)));
    outputs(5260) <= layer4_outputs(955);
    outputs(5261) <= not((layer4_outputs(7249)) xor (layer4_outputs(5256)));
    outputs(5262) <= (layer4_outputs(4248)) xor (layer4_outputs(2179));
    outputs(5263) <= not(layer4_outputs(505));
    outputs(5264) <= (layer4_outputs(6360)) xor (layer4_outputs(8129));
    outputs(5265) <= (layer4_outputs(2288)) xor (layer4_outputs(6216));
    outputs(5266) <= (layer4_outputs(9553)) or (layer4_outputs(1548));
    outputs(5267) <= (layer4_outputs(2072)) xor (layer4_outputs(6085));
    outputs(5268) <= not((layer4_outputs(6683)) or (layer4_outputs(6547)));
    outputs(5269) <= not((layer4_outputs(6418)) xor (layer4_outputs(8172)));
    outputs(5270) <= not(layer4_outputs(33));
    outputs(5271) <= (layer4_outputs(4643)) xor (layer4_outputs(3717));
    outputs(5272) <= not((layer4_outputs(153)) or (layer4_outputs(8380)));
    outputs(5273) <= (layer4_outputs(10179)) or (layer4_outputs(9961));
    outputs(5274) <= (layer4_outputs(6918)) xor (layer4_outputs(2852));
    outputs(5275) <= not(layer4_outputs(1216));
    outputs(5276) <= not(layer4_outputs(2455));
    outputs(5277) <= not(layer4_outputs(4862));
    outputs(5278) <= layer4_outputs(3295);
    outputs(5279) <= layer4_outputs(8634);
    outputs(5280) <= not(layer4_outputs(5340));
    outputs(5281) <= not((layer4_outputs(2173)) xor (layer4_outputs(2372)));
    outputs(5282) <= not((layer4_outputs(1152)) or (layer4_outputs(5941)));
    outputs(5283) <= not((layer4_outputs(6214)) xor (layer4_outputs(9507)));
    outputs(5284) <= layer4_outputs(4593);
    outputs(5285) <= layer4_outputs(6951);
    outputs(5286) <= not(layer4_outputs(6117));
    outputs(5287) <= (layer4_outputs(7041)) xor (layer4_outputs(2818));
    outputs(5288) <= not((layer4_outputs(1905)) xor (layer4_outputs(555)));
    outputs(5289) <= not(layer4_outputs(9864));
    outputs(5290) <= layer4_outputs(7921);
    outputs(5291) <= not(layer4_outputs(2982));
    outputs(5292) <= (layer4_outputs(6090)) or (layer4_outputs(4097));
    outputs(5293) <= (layer4_outputs(9500)) xor (layer4_outputs(3475));
    outputs(5294) <= '1';
    outputs(5295) <= not(layer4_outputs(403));
    outputs(5296) <= not((layer4_outputs(9325)) xor (layer4_outputs(244)));
    outputs(5297) <= not((layer4_outputs(4955)) xor (layer4_outputs(9729)));
    outputs(5298) <= not(layer4_outputs(1854));
    outputs(5299) <= layer4_outputs(156);
    outputs(5300) <= layer4_outputs(10057);
    outputs(5301) <= not(layer4_outputs(6513));
    outputs(5302) <= (layer4_outputs(1678)) xor (layer4_outputs(515));
    outputs(5303) <= not((layer4_outputs(5222)) xor (layer4_outputs(294)));
    outputs(5304) <= not((layer4_outputs(3608)) xor (layer4_outputs(3789)));
    outputs(5305) <= not(layer4_outputs(2901));
    outputs(5306) <= layer4_outputs(8163);
    outputs(5307) <= not((layer4_outputs(6136)) xor (layer4_outputs(3074)));
    outputs(5308) <= not(layer4_outputs(4943));
    outputs(5309) <= (layer4_outputs(4110)) or (layer4_outputs(6465));
    outputs(5310) <= not((layer4_outputs(5501)) xor (layer4_outputs(8259)));
    outputs(5311) <= not((layer4_outputs(2403)) xor (layer4_outputs(9884)));
    outputs(5312) <= not(layer4_outputs(2786));
    outputs(5313) <= not(layer4_outputs(343));
    outputs(5314) <= (layer4_outputs(1969)) and (layer4_outputs(8502));
    outputs(5315) <= (layer4_outputs(836)) xor (layer4_outputs(796));
    outputs(5316) <= layer4_outputs(3085);
    outputs(5317) <= (layer4_outputs(5054)) xor (layer4_outputs(5770));
    outputs(5318) <= not((layer4_outputs(3209)) and (layer4_outputs(9365)));
    outputs(5319) <= (layer4_outputs(1565)) xor (layer4_outputs(3656));
    outputs(5320) <= layer4_outputs(3328);
    outputs(5321) <= not((layer4_outputs(7924)) xor (layer4_outputs(4554)));
    outputs(5322) <= layer4_outputs(8085);
    outputs(5323) <= layer4_outputs(18);
    outputs(5324) <= not(layer4_outputs(5773));
    outputs(5325) <= layer4_outputs(4045);
    outputs(5326) <= layer4_outputs(1901);
    outputs(5327) <= layer4_outputs(5354);
    outputs(5328) <= not(layer4_outputs(4752));
    outputs(5329) <= not(layer4_outputs(6663));
    outputs(5330) <= (layer4_outputs(3475)) xor (layer4_outputs(2159));
    outputs(5331) <= '1';
    outputs(5332) <= not((layer4_outputs(5777)) xor (layer4_outputs(2282)));
    outputs(5333) <= not(layer4_outputs(3939));
    outputs(5334) <= (layer4_outputs(518)) and (layer4_outputs(1800));
    outputs(5335) <= not((layer4_outputs(1220)) xor (layer4_outputs(2706)));
    outputs(5336) <= not(layer4_outputs(8994));
    outputs(5337) <= not(layer4_outputs(3977));
    outputs(5338) <= not(layer4_outputs(6402));
    outputs(5339) <= (layer4_outputs(5629)) xor (layer4_outputs(2354));
    outputs(5340) <= layer4_outputs(3318);
    outputs(5341) <= not(layer4_outputs(1454)) or (layer4_outputs(6876));
    outputs(5342) <= not(layer4_outputs(6761));
    outputs(5343) <= not(layer4_outputs(4226));
    outputs(5344) <= not((layer4_outputs(4947)) xor (layer4_outputs(8303)));
    outputs(5345) <= not((layer4_outputs(2330)) xor (layer4_outputs(9626)));
    outputs(5346) <= (layer4_outputs(7405)) xor (layer4_outputs(1185));
    outputs(5347) <= (layer4_outputs(3464)) xor (layer4_outputs(2825));
    outputs(5348) <= not(layer4_outputs(4113));
    outputs(5349) <= layer4_outputs(3862);
    outputs(5350) <= layer4_outputs(5078);
    outputs(5351) <= not(layer4_outputs(5917));
    outputs(5352) <= layer4_outputs(79);
    outputs(5353) <= not(layer4_outputs(6858));
    outputs(5354) <= (layer4_outputs(2060)) xor (layer4_outputs(1527));
    outputs(5355) <= (layer4_outputs(8642)) xor (layer4_outputs(3613));
    outputs(5356) <= not(layer4_outputs(2827)) or (layer4_outputs(4036));
    outputs(5357) <= (layer4_outputs(7490)) xor (layer4_outputs(9164));
    outputs(5358) <= not((layer4_outputs(9928)) xor (layer4_outputs(5282)));
    outputs(5359) <= (layer4_outputs(1295)) xor (layer4_outputs(6755));
    outputs(5360) <= layer4_outputs(9013);
    outputs(5361) <= layer4_outputs(8905);
    outputs(5362) <= not(layer4_outputs(4756));
    outputs(5363) <= not(layer4_outputs(4065)) or (layer4_outputs(5675));
    outputs(5364) <= layer4_outputs(444);
    outputs(5365) <= layer4_outputs(9459);
    outputs(5366) <= layer4_outputs(7477);
    outputs(5367) <= not((layer4_outputs(3573)) xor (layer4_outputs(3367)));
    outputs(5368) <= not((layer4_outputs(3077)) xor (layer4_outputs(1480)));
    outputs(5369) <= (layer4_outputs(8407)) xor (layer4_outputs(9988));
    outputs(5370) <= layer4_outputs(8946);
    outputs(5371) <= layer4_outputs(5672);
    outputs(5372) <= not(layer4_outputs(8747));
    outputs(5373) <= '1';
    outputs(5374) <= not((layer4_outputs(4539)) or (layer4_outputs(9632)));
    outputs(5375) <= layer4_outputs(8474);
    outputs(5376) <= (layer4_outputs(7527)) xor (layer4_outputs(6045));
    outputs(5377) <= not(layer4_outputs(2176));
    outputs(5378) <= not(layer4_outputs(9642));
    outputs(5379) <= layer4_outputs(7788);
    outputs(5380) <= not((layer4_outputs(5082)) xor (layer4_outputs(9871)));
    outputs(5381) <= not(layer4_outputs(8876));
    outputs(5382) <= not((layer4_outputs(3410)) xor (layer4_outputs(1265)));
    outputs(5383) <= not(layer4_outputs(9326));
    outputs(5384) <= not(layer4_outputs(8848));
    outputs(5385) <= not(layer4_outputs(1448));
    outputs(5386) <= not((layer4_outputs(8102)) xor (layer4_outputs(787)));
    outputs(5387) <= layer4_outputs(9086);
    outputs(5388) <= layer4_outputs(3330);
    outputs(5389) <= layer4_outputs(1341);
    outputs(5390) <= not((layer4_outputs(5595)) xor (layer4_outputs(4563)));
    outputs(5391) <= (layer4_outputs(210)) and not (layer4_outputs(7650));
    outputs(5392) <= (layer4_outputs(4915)) xor (layer4_outputs(5707));
    outputs(5393) <= not((layer4_outputs(7683)) xor (layer4_outputs(1883)));
    outputs(5394) <= not((layer4_outputs(8448)) and (layer4_outputs(8743)));
    outputs(5395) <= (layer4_outputs(5522)) or (layer4_outputs(4908));
    outputs(5396) <= layer4_outputs(758);
    outputs(5397) <= layer4_outputs(3478);
    outputs(5398) <= layer4_outputs(4449);
    outputs(5399) <= not(layer4_outputs(6989));
    outputs(5400) <= not(layer4_outputs(6810));
    outputs(5401) <= (layer4_outputs(7237)) and (layer4_outputs(3589));
    outputs(5402) <= not(layer4_outputs(9177));
    outputs(5403) <= layer4_outputs(5415);
    outputs(5404) <= (layer4_outputs(4605)) xor (layer4_outputs(6210));
    outputs(5405) <= (layer4_outputs(10036)) and not (layer4_outputs(8479));
    outputs(5406) <= layer4_outputs(7210);
    outputs(5407) <= (layer4_outputs(8364)) xor (layer4_outputs(9960));
    outputs(5408) <= not(layer4_outputs(420));
    outputs(5409) <= not(layer4_outputs(8446));
    outputs(5410) <= (layer4_outputs(7506)) xor (layer4_outputs(9190));
    outputs(5411) <= not(layer4_outputs(496)) or (layer4_outputs(4120));
    outputs(5412) <= not((layer4_outputs(4962)) xor (layer4_outputs(7955)));
    outputs(5413) <= not((layer4_outputs(2549)) and (layer4_outputs(9730)));
    outputs(5414) <= not(layer4_outputs(4114));
    outputs(5415) <= (layer4_outputs(9823)) xor (layer4_outputs(5855));
    outputs(5416) <= (layer4_outputs(2580)) xor (layer4_outputs(9712));
    outputs(5417) <= layer4_outputs(7653);
    outputs(5418) <= layer4_outputs(1348);
    outputs(5419) <= not((layer4_outputs(4706)) and (layer4_outputs(8236)));
    outputs(5420) <= not(layer4_outputs(8238));
    outputs(5421) <= not(layer4_outputs(3913)) or (layer4_outputs(379));
    outputs(5422) <= layer4_outputs(2038);
    outputs(5423) <= not(layer4_outputs(2917));
    outputs(5424) <= layer4_outputs(6028);
    outputs(5425) <= (layer4_outputs(2465)) or (layer4_outputs(999));
    outputs(5426) <= not(layer4_outputs(8590)) or (layer4_outputs(3665));
    outputs(5427) <= layer4_outputs(8051);
    outputs(5428) <= (layer4_outputs(7290)) xor (layer4_outputs(6115));
    outputs(5429) <= (layer4_outputs(6831)) and (layer4_outputs(7883));
    outputs(5430) <= (layer4_outputs(10172)) and not (layer4_outputs(1069));
    outputs(5431) <= layer4_outputs(7236);
    outputs(5432) <= not(layer4_outputs(2712));
    outputs(5433) <= layer4_outputs(4968);
    outputs(5434) <= layer4_outputs(9305);
    outputs(5435) <= layer4_outputs(7986);
    outputs(5436) <= layer4_outputs(3834);
    outputs(5437) <= not((layer4_outputs(7737)) xor (layer4_outputs(6225)));
    outputs(5438) <= (layer4_outputs(6042)) or (layer4_outputs(1810));
    outputs(5439) <= (layer4_outputs(1553)) xor (layer4_outputs(9454));
    outputs(5440) <= (layer4_outputs(7077)) and (layer4_outputs(7935));
    outputs(5441) <= (layer4_outputs(3136)) and (layer4_outputs(5836));
    outputs(5442) <= not((layer4_outputs(4952)) xor (layer4_outputs(10070)));
    outputs(5443) <= not((layer4_outputs(2957)) and (layer4_outputs(5464)));
    outputs(5444) <= layer4_outputs(282);
    outputs(5445) <= not(layer4_outputs(3945));
    outputs(5446) <= (layer4_outputs(6558)) xor (layer4_outputs(7022));
    outputs(5447) <= layer4_outputs(2016);
    outputs(5448) <= not((layer4_outputs(6654)) xor (layer4_outputs(9801)));
    outputs(5449) <= not((layer4_outputs(4422)) xor (layer4_outputs(8584)));
    outputs(5450) <= layer4_outputs(1558);
    outputs(5451) <= not((layer4_outputs(10098)) xor (layer4_outputs(4317)));
    outputs(5452) <= (layer4_outputs(2375)) xor (layer4_outputs(4376));
    outputs(5453) <= not(layer4_outputs(6059)) or (layer4_outputs(5318));
    outputs(5454) <= (layer4_outputs(3845)) xor (layer4_outputs(5022));
    outputs(5455) <= not(layer4_outputs(4169));
    outputs(5456) <= (layer4_outputs(5260)) and (layer4_outputs(199));
    outputs(5457) <= layer4_outputs(8542);
    outputs(5458) <= not(layer4_outputs(4059));
    outputs(5459) <= (layer4_outputs(1428)) xor (layer4_outputs(5161));
    outputs(5460) <= not((layer4_outputs(10095)) xor (layer4_outputs(9940)));
    outputs(5461) <= not((layer4_outputs(4399)) xor (layer4_outputs(1284)));
    outputs(5462) <= (layer4_outputs(2939)) xor (layer4_outputs(7518));
    outputs(5463) <= not((layer4_outputs(7740)) xor (layer4_outputs(2627)));
    outputs(5464) <= layer4_outputs(3412);
    outputs(5465) <= not(layer4_outputs(6809));
    outputs(5466) <= layer4_outputs(6329);
    outputs(5467) <= not(layer4_outputs(7250));
    outputs(5468) <= not(layer4_outputs(348));
    outputs(5469) <= not(layer4_outputs(5382));
    outputs(5470) <= layer4_outputs(1869);
    outputs(5471) <= not(layer4_outputs(4907));
    outputs(5472) <= (layer4_outputs(8374)) and not (layer4_outputs(9250));
    outputs(5473) <= layer4_outputs(4433);
    outputs(5474) <= layer4_outputs(4591);
    outputs(5475) <= layer4_outputs(2790);
    outputs(5476) <= layer4_outputs(8887);
    outputs(5477) <= not(layer4_outputs(459));
    outputs(5478) <= (layer4_outputs(7526)) and not (layer4_outputs(7611));
    outputs(5479) <= (layer4_outputs(4695)) xor (layer4_outputs(6314));
    outputs(5480) <= layer4_outputs(9814);
    outputs(5481) <= not((layer4_outputs(8464)) xor (layer4_outputs(1239)));
    outputs(5482) <= (layer4_outputs(3132)) xor (layer4_outputs(4346));
    outputs(5483) <= not(layer4_outputs(8834));
    outputs(5484) <= not(layer4_outputs(2775));
    outputs(5485) <= layer4_outputs(3493);
    outputs(5486) <= not(layer4_outputs(9370));
    outputs(5487) <= layer4_outputs(6159);
    outputs(5488) <= not((layer4_outputs(3113)) xor (layer4_outputs(4275)));
    outputs(5489) <= not(layer4_outputs(5058));
    outputs(5490) <= not(layer4_outputs(2586));
    outputs(5491) <= not(layer4_outputs(1316));
    outputs(5492) <= not((layer4_outputs(5826)) xor (layer4_outputs(2287)));
    outputs(5493) <= (layer4_outputs(9360)) and not (layer4_outputs(5949));
    outputs(5494) <= (layer4_outputs(9328)) xor (layer4_outputs(694));
    outputs(5495) <= not(layer4_outputs(384));
    outputs(5496) <= not(layer4_outputs(3984));
    outputs(5497) <= not(layer4_outputs(14));
    outputs(5498) <= not(layer4_outputs(8797));
    outputs(5499) <= (layer4_outputs(4273)) xor (layer4_outputs(6614));
    outputs(5500) <= layer4_outputs(2795);
    outputs(5501) <= (layer4_outputs(10116)) xor (layer4_outputs(1354));
    outputs(5502) <= not(layer4_outputs(875));
    outputs(5503) <= layer4_outputs(6007);
    outputs(5504) <= not(layer4_outputs(5701)) or (layer4_outputs(73));
    outputs(5505) <= (layer4_outputs(5937)) xor (layer4_outputs(9511));
    outputs(5506) <= not((layer4_outputs(6759)) xor (layer4_outputs(5672)));
    outputs(5507) <= not((layer4_outputs(4488)) xor (layer4_outputs(6329)));
    outputs(5508) <= (layer4_outputs(5906)) xor (layer4_outputs(8145));
    outputs(5509) <= not(layer4_outputs(3836));
    outputs(5510) <= (layer4_outputs(574)) and not (layer4_outputs(1496));
    outputs(5511) <= not((layer4_outputs(2748)) and (layer4_outputs(5220)));
    outputs(5512) <= not(layer4_outputs(4796));
    outputs(5513) <= not((layer4_outputs(6239)) xor (layer4_outputs(2317)));
    outputs(5514) <= (layer4_outputs(1975)) and not (layer4_outputs(1622));
    outputs(5515) <= (layer4_outputs(3876)) and (layer4_outputs(3271));
    outputs(5516) <= layer4_outputs(4534);
    outputs(5517) <= layer4_outputs(1828);
    outputs(5518) <= not(layer4_outputs(7639)) or (layer4_outputs(6855));
    outputs(5519) <= not(layer4_outputs(4338));
    outputs(5520) <= not((layer4_outputs(9685)) xor (layer4_outputs(2080)));
    outputs(5521) <= not((layer4_outputs(2920)) and (layer4_outputs(2425)));
    outputs(5522) <= layer4_outputs(9762);
    outputs(5523) <= (layer4_outputs(9335)) xor (layer4_outputs(10117));
    outputs(5524) <= not(layer4_outputs(402));
    outputs(5525) <= (layer4_outputs(7200)) and (layer4_outputs(6091));
    outputs(5526) <= not(layer4_outputs(716));
    outputs(5527) <= (layer4_outputs(5168)) and not (layer4_outputs(4548));
    outputs(5528) <= layer4_outputs(2590);
    outputs(5529) <= not(layer4_outputs(5537));
    outputs(5530) <= not((layer4_outputs(7234)) xor (layer4_outputs(3219)));
    outputs(5531) <= not((layer4_outputs(8111)) xor (layer4_outputs(6002)));
    outputs(5532) <= not((layer4_outputs(8037)) xor (layer4_outputs(901)));
    outputs(5533) <= not(layer4_outputs(7049));
    outputs(5534) <= layer4_outputs(1677);
    outputs(5535) <= layer4_outputs(2031);
    outputs(5536) <= (layer4_outputs(5114)) and not (layer4_outputs(1843));
    outputs(5537) <= not((layer4_outputs(9120)) xor (layer4_outputs(7215)));
    outputs(5538) <= (layer4_outputs(5411)) and not (layer4_outputs(7330));
    outputs(5539) <= (layer4_outputs(7000)) xor (layer4_outputs(1270));
    outputs(5540) <= (layer4_outputs(6548)) xor (layer4_outputs(3536));
    outputs(5541) <= not(layer4_outputs(5963));
    outputs(5542) <= not(layer4_outputs(4001));
    outputs(5543) <= (layer4_outputs(4458)) or (layer4_outputs(6390));
    outputs(5544) <= not((layer4_outputs(2382)) and (layer4_outputs(261)));
    outputs(5545) <= layer4_outputs(4351);
    outputs(5546) <= layer4_outputs(8151);
    outputs(5547) <= not((layer4_outputs(8659)) xor (layer4_outputs(4382)));
    outputs(5548) <= not((layer4_outputs(3217)) xor (layer4_outputs(4657)));
    outputs(5549) <= layer4_outputs(7341);
    outputs(5550) <= not(layer4_outputs(9652));
    outputs(5551) <= layer4_outputs(917);
    outputs(5552) <= not((layer4_outputs(2937)) xor (layer4_outputs(8365)));
    outputs(5553) <= not(layer4_outputs(6119));
    outputs(5554) <= not((layer4_outputs(8042)) xor (layer4_outputs(853)));
    outputs(5555) <= not((layer4_outputs(9503)) or (layer4_outputs(2749)));
    outputs(5556) <= not(layer4_outputs(4018));
    outputs(5557) <= not((layer4_outputs(2443)) xor (layer4_outputs(1233)));
    outputs(5558) <= not((layer4_outputs(6147)) xor (layer4_outputs(784)));
    outputs(5559) <= layer4_outputs(4887);
    outputs(5560) <= layer4_outputs(5207);
    outputs(5561) <= not(layer4_outputs(8309));
    outputs(5562) <= not(layer4_outputs(6118));
    outputs(5563) <= not(layer4_outputs(6309)) or (layer4_outputs(3740));
    outputs(5564) <= (layer4_outputs(1176)) or (layer4_outputs(1606));
    outputs(5565) <= layer4_outputs(2606);
    outputs(5566) <= (layer4_outputs(5399)) xor (layer4_outputs(2666));
    outputs(5567) <= not((layer4_outputs(2532)) xor (layer4_outputs(8463)));
    outputs(5568) <= not((layer4_outputs(4914)) xor (layer4_outputs(7466)));
    outputs(5569) <= (layer4_outputs(8979)) xor (layer4_outputs(302));
    outputs(5570) <= layer4_outputs(2773);
    outputs(5571) <= not(layer4_outputs(8914));
    outputs(5572) <= (layer4_outputs(5988)) xor (layer4_outputs(7698));
    outputs(5573) <= not(layer4_outputs(5042));
    outputs(5574) <= layer4_outputs(9998);
    outputs(5575) <= layer4_outputs(1644);
    outputs(5576) <= layer4_outputs(1920);
    outputs(5577) <= not((layer4_outputs(7967)) and (layer4_outputs(8088)));
    outputs(5578) <= not(layer4_outputs(5165));
    outputs(5579) <= (layer4_outputs(3753)) and not (layer4_outputs(3031));
    outputs(5580) <= (layer4_outputs(7255)) and (layer4_outputs(9189));
    outputs(5581) <= not(layer4_outputs(3397));
    outputs(5582) <= (layer4_outputs(6576)) xor (layer4_outputs(7346));
    outputs(5583) <= (layer4_outputs(4972)) xor (layer4_outputs(5700));
    outputs(5584) <= layer4_outputs(3270);
    outputs(5585) <= (layer4_outputs(6446)) xor (layer4_outputs(1607));
    outputs(5586) <= not(layer4_outputs(5192));
    outputs(5587) <= not((layer4_outputs(5723)) xor (layer4_outputs(4540)));
    outputs(5588) <= not(layer4_outputs(1419));
    outputs(5589) <= layer4_outputs(9835);
    outputs(5590) <= not((layer4_outputs(9654)) xor (layer4_outputs(9775)));
    outputs(5591) <= layer4_outputs(617);
    outputs(5592) <= (layer4_outputs(5445)) xor (layer4_outputs(8993));
    outputs(5593) <= (layer4_outputs(7407)) xor (layer4_outputs(6211));
    outputs(5594) <= not((layer4_outputs(1244)) xor (layer4_outputs(2829)));
    outputs(5595) <= not((layer4_outputs(972)) xor (layer4_outputs(2896)));
    outputs(5596) <= (layer4_outputs(5924)) xor (layer4_outputs(8387));
    outputs(5597) <= not(layer4_outputs(565));
    outputs(5598) <= not((layer4_outputs(4670)) xor (layer4_outputs(6607)));
    outputs(5599) <= (layer4_outputs(6326)) xor (layer4_outputs(9017));
    outputs(5600) <= not(layer4_outputs(9393));
    outputs(5601) <= not((layer4_outputs(2048)) or (layer4_outputs(2649)));
    outputs(5602) <= not((layer4_outputs(2680)) xor (layer4_outputs(6561)));
    outputs(5603) <= not(layer4_outputs(1914)) or (layer4_outputs(7350));
    outputs(5604) <= layer4_outputs(7251);
    outputs(5605) <= (layer4_outputs(5149)) and not (layer4_outputs(2930));
    outputs(5606) <= layer4_outputs(5430);
    outputs(5607) <= (layer4_outputs(1085)) or (layer4_outputs(6930));
    outputs(5608) <= not(layer4_outputs(6769));
    outputs(5609) <= not(layer4_outputs(5492));
    outputs(5610) <= (layer4_outputs(8021)) and (layer4_outputs(5923));
    outputs(5611) <= (layer4_outputs(1902)) or (layer4_outputs(3856));
    outputs(5612) <= not(layer4_outputs(7580));
    outputs(5613) <= (layer4_outputs(6721)) xor (layer4_outputs(7660));
    outputs(5614) <= (layer4_outputs(5992)) and (layer4_outputs(6202));
    outputs(5615) <= (layer4_outputs(731)) xor (layer4_outputs(1855));
    outputs(5616) <= layer4_outputs(6046);
    outputs(5617) <= layer4_outputs(8171);
    outputs(5618) <= not((layer4_outputs(7451)) xor (layer4_outputs(7087)));
    outputs(5619) <= layer4_outputs(3494);
    outputs(5620) <= not((layer4_outputs(1643)) xor (layer4_outputs(4522)));
    outputs(5621) <= not(layer4_outputs(5687));
    outputs(5622) <= layer4_outputs(2756);
    outputs(5623) <= layer4_outputs(7109);
    outputs(5624) <= not(layer4_outputs(2633));
    outputs(5625) <= not((layer4_outputs(4561)) and (layer4_outputs(8222)));
    outputs(5626) <= not((layer4_outputs(5343)) xor (layer4_outputs(9050)));
    outputs(5627) <= layer4_outputs(518);
    outputs(5628) <= layer4_outputs(4809);
    outputs(5629) <= not((layer4_outputs(6634)) xor (layer4_outputs(124)));
    outputs(5630) <= (layer4_outputs(2977)) or (layer4_outputs(3205));
    outputs(5631) <= (layer4_outputs(6417)) xor (layer4_outputs(5192));
    outputs(5632) <= layer4_outputs(5487);
    outputs(5633) <= not((layer4_outputs(5953)) xor (layer4_outputs(1307)));
    outputs(5634) <= not(layer4_outputs(225));
    outputs(5635) <= layer4_outputs(3885);
    outputs(5636) <= not(layer4_outputs(2564));
    outputs(5637) <= not(layer4_outputs(3641));
    outputs(5638) <= (layer4_outputs(4389)) xor (layer4_outputs(4527));
    outputs(5639) <= layer4_outputs(8258);
    outputs(5640) <= (layer4_outputs(2515)) xor (layer4_outputs(8405));
    outputs(5641) <= not(layer4_outputs(4619)) or (layer4_outputs(3277));
    outputs(5642) <= layer4_outputs(7688);
    outputs(5643) <= (layer4_outputs(9769)) xor (layer4_outputs(2106));
    outputs(5644) <= (layer4_outputs(3176)) or (layer4_outputs(991));
    outputs(5645) <= not((layer4_outputs(9887)) xor (layer4_outputs(393)));
    outputs(5646) <= layer4_outputs(1236);
    outputs(5647) <= not(layer4_outputs(6110));
    outputs(5648) <= not((layer4_outputs(9641)) xor (layer4_outputs(9605)));
    outputs(5649) <= (layer4_outputs(7085)) or (layer4_outputs(728));
    outputs(5650) <= not(layer4_outputs(1361)) or (layer4_outputs(1334));
    outputs(5651) <= layer4_outputs(8664);
    outputs(5652) <= layer4_outputs(74);
    outputs(5653) <= not((layer4_outputs(4519)) and (layer4_outputs(9119)));
    outputs(5654) <= not(layer4_outputs(6177));
    outputs(5655) <= (layer4_outputs(8254)) and not (layer4_outputs(6716));
    outputs(5656) <= not(layer4_outputs(5210));
    outputs(5657) <= (layer4_outputs(4500)) xor (layer4_outputs(9774));
    outputs(5658) <= not(layer4_outputs(1462)) or (layer4_outputs(5562));
    outputs(5659) <= layer4_outputs(6659);
    outputs(5660) <= layer4_outputs(8616);
    outputs(5661) <= (layer4_outputs(3244)) xor (layer4_outputs(9898));
    outputs(5662) <= not((layer4_outputs(2832)) xor (layer4_outputs(5135)));
    outputs(5663) <= not(layer4_outputs(8713));
    outputs(5664) <= not(layer4_outputs(5049));
    outputs(5665) <= (layer4_outputs(9118)) and not (layer4_outputs(4784));
    outputs(5666) <= not(layer4_outputs(3952));
    outputs(5667) <= (layer4_outputs(6505)) xor (layer4_outputs(6259));
    outputs(5668) <= not(layer4_outputs(3719));
    outputs(5669) <= (layer4_outputs(8539)) or (layer4_outputs(6658));
    outputs(5670) <= layer4_outputs(2233);
    outputs(5671) <= not(layer4_outputs(4985)) or (layer4_outputs(5634));
    outputs(5672) <= layer4_outputs(3049);
    outputs(5673) <= not(layer4_outputs(2679));
    outputs(5674) <= not(layer4_outputs(1680));
    outputs(5675) <= not(layer4_outputs(4966));
    outputs(5676) <= not(layer4_outputs(4103));
    outputs(5677) <= layer4_outputs(864);
    outputs(5678) <= not(layer4_outputs(4976));
    outputs(5679) <= (layer4_outputs(1519)) and not (layer4_outputs(745));
    outputs(5680) <= not(layer4_outputs(1638)) or (layer4_outputs(8864));
    outputs(5681) <= not(layer4_outputs(732));
    outputs(5682) <= layer4_outputs(7113);
    outputs(5683) <= not(layer4_outputs(6727));
    outputs(5684) <= layer4_outputs(6560);
    outputs(5685) <= layer4_outputs(9490);
    outputs(5686) <= not((layer4_outputs(5365)) and (layer4_outputs(8071)));
    outputs(5687) <= not((layer4_outputs(5296)) xor (layer4_outputs(9477)));
    outputs(5688) <= not((layer4_outputs(9959)) xor (layer4_outputs(5785)));
    outputs(5689) <= not(layer4_outputs(4185));
    outputs(5690) <= layer4_outputs(4252);
    outputs(5691) <= not(layer4_outputs(4557));
    outputs(5692) <= layer4_outputs(9110);
    outputs(5693) <= layer4_outputs(10121);
    outputs(5694) <= not(layer4_outputs(3994));
    outputs(5695) <= layer4_outputs(8710);
    outputs(5696) <= layer4_outputs(818);
    outputs(5697) <= not(layer4_outputs(1938));
    outputs(5698) <= layer4_outputs(5236);
    outputs(5699) <= (layer4_outputs(9458)) xor (layer4_outputs(8677));
    outputs(5700) <= (layer4_outputs(2897)) xor (layer4_outputs(5169));
    outputs(5701) <= layer4_outputs(1718);
    outputs(5702) <= layer4_outputs(3552);
    outputs(5703) <= not((layer4_outputs(4745)) xor (layer4_outputs(9609)));
    outputs(5704) <= (layer4_outputs(21)) or (layer4_outputs(8365));
    outputs(5705) <= layer4_outputs(4818);
    outputs(5706) <= (layer4_outputs(4833)) xor (layer4_outputs(6356));
    outputs(5707) <= layer4_outputs(7445);
    outputs(5708) <= layer4_outputs(6305);
    outputs(5709) <= not(layer4_outputs(5113));
    outputs(5710) <= not((layer4_outputs(6548)) xor (layer4_outputs(556)));
    outputs(5711) <= not(layer4_outputs(8657)) or (layer4_outputs(3356));
    outputs(5712) <= (layer4_outputs(5768)) xor (layer4_outputs(2481));
    outputs(5713) <= (layer4_outputs(874)) xor (layer4_outputs(8076));
    outputs(5714) <= not(layer4_outputs(7275));
    outputs(5715) <= (layer4_outputs(2244)) or (layer4_outputs(5827));
    outputs(5716) <= (layer4_outputs(6579)) xor (layer4_outputs(3786));
    outputs(5717) <= not(layer4_outputs(8023));
    outputs(5718) <= not(layer4_outputs(808));
    outputs(5719) <= not((layer4_outputs(5764)) xor (layer4_outputs(5212)));
    outputs(5720) <= not(layer4_outputs(5551));
    outputs(5721) <= layer4_outputs(3657);
    outputs(5722) <= (layer4_outputs(6936)) xor (layer4_outputs(3664));
    outputs(5723) <= layer4_outputs(8608);
    outputs(5724) <= (layer4_outputs(6830)) xor (layer4_outputs(5690));
    outputs(5725) <= layer4_outputs(3764);
    outputs(5726) <= not(layer4_outputs(10061));
    outputs(5727) <= not((layer4_outputs(9881)) xor (layer4_outputs(1534)));
    outputs(5728) <= not((layer4_outputs(9640)) and (layer4_outputs(3531)));
    outputs(5729) <= (layer4_outputs(7416)) xor (layer4_outputs(2463));
    outputs(5730) <= not(layer4_outputs(6507));
    outputs(5731) <= not(layer4_outputs(9555));
    outputs(5732) <= layer4_outputs(9629);
    outputs(5733) <= not(layer4_outputs(9003));
    outputs(5734) <= layer4_outputs(3966);
    outputs(5735) <= layer4_outputs(1591);
    outputs(5736) <= not(layer4_outputs(505));
    outputs(5737) <= (layer4_outputs(6609)) xor (layer4_outputs(8851));
    outputs(5738) <= not(layer4_outputs(6004));
    outputs(5739) <= layer4_outputs(9160);
    outputs(5740) <= (layer4_outputs(2146)) xor (layer4_outputs(8885));
    outputs(5741) <= layer4_outputs(4188);
    outputs(5742) <= layer4_outputs(7875);
    outputs(5743) <= (layer4_outputs(919)) xor (layer4_outputs(5193));
    outputs(5744) <= not(layer4_outputs(3433));
    outputs(5745) <= not(layer4_outputs(3447));
    outputs(5746) <= layer4_outputs(8219);
    outputs(5747) <= layer4_outputs(1618);
    outputs(5748) <= not(layer4_outputs(2762));
    outputs(5749) <= layer4_outputs(2642);
    outputs(5750) <= not(layer4_outputs(635));
    outputs(5751) <= not(layer4_outputs(4466));
    outputs(5752) <= (layer4_outputs(1756)) and (layer4_outputs(6091));
    outputs(5753) <= (layer4_outputs(2610)) xor (layer4_outputs(1121));
    outputs(5754) <= layer4_outputs(8547);
    outputs(5755) <= not((layer4_outputs(1151)) xor (layer4_outputs(1780)));
    outputs(5756) <= not((layer4_outputs(5632)) xor (layer4_outputs(5535)));
    outputs(5757) <= not((layer4_outputs(9732)) and (layer4_outputs(9863)));
    outputs(5758) <= layer4_outputs(243);
    outputs(5759) <= layer4_outputs(6228);
    outputs(5760) <= not(layer4_outputs(6372));
    outputs(5761) <= (layer4_outputs(7749)) xor (layer4_outputs(172));
    outputs(5762) <= (layer4_outputs(2902)) or (layer4_outputs(67));
    outputs(5763) <= (layer4_outputs(1254)) xor (layer4_outputs(3874));
    outputs(5764) <= not((layer4_outputs(5594)) xor (layer4_outputs(1660)));
    outputs(5765) <= not(layer4_outputs(1917));
    outputs(5766) <= layer4_outputs(9004);
    outputs(5767) <= not((layer4_outputs(1863)) xor (layer4_outputs(4267)));
    outputs(5768) <= layer4_outputs(2840);
    outputs(5769) <= layer4_outputs(2958);
    outputs(5770) <= layer4_outputs(9372);
    outputs(5771) <= not((layer4_outputs(8212)) and (layer4_outputs(1027)));
    outputs(5772) <= layer4_outputs(8982);
    outputs(5773) <= (layer4_outputs(9914)) xor (layer4_outputs(9435));
    outputs(5774) <= (layer4_outputs(5527)) xor (layer4_outputs(1161));
    outputs(5775) <= not(layer4_outputs(7453));
    outputs(5776) <= (layer4_outputs(9004)) xor (layer4_outputs(3019));
    outputs(5777) <= not(layer4_outputs(2604));
    outputs(5778) <= not(layer4_outputs(6155)) or (layer4_outputs(5170));
    outputs(5779) <= not(layer4_outputs(3520));
    outputs(5780) <= layer4_outputs(7758);
    outputs(5781) <= layer4_outputs(6351);
    outputs(5782) <= (layer4_outputs(84)) xor (layer4_outputs(3391));
    outputs(5783) <= (layer4_outputs(7654)) xor (layer4_outputs(1265));
    outputs(5784) <= not((layer4_outputs(2149)) xor (layer4_outputs(1770)));
    outputs(5785) <= not(layer4_outputs(6507));
    outputs(5786) <= layer4_outputs(3420);
    outputs(5787) <= not((layer4_outputs(8158)) and (layer4_outputs(9317)));
    outputs(5788) <= layer4_outputs(453);
    outputs(5789) <= not((layer4_outputs(413)) xor (layer4_outputs(3369)));
    outputs(5790) <= (layer4_outputs(2764)) and not (layer4_outputs(2122));
    outputs(5791) <= not(layer4_outputs(7998));
    outputs(5792) <= (layer4_outputs(1003)) xor (layer4_outputs(5925));
    outputs(5793) <= layer4_outputs(5457);
    outputs(5794) <= layer4_outputs(2730);
    outputs(5795) <= not(layer4_outputs(10212));
    outputs(5796) <= layer4_outputs(2772);
    outputs(5797) <= layer4_outputs(9726);
    outputs(5798) <= not(layer4_outputs(3089));
    outputs(5799) <= (layer4_outputs(4294)) and not (layer4_outputs(3036));
    outputs(5800) <= (layer4_outputs(1908)) and not (layer4_outputs(1));
    outputs(5801) <= (layer4_outputs(5524)) xor (layer4_outputs(4848));
    outputs(5802) <= layer4_outputs(7699);
    outputs(5803) <= not((layer4_outputs(7188)) xor (layer4_outputs(5016)));
    outputs(5804) <= not((layer4_outputs(6790)) xor (layer4_outputs(6619)));
    outputs(5805) <= layer4_outputs(8325);
    outputs(5806) <= layer4_outputs(6290);
    outputs(5807) <= layer4_outputs(5332);
    outputs(5808) <= not(layer4_outputs(2078));
    outputs(5809) <= layer4_outputs(743);
    outputs(5810) <= not(layer4_outputs(1522));
    outputs(5811) <= layer4_outputs(9756);
    outputs(5812) <= not(layer4_outputs(8025));
    outputs(5813) <= not((layer4_outputs(5978)) xor (layer4_outputs(6064)));
    outputs(5814) <= layer4_outputs(5473);
    outputs(5815) <= not((layer4_outputs(2175)) xor (layer4_outputs(2527)));
    outputs(5816) <= not((layer4_outputs(9528)) xor (layer4_outputs(10153)));
    outputs(5817) <= not(layer4_outputs(1657));
    outputs(5818) <= not(layer4_outputs(1782));
    outputs(5819) <= not(layer4_outputs(9843)) or (layer4_outputs(5213));
    outputs(5820) <= not((layer4_outputs(477)) and (layer4_outputs(7082)));
    outputs(5821) <= not((layer4_outputs(7845)) xor (layer4_outputs(6458)));
    outputs(5822) <= layer4_outputs(831);
    outputs(5823) <= (layer4_outputs(2510)) xor (layer4_outputs(2553));
    outputs(5824) <= layer4_outputs(6233);
    outputs(5825) <= (layer4_outputs(8251)) xor (layer4_outputs(3613));
    outputs(5826) <= layer4_outputs(9239);
    outputs(5827) <= not(layer4_outputs(586));
    outputs(5828) <= (layer4_outputs(1552)) or (layer4_outputs(8059));
    outputs(5829) <= (layer4_outputs(831)) and not (layer4_outputs(5477));
    outputs(5830) <= not(layer4_outputs(5868));
    outputs(5831) <= not((layer4_outputs(8149)) xor (layer4_outputs(2271)));
    outputs(5832) <= not(layer4_outputs(9570));
    outputs(5833) <= (layer4_outputs(6998)) xor (layer4_outputs(5350));
    outputs(5834) <= not(layer4_outputs(1324));
    outputs(5835) <= not(layer4_outputs(2552));
    outputs(5836) <= not(layer4_outputs(5334));
    outputs(5837) <= (layer4_outputs(9549)) xor (layer4_outputs(9904));
    outputs(5838) <= layer4_outputs(6954);
    outputs(5839) <= not(layer4_outputs(7323));
    outputs(5840) <= not(layer4_outputs(4297));
    outputs(5841) <= not(layer4_outputs(9048));
    outputs(5842) <= layer4_outputs(10100);
    outputs(5843) <= layer4_outputs(4957);
    outputs(5844) <= (layer4_outputs(7105)) and (layer4_outputs(9836));
    outputs(5845) <= not((layer4_outputs(4330)) xor (layer4_outputs(3132)));
    outputs(5846) <= not(layer4_outputs(6870));
    outputs(5847) <= not((layer4_outputs(9472)) xor (layer4_outputs(6786)));
    outputs(5848) <= not(layer4_outputs(1850));
    outputs(5849) <= not((layer4_outputs(5273)) xor (layer4_outputs(4583)));
    outputs(5850) <= (layer4_outputs(8671)) or (layer4_outputs(1033));
    outputs(5851) <= (layer4_outputs(5638)) xor (layer4_outputs(7928));
    outputs(5852) <= layer4_outputs(7051);
    outputs(5853) <= not(layer4_outputs(3859));
    outputs(5854) <= layer4_outputs(7084);
    outputs(5855) <= not(layer4_outputs(7907));
    outputs(5856) <= layer4_outputs(9618);
    outputs(5857) <= (layer4_outputs(5045)) and not (layer4_outputs(2832));
    outputs(5858) <= (layer4_outputs(1078)) and (layer4_outputs(5661));
    outputs(5859) <= not(layer4_outputs(7578));
    outputs(5860) <= layer4_outputs(7268);
    outputs(5861) <= not(layer4_outputs(9523));
    outputs(5862) <= '1';
    outputs(5863) <= not(layer4_outputs(196));
    outputs(5864) <= layer4_outputs(6275);
    outputs(5865) <= not(layer4_outputs(5404));
    outputs(5866) <= not((layer4_outputs(2683)) xor (layer4_outputs(7627)));
    outputs(5867) <= layer4_outputs(6709);
    outputs(5868) <= not((layer4_outputs(9419)) xor (layer4_outputs(5434)));
    outputs(5869) <= (layer4_outputs(781)) xor (layer4_outputs(2783));
    outputs(5870) <= not(layer4_outputs(1757));
    outputs(5871) <= layer4_outputs(7542);
    outputs(5872) <= layer4_outputs(425);
    outputs(5873) <= layer4_outputs(7125);
    outputs(5874) <= not(layer4_outputs(1506));
    outputs(5875) <= not(layer4_outputs(3334));
    outputs(5876) <= not((layer4_outputs(6057)) xor (layer4_outputs(6125)));
    outputs(5877) <= (layer4_outputs(1014)) xor (layer4_outputs(9024));
    outputs(5878) <= (layer4_outputs(9100)) xor (layer4_outputs(7953));
    outputs(5879) <= not((layer4_outputs(9530)) and (layer4_outputs(7960)));
    outputs(5880) <= not(layer4_outputs(8681));
    outputs(5881) <= (layer4_outputs(9394)) and not (layer4_outputs(4906));
    outputs(5882) <= (layer4_outputs(9992)) or (layer4_outputs(2184));
    outputs(5883) <= layer4_outputs(759);
    outputs(5884) <= not((layer4_outputs(454)) xor (layer4_outputs(7490)));
    outputs(5885) <= layer4_outputs(7802);
    outputs(5886) <= not(layer4_outputs(5250));
    outputs(5887) <= not((layer4_outputs(9414)) and (layer4_outputs(313)));
    outputs(5888) <= (layer4_outputs(7463)) xor (layer4_outputs(204));
    outputs(5889) <= not(layer4_outputs(1542)) or (layer4_outputs(7464));
    outputs(5890) <= (layer4_outputs(6223)) or (layer4_outputs(6629));
    outputs(5891) <= not(layer4_outputs(4715));
    outputs(5892) <= not(layer4_outputs(5465));
    outputs(5893) <= layer4_outputs(9504);
    outputs(5894) <= not(layer4_outputs(7565));
    outputs(5895) <= not((layer4_outputs(9799)) xor (layer4_outputs(107)));
    outputs(5896) <= (layer4_outputs(2909)) or (layer4_outputs(5337));
    outputs(5897) <= layer4_outputs(7375);
    outputs(5898) <= layer4_outputs(9954);
    outputs(5899) <= layer4_outputs(5040);
    outputs(5900) <= (layer4_outputs(3456)) xor (layer4_outputs(7114));
    outputs(5901) <= not(layer4_outputs(722));
    outputs(5902) <= not(layer4_outputs(8644)) or (layer4_outputs(4492));
    outputs(5903) <= (layer4_outputs(6295)) xor (layer4_outputs(5375));
    outputs(5904) <= not(layer4_outputs(8292));
    outputs(5905) <= layer4_outputs(9020);
    outputs(5906) <= not(layer4_outputs(33));
    outputs(5907) <= layer4_outputs(6522);
    outputs(5908) <= (layer4_outputs(1799)) or (layer4_outputs(4339));
    outputs(5909) <= not(layer4_outputs(6864));
    outputs(5910) <= not((layer4_outputs(5414)) xor (layer4_outputs(4186)));
    outputs(5911) <= (layer4_outputs(8460)) and not (layer4_outputs(5310));
    outputs(5912) <= layer4_outputs(5141);
    outputs(5913) <= layer4_outputs(7633);
    outputs(5914) <= (layer4_outputs(6277)) and not (layer4_outputs(8782));
    outputs(5915) <= not(layer4_outputs(4851));
    outputs(5916) <= layer4_outputs(9580);
    outputs(5917) <= layer4_outputs(6883);
    outputs(5918) <= not((layer4_outputs(9663)) and (layer4_outputs(5757)));
    outputs(5919) <= layer4_outputs(187);
    outputs(5920) <= (layer4_outputs(2492)) or (layer4_outputs(7317));
    outputs(5921) <= layer4_outputs(1298);
    outputs(5922) <= (layer4_outputs(8724)) xor (layer4_outputs(484));
    outputs(5923) <= not((layer4_outputs(7084)) xor (layer4_outputs(2797)));
    outputs(5924) <= layer4_outputs(8676);
    outputs(5925) <= not(layer4_outputs(887));
    outputs(5926) <= not(layer4_outputs(9848));
    outputs(5927) <= (layer4_outputs(5970)) xor (layer4_outputs(4151));
    outputs(5928) <= not((layer4_outputs(1418)) or (layer4_outputs(1123)));
    outputs(5929) <= layer4_outputs(3073);
    outputs(5930) <= (layer4_outputs(449)) xor (layer4_outputs(7100));
    outputs(5931) <= layer4_outputs(4310);
    outputs(5932) <= not(layer4_outputs(9707));
    outputs(5933) <= not(layer4_outputs(1688));
    outputs(5934) <= (layer4_outputs(5997)) xor (layer4_outputs(803));
    outputs(5935) <= not((layer4_outputs(5321)) and (layer4_outputs(2525)));
    outputs(5936) <= not(layer4_outputs(7314));
    outputs(5937) <= not(layer4_outputs(5936)) or (layer4_outputs(3443));
    outputs(5938) <= (layer4_outputs(6857)) xor (layer4_outputs(3582));
    outputs(5939) <= not(layer4_outputs(6385));
    outputs(5940) <= not(layer4_outputs(9343));
    outputs(5941) <= layer4_outputs(622);
    outputs(5942) <= not(layer4_outputs(3585));
    outputs(5943) <= layer4_outputs(2753);
    outputs(5944) <= layer4_outputs(193);
    outputs(5945) <= (layer4_outputs(9123)) xor (layer4_outputs(3326));
    outputs(5946) <= not(layer4_outputs(7614));
    outputs(5947) <= not(layer4_outputs(4440));
    outputs(5948) <= not((layer4_outputs(5119)) xor (layer4_outputs(2148)));
    outputs(5949) <= not((layer4_outputs(1645)) and (layer4_outputs(7656)));
    outputs(5950) <= not(layer4_outputs(4844)) or (layer4_outputs(954));
    outputs(5951) <= not(layer4_outputs(1928));
    outputs(5952) <= not(layer4_outputs(2679));
    outputs(5953) <= not((layer4_outputs(63)) xor (layer4_outputs(1717)));
    outputs(5954) <= (layer4_outputs(7109)) xor (layer4_outputs(3284));
    outputs(5955) <= layer4_outputs(7961);
    outputs(5956) <= not((layer4_outputs(4999)) and (layer4_outputs(7033)));
    outputs(5957) <= not((layer4_outputs(439)) xor (layer4_outputs(8575)));
    outputs(5958) <= not((layer4_outputs(3391)) xor (layer4_outputs(5159)));
    outputs(5959) <= (layer4_outputs(2209)) xor (layer4_outputs(4079));
    outputs(5960) <= layer4_outputs(8645);
    outputs(5961) <= not((layer4_outputs(2427)) xor (layer4_outputs(1260)));
    outputs(5962) <= (layer4_outputs(4239)) or (layer4_outputs(1041));
    outputs(5963) <= not(layer4_outputs(4528));
    outputs(5964) <= layer4_outputs(6320);
    outputs(5965) <= not(layer4_outputs(8708));
    outputs(5966) <= (layer4_outputs(8918)) xor (layer4_outputs(3225));
    outputs(5967) <= not(layer4_outputs(9450));
    outputs(5968) <= (layer4_outputs(4491)) xor (layer4_outputs(1302));
    outputs(5969) <= layer4_outputs(8579);
    outputs(5970) <= layer4_outputs(1869);
    outputs(5971) <= not(layer4_outputs(4335)) or (layer4_outputs(1061));
    outputs(5972) <= (layer4_outputs(9039)) xor (layer4_outputs(1852));
    outputs(5973) <= (layer4_outputs(7952)) xor (layer4_outputs(2522));
    outputs(5974) <= (layer4_outputs(9211)) xor (layer4_outputs(9289));
    outputs(5975) <= (layer4_outputs(7434)) xor (layer4_outputs(6860));
    outputs(5976) <= layer4_outputs(7238);
    outputs(5977) <= not((layer4_outputs(3290)) xor (layer4_outputs(4896)));
    outputs(5978) <= not((layer4_outputs(2460)) xor (layer4_outputs(8719)));
    outputs(5979) <= layer4_outputs(7815);
    outputs(5980) <= (layer4_outputs(1499)) or (layer4_outputs(646));
    outputs(5981) <= layer4_outputs(6121);
    outputs(5982) <= not(layer4_outputs(8123));
    outputs(5983) <= (layer4_outputs(781)) and (layer4_outputs(125));
    outputs(5984) <= layer4_outputs(845);
    outputs(5985) <= layer4_outputs(4303);
    outputs(5986) <= not((layer4_outputs(6982)) xor (layer4_outputs(4209)));
    outputs(5987) <= (layer4_outputs(448)) xor (layer4_outputs(9804));
    outputs(5988) <= not(layer4_outputs(1689));
    outputs(5989) <= (layer4_outputs(6411)) xor (layer4_outputs(3584));
    outputs(5990) <= not(layer4_outputs(4003)) or (layer4_outputs(3944));
    outputs(5991) <= not((layer4_outputs(8483)) xor (layer4_outputs(7000)));
    outputs(5992) <= layer4_outputs(2229);
    outputs(5993) <= not(layer4_outputs(5074));
    outputs(5994) <= (layer4_outputs(2877)) xor (layer4_outputs(6596));
    outputs(5995) <= (layer4_outputs(6168)) xor (layer4_outputs(5812));
    outputs(5996) <= not(layer4_outputs(262)) or (layer4_outputs(1273));
    outputs(5997) <= not((layer4_outputs(2022)) xor (layer4_outputs(1189)));
    outputs(5998) <= not((layer4_outputs(4438)) xor (layer4_outputs(6802)));
    outputs(5999) <= not(layer4_outputs(1487));
    outputs(6000) <= not(layer4_outputs(4306));
    outputs(6001) <= not(layer4_outputs(9126));
    outputs(6002) <= not((layer4_outputs(5881)) xor (layer4_outputs(1650)));
    outputs(6003) <= layer4_outputs(3252);
    outputs(6004) <= (layer4_outputs(6798)) and (layer4_outputs(6666));
    outputs(6005) <= not(layer4_outputs(941));
    outputs(6006) <= (layer4_outputs(3285)) xor (layer4_outputs(2050));
    outputs(6007) <= not((layer4_outputs(9477)) xor (layer4_outputs(5749)));
    outputs(6008) <= not(layer4_outputs(2655));
    outputs(6009) <= not(layer4_outputs(575));
    outputs(6010) <= not(layer4_outputs(1893));
    outputs(6011) <= layer4_outputs(9408);
    outputs(6012) <= layer4_outputs(6393);
    outputs(6013) <= not(layer4_outputs(2463));
    outputs(6014) <= layer4_outputs(8665);
    outputs(6015) <= not((layer4_outputs(2256)) and (layer4_outputs(5003)));
    outputs(6016) <= not(layer4_outputs(9191));
    outputs(6017) <= not((layer4_outputs(6431)) xor (layer4_outputs(6251)));
    outputs(6018) <= layer4_outputs(9221);
    outputs(6019) <= '1';
    outputs(6020) <= not(layer4_outputs(2216));
    outputs(6021) <= not(layer4_outputs(8392));
    outputs(6022) <= (layer4_outputs(2700)) xor (layer4_outputs(6231));
    outputs(6023) <= (layer4_outputs(6993)) xor (layer4_outputs(7299));
    outputs(6024) <= (layer4_outputs(8196)) xor (layer4_outputs(8074));
    outputs(6025) <= not(layer4_outputs(7714));
    outputs(6026) <= not((layer4_outputs(5542)) xor (layer4_outputs(8459)));
    outputs(6027) <= (layer4_outputs(2190)) xor (layer4_outputs(7312));
    outputs(6028) <= (layer4_outputs(2423)) xor (layer4_outputs(8999));
    outputs(6029) <= (layer4_outputs(9913)) and (layer4_outputs(1045));
    outputs(6030) <= layer4_outputs(58);
    outputs(6031) <= not((layer4_outputs(202)) xor (layer4_outputs(9715)));
    outputs(6032) <= not(layer4_outputs(3096));
    outputs(6033) <= not(layer4_outputs(2913));
    outputs(6034) <= layer4_outputs(2840);
    outputs(6035) <= layer4_outputs(7474);
    outputs(6036) <= (layer4_outputs(3660)) xor (layer4_outputs(2950));
    outputs(6037) <= layer4_outputs(4684);
    outputs(6038) <= (layer4_outputs(6455)) and not (layer4_outputs(9918));
    outputs(6039) <= not((layer4_outputs(6337)) xor (layer4_outputs(4069)));
    outputs(6040) <= layer4_outputs(10029);
    outputs(6041) <= not(layer4_outputs(8497));
    outputs(6042) <= layer4_outputs(5383);
    outputs(6043) <= (layer4_outputs(4121)) xor (layer4_outputs(3842));
    outputs(6044) <= not((layer4_outputs(8723)) xor (layer4_outputs(6036)));
    outputs(6045) <= (layer4_outputs(6396)) xor (layer4_outputs(4781));
    outputs(6046) <= not(layer4_outputs(6692));
    outputs(6047) <= not((layer4_outputs(7048)) xor (layer4_outputs(5166)));
    outputs(6048) <= layer4_outputs(2067);
    outputs(6049) <= not((layer4_outputs(2166)) or (layer4_outputs(6521)));
    outputs(6050) <= layer4_outputs(2592);
    outputs(6051) <= (layer4_outputs(2696)) or (layer4_outputs(6950));
    outputs(6052) <= not(layer4_outputs(6380));
    outputs(6053) <= not((layer4_outputs(1804)) and (layer4_outputs(274)));
    outputs(6054) <= not(layer4_outputs(3637)) or (layer4_outputs(4087));
    outputs(6055) <= not(layer4_outputs(8521));
    outputs(6056) <= layer4_outputs(9221);
    outputs(6057) <= not(layer4_outputs(1256)) or (layer4_outputs(9758));
    outputs(6058) <= layer4_outputs(227);
    outputs(6059) <= not((layer4_outputs(7923)) or (layer4_outputs(6301)));
    outputs(6060) <= not(layer4_outputs(3929)) or (layer4_outputs(7957));
    outputs(6061) <= not((layer4_outputs(6262)) xor (layer4_outputs(8546)));
    outputs(6062) <= not(layer4_outputs(4205));
    outputs(6063) <= not(layer4_outputs(1007));
    outputs(6064) <= not((layer4_outputs(224)) xor (layer4_outputs(6100)));
    outputs(6065) <= not((layer4_outputs(8288)) xor (layer4_outputs(1084)));
    outputs(6066) <= (layer4_outputs(5376)) xor (layer4_outputs(4114));
    outputs(6067) <= not((layer4_outputs(7937)) xor (layer4_outputs(3284)));
    outputs(6068) <= not((layer4_outputs(8612)) or (layer4_outputs(9782)));
    outputs(6069) <= layer4_outputs(8012);
    outputs(6070) <= not(layer4_outputs(4759));
    outputs(6071) <= not((layer4_outputs(7536)) xor (layer4_outputs(5806)));
    outputs(6072) <= (layer4_outputs(2704)) xor (layer4_outputs(8466));
    outputs(6073) <= not(layer4_outputs(3526));
    outputs(6074) <= '1';
    outputs(6075) <= (layer4_outputs(8528)) and not (layer4_outputs(7278));
    outputs(6076) <= layer4_outputs(668);
    outputs(6077) <= not((layer4_outputs(5845)) xor (layer4_outputs(3651)));
    outputs(6078) <= (layer4_outputs(5921)) xor (layer4_outputs(5162));
    outputs(6079) <= not(layer4_outputs(9107));
    outputs(6080) <= not(layer4_outputs(3851)) or (layer4_outputs(1774));
    outputs(6081) <= (layer4_outputs(7417)) xor (layer4_outputs(9800));
    outputs(6082) <= (layer4_outputs(5298)) xor (layer4_outputs(381));
    outputs(6083) <= not((layer4_outputs(6193)) and (layer4_outputs(1680)));
    outputs(6084) <= not((layer4_outputs(8870)) xor (layer4_outputs(1656)));
    outputs(6085) <= not(layer4_outputs(9165));
    outputs(6086) <= not(layer4_outputs(6386));
    outputs(6087) <= (layer4_outputs(3)) and not (layer4_outputs(2145));
    outputs(6088) <= layer4_outputs(4111);
    outputs(6089) <= (layer4_outputs(7058)) or (layer4_outputs(2904));
    outputs(6090) <= (layer4_outputs(6414)) and (layer4_outputs(5418));
    outputs(6091) <= (layer4_outputs(9173)) xor (layer4_outputs(4724));
    outputs(6092) <= not((layer4_outputs(3092)) and (layer4_outputs(1218)));
    outputs(6093) <= not(layer4_outputs(8812));
    outputs(6094) <= (layer4_outputs(8255)) xor (layer4_outputs(4456));
    outputs(6095) <= not((layer4_outputs(3294)) xor (layer4_outputs(2899)));
    outputs(6096) <= not((layer4_outputs(8170)) or (layer4_outputs(5022)));
    outputs(6097) <= not((layer4_outputs(8895)) xor (layer4_outputs(8021)));
    outputs(6098) <= not(layer4_outputs(4032));
    outputs(6099) <= not((layer4_outputs(7110)) xor (layer4_outputs(2377)));
    outputs(6100) <= not(layer4_outputs(3495));
    outputs(6101) <= (layer4_outputs(5421)) and (layer4_outputs(4432));
    outputs(6102) <= not(layer4_outputs(5686));
    outputs(6103) <= not(layer4_outputs(2733));
    outputs(6104) <= not(layer4_outputs(430));
    outputs(6105) <= layer4_outputs(1198);
    outputs(6106) <= layer4_outputs(1626);
    outputs(6107) <= layer4_outputs(7424);
    outputs(6108) <= not(layer4_outputs(135)) or (layer4_outputs(949));
    outputs(6109) <= not(layer4_outputs(9312));
    outputs(6110) <= not((layer4_outputs(7573)) and (layer4_outputs(458)));
    outputs(6111) <= (layer4_outputs(1790)) xor (layer4_outputs(2171));
    outputs(6112) <= (layer4_outputs(3951)) and not (layer4_outputs(9087));
    outputs(6113) <= layer4_outputs(2054);
    outputs(6114) <= not((layer4_outputs(7954)) or (layer4_outputs(1282)));
    outputs(6115) <= not((layer4_outputs(7517)) xor (layer4_outputs(9291)));
    outputs(6116) <= layer4_outputs(3088);
    outputs(6117) <= (layer4_outputs(7143)) xor (layer4_outputs(3111));
    outputs(6118) <= (layer4_outputs(8343)) xor (layer4_outputs(8492));
    outputs(6119) <= not((layer4_outputs(5115)) xor (layer4_outputs(1425)));
    outputs(6120) <= layer4_outputs(7615);
    outputs(6121) <= not(layer4_outputs(4687)) or (layer4_outputs(2579));
    outputs(6122) <= (layer4_outputs(4899)) xor (layer4_outputs(1696));
    outputs(6123) <= not((layer4_outputs(8091)) or (layer4_outputs(2170)));
    outputs(6124) <= not((layer4_outputs(1612)) xor (layer4_outputs(4096)));
    outputs(6125) <= layer4_outputs(3055);
    outputs(6126) <= layer4_outputs(6757);
    outputs(6127) <= not(layer4_outputs(8724)) or (layer4_outputs(5976));
    outputs(6128) <= (layer4_outputs(9163)) xor (layer4_outputs(2629));
    outputs(6129) <= not(layer4_outputs(8216));
    outputs(6130) <= not(layer4_outputs(8168));
    outputs(6131) <= not(layer4_outputs(4040));
    outputs(6132) <= (layer4_outputs(5848)) xor (layer4_outputs(6902));
    outputs(6133) <= (layer4_outputs(4641)) xor (layer4_outputs(4891));
    outputs(6134) <= not(layer4_outputs(324));
    outputs(6135) <= not(layer4_outputs(5649));
    outputs(6136) <= (layer4_outputs(9341)) xor (layer4_outputs(7151));
    outputs(6137) <= (layer4_outputs(5489)) xor (layer4_outputs(6526));
    outputs(6138) <= layer4_outputs(445);
    outputs(6139) <= not(layer4_outputs(3787));
    outputs(6140) <= not(layer4_outputs(833));
    outputs(6141) <= layer4_outputs(6581);
    outputs(6142) <= not(layer4_outputs(252));
    outputs(6143) <= not(layer4_outputs(1822));
    outputs(6144) <= not(layer4_outputs(8107));
    outputs(6145) <= (layer4_outputs(1426)) and not (layer4_outputs(3115));
    outputs(6146) <= not((layer4_outputs(6447)) xor (layer4_outputs(9635)));
    outputs(6147) <= (layer4_outputs(3234)) or (layer4_outputs(6332));
    outputs(6148) <= layer4_outputs(3886);
    outputs(6149) <= not(layer4_outputs(6805));
    outputs(6150) <= layer4_outputs(3571);
    outputs(6151) <= not(layer4_outputs(9271)) or (layer4_outputs(9519));
    outputs(6152) <= not((layer4_outputs(928)) or (layer4_outputs(9781)));
    outputs(6153) <= layer4_outputs(5872);
    outputs(6154) <= (layer4_outputs(10126)) and not (layer4_outputs(9628));
    outputs(6155) <= not(layer4_outputs(2211));
    outputs(6156) <= (layer4_outputs(9524)) and (layer4_outputs(3167));
    outputs(6157) <= not(layer4_outputs(3097));
    outputs(6158) <= layer4_outputs(4282);
    outputs(6159) <= not(layer4_outputs(6006));
    outputs(6160) <= layer4_outputs(5467);
    outputs(6161) <= layer4_outputs(7447);
    outputs(6162) <= not(layer4_outputs(8138)) or (layer4_outputs(4821));
    outputs(6163) <= not(layer4_outputs(5184));
    outputs(6164) <= not((layer4_outputs(6531)) xor (layer4_outputs(1608)));
    outputs(6165) <= not(layer4_outputs(4951));
    outputs(6166) <= (layer4_outputs(8204)) xor (layer4_outputs(8173));
    outputs(6167) <= (layer4_outputs(3228)) or (layer4_outputs(2946));
    outputs(6168) <= layer4_outputs(2766);
    outputs(6169) <= layer4_outputs(2089);
    outputs(6170) <= layer4_outputs(6748);
    outputs(6171) <= not((layer4_outputs(350)) xor (layer4_outputs(10084)));
    outputs(6172) <= not((layer4_outputs(5351)) and (layer4_outputs(10192)));
    outputs(6173) <= (layer4_outputs(9001)) xor (layer4_outputs(8560));
    outputs(6174) <= layer4_outputs(7379);
    outputs(6175) <= layer4_outputs(1660);
    outputs(6176) <= layer4_outputs(6859);
    outputs(6177) <= layer4_outputs(3812);
    outputs(6178) <= layer4_outputs(5560);
    outputs(6179) <= not(layer4_outputs(1670));
    outputs(6180) <= (layer4_outputs(1288)) xor (layer4_outputs(1482));
    outputs(6181) <= layer4_outputs(6747);
    outputs(6182) <= not((layer4_outputs(2127)) and (layer4_outputs(4445)));
    outputs(6183) <= (layer4_outputs(8385)) xor (layer4_outputs(7511));
    outputs(6184) <= layer4_outputs(8391);
    outputs(6185) <= layer4_outputs(6598);
    outputs(6186) <= not(layer4_outputs(10146));
    outputs(6187) <= not((layer4_outputs(578)) xor (layer4_outputs(9216)));
    outputs(6188) <= layer4_outputs(9161);
    outputs(6189) <= layer4_outputs(5494);
    outputs(6190) <= not((layer4_outputs(9831)) xor (layer4_outputs(5845)));
    outputs(6191) <= not(layer4_outputs(4900));
    outputs(6192) <= not(layer4_outputs(6317));
    outputs(6193) <= (layer4_outputs(1456)) or (layer4_outputs(8265));
    outputs(6194) <= not(layer4_outputs(346));
    outputs(6195) <= not(layer4_outputs(8892));
    outputs(6196) <= layer4_outputs(9070);
    outputs(6197) <= layer4_outputs(10162);
    outputs(6198) <= layer4_outputs(9182);
    outputs(6199) <= not(layer4_outputs(6773));
    outputs(6200) <= not(layer4_outputs(8629));
    outputs(6201) <= layer4_outputs(553);
    outputs(6202) <= not(layer4_outputs(9044));
    outputs(6203) <= not(layer4_outputs(7380));
    outputs(6204) <= layer4_outputs(4683);
    outputs(6205) <= layer4_outputs(3371);
    outputs(6206) <= layer4_outputs(647);
    outputs(6207) <= not(layer4_outputs(5648));
    outputs(6208) <= layer4_outputs(3138);
    outputs(6209) <= layer4_outputs(67);
    outputs(6210) <= (layer4_outputs(7613)) and not (layer4_outputs(9489));
    outputs(6211) <= layer4_outputs(9149);
    outputs(6212) <= layer4_outputs(8156);
    outputs(6213) <= not(layer4_outputs(9788)) or (layer4_outputs(852));
    outputs(6214) <= layer4_outputs(2963);
    outputs(6215) <= layer4_outputs(7011);
    outputs(6216) <= (layer4_outputs(4493)) xor (layer4_outputs(429));
    outputs(6217) <= (layer4_outputs(3185)) xor (layer4_outputs(4474));
    outputs(6218) <= not((layer4_outputs(7103)) xor (layer4_outputs(6960)));
    outputs(6219) <= (layer4_outputs(9682)) and not (layer4_outputs(6658));
    outputs(6220) <= (layer4_outputs(1535)) xor (layer4_outputs(5255));
    outputs(6221) <= layer4_outputs(3559);
    outputs(6222) <= not(layer4_outputs(3902));
    outputs(6223) <= not(layer4_outputs(8555));
    outputs(6224) <= not((layer4_outputs(9316)) xor (layer4_outputs(4824)));
    outputs(6225) <= not(layer4_outputs(9552));
    outputs(6226) <= not(layer4_outputs(9278));
    outputs(6227) <= not(layer4_outputs(8090));
    outputs(6228) <= not(layer4_outputs(2658));
    outputs(6229) <= not(layer4_outputs(1790));
    outputs(6230) <= (layer4_outputs(3855)) or (layer4_outputs(8853));
    outputs(6231) <= not(layer4_outputs(7488));
    outputs(6232) <= layer4_outputs(1682);
    outputs(6233) <= not(layer4_outputs(5077));
    outputs(6234) <= not(layer4_outputs(2851));
    outputs(6235) <= layer4_outputs(3624);
    outputs(6236) <= (layer4_outputs(7594)) xor (layer4_outputs(3370));
    outputs(6237) <= not(layer4_outputs(10075));
    outputs(6238) <= layer4_outputs(3990);
    outputs(6239) <= not(layer4_outputs(4614));
    outputs(6240) <= layer4_outputs(4766);
    outputs(6241) <= not(layer4_outputs(5729));
    outputs(6242) <= layer4_outputs(6536);
    outputs(6243) <= not(layer4_outputs(2632));
    outputs(6244) <= layer4_outputs(3082);
    outputs(6245) <= not(layer4_outputs(35));
    outputs(6246) <= (layer4_outputs(8838)) and not (layer4_outputs(880));
    outputs(6247) <= layer4_outputs(4722);
    outputs(6248) <= not(layer4_outputs(3897));
    outputs(6249) <= (layer4_outputs(7018)) xor (layer4_outputs(2126));
    outputs(6250) <= not((layer4_outputs(3543)) xor (layer4_outputs(80)));
    outputs(6251) <= layer4_outputs(4483);
    outputs(6252) <= not(layer4_outputs(3565));
    outputs(6253) <= (layer4_outputs(7851)) xor (layer4_outputs(3745));
    outputs(6254) <= layer4_outputs(9151);
    outputs(6255) <= layer4_outputs(6177);
    outputs(6256) <= not((layer4_outputs(216)) or (layer4_outputs(3662)));
    outputs(6257) <= not((layer4_outputs(4461)) xor (layer4_outputs(6781)));
    outputs(6258) <= (layer4_outputs(9386)) xor (layer4_outputs(7461));
    outputs(6259) <= layer4_outputs(7092);
    outputs(6260) <= layer4_outputs(9979);
    outputs(6261) <= not(layer4_outputs(6315));
    outputs(6262) <= not(layer4_outputs(3454));
    outputs(6263) <= not(layer4_outputs(4833));
    outputs(6264) <= (layer4_outputs(674)) xor (layer4_outputs(6364));
    outputs(6265) <= layer4_outputs(2770);
    outputs(6266) <= not(layer4_outputs(5019));
    outputs(6267) <= (layer4_outputs(5315)) and not (layer4_outputs(9779));
    outputs(6268) <= not(layer4_outputs(7450));
    outputs(6269) <= layer4_outputs(9973);
    outputs(6270) <= layer4_outputs(1694);
    outputs(6271) <= not(layer4_outputs(7397));
    outputs(6272) <= layer4_outputs(4363);
    outputs(6273) <= not((layer4_outputs(9584)) xor (layer4_outputs(2934)));
    outputs(6274) <= not(layer4_outputs(8911));
    outputs(6275) <= not(layer4_outputs(6756));
    outputs(6276) <= not(layer4_outputs(1813));
    outputs(6277) <= (layer4_outputs(1369)) or (layer4_outputs(8544));
    outputs(6278) <= (layer4_outputs(9903)) xor (layer4_outputs(9661));
    outputs(6279) <= not(layer4_outputs(6226));
    outputs(6280) <= not((layer4_outputs(6829)) or (layer4_outputs(7057)));
    outputs(6281) <= layer4_outputs(8139);
    outputs(6282) <= layer4_outputs(3775);
    outputs(6283) <= layer4_outputs(9939);
    outputs(6284) <= layer4_outputs(2533);
    outputs(6285) <= layer4_outputs(5810);
    outputs(6286) <= not(layer4_outputs(8301));
    outputs(6287) <= layer4_outputs(4140);
    outputs(6288) <= not(layer4_outputs(8038));
    outputs(6289) <= not(layer4_outputs(5362));
    outputs(6290) <= (layer4_outputs(4382)) and not (layer4_outputs(3666));
    outputs(6291) <= layer4_outputs(3012);
    outputs(6292) <= layer4_outputs(7326);
    outputs(6293) <= layer4_outputs(8092);
    outputs(6294) <= layer4_outputs(2037);
    outputs(6295) <= layer4_outputs(8202);
    outputs(6296) <= not(layer4_outputs(5849));
    outputs(6297) <= not(layer4_outputs(2221));
    outputs(6298) <= layer4_outputs(8817);
    outputs(6299) <= not((layer4_outputs(9223)) and (layer4_outputs(6901)));
    outputs(6300) <= not(layer4_outputs(4052)) or (layer4_outputs(4624));
    outputs(6301) <= (layer4_outputs(3004)) and not (layer4_outputs(34));
    outputs(6302) <= layer4_outputs(7231);
    outputs(6303) <= not((layer4_outputs(10184)) xor (layer4_outputs(5027)));
    outputs(6304) <= layer4_outputs(8730);
    outputs(6305) <= not(layer4_outputs(3211));
    outputs(6306) <= layer4_outputs(7310);
    outputs(6307) <= not(layer4_outputs(920));
    outputs(6308) <= (layer4_outputs(8384)) and not (layer4_outputs(9953));
    outputs(6309) <= not((layer4_outputs(7982)) or (layer4_outputs(588)));
    outputs(6310) <= not(layer4_outputs(5228));
    outputs(6311) <= not(layer4_outputs(6028));
    outputs(6312) <= not(layer4_outputs(10214));
    outputs(6313) <= layer4_outputs(3868);
    outputs(6314) <= not(layer4_outputs(6712));
    outputs(6315) <= layer4_outputs(8668);
    outputs(6316) <= layer4_outputs(1947);
    outputs(6317) <= (layer4_outputs(2849)) xor (layer4_outputs(5911));
    outputs(6318) <= layer4_outputs(1308);
    outputs(6319) <= (layer4_outputs(6200)) or (layer4_outputs(5127));
    outputs(6320) <= layer4_outputs(2834);
    outputs(6321) <= layer4_outputs(4779);
    outputs(6322) <= layer4_outputs(4448);
    outputs(6323) <= not((layer4_outputs(1752)) xor (layer4_outputs(6699)));
    outputs(6324) <= not(layer4_outputs(9226));
    outputs(6325) <= layer4_outputs(1884);
    outputs(6326) <= layer4_outputs(7224);
    outputs(6327) <= not(layer4_outputs(9145));
    outputs(6328) <= layer4_outputs(2045);
    outputs(6329) <= (layer4_outputs(9729)) and not (layer4_outputs(4062));
    outputs(6330) <= layer4_outputs(663);
    outputs(6331) <= not(layer4_outputs(112));
    outputs(6332) <= not(layer4_outputs(3125)) or (layer4_outputs(9792));
    outputs(6333) <= not(layer4_outputs(3207));
    outputs(6334) <= layer4_outputs(16);
    outputs(6335) <= layer4_outputs(8399);
    outputs(6336) <= not((layer4_outputs(8063)) xor (layer4_outputs(4123)));
    outputs(6337) <= layer4_outputs(937);
    outputs(6338) <= not((layer4_outputs(8912)) or (layer4_outputs(10097)));
    outputs(6339) <= not(layer4_outputs(6424));
    outputs(6340) <= layer4_outputs(5727);
    outputs(6341) <= (layer4_outputs(7600)) and not (layer4_outputs(5688));
    outputs(6342) <= (layer4_outputs(4146)) xor (layer4_outputs(9048));
    outputs(6343) <= not((layer4_outputs(7721)) xor (layer4_outputs(1073)));
    outputs(6344) <= not(layer4_outputs(8103));
    outputs(6345) <= (layer4_outputs(4455)) and (layer4_outputs(1109));
    outputs(6346) <= layer4_outputs(525);
    outputs(6347) <= not(layer4_outputs(2435));
    outputs(6348) <= not(layer4_outputs(7135));
    outputs(6349) <= not(layer4_outputs(5374)) or (layer4_outputs(2158));
    outputs(6350) <= not(layer4_outputs(3375));
    outputs(6351) <= not(layer4_outputs(261));
    outputs(6352) <= not(layer4_outputs(7277));
    outputs(6353) <= not(layer4_outputs(8821));
    outputs(6354) <= layer4_outputs(6118);
    outputs(6355) <= (layer4_outputs(517)) xor (layer4_outputs(10120));
    outputs(6356) <= not((layer4_outputs(6813)) or (layer4_outputs(2544)));
    outputs(6357) <= layer4_outputs(9424);
    outputs(6358) <= layer4_outputs(9607);
    outputs(6359) <= not(layer4_outputs(2464));
    outputs(6360) <= not((layer4_outputs(7104)) or (layer4_outputs(3248)));
    outputs(6361) <= not(layer4_outputs(8537));
    outputs(6362) <= (layer4_outputs(7032)) xor (layer4_outputs(4184));
    outputs(6363) <= not(layer4_outputs(741));
    outputs(6364) <= layer4_outputs(8457);
    outputs(6365) <= layer4_outputs(10126);
    outputs(6366) <= not(layer4_outputs(2462));
    outputs(6367) <= (layer4_outputs(1641)) xor (layer4_outputs(8277));
    outputs(6368) <= layer4_outputs(9610);
    outputs(6369) <= not(layer4_outputs(7932));
    outputs(6370) <= layer4_outputs(3720);
    outputs(6371) <= not(layer4_outputs(3330)) or (layer4_outputs(1386));
    outputs(6372) <= not(layer4_outputs(7420)) or (layer4_outputs(9469));
    outputs(6373) <= not(layer4_outputs(1229));
    outputs(6374) <= layer4_outputs(7695);
    outputs(6375) <= (layer4_outputs(3602)) or (layer4_outputs(2442));
    outputs(6376) <= (layer4_outputs(2203)) xor (layer4_outputs(2650));
    outputs(6377) <= not(layer4_outputs(8659));
    outputs(6378) <= '1';
    outputs(6379) <= layer4_outputs(1797);
    outputs(6380) <= layer4_outputs(1115);
    outputs(6381) <= layer4_outputs(1486);
    outputs(6382) <= not(layer4_outputs(8749));
    outputs(6383) <= layer4_outputs(40);
    outputs(6384) <= not(layer4_outputs(8002));
    outputs(6385) <= not(layer4_outputs(5640));
    outputs(6386) <= not(layer4_outputs(549));
    outputs(6387) <= layer4_outputs(4655);
    outputs(6388) <= not((layer4_outputs(4832)) xor (layer4_outputs(8329)));
    outputs(6389) <= layer4_outputs(1372);
    outputs(6390) <= not(layer4_outputs(3918));
    outputs(6391) <= not(layer4_outputs(7854));
    outputs(6392) <= not(layer4_outputs(3074));
    outputs(6393) <= not(layer4_outputs(3127));
    outputs(6394) <= not(layer4_outputs(3778));
    outputs(6395) <= (layer4_outputs(5406)) xor (layer4_outputs(5891));
    outputs(6396) <= not((layer4_outputs(6762)) xor (layer4_outputs(108)));
    outputs(6397) <= not(layer4_outputs(9402));
    outputs(6398) <= layer4_outputs(8010);
    outputs(6399) <= layer4_outputs(2518);
    outputs(6400) <= not(layer4_outputs(5519));
    outputs(6401) <= not(layer4_outputs(8106)) or (layer4_outputs(9423));
    outputs(6402) <= layer4_outputs(5716);
    outputs(6403) <= layer4_outputs(4794);
    outputs(6404) <= layer4_outputs(2925);
    outputs(6405) <= not(layer4_outputs(9255));
    outputs(6406) <= not(layer4_outputs(10107)) or (layer4_outputs(1427));
    outputs(6407) <= layer4_outputs(8461);
    outputs(6408) <= layer4_outputs(1586);
    outputs(6409) <= not((layer4_outputs(3587)) xor (layer4_outputs(7029)));
    outputs(6410) <= layer4_outputs(8194);
    outputs(6411) <= not(layer4_outputs(2782));
    outputs(6412) <= not(layer4_outputs(1594));
    outputs(6413) <= not(layer4_outputs(9604));
    outputs(6414) <= not(layer4_outputs(3912));
    outputs(6415) <= not(layer4_outputs(359));
    outputs(6416) <= layer4_outputs(2552);
    outputs(6417) <= not((layer4_outputs(4401)) xor (layer4_outputs(6213)));
    outputs(6418) <= (layer4_outputs(9237)) and (layer4_outputs(2234));
    outputs(6419) <= not(layer4_outputs(8192)) or (layer4_outputs(9463));
    outputs(6420) <= not(layer4_outputs(7735));
    outputs(6421) <= (layer4_outputs(9646)) and not (layer4_outputs(7760));
    outputs(6422) <= not((layer4_outputs(3649)) and (layer4_outputs(6469)));
    outputs(6423) <= not(layer4_outputs(6119));
    outputs(6424) <= layer4_outputs(5175);
    outputs(6425) <= layer4_outputs(8780);
    outputs(6426) <= layer4_outputs(8496);
    outputs(6427) <= not((layer4_outputs(1232)) or (layer4_outputs(2227)));
    outputs(6428) <= (layer4_outputs(8690)) xor (layer4_outputs(1089));
    outputs(6429) <= layer4_outputs(7448);
    outputs(6430) <= layer4_outputs(472);
    outputs(6431) <= layer4_outputs(357);
    outputs(6432) <= not(layer4_outputs(1667));
    outputs(6433) <= not((layer4_outputs(9989)) xor (layer4_outputs(7522)));
    outputs(6434) <= layer4_outputs(4739);
    outputs(6435) <= not((layer4_outputs(5989)) xor (layer4_outputs(4602)));
    outputs(6436) <= (layer4_outputs(3014)) xor (layer4_outputs(9885));
    outputs(6437) <= layer4_outputs(3142);
    outputs(6438) <= not(layer4_outputs(7858));
    outputs(6439) <= not(layer4_outputs(8338));
    outputs(6440) <= layer4_outputs(9316);
    outputs(6441) <= not(layer4_outputs(4808));
    outputs(6442) <= (layer4_outputs(9795)) and not (layer4_outputs(2348));
    outputs(6443) <= not((layer4_outputs(8157)) or (layer4_outputs(2771)));
    outputs(6444) <= layer4_outputs(2523);
    outputs(6445) <= not((layer4_outputs(5210)) xor (layer4_outputs(7209)));
    outputs(6446) <= layer4_outputs(3837);
    outputs(6447) <= not(layer4_outputs(3931));
    outputs(6448) <= (layer4_outputs(9224)) xor (layer4_outputs(4489));
    outputs(6449) <= layer4_outputs(6196);
    outputs(6450) <= not(layer4_outputs(9615));
    outputs(6451) <= layer4_outputs(1973);
    outputs(6452) <= (layer4_outputs(9505)) xor (layer4_outputs(8507));
    outputs(6453) <= layer4_outputs(2022);
    outputs(6454) <= not((layer4_outputs(485)) xor (layer4_outputs(1501)));
    outputs(6455) <= layer4_outputs(4024);
    outputs(6456) <= layer4_outputs(4770);
    outputs(6457) <= layer4_outputs(1486);
    outputs(6458) <= (layer4_outputs(8794)) xor (layer4_outputs(826));
    outputs(6459) <= not(layer4_outputs(8771));
    outputs(6460) <= not(layer4_outputs(1522));
    outputs(6461) <= layer4_outputs(8144);
    outputs(6462) <= layer4_outputs(746);
    outputs(6463) <= (layer4_outputs(9640)) xor (layer4_outputs(4870));
    outputs(6464) <= layer4_outputs(3647);
    outputs(6465) <= not(layer4_outputs(4392));
    outputs(6466) <= not(layer4_outputs(5503)) or (layer4_outputs(3583));
    outputs(6467) <= layer4_outputs(1338);
    outputs(6468) <= layer4_outputs(8510);
    outputs(6469) <= not(layer4_outputs(3044));
    outputs(6470) <= not(layer4_outputs(5405));
    outputs(6471) <= not(layer4_outputs(6330));
    outputs(6472) <= not(layer4_outputs(2023));
    outputs(6473) <= layer4_outputs(2600);
    outputs(6474) <= not(layer4_outputs(4725));
    outputs(6475) <= layer4_outputs(3477);
    outputs(6476) <= (layer4_outputs(9089)) xor (layer4_outputs(3437));
    outputs(6477) <= not((layer4_outputs(5952)) xor (layer4_outputs(1350)));
    outputs(6478) <= (layer4_outputs(8296)) xor (layer4_outputs(8235));
    outputs(6479) <= not(layer4_outputs(6195));
    outputs(6480) <= (layer4_outputs(5417)) xor (layer4_outputs(344));
    outputs(6481) <= layer4_outputs(4030);
    outputs(6482) <= not((layer4_outputs(8519)) xor (layer4_outputs(2150)));
    outputs(6483) <= (layer4_outputs(3987)) and (layer4_outputs(1055));
    outputs(6484) <= not(layer4_outputs(834)) or (layer4_outputs(3928));
    outputs(6485) <= not((layer4_outputs(7625)) and (layer4_outputs(3832)));
    outputs(6486) <= not(layer4_outputs(2884));
    outputs(6487) <= (layer4_outputs(1504)) xor (layer4_outputs(6166));
    outputs(6488) <= layer4_outputs(1728);
    outputs(6489) <= layer4_outputs(6475);
    outputs(6490) <= not((layer4_outputs(8346)) xor (layer4_outputs(7013)));
    outputs(6491) <= (layer4_outputs(408)) xor (layer4_outputs(7365));
    outputs(6492) <= not((layer4_outputs(2123)) or (layer4_outputs(8415)));
    outputs(6493) <= not((layer4_outputs(9906)) xor (layer4_outputs(4137)));
    outputs(6494) <= not(layer4_outputs(1964));
    outputs(6495) <= (layer4_outputs(3289)) and not (layer4_outputs(799));
    outputs(6496) <= (layer4_outputs(3040)) xor (layer4_outputs(5199));
    outputs(6497) <= not(layer4_outputs(2571));
    outputs(6498) <= not((layer4_outputs(397)) xor (layer4_outputs(9831)));
    outputs(6499) <= layer4_outputs(5441);
    outputs(6500) <= not(layer4_outputs(7824));
    outputs(6501) <= not(layer4_outputs(2772));
    outputs(6502) <= layer4_outputs(8004);
    outputs(6503) <= (layer4_outputs(6875)) and not (layer4_outputs(8729));
    outputs(6504) <= not(layer4_outputs(4056));
    outputs(6505) <= not(layer4_outputs(8287));
    outputs(6506) <= layer4_outputs(5176);
    outputs(6507) <= not(layer4_outputs(3353));
    outputs(6508) <= layer4_outputs(7108);
    outputs(6509) <= not((layer4_outputs(1695)) xor (layer4_outputs(6560)));
    outputs(6510) <= layer4_outputs(2751);
    outputs(6511) <= (layer4_outputs(9499)) or (layer4_outputs(3122));
    outputs(6512) <= (layer4_outputs(8116)) and (layer4_outputs(6700));
    outputs(6513) <= layer4_outputs(9683);
    outputs(6514) <= not(layer4_outputs(9874));
    outputs(6515) <= not((layer4_outputs(173)) xor (layer4_outputs(9864)));
    outputs(6516) <= layer4_outputs(4455);
    outputs(6517) <= not(layer4_outputs(1820));
    outputs(6518) <= not((layer4_outputs(1842)) xor (layer4_outputs(2796)));
    outputs(6519) <= not((layer4_outputs(1146)) xor (layer4_outputs(8442)));
    outputs(6520) <= layer4_outputs(2134);
    outputs(6521) <= not(layer4_outputs(4437));
    outputs(6522) <= not(layer4_outputs(5831));
    outputs(6523) <= not(layer4_outputs(4219));
    outputs(6524) <= not((layer4_outputs(1932)) and (layer4_outputs(2878)));
    outputs(6525) <= not(layer4_outputs(8523));
    outputs(6526) <= not(layer4_outputs(6235));
    outputs(6527) <= layer4_outputs(3590);
    outputs(6528) <= layer4_outputs(8201);
    outputs(6529) <= not((layer4_outputs(5803)) xor (layer4_outputs(2125)));
    outputs(6530) <= not(layer4_outputs(914)) or (layer4_outputs(9181));
    outputs(6531) <= layer4_outputs(2596);
    outputs(6532) <= layer4_outputs(9320);
    outputs(6533) <= layer4_outputs(7338);
    outputs(6534) <= not(layer4_outputs(3267));
    outputs(6535) <= not(layer4_outputs(2123));
    outputs(6536) <= layer4_outputs(6986);
    outputs(6537) <= layer4_outputs(6551);
    outputs(6538) <= not((layer4_outputs(6602)) xor (layer4_outputs(883)));
    outputs(6539) <= layer4_outputs(6899);
    outputs(6540) <= layer4_outputs(3967);
    outputs(6541) <= layer4_outputs(5571);
    outputs(6542) <= (layer4_outputs(9757)) or (layer4_outputs(9301));
    outputs(6543) <= not(layer4_outputs(9231));
    outputs(6544) <= not(layer4_outputs(6351));
    outputs(6545) <= not((layer4_outputs(7136)) and (layer4_outputs(9971)));
    outputs(6546) <= (layer4_outputs(9233)) and not (layer4_outputs(3651));
    outputs(6547) <= not(layer4_outputs(7154)) or (layer4_outputs(2124));
    outputs(6548) <= (layer4_outputs(3465)) and not (layer4_outputs(3044));
    outputs(6549) <= not(layer4_outputs(2212));
    outputs(6550) <= not(layer4_outputs(2109));
    outputs(6551) <= layer4_outputs(6884);
    outputs(6552) <= not(layer4_outputs(2571));
    outputs(6553) <= not(layer4_outputs(6305));
    outputs(6554) <= not((layer4_outputs(3722)) xor (layer4_outputs(7285)));
    outputs(6555) <= not((layer4_outputs(8877)) xor (layer4_outputs(1349)));
    outputs(6556) <= not(layer4_outputs(1406));
    outputs(6557) <= not((layer4_outputs(2010)) and (layer4_outputs(2049)));
    outputs(6558) <= (layer4_outputs(1233)) xor (layer4_outputs(9242));
    outputs(6559) <= layer4_outputs(2800);
    outputs(6560) <= not((layer4_outputs(192)) xor (layer4_outputs(5536)));
    outputs(6561) <= not(layer4_outputs(2999));
    outputs(6562) <= not(layer4_outputs(7048));
    outputs(6563) <= not(layer4_outputs(6286));
    outputs(6564) <= layer4_outputs(5460);
    outputs(6565) <= not(layer4_outputs(10209));
    outputs(6566) <= not(layer4_outputs(5274));
    outputs(6567) <= layer4_outputs(4719);
    outputs(6568) <= not(layer4_outputs(1167));
    outputs(6569) <= (layer4_outputs(9999)) xor (layer4_outputs(1166));
    outputs(6570) <= layer4_outputs(2834);
    outputs(6571) <= layer4_outputs(9822);
    outputs(6572) <= not((layer4_outputs(361)) xor (layer4_outputs(6484)));
    outputs(6573) <= layer4_outputs(5781);
    outputs(6574) <= layer4_outputs(4784);
    outputs(6575) <= layer4_outputs(528);
    outputs(6576) <= not((layer4_outputs(9352)) xor (layer4_outputs(10195)));
    outputs(6577) <= not(layer4_outputs(9274));
    outputs(6578) <= layer4_outputs(8030);
    outputs(6579) <= not(layer4_outputs(7341));
    outputs(6580) <= layer4_outputs(3572);
    outputs(6581) <= (layer4_outputs(3090)) xor (layer4_outputs(9111));
    outputs(6582) <= not(layer4_outputs(8486));
    outputs(6583) <= not(layer4_outputs(187));
    outputs(6584) <= not((layer4_outputs(10104)) xor (layer4_outputs(161)));
    outputs(6585) <= layer4_outputs(3144);
    outputs(6586) <= (layer4_outputs(3103)) and (layer4_outputs(7543));
    outputs(6587) <= not((layer4_outputs(5493)) xor (layer4_outputs(2758)));
    outputs(6588) <= (layer4_outputs(8955)) or (layer4_outputs(3619));
    outputs(6589) <= (layer4_outputs(6175)) xor (layer4_outputs(5507));
    outputs(6590) <= not(layer4_outputs(4743));
    outputs(6591) <= not((layer4_outputs(9544)) xor (layer4_outputs(2514)));
    outputs(6592) <= not(layer4_outputs(7017)) or (layer4_outputs(2670));
    outputs(6593) <= layer4_outputs(1434);
    outputs(6594) <= not(layer4_outputs(9857));
    outputs(6595) <= layer4_outputs(2940);
    outputs(6596) <= layer4_outputs(843);
    outputs(6597) <= layer4_outputs(2096);
    outputs(6598) <= not(layer4_outputs(7792));
    outputs(6599) <= not((layer4_outputs(7682)) xor (layer4_outputs(6694)));
    outputs(6600) <= layer4_outputs(3008);
    outputs(6601) <= (layer4_outputs(9895)) or (layer4_outputs(2005));
    outputs(6602) <= not(layer4_outputs(634));
    outputs(6603) <= (layer4_outputs(1134)) xor (layer4_outputs(3650));
    outputs(6604) <= not(layer4_outputs(9564));
    outputs(6605) <= layer4_outputs(4173);
    outputs(6606) <= not(layer4_outputs(5145));
    outputs(6607) <= (layer4_outputs(10056)) and not (layer4_outputs(1445));
    outputs(6608) <= layer4_outputs(1769);
    outputs(6609) <= layer4_outputs(6667);
    outputs(6610) <= layer4_outputs(471);
    outputs(6611) <= (layer4_outputs(8060)) and (layer4_outputs(2853));
    outputs(6612) <= not(layer4_outputs(5707));
    outputs(6613) <= (layer4_outputs(5746)) and not (layer4_outputs(9513));
    outputs(6614) <= layer4_outputs(1683);
    outputs(6615) <= not(layer4_outputs(5968));
    outputs(6616) <= not(layer4_outputs(9753));
    outputs(6617) <= not((layer4_outputs(2975)) and (layer4_outputs(7800)));
    outputs(6618) <= not((layer4_outputs(2036)) xor (layer4_outputs(2612)));
    outputs(6619) <= not((layer4_outputs(7167)) xor (layer4_outputs(6702)));
    outputs(6620) <= layer4_outputs(4927);
    outputs(6621) <= layer4_outputs(7467);
    outputs(6622) <= layer4_outputs(3621);
    outputs(6623) <= not(layer4_outputs(1209));
    outputs(6624) <= not((layer4_outputs(3429)) xor (layer4_outputs(8793)));
    outputs(6625) <= not(layer4_outputs(5915));
    outputs(6626) <= layer4_outputs(8853);
    outputs(6627) <= not((layer4_outputs(195)) xor (layer4_outputs(4933)));
    outputs(6628) <= not(layer4_outputs(7816));
    outputs(6629) <= layer4_outputs(351);
    outputs(6630) <= (layer4_outputs(218)) and not (layer4_outputs(4292));
    outputs(6631) <= not(layer4_outputs(8249));
    outputs(6632) <= not(layer4_outputs(4006));
    outputs(6633) <= layer4_outputs(37);
    outputs(6634) <= not(layer4_outputs(270));
    outputs(6635) <= not((layer4_outputs(557)) xor (layer4_outputs(5483)));
    outputs(6636) <= not(layer4_outputs(10029));
    outputs(6637) <= (layer4_outputs(8959)) xor (layer4_outputs(2738));
    outputs(6638) <= (layer4_outputs(1610)) xor (layer4_outputs(9301));
    outputs(6639) <= not(layer4_outputs(1629));
    outputs(6640) <= (layer4_outputs(4269)) or (layer4_outputs(1699));
    outputs(6641) <= (layer4_outputs(4499)) xor (layer4_outputs(3390));
    outputs(6642) <= not(layer4_outputs(6684));
    outputs(6643) <= layer4_outputs(5476);
    outputs(6644) <= not(layer4_outputs(896));
    outputs(6645) <= not(layer4_outputs(8944));
    outputs(6646) <= not(layer4_outputs(1371)) or (layer4_outputs(6697));
    outputs(6647) <= (layer4_outputs(2364)) and (layer4_outputs(289));
    outputs(6648) <= (layer4_outputs(3033)) xor (layer4_outputs(8165));
    outputs(6649) <= (layer4_outputs(4705)) xor (layer4_outputs(2275));
    outputs(6650) <= layer4_outputs(1493);
    outputs(6651) <= not(layer4_outputs(4407));
    outputs(6652) <= not(layer4_outputs(7044));
    outputs(6653) <= not((layer4_outputs(7364)) xor (layer4_outputs(5619)));
    outputs(6654) <= not((layer4_outputs(9955)) and (layer4_outputs(2052)));
    outputs(6655) <= (layer4_outputs(8337)) and not (layer4_outputs(1783));
    outputs(6656) <= (layer4_outputs(3067)) xor (layer4_outputs(5406));
    outputs(6657) <= not(layer4_outputs(5880));
    outputs(6658) <= layer4_outputs(9915);
    outputs(6659) <= not(layer4_outputs(924));
    outputs(6660) <= (layer4_outputs(6217)) and not (layer4_outputs(9015));
    outputs(6661) <= (layer4_outputs(7124)) xor (layer4_outputs(7787));
    outputs(6662) <= (layer4_outputs(8627)) xor (layer4_outputs(10221));
    outputs(6663) <= not(layer4_outputs(3210));
    outputs(6664) <= layer4_outputs(3251);
    outputs(6665) <= not(layer4_outputs(9767));
    outputs(6666) <= not(layer4_outputs(8541));
    outputs(6667) <= (layer4_outputs(7155)) and not (layer4_outputs(7327));
    outputs(6668) <= not((layer4_outputs(7015)) or (layer4_outputs(737)));
    outputs(6669) <= not((layer4_outputs(2101)) and (layer4_outputs(5428)));
    outputs(6670) <= not(layer4_outputs(5756));
    outputs(6671) <= layer4_outputs(2659);
    outputs(6672) <= layer4_outputs(5041);
    outputs(6673) <= (layer4_outputs(5808)) xor (layer4_outputs(590));
    outputs(6674) <= layer4_outputs(5176);
    outputs(6675) <= (layer4_outputs(2812)) and not (layer4_outputs(8319));
    outputs(6676) <= not(layer4_outputs(5715));
    outputs(6677) <= not((layer4_outputs(1949)) xor (layer4_outputs(5276)));
    outputs(6678) <= not(layer4_outputs(1789));
    outputs(6679) <= not((layer4_outputs(7477)) xor (layer4_outputs(5430)));
    outputs(6680) <= (layer4_outputs(5212)) xor (layer4_outputs(1141));
    outputs(6681) <= (layer4_outputs(6453)) and not (layer4_outputs(9920));
    outputs(6682) <= not((layer4_outputs(7875)) xor (layer4_outputs(4583)));
    outputs(6683) <= not((layer4_outputs(7374)) xor (layer4_outputs(903)));
    outputs(6684) <= layer4_outputs(6787);
    outputs(6685) <= not((layer4_outputs(9493)) or (layer4_outputs(5140)));
    outputs(6686) <= layer4_outputs(8435);
    outputs(6687) <= not(layer4_outputs(6626));
    outputs(6688) <= not(layer4_outputs(1240));
    outputs(6689) <= (layer4_outputs(1795)) xor (layer4_outputs(1069));
    outputs(6690) <= not(layer4_outputs(386));
    outputs(6691) <= layer4_outputs(576);
    outputs(6692) <= (layer4_outputs(8390)) and not (layer4_outputs(5470));
    outputs(6693) <= not(layer4_outputs(2779));
    outputs(6694) <= layer4_outputs(7969);
    outputs(6695) <= not((layer4_outputs(2149)) xor (layer4_outputs(3302)));
    outputs(6696) <= layer4_outputs(7463);
    outputs(6697) <= (layer4_outputs(7840)) and not (layer4_outputs(2291));
    outputs(6698) <= not(layer4_outputs(6053));
    outputs(6699) <= not(layer4_outputs(4516));
    outputs(6700) <= layer4_outputs(9964);
    outputs(6701) <= not(layer4_outputs(7070));
    outputs(6702) <= not(layer4_outputs(8888));
    outputs(6703) <= not(layer4_outputs(8027)) or (layer4_outputs(597));
    outputs(6704) <= layer4_outputs(1749);
    outputs(6705) <= not(layer4_outputs(9297));
    outputs(6706) <= not(layer4_outputs(8595));
    outputs(6707) <= (layer4_outputs(615)) xor (layer4_outputs(2980));
    outputs(6708) <= (layer4_outputs(9558)) and not (layer4_outputs(7053));
    outputs(6709) <= not(layer4_outputs(5071));
    outputs(6710) <= layer4_outputs(7244);
    outputs(6711) <= not((layer4_outputs(1667)) xor (layer4_outputs(6843)));
    outputs(6712) <= not(layer4_outputs(364));
    outputs(6713) <= not((layer4_outputs(2531)) xor (layer4_outputs(1646)));
    outputs(6714) <= layer4_outputs(2688);
    outputs(6715) <= layer4_outputs(8842);
    outputs(6716) <= not(layer4_outputs(8326));
    outputs(6717) <= layer4_outputs(3079);
    outputs(6718) <= not(layer4_outputs(9738));
    outputs(6719) <= not((layer4_outputs(5547)) xor (layer4_outputs(1180)));
    outputs(6720) <= not((layer4_outputs(5809)) xor (layer4_outputs(8242)));
    outputs(6721) <= layer4_outputs(3343);
    outputs(6722) <= not(layer4_outputs(5202));
    outputs(6723) <= not(layer4_outputs(9872));
    outputs(6724) <= layer4_outputs(4315);
    outputs(6725) <= not((layer4_outputs(2210)) xor (layer4_outputs(1714)));
    outputs(6726) <= (layer4_outputs(7480)) and not (layer4_outputs(5602));
    outputs(6727) <= not(layer4_outputs(7336));
    outputs(6728) <= (layer4_outputs(8818)) xor (layer4_outputs(3174));
    outputs(6729) <= not((layer4_outputs(5573)) or (layer4_outputs(6407)));
    outputs(6730) <= (layer4_outputs(3170)) xor (layer4_outputs(4094));
    outputs(6731) <= not((layer4_outputs(4196)) xor (layer4_outputs(4772)));
    outputs(6732) <= not(layer4_outputs(2617));
    outputs(6733) <= layer4_outputs(7745);
    outputs(6734) <= layer4_outputs(5400);
    outputs(6735) <= (layer4_outputs(9678)) xor (layer4_outputs(9299));
    outputs(6736) <= not((layer4_outputs(5946)) xor (layer4_outputs(3876)));
    outputs(6737) <= not(layer4_outputs(8005));
    outputs(6738) <= not(layer4_outputs(8007));
    outputs(6739) <= not((layer4_outputs(8709)) xor (layer4_outputs(6438)));
    outputs(6740) <= not((layer4_outputs(5161)) xor (layer4_outputs(1451)));
    outputs(6741) <= layer4_outputs(2355);
    outputs(6742) <= not(layer4_outputs(5462));
    outputs(6743) <= (layer4_outputs(7323)) xor (layer4_outputs(4276));
    outputs(6744) <= not(layer4_outputs(3261));
    outputs(6745) <= not(layer4_outputs(4629));
    outputs(6746) <= not(layer4_outputs(623));
    outputs(6747) <= not(layer4_outputs(6906));
    outputs(6748) <= not(layer4_outputs(7110));
    outputs(6749) <= (layer4_outputs(7153)) xor (layer4_outputs(7352));
    outputs(6750) <= layer4_outputs(5139);
    outputs(6751) <= layer4_outputs(972);
    outputs(6752) <= (layer4_outputs(2358)) or (layer4_outputs(6021));
    outputs(6753) <= not(layer4_outputs(5645));
    outputs(6754) <= not(layer4_outputs(7333)) or (layer4_outputs(6969));
    outputs(6755) <= not(layer4_outputs(1909));
    outputs(6756) <= not(layer4_outputs(5884));
    outputs(6757) <= (layer4_outputs(7128)) xor (layer4_outputs(5694));
    outputs(6758) <= not(layer4_outputs(10077));
    outputs(6759) <= not(layer4_outputs(2490));
    outputs(6760) <= (layer4_outputs(7947)) xor (layer4_outputs(9586));
    outputs(6761) <= layer4_outputs(795);
    outputs(6762) <= not(layer4_outputs(2699));
    outputs(6763) <= layer4_outputs(2611);
    outputs(6764) <= not(layer4_outputs(9710)) or (layer4_outputs(3566));
    outputs(6765) <= not(layer4_outputs(4518));
    outputs(6766) <= layer4_outputs(8257);
    outputs(6767) <= not(layer4_outputs(1960));
    outputs(6768) <= not(layer4_outputs(6785));
    outputs(6769) <= layer4_outputs(7775);
    outputs(6770) <= layer4_outputs(9942);
    outputs(6771) <= not(layer4_outputs(5729));
    outputs(6772) <= layer4_outputs(3446);
    outputs(6773) <= (layer4_outputs(8823)) xor (layer4_outputs(7315));
    outputs(6774) <= not(layer4_outputs(6143));
    outputs(6775) <= not(layer4_outputs(6698));
    outputs(6776) <= layer4_outputs(6768);
    outputs(6777) <= (layer4_outputs(6539)) xor (layer4_outputs(9707));
    outputs(6778) <= layer4_outputs(663);
    outputs(6779) <= not(layer4_outputs(1805)) or (layer4_outputs(5371));
    outputs(6780) <= (layer4_outputs(116)) xor (layer4_outputs(7917));
    outputs(6781) <= layer4_outputs(3634);
    outputs(6782) <= layer4_outputs(6392);
    outputs(6783) <= not(layer4_outputs(2446));
    outputs(6784) <= not(layer4_outputs(9253));
    outputs(6785) <= (layer4_outputs(7120)) xor (layer4_outputs(1567));
    outputs(6786) <= not(layer4_outputs(871));
    outputs(6787) <= not((layer4_outputs(4855)) xor (layer4_outputs(558)));
    outputs(6788) <= (layer4_outputs(3711)) and not (layer4_outputs(9176));
    outputs(6789) <= layer4_outputs(2245);
    outputs(6790) <= not(layer4_outputs(107));
    outputs(6791) <= not((layer4_outputs(8919)) xor (layer4_outputs(4840)));
    outputs(6792) <= not((layer4_outputs(1028)) xor (layer4_outputs(2975)));
    outputs(6793) <= layer4_outputs(7832);
    outputs(6794) <= layer4_outputs(5186);
    outputs(6795) <= layer4_outputs(2508);
    outputs(6796) <= not((layer4_outputs(7706)) xor (layer4_outputs(2660)));
    outputs(6797) <= (layer4_outputs(3371)) or (layer4_outputs(8136));
    outputs(6798) <= not(layer4_outputs(752));
    outputs(6799) <= layer4_outputs(5793);
    outputs(6800) <= not(layer4_outputs(9201));
    outputs(6801) <= not(layer4_outputs(389));
    outputs(6802) <= (layer4_outputs(5781)) xor (layer4_outputs(2041));
    outputs(6803) <= not((layer4_outputs(4093)) xor (layer4_outputs(179)));
    outputs(6804) <= (layer4_outputs(2883)) and not (layer4_outputs(2998));
    outputs(6805) <= '1';
    outputs(6806) <= (layer4_outputs(8697)) or (layer4_outputs(3470));
    outputs(6807) <= not(layer4_outputs(5438));
    outputs(6808) <= not(layer4_outputs(4355));
    outputs(6809) <= layer4_outputs(609);
    outputs(6810) <= layer4_outputs(4401);
    outputs(6811) <= not((layer4_outputs(6263)) and (layer4_outputs(7363)));
    outputs(6812) <= layer4_outputs(3404);
    outputs(6813) <= not(layer4_outputs(1889));
    outputs(6814) <= layer4_outputs(5477);
    outputs(6815) <= layer4_outputs(10056);
    outputs(6816) <= '0';
    outputs(6817) <= not((layer4_outputs(8983)) xor (layer4_outputs(7499)));
    outputs(6818) <= layer4_outputs(6173);
    outputs(6819) <= layer4_outputs(8657);
    outputs(6820) <= layer4_outputs(9815);
    outputs(6821) <= not(layer4_outputs(234));
    outputs(6822) <= layer4_outputs(1640);
    outputs(6823) <= (layer4_outputs(7836)) xor (layer4_outputs(9719));
    outputs(6824) <= not((layer4_outputs(8339)) xor (layer4_outputs(2841)));
    outputs(6825) <= (layer4_outputs(946)) xor (layer4_outputs(8132));
    outputs(6826) <= not((layer4_outputs(6324)) xor (layer4_outputs(5819)));
    outputs(6827) <= layer4_outputs(10028);
    outputs(6828) <= not((layer4_outputs(2411)) xor (layer4_outputs(1004)));
    outputs(6829) <= layer4_outputs(5862);
    outputs(6830) <= (layer4_outputs(8745)) and (layer4_outputs(1267));
    outputs(6831) <= layer4_outputs(2916);
    outputs(6832) <= layer4_outputs(2071);
    outputs(6833) <= layer4_outputs(5975);
    outputs(6834) <= not((layer4_outputs(7052)) xor (layer4_outputs(3147)));
    outputs(6835) <= not((layer4_outputs(819)) xor (layer4_outputs(6613)));
    outputs(6836) <= layer4_outputs(1448);
    outputs(6837) <= layer4_outputs(171);
    outputs(6838) <= not(layer4_outputs(7808));
    outputs(6839) <= not((layer4_outputs(8768)) xor (layer4_outputs(80)));
    outputs(6840) <= not(layer4_outputs(6139));
    outputs(6841) <= layer4_outputs(7196);
    outputs(6842) <= '1';
    outputs(6843) <= not(layer4_outputs(8475));
    outputs(6844) <= (layer4_outputs(5885)) and not (layer4_outputs(6081));
    outputs(6845) <= not(layer4_outputs(8627)) or (layer4_outputs(4783));
    outputs(6846) <= layer4_outputs(1721);
    outputs(6847) <= not(layer4_outputs(7777));
    outputs(6848) <= not(layer4_outputs(8830));
    outputs(6849) <= (layer4_outputs(4777)) xor (layer4_outputs(3405));
    outputs(6850) <= not(layer4_outputs(9071));
    outputs(6851) <= not(layer4_outputs(2192));
    outputs(6852) <= (layer4_outputs(3609)) xor (layer4_outputs(9327));
    outputs(6853) <= not(layer4_outputs(6525));
    outputs(6854) <= not(layer4_outputs(3083));
    outputs(6855) <= (layer4_outputs(9986)) xor (layer4_outputs(2964));
    outputs(6856) <= not(layer4_outputs(7702));
    outputs(6857) <= layer4_outputs(4996);
    outputs(6858) <= (layer4_outputs(2941)) xor (layer4_outputs(9778));
    outputs(6859) <= not(layer4_outputs(1263));
    outputs(6860) <= not(layer4_outputs(5769));
    outputs(6861) <= not(layer4_outputs(1560));
    outputs(6862) <= not((layer4_outputs(1418)) xor (layer4_outputs(9681)));
    outputs(6863) <= layer4_outputs(9122);
    outputs(6864) <= not(layer4_outputs(7891));
    outputs(6865) <= (layer4_outputs(1874)) and not (layer4_outputs(5345));
    outputs(6866) <= (layer4_outputs(4058)) xor (layer4_outputs(8478));
    outputs(6867) <= (layer4_outputs(9656)) and not (layer4_outputs(2624));
    outputs(6868) <= not(layer4_outputs(6003));
    outputs(6869) <= layer4_outputs(8137);
    outputs(6870) <= layer4_outputs(3334);
    outputs(6871) <= (layer4_outputs(9065)) xor (layer4_outputs(6278));
    outputs(6872) <= (layer4_outputs(6783)) xor (layer4_outputs(52));
    outputs(6873) <= (layer4_outputs(1583)) xor (layer4_outputs(2701));
    outputs(6874) <= not(layer4_outputs(4541));
    outputs(6875) <= not((layer4_outputs(5832)) xor (layer4_outputs(6777)));
    outputs(6876) <= not(layer4_outputs(429));
    outputs(6877) <= not(layer4_outputs(9977)) or (layer4_outputs(6397));
    outputs(6878) <= not(layer4_outputs(10136));
    outputs(6879) <= layer4_outputs(8967);
    outputs(6880) <= layer4_outputs(2558);
    outputs(6881) <= layer4_outputs(5901);
    outputs(6882) <= not((layer4_outputs(1980)) and (layer4_outputs(6912)));
    outputs(6883) <= not(layer4_outputs(1333));
    outputs(6884) <= (layer4_outputs(5154)) xor (layer4_outputs(91));
    outputs(6885) <= not(layer4_outputs(6487));
    outputs(6886) <= layer4_outputs(1463);
    outputs(6887) <= not(layer4_outputs(5780));
    outputs(6888) <= not(layer4_outputs(4446));
    outputs(6889) <= not(layer4_outputs(5344));
    outputs(6890) <= (layer4_outputs(5123)) and not (layer4_outputs(6854));
    outputs(6891) <= not(layer4_outputs(2741));
    outputs(6892) <= layer4_outputs(4258);
    outputs(6893) <= not(layer4_outputs(3410));
    outputs(6894) <= layer4_outputs(7694);
    outputs(6895) <= layer4_outputs(4905);
    outputs(6896) <= not(layer4_outputs(983));
    outputs(6897) <= (layer4_outputs(8455)) xor (layer4_outputs(7313));
    outputs(6898) <= not((layer4_outputs(390)) or (layer4_outputs(2189)));
    outputs(6899) <= layer4_outputs(8871);
    outputs(6900) <= not(layer4_outputs(5532));
    outputs(6901) <= layer4_outputs(8756);
    outputs(6902) <= not(layer4_outputs(8924));
    outputs(6903) <= layer4_outputs(3116);
    outputs(6904) <= layer4_outputs(6784);
    outputs(6905) <= not((layer4_outputs(813)) xor (layer4_outputs(4079)));
    outputs(6906) <= not(layer4_outputs(3052)) or (layer4_outputs(4349));
    outputs(6907) <= not(layer4_outputs(6543));
    outputs(6908) <= not(layer4_outputs(4348));
    outputs(6909) <= not((layer4_outputs(4885)) xor (layer4_outputs(6383)));
    outputs(6910) <= not(layer4_outputs(4391));
    outputs(6911) <= not(layer4_outputs(6424));
    outputs(6912) <= not((layer4_outputs(1502)) xor (layer4_outputs(10083)));
    outputs(6913) <= layer4_outputs(6629);
    outputs(6914) <= not(layer4_outputs(3170)) or (layer4_outputs(8960));
    outputs(6915) <= not(layer4_outputs(7212));
    outputs(6916) <= not(layer4_outputs(7891));
    outputs(6917) <= not(layer4_outputs(9123));
    outputs(6918) <= not(layer4_outputs(10173));
    outputs(6919) <= not((layer4_outputs(787)) or (layer4_outputs(2715)));
    outputs(6920) <= not(layer4_outputs(392));
    outputs(6921) <= layer4_outputs(6238);
    outputs(6922) <= (layer4_outputs(5867)) xor (layer4_outputs(3898));
    outputs(6923) <= layer4_outputs(7606);
    outputs(6924) <= not((layer4_outputs(1386)) xor (layer4_outputs(4749)));
    outputs(6925) <= not(layer4_outputs(3677));
    outputs(6926) <= (layer4_outputs(2327)) and (layer4_outputs(6385));
    outputs(6927) <= not(layer4_outputs(2643)) or (layer4_outputs(8432));
    outputs(6928) <= (layer4_outputs(3332)) xor (layer4_outputs(7811));
    outputs(6929) <= layer4_outputs(7788);
    outputs(6930) <= not(layer4_outputs(7537));
    outputs(6931) <= (layer4_outputs(7612)) or (layer4_outputs(2566));
    outputs(6932) <= not(layer4_outputs(263));
    outputs(6933) <= layer4_outputs(5269);
    outputs(6934) <= not(layer4_outputs(4635));
    outputs(6935) <= (layer4_outputs(3124)) xor (layer4_outputs(3322));
    outputs(6936) <= (layer4_outputs(270)) xor (layer4_outputs(4179));
    outputs(6937) <= layer4_outputs(1870);
    outputs(6938) <= not(layer4_outputs(8268)) or (layer4_outputs(1814));
    outputs(6939) <= layer4_outputs(6258);
    outputs(6940) <= not((layer4_outputs(7916)) or (layer4_outputs(6013)));
    outputs(6941) <= not(layer4_outputs(2117));
    outputs(6942) <= (layer4_outputs(3037)) or (layer4_outputs(4624));
    outputs(6943) <= layer4_outputs(2297);
    outputs(6944) <= not(layer4_outputs(4735));
    outputs(6945) <= (layer4_outputs(2811)) xor (layer4_outputs(277));
    outputs(6946) <= not(layer4_outputs(2901));
    outputs(6947) <= layer4_outputs(9051);
    outputs(6948) <= not(layer4_outputs(6712));
    outputs(6949) <= layer4_outputs(9534);
    outputs(6950) <= not(layer4_outputs(300)) or (layer4_outputs(4200));
    outputs(6951) <= not(layer4_outputs(1243));
    outputs(6952) <= layer4_outputs(8780);
    outputs(6953) <= layer4_outputs(8045);
    outputs(6954) <= layer4_outputs(8229);
    outputs(6955) <= not(layer4_outputs(7696));
    outputs(6956) <= (layer4_outputs(341)) xor (layer4_outputs(3828));
    outputs(6957) <= not(layer4_outputs(217));
    outputs(6958) <= layer4_outputs(9254);
    outputs(6959) <= not(layer4_outputs(7916));
    outputs(6960) <= layer4_outputs(7467);
    outputs(6961) <= not(layer4_outputs(5267)) or (layer4_outputs(1122));
    outputs(6962) <= not(layer4_outputs(3054));
    outputs(6963) <= not(layer4_outputs(6525));
    outputs(6964) <= layer4_outputs(6197);
    outputs(6965) <= (layer4_outputs(6173)) or (layer4_outputs(8955));
    outputs(6966) <= not((layer4_outputs(9950)) xor (layer4_outputs(8013)));
    outputs(6967) <= (layer4_outputs(2497)) xor (layer4_outputs(7661));
    outputs(6968) <= (layer4_outputs(6902)) and not (layer4_outputs(34));
    outputs(6969) <= not(layer4_outputs(2496));
    outputs(6970) <= (layer4_outputs(5865)) and not (layer4_outputs(535));
    outputs(6971) <= not(layer4_outputs(6771));
    outputs(6972) <= not((layer4_outputs(5984)) xor (layer4_outputs(3601)));
    outputs(6973) <= not(layer4_outputs(4990));
    outputs(6974) <= layer4_outputs(6607);
    outputs(6975) <= layer4_outputs(8244);
    outputs(6976) <= layer4_outputs(6534);
    outputs(6977) <= not(layer4_outputs(712));
    outputs(6978) <= not((layer4_outputs(2082)) xor (layer4_outputs(4558)));
    outputs(6979) <= not(layer4_outputs(8802)) or (layer4_outputs(3674));
    outputs(6980) <= layer4_outputs(241);
    outputs(6981) <= not(layer4_outputs(6874));
    outputs(6982) <= (layer4_outputs(341)) and (layer4_outputs(9198));
    outputs(6983) <= layer4_outputs(3977);
    outputs(6984) <= (layer4_outputs(7459)) and (layer4_outputs(4684));
    outputs(6985) <= layer4_outputs(8685);
    outputs(6986) <= not(layer4_outputs(2478));
    outputs(6987) <= layer4_outputs(8726);
    outputs(6988) <= not(layer4_outputs(3535));
    outputs(6989) <= not(layer4_outputs(2368));
    outputs(6990) <= layer4_outputs(7189);
    outputs(6991) <= not(layer4_outputs(3562));
    outputs(6992) <= not(layer4_outputs(2337));
    outputs(6993) <= not(layer4_outputs(9509));
    outputs(6994) <= (layer4_outputs(6230)) and (layer4_outputs(5304));
    outputs(6995) <= not((layer4_outputs(9306)) xor (layer4_outputs(3399)));
    outputs(6996) <= not((layer4_outputs(7819)) xor (layer4_outputs(8910)));
    outputs(6997) <= not((layer4_outputs(9007)) xor (layer4_outputs(9934)));
    outputs(6998) <= (layer4_outputs(8282)) xor (layer4_outputs(9227));
    outputs(6999) <= layer4_outputs(8813);
    outputs(7000) <= (layer4_outputs(4406)) xor (layer4_outputs(4889));
    outputs(7001) <= not(layer4_outputs(932));
    outputs(7002) <= (layer4_outputs(8193)) xor (layer4_outputs(7215));
    outputs(7003) <= not(layer4_outputs(9924));
    outputs(7004) <= not(layer4_outputs(7705));
    outputs(7005) <= (layer4_outputs(129)) and not (layer4_outputs(2301));
    outputs(7006) <= not(layer4_outputs(7406)) or (layer4_outputs(2681));
    outputs(7007) <= not((layer4_outputs(1043)) or (layer4_outputs(6975)));
    outputs(7008) <= layer4_outputs(27);
    outputs(7009) <= layer4_outputs(3098);
    outputs(7010) <= not(layer4_outputs(5061));
    outputs(7011) <= layer4_outputs(5454);
    outputs(7012) <= layer4_outputs(6440);
    outputs(7013) <= layer4_outputs(10062);
    outputs(7014) <= not((layer4_outputs(1985)) xor (layer4_outputs(701)));
    outputs(7015) <= (layer4_outputs(4165)) xor (layer4_outputs(9392));
    outputs(7016) <= layer4_outputs(6428);
    outputs(7017) <= layer4_outputs(5521);
    outputs(7018) <= not(layer4_outputs(3329));
    outputs(7019) <= not(layer4_outputs(9991));
    outputs(7020) <= (layer4_outputs(3365)) xor (layer4_outputs(3909));
    outputs(7021) <= not((layer4_outputs(4589)) or (layer4_outputs(3702)));
    outputs(7022) <= layer4_outputs(5047);
    outputs(7023) <= (layer4_outputs(5064)) xor (layer4_outputs(4045));
    outputs(7024) <= (layer4_outputs(3431)) and (layer4_outputs(5643));
    outputs(7025) <= not(layer4_outputs(5796));
    outputs(7026) <= (layer4_outputs(2324)) or (layer4_outputs(4178));
    outputs(7027) <= not(layer4_outputs(5807)) or (layer4_outputs(3076));
    outputs(7028) <= layer4_outputs(2520);
    outputs(7029) <= layer4_outputs(8154);
    outputs(7030) <= not((layer4_outputs(8974)) xor (layer4_outputs(1347)));
    outputs(7031) <= not(layer4_outputs(4473));
    outputs(7032) <= layer4_outputs(1817);
    outputs(7033) <= not(layer4_outputs(9498));
    outputs(7034) <= layer4_outputs(8744);
    outputs(7035) <= not(layer4_outputs(8318)) or (layer4_outputs(3137));
    outputs(7036) <= not(layer4_outputs(3068)) or (layer4_outputs(9021));
    outputs(7037) <= not(layer4_outputs(6705));
    outputs(7038) <= not(layer4_outputs(512));
    outputs(7039) <= layer4_outputs(1743);
    outputs(7040) <= not(layer4_outputs(6194));
    outputs(7041) <= not(layer4_outputs(9184));
    outputs(7042) <= not(layer4_outputs(9047));
    outputs(7043) <= not(layer4_outputs(7604));
    outputs(7044) <= not(layer4_outputs(4423));
    outputs(7045) <= not(layer4_outputs(7334));
    outputs(7046) <= (layer4_outputs(3827)) xor (layer4_outputs(7874));
    outputs(7047) <= not(layer4_outputs(8727));
    outputs(7048) <= not(layer4_outputs(5171));
    outputs(7049) <= '1';
    outputs(7050) <= layer4_outputs(4144);
    outputs(7051) <= (layer4_outputs(8997)) xor (layer4_outputs(5611));
    outputs(7052) <= not(layer4_outputs(3733));
    outputs(7053) <= not(layer4_outputs(10130));
    outputs(7054) <= layer4_outputs(6776);
    outputs(7055) <= not(layer4_outputs(3016));
    outputs(7056) <= (layer4_outputs(404)) xor (layer4_outputs(9675));
    outputs(7057) <= layer4_outputs(3343);
    outputs(7058) <= not(layer4_outputs(8884));
    outputs(7059) <= not(layer4_outputs(9102));
    outputs(7060) <= layer4_outputs(8148);
    outputs(7061) <= (layer4_outputs(7528)) xor (layer4_outputs(7674));
    outputs(7062) <= not(layer4_outputs(8962));
    outputs(7063) <= not(layer4_outputs(1925));
    outputs(7064) <= not(layer4_outputs(2068));
    outputs(7065) <= not(layer4_outputs(3463));
    outputs(7066) <= (layer4_outputs(3739)) xor (layer4_outputs(5968));
    outputs(7067) <= layer4_outputs(9995);
    outputs(7068) <= not((layer4_outputs(2250)) xor (layer4_outputs(5293)));
    outputs(7069) <= layer4_outputs(4750);
    outputs(7070) <= not(layer4_outputs(9380));
    outputs(7071) <= not(layer4_outputs(203));
    outputs(7072) <= layer4_outputs(3385);
    outputs(7073) <= not((layer4_outputs(4305)) xor (layer4_outputs(912)));
    outputs(7074) <= not(layer4_outputs(9516)) or (layer4_outputs(5187));
    outputs(7075) <= layer4_outputs(7436);
    outputs(7076) <= not(layer4_outputs(3329));
    outputs(7077) <= not((layer4_outputs(6669)) or (layer4_outputs(6204)));
    outputs(7078) <= layer4_outputs(6961);
    outputs(7079) <= not((layer4_outputs(9596)) or (layer4_outputs(5189)));
    outputs(7080) <= '0';
    outputs(7081) <= not(layer4_outputs(6592));
    outputs(7082) <= (layer4_outputs(8585)) xor (layer4_outputs(7460));
    outputs(7083) <= layer4_outputs(7941);
    outputs(7084) <= (layer4_outputs(2098)) and (layer4_outputs(8359));
    outputs(7085) <= (layer4_outputs(72)) xor (layer4_outputs(5800));
    outputs(7086) <= not(layer4_outputs(2943));
    outputs(7087) <= not(layer4_outputs(6553));
    outputs(7088) <= not(layer4_outputs(2515));
    outputs(7089) <= layer4_outputs(1743);
    outputs(7090) <= layer4_outputs(8015);
    outputs(7091) <= not(layer4_outputs(10042));
    outputs(7092) <= not(layer4_outputs(557)) or (layer4_outputs(7617));
    outputs(7093) <= not(layer4_outputs(2171));
    outputs(7094) <= layer4_outputs(7622);
    outputs(7095) <= (layer4_outputs(2162)) xor (layer4_outputs(3980));
    outputs(7096) <= layer4_outputs(529);
    outputs(7097) <= (layer4_outputs(2548)) xor (layer4_outputs(935));
    outputs(7098) <= (layer4_outputs(5588)) xor (layer4_outputs(2174));
    outputs(7099) <= (layer4_outputs(4311)) xor (layer4_outputs(3572));
    outputs(7100) <= not((layer4_outputs(547)) xor (layer4_outputs(4810)));
    outputs(7101) <= layer4_outputs(8847);
    outputs(7102) <= not(layer4_outputs(79));
    outputs(7103) <= (layer4_outputs(3895)) or (layer4_outputs(8246));
    outputs(7104) <= (layer4_outputs(687)) xor (layer4_outputs(6328));
    outputs(7105) <= not(layer4_outputs(7764));
    outputs(7106) <= (layer4_outputs(6468)) and not (layer4_outputs(5230));
    outputs(7107) <= not(layer4_outputs(5663));
    outputs(7108) <= not(layer4_outputs(9909));
    outputs(7109) <= layer4_outputs(6069);
    outputs(7110) <= not((layer4_outputs(5452)) xor (layer4_outputs(1952)));
    outputs(7111) <= layer4_outputs(537);
    outputs(7112) <= not(layer4_outputs(2414));
    outputs(7113) <= not(layer4_outputs(2421));
    outputs(7114) <= not((layer4_outputs(5014)) xor (layer4_outputs(225)));
    outputs(7115) <= not((layer4_outputs(1954)) xor (layer4_outputs(149)));
    outputs(7116) <= not(layer4_outputs(888));
    outputs(7117) <= (layer4_outputs(1224)) xor (layer4_outputs(7821));
    outputs(7118) <= layer4_outputs(487);
    outputs(7119) <= layer4_outputs(7281);
    outputs(7120) <= layer4_outputs(9214);
    outputs(7121) <= (layer4_outputs(10119)) xor (layer4_outputs(8880));
    outputs(7122) <= not(layer4_outputs(1709)) or (layer4_outputs(5188));
    outputs(7123) <= not(layer4_outputs(7787));
    outputs(7124) <= layer4_outputs(6152);
    outputs(7125) <= not(layer4_outputs(5497));
    outputs(7126) <= (layer4_outputs(7276)) xor (layer4_outputs(813));
    outputs(7127) <= not(layer4_outputs(3395));
    outputs(7128) <= not((layer4_outputs(6338)) xor (layer4_outputs(7054)));
    outputs(7129) <= layer4_outputs(7366);
    outputs(7130) <= not(layer4_outputs(10080)) or (layer4_outputs(9067));
    outputs(7131) <= layer4_outputs(9557);
    outputs(7132) <= not(layer4_outputs(5829)) or (layer4_outputs(9227));
    outputs(7133) <= layer4_outputs(6898);
    outputs(7134) <= not(layer4_outputs(3235));
    outputs(7135) <= layer4_outputs(1035);
    outputs(7136) <= not(layer4_outputs(3594));
    outputs(7137) <= not(layer4_outputs(8444));
    outputs(7138) <= layer4_outputs(1270);
    outputs(7139) <= layer4_outputs(10071);
    outputs(7140) <= layer4_outputs(1354);
    outputs(7141) <= not(layer4_outputs(2577));
    outputs(7142) <= not(layer4_outputs(2090));
    outputs(7143) <= (layer4_outputs(6581)) and not (layer4_outputs(3561));
    outputs(7144) <= not(layer4_outputs(6588));
    outputs(7145) <= not(layer4_outputs(7279));
    outputs(7146) <= (layer4_outputs(72)) and not (layer4_outputs(3094));
    outputs(7147) <= not(layer4_outputs(5964));
    outputs(7148) <= (layer4_outputs(8386)) xor (layer4_outputs(8344));
    outputs(7149) <= not(layer4_outputs(3988));
    outputs(7150) <= layer4_outputs(2385);
    outputs(7151) <= layer4_outputs(3799);
    outputs(7152) <= not(layer4_outputs(3712));
    outputs(7153) <= (layer4_outputs(4985)) and not (layer4_outputs(8413));
    outputs(7154) <= layer4_outputs(7452);
    outputs(7155) <= (layer4_outputs(5697)) and (layer4_outputs(6456));
    outputs(7156) <= layer4_outputs(8147);
    outputs(7157) <= not(layer4_outputs(1886));
    outputs(7158) <= not((layer4_outputs(3182)) xor (layer4_outputs(3028)));
    outputs(7159) <= (layer4_outputs(2218)) xor (layer4_outputs(9724));
    outputs(7160) <= layer4_outputs(3647);
    outputs(7161) <= not(layer4_outputs(8835));
    outputs(7162) <= layer4_outputs(9104);
    outputs(7163) <= not(layer4_outputs(8347));
    outputs(7164) <= not((layer4_outputs(1546)) xor (layer4_outputs(9448)));
    outputs(7165) <= not(layer4_outputs(9262));
    outputs(7166) <= layer4_outputs(7431);
    outputs(7167) <= (layer4_outputs(1395)) and not (layer4_outputs(8415));
    outputs(7168) <= layer4_outputs(7437);
    outputs(7169) <= not(layer4_outputs(3653));
    outputs(7170) <= (layer4_outputs(8121)) xor (layer4_outputs(3481));
    outputs(7171) <= not(layer4_outputs(12));
    outputs(7172) <= not(layer4_outputs(504));
    outputs(7173) <= layer4_outputs(5321);
    outputs(7174) <= not(layer4_outputs(316));
    outputs(7175) <= not((layer4_outputs(6641)) xor (layer4_outputs(8136)));
    outputs(7176) <= not(layer4_outputs(1125));
    outputs(7177) <= not(layer4_outputs(1439));
    outputs(7178) <= layer4_outputs(7234);
    outputs(7179) <= '0';
    outputs(7180) <= layer4_outputs(4357);
    outputs(7181) <= not((layer4_outputs(8245)) or (layer4_outputs(1334)));
    outputs(7182) <= (layer4_outputs(2871)) and not (layer4_outputs(9083));
    outputs(7183) <= layer4_outputs(7055);
    outputs(7184) <= (layer4_outputs(9809)) xor (layer4_outputs(4946));
    outputs(7185) <= layer4_outputs(4742);
    outputs(7186) <= not(layer4_outputs(5136));
    outputs(7187) <= (layer4_outputs(1503)) or (layer4_outputs(9438));
    outputs(7188) <= (layer4_outputs(8885)) xor (layer4_outputs(7370));
    outputs(7189) <= (layer4_outputs(8894)) or (layer4_outputs(839));
    outputs(7190) <= layer4_outputs(2934);
    outputs(7191) <= layer4_outputs(8003);
    outputs(7192) <= (layer4_outputs(4066)) and not (layer4_outputs(6354));
    outputs(7193) <= not(layer4_outputs(9195));
    outputs(7194) <= not(layer4_outputs(488));
    outputs(7195) <= not(layer4_outputs(6255));
    outputs(7196) <= not(layer4_outputs(1205));
    outputs(7197) <= (layer4_outputs(6044)) xor (layer4_outputs(8124));
    outputs(7198) <= not(layer4_outputs(6050));
    outputs(7199) <= layer4_outputs(2976);
    outputs(7200) <= not(layer4_outputs(579));
    outputs(7201) <= layer4_outputs(9572);
    outputs(7202) <= not(layer4_outputs(8340));
    outputs(7203) <= layer4_outputs(2087);
    outputs(7204) <= not(layer4_outputs(5899)) or (layer4_outputs(3361));
    outputs(7205) <= layer4_outputs(4668);
    outputs(7206) <= layer4_outputs(6766);
    outputs(7207) <= layer4_outputs(4613);
    outputs(7208) <= layer4_outputs(5916);
    outputs(7209) <= not(layer4_outputs(164));
    outputs(7210) <= not(layer4_outputs(2524));
    outputs(7211) <= not(layer4_outputs(8044));
    outputs(7212) <= not(layer4_outputs(7284));
    outputs(7213) <= not(layer4_outputs(2864));
    outputs(7214) <= layer4_outputs(4687);
    outputs(7215) <= layer4_outputs(9295);
    outputs(7216) <= not(layer4_outputs(9807));
    outputs(7217) <= layer4_outputs(8117);
    outputs(7218) <= layer4_outputs(43);
    outputs(7219) <= layer4_outputs(649);
    outputs(7220) <= layer4_outputs(9925);
    outputs(7221) <= not(layer4_outputs(2672));
    outputs(7222) <= layer4_outputs(1707);
    outputs(7223) <= not(layer4_outputs(53));
    outputs(7224) <= layer4_outputs(9621);
    outputs(7225) <= not(layer4_outputs(2130));
    outputs(7226) <= not(layer4_outputs(802));
    outputs(7227) <= (layer4_outputs(2318)) and not (layer4_outputs(2648));
    outputs(7228) <= (layer4_outputs(3501)) xor (layer4_outputs(9855));
    outputs(7229) <= layer4_outputs(5636);
    outputs(7230) <= not((layer4_outputs(1048)) and (layer4_outputs(3040)));
    outputs(7231) <= layer4_outputs(2914);
    outputs(7232) <= layer4_outputs(4968);
    outputs(7233) <= layer4_outputs(9555);
    outputs(7234) <= not(layer4_outputs(8760));
    outputs(7235) <= layer4_outputs(6626);
    outputs(7236) <= not(layer4_outputs(2411));
    outputs(7237) <= layer4_outputs(9218);
    outputs(7238) <= not((layer4_outputs(3687)) xor (layer4_outputs(6774)));
    outputs(7239) <= not(layer4_outputs(2297));
    outputs(7240) <= (layer4_outputs(9496)) and not (layer4_outputs(7266));
    outputs(7241) <= not(layer4_outputs(981));
    outputs(7242) <= not((layer4_outputs(9161)) xor (layer4_outputs(5347)));
    outputs(7243) <= (layer4_outputs(10189)) and (layer4_outputs(5586));
    outputs(7244) <= not((layer4_outputs(2237)) xor (layer4_outputs(2579)));
    outputs(7245) <= not((layer4_outputs(8695)) xor (layer4_outputs(6051)));
    outputs(7246) <= (layer4_outputs(104)) xor (layer4_outputs(4039));
    outputs(7247) <= not(layer4_outputs(1797));
    outputs(7248) <= (layer4_outputs(3939)) xor (layer4_outputs(5));
    outputs(7249) <= layer4_outputs(5721);
    outputs(7250) <= not(layer4_outputs(8600));
    outputs(7251) <= not(layer4_outputs(7765));
    outputs(7252) <= layer4_outputs(1219);
    outputs(7253) <= (layer4_outputs(9622)) or (layer4_outputs(753));
    outputs(7254) <= layer4_outputs(1417);
    outputs(7255) <= (layer4_outputs(2882)) xor (layer4_outputs(8130));
    outputs(7256) <= (layer4_outputs(8168)) xor (layer4_outputs(3758));
    outputs(7257) <= not(layer4_outputs(7712));
    outputs(7258) <= layer4_outputs(3509);
    outputs(7259) <= not(layer4_outputs(7944));
    outputs(7260) <= not(layer4_outputs(2332));
    outputs(7261) <= not(layer4_outputs(5657));
    outputs(7262) <= layer4_outputs(3504);
    outputs(7263) <= not(layer4_outputs(5609));
    outputs(7264) <= not(layer4_outputs(9610));
    outputs(7265) <= not(layer4_outputs(7061)) or (layer4_outputs(3485));
    outputs(7266) <= (layer4_outputs(7521)) and (layer4_outputs(8118));
    outputs(7267) <= not(layer4_outputs(5172));
    outputs(7268) <= not(layer4_outputs(6397));
    outputs(7269) <= not(layer4_outputs(1706));
    outputs(7270) <= layer4_outputs(9658);
    outputs(7271) <= not((layer4_outputs(360)) xor (layer4_outputs(1719)));
    outputs(7272) <= not((layer4_outputs(5003)) xor (layer4_outputs(9967)));
    outputs(7273) <= not(layer4_outputs(8753));
    outputs(7274) <= layer4_outputs(3727);
    outputs(7275) <= layer4_outputs(7975);
    outputs(7276) <= (layer4_outputs(4025)) and not (layer4_outputs(1525));
    outputs(7277) <= layer4_outputs(9748);
    outputs(7278) <= (layer4_outputs(4470)) or (layer4_outputs(2641));
    outputs(7279) <= (layer4_outputs(5295)) xor (layer4_outputs(7462));
    outputs(7280) <= (layer4_outputs(7918)) xor (layer4_outputs(8262));
    outputs(7281) <= not(layer4_outputs(3921));
    outputs(7282) <= layer4_outputs(5957);
    outputs(7283) <= (layer4_outputs(4288)) xor (layer4_outputs(6216));
    outputs(7284) <= layer4_outputs(6132);
    outputs(7285) <= layer4_outputs(4370);
    outputs(7286) <= layer4_outputs(9404);
    outputs(7287) <= not(layer4_outputs(10081));
    outputs(7288) <= not((layer4_outputs(6269)) xor (layer4_outputs(10101)));
    outputs(7289) <= layer4_outputs(8049);
    outputs(7290) <= layer4_outputs(7054);
    outputs(7291) <= layer4_outputs(5386);
    outputs(7292) <= layer4_outputs(8535);
    outputs(7293) <= (layer4_outputs(3683)) and not (layer4_outputs(8011));
    outputs(7294) <= not(layer4_outputs(530));
    outputs(7295) <= (layer4_outputs(6083)) xor (layer4_outputs(2522));
    outputs(7296) <= layer4_outputs(8561);
    outputs(7297) <= not((layer4_outputs(4856)) xor (layer4_outputs(2079)));
    outputs(7298) <= not(layer4_outputs(5317));
    outputs(7299) <= layer4_outputs(9244);
    outputs(7300) <= not(layer4_outputs(9320));
    outputs(7301) <= layer4_outputs(9175);
    outputs(7302) <= not((layer4_outputs(8730)) and (layer4_outputs(3212)));
    outputs(7303) <= not((layer4_outputs(850)) xor (layer4_outputs(3919)));
    outputs(7304) <= not((layer4_outputs(5143)) xor (layer4_outputs(10059)));
    outputs(7305) <= (layer4_outputs(8676)) and not (layer4_outputs(7409));
    outputs(7306) <= not(layer4_outputs(6086));
    outputs(7307) <= not((layer4_outputs(7338)) or (layer4_outputs(2910)));
    outputs(7308) <= (layer4_outputs(1294)) and not (layer4_outputs(3685));
    outputs(7309) <= not(layer4_outputs(3365));
    outputs(7310) <= layer4_outputs(1289);
    outputs(7311) <= layer4_outputs(3960);
    outputs(7312) <= not(layer4_outputs(4334));
    outputs(7313) <= not((layer4_outputs(9877)) xor (layer4_outputs(2144)));
    outputs(7314) <= (layer4_outputs(9112)) and not (layer4_outputs(1408));
    outputs(7315) <= layer4_outputs(8751);
    outputs(7316) <= (layer4_outputs(1092)) xor (layer4_outputs(710));
    outputs(7317) <= not((layer4_outputs(3472)) xor (layer4_outputs(7258)));
    outputs(7318) <= not(layer4_outputs(3989));
    outputs(7319) <= not(layer4_outputs(3995));
    outputs(7320) <= (layer4_outputs(6082)) and (layer4_outputs(4424));
    outputs(7321) <= not(layer4_outputs(3986));
    outputs(7322) <= layer4_outputs(414);
    outputs(7323) <= layer4_outputs(5859);
    outputs(7324) <= layer4_outputs(477);
    outputs(7325) <= layer4_outputs(840);
    outputs(7326) <= not((layer4_outputs(4852)) xor (layer4_outputs(1662)));
    outputs(7327) <= not(layer4_outputs(196));
    outputs(7328) <= not(layer4_outputs(992));
    outputs(7329) <= layer4_outputs(4216);
    outputs(7330) <= not((layer4_outputs(3788)) or (layer4_outputs(4676)));
    outputs(7331) <= (layer4_outputs(8485)) xor (layer4_outputs(2989));
    outputs(7332) <= not(layer4_outputs(9422));
    outputs(7333) <= not(layer4_outputs(8097));
    outputs(7334) <= not((layer4_outputs(8966)) xor (layer4_outputs(7835)));
    outputs(7335) <= not((layer4_outputs(8702)) or (layer4_outputs(3517)));
    outputs(7336) <= not(layer4_outputs(5146));
    outputs(7337) <= layer4_outputs(1962);
    outputs(7338) <= not(layer4_outputs(1729));
    outputs(7339) <= (layer4_outputs(7414)) xor (layer4_outputs(5949));
    outputs(7340) <= layer4_outputs(8084);
    outputs(7341) <= not(layer4_outputs(6856));
    outputs(7342) <= not((layer4_outputs(7094)) xor (layer4_outputs(3136)));
    outputs(7343) <= not(layer4_outputs(10099));
    outputs(7344) <= not((layer4_outputs(1632)) or (layer4_outputs(628)));
    outputs(7345) <= (layer4_outputs(2724)) xor (layer4_outputs(2892));
    outputs(7346) <= (layer4_outputs(4189)) and not (layer4_outputs(7145));
    outputs(7347) <= layer4_outputs(4446);
    outputs(7348) <= layer4_outputs(8081);
    outputs(7349) <= not((layer4_outputs(7472)) xor (layer4_outputs(4933)));
    outputs(7350) <= (layer4_outputs(9616)) xor (layer4_outputs(8617));
    outputs(7351) <= not((layer4_outputs(10158)) xor (layer4_outputs(7518)));
    outputs(7352) <= layer4_outputs(3553);
    outputs(7353) <= not((layer4_outputs(670)) xor (layer4_outputs(9780)));
    outputs(7354) <= not(layer4_outputs(7309)) or (layer4_outputs(10134));
    outputs(7355) <= (layer4_outputs(2716)) xor (layer4_outputs(2849));
    outputs(7356) <= not(layer4_outputs(4597));
    outputs(7357) <= not((layer4_outputs(685)) xor (layer4_outputs(8775)));
    outputs(7358) <= layer4_outputs(7107);
    outputs(7359) <= (layer4_outputs(7893)) and not (layer4_outputs(6959));
    outputs(7360) <= not(layer4_outputs(4291));
    outputs(7361) <= not(layer4_outputs(5644));
    outputs(7362) <= not(layer4_outputs(3529));
    outputs(7363) <= layer4_outputs(5937);
    outputs(7364) <= not(layer4_outputs(1331));
    outputs(7365) <= not((layer4_outputs(4254)) or (layer4_outputs(6779)));
    outputs(7366) <= not(layer4_outputs(9377));
    outputs(7367) <= layer4_outputs(9193);
    outputs(7368) <= not((layer4_outputs(3575)) xor (layer4_outputs(9987)));
    outputs(7369) <= layer4_outputs(8322);
    outputs(7370) <= (layer4_outputs(1854)) xor (layer4_outputs(2266));
    outputs(7371) <= (layer4_outputs(2308)) xor (layer4_outputs(9520));
    outputs(7372) <= not(layer4_outputs(8778));
    outputs(7373) <= not(layer4_outputs(3318));
    outputs(7374) <= not(layer4_outputs(8008));
    outputs(7375) <= not(layer4_outputs(2658));
    outputs(7376) <= not(layer4_outputs(1412)) or (layer4_outputs(4816));
    outputs(7377) <= layer4_outputs(3791);
    outputs(7378) <= not(layer4_outputs(4871));
    outputs(7379) <= layer4_outputs(9811);
    outputs(7380) <= layer4_outputs(1116);
    outputs(7381) <= (layer4_outputs(6088)) xor (layer4_outputs(3234));
    outputs(7382) <= layer4_outputs(7584);
    outputs(7383) <= not((layer4_outputs(7715)) xor (layer4_outputs(2376)));
    outputs(7384) <= layer4_outputs(8078);
    outputs(7385) <= not((layer4_outputs(6105)) xor (layer4_outputs(3304)));
    outputs(7386) <= layer4_outputs(5691);
    outputs(7387) <= (layer4_outputs(3751)) and not (layer4_outputs(6533));
    outputs(7388) <= layer4_outputs(1792);
    outputs(7389) <= layer4_outputs(8809);
    outputs(7390) <= not(layer4_outputs(2299));
    outputs(7391) <= not((layer4_outputs(5548)) or (layer4_outputs(9526)));
    outputs(7392) <= layer4_outputs(9188);
    outputs(7393) <= not(layer4_outputs(8720));
    outputs(7394) <= layer4_outputs(5626);
    outputs(7395) <= not(layer4_outputs(399));
    outputs(7396) <= (layer4_outputs(5967)) xor (layer4_outputs(4019));
    outputs(7397) <= (layer4_outputs(751)) xor (layer4_outputs(9315));
    outputs(7398) <= not(layer4_outputs(4252));
    outputs(7399) <= layer4_outputs(4709);
    outputs(7400) <= layer4_outputs(3704);
    outputs(7401) <= layer4_outputs(7716);
    outputs(7402) <= not(layer4_outputs(1484));
    outputs(7403) <= layer4_outputs(1575);
    outputs(7404) <= layer4_outputs(9117);
    outputs(7405) <= not(layer4_outputs(9679));
    outputs(7406) <= not((layer4_outputs(616)) xor (layer4_outputs(5860)));
    outputs(7407) <= (layer4_outputs(3177)) and (layer4_outputs(9483));
    outputs(7408) <= layer4_outputs(7852);
    outputs(7409) <= layer4_outputs(1309);
    outputs(7410) <= layer4_outputs(4576);
    outputs(7411) <= not(layer4_outputs(5172));
    outputs(7412) <= not((layer4_outputs(7447)) xor (layer4_outputs(2351)));
    outputs(7413) <= layer4_outputs(3421);
    outputs(7414) <= layer4_outputs(4431);
    outputs(7415) <= not((layer4_outputs(4669)) xor (layer4_outputs(971)));
    outputs(7416) <= (layer4_outputs(4767)) xor (layer4_outputs(503));
    outputs(7417) <= not((layer4_outputs(3385)) or (layer4_outputs(1068)));
    outputs(7418) <= layer4_outputs(3071);
    outputs(7419) <= not(layer4_outputs(4789));
    outputs(7420) <= not(layer4_outputs(471));
    outputs(7421) <= not(layer4_outputs(7936));
    outputs(7422) <= (layer4_outputs(8356)) and not (layer4_outputs(8155));
    outputs(7423) <= not(layer4_outputs(6024));
    outputs(7424) <= not(layer4_outputs(2504));
    outputs(7425) <= layer4_outputs(3457);
    outputs(7426) <= not((layer4_outputs(230)) or (layer4_outputs(7429)));
    outputs(7427) <= (layer4_outputs(4472)) xor (layer4_outputs(476));
    outputs(7428) <= (layer4_outputs(2318)) and (layer4_outputs(9696));
    outputs(7429) <= not(layer4_outputs(9740));
    outputs(7430) <= not(layer4_outputs(6652)) or (layer4_outputs(5278));
    outputs(7431) <= not(layer4_outputs(6311));
    outputs(7432) <= layer4_outputs(2919);
    outputs(7433) <= not((layer4_outputs(1543)) xor (layer4_outputs(4369)));
    outputs(7434) <= (layer4_outputs(4426)) xor (layer4_outputs(1483));
    outputs(7435) <= not(layer4_outputs(1175));
    outputs(7436) <= (layer4_outputs(4761)) xor (layer4_outputs(221));
    outputs(7437) <= (layer4_outputs(329)) and (layer4_outputs(6357));
    outputs(7438) <= not(layer4_outputs(115));
    outputs(7439) <= not(layer4_outputs(1333)) or (layer4_outputs(2396));
    outputs(7440) <= layer4_outputs(6763);
    outputs(7441) <= not(layer4_outputs(9603));
    outputs(7442) <= not((layer4_outputs(603)) or (layer4_outputs(3142)));
    outputs(7443) <= not(layer4_outputs(8996));
    outputs(7444) <= not(layer4_outputs(9976)) or (layer4_outputs(2000));
    outputs(7445) <= layer4_outputs(7680);
    outputs(7446) <= layer4_outputs(2185);
    outputs(7447) <= layer4_outputs(7306);
    outputs(7448) <= (layer4_outputs(1830)) xor (layer4_outputs(9823));
    outputs(7449) <= layer4_outputs(6451);
    outputs(7450) <= layer4_outputs(9037);
    outputs(7451) <= layer4_outputs(8401);
    outputs(7452) <= not((layer4_outputs(654)) or (layer4_outputs(3218)));
    outputs(7453) <= (layer4_outputs(5183)) xor (layer4_outputs(5409));
    outputs(7454) <= (layer4_outputs(1841)) xor (layer4_outputs(1801));
    outputs(7455) <= not((layer4_outputs(9318)) xor (layer4_outputs(4342)));
    outputs(7456) <= layer4_outputs(1424);
    outputs(7457) <= (layer4_outputs(9750)) and (layer4_outputs(3502));
    outputs(7458) <= layer4_outputs(7974);
    outputs(7459) <= not(layer4_outputs(8299));
    outputs(7460) <= layer4_outputs(1710);
    outputs(7461) <= not((layer4_outputs(7508)) xor (layer4_outputs(8984)));
    outputs(7462) <= not(layer4_outputs(470));
    outputs(7463) <= not((layer4_outputs(2169)) xor (layer4_outputs(2089)));
    outputs(7464) <= (layer4_outputs(416)) xor (layer4_outputs(1389));
    outputs(7465) <= (layer4_outputs(5824)) xor (layer4_outputs(6365));
    outputs(7466) <= layer4_outputs(8787);
    outputs(7467) <= (layer4_outputs(6055)) and not (layer4_outputs(2809));
    outputs(7468) <= layer4_outputs(3324);
    outputs(7469) <= not((layer4_outputs(7367)) xor (layer4_outputs(2768)));
    outputs(7470) <= not((layer4_outputs(4244)) xor (layer4_outputs(1400)));
    outputs(7471) <= layer4_outputs(1494);
    outputs(7472) <= (layer4_outputs(9276)) xor (layer4_outputs(6145));
    outputs(7473) <= not(layer4_outputs(584));
    outputs(7474) <= (layer4_outputs(2964)) and (layer4_outputs(5880));
    outputs(7475) <= (layer4_outputs(2312)) and not (layer4_outputs(609));
    outputs(7476) <= layer4_outputs(2128);
    outputs(7477) <= not(layer4_outputs(3767));
    outputs(7478) <= layer4_outputs(6992);
    outputs(7479) <= layer4_outputs(4148);
    outputs(7480) <= layer4_outputs(5762);
    outputs(7481) <= layer4_outputs(7748);
    outputs(7482) <= not(layer4_outputs(4760));
    outputs(7483) <= not((layer4_outputs(10174)) xor (layer4_outputs(3761)));
    outputs(7484) <= layer4_outputs(3969);
    outputs(7485) <= (layer4_outputs(4832)) xor (layer4_outputs(6977));
    outputs(7486) <= not(layer4_outputs(8635)) or (layer4_outputs(1950));
    outputs(7487) <= not(layer4_outputs(98));
    outputs(7488) <= layer4_outputs(9901);
    outputs(7489) <= not(layer4_outputs(4037));
    outputs(7490) <= not(layer4_outputs(7271));
    outputs(7491) <= (layer4_outputs(1829)) and not (layer4_outputs(9139));
    outputs(7492) <= not((layer4_outputs(2068)) xor (layer4_outputs(6908)));
    outputs(7493) <= not((layer4_outputs(8524)) xor (layer4_outputs(5737)));
    outputs(7494) <= layer4_outputs(2018);
    outputs(7495) <= not(layer4_outputs(636));
    outputs(7496) <= (layer4_outputs(594)) and not (layer4_outputs(3609));
    outputs(7497) <= not((layer4_outputs(8858)) xor (layer4_outputs(2675)));
    outputs(7498) <= not((layer4_outputs(3207)) xor (layer4_outputs(1874)));
    outputs(7499) <= layer4_outputs(8381);
    outputs(7500) <= not(layer4_outputs(1936));
    outputs(7501) <= not(layer4_outputs(925));
    outputs(7502) <= (layer4_outputs(2841)) xor (layer4_outputs(2858));
    outputs(7503) <= not(layer4_outputs(7123));
    outputs(7504) <= not(layer4_outputs(8417));
    outputs(7505) <= not((layer4_outputs(10115)) or (layer4_outputs(6645)));
    outputs(7506) <= (layer4_outputs(10103)) xor (layer4_outputs(8696));
    outputs(7507) <= not((layer4_outputs(8861)) xor (layer4_outputs(9561)));
    outputs(7508) <= (layer4_outputs(4345)) and not (layer4_outputs(7771));
    outputs(7509) <= not((layer4_outputs(1013)) xor (layer4_outputs(8161)));
    outputs(7510) <= layer4_outputs(9461);
    outputs(7511) <= (layer4_outputs(1145)) or (layer4_outputs(6394));
    outputs(7512) <= (layer4_outputs(708)) xor (layer4_outputs(6434));
    outputs(7513) <= not(layer4_outputs(573));
    outputs(7514) <= not(layer4_outputs(1329));
    outputs(7515) <= (layer4_outputs(2383)) xor (layer4_outputs(1163));
    outputs(7516) <= not((layer4_outputs(9406)) xor (layer4_outputs(4595)));
    outputs(7517) <= layer4_outputs(1890);
    outputs(7518) <= layer4_outputs(6932);
    outputs(7519) <= layer4_outputs(3768);
    outputs(7520) <= (layer4_outputs(3846)) xor (layer4_outputs(4208));
    outputs(7521) <= (layer4_outputs(3084)) and not (layer4_outputs(882));
    outputs(7522) <= not(layer4_outputs(9495));
    outputs(7523) <= not(layer4_outputs(8908));
    outputs(7524) <= not((layer4_outputs(2737)) xor (layer4_outputs(5821)));
    outputs(7525) <= layer4_outputs(9972);
    outputs(7526) <= layer4_outputs(1756);
    outputs(7527) <= not(layer4_outputs(8248));
    outputs(7528) <= (layer4_outputs(6183)) and (layer4_outputs(8799));
    outputs(7529) <= (layer4_outputs(3743)) and not (layer4_outputs(8873));
    outputs(7530) <= (layer4_outputs(1574)) and not (layer4_outputs(3797));
    outputs(7531) <= not(layer4_outputs(9468));
    outputs(7532) <= (layer4_outputs(8899)) xor (layer4_outputs(4202));
    outputs(7533) <= layer4_outputs(5479);
    outputs(7534) <= not((layer4_outputs(5222)) xor (layer4_outputs(9588)));
    outputs(7535) <= (layer4_outputs(2075)) xor (layer4_outputs(3080));
    outputs(7536) <= layer4_outputs(5234);
    outputs(7537) <= not((layer4_outputs(8459)) xor (layer4_outputs(5456)));
    outputs(7538) <= (layer4_outputs(8914)) xor (layer4_outputs(8997));
    outputs(7539) <= not(layer4_outputs(1587)) or (layer4_outputs(4517));
    outputs(7540) <= not((layer4_outputs(9557)) xor (layer4_outputs(7956)));
    outputs(7541) <= (layer4_outputs(2997)) and not (layer4_outputs(7938));
    outputs(7542) <= not((layer4_outputs(994)) xor (layer4_outputs(9671)));
    outputs(7543) <= not(layer4_outputs(6885));
    outputs(7544) <= not((layer4_outputs(7881)) xor (layer4_outputs(4634)));
    outputs(7545) <= not((layer4_outputs(8651)) or (layer4_outputs(7139)));
    outputs(7546) <= (layer4_outputs(1745)) xor (layer4_outputs(2941));
    outputs(7547) <= not((layer4_outputs(1925)) xor (layer4_outputs(9339)));
    outputs(7548) <= not(layer4_outputs(9325));
    outputs(7549) <= not(layer4_outputs(4211));
    outputs(7550) <= layer4_outputs(5525);
    outputs(7551) <= (layer4_outputs(5039)) xor (layer4_outputs(3281));
    outputs(7552) <= not(layer4_outputs(7758));
    outputs(7553) <= (layer4_outputs(100)) and not (layer4_outputs(4195));
    outputs(7554) <= layer4_outputs(3499);
    outputs(7555) <= layer4_outputs(2944);
    outputs(7556) <= not((layer4_outputs(3303)) or (layer4_outputs(6494)));
    outputs(7557) <= not(layer4_outputs(5377));
    outputs(7558) <= not((layer4_outputs(6405)) xor (layer4_outputs(3989)));
    outputs(7559) <= '0';
    outputs(7560) <= layer4_outputs(4945);
    outputs(7561) <= not((layer4_outputs(9518)) xor (layer4_outputs(8351)));
    outputs(7562) <= layer4_outputs(3157);
    outputs(7563) <= not(layer4_outputs(9213));
    outputs(7564) <= not((layer4_outputs(8424)) xor (layer4_outputs(6472)));
    outputs(7565) <= layer4_outputs(246);
    outputs(7566) <= not((layer4_outputs(2843)) xor (layer4_outputs(2752)));
    outputs(7567) <= (layer4_outputs(152)) xor (layer4_outputs(688));
    outputs(7568) <= layer4_outputs(4279);
    outputs(7569) <= (layer4_outputs(554)) xor (layer4_outputs(10232));
    outputs(7570) <= layer4_outputs(4151);
    outputs(7571) <= layer4_outputs(7803);
    outputs(7572) <= not(layer4_outputs(6845));
    outputs(7573) <= not(layer4_outputs(4970));
    outputs(7574) <= not((layer4_outputs(4884)) xor (layer4_outputs(10065)));
    outputs(7575) <= not(layer4_outputs(577)) or (layer4_outputs(1323));
    outputs(7576) <= (layer4_outputs(3435)) and (layer4_outputs(6034));
    outputs(7577) <= (layer4_outputs(9926)) and not (layer4_outputs(6244));
    outputs(7578) <= layer4_outputs(2356);
    outputs(7579) <= (layer4_outputs(668)) and (layer4_outputs(4854));
    outputs(7580) <= not(layer4_outputs(191));
    outputs(7581) <= layer4_outputs(9102);
    outputs(7582) <= layer4_outputs(5526);
    outputs(7583) <= not((layer4_outputs(8145)) xor (layer4_outputs(7950)));
    outputs(7584) <= not((layer4_outputs(2115)) xor (layer4_outputs(2837)));
    outputs(7585) <= not(layer4_outputs(5307));
    outputs(7586) <= layer4_outputs(95);
    outputs(7587) <= (layer4_outputs(8507)) and not (layer4_outputs(1019));
    outputs(7588) <= not(layer4_outputs(2444));
    outputs(7589) <= not((layer4_outputs(5652)) xor (layer4_outputs(6126)));
    outputs(7590) <= layer4_outputs(9893);
    outputs(7591) <= not(layer4_outputs(180));
    outputs(7592) <= layer4_outputs(10112);
    outputs(7593) <= not((layer4_outputs(1647)) and (layer4_outputs(8018)));
    outputs(7594) <= not(layer4_outputs(5033));
    outputs(7595) <= not(layer4_outputs(1514));
    outputs(7596) <= not(layer4_outputs(6778));
    outputs(7597) <= (layer4_outputs(1240)) xor (layer4_outputs(3068));
    outputs(7598) <= layer4_outputs(7629);
    outputs(7599) <= layer4_outputs(757);
    outputs(7600) <= layer4_outputs(9647);
    outputs(7601) <= layer4_outputs(4417);
    outputs(7602) <= not((layer4_outputs(4902)) xor (layer4_outputs(8042)));
    outputs(7603) <= (layer4_outputs(10021)) xor (layer4_outputs(726));
    outputs(7604) <= layer4_outputs(9554);
    outputs(7605) <= layer4_outputs(8693);
    outputs(7606) <= (layer4_outputs(2195)) and not (layer4_outputs(2806));
    outputs(7607) <= layer4_outputs(1930);
    outputs(7608) <= layer4_outputs(259);
    outputs(7609) <= (layer4_outputs(6728)) and (layer4_outputs(5042));
    outputs(7610) <= (layer4_outputs(4301)) xor (layer4_outputs(6967));
    outputs(7611) <= layer4_outputs(3924);
    outputs(7612) <= layer4_outputs(2499);
    outputs(7613) <= layer4_outputs(75);
    outputs(7614) <= not(layer4_outputs(3048));
    outputs(7615) <= not(layer4_outputs(2821));
    outputs(7616) <= layer4_outputs(7902);
    outputs(7617) <= (layer4_outputs(7964)) xor (layer4_outputs(1753));
    outputs(7618) <= (layer4_outputs(9464)) xor (layer4_outputs(8621));
    outputs(7619) <= (layer4_outputs(5854)) xor (layer4_outputs(7176));
    outputs(7620) <= layer4_outputs(3565);
    outputs(7621) <= layer4_outputs(3839);
    outputs(7622) <= layer4_outputs(9830);
    outputs(7623) <= not(layer4_outputs(6740));
    outputs(7624) <= not(layer4_outputs(3690));
    outputs(7625) <= not(layer4_outputs(755));
    outputs(7626) <= layer4_outputs(1672);
    outputs(7627) <= not(layer4_outputs(3250));
    outputs(7628) <= layer4_outputs(4407);
    outputs(7629) <= (layer4_outputs(1910)) xor (layer4_outputs(804));
    outputs(7630) <= (layer4_outputs(3051)) and not (layer4_outputs(360));
    outputs(7631) <= not(layer4_outputs(5151));
    outputs(7632) <= not(layer4_outputs(5057));
    outputs(7633) <= not((layer4_outputs(3846)) xor (layer4_outputs(7834)));
    outputs(7634) <= layer4_outputs(6830);
    outputs(7635) <= layer4_outputs(6512);
    outputs(7636) <= (layer4_outputs(6775)) xor (layer4_outputs(212));
    outputs(7637) <= layer4_outputs(4742);
    outputs(7638) <= not(layer4_outputs(2962));
    outputs(7639) <= layer4_outputs(3879);
    outputs(7640) <= layer4_outputs(3704);
    outputs(7641) <= not(layer4_outputs(9077));
    outputs(7642) <= not(layer4_outputs(8375));
    outputs(7643) <= layer4_outputs(8239);
    outputs(7644) <= (layer4_outputs(9591)) or (layer4_outputs(8912));
    outputs(7645) <= layer4_outputs(1992);
    outputs(7646) <= layer4_outputs(4437);
    outputs(7647) <= not(layer4_outputs(3172));
    outputs(7648) <= not(layer4_outputs(4954));
    outputs(7649) <= layer4_outputs(3765);
    outputs(7650) <= layer4_outputs(863);
    outputs(7651) <= not((layer4_outputs(8884)) xor (layer4_outputs(2029)));
    outputs(7652) <= (layer4_outputs(6482)) xor (layer4_outputs(5813));
    outputs(7653) <= (layer4_outputs(1404)) or (layer4_outputs(874));
    outputs(7654) <= not(layer4_outputs(5018));
    outputs(7655) <= (layer4_outputs(1377)) and not (layer4_outputs(1394));
    outputs(7656) <= layer4_outputs(6926);
    outputs(7657) <= (layer4_outputs(8052)) and not (layer4_outputs(60));
    outputs(7658) <= not(layer4_outputs(308));
    outputs(7659) <= not((layer4_outputs(2429)) xor (layer4_outputs(102)));
    outputs(7660) <= (layer4_outputs(3866)) xor (layer4_outputs(6976));
    outputs(7661) <= not(layer4_outputs(10210));
    outputs(7662) <= layer4_outputs(4616);
    outputs(7663) <= not((layer4_outputs(9530)) xor (layer4_outputs(4505)));
    outputs(7664) <= not(layer4_outputs(3524)) or (layer4_outputs(2989));
    outputs(7665) <= (layer4_outputs(9978)) and (layer4_outputs(8135));
    outputs(7666) <= not(layer4_outputs(3297));
    outputs(7667) <= (layer4_outputs(7529)) xor (layer4_outputs(5932));
    outputs(7668) <= layer4_outputs(1833);
    outputs(7669) <= not((layer4_outputs(1399)) xor (layer4_outputs(7692)));
    outputs(7670) <= layer4_outputs(7199);
    outputs(7671) <= not((layer4_outputs(7147)) or (layer4_outputs(8801)));
    outputs(7672) <= not((layer4_outputs(1010)) xor (layer4_outputs(958)));
    outputs(7673) <= not((layer4_outputs(6796)) xor (layer4_outputs(4949)));
    outputs(7674) <= not(layer4_outputs(4568));
    outputs(7675) <= layer4_outputs(3406);
    outputs(7676) <= not(layer4_outputs(7504));
    outputs(7677) <= layer4_outputs(2155);
    outputs(7678) <= not(layer4_outputs(6072));
    outputs(7679) <= not(layer4_outputs(7548)) or (layer4_outputs(5699));
    outputs(7680) <= (layer4_outputs(1403)) and (layer4_outputs(8358));
    outputs(7681) <= not(layer4_outputs(2793));
    outputs(7682) <= (layer4_outputs(7741)) and not (layer4_outputs(1978));
    outputs(7683) <= (layer4_outputs(2424)) xor (layer4_outputs(3969));
    outputs(7684) <= layer4_outputs(5382);
    outputs(7685) <= not((layer4_outputs(522)) and (layer4_outputs(851)));
    outputs(7686) <= not(layer4_outputs(1248));
    outputs(7687) <= not(layer4_outputs(822));
    outputs(7688) <= not(layer4_outputs(8692));
    outputs(7689) <= layer4_outputs(6349);
    outputs(7690) <= not(layer4_outputs(1125));
    outputs(7691) <= layer4_outputs(3650);
    outputs(7692) <= (layer4_outputs(2025)) and not (layer4_outputs(7734));
    outputs(7693) <= not(layer4_outputs(2794));
    outputs(7694) <= not(layer4_outputs(7402));
    outputs(7695) <= layer4_outputs(8603);
    outputs(7696) <= (layer4_outputs(8967)) xor (layer4_outputs(1878));
    outputs(7697) <= not(layer4_outputs(1432));
    outputs(7698) <= not((layer4_outputs(9817)) or (layer4_outputs(6947)));
    outputs(7699) <= not(layer4_outputs(948));
    outputs(7700) <= not((layer4_outputs(9282)) xor (layer4_outputs(602)));
    outputs(7701) <= (layer4_outputs(5868)) and not (layer4_outputs(1379));
    outputs(7702) <= (layer4_outputs(5111)) and (layer4_outputs(2656));
    outputs(7703) <= not((layer4_outputs(7984)) or (layer4_outputs(6039)));
    outputs(7704) <= not(layer4_outputs(3378));
    outputs(7705) <= not(layer4_outputs(6420));
    outputs(7706) <= not(layer4_outputs(3638));
    outputs(7707) <= layer4_outputs(367);
    outputs(7708) <= (layer4_outputs(993)) and (layer4_outputs(5770));
    outputs(7709) <= (layer4_outputs(8891)) xor (layer4_outputs(6109));
    outputs(7710) <= layer4_outputs(182);
    outputs(7711) <= layer4_outputs(7363);
    outputs(7712) <= (layer4_outputs(1068)) xor (layer4_outputs(10066));
    outputs(7713) <= not(layer4_outputs(3095));
    outputs(7714) <= layer4_outputs(10006);
    outputs(7715) <= (layer4_outputs(7035)) and (layer4_outputs(8708));
    outputs(7716) <= not(layer4_outputs(7730));
    outputs(7717) <= not(layer4_outputs(2));
    outputs(7718) <= layer4_outputs(8707);
    outputs(7719) <= not(layer4_outputs(4498));
    outputs(7720) <= layer4_outputs(3091);
    outputs(7721) <= (layer4_outputs(9879)) xor (layer4_outputs(7710));
    outputs(7722) <= layer4_outputs(1266);
    outputs(7723) <= not(layer4_outputs(3199));
    outputs(7724) <= not((layer4_outputs(5644)) xor (layer4_outputs(1540)));
    outputs(7725) <= layer4_outputs(460);
    outputs(7726) <= not(layer4_outputs(7470));
    outputs(7727) <= (layer4_outputs(4785)) and (layer4_outputs(6895));
    outputs(7728) <= not(layer4_outputs(9370));
    outputs(7729) <= not((layer4_outputs(5776)) xor (layer4_outputs(7877)));
    outputs(7730) <= (layer4_outputs(9079)) xor (layer4_outputs(1599));
    outputs(7731) <= layer4_outputs(7242);
    outputs(7732) <= layer4_outputs(4168);
    outputs(7733) <= layer4_outputs(6827);
    outputs(7734) <= layer4_outputs(3406);
    outputs(7735) <= not(layer4_outputs(8599));
    outputs(7736) <= (layer4_outputs(8377)) and (layer4_outputs(7910));
    outputs(7737) <= (layer4_outputs(5128)) and (layer4_outputs(8165));
    outputs(7738) <= layer4_outputs(2584);
    outputs(7739) <= (layer4_outputs(4080)) and not (layer4_outputs(3812));
    outputs(7740) <= not(layer4_outputs(5571));
    outputs(7741) <= not((layer4_outputs(2886)) xor (layer4_outputs(1250)));
    outputs(7742) <= not(layer4_outputs(10129));
    outputs(7743) <= (layer4_outputs(7785)) xor (layer4_outputs(10173));
    outputs(7744) <= not((layer4_outputs(5947)) xor (layer4_outputs(1466)));
    outputs(7745) <= layer4_outputs(8305);
    outputs(7746) <= layer4_outputs(9593);
    outputs(7747) <= not(layer4_outputs(5141));
    outputs(7748) <= not(layer4_outputs(6760));
    outputs(7749) <= not(layer4_outputs(9390));
    outputs(7750) <= layer4_outputs(911);
    outputs(7751) <= (layer4_outputs(8629)) xor (layer4_outputs(6365));
    outputs(7752) <= not(layer4_outputs(5914));
    outputs(7753) <= layer4_outputs(2122);
    outputs(7754) <= (layer4_outputs(1690)) and (layer4_outputs(1023));
    outputs(7755) <= not((layer4_outputs(5270)) xor (layer4_outputs(1708)));
    outputs(7756) <= not(layer4_outputs(2444));
    outputs(7757) <= not((layer4_outputs(4895)) xor (layer4_outputs(1725)));
    outputs(7758) <= layer4_outputs(883);
    outputs(7759) <= not(layer4_outputs(884));
    outputs(7760) <= (layer4_outputs(4447)) xor (layer4_outputs(4362));
    outputs(7761) <= (layer4_outputs(3811)) and not (layer4_outputs(3912));
    outputs(7762) <= not((layer4_outputs(5448)) or (layer4_outputs(5311)));
    outputs(7763) <= (layer4_outputs(3920)) xor (layer4_outputs(7290));
    outputs(7764) <= not(layer4_outputs(1942));
    outputs(7765) <= layer4_outputs(5254);
    outputs(7766) <= layer4_outputs(7767);
    outputs(7767) <= not(layer4_outputs(5245));
    outputs(7768) <= not((layer4_outputs(4256)) xor (layer4_outputs(8645)));
    outputs(7769) <= not(layer4_outputs(8929));
    outputs(7770) <= layer4_outputs(9324);
    outputs(7771) <= not(layer4_outputs(2074));
    outputs(7772) <= (layer4_outputs(3253)) and not (layer4_outputs(2433));
    outputs(7773) <= '0';
    outputs(7774) <= not(layer4_outputs(1944));
    outputs(7775) <= (layer4_outputs(8434)) xor (layer4_outputs(6941));
    outputs(7776) <= not(layer4_outputs(1329));
    outputs(7777) <= not((layer4_outputs(8678)) xor (layer4_outputs(2811)));
    outputs(7778) <= not((layer4_outputs(9305)) xor (layer4_outputs(6277)));
    outputs(7779) <= layer4_outputs(4162);
    outputs(7780) <= not((layer4_outputs(10164)) xor (layer4_outputs(5678)));
    outputs(7781) <= (layer4_outputs(5881)) xor (layer4_outputs(103));
    outputs(7782) <= (layer4_outputs(1926)) xor (layer4_outputs(8454));
    outputs(7783) <= (layer4_outputs(5439)) and not (layer4_outputs(9742));
    outputs(7784) <= layer4_outputs(5572);
    outputs(7785) <= not((layer4_outputs(2172)) or (layer4_outputs(266)));
    outputs(7786) <= (layer4_outputs(3166)) and not (layer4_outputs(9300));
    outputs(7787) <= not(layer4_outputs(6694));
    outputs(7788) <= not(layer4_outputs(4750)) or (layer4_outputs(6955));
    outputs(7789) <= layer4_outputs(9937);
    outputs(7790) <= layer4_outputs(6741);
    outputs(7791) <= (layer4_outputs(2350)) xor (layer4_outputs(6061));
    outputs(7792) <= not(layer4_outputs(9668));
    outputs(7793) <= layer4_outputs(3411);
    outputs(7794) <= (layer4_outputs(301)) xor (layer4_outputs(4889));
    outputs(7795) <= not((layer4_outputs(3530)) xor (layer4_outputs(7118)));
    outputs(7796) <= not(layer4_outputs(3110));
    outputs(7797) <= not(layer4_outputs(5730)) or (layer4_outputs(1630));
    outputs(7798) <= layer4_outputs(3597);
    outputs(7799) <= layer4_outputs(2309);
    outputs(7800) <= (layer4_outputs(2222)) xor (layer4_outputs(86));
    outputs(7801) <= not((layer4_outputs(4119)) xor (layer4_outputs(5055)));
    outputs(7802) <= not((layer4_outputs(6850)) xor (layer4_outputs(1355)));
    outputs(7803) <= (layer4_outputs(8843)) and not (layer4_outputs(2336));
    outputs(7804) <= not(layer4_outputs(7144));
    outputs(7805) <= not(layer4_outputs(7332));
    outputs(7806) <= (layer4_outputs(1690)) xor (layer4_outputs(5084));
    outputs(7807) <= layer4_outputs(9146);
    outputs(7808) <= not(layer4_outputs(6303));
    outputs(7809) <= not((layer4_outputs(8902)) xor (layer4_outputs(5110)));
    outputs(7810) <= (layer4_outputs(1406)) xor (layer4_outputs(2622));
    outputs(7811) <= layer4_outputs(6787);
    outputs(7812) <= not((layer4_outputs(4324)) xor (layer4_outputs(5340)));
    outputs(7813) <= not((layer4_outputs(10113)) xor (layer4_outputs(3618)));
    outputs(7814) <= (layer4_outputs(4359)) or (layer4_outputs(1723));
    outputs(7815) <= not(layer4_outputs(6509));
    outputs(7816) <= not(layer4_outputs(9564));
    outputs(7817) <= layer4_outputs(10172);
    outputs(7818) <= layer4_outputs(6890);
    outputs(7819) <= not(layer4_outputs(907));
    outputs(7820) <= not(layer4_outputs(2343));
    outputs(7821) <= not(layer4_outputs(6657));
    outputs(7822) <= layer4_outputs(9688);
    outputs(7823) <= not(layer4_outputs(5793));
    outputs(7824) <= (layer4_outputs(4873)) or (layer4_outputs(8790));
    outputs(7825) <= not((layer4_outputs(5081)) xor (layer4_outputs(5476)));
    outputs(7826) <= not(layer4_outputs(4793));
    outputs(7827) <= (layer4_outputs(9407)) and not (layer4_outputs(4333));
    outputs(7828) <= not((layer4_outputs(8925)) xor (layer4_outputs(8648)));
    outputs(7829) <= not(layer4_outputs(3333));
    outputs(7830) <= not(layer4_outputs(5481));
    outputs(7831) <= not(layer4_outputs(6551));
    outputs(7832) <= not(layer4_outputs(9603));
    outputs(7833) <= not(layer4_outputs(9782));
    outputs(7834) <= (layer4_outputs(478)) and (layer4_outputs(4897));
    outputs(7835) <= not(layer4_outputs(4965));
    outputs(7836) <= layer4_outputs(9208);
    outputs(7837) <= (layer4_outputs(8096)) and not (layer4_outputs(3720));
    outputs(7838) <= not(layer4_outputs(3223));
    outputs(7839) <= not(layer4_outputs(9776));
    outputs(7840) <= layer4_outputs(2702);
    outputs(7841) <= (layer4_outputs(2386)) and not (layer4_outputs(10220));
    outputs(7842) <= (layer4_outputs(698)) and (layer4_outputs(92));
    outputs(7843) <= (layer4_outputs(1379)) xor (layer4_outputs(9010));
    outputs(7844) <= (layer4_outputs(10114)) xor (layer4_outputs(856));
    outputs(7845) <= (layer4_outputs(4283)) and not (layer4_outputs(323));
    outputs(7846) <= (layer4_outputs(2687)) xor (layer4_outputs(9830));
    outputs(7847) <= not((layer4_outputs(9508)) or (layer4_outputs(9179)));
    outputs(7848) <= not(layer4_outputs(256));
    outputs(7849) <= layer4_outputs(6324);
    outputs(7850) <= (layer4_outputs(2047)) and (layer4_outputs(9948));
    outputs(7851) <= layer4_outputs(6452);
    outputs(7852) <= not((layer4_outputs(7193)) or (layer4_outputs(6039)));
    outputs(7853) <= not((layer4_outputs(9573)) xor (layer4_outputs(5698)));
    outputs(7854) <= not(layer4_outputs(564));
    outputs(7855) <= not(layer4_outputs(6395));
    outputs(7856) <= not(layer4_outputs(5988)) or (layer4_outputs(7669));
    outputs(7857) <= layer4_outputs(5787);
    outputs(7858) <= layer4_outputs(7943);
    outputs(7859) <= not(layer4_outputs(9643));
    outputs(7860) <= not(layer4_outputs(6096));
    outputs(7861) <= not(layer4_outputs(1306));
    outputs(7862) <= not(layer4_outputs(7239));
    outputs(7863) <= layer4_outputs(9251);
    outputs(7864) <= not(layer4_outputs(8758));
    outputs(7865) <= not((layer4_outputs(1509)) or (layer4_outputs(6440)));
    outputs(7866) <= not(layer4_outputs(6421));
    outputs(7867) <= not(layer4_outputs(8295));
    outputs(7868) <= not((layer4_outputs(10073)) xor (layer4_outputs(4767)));
    outputs(7869) <= not((layer4_outputs(2724)) and (layer4_outputs(8490)));
    outputs(7870) <= not(layer4_outputs(661));
    outputs(7871) <= not(layer4_outputs(3661));
    outputs(7872) <= layer4_outputs(10201);
    outputs(7873) <= not(layer4_outputs(7602));
    outputs(7874) <= (layer4_outputs(1832)) xor (layer4_outputs(5173));
    outputs(7875) <= not(layer4_outputs(180));
    outputs(7876) <= not(layer4_outputs(2750));
    outputs(7877) <= not(layer4_outputs(4553));
    outputs(7878) <= (layer4_outputs(494)) xor (layer4_outputs(298));
    outputs(7879) <= not((layer4_outputs(9209)) xor (layer4_outputs(9387)));
    outputs(7880) <= layer4_outputs(1378);
    outputs(7881) <= (layer4_outputs(1210)) and not (layer4_outputs(5379));
    outputs(7882) <= not((layer4_outputs(4612)) xor (layer4_outputs(2491)));
    outputs(7883) <= (layer4_outputs(2926)) xor (layer4_outputs(9594));
    outputs(7884) <= layer4_outputs(9533);
    outputs(7885) <= layer4_outputs(6408);
    outputs(7886) <= not(layer4_outputs(9023));
    outputs(7887) <= layer4_outputs(10142);
    outputs(7888) <= layer4_outputs(6133);
    outputs(7889) <= not(layer4_outputs(7028)) or (layer4_outputs(1930));
    outputs(7890) <= layer4_outputs(7633);
    outputs(7891) <= (layer4_outputs(206)) xor (layer4_outputs(10224));
    outputs(7892) <= layer4_outputs(4762);
    outputs(7893) <= (layer4_outputs(3159)) and not (layer4_outputs(964));
    outputs(7894) <= layer4_outputs(3585);
    outputs(7895) <= layer4_outputs(4805);
    outputs(7896) <= not(layer4_outputs(5746));
    outputs(7897) <= not(layer4_outputs(1017));
    outputs(7898) <= not(layer4_outputs(1469));
    outputs(7899) <= layer4_outputs(4071);
    outputs(7900) <= layer4_outputs(7002);
    outputs(7901) <= (layer4_outputs(7549)) xor (layer4_outputs(6945));
    outputs(7902) <= not(layer4_outputs(4178)) or (layer4_outputs(2108));
    outputs(7903) <= not(layer4_outputs(4547));
    outputs(7904) <= not(layer4_outputs(3897));
    outputs(7905) <= layer4_outputs(2442);
    outputs(7906) <= (layer4_outputs(5614)) xor (layer4_outputs(3245));
    outputs(7907) <= not(layer4_outputs(2538));
    outputs(7908) <= (layer4_outputs(9764)) and (layer4_outputs(1898));
    outputs(7909) <= layer4_outputs(4192);
    outputs(7910) <= not((layer4_outputs(2020)) xor (layer4_outputs(6935)));
    outputs(7911) <= layer4_outputs(10175);
    outputs(7912) <= not((layer4_outputs(6078)) xor (layer4_outputs(9362)));
    outputs(7913) <= not(layer4_outputs(8828));
    outputs(7914) <= not((layer4_outputs(6032)) or (layer4_outputs(5407)));
    outputs(7915) <= not(layer4_outputs(6996));
    outputs(7916) <= (layer4_outputs(5355)) and not (layer4_outputs(211));
    outputs(7917) <= (layer4_outputs(7529)) xor (layer4_outputs(1782));
    outputs(7918) <= not(layer4_outputs(1967));
    outputs(7919) <= not(layer4_outputs(257));
    outputs(7920) <= layer4_outputs(5579);
    outputs(7921) <= (layer4_outputs(827)) and (layer4_outputs(7096));
    outputs(7922) <= not((layer4_outputs(3825)) xor (layer4_outputs(7067)));
    outputs(7923) <= not(layer4_outputs(9400));
    outputs(7924) <= not(layer4_outputs(2349));
    outputs(7925) <= '1';
    outputs(7926) <= layer4_outputs(6707);
    outputs(7927) <= not(layer4_outputs(3941));
    outputs(7928) <= layer4_outputs(8883);
    outputs(7929) <= (layer4_outputs(7014)) xor (layer4_outputs(3851));
    outputs(7930) <= not((layer4_outputs(4632)) or (layer4_outputs(6958)));
    outputs(7931) <= not(layer4_outputs(7508));
    outputs(7932) <= layer4_outputs(10163);
    outputs(7933) <= layer4_outputs(1764);
    outputs(7934) <= layer4_outputs(1579);
    outputs(7935) <= not(layer4_outputs(9047));
    outputs(7936) <= (layer4_outputs(6642)) and (layer4_outputs(6128));
    outputs(7937) <= not((layer4_outputs(5548)) or (layer4_outputs(5394)));
    outputs(7938) <= (layer4_outputs(8525)) xor (layer4_outputs(2131));
    outputs(7939) <= (layer4_outputs(7948)) or (layer4_outputs(9896));
    outputs(7940) <= not((layer4_outputs(9788)) xor (layer4_outputs(1593)));
    outputs(7941) <= (layer4_outputs(5723)) xor (layer4_outputs(2308));
    outputs(7942) <= layer4_outputs(1910);
    outputs(7943) <= not((layer4_outputs(7652)) xor (layer4_outputs(8624)));
    outputs(7944) <= not(layer4_outputs(3120));
    outputs(7945) <= layer4_outputs(9566);
    outputs(7946) <= not((layer4_outputs(4177)) xor (layer4_outputs(2331)));
    outputs(7947) <= not((layer4_outputs(1371)) xor (layer4_outputs(5037)));
    outputs(7948) <= layer4_outputs(5932);
    outputs(7949) <= layer4_outputs(2958);
    outputs(7950) <= not((layer4_outputs(9990)) xor (layer4_outputs(5839)));
    outputs(7951) <= (layer4_outputs(848)) xor (layer4_outputs(9791));
    outputs(7952) <= layer4_outputs(6387);
    outputs(7953) <= not(layer4_outputs(7678));
    outputs(7954) <= layer4_outputs(490);
    outputs(7955) <= layer4_outputs(7523);
    outputs(7956) <= not(layer4_outputs(4885));
    outputs(7957) <= not(layer4_outputs(6597));
    outputs(7958) <= layer4_outputs(8588);
    outputs(7959) <= not(layer4_outputs(4991));
    outputs(7960) <= (layer4_outputs(3632)) and not (layer4_outputs(8420));
    outputs(7961) <= layer4_outputs(6030);
    outputs(7962) <= not(layer4_outputs(8536));
    outputs(7963) <= not(layer4_outputs(3246));
    outputs(7964) <= layer4_outputs(3146);
    outputs(7965) <= not(layer4_outputs(1017));
    outputs(7966) <= not(layer4_outputs(3383));
    outputs(7967) <= not(layer4_outputs(7123));
    outputs(7968) <= not((layer4_outputs(52)) xor (layer4_outputs(8913)));
    outputs(7969) <= not(layer4_outputs(1306));
    outputs(7970) <= layer4_outputs(76);
    outputs(7971) <= layer4_outputs(1207);
    outputs(7972) <= not((layer4_outputs(6979)) xor (layer4_outputs(548)));
    outputs(7973) <= layer4_outputs(5312);
    outputs(7974) <= not(layer4_outputs(9055));
    outputs(7975) <= layer4_outputs(10091);
    outputs(7976) <= layer4_outputs(3607);
    outputs(7977) <= (layer4_outputs(5900)) and (layer4_outputs(7416));
    outputs(7978) <= not((layer4_outputs(9401)) and (layer4_outputs(2139)));
    outputs(7979) <= (layer4_outputs(1430)) xor (layer4_outputs(571));
    outputs(7980) <= layer4_outputs(4690);
    outputs(7981) <= not(layer4_outputs(6676));
    outputs(7982) <= (layer4_outputs(7646)) xor (layer4_outputs(4379));
    outputs(7983) <= not(layer4_outputs(5007));
    outputs(7984) <= layer4_outputs(8096);
    outputs(7985) <= layer4_outputs(3166);
    outputs(7986) <= (layer4_outputs(7218)) and (layer4_outputs(89));
    outputs(7987) <= (layer4_outputs(5546)) and (layer4_outputs(640));
    outputs(7988) <= not(layer4_outputs(1781));
    outputs(7989) <= layer4_outputs(2885);
    outputs(7990) <= layer4_outputs(3243);
    outputs(7991) <= layer4_outputs(1116);
    outputs(7992) <= (layer4_outputs(480)) xor (layer4_outputs(1476));
    outputs(7993) <= layer4_outputs(5425);
    outputs(7994) <= not(layer4_outputs(5645));
    outputs(7995) <= (layer4_outputs(5942)) and not (layer4_outputs(4306));
    outputs(7996) <= not((layer4_outputs(7804)) or (layer4_outputs(164)));
    outputs(7997) <= (layer4_outputs(2404)) xor (layer4_outputs(985));
    outputs(7998) <= layer4_outputs(7951);
    outputs(7999) <= not(layer4_outputs(3432));
    outputs(8000) <= (layer4_outputs(5080)) xor (layer4_outputs(3771));
    outputs(8001) <= (layer4_outputs(3450)) xor (layer4_outputs(8580));
    outputs(8002) <= layer4_outputs(3670);
    outputs(8003) <= layer4_outputs(2061);
    outputs(8004) <= not(layer4_outputs(3805));
    outputs(8005) <= not((layer4_outputs(1921)) xor (layer4_outputs(1202)));
    outputs(8006) <= layer4_outputs(3762);
    outputs(8007) <= not((layer4_outputs(6226)) xor (layer4_outputs(6643)));
    outputs(8008) <= (layer4_outputs(8271)) xor (layer4_outputs(1990));
    outputs(8009) <= layer4_outputs(5490);
    outputs(8010) <= not((layer4_outputs(998)) xor (layer4_outputs(8934)));
    outputs(8011) <= not(layer4_outputs(4281));
    outputs(8012) <= not(layer4_outputs(1038));
    outputs(8013) <= not(layer4_outputs(240));
    outputs(8014) <= not((layer4_outputs(1498)) xor (layer4_outputs(4152)));
    outputs(8015) <= (layer4_outputs(6686)) and (layer4_outputs(3361));
    outputs(8016) <= not((layer4_outputs(4819)) or (layer4_outputs(8445)));
    outputs(8017) <= not(layer4_outputs(9493));
    outputs(8018) <= layer4_outputs(6339);
    outputs(8019) <= not((layer4_outputs(2718)) xor (layer4_outputs(7413)));
    outputs(8020) <= not(layer4_outputs(5297));
    outputs(8021) <= not(layer4_outputs(5598));
    outputs(8022) <= not(layer4_outputs(6103));
    outputs(8023) <= not(layer4_outputs(6031));
    outputs(8024) <= not(layer4_outputs(3256));
    outputs(8025) <= not(layer4_outputs(3035));
    outputs(8026) <= not(layer4_outputs(4288));
    outputs(8027) <= not(layer4_outputs(5809));
    outputs(8028) <= layer4_outputs(9252);
    outputs(8029) <= (layer4_outputs(4182)) or (layer4_outputs(6834));
    outputs(8030) <= not(layer4_outputs(6254));
    outputs(8031) <= (layer4_outputs(1321)) and not (layer4_outputs(6861));
    outputs(8032) <= layer4_outputs(5167);
    outputs(8033) <= layer4_outputs(1804);
    outputs(8034) <= (layer4_outputs(2180)) xor (layer4_outputs(10001));
    outputs(8035) <= layer4_outputs(8683);
    outputs(8036) <= not((layer4_outputs(621)) xor (layer4_outputs(2714)));
    outputs(8037) <= layer4_outputs(8469);
    outputs(8038) <= not((layer4_outputs(1049)) xor (layer4_outputs(6285)));
    outputs(8039) <= layer4_outputs(1744);
    outputs(8040) <= not(layer4_outputs(4871));
    outputs(8041) <= (layer4_outputs(4399)) and not (layer4_outputs(1788));
    outputs(8042) <= not((layer4_outputs(495)) xor (layer4_outputs(3096)));
    outputs(8043) <= (layer4_outputs(7157)) and not (layer4_outputs(2103));
    outputs(8044) <= (layer4_outputs(4661)) xor (layer4_outputs(1761));
    outputs(8045) <= not(layer4_outputs(656));
    outputs(8046) <= not((layer4_outputs(8465)) xor (layer4_outputs(3596)));
    outputs(8047) <= layer4_outputs(7390);
    outputs(8048) <= not(layer4_outputs(1160));
    outputs(8049) <= not(layer4_outputs(1407));
    outputs(8050) <= not((layer4_outputs(543)) xor (layer4_outputs(3547)));
    outputs(8051) <= not((layer4_outputs(2718)) xor (layer4_outputs(4366)));
    outputs(8052) <= (layer4_outputs(2812)) xor (layer4_outputs(817));
    outputs(8053) <= layer4_outputs(690);
    outputs(8054) <= not(layer4_outputs(7178));
    outputs(8055) <= layer4_outputs(8774);
    outputs(8056) <= (layer4_outputs(907)) xor (layer4_outputs(588));
    outputs(8057) <= (layer4_outputs(2636)) or (layer4_outputs(9298));
    outputs(8058) <= not(layer4_outputs(6736));
    outputs(8059) <= not(layer4_outputs(7697));
    outputs(8060) <= layer4_outputs(2356);
    outputs(8061) <= not(layer4_outputs(701));
    outputs(8062) <= (layer4_outputs(8746)) xor (layer4_outputs(1008));
    outputs(8063) <= layer4_outputs(2719);
    outputs(8064) <= not(layer4_outputs(655));
    outputs(8065) <= layer4_outputs(556);
    outputs(8066) <= layer4_outputs(1262);
    outputs(8067) <= not((layer4_outputs(2860)) xor (layer4_outputs(2037)));
    outputs(8068) <= layer4_outputs(1305);
    outputs(8069) <= layer4_outputs(7593);
    outputs(8070) <= not(layer4_outputs(8846));
    outputs(8071) <= not(layer4_outputs(2817));
    outputs(8072) <= not(layer4_outputs(497)) or (layer4_outputs(6056));
    outputs(8073) <= layer4_outputs(1653);
    outputs(8074) <= not(layer4_outputs(1259));
    outputs(8075) <= (layer4_outputs(4497)) and not (layer4_outputs(857));
    outputs(8076) <= (layer4_outputs(5879)) xor (layer4_outputs(9288));
    outputs(8077) <= not(layer4_outputs(4797));
    outputs(8078) <= not(layer4_outputs(9424));
    outputs(8079) <= not(layer4_outputs(3931));
    outputs(8080) <= (layer4_outputs(8920)) and (layer4_outputs(3819));
    outputs(8081) <= not(layer4_outputs(6373));
    outputs(8082) <= (layer4_outputs(119)) xor (layer4_outputs(1229));
    outputs(8083) <= not(layer4_outputs(4643));
    outputs(8084) <= not((layer4_outputs(2646)) and (layer4_outputs(5070)));
    outputs(8085) <= layer4_outputs(4686);
    outputs(8086) <= not(layer4_outputs(1913));
    outputs(8087) <= layer4_outputs(2555);
    outputs(8088) <= layer4_outputs(657);
    outputs(8089) <= (layer4_outputs(7585)) or (layer4_outputs(5652));
    outputs(8090) <= not((layer4_outputs(5779)) or (layer4_outputs(4633)));
    outputs(8091) <= not((layer4_outputs(7380)) xor (layer4_outputs(5716)));
    outputs(8092) <= (layer4_outputs(4800)) and (layer4_outputs(10074));
    outputs(8093) <= not((layer4_outputs(7094)) xor (layer4_outputs(1221)));
    outputs(8094) <= not(layer4_outputs(8452));
    outputs(8095) <= not((layer4_outputs(10186)) xor (layer4_outputs(5101)));
    outputs(8096) <= not((layer4_outputs(5961)) xor (layer4_outputs(3874)));
    outputs(8097) <= layer4_outputs(3435);
    outputs(8098) <= not(layer4_outputs(373));
    outputs(8099) <= (layer4_outputs(7798)) and (layer4_outputs(2669));
    outputs(8100) <= (layer4_outputs(2365)) and not (layer4_outputs(3814));
    outputs(8101) <= not(layer4_outputs(7116));
    outputs(8102) <= not(layer4_outputs(375));
    outputs(8103) <= not((layer4_outputs(10216)) xor (layer4_outputs(5170)));
    outputs(8104) <= not((layer4_outputs(2484)) xor (layer4_outputs(5451)));
    outputs(8105) <= not(layer4_outputs(5909));
    outputs(8106) <= not(layer4_outputs(2743));
    outputs(8107) <= layer4_outputs(1900);
    outputs(8108) <= not((layer4_outputs(7043)) xor (layer4_outputs(9190)));
    outputs(8109) <= not((layer4_outputs(8516)) xor (layer4_outputs(2170)));
    outputs(8110) <= not((layer4_outputs(1681)) xor (layer4_outputs(9591)));
    outputs(8111) <= not((layer4_outputs(4811)) and (layer4_outputs(3402)));
    outputs(8112) <= layer4_outputs(3307);
    outputs(8113) <= not((layer4_outputs(4323)) xor (layer4_outputs(7760)));
    outputs(8114) <= layer4_outputs(6441);
    outputs(8115) <= not(layer4_outputs(4763));
    outputs(8116) <= not(layer4_outputs(8906));
    outputs(8117) <= layer4_outputs(1620);
    outputs(8118) <= layer4_outputs(620);
    outputs(8119) <= layer4_outputs(2428);
    outputs(8120) <= not(layer4_outputs(1917));
    outputs(8121) <= not(layer4_outputs(3620));
    outputs(8122) <= not((layer4_outputs(6179)) xor (layer4_outputs(8209)));
    outputs(8123) <= not(layer4_outputs(3773));
    outputs(8124) <= (layer4_outputs(253)) xor (layer4_outputs(7033));
    outputs(8125) <= layer4_outputs(6763);
    outputs(8126) <= not(layer4_outputs(6206));
    outputs(8127) <= not(layer4_outputs(9239));
    outputs(8128) <= layer4_outputs(7298);
    outputs(8129) <= not(layer4_outputs(1978));
    outputs(8130) <= not(layer4_outputs(3776));
    outputs(8131) <= (layer4_outputs(9337)) or (layer4_outputs(6674));
    outputs(8132) <= not(layer4_outputs(407));
    outputs(8133) <= layer4_outputs(8328);
    outputs(8134) <= layer4_outputs(1731);
    outputs(8135) <= not(layer4_outputs(9348));
    outputs(8136) <= not(layer4_outputs(5143));
    outputs(8137) <= (layer4_outputs(7165)) xor (layer4_outputs(7667));
    outputs(8138) <= layer4_outputs(2480);
    outputs(8139) <= not(layer4_outputs(3383));
    outputs(8140) <= not(layer4_outputs(9734));
    outputs(8141) <= not(layer4_outputs(10154));
    outputs(8142) <= layer4_outputs(26);
    outputs(8143) <= (layer4_outputs(1226)) xor (layer4_outputs(1131));
    outputs(8144) <= not(layer4_outputs(3286));
    outputs(8145) <= (layer4_outputs(5915)) and (layer4_outputs(4404));
    outputs(8146) <= not(layer4_outputs(6208));
    outputs(8147) <= '0';
    outputs(8148) <= (layer4_outputs(5020)) or (layer4_outputs(8648));
    outputs(8149) <= (layer4_outputs(9441)) xor (layer4_outputs(3629));
    outputs(8150) <= not(layer4_outputs(8887)) or (layer4_outputs(1168));
    outputs(8151) <= layer4_outputs(1345);
    outputs(8152) <= not(layer4_outputs(6878));
    outputs(8153) <= not(layer4_outputs(8752));
    outputs(8154) <= (layer4_outputs(1129)) xor (layer4_outputs(597));
    outputs(8155) <= layer4_outputs(1107);
    outputs(8156) <= not(layer4_outputs(482));
    outputs(8157) <= not(layer4_outputs(7474));
    outputs(8158) <= layer4_outputs(4577);
    outputs(8159) <= layer4_outputs(8681);
    outputs(8160) <= not(layer4_outputs(9714));
    outputs(8161) <= (layer4_outputs(5636)) and (layer4_outputs(1133));
    outputs(8162) <= layer4_outputs(6000);
    outputs(8163) <= layer4_outputs(6832);
    outputs(8164) <= not(layer4_outputs(5929));
    outputs(8165) <= layer4_outputs(6272);
    outputs(8166) <= not(layer4_outputs(7542));
    outputs(8167) <= (layer4_outputs(7345)) or (layer4_outputs(5227));
    outputs(8168) <= not(layer4_outputs(6636));
    outputs(8169) <= not(layer4_outputs(4394));
    outputs(8170) <= (layer4_outputs(5071)) xor (layer4_outputs(3315));
    outputs(8171) <= (layer4_outputs(5926)) and not (layer4_outputs(418));
    outputs(8172) <= layer4_outputs(5301);
    outputs(8173) <= layer4_outputs(4717);
    outputs(8174) <= (layer4_outputs(662)) and (layer4_outputs(5792));
    outputs(8175) <= (layer4_outputs(8621)) xor (layer4_outputs(2907));
    outputs(8176) <= not((layer4_outputs(8215)) xor (layer4_outputs(5197)));
    outputs(8177) <= layer4_outputs(2736);
    outputs(8178) <= (layer4_outputs(2085)) xor (layer4_outputs(2343));
    outputs(8179) <= layer4_outputs(6049);
    outputs(8180) <= layer4_outputs(5329);
    outputs(8181) <= not(layer4_outputs(2545));
    outputs(8182) <= layer4_outputs(9251);
    outputs(8183) <= (layer4_outputs(9893)) and (layer4_outputs(10037));
    outputs(8184) <= layer4_outputs(7262);
    outputs(8185) <= (layer4_outputs(5828)) and not (layer4_outputs(7870));
    outputs(8186) <= not(layer4_outputs(9398));
    outputs(8187) <= not(layer4_outputs(7232));
    outputs(8188) <= not((layer4_outputs(1533)) xor (layer4_outputs(7286)));
    outputs(8189) <= not(layer4_outputs(5091));
    outputs(8190) <= not((layer4_outputs(10009)) xor (layer4_outputs(4390)));
    outputs(8191) <= not(layer4_outputs(5226));
    outputs(8192) <= (layer4_outputs(8757)) xor (layer4_outputs(1654));
    outputs(8193) <= not((layer4_outputs(10124)) or (layer4_outputs(4064)));
    outputs(8194) <= not(layer4_outputs(6321)) or (layer4_outputs(1592));
    outputs(8195) <= not(layer4_outputs(1234));
    outputs(8196) <= layer4_outputs(9066);
    outputs(8197) <= layer4_outputs(8553);
    outputs(8198) <= layer4_outputs(6750);
    outputs(8199) <= (layer4_outputs(3163)) xor (layer4_outputs(6975));
    outputs(8200) <= layer4_outputs(8851);
    outputs(8201) <= (layer4_outputs(738)) or (layer4_outputs(8667));
    outputs(8202) <= not(layer4_outputs(6184));
    outputs(8203) <= (layer4_outputs(4381)) xor (layer4_outputs(723));
    outputs(8204) <= (layer4_outputs(8957)) xor (layer4_outputs(6824));
    outputs(8205) <= (layer4_outputs(664)) xor (layer4_outputs(6729));
    outputs(8206) <= (layer4_outputs(5248)) xor (layer4_outputs(5917));
    outputs(8207) <= not((layer4_outputs(3831)) xor (layer4_outputs(7354)));
    outputs(8208) <= not((layer4_outputs(2015)) xor (layer4_outputs(4166)));
    outputs(8209) <= (layer4_outputs(145)) xor (layer4_outputs(6754));
    outputs(8210) <= (layer4_outputs(3024)) and (layer4_outputs(2416));
    outputs(8211) <= not(layer4_outputs(4920)) or (layer4_outputs(6160));
    outputs(8212) <= (layer4_outputs(1435)) xor (layer4_outputs(8783));
    outputs(8213) <= layer4_outputs(436);
    outputs(8214) <= not(layer4_outputs(7282)) or (layer4_outputs(6688));
    outputs(8215) <= (layer4_outputs(395)) xor (layer4_outputs(9617));
    outputs(8216) <= layer4_outputs(4418);
    outputs(8217) <= not((layer4_outputs(8714)) xor (layer4_outputs(4211)));
    outputs(8218) <= layer4_outputs(5051);
    outputs(8219) <= layer4_outputs(6116);
    outputs(8220) <= not((layer4_outputs(132)) xor (layer4_outputs(4505)));
    outputs(8221) <= not(layer4_outputs(9481));
    outputs(8222) <= layer4_outputs(5863);
    outputs(8223) <= not(layer4_outputs(9916));
    outputs(8224) <= layer4_outputs(6584);
    outputs(8225) <= layer4_outputs(474);
    outputs(8226) <= not((layer4_outputs(276)) xor (layer4_outputs(6977)));
    outputs(8227) <= layer4_outputs(3732);
    outputs(8228) <= not(layer4_outputs(7997));
    outputs(8229) <= not(layer4_outputs(508));
    outputs(8230) <= not(layer4_outputs(9813));
    outputs(8231) <= not(layer4_outputs(350)) or (layer4_outputs(5991));
    outputs(8232) <= layer4_outputs(2591);
    outputs(8233) <= not(layer4_outputs(1973));
    outputs(8234) <= (layer4_outputs(3992)) and not (layer4_outputs(5668));
    outputs(8235) <= not(layer4_outputs(3459));
    outputs(8236) <= layer4_outputs(6307);
    outputs(8237) <= layer4_outputs(5998);
    outputs(8238) <= not((layer4_outputs(5670)) xor (layer4_outputs(3005)));
    outputs(8239) <= layer4_outputs(9332);
    outputs(8240) <= layer4_outputs(5607);
    outputs(8241) <= not((layer4_outputs(4377)) xor (layer4_outputs(8867)));
    outputs(8242) <= (layer4_outputs(2328)) xor (layer4_outputs(4150));
    outputs(8243) <= not(layer4_outputs(2302));
    outputs(8244) <= not(layer4_outputs(6934));
    outputs(8245) <= not(layer4_outputs(4559)) or (layer4_outputs(5279));
    outputs(8246) <= not(layer4_outputs(605));
    outputs(8247) <= not(layer4_outputs(7978));
    outputs(8248) <= not(layer4_outputs(5008)) or (layer4_outputs(8779));
    outputs(8249) <= not((layer4_outputs(9586)) and (layer4_outputs(8893)));
    outputs(8250) <= (layer4_outputs(3617)) xor (layer4_outputs(7085));
    outputs(8251) <= not(layer4_outputs(409));
    outputs(8252) <= layer4_outputs(9630);
    outputs(8253) <= (layer4_outputs(724)) or (layer4_outputs(7063));
    outputs(8254) <= not((layer4_outputs(1299)) xor (layer4_outputs(5073)));
    outputs(8255) <= layer4_outputs(8492);
    outputs(8256) <= layer4_outputs(3580);
    outputs(8257) <= not((layer4_outputs(6523)) xor (layer4_outputs(4191)));
    outputs(8258) <= not(layer4_outputs(7620));
    outputs(8259) <= not((layer4_outputs(8617)) xor (layer4_outputs(8148)));
    outputs(8260) <= not(layer4_outputs(2225));
    outputs(8261) <= not((layer4_outputs(2379)) xor (layer4_outputs(6017)));
    outputs(8262) <= not(layer4_outputs(9959)) or (layer4_outputs(4689));
    outputs(8263) <= not(layer4_outputs(8793));
    outputs(8264) <= (layer4_outputs(2001)) xor (layer4_outputs(6708));
    outputs(8265) <= layer4_outputs(3800);
    outputs(8266) <= not((layer4_outputs(542)) xor (layer4_outputs(2466)));
    outputs(8267) <= layer4_outputs(2182);
    outputs(8268) <= layer4_outputs(5432);
    outputs(8269) <= not(layer4_outputs(7095)) or (layer4_outputs(1444));
    outputs(8270) <= not(layer4_outputs(5979));
    outputs(8271) <= not((layer4_outputs(10105)) xor (layer4_outputs(6735)));
    outputs(8272) <= not(layer4_outputs(8965));
    outputs(8273) <= not(layer4_outputs(3279)) or (layer4_outputs(9932));
    outputs(8274) <= layer4_outputs(9507);
    outputs(8275) <= (layer4_outputs(4133)) and (layer4_outputs(5300));
    outputs(8276) <= (layer4_outputs(8504)) and (layer4_outputs(4904));
    outputs(8277) <= not(layer4_outputs(2490));
    outputs(8278) <= not(layer4_outputs(2523));
    outputs(8279) <= layer4_outputs(1286);
    outputs(8280) <= not(layer4_outputs(6645));
    outputs(8281) <= (layer4_outputs(5970)) xor (layer4_outputs(7366));
    outputs(8282) <= not(layer4_outputs(4831));
    outputs(8283) <= not(layer4_outputs(9362));
    outputs(8284) <= not(layer4_outputs(4138));
    outputs(8285) <= layer4_outputs(1420);
    outputs(8286) <= not(layer4_outputs(6368));
    outputs(8287) <= (layer4_outputs(3894)) or (layer4_outputs(10207));
    outputs(8288) <= (layer4_outputs(2117)) or (layer4_outputs(5130));
    outputs(8289) <= not((layer4_outputs(646)) xor (layer4_outputs(4020)));
    outputs(8290) <= layer4_outputs(968);
    outputs(8291) <= layer4_outputs(6151);
    outputs(8292) <= not(layer4_outputs(4798)) or (layer4_outputs(7031));
    outputs(8293) <= layer4_outputs(5148);
    outputs(8294) <= '1';
    outputs(8295) <= layer4_outputs(1840);
    outputs(8296) <= not(layer4_outputs(3736)) or (layer4_outputs(4244));
    outputs(8297) <= layer4_outputs(2006);
    outputs(8298) <= not(layer4_outputs(7657)) or (layer4_outputs(9607));
    outputs(8299) <= layer4_outputs(6463);
    outputs(8300) <= layer4_outputs(2842);
    outputs(8301) <= not((layer4_outputs(5086)) or (layer4_outputs(4261)));
    outputs(8302) <= (layer4_outputs(6221)) xor (layer4_outputs(9387));
    outputs(8303) <= not((layer4_outputs(9917)) and (layer4_outputs(8823)));
    outputs(8304) <= layer4_outputs(2083);
    outputs(8305) <= layer4_outputs(3225);
    outputs(8306) <= not(layer4_outputs(4920));
    outputs(8307) <= (layer4_outputs(7846)) xor (layer4_outputs(2003));
    outputs(8308) <= layer4_outputs(5903);
    outputs(8309) <= (layer4_outputs(1914)) and not (layer4_outputs(7276));
    outputs(8310) <= layer4_outputs(9983);
    outputs(8311) <= not(layer4_outputs(6155));
    outputs(8312) <= not(layer4_outputs(6338));
    outputs(8313) <= not(layer4_outputs(1715));
    outputs(8314) <= (layer4_outputs(642)) xor (layer4_outputs(8765));
    outputs(8315) <= layer4_outputs(1091);
    outputs(8316) <= layer4_outputs(764);
    outputs(8317) <= (layer4_outputs(6186)) or (layer4_outputs(2876));
    outputs(8318) <= layer4_outputs(62);
    outputs(8319) <= not((layer4_outputs(9922)) xor (layer4_outputs(4116)));
    outputs(8320) <= not((layer4_outputs(2848)) xor (layer4_outputs(2846)));
    outputs(8321) <= layer4_outputs(6783);
    outputs(8322) <= not(layer4_outputs(3974));
    outputs(8323) <= layer4_outputs(8950);
    outputs(8324) <= not(layer4_outputs(2069));
    outputs(8325) <= layer4_outputs(5435);
    outputs(8326) <= not((layer4_outputs(2489)) xor (layer4_outputs(335)));
    outputs(8327) <= (layer4_outputs(291)) or (layer4_outputs(7640));
    outputs(8328) <= not(layer4_outputs(3924)) or (layer4_outputs(5631));
    outputs(8329) <= not(layer4_outputs(676)) or (layer4_outputs(8378));
    outputs(8330) <= not(layer4_outputs(205)) or (layer4_outputs(8053));
    outputs(8331) <= not(layer4_outputs(1067));
    outputs(8332) <= '0';
    outputs(8333) <= not((layer4_outputs(861)) xor (layer4_outputs(5173)));
    outputs(8334) <= layer4_outputs(9836);
    outputs(8335) <= layer4_outputs(6423);
    outputs(8336) <= not((layer4_outputs(6061)) and (layer4_outputs(9415)));
    outputs(8337) <= (layer4_outputs(1373)) xor (layer4_outputs(8512));
    outputs(8338) <= not(layer4_outputs(9859));
    outputs(8339) <= not(layer4_outputs(9342)) or (layer4_outputs(8134));
    outputs(8340) <= layer4_outputs(6083);
    outputs(8341) <= (layer4_outputs(7514)) xor (layer4_outputs(6917));
    outputs(8342) <= not((layer4_outputs(3626)) xor (layer4_outputs(1402)));
    outputs(8343) <= layer4_outputs(5214);
    outputs(8344) <= layer4_outputs(2050);
    outputs(8345) <= (layer4_outputs(3938)) xor (layer4_outputs(5190));
    outputs(8346) <= (layer4_outputs(2844)) and (layer4_outputs(1101));
    outputs(8347) <= not((layer4_outputs(879)) xor (layer4_outputs(7172)));
    outputs(8348) <= layer4_outputs(5268);
    outputs(8349) <= not((layer4_outputs(256)) xor (layer4_outputs(123)));
    outputs(8350) <= layer4_outputs(6164);
    outputs(8351) <= not(layer4_outputs(8815));
    outputs(8352) <= not(layer4_outputs(6799));
    outputs(8353) <= not((layer4_outputs(8943)) xor (layer4_outputs(6209)));
    outputs(8354) <= layer4_outputs(2668);
    outputs(8355) <= (layer4_outputs(1544)) or (layer4_outputs(8697));
    outputs(8356) <= not(layer4_outputs(3189));
    outputs(8357) <= (layer4_outputs(4635)) and (layer4_outputs(8178));
    outputs(8358) <= not((layer4_outputs(9912)) xor (layer4_outputs(8183)));
    outputs(8359) <= layer4_outputs(9294);
    outputs(8360) <= layer4_outputs(6243);
    outputs(8361) <= not(layer4_outputs(4744));
    outputs(8362) <= not(layer4_outputs(5189));
    outputs(8363) <= layer4_outputs(5075);
    outputs(8364) <= layer4_outputs(3558);
    outputs(8365) <= not(layer4_outputs(2751));
    outputs(8366) <= layer4_outputs(2798);
    outputs(8367) <= (layer4_outputs(5339)) xor (layer4_outputs(9220));
    outputs(8368) <= not((layer4_outputs(289)) and (layer4_outputs(7822)));
    outputs(8369) <= (layer4_outputs(5869)) and (layer4_outputs(6485));
    outputs(8370) <= (layer4_outputs(9862)) or (layer4_outputs(4384));
    outputs(8371) <= not(layer4_outputs(6707));
    outputs(8372) <= (layer4_outputs(4638)) and (layer4_outputs(3731));
    outputs(8373) <= (layer4_outputs(9303)) xor (layer4_outputs(9780));
    outputs(8374) <= layer4_outputs(5442);
    outputs(8375) <= layer4_outputs(1179);
    outputs(8376) <= not(layer4_outputs(8635)) or (layer4_outputs(461));
    outputs(8377) <= layer4_outputs(8044);
    outputs(8378) <= layer4_outputs(3030);
    outputs(8379) <= layer4_outputs(7114);
    outputs(8380) <= layer4_outputs(1818);
    outputs(8381) <= (layer4_outputs(1956)) and not (layer4_outputs(9829));
    outputs(8382) <= (layer4_outputs(4135)) xor (layer4_outputs(614));
    outputs(8383) <= not(layer4_outputs(1742));
    outputs(8384) <= (layer4_outputs(3638)) and not (layer4_outputs(455));
    outputs(8385) <= not(layer4_outputs(3616)) or (layer4_outputs(1410));
    outputs(8386) <= not(layer4_outputs(66));
    outputs(8387) <= not(layer4_outputs(1005));
    outputs(8388) <= not(layer4_outputs(4761)) or (layer4_outputs(5066));
    outputs(8389) <= not((layer4_outputs(6170)) or (layer4_outputs(8407)));
    outputs(8390) <= not((layer4_outputs(1998)) or (layer4_outputs(9115)));
    outputs(8391) <= not(layer4_outputs(2987));
    outputs(8392) <= not((layer4_outputs(8356)) and (layer4_outputs(3543)));
    outputs(8393) <= not(layer4_outputs(2808));
    outputs(8394) <= not(layer4_outputs(8357)) or (layer4_outputs(8903));
    outputs(8395) <= layer4_outputs(8705);
    outputs(8396) <= layer4_outputs(1595);
    outputs(8397) <= '0';
    outputs(8398) <= (layer4_outputs(5203)) xor (layer4_outputs(3771));
    outputs(8399) <= (layer4_outputs(4806)) xor (layer4_outputs(10090));
    outputs(8400) <= not(layer4_outputs(6248));
    outputs(8401) <= not(layer4_outputs(6112));
    outputs(8402) <= layer4_outputs(2214);
    outputs(8403) <= layer4_outputs(1997);
    outputs(8404) <= not((layer4_outputs(1359)) xor (layer4_outputs(9214)));
    outputs(8405) <= not(layer4_outputs(450));
    outputs(8406) <= not(layer4_outputs(4743));
    outputs(8407) <= layer4_outputs(2683);
    outputs(8408) <= not(layer4_outputs(7917));
    outputs(8409) <= not(layer4_outputs(9107)) or (layer4_outputs(2903));
    outputs(8410) <= (layer4_outputs(5911)) xor (layer4_outputs(798));
    outputs(8411) <= (layer4_outputs(5416)) xor (layer4_outputs(6106));
    outputs(8412) <= not(layer4_outputs(3120));
    outputs(8413) <= layer4_outputs(2066);
    outputs(8414) <= layer4_outputs(5990);
    outputs(8415) <= not(layer4_outputs(7142));
    outputs(8416) <= '0';
    outputs(8417) <= not(layer4_outputs(8080));
    outputs(8418) <= (layer4_outputs(9204)) xor (layer4_outputs(6614));
    outputs(8419) <= not((layer4_outputs(6853)) and (layer4_outputs(1607)));
    outputs(8420) <= not(layer4_outputs(6354));
    outputs(8421) <= (layer4_outputs(2074)) and not (layer4_outputs(7140));
    outputs(8422) <= layer4_outputs(35);
    outputs(8423) <= not((layer4_outputs(3802)) and (layer4_outputs(684)));
    outputs(8424) <= not(layer4_outputs(9105));
    outputs(8425) <= not(layer4_outputs(7330));
    outputs(8426) <= layer4_outputs(8186);
    outputs(8427) <= layer4_outputs(7942);
    outputs(8428) <= not((layer4_outputs(6199)) xor (layer4_outputs(10213)));
    outputs(8429) <= not(layer4_outputs(9929)) or (layer4_outputs(7356));
    outputs(8430) <= layer4_outputs(5974);
    outputs(8431) <= not((layer4_outputs(2075)) or (layer4_outputs(9464)));
    outputs(8432) <= layer4_outputs(7681);
    outputs(8433) <= not(layer4_outputs(4699));
    outputs(8434) <= not(layer4_outputs(2510));
    outputs(8435) <= layer4_outputs(1332);
    outputs(8436) <= (layer4_outputs(3907)) xor (layer4_outputs(892));
    outputs(8437) <= not(layer4_outputs(8322));
    outputs(8438) <= (layer4_outputs(188)) or (layer4_outputs(2722));
    outputs(8439) <= (layer4_outputs(5680)) xor (layer4_outputs(7551));
    outputs(8440) <= (layer4_outputs(1700)) xor (layer4_outputs(3045));
    outputs(8441) <= (layer4_outputs(10096)) and (layer4_outputs(6801));
    outputs(8442) <= (layer4_outputs(4389)) or (layer4_outputs(5084));
    outputs(8443) <= layer4_outputs(6208);
    outputs(8444) <= (layer4_outputs(10118)) xor (layer4_outputs(8256));
    outputs(8445) <= not((layer4_outputs(6851)) and (layer4_outputs(9357)));
    outputs(8446) <= layer4_outputs(1965);
    outputs(8447) <= not(layer4_outputs(8906)) or (layer4_outputs(678));
    outputs(8448) <= not((layer4_outputs(9882)) xor (layer4_outputs(4954)));
    outputs(8449) <= (layer4_outputs(3117)) or (layer4_outputs(8932));
    outputs(8450) <= not(layer4_outputs(5252));
    outputs(8451) <= layer4_outputs(3255);
    outputs(8452) <= (layer4_outputs(8886)) xor (layer4_outputs(1543));
    outputs(8453) <= (layer4_outputs(3605)) xor (layer4_outputs(4828));
    outputs(8454) <= not((layer4_outputs(5759)) xor (layer4_outputs(4088)));
    outputs(8455) <= not(layer4_outputs(3299));
    outputs(8456) <= layer4_outputs(8206);
    outputs(8457) <= not(layer4_outputs(7619));
    outputs(8458) <= not((layer4_outputs(10213)) xor (layer4_outputs(7816)));
    outputs(8459) <= layer4_outputs(5427);
    outputs(8460) <= not((layer4_outputs(6816)) and (layer4_outputs(9843)));
    outputs(8461) <= not(layer4_outputs(9785));
    outputs(8462) <= (layer4_outputs(9544)) xor (layer4_outputs(4008));
    outputs(8463) <= layer4_outputs(2725);
    outputs(8464) <= not((layer4_outputs(6092)) and (layer4_outputs(525)));
    outputs(8465) <= (layer4_outputs(2758)) xor (layer4_outputs(8487));
    outputs(8466) <= not(layer4_outputs(2889));
    outputs(8467) <= layer4_outputs(4793);
    outputs(8468) <= not((layer4_outputs(1096)) and (layer4_outputs(4014)));
    outputs(8469) <= layer4_outputs(3881);
    outputs(8470) <= not(layer4_outputs(5739));
    outputs(8471) <= (layer4_outputs(9358)) xor (layer4_outputs(1196));
    outputs(8472) <= layer4_outputs(6215);
    outputs(8473) <= layer4_outputs(9170);
    outputs(8474) <= not(layer4_outputs(6023)) or (layer4_outputs(4513));
    outputs(8475) <= not(layer4_outputs(1894));
    outputs(8476) <= layer4_outputs(62);
    outputs(8477) <= layer4_outputs(3108);
    outputs(8478) <= not(layer4_outputs(6987));
    outputs(8479) <= (layer4_outputs(5285)) xor (layer4_outputs(232));
    outputs(8480) <= not(layer4_outputs(5609));
    outputs(8481) <= not((layer4_outputs(9226)) xor (layer4_outputs(5043)));
    outputs(8482) <= layer4_outputs(5429);
    outputs(8483) <= not(layer4_outputs(8836));
    outputs(8484) <= not((layer4_outputs(4077)) xor (layer4_outputs(5216)));
    outputs(8485) <= layer4_outputs(7325);
    outputs(8486) <= layer4_outputs(9536);
    outputs(8487) <= layer4_outputs(3512);
    outputs(8488) <= not((layer4_outputs(2582)) and (layer4_outputs(9427)));
    outputs(8489) <= layer4_outputs(7271);
    outputs(8490) <= layer4_outputs(6682);
    outputs(8491) <= not((layer4_outputs(8613)) xor (layer4_outputs(9642)));
    outputs(8492) <= layer4_outputs(2498);
    outputs(8493) <= not((layer4_outputs(3854)) and (layer4_outputs(730)));
    outputs(8494) <= layer4_outputs(5219);
    outputs(8495) <= not(layer4_outputs(766));
    outputs(8496) <= layer4_outputs(8769);
    outputs(8497) <= not((layer4_outputs(1215)) xor (layer4_outputs(2330)));
    outputs(8498) <= (layer4_outputs(4356)) or (layer4_outputs(4248));
    outputs(8499) <= not((layer4_outputs(7828)) xor (layer4_outputs(4233)));
    outputs(8500) <= layer4_outputs(3291);
    outputs(8501) <= layer4_outputs(7278);
    outputs(8502) <= layer4_outputs(5278);
    outputs(8503) <= not(layer4_outputs(9994));
    outputs(8504) <= (layer4_outputs(6315)) and not (layer4_outputs(2540));
    outputs(8505) <= not((layer4_outputs(536)) xor (layer4_outputs(6953)));
    outputs(8506) <= layer4_outputs(1150);
    outputs(8507) <= layer4_outputs(2843);
    outputs(8508) <= not((layer4_outputs(6185)) xor (layer4_outputs(1136)));
    outputs(8509) <= layer4_outputs(4842);
    outputs(8510) <= not(layer4_outputs(2647));
    outputs(8511) <= layer4_outputs(7219);
    outputs(8512) <= not(layer4_outputs(568));
    outputs(8513) <= layer4_outputs(1245);
    outputs(8514) <= (layer4_outputs(4795)) and not (layer4_outputs(8320));
    outputs(8515) <= not(layer4_outputs(2500)) or (layer4_outputs(1053));
    outputs(8516) <= not(layer4_outputs(8318));
    outputs(8517) <= not(layer4_outputs(876));
    outputs(8518) <= not(layer4_outputs(4698));
    outputs(8519) <= not(layer4_outputs(2004));
    outputs(8520) <= not(layer4_outputs(4843));
    outputs(8521) <= not(layer4_outputs(861));
    outputs(8522) <= (layer4_outputs(3420)) xor (layer4_outputs(5569));
    outputs(8523) <= layer4_outputs(1665);
    outputs(8524) <= (layer4_outputs(6432)) and not (layer4_outputs(3942));
    outputs(8525) <= (layer4_outputs(4187)) or (layer4_outputs(8245));
    outputs(8526) <= not(layer4_outputs(899));
    outputs(8527) <= layer4_outputs(6638);
    outputs(8528) <= layer4_outputs(4017);
    outputs(8529) <= not(layer4_outputs(6310));
    outputs(8530) <= not(layer4_outputs(2004));
    outputs(8531) <= (layer4_outputs(4074)) xor (layer4_outputs(7847));
    outputs(8532) <= (layer4_outputs(3133)) or (layer4_outputs(6595));
    outputs(8533) <= not((layer4_outputs(4606)) xor (layer4_outputs(532)));
    outputs(8534) <= layer4_outputs(4498);
    outputs(8535) <= not((layer4_outputs(9813)) and (layer4_outputs(7627)));
    outputs(8536) <= (layer4_outputs(619)) xor (layer4_outputs(2279));
    outputs(8537) <= (layer4_outputs(3893)) and not (layer4_outputs(5083));
    outputs(8538) <= not(layer4_outputs(487));
    outputs(8539) <= (layer4_outputs(2574)) and not (layer4_outputs(4157));
    outputs(8540) <= layer4_outputs(5816);
    outputs(8541) <= not((layer4_outputs(5345)) xor (layer4_outputs(1062)));
    outputs(8542) <= not((layer4_outputs(2785)) xor (layer4_outputs(10160)));
    outputs(8543) <= (layer4_outputs(3680)) or (layer4_outputs(6015));
    outputs(8544) <= not(layer4_outputs(7358));
    outputs(8545) <= (layer4_outputs(7849)) or (layer4_outputs(1998));
    outputs(8546) <= layer4_outputs(8338);
    outputs(8547) <= layer4_outputs(9277);
    outputs(8548) <= layer4_outputs(5755);
    outputs(8549) <= (layer4_outputs(8169)) xor (layer4_outputs(6453));
    outputs(8550) <= not(layer4_outputs(4751));
    outputs(8551) <= not((layer4_outputs(2118)) xor (layer4_outputs(1071)));
    outputs(8552) <= not((layer4_outputs(117)) xor (layer4_outputs(4105)));
    outputs(8553) <= not(layer4_outputs(8784));
    outputs(8554) <= not((layer4_outputs(4640)) xor (layer4_outputs(1113)));
    outputs(8555) <= not((layer4_outputs(6918)) xor (layer4_outputs(9439)));
    outputs(8556) <= not(layer4_outputs(6806)) or (layer4_outputs(8481));
    outputs(8557) <= (layer4_outputs(9053)) xor (layer4_outputs(7526));
    outputs(8558) <= layer4_outputs(10169);
    outputs(8559) <= layer4_outputs(7026);
    outputs(8560) <= (layer4_outputs(4260)) or (layer4_outputs(1918));
    outputs(8561) <= not(layer4_outputs(3272)) or (layer4_outputs(2231));
    outputs(8562) <= layer4_outputs(8284);
    outputs(8563) <= layer4_outputs(7538);
    outputs(8564) <= layer4_outputs(1101);
    outputs(8565) <= not(layer4_outputs(6350));
    outputs(8566) <= (layer4_outputs(1987)) xor (layer4_outputs(3899));
    outputs(8567) <= layer4_outputs(4155);
    outputs(8568) <= layer4_outputs(7122);
    outputs(8569) <= not((layer4_outputs(4327)) or (layer4_outputs(9484)));
    outputs(8570) <= layer4_outputs(1245);
    outputs(8571) <= not(layer4_outputs(1309));
    outputs(8572) <= not(layer4_outputs(3374));
    outputs(8573) <= not(layer4_outputs(5129)) or (layer4_outputs(4269));
    outputs(8574) <= layer4_outputs(6524);
    outputs(8575) <= layer4_outputs(5967);
    outputs(8576) <= not(layer4_outputs(1005));
    outputs(8577) <= (layer4_outputs(6587)) xor (layer4_outputs(133));
    outputs(8578) <= not((layer4_outputs(7839)) xor (layer4_outputs(2208)));
    outputs(8579) <= layer4_outputs(8772);
    outputs(8580) <= (layer4_outputs(5379)) or (layer4_outputs(2272));
    outputs(8581) <= not(layer4_outputs(4157));
    outputs(8582) <= not((layer4_outputs(1472)) and (layer4_outputs(9918)));
    outputs(8583) <= not(layer4_outputs(3773)) or (layer4_outputs(8733));
    outputs(8584) <= not((layer4_outputs(340)) xor (layer4_outputs(5815)));
    outputs(8585) <= layer4_outputs(4474);
    outputs(8586) <= not(layer4_outputs(8552)) or (layer4_outputs(9075));
    outputs(8587) <= not((layer4_outputs(7411)) xor (layer4_outputs(2206)));
    outputs(8588) <= not(layer4_outputs(6230));
    outputs(8589) <= not(layer4_outputs(5625));
    outputs(8590) <= not(layer4_outputs(5893));
    outputs(8591) <= not((layer4_outputs(4417)) xor (layer4_outputs(1410)));
    outputs(8592) <= not(layer4_outputs(2754));
    outputs(8593) <= layer4_outputs(2006);
    outputs(8594) <= (layer4_outputs(6785)) and (layer4_outputs(10040));
    outputs(8595) <= not((layer4_outputs(1880)) xor (layer4_outputs(8331)));
    outputs(8596) <= not(layer4_outputs(7763));
    outputs(8597) <= layer4_outputs(5178);
    outputs(8598) <= not((layer4_outputs(8518)) xor (layer4_outputs(4320)));
    outputs(8599) <= layer4_outputs(2101);
    outputs(8600) <= not(layer4_outputs(3675));
    outputs(8601) <= not(layer4_outputs(5433)) or (layer4_outputs(7027));
    outputs(8602) <= layer4_outputs(1955);
    outputs(8603) <= not(layer4_outputs(4841));
    outputs(8604) <= not(layer4_outputs(7002));
    outputs(8605) <= not((layer4_outputs(7634)) xor (layer4_outputs(5647)));
    outputs(8606) <= layer4_outputs(961);
    outputs(8607) <= (layer4_outputs(4865)) xor (layer4_outputs(1445));
    outputs(8608) <= layer4_outputs(1827);
    outputs(8609) <= layer4_outputs(9063);
    outputs(8610) <= layer4_outputs(6245);
    outputs(8611) <= not(layer4_outputs(281));
    outputs(8612) <= not(layer4_outputs(2227)) or (layer4_outputs(2394));
    outputs(8613) <= (layer4_outputs(3784)) xor (layer4_outputs(7595));
    outputs(8614) <= not((layer4_outputs(8975)) xor (layer4_outputs(7112)));
    outputs(8615) <= layer4_outputs(9380);
    outputs(8616) <= not(layer4_outputs(7864));
    outputs(8617) <= not(layer4_outputs(6973));
    outputs(8618) <= not((layer4_outputs(4081)) xor (layer4_outputs(672)));
    outputs(8619) <= layer4_outputs(5630);
    outputs(8620) <= layer4_outputs(1859);
    outputs(8621) <= not(layer4_outputs(6300));
    outputs(8622) <= layer4_outputs(2251);
    outputs(8623) <= not((layer4_outputs(767)) or (layer4_outputs(10155)));
    outputs(8624) <= not((layer4_outputs(4808)) xor (layer4_outputs(5934)));
    outputs(8625) <= layer4_outputs(2445);
    outputs(8626) <= not(layer4_outputs(9475));
    outputs(8627) <= (layer4_outputs(8382)) xor (layer4_outputs(1988));
    outputs(8628) <= (layer4_outputs(9363)) xor (layer4_outputs(9364));
    outputs(8629) <= layer4_outputs(8766);
    outputs(8630) <= layer4_outputs(6474);
    outputs(8631) <= not(layer4_outputs(4836)) or (layer4_outputs(5898));
    outputs(8632) <= not(layer4_outputs(4201));
    outputs(8633) <= not(layer4_outputs(1056));
    outputs(8634) <= not(layer4_outputs(5530));
    outputs(8635) <= not(layer4_outputs(8494));
    outputs(8636) <= layer4_outputs(2745);
    outputs(8637) <= not(layer4_outputs(8725)) or (layer4_outputs(854));
    outputs(8638) <= not(layer4_outputs(3539));
    outputs(8639) <= not(layer4_outputs(5627));
    outputs(8640) <= layer4_outputs(5667);
    outputs(8641) <= not(layer4_outputs(9861)) or (layer4_outputs(2451));
    outputs(8642) <= (layer4_outputs(1483)) xor (layer4_outputs(9135));
    outputs(8643) <= not(layer4_outputs(4690));
    outputs(8644) <= (layer4_outputs(7190)) xor (layer4_outputs(7745));
    outputs(8645) <= not((layer4_outputs(7933)) or (layer4_outputs(9075)));
    outputs(8646) <= layer4_outputs(4464);
    outputs(8647) <= not(layer4_outputs(9087));
    outputs(8648) <= not(layer4_outputs(1518));
    outputs(8649) <= (layer4_outputs(2678)) xor (layer4_outputs(3982));
    outputs(8650) <= not(layer4_outputs(844));
    outputs(8651) <= layer4_outputs(5293);
    outputs(8652) <= (layer4_outputs(8088)) or (layer4_outputs(3564));
    outputs(8653) <= layer4_outputs(10058);
    outputs(8654) <= layer4_outputs(2675);
    outputs(8655) <= layer4_outputs(3359);
    outputs(8656) <= (layer4_outputs(4125)) or (layer4_outputs(4521));
    outputs(8657) <= not(layer4_outputs(7675));
    outputs(8658) <= not(layer4_outputs(5739));
    outputs(8659) <= not(layer4_outputs(9632)) or (layer4_outputs(5733));
    outputs(8660) <= not((layer4_outputs(9391)) xor (layer4_outputs(1376)));
    outputs(8661) <= (layer4_outputs(9717)) and not (layer4_outputs(10068));
    outputs(8662) <= not((layer4_outputs(9742)) xor (layer4_outputs(9372)));
    outputs(8663) <= (layer4_outputs(895)) xor (layer4_outputs(10016));
    outputs(8664) <= (layer4_outputs(9270)) xor (layer4_outputs(10047));
    outputs(8665) <= layer4_outputs(7651);
    outputs(8666) <= layer4_outputs(60);
    outputs(8667) <= not(layer4_outputs(163));
    outputs(8668) <= layer4_outputs(2996);
    outputs(8669) <= (layer4_outputs(10064)) or (layer4_outputs(105));
    outputs(8670) <= not((layer4_outputs(1370)) xor (layer4_outputs(1046)));
    outputs(8671) <= not((layer4_outputs(1465)) xor (layer4_outputs(5469)));
    outputs(8672) <= layer4_outputs(3715);
    outputs(8673) <= layer4_outputs(48);
    outputs(8674) <= not((layer4_outputs(4353)) xor (layer4_outputs(5349)));
    outputs(8675) <= (layer4_outputs(9220)) or (layer4_outputs(4247));
    outputs(8676) <= layer4_outputs(6410);
    outputs(8677) <= not((layer4_outputs(1097)) xor (layer4_outputs(9870)));
    outputs(8678) <= not(layer4_outputs(6047));
    outputs(8679) <= not(layer4_outputs(208)) or (layer4_outputs(5109));
    outputs(8680) <= not((layer4_outputs(130)) xor (layer4_outputs(9672)));
    outputs(8681) <= not(layer4_outputs(9860));
    outputs(8682) <= not((layer4_outputs(2061)) xor (layer4_outputs(5972)));
    outputs(8683) <= layer4_outputs(2537);
    outputs(8684) <= not(layer4_outputs(7639));
    outputs(8685) <= (layer4_outputs(9359)) xor (layer4_outputs(1554));
    outputs(8686) <= not(layer4_outputs(1212)) or (layer4_outputs(2441));
    outputs(8687) <= (layer4_outputs(4349)) xor (layer4_outputs(2254));
    outputs(8688) <= not(layer4_outputs(4208));
    outputs(8689) <= not((layer4_outputs(5825)) xor (layer4_outputs(5389)));
    outputs(8690) <= not(layer4_outputs(956));
    outputs(8691) <= not((layer4_outputs(456)) xor (layer4_outputs(8203)));
    outputs(8692) <= layer4_outputs(5575);
    outputs(8693) <= not(layer4_outputs(6906));
    outputs(8694) <= layer4_outputs(4517);
    outputs(8695) <= layer4_outputs(7251);
    outputs(8696) <= layer4_outputs(5790);
    outputs(8697) <= (layer4_outputs(8250)) or (layer4_outputs(1159));
    outputs(8698) <= not((layer4_outputs(7328)) xor (layer4_outputs(3201)));
    outputs(8699) <= not((layer4_outputs(1881)) xor (layer4_outputs(9231)));
    outputs(8700) <= layer4_outputs(8019);
    outputs(8701) <= layer4_outputs(218);
    outputs(8702) <= not(layer4_outputs(8516)) or (layer4_outputs(1648));
    outputs(8703) <= layer4_outputs(4084);
    outputs(8704) <= not((layer4_outputs(2959)) xor (layer4_outputs(4325)));
    outputs(8705) <= not(layer4_outputs(136));
    outputs(8706) <= layer4_outputs(6294);
    outputs(8707) <= not(layer4_outputs(704));
    outputs(8708) <= not((layer4_outputs(7320)) and (layer4_outputs(4438)));
    outputs(8709) <= not(layer4_outputs(8589));
    outputs(8710) <= not(layer4_outputs(5851));
    outputs(8711) <= layer4_outputs(1669);
    outputs(8712) <= layer4_outputs(9395);
    outputs(8713) <= (layer4_outputs(6826)) xor (layer4_outputs(807));
    outputs(8714) <= (layer4_outputs(9026)) xor (layer4_outputs(9103));
    outputs(8715) <= layer4_outputs(8241);
    outputs(8716) <= not((layer4_outputs(6470)) xor (layer4_outputs(4482)));
    outputs(8717) <= not((layer4_outputs(1390)) xor (layer4_outputs(7381)));
    outputs(8718) <= layer4_outputs(1255);
    outputs(8719) <= not(layer4_outputs(9789));
    outputs(8720) <= layer4_outputs(9399);
    outputs(8721) <= not(layer4_outputs(893)) or (layer4_outputs(5471));
    outputs(8722) <= not(layer4_outputs(8624));
    outputs(8723) <= not((layer4_outputs(5536)) xor (layer4_outputs(8209)));
    outputs(8724) <= layer4_outputs(2502);
    outputs(8725) <= layer4_outputs(2684);
    outputs(8726) <= not(layer4_outputs(3918));
    outputs(8727) <= layer4_outputs(8183);
    outputs(8728) <= not(layer4_outputs(6449)) or (layer4_outputs(2578));
    outputs(8729) <= layer4_outputs(170);
    outputs(8730) <= not(layer4_outputs(4790));
    outputs(8731) <= (layer4_outputs(8604)) xor (layer4_outputs(1223));
    outputs(8732) <= layer4_outputs(2750);
    outputs(8733) <= (layer4_outputs(8110)) and not (layer4_outputs(3780));
    outputs(8734) <= not(layer4_outputs(7964));
    outputs(8735) <= not(layer4_outputs(24)) or (layer4_outputs(4997));
    outputs(8736) <= not(layer4_outputs(3102));
    outputs(8737) <= not(layer4_outputs(5225)) or (layer4_outputs(296));
    outputs(8738) <= (layer4_outputs(1662)) and (layer4_outputs(7965));
    outputs(8739) <= (layer4_outputs(6327)) xor (layer4_outputs(9806));
    outputs(8740) <= not((layer4_outputs(7493)) xor (layer4_outputs(7224)));
    outputs(8741) <= (layer4_outputs(719)) or (layer4_outputs(4131));
    outputs(8742) <= not(layer4_outputs(9984)) or (layer4_outputs(6323));
    outputs(8743) <= (layer4_outputs(10151)) or (layer4_outputs(8728));
    outputs(8744) <= (layer4_outputs(5313)) xor (layer4_outputs(466));
    outputs(8745) <= (layer4_outputs(6025)) and not (layer4_outputs(5496));
    outputs(8746) <= (layer4_outputs(2743)) and (layer4_outputs(9749));
    outputs(8747) <= not((layer4_outputs(3658)) or (layer4_outputs(9917)));
    outputs(8748) <= (layer4_outputs(3853)) and not (layer4_outputs(3577));
    outputs(8749) <= not(layer4_outputs(1777));
    outputs(8750) <= not(layer4_outputs(6259)) or (layer4_outputs(275));
    outputs(8751) <= not((layer4_outputs(5580)) or (layer4_outputs(1400)));
    outputs(8752) <= not((layer4_outputs(8520)) xor (layer4_outputs(8439)));
    outputs(8753) <= '1';
    outputs(8754) <= not(layer4_outputs(7078));
    outputs(8755) <= not((layer4_outputs(2647)) xor (layer4_outputs(9353)));
    outputs(8756) <= (layer4_outputs(7455)) xor (layer4_outputs(4064));
    outputs(8757) <= not(layer4_outputs(8985));
    outputs(8758) <= not(layer4_outputs(6892)) or (layer4_outputs(8151));
    outputs(8759) <= layer4_outputs(4358);
    outputs(8760) <= layer4_outputs(7805);
    outputs(8761) <= layer4_outputs(5169);
    outputs(8762) <= not(layer4_outputs(5431)) or (layer4_outputs(5116));
    outputs(8763) <= not(layer4_outputs(1337));
    outputs(8764) <= (layer4_outputs(5908)) xor (layer4_outputs(3889));
    outputs(8765) <= not(layer4_outputs(1258));
    outputs(8766) <= not(layer4_outputs(8001));
    outputs(8767) <= layer4_outputs(3065);
    outputs(8768) <= layer4_outputs(7144);
    outputs(8769) <= layer4_outputs(1706);
    outputs(8770) <= not(layer4_outputs(6973));
    outputs(8771) <= layer4_outputs(5524);
    outputs(8772) <= layer4_outputs(6169);
    outputs(8773) <= not(layer4_outputs(1191));
    outputs(8774) <= not(layer4_outputs(3634));
    outputs(8775) <= not(layer4_outputs(4740));
    outputs(8776) <= layer4_outputs(1876);
    outputs(8777) <= layer4_outputs(9598);
    outputs(8778) <= not((layer4_outputs(3374)) and (layer4_outputs(8375)));
    outputs(8779) <= (layer4_outputs(9225)) or (layer4_outputs(8068));
    outputs(8780) <= not(layer4_outputs(679));
    outputs(8781) <= layer4_outputs(3430);
    outputs(8782) <= layer4_outputs(43);
    outputs(8783) <= (layer4_outputs(2973)) and not (layer4_outputs(1734));
    outputs(8784) <= not((layer4_outputs(2765)) xor (layer4_outputs(7252)));
    outputs(8785) <= not(layer4_outputs(8596));
    outputs(8786) <= layer4_outputs(3172);
    outputs(8787) <= layer4_outputs(1120);
    outputs(8788) <= (layer4_outputs(5374)) xor (layer4_outputs(8126));
    outputs(8789) <= not((layer4_outputs(7065)) and (layer4_outputs(6862)));
    outputs(8790) <= not(layer4_outputs(452));
    outputs(8791) <= (layer4_outputs(8611)) xor (layer4_outputs(4299));
    outputs(8792) <= not(layer4_outputs(5254)) or (layer4_outputs(4542));
    outputs(8793) <= (layer4_outputs(636)) and not (layer4_outputs(4122));
    outputs(8794) <= (layer4_outputs(1932)) xor (layer4_outputs(3399));
    outputs(8795) <= layer4_outputs(1661);
    outputs(8796) <= not(layer4_outputs(4484));
    outputs(8797) <= not(layer4_outputs(740));
    outputs(8798) <= (layer4_outputs(7373)) or (layer4_outputs(3321));
    outputs(8799) <= not(layer4_outputs(7895));
    outputs(8800) <= layer4_outputs(4928);
    outputs(8801) <= not((layer4_outputs(9725)) and (layer4_outputs(7175)));
    outputs(8802) <= (layer4_outputs(8205)) xor (layer4_outputs(7262));
    outputs(8803) <= not(layer4_outputs(752));
    outputs(8804) <= not(layer4_outputs(4698));
    outputs(8805) <= not(layer4_outputs(3203));
    outputs(8806) <= (layer4_outputs(7241)) and (layer4_outputs(405));
    outputs(8807) <= not(layer4_outputs(1364));
    outputs(8808) <= not((layer4_outputs(5059)) and (layer4_outputs(8893)));
    outputs(8809) <= layer4_outputs(4276);
    outputs(8810) <= not(layer4_outputs(503)) or (layer4_outputs(2470));
    outputs(8811) <= not(layer4_outputs(5962));
    outputs(8812) <= not(layer4_outputs(7065)) or (layer4_outputs(5265));
    outputs(8813) <= not(layer4_outputs(6218)) or (layer4_outputs(7161));
    outputs(8814) <= not((layer4_outputs(2138)) xor (layer4_outputs(5955)));
    outputs(8815) <= not(layer4_outputs(7242));
    outputs(8816) <= not((layer4_outputs(1863)) xor (layer4_outputs(765)));
    outputs(8817) <= layer4_outputs(8587);
    outputs(8818) <= not(layer4_outputs(8179));
    outputs(8819) <= layer4_outputs(6103);
    outputs(8820) <= not(layer4_outputs(8279));
    outputs(8821) <= not(layer4_outputs(6393));
    outputs(8822) <= layer4_outputs(6318);
    outputs(8823) <= not(layer4_outputs(1144));
    outputs(8824) <= not(layer4_outputs(6733));
    outputs(8825) <= not((layer4_outputs(5799)) xor (layer4_outputs(7925)));
    outputs(8826) <= (layer4_outputs(2032)) and not (layer4_outputs(9627));
    outputs(8827) <= not(layer4_outputs(8386)) or (layer4_outputs(9396));
    outputs(8828) <= not(layer4_outputs(1614));
    outputs(8829) <= layer4_outputs(8901);
    outputs(8830) <= not(layer4_outputs(1387));
    outputs(8831) <= not((layer4_outputs(8984)) or (layer4_outputs(1475)));
    outputs(8832) <= (layer4_outputs(6520)) and not (layer4_outputs(4852));
    outputs(8833) <= not(layer4_outputs(846));
    outputs(8834) <= (layer4_outputs(2966)) xor (layer4_outputs(758));
    outputs(8835) <= layer4_outputs(1324);
    outputs(8836) <= not(layer4_outputs(3505)) or (layer4_outputs(10110));
    outputs(8837) <= not((layer4_outputs(6131)) xor (layer4_outputs(4723)));
    outputs(8838) <= not(layer4_outputs(273));
    outputs(8839) <= layer4_outputs(54);
    outputs(8840) <= not((layer4_outputs(7222)) or (layer4_outputs(10)));
    outputs(8841) <= not(layer4_outputs(2867));
    outputs(8842) <= not(layer4_outputs(5010));
    outputs(8843) <= not(layer4_outputs(3726));
    outputs(8844) <= (layer4_outputs(4419)) xor (layer4_outputs(6565));
    outputs(8845) <= layer4_outputs(2246);
    outputs(8846) <= layer4_outputs(8742);
    outputs(8847) <= layer4_outputs(6636);
    outputs(8848) <= not((layer4_outputs(5014)) and (layer4_outputs(9648)));
    outputs(8849) <= (layer4_outputs(3007)) xor (layer4_outputs(7540));
    outputs(8850) <= not(layer4_outputs(8428));
    outputs(8851) <= (layer4_outputs(6775)) and not (layer4_outputs(868));
    outputs(8852) <= not(layer4_outputs(8298));
    outputs(8853) <= not((layer4_outputs(4167)) and (layer4_outputs(9274)));
    outputs(8854) <= layer4_outputs(4658);
    outputs(8855) <= layer4_outputs(5754);
    outputs(8856) <= not(layer4_outputs(6685));
    outputs(8857) <= not(layer4_outputs(7348));
    outputs(8858) <= not(layer4_outputs(3382));
    outputs(8859) <= layer4_outputs(6370);
    outputs(8860) <= layer4_outputs(10004);
    outputs(8861) <= layer4_outputs(3135);
    outputs(8862) <= layer4_outputs(9794);
    outputs(8863) <= not((layer4_outputs(3750)) xor (layer4_outputs(1949)));
    outputs(8864) <= '1';
    outputs(8865) <= not(layer4_outputs(10175));
    outputs(8866) <= (layer4_outputs(4711)) or (layer4_outputs(4888));
    outputs(8867) <= layer4_outputs(9125);
    outputs(8868) <= not(layer4_outputs(1577));
    outputs(8869) <= (layer4_outputs(3378)) and not (layer4_outputs(9391));
    outputs(8870) <= (layer4_outputs(8808)) xor (layer4_outputs(6224));
    outputs(8871) <= not((layer4_outputs(5502)) and (layer4_outputs(6928)));
    outputs(8872) <= not((layer4_outputs(4047)) xor (layer4_outputs(3751)));
    outputs(8873) <= not(layer4_outputs(30)) or (layer4_outputs(8685));
    outputs(8874) <= layer4_outputs(8041);
    outputs(8875) <= (layer4_outputs(4344)) xor (layer4_outputs(4878));
    outputs(8876) <= not(layer4_outputs(10019)) or (layer4_outputs(1676));
    outputs(8877) <= not((layer4_outputs(9479)) and (layer4_outputs(8952)));
    outputs(8878) <= (layer4_outputs(7137)) and not (layer4_outputs(1403));
    outputs(8879) <= not(layer4_outputs(9838));
    outputs(8880) <= layer4_outputs(8034);
    outputs(8881) <= layer4_outputs(6751);
    outputs(8882) <= (layer4_outputs(9344)) or (layer4_outputs(1588));
    outputs(8883) <= not(layer4_outputs(2201));
    outputs(8884) <= (layer4_outputs(6519)) xor (layer4_outputs(5121));
    outputs(8885) <= not(layer4_outputs(1076));
    outputs(8886) <= not(layer4_outputs(2136));
    outputs(8887) <= (layer4_outputs(9411)) xor (layer4_outputs(8631));
    outputs(8888) <= (layer4_outputs(1749)) xor (layer4_outputs(3305));
    outputs(8889) <= (layer4_outputs(5650)) xor (layer4_outputs(7050));
    outputs(8890) <= layer4_outputs(6675);
    outputs(8891) <= not(layer4_outputs(6746));
    outputs(8892) <= not((layer4_outputs(7744)) xor (layer4_outputs(9344)));
    outputs(8893) <= layer4_outputs(7555);
    outputs(8894) <= layer4_outputs(5408);
    outputs(8895) <= (layer4_outputs(2512)) xor (layer4_outputs(8372));
    outputs(8896) <= not(layer4_outputs(251));
    outputs(8897) <= not((layer4_outputs(10238)) and (layer4_outputs(1611)));
    outputs(8898) <= not(layer4_outputs(7823));
    outputs(8899) <= layer4_outputs(2329);
    outputs(8900) <= not((layer4_outputs(6599)) or (layer4_outputs(2985)));
    outputs(8901) <= not(layer4_outputs(9987)) or (layer4_outputs(6490));
    outputs(8902) <= layer4_outputs(1336);
    outputs(8903) <= not(layer4_outputs(5303));
    outputs(8904) <= not((layer4_outputs(5581)) and (layer4_outputs(8218)));
    outputs(8905) <= (layer4_outputs(2207)) and not (layer4_outputs(9064));
    outputs(8906) <= (layer4_outputs(5610)) or (layer4_outputs(4940));
    outputs(8907) <= (layer4_outputs(430)) xor (layer4_outputs(2505));
    outputs(8908) <= (layer4_outputs(6257)) xor (layer4_outputs(6282));
    outputs(8909) <= not(layer4_outputs(9463));
    outputs(8910) <= layer4_outputs(7269);
    outputs(8911) <= not(layer4_outputs(973));
    outputs(8912) <= not(layer4_outputs(2345)) or (layer4_outputs(8020));
    outputs(8913) <= (layer4_outputs(231)) xor (layer4_outputs(1230));
    outputs(8914) <= not(layer4_outputs(2076)) or (layer4_outputs(10200));
    outputs(8915) <= (layer4_outputs(10187)) and (layer4_outputs(5811));
    outputs(8916) <= layer4_outputs(1335);
    outputs(8917) <= layer4_outputs(8087);
    outputs(8918) <= not((layer4_outputs(7090)) xor (layer4_outputs(6652)));
    outputs(8919) <= not(layer4_outputs(9355));
    outputs(8920) <= not(layer4_outputs(3204));
    outputs(8921) <= layer4_outputs(4650);
    outputs(8922) <= not(layer4_outputs(5381));
    outputs(8923) <= (layer4_outputs(1030)) xor (layer4_outputs(3669));
    outputs(8924) <= not(layer4_outputs(8432)) or (layer4_outputs(8478));
    outputs(8925) <= not((layer4_outputs(7814)) xor (layer4_outputs(6833)));
    outputs(8926) <= not((layer4_outputs(9146)) and (layer4_outputs(4029)));
    outputs(8927) <= not(layer4_outputs(1316));
    outputs(8928) <= not(layer4_outputs(7245));
    outputs(8929) <= layer4_outputs(2481);
    outputs(8930) <= not((layer4_outputs(8636)) xor (layer4_outputs(5415)));
    outputs(8931) <= not(layer4_outputs(9194));
    outputs(8932) <= not((layer4_outputs(7)) and (layer4_outputs(7240)));
    outputs(8933) <= not(layer4_outputs(9459));
    outputs(8934) <= not((layer4_outputs(3685)) xor (layer4_outputs(10223)));
    outputs(8935) <= layer4_outputs(4005);
    outputs(8936) <= not(layer4_outputs(4824));
    outputs(8937) <= layer4_outputs(8813);
    outputs(8938) <= not((layer4_outputs(7598)) and (layer4_outputs(8428)));
    outputs(8939) <= layer4_outputs(7379);
    outputs(8940) <= (layer4_outputs(3904)) xor (layer4_outputs(2927));
    outputs(8941) <= not((layer4_outputs(9981)) xor (layer4_outputs(7386)));
    outputs(8942) <= layer4_outputs(6831);
    outputs(8943) <= not(layer4_outputs(5549));
    outputs(8944) <= not(layer4_outputs(6163)) or (layer4_outputs(6286));
    outputs(8945) <= not((layer4_outputs(5633)) or (layer4_outputs(8660)));
    outputs(8946) <= not((layer4_outputs(6940)) xor (layer4_outputs(1953)));
    outputs(8947) <= not((layer4_outputs(3887)) and (layer4_outputs(4537)));
    outputs(8948) <= not((layer4_outputs(10069)) xor (layer4_outputs(2395)));
    outputs(8949) <= not((layer4_outputs(4578)) and (layer4_outputs(318)));
    outputs(8950) <= (layer4_outputs(8262)) and not (layer4_outputs(2466));
    outputs(8951) <= not((layer4_outputs(6970)) xor (layer4_outputs(4562)));
    outputs(8952) <= not((layer4_outputs(4162)) xor (layer4_outputs(2067)));
    outputs(8953) <= (layer4_outputs(7708)) xor (layer4_outputs(1407));
    outputs(8954) <= layer4_outputs(8682);
    outputs(8955) <= layer4_outputs(7344);
    outputs(8956) <= not((layer4_outputs(5713)) xor (layer4_outputs(8991)));
    outputs(8957) <= not(layer4_outputs(5544));
    outputs(8958) <= (layer4_outputs(8277)) xor (layer4_outputs(4543));
    outputs(8959) <= not(layer4_outputs(5865));
    outputs(8960) <= layer4_outputs(6362);
    outputs(8961) <= (layer4_outputs(8607)) xor (layer4_outputs(8927));
    outputs(8962) <= not(layer4_outputs(1966));
    outputs(8963) <= (layer4_outputs(2043)) xor (layer4_outputs(7443));
    outputs(8964) <= not(layer4_outputs(4194));
    outputs(8965) <= not((layer4_outputs(6796)) xor (layer4_outputs(2792)));
    outputs(8966) <= not(layer4_outputs(1570));
    outputs(8967) <= '1';
    outputs(8968) <= layer4_outputs(61);
    outputs(8969) <= layer4_outputs(8798);
    outputs(8970) <= not(layer4_outputs(1404));
    outputs(8971) <= (layer4_outputs(131)) and not (layer4_outputs(5508));
    outputs(8972) <= layer4_outputs(8560);
    outputs(8973) <= layer4_outputs(9132);
    outputs(8974) <= not(layer4_outputs(2235));
    outputs(8975) <= not((layer4_outputs(1969)) xor (layer4_outputs(2617)));
    outputs(8976) <= (layer4_outputs(5607)) and (layer4_outputs(842));
    outputs(8977) <= layer4_outputs(2598);
    outputs(8978) <= not(layer4_outputs(9525));
    outputs(8979) <= layer4_outputs(7444);
    outputs(8980) <= layer4_outputs(2947);
    outputs(8981) <= not((layer4_outputs(926)) and (layer4_outputs(2671)));
    outputs(8982) <= (layer4_outputs(8701)) and not (layer4_outputs(6093));
    outputs(8983) <= layer4_outputs(8072);
    outputs(8984) <= not((layer4_outputs(7781)) xor (layer4_outputs(4298)));
    outputs(8985) <= not(layer4_outputs(4268));
    outputs(8986) <= not(layer4_outputs(8291));
    outputs(8987) <= layer4_outputs(8225);
    outputs(8988) <= (layer4_outputs(7590)) xor (layer4_outputs(8231));
    outputs(8989) <= (layer4_outputs(2859)) xor (layer4_outputs(6443));
    outputs(8990) <= not(layer4_outputs(7550)) or (layer4_outputs(1732));
    outputs(8991) <= (layer4_outputs(6907)) and (layer4_outputs(7692));
    outputs(8992) <= layer4_outputs(5463);
    outputs(8993) <= layer4_outputs(4262);
    outputs(8994) <= not(layer4_outputs(355));
    outputs(8995) <= layer4_outputs(8473);
    outputs(8996) <= not(layer4_outputs(3506));
    outputs(8997) <= not(layer4_outputs(37));
    outputs(8998) <= layer4_outputs(5055);
    outputs(8999) <= (layer4_outputs(1459)) and not (layer4_outputs(5306));
    outputs(9000) <= layer4_outputs(2241);
    outputs(9001) <= layer4_outputs(1292);
    outputs(9002) <= not(layer4_outputs(9248)) or (layer4_outputs(2847));
    outputs(9003) <= (layer4_outputs(2722)) or (layer4_outputs(2893));
    outputs(9004) <= (layer4_outputs(4215)) xor (layer4_outputs(4888));
    outputs(9005) <= not(layer4_outputs(9760)) or (layer4_outputs(9345));
    outputs(9006) <= layer4_outputs(877);
    outputs(9007) <= not(layer4_outputs(6997));
    outputs(9008) <= not(layer4_outputs(4771));
    outputs(9009) <= not((layer4_outputs(9514)) xor (layer4_outputs(9271)));
    outputs(9010) <= (layer4_outputs(3627)) xor (layer4_outputs(4176));
    outputs(9011) <= not(layer4_outputs(2949));
    outputs(9012) <= layer4_outputs(5289);
    outputs(9013) <= not(layer4_outputs(9133));
    outputs(9014) <= layer4_outputs(6220);
    outputs(9015) <= (layer4_outputs(5135)) xor (layer4_outputs(4143));
    outputs(9016) <= not(layer4_outputs(7443));
    outputs(9017) <= not(layer4_outputs(4109));
    outputs(9018) <= layer4_outputs(3202);
    outputs(9019) <= (layer4_outputs(3231)) or (layer4_outputs(3716));
    outputs(9020) <= layer4_outputs(3462);
    outputs(9021) <= not((layer4_outputs(8330)) xor (layer4_outputs(673)));
    outputs(9022) <= layer4_outputs(2338);
    outputs(9023) <= (layer4_outputs(19)) and not (layer4_outputs(9172));
    outputs(9024) <= layer4_outputs(1825);
    outputs(9025) <= not(layer4_outputs(4826)) or (layer4_outputs(7682));
    outputs(9026) <= layer4_outputs(1346);
    outputs(9027) <= layer4_outputs(5168);
    outputs(9028) <= not(layer4_outputs(5413));
    outputs(9029) <= not(layer4_outputs(8031));
    outputs(9030) <= (layer4_outputs(5435)) or (layer4_outputs(8859));
    outputs(9031) <= (layer4_outputs(4360)) xor (layer4_outputs(4725));
    outputs(9032) <= not(layer4_outputs(5095));
    outputs(9033) <= (layer4_outputs(2781)) or (layer4_outputs(1586));
    outputs(9034) <= not(layer4_outputs(7579));
    outputs(9035) <= layer4_outputs(10057);
    outputs(9036) <= not(layer4_outputs(9219));
    outputs(9037) <= not(layer4_outputs(28));
    outputs(9038) <= not(layer4_outputs(2114));
    outputs(9039) <= (layer4_outputs(15)) xor (layer4_outputs(6817));
    outputs(9040) <= not(layer4_outputs(5914)) or (layer4_outputs(2624));
    outputs(9041) <= not(layer4_outputs(5706));
    outputs(9042) <= not(layer4_outputs(8662));
    outputs(9043) <= not(layer4_outputs(6384)) or (layer4_outputs(1950));
    outputs(9044) <= layer4_outputs(6206);
    outputs(9045) <= not((layer4_outputs(7096)) xor (layer4_outputs(3076)));
    outputs(9046) <= layer4_outputs(380);
    outputs(9047) <= layer4_outputs(2066);
    outputs(9048) <= not(layer4_outputs(559));
    outputs(9049) <= layer4_outputs(6492);
    outputs(9050) <= layer4_outputs(115);
    outputs(9051) <= (layer4_outputs(6441)) xor (layer4_outputs(9657));
    outputs(9052) <= layer4_outputs(5597);
    outputs(9053) <= not(layer4_outputs(1100));
    outputs(9054) <= not((layer4_outputs(10184)) and (layer4_outputs(6460)));
    outputs(9055) <= layer4_outputs(6203);
    outputs(9056) <= not(layer4_outputs(3085));
    outputs(9057) <= layer4_outputs(6834);
    outputs(9058) <= not((layer4_outputs(2053)) xor (layer4_outputs(8080)));
    outputs(9059) <= (layer4_outputs(5465)) xor (layer4_outputs(9739));
    outputs(9060) <= layer4_outputs(5696);
    outputs(9061) <= (layer4_outputs(9598)) and (layer4_outputs(6539));
    outputs(9062) <= not(layer4_outputs(2044));
    outputs(9063) <= not(layer4_outputs(3550));
    outputs(9064) <= not(layer4_outputs(8580));
    outputs(9065) <= layer4_outputs(9491);
    outputs(9066) <= (layer4_outputs(7162)) and (layer4_outputs(3817));
    outputs(9067) <= (layer4_outputs(7996)) xor (layer4_outputs(9748));
    outputs(9068) <= not(layer4_outputs(2838));
    outputs(9069) <= not((layer4_outputs(1728)) xor (layer4_outputs(9822)));
    outputs(9070) <= not((layer4_outputs(9545)) or (layer4_outputs(6586)));
    outputs(9071) <= not(layer4_outputs(5674));
    outputs(9072) <= layer4_outputs(143);
    outputs(9073) <= not(layer4_outputs(1966)) or (layer4_outputs(7308));
    outputs(9074) <= (layer4_outputs(8898)) xor (layer4_outputs(6745));
    outputs(9075) <= not((layer4_outputs(2376)) xor (layer4_outputs(866)));
    outputs(9076) <= not((layer4_outputs(8210)) xor (layer4_outputs(3555)));
    outputs(9077) <= not(layer4_outputs(7582)) or (layer4_outputs(267));
    outputs(9078) <= (layer4_outputs(4532)) and not (layer4_outputs(8099));
    outputs(9079) <= layer4_outputs(7177);
    outputs(9080) <= (layer4_outputs(8048)) and not (layer4_outputs(144));
    outputs(9081) <= layer4_outputs(3215);
    outputs(9082) <= layer4_outputs(1857);
    outputs(9083) <= not(layer4_outputs(3595));
    outputs(9084) <= not((layer4_outputs(128)) xor (layer4_outputs(7401)));
    outputs(9085) <= (layer4_outputs(6657)) and (layer4_outputs(3065));
    outputs(9086) <= layer4_outputs(7024);
    outputs(9087) <= not((layer4_outputs(7582)) xor (layer4_outputs(4639)));
    outputs(9088) <= not(layer4_outputs(6502)) or (layer4_outputs(2820));
    outputs(9089) <= layer4_outputs(6434);
    outputs(9090) <= not(layer4_outputs(2085));
    outputs(9091) <= not(layer4_outputs(2754)) or (layer4_outputs(9716));
    outputs(9092) <= not(layer4_outputs(6932)) or (layer4_outputs(6662));
    outputs(9093) <= not((layer4_outputs(4478)) and (layer4_outputs(4039)));
    outputs(9094) <= not((layer4_outputs(4513)) xor (layer4_outputs(4365)));
    outputs(9095) <= not(layer4_outputs(8358));
    outputs(9096) <= layer4_outputs(9716);
    outputs(9097) <= not((layer4_outputs(1664)) xor (layer4_outputs(6580)));
    outputs(9098) <= '1';
    outputs(9099) <= not((layer4_outputs(3625)) xor (layer4_outputs(947)));
    outputs(9100) <= not(layer4_outputs(10193)) or (layer4_outputs(5386));
    outputs(9101) <= layer4_outputs(8506);
    outputs(9102) <= (layer4_outputs(181)) or (layer4_outputs(3502));
    outputs(9103) <= not(layer4_outputs(9163)) or (layer4_outputs(8385));
    outputs(9104) <= not(layer4_outputs(2559)) or (layer4_outputs(1795));
    outputs(9105) <= not(layer4_outputs(5857));
    outputs(9106) <= (layer4_outputs(7702)) xor (layer4_outputs(8488));
    outputs(9107) <= not(layer4_outputs(9657));
    outputs(9108) <= not(layer4_outputs(1899));
    outputs(9109) <= layer4_outputs(244);
    outputs(9110) <= (layer4_outputs(5360)) xor (layer4_outputs(984));
    outputs(9111) <= not((layer4_outputs(2699)) or (layer4_outputs(5539)));
    outputs(9112) <= not(layer4_outputs(860)) or (layer4_outputs(1184));
    outputs(9113) <= not((layer4_outputs(2286)) and (layer4_outputs(3069)));
    outputs(9114) <= not(layer4_outputs(10182));
    outputs(9115) <= not(layer4_outputs(8741));
    outputs(9116) <= layer4_outputs(7949);
    outputs(9117) <= not(layer4_outputs(6723));
    outputs(9118) <= layer4_outputs(3296);
    outputs(9119) <= not(layer4_outputs(258));
    outputs(9120) <= not(layer4_outputs(847));
    outputs(9121) <= layer4_outputs(3800);
    outputs(9122) <= (layer4_outputs(4381)) and (layer4_outputs(1135));
    outputs(9123) <= not(layer4_outputs(2918));
    outputs(9124) <= layer4_outputs(6052);
    outputs(9125) <= (layer4_outputs(9188)) xor (layer4_outputs(7830));
    outputs(9126) <= (layer4_outputs(2778)) xor (layer4_outputs(5952));
    outputs(9127) <= (layer4_outputs(8500)) or (layer4_outputs(4912));
    outputs(9128) <= (layer4_outputs(7043)) or (layer4_outputs(1853));
    outputs(9129) <= not((layer4_outputs(7641)) xor (layer4_outputs(5420)));
    outputs(9130) <= layer4_outputs(9997);
    outputs(9131) <= layer4_outputs(4766);
    outputs(9132) <= not((layer4_outputs(7672)) or (layer4_outputs(976)));
    outputs(9133) <= layer4_outputs(7499);
    outputs(9134) <= not((layer4_outputs(683)) xor (layer4_outputs(5986)));
    outputs(9135) <= layer4_outputs(2660);
    outputs(9136) <= layer4_outputs(10020);
    outputs(9137) <= (layer4_outputs(855)) xor (layer4_outputs(6814));
    outputs(9138) <= (layer4_outputs(7926)) xor (layer4_outputs(9283));
    outputs(9139) <= not(layer4_outputs(8732));
    outputs(9140) <= not(layer4_outputs(3443));
    outputs(9141) <= (layer4_outputs(7739)) xor (layer4_outputs(9892));
    outputs(9142) <= not((layer4_outputs(3903)) and (layer4_outputs(3124)));
    outputs(9143) <= not(layer4_outputs(2546));
    outputs(9144) <= not(layer4_outputs(6178));
    outputs(9145) <= (layer4_outputs(3269)) xor (layer4_outputs(6308));
    outputs(9146) <= not(layer4_outputs(7392)) or (layer4_outputs(1806));
    outputs(9147) <= (layer4_outputs(2208)) and not (layer4_outputs(1312));
    outputs(9148) <= layer4_outputs(9334);
    outputs(9149) <= not((layer4_outputs(7631)) xor (layer4_outputs(1671)));
    outputs(9150) <= (layer4_outputs(6040)) and not (layer4_outputs(4662));
    outputs(9151) <= layer4_outputs(3080);
    outputs(9152) <= not(layer4_outputs(916));
    outputs(9153) <= layer4_outputs(2488);
    outputs(9154) <= layer4_outputs(8719);
    outputs(9155) <= not((layer4_outputs(1698)) or (layer4_outputs(4204)));
    outputs(9156) <= not(layer4_outputs(4544));
    outputs(9157) <= not((layer4_outputs(5223)) xor (layer4_outputs(8742)));
    outputs(9158) <= layer4_outputs(3138);
    outputs(9159) <= layer4_outputs(4516);
    outputs(9160) <= not((layer4_outputs(7647)) or (layer4_outputs(9012)));
    outputs(9161) <= not(layer4_outputs(8896));
    outputs(9162) <= not((layer4_outputs(10193)) and (layer4_outputs(2857)));
    outputs(9163) <= '1';
    outputs(9164) <= not(layer4_outputs(5082));
    outputs(9165) <= not(layer4_outputs(7999));
    outputs(9166) <= not(layer4_outputs(1888)) or (layer4_outputs(6410));
    outputs(9167) <= not(layer4_outputs(90)) or (layer4_outputs(5296));
    outputs(9168) <= not(layer4_outputs(5658));
    outputs(9169) <= layer4_outputs(6051);
    outputs(9170) <= layer4_outputs(9767);
    outputs(9171) <= (layer4_outputs(7030)) or (layer4_outputs(1591));
    outputs(9172) <= not(layer4_outputs(7335));
    outputs(9173) <= not((layer4_outputs(3909)) xor (layer4_outputs(6933)));
    outputs(9174) <= (layer4_outputs(3188)) xor (layer4_outputs(3514));
    outputs(9175) <= (layer4_outputs(5498)) xor (layer4_outputs(2025));
    outputs(9176) <= not(layer4_outputs(1502));
    outputs(9177) <= not(layer4_outputs(7136)) or (layer4_outputs(4408));
    outputs(9178) <= (layer4_outputs(7488)) xor (layer4_outputs(2769));
    outputs(9179) <= not(layer4_outputs(6392));
    outputs(9180) <= not(layer4_outputs(2509));
    outputs(9181) <= not(layer4_outputs(1143));
    outputs(9182) <= layer4_outputs(2176);
    outputs(9183) <= layer4_outputs(5369);
    outputs(9184) <= (layer4_outputs(1738)) xor (layer4_outputs(773));
    outputs(9185) <= not((layer4_outputs(2504)) xor (layer4_outputs(4134)));
    outputs(9186) <= not(layer4_outputs(563));
    outputs(9187) <= not(layer4_outputs(443));
    outputs(9188) <= not((layer4_outputs(5801)) and (layer4_outputs(1342)));
    outputs(9189) <= not(layer4_outputs(2423)) or (layer4_outputs(2034));
    outputs(9190) <= layer4_outputs(10212);
    outputs(9191) <= (layer4_outputs(328)) xor (layer4_outputs(5957));
    outputs(9192) <= layer4_outputs(3087);
    outputs(9193) <= (layer4_outputs(5554)) xor (layer4_outputs(8109));
    outputs(9194) <= not((layer4_outputs(7546)) xor (layer4_outputs(1551)));
    outputs(9195) <= layer4_outputs(10228);
    outputs(9196) <= (layer4_outputs(9787)) xor (layer4_outputs(7455));
    outputs(9197) <= not((layer4_outputs(3940)) xor (layer4_outputs(3455)));
    outputs(9198) <= (layer4_outputs(7605)) xor (layer4_outputs(4592));
    outputs(9199) <= (layer4_outputs(5983)) xor (layer4_outputs(8864));
    outputs(9200) <= not(layer4_outputs(9999));
    outputs(9201) <= (layer4_outputs(947)) xor (layer4_outputs(8504));
    outputs(9202) <= not(layer4_outputs(8583)) or (layer4_outputs(8188));
    outputs(9203) <= not((layer4_outputs(4518)) xor (layer4_outputs(230)));
    outputs(9204) <= layer4_outputs(8675);
    outputs(9205) <= not(layer4_outputs(8039));
    outputs(9206) <= (layer4_outputs(345)) or (layer4_outputs(2371));
    outputs(9207) <= not(layer4_outputs(6604));
    outputs(9208) <= (layer4_outputs(5280)) or (layer4_outputs(6140));
    outputs(9209) <= '1';
    outputs(9210) <= not((layer4_outputs(8981)) xor (layer4_outputs(3793)));
    outputs(9211) <= layer4_outputs(7277);
    outputs(9212) <= not(layer4_outputs(2570));
    outputs(9213) <= layer4_outputs(5543);
    outputs(9214) <= (layer4_outputs(7601)) or (layer4_outputs(8040));
    outputs(9215) <= layer4_outputs(2320);
    outputs(9216) <= not((layer4_outputs(7580)) xor (layer4_outputs(7034)));
    outputs(9217) <= not(layer4_outputs(5541)) or (layer4_outputs(8072));
    outputs(9218) <= not((layer4_outputs(845)) xor (layer4_outputs(3891)));
    outputs(9219) <= layer4_outputs(1701);
    outputs(9220) <= (layer4_outputs(4144)) xor (layer4_outputs(5951));
    outputs(9221) <= not((layer4_outputs(5637)) xor (layer4_outputs(2467)));
    outputs(9222) <= not((layer4_outputs(2983)) or (layer4_outputs(4514)));
    outputs(9223) <= not((layer4_outputs(4749)) xor (layer4_outputs(36)));
    outputs(9224) <= layer4_outputs(592);
    outputs(9225) <= (layer4_outputs(865)) xor (layer4_outputs(2347));
    outputs(9226) <= (layer4_outputs(5096)) xor (layer4_outputs(6920));
    outputs(9227) <= layer4_outputs(358);
    outputs(9228) <= layer4_outputs(2705);
    outputs(9229) <= not(layer4_outputs(3106));
    outputs(9230) <= (layer4_outputs(3275)) xor (layer4_outputs(7538));
    outputs(9231) <= layer4_outputs(1073);
    outputs(9232) <= (layer4_outputs(2200)) and not (layer4_outputs(3901));
    outputs(9233) <= layer4_outputs(428);
    outputs(9234) <= (layer4_outputs(7098)) and (layer4_outputs(7292));
    outputs(9235) <= layer4_outputs(8367);
    outputs(9236) <= not((layer4_outputs(7227)) xor (layer4_outputs(7628)));
    outputs(9237) <= not(layer4_outputs(4212));
    outputs(9238) <= layer4_outputs(8128);
    outputs(9239) <= (layer4_outputs(8501)) xor (layer4_outputs(8231));
    outputs(9240) <= layer4_outputs(1376);
    outputs(9241) <= not(layer4_outputs(9388));
    outputs(9242) <= layer4_outputs(5610);
    outputs(9243) <= layer4_outputs(676);
    outputs(9244) <= not(layer4_outputs(6237));
    outputs(9245) <= not((layer4_outputs(9543)) and (layer4_outputs(5393)));
    outputs(9246) <= not(layer4_outputs(3516));
    outputs(9247) <= layer4_outputs(2309);
    outputs(9248) <= not((layer4_outputs(8414)) xor (layer4_outputs(7182)));
    outputs(9249) <= layer4_outputs(1821);
    outputs(9250) <= not((layer4_outputs(434)) xor (layer4_outputs(1521)));
    outputs(9251) <= not((layer4_outputs(9382)) xor (layer4_outputs(6408)));
    outputs(9252) <= not(layer4_outputs(9229));
    outputs(9253) <= layer4_outputs(7879);
    outputs(9254) <= not((layer4_outputs(6501)) xor (layer4_outputs(5112)));
    outputs(9255) <= layer4_outputs(8526);
    outputs(9256) <= not(layer4_outputs(5478));
    outputs(9257) <= layer4_outputs(6495);
    outputs(9258) <= not((layer4_outputs(9095)) xor (layer4_outputs(772)));
    outputs(9259) <= layer4_outputs(9247);
    outputs(9260) <= not((layer4_outputs(5719)) or (layer4_outputs(96)));
    outputs(9261) <= (layer4_outputs(9366)) and not (layer4_outputs(9526));
    outputs(9262) <= not((layer4_outputs(625)) xor (layer4_outputs(3003)));
    outputs(9263) <= not(layer4_outputs(7080));
    outputs(9264) <= not((layer4_outputs(8181)) xor (layer4_outputs(1440)));
    outputs(9265) <= not(layer4_outputs(2657));
    outputs(9266) <= layer4_outputs(4388);
    outputs(9267) <= not(layer4_outputs(7182));
    outputs(9268) <= (layer4_outputs(3366)) xor (layer4_outputs(235));
    outputs(9269) <= layer4_outputs(4805);
    outputs(9270) <= (layer4_outputs(6917)) xor (layer4_outputs(4646));
    outputs(9271) <= (layer4_outputs(6059)) and not (layer4_outputs(2391));
    outputs(9272) <= not(layer4_outputs(9514));
    outputs(9273) <= not(layer4_outputs(3347));
    outputs(9274) <= (layer4_outputs(2278)) xor (layer4_outputs(6258));
    outputs(9275) <= layer4_outputs(941);
    outputs(9276) <= layer4_outputs(9938);
    outputs(9277) <= not(layer4_outputs(1280));
    outputs(9278) <= layer4_outputs(1050);
    outputs(9279) <= not(layer4_outputs(5718));
    outputs(9280) <= not(layer4_outputs(6947));
    outputs(9281) <= layer4_outputs(3765);
    outputs(9282) <= layer4_outputs(7823);
    outputs(9283) <= not((layer4_outputs(1110)) xor (layer4_outputs(3030)));
    outputs(9284) <= layer4_outputs(494);
    outputs(9285) <= (layer4_outputs(9501)) xor (layer4_outputs(4735));
    outputs(9286) <= (layer4_outputs(3849)) xor (layer4_outputs(6664));
    outputs(9287) <= not(layer4_outputs(4637));
    outputs(9288) <= (layer4_outputs(4713)) and not (layer4_outputs(560));
    outputs(9289) <= layer4_outputs(2974);
    outputs(9290) <= not((layer4_outputs(2191)) xor (layer4_outputs(1218)));
    outputs(9291) <= not(layer4_outputs(3171));
    outputs(9292) <= (layer4_outputs(940)) xor (layer4_outputs(8786));
    outputs(9293) <= layer4_outputs(7901);
    outputs(9294) <= layer4_outputs(410);
    outputs(9295) <= not(layer4_outputs(733));
    outputs(9296) <= not(layer4_outputs(704));
    outputs(9297) <= layer4_outputs(2152);
    outputs(9298) <= not(layer4_outputs(3018));
    outputs(9299) <= layer4_outputs(4709);
    outputs(9300) <= (layer4_outputs(1943)) xor (layer4_outputs(2383));
    outputs(9301) <= not((layer4_outputs(9869)) xor (layer4_outputs(8065)));
    outputs(9302) <= layer4_outputs(5531);
    outputs(9303) <= layer4_outputs(496);
    outputs(9304) <= layer4_outputs(9633);
    outputs(9305) <= not(layer4_outputs(6473));
    outputs(9306) <= not((layer4_outputs(5553)) or (layer4_outputs(5631)));
    outputs(9307) <= layer4_outputs(4348);
    outputs(9308) <= not((layer4_outputs(10084)) xor (layer4_outputs(1876)));
    outputs(9309) <= not(layer4_outputs(2608));
    outputs(9310) <= not(layer4_outputs(1506));
    outputs(9311) <= not(layer4_outputs(2763));
    outputs(9312) <= not(layer4_outputs(9122));
    outputs(9313) <= layer4_outputs(1480);
    outputs(9314) <= layer4_outputs(7319);
    outputs(9315) <= not((layer4_outputs(7525)) xor (layer4_outputs(777)));
    outputs(9316) <= not((layer4_outputs(8337)) xor (layer4_outputs(3262)));
    outputs(9317) <= (layer4_outputs(1183)) and (layer4_outputs(8180));
    outputs(9318) <= layer4_outputs(648);
    outputs(9319) <= (layer4_outputs(1238)) xor (layer4_outputs(649));
    outputs(9320) <= not((layer4_outputs(8237)) xor (layer4_outputs(8387)));
    outputs(9321) <= not((layer4_outputs(10028)) xor (layer4_outputs(9280)));
    outputs(9322) <= not(layer4_outputs(2217));
    outputs(9323) <= not(layer4_outputs(2630));
    outputs(9324) <= not((layer4_outputs(3723)) xor (layer4_outputs(5618)));
    outputs(9325) <= (layer4_outputs(3604)) and not (layer4_outputs(9));
    outputs(9326) <= layer4_outputs(2565);
    outputs(9327) <= (layer4_outputs(2270)) xor (layer4_outputs(7173));
    outputs(9328) <= not(layer4_outputs(5068));
    outputs(9329) <= not(layer4_outputs(7728));
    outputs(9330) <= (layer4_outputs(2878)) xor (layer4_outputs(4345));
    outputs(9331) <= (layer4_outputs(1718)) xor (layer4_outputs(8910));
    outputs(9332) <= layer4_outputs(6572);
    outputs(9333) <= not((layer4_outputs(568)) xor (layer4_outputs(6390)));
    outputs(9334) <= layer4_outputs(9573);
    outputs(9335) <= not(layer4_outputs(4153));
    outputs(9336) <= (layer4_outputs(8622)) and not (layer4_outputs(9409));
    outputs(9337) <= not((layer4_outputs(8785)) xor (layer4_outputs(9234)));
    outputs(9338) <= (layer4_outputs(9285)) xor (layer4_outputs(8879));
    outputs(9339) <= (layer4_outputs(6125)) and not (layer4_outputs(5459));
    outputs(9340) <= (layer4_outputs(5815)) and not (layer4_outputs(1053));
    outputs(9341) <= not(layer4_outputs(3882));
    outputs(9342) <= layer4_outputs(8637);
    outputs(9343) <= (layer4_outputs(7774)) xor (layer4_outputs(9722));
    outputs(9344) <= not((layer4_outputs(8532)) or (layer4_outputs(1891)));
    outputs(9345) <= (layer4_outputs(600)) and (layer4_outputs(3456));
    outputs(9346) <= (layer4_outputs(849)) xor (layer4_outputs(1848));
    outputs(9347) <= (layer4_outputs(7904)) or (layer4_outputs(2570));
    outputs(9348) <= not(layer4_outputs(2469));
    outputs(9349) <= not(layer4_outputs(5454));
    outputs(9350) <= layer4_outputs(4738);
    outputs(9351) <= not((layer4_outputs(5685)) and (layer4_outputs(7686)));
    outputs(9352) <= layer4_outputs(2875);
    outputs(9353) <= not(layer4_outputs(7372));
    outputs(9354) <= not((layer4_outputs(283)) xor (layer4_outputs(7995)));
    outputs(9355) <= layer4_outputs(502);
    outputs(9356) <= not(layer4_outputs(2077));
    outputs(9357) <= not(layer4_outputs(2518)) or (layer4_outputs(9532));
    outputs(9358) <= layer4_outputs(748);
    outputs(9359) <= layer4_outputs(666);
    outputs(9360) <= (layer4_outputs(6988)) xor (layer4_outputs(8846));
    outputs(9361) <= not(layer4_outputs(1461));
    outputs(9362) <= not(layer4_outputs(7920));
    outputs(9363) <= not((layer4_outputs(1570)) xor (layer4_outputs(282)));
    outputs(9364) <= not(layer4_outputs(3640)) or (layer4_outputs(6939));
    outputs(9365) <= not(layer4_outputs(4024));
    outputs(9366) <= not((layer4_outputs(3482)) xor (layer4_outputs(4652)));
    outputs(9367) <= not(layer4_outputs(9500));
    outputs(9368) <= not((layer4_outputs(9410)) xor (layer4_outputs(3963)));
    outputs(9369) <= not(layer4_outputs(3880));
    outputs(9370) <= layer4_outputs(9520);
    outputs(9371) <= layer4_outputs(4295);
    outputs(9372) <= '1';
    outputs(9373) <= layer4_outputs(5666);
    outputs(9374) <= not(layer4_outputs(5115));
    outputs(9375) <= not(layer4_outputs(8060));
    outputs(9376) <= (layer4_outputs(3457)) or (layer4_outputs(386));
    outputs(9377) <= (layer4_outputs(9443)) or (layer4_outputs(6894));
    outputs(9378) <= (layer4_outputs(9429)) xor (layer4_outputs(5327));
    outputs(9379) <= not(layer4_outputs(5894));
    outputs(9380) <= layer4_outputs(7784);
    outputs(9381) <= (layer4_outputs(3942)) or (layer4_outputs(7184));
    outputs(9382) <= not((layer4_outputs(475)) xor (layer4_outputs(6022)));
    outputs(9383) <= not(layer4_outputs(6996));
    outputs(9384) <= (layer4_outputs(8949)) xor (layer4_outputs(9430));
    outputs(9385) <= not(layer4_outputs(8761));
    outputs(9386) <= layer4_outputs(3260);
    outputs(9387) <= not((layer4_outputs(9585)) xor (layer4_outputs(7184)));
    outputs(9388) <= not(layer4_outputs(3837));
    outputs(9389) <= (layer4_outputs(7351)) and not (layer4_outputs(7861));
    outputs(9390) <= (layer4_outputs(1304)) xor (layer4_outputs(4622));
    outputs(9391) <= layer4_outputs(7270);
    outputs(9392) <= layer4_outputs(9487);
    outputs(9393) <= not(layer4_outputs(278));
    outputs(9394) <= layer4_outputs(8554);
    outputs(9395) <= not(layer4_outputs(5181));
    outputs(9396) <= layer4_outputs(7397);
    outputs(9397) <= not(layer4_outputs(447));
    outputs(9398) <= (layer4_outputs(4597)) xor (layer4_outputs(7645));
    outputs(9399) <= not(layer4_outputs(6021)) or (layer4_outputs(8503));
    outputs(9400) <= not(layer4_outputs(4453));
    outputs(9401) <= (layer4_outputs(9798)) xor (layer4_outputs(8223));
    outputs(9402) <= layer4_outputs(2053);
    outputs(9403) <= layer4_outputs(7457);
    outputs(9404) <= (layer4_outputs(4176)) xor (layer4_outputs(4488));
    outputs(9405) <= not(layer4_outputs(6018)) or (layer4_outputs(9744));
    outputs(9406) <= not(layer4_outputs(174));
    outputs(9407) <= layer4_outputs(4710);
    outputs(9408) <= not(layer4_outputs(4179));
    outputs(9409) <= layer4_outputs(605);
    outputs(9410) <= layer4_outputs(4685);
    outputs(9411) <= layer4_outputs(6047);
    outputs(9412) <= layer4_outputs(7983);
    outputs(9413) <= not(layer4_outputs(4297));
    outputs(9414) <= layer4_outputs(4542);
    outputs(9415) <= not((layer4_outputs(8927)) xor (layer4_outputs(6983)));
    outputs(9416) <= not(layer4_outputs(4449));
    outputs(9417) <= layer4_outputs(8292);
    outputs(9418) <= (layer4_outputs(3595)) xor (layer4_outputs(9012));
    outputs(9419) <= not((layer4_outputs(862)) xor (layer4_outputs(939)));
    outputs(9420) <= layer4_outputs(8833);
    outputs(9421) <= (layer4_outputs(1488)) and not (layer4_outputs(857));
    outputs(9422) <= (layer4_outputs(8083)) and not (layer4_outputs(8566));
    outputs(9423) <= not(layer4_outputs(8275));
    outputs(9424) <= layer4_outputs(8674);
    outputs(9425) <= (layer4_outputs(1011)) and (layer4_outputs(997));
    outputs(9426) <= not(layer4_outputs(8597));
    outputs(9427) <= layer4_outputs(6532);
    outputs(9428) <= not((layer4_outputs(6234)) xor (layer4_outputs(8366)));
    outputs(9429) <= not((layer4_outputs(6553)) xor (layer4_outputs(2576)));
    outputs(9430) <= (layer4_outputs(8220)) or (layer4_outputs(1786));
    outputs(9431) <= (layer4_outputs(2912)) xor (layer4_outputs(729));
    outputs(9432) <= (layer4_outputs(7250)) xor (layer4_outputs(6556));
    outputs(9433) <= not((layer4_outputs(4942)) xor (layer4_outputs(7461)));
    outputs(9434) <= (layer4_outputs(4529)) and not (layer4_outputs(8791));
    outputs(9435) <= '0';
    outputs(9436) <= (layer4_outputs(46)) and not (layer4_outputs(2673));
    outputs(9437) <= not((layer4_outputs(1094)) xor (layer4_outputs(6279)));
    outputs(9438) <= not(layer4_outputs(6146));
    outputs(9439) <= (layer4_outputs(1754)) or (layer4_outputs(4647));
    outputs(9440) <= not(layer4_outputs(2521));
    outputs(9441) <= not(layer4_outputs(8626));
    outputs(9442) <= layer4_outputs(7507);
    outputs(9443) <= not(layer4_outputs(366));
    outputs(9444) <= not((layer4_outputs(8119)) xor (layer4_outputs(906)));
    outputs(9445) <= layer4_outputs(1893);
    outputs(9446) <= layer4_outputs(9015);
    outputs(9447) <= not((layer4_outputs(6436)) or (layer4_outputs(3713)));
    outputs(9448) <= (layer4_outputs(8542)) and (layer4_outputs(306));
    outputs(9449) <= '0';
    outputs(9450) <= not(layer4_outputs(2429));
    outputs(9451) <= (layer4_outputs(6587)) xor (layer4_outputs(2003));
    outputs(9452) <= (layer4_outputs(71)) xor (layer4_outputs(1193));
    outputs(9453) <= layer4_outputs(5891);
    outputs(9454) <= not((layer4_outputs(7636)) or (layer4_outputs(8567)));
    outputs(9455) <= layer4_outputs(8576);
    outputs(9456) <= not(layer4_outputs(520));
    outputs(9457) <= '1';
    outputs(9458) <= not(layer4_outputs(8006));
    outputs(9459) <= not(layer4_outputs(4790));
    outputs(9460) <= layer4_outputs(604);
    outputs(9461) <= not(layer4_outputs(4188));
    outputs(9462) <= layer4_outputs(1185);
    outputs(9463) <= layer4_outputs(10158);
    outputs(9464) <= not(layer4_outputs(7289));
    outputs(9465) <= not((layer4_outputs(3967)) or (layer4_outputs(2503)));
    outputs(9466) <= (layer4_outputs(5233)) and not (layer4_outputs(7220));
    outputs(9467) <= not((layer4_outputs(6719)) xor (layer4_outputs(1605)));
    outputs(9468) <= (layer4_outputs(6722)) xor (layer4_outputs(8744));
    outputs(9469) <= not(layer4_outputs(48));
    outputs(9470) <= not((layer4_outputs(2990)) xor (layer4_outputs(3243)));
    outputs(9471) <= layer4_outputs(3670);
    outputs(9472) <= layer4_outputs(5717);
    outputs(9473) <= layer4_outputs(2645);
    outputs(9474) <= not(layer4_outputs(3291));
    outputs(9475) <= not(layer4_outputs(231));
    outputs(9476) <= (layer4_outputs(5050)) xor (layer4_outputs(6578));
    outputs(9477) <= not(layer4_outputs(5045));
    outputs(9478) <= layer4_outputs(8792);
    outputs(9479) <= layer4_outputs(9338);
    outputs(9480) <= not((layer4_outputs(709)) xor (layer4_outputs(4913)));
    outputs(9481) <= layer4_outputs(546);
    outputs(9482) <= layer4_outputs(9727);
    outputs(9483) <= layer4_outputs(4044);
    outputs(9484) <= not(layer4_outputs(7717));
    outputs(9485) <= not(layer4_outputs(1911));
    outputs(9486) <= not((layer4_outputs(4799)) xor (layer4_outputs(6342)));
    outputs(9487) <= not(layer4_outputs(6515));
    outputs(9488) <= (layer4_outputs(10065)) xor (layer4_outputs(159));
    outputs(9489) <= not((layer4_outputs(2366)) xor (layer4_outputs(1835)));
    outputs(9490) <= (layer4_outputs(372)) xor (layer4_outputs(8003));
    outputs(9491) <= (layer4_outputs(2306)) and not (layer4_outputs(9290));
    outputs(9492) <= not((layer4_outputs(6224)) xor (layer4_outputs(9919)));
    outputs(9493) <= not(layer4_outputs(28));
    outputs(9494) <= layer4_outputs(4497);
    outputs(9495) <= not(layer4_outputs(1468));
    outputs(9496) <= not(layer4_outputs(6725));
    outputs(9497) <= (layer4_outputs(7322)) and not (layer4_outputs(4378));
    outputs(9498) <= (layer4_outputs(7547)) xor (layer4_outputs(8714));
    outputs(9499) <= not(layer4_outputs(8157));
    outputs(9500) <= not(layer4_outputs(7843));
    outputs(9501) <= not(layer4_outputs(1651));
    outputs(9502) <= (layer4_outputs(10139)) xor (layer4_outputs(9240));
    outputs(9503) <= layer4_outputs(9852);
    outputs(9504) <= (layer4_outputs(6358)) and not (layer4_outputs(3363));
    outputs(9505) <= not((layer4_outputs(4884)) xor (layer4_outputs(1642)));
    outputs(9506) <= not((layer4_outputs(3331)) xor (layer4_outputs(3740)));
    outputs(9507) <= '0';
    outputs(9508) <= layer4_outputs(5843);
    outputs(9509) <= not((layer4_outputs(6458)) xor (layer4_outputs(1589)));
    outputs(9510) <= not(layer4_outputs(5761)) or (layer4_outputs(6742));
    outputs(9511) <= layer4_outputs(4009);
    outputs(9512) <= not(layer4_outputs(3445));
    outputs(9513) <= not(layer4_outputs(9329));
    outputs(9514) <= not((layer4_outputs(3748)) xor (layer4_outputs(7884)));
    outputs(9515) <= not(layer4_outputs(866));
    outputs(9516) <= layer4_outputs(3324);
    outputs(9517) <= (layer4_outputs(7826)) xor (layer4_outputs(4912));
    outputs(9518) <= layer4_outputs(4769);
    outputs(9519) <= layer4_outputs(7010);
    outputs(9520) <= not((layer4_outputs(8554)) xor (layer4_outputs(9576)));
    outputs(9521) <= (layer4_outputs(252)) xor (layer4_outputs(3428));
    outputs(9522) <= not((layer4_outputs(7317)) xor (layer4_outputs(3408)));
    outputs(9523) <= not((layer4_outputs(1177)) or (layer4_outputs(8915)));
    outputs(9524) <= layer4_outputs(7624);
    outputs(9525) <= not(layer4_outputs(658)) or (layer4_outputs(8623));
    outputs(9526) <= not(layer4_outputs(7551)) or (layer4_outputs(9466));
    outputs(9527) <= not(layer4_outputs(4552));
    outputs(9528) <= layer4_outputs(8709);
    outputs(9529) <= (layer4_outputs(2002)) xor (layer4_outputs(677));
    outputs(9530) <= layer4_outputs(2654);
    outputs(9531) <= layer4_outputs(7895);
    outputs(9532) <= layer4_outputs(6651);
    outputs(9533) <= not(layer4_outputs(4061));
    outputs(9534) <= layer4_outputs(5266);
    outputs(9535) <= not((layer4_outputs(419)) xor (layer4_outputs(3684)));
    outputs(9536) <= not(layer4_outputs(7722));
    outputs(9537) <= layer4_outputs(2456);
    outputs(9538) <= layer4_outputs(5511);
    outputs(9539) <= not((layer4_outputs(3525)) xor (layer4_outputs(154)));
    outputs(9540) <= (layer4_outputs(2381)) and (layer4_outputs(3654));
    outputs(9541) <= (layer4_outputs(6610)) xor (layer4_outputs(5856));
    outputs(9542) <= (layer4_outputs(6986)) and (layer4_outputs(1720));
    outputs(9543) <= layer4_outputs(527);
    outputs(9544) <= layer4_outputs(445);
    outputs(9545) <= (layer4_outputs(7261)) or (layer4_outputs(7749));
    outputs(9546) <= layer4_outputs(3211);
    outputs(9547) <= layer4_outputs(789);
    outputs(9548) <= not((layer4_outputs(9022)) xor (layer4_outputs(1366)));
    outputs(9549) <= layer4_outputs(3312);
    outputs(9550) <= not((layer4_outputs(10237)) xor (layer4_outputs(6138)));
    outputs(9551) <= not(layer4_outputs(8113));
    outputs(9552) <= (layer4_outputs(5039)) and not (layer4_outputs(5789));
    outputs(9553) <= (layer4_outputs(1079)) and not (layer4_outputs(3240));
    outputs(9554) <= (layer4_outputs(2213)) xor (layer4_outputs(7981));
    outputs(9555) <= (layer4_outputs(7989)) xor (layer4_outputs(13));
    outputs(9556) <= layer4_outputs(109);
    outputs(9557) <= not(layer4_outputs(791));
    outputs(9558) <= layer4_outputs(6272);
    outputs(9559) <= not((layer4_outputs(665)) xor (layer4_outputs(901)));
    outputs(9560) <= not(layer4_outputs(9568));
    outputs(9561) <= (layer4_outputs(4022)) xor (layer4_outputs(366));
    outputs(9562) <= layer4_outputs(3803);
    outputs(9563) <= not(layer4_outputs(7429));
    outputs(9564) <= not(layer4_outputs(8227));
    outputs(9565) <= not((layer4_outputs(10027)) or (layer4_outputs(7610)));
    outputs(9566) <= (layer4_outputs(9527)) xor (layer4_outputs(3472));
    outputs(9567) <= not((layer4_outputs(4427)) xor (layer4_outputs(1826)));
    outputs(9568) <= (layer4_outputs(9462)) xor (layer4_outputs(5965));
    outputs(9569) <= layer4_outputs(5745);
    outputs(9570) <= layer4_outputs(3454);
    outputs(9571) <= layer4_outputs(9861);
    outputs(9572) <= layer4_outputs(7585);
    outputs(9573) <= not(layer4_outputs(6733));
    outputs(9574) <= layer4_outputs(5780);
    outputs(9575) <= not((layer4_outputs(7140)) xor (layer4_outputs(4839)));
    outputs(9576) <= not(layer4_outputs(6535));
    outputs(9577) <= not(layer4_outputs(2441)) or (layer4_outputs(7069));
    outputs(9578) <= layer4_outputs(6713);
    outputs(9579) <= (layer4_outputs(5015)) xor (layer4_outputs(9731));
    outputs(9580) <= not(layer4_outputs(5861));
    outputs(9581) <= not((layer4_outputs(146)) xor (layer4_outputs(8972)));
    outputs(9582) <= (layer4_outputs(4492)) xor (layer4_outputs(5923));
    outputs(9583) <= layer4_outputs(1533);
    outputs(9584) <= not((layer4_outputs(8014)) and (layer4_outputs(1363)));
    outputs(9585) <= layer4_outputs(6081);
    outputs(9586) <= layer4_outputs(2543);
    outputs(9587) <= layer4_outputs(674);
    outputs(9588) <= layer4_outputs(3248);
    outputs(9589) <= not(layer4_outputs(1450));
    outputs(9590) <= layer4_outputs(155);
    outputs(9591) <= not(layer4_outputs(7780));
    outputs(9592) <= (layer4_outputs(8284)) xor (layer4_outputs(238));
    outputs(9593) <= not(layer4_outputs(5620));
    outputs(9594) <= not((layer4_outputs(3606)) xor (layer4_outputs(1984)));
    outputs(9595) <= (layer4_outputs(5344)) and (layer4_outputs(154));
    outputs(9596) <= not(layer4_outputs(8097));
    outputs(9597) <= not(layer4_outputs(2405));
    outputs(9598) <= (layer4_outputs(8913)) xor (layer4_outputs(3398));
    outputs(9599) <= layer4_outputs(3966);
    outputs(9600) <= layer4_outputs(1572);
    outputs(9601) <= not(layer4_outputs(799));
    outputs(9602) <= layer4_outputs(6076);
    outputs(9603) <= layer4_outputs(1466);
    outputs(9604) <= (layer4_outputs(689)) xor (layer4_outputs(2347));
    outputs(9605) <= not(layer4_outputs(1070));
    outputs(9606) <= (layer4_outputs(6090)) and not (layer4_outputs(5323));
    outputs(9607) <= not(layer4_outputs(5557));
    outputs(9608) <= layer4_outputs(877);
    outputs(9609) <= not(layer4_outputs(4995)) or (layer4_outputs(598));
    outputs(9610) <= (layer4_outputs(4111)) xor (layer4_outputs(4836));
    outputs(9611) <= (layer4_outputs(9156)) and not (layer4_outputs(6019));
    outputs(9612) <= layer4_outputs(5871);
    outputs(9613) <= not(layer4_outputs(9621));
    outputs(9614) <= not(layer4_outputs(9637));
    outputs(9615) <= not(layer4_outputs(5053));
    outputs(9616) <= layer4_outputs(1945);
    outputs(9617) <= layer4_outputs(6283);
    outputs(9618) <= not((layer4_outputs(5929)) xor (layer4_outputs(4858)));
    outputs(9619) <= layer4_outputs(5338);
    outputs(9620) <= layer4_outputs(7418);
    outputs(9621) <= not(layer4_outputs(8348));
    outputs(9622) <= not((layer4_outputs(3998)) xor (layer4_outputs(3394)));
    outputs(9623) <= layer4_outputs(4931);
    outputs(9624) <= layer4_outputs(10190);
    outputs(9625) <= not(layer4_outputs(5554)) or (layer4_outputs(7897));
    outputs(9626) <= not(layer4_outputs(1611));
    outputs(9627) <= not(layer4_outputs(2129));
    outputs(9628) <= layer4_outputs(8736);
    outputs(9629) <= not(layer4_outputs(889));
    outputs(9630) <= not(layer4_outputs(2451));
    outputs(9631) <= not(layer4_outputs(2685));
    outputs(9632) <= layer4_outputs(9415);
    outputs(9633) <= (layer4_outputs(4782)) and not (layer4_outputs(1314));
    outputs(9634) <= layer4_outputs(1873);
    outputs(9635) <= not(layer4_outputs(6459));
    outputs(9636) <= (layer4_outputs(9082)) xor (layer4_outputs(8509));
    outputs(9637) <= not(layer4_outputs(5419));
    outputs(9638) <= not(layer4_outputs(9400));
    outputs(9639) <= not(layer4_outputs(735));
    outputs(9640) <= not((layer4_outputs(4286)) xor (layer4_outputs(8502)));
    outputs(9641) <= (layer4_outputs(3878)) xor (layer4_outputs(8840));
    outputs(9642) <= not((layer4_outputs(6304)) xor (layer4_outputs(3341)));
    outputs(9643) <= (layer4_outputs(8715)) and not (layer4_outputs(6335));
    outputs(9644) <= layer4_outputs(3937);
    outputs(9645) <= not(layer4_outputs(349));
    outputs(9646) <= not((layer4_outputs(2651)) xor (layer4_outputs(389)));
    outputs(9647) <= not(layer4_outputs(9286));
    outputs(9648) <= not(layer4_outputs(9997));
    outputs(9649) <= not(layer4_outputs(1330));
    outputs(9650) <= layer4_outputs(5567);
    outputs(9651) <= not(layer4_outputs(1396));
    outputs(9652) <= layer4_outputs(3061);
    outputs(9653) <= layer4_outputs(7056);
    outputs(9654) <= layer4_outputs(7684);
    outputs(9655) <= not(layer4_outputs(3933));
    outputs(9656) <= not((layer4_outputs(938)) xor (layer4_outputs(3348)));
    outputs(9657) <= (layer4_outputs(3938)) xor (layer4_outputs(9697));
    outputs(9658) <= not(layer4_outputs(2973));
    outputs(9659) <= (layer4_outputs(10203)) xor (layer4_outputs(9073));
    outputs(9660) <= not(layer4_outputs(1681));
    outputs(9661) <= not(layer4_outputs(88));
    outputs(9662) <= layer4_outputs(10191);
    outputs(9663) <= layer4_outputs(4396);
    outputs(9664) <= layer4_outputs(5958);
    outputs(9665) <= not(layer4_outputs(4930)) or (layer4_outputs(2520));
    outputs(9666) <= (layer4_outputs(4789)) xor (layer4_outputs(2166));
    outputs(9667) <= (layer4_outputs(9428)) or (layer4_outputs(3430));
    outputs(9668) <= not((layer4_outputs(1018)) xor (layer4_outputs(1592)));
    outputs(9669) <= layer4_outputs(5664);
    outputs(9670) <= layer4_outputs(5171);
    outputs(9671) <= not(layer4_outputs(1692));
    outputs(9672) <= layer4_outputs(5134);
    outputs(9673) <= (layer4_outputs(5277)) xor (layer4_outputs(5516));
    outputs(9674) <= not(layer4_outputs(7060));
    outputs(9675) <= (layer4_outputs(4463)) xor (layer4_outputs(3087));
    outputs(9676) <= not(layer4_outputs(2507));
    outputs(9677) <= not((layer4_outputs(1504)) xor (layer4_outputs(9761)));
    outputs(9678) <= not(layer4_outputs(547));
    outputs(9679) <= (layer4_outputs(6074)) xor (layer4_outputs(4022));
    outputs(9680) <= not((layer4_outputs(5165)) xor (layer4_outputs(7616)));
    outputs(9681) <= not((layer4_outputs(258)) xor (layer4_outputs(4214)));
    outputs(9682) <= (layer4_outputs(9720)) and not (layer4_outputs(6517));
    outputs(9683) <= not(layer4_outputs(4142));
    outputs(9684) <= not(layer4_outputs(10014));
    outputs(9685) <= not(layer4_outputs(6616));
    outputs(9686) <= not((layer4_outputs(9680)) xor (layer4_outputs(1582)));
    outputs(9687) <= layer4_outputs(1711);
    outputs(9688) <= not(layer4_outputs(9232));
    outputs(9689) <= not((layer4_outputs(810)) xor (layer4_outputs(6543)));
    outputs(9690) <= not((layer4_outputs(7347)) xor (layer4_outputs(7547)));
    outputs(9691) <= layer4_outputs(6992);
    outputs(9692) <= not(layer4_outputs(5562));
    outputs(9693) <= layer4_outputs(6971);
    outputs(9694) <= not(layer4_outputs(3496));
    outputs(9695) <= not(layer4_outputs(1258));
    outputs(9696) <= (layer4_outputs(1576)) and not (layer4_outputs(8759));
    outputs(9697) <= not(layer4_outputs(1238));
    outputs(9698) <= layer4_outputs(6780);
    outputs(9699) <= (layer4_outputs(9183)) xor (layer4_outputs(1873));
    outputs(9700) <= not(layer4_outputs(5712));
    outputs(9701) <= layer4_outputs(6955);
    outputs(9702) <= layer4_outputs(6005);
    outputs(9703) <= layer4_outputs(9785);
    outputs(9704) <= not(layer4_outputs(7764));
    outputs(9705) <= layer4_outputs(6832);
    outputs(9706) <= not((layer4_outputs(3596)) or (layer4_outputs(4411)));
    outputs(9707) <= (layer4_outputs(6818)) xor (layer4_outputs(3050));
    outputs(9708) <= not((layer4_outputs(5347)) xor (layer4_outputs(9783)));
    outputs(9709) <= not(layer4_outputs(4965));
    outputs(9710) <= not((layer4_outputs(10001)) or (layer4_outputs(7997)));
    outputs(9711) <= not(layer4_outputs(1457));
    outputs(9712) <= layer4_outputs(2109);
    outputs(9713) <= not((layer4_outputs(7260)) xor (layer4_outputs(5250)));
    outputs(9714) <= layer4_outputs(8573);
    outputs(9715) <= (layer4_outputs(5018)) and (layer4_outputs(4484));
    outputs(9716) <= (layer4_outputs(493)) xor (layer4_outputs(6907));
    outputs(9717) <= (layer4_outputs(10038)) and not (layer4_outputs(8400));
    outputs(9718) <= not((layer4_outputs(2437)) xor (layer4_outputs(8881)));
    outputs(9719) <= not((layer4_outputs(2739)) xor (layer4_outputs(5812)));
    outputs(9720) <= not(layer4_outputs(4875));
    outputs(9721) <= layer4_outputs(3487);
    outputs(9722) <= not(layer4_outputs(9420));
    outputs(9723) <= layer4_outputs(2775);
    outputs(9724) <= (layer4_outputs(2339)) xor (layer4_outputs(1365));
    outputs(9725) <= (layer4_outputs(5442)) xor (layer4_outputs(8467));
    outputs(9726) <= not(layer4_outputs(4258));
    outputs(9727) <= not(layer4_outputs(58));
    outputs(9728) <= layer4_outputs(2361);
    outputs(9729) <= not(layer4_outputs(1918));
    outputs(9730) <= not(layer4_outputs(805));
    outputs(9731) <= (layer4_outputs(583)) or (layer4_outputs(1439));
    outputs(9732) <= not(layer4_outputs(5944));
    outputs(9733) <= not(layer4_outputs(3101));
    outputs(9734) <= not(layer4_outputs(3335));
    outputs(9735) <= layer4_outputs(5561);
    outputs(9736) <= layer4_outputs(10033);
    outputs(9737) <= not(layer4_outputs(8765));
    outputs(9738) <= layer4_outputs(6681);
    outputs(9739) <= not(layer4_outputs(7125));
    outputs(9740) <= not((layer4_outputs(1381)) and (layer4_outputs(1838)));
    outputs(9741) <= not(layer4_outputs(4525));
    outputs(9742) <= not((layer4_outputs(7833)) xor (layer4_outputs(6227)));
    outputs(9743) <= not(layer4_outputs(1305));
    outputs(9744) <= not((layer4_outputs(3051)) xor (layer4_outputs(7237)));
    outputs(9745) <= (layer4_outputs(10140)) and not (layer4_outputs(1179));
    outputs(9746) <= not(layer4_outputs(7160)) or (layer4_outputs(7014));
    outputs(9747) <= layer4_outputs(5727);
    outputs(9748) <= layer4_outputs(643);
    outputs(9749) <= not(layer4_outputs(8031));
    outputs(9750) <= (layer4_outputs(4670)) xor (layer4_outputs(3959));
    outputs(9751) <= not((layer4_outputs(7527)) or (layer4_outputs(8196)));
    outputs(9752) <= not(layer4_outputs(7185));
    outputs(9753) <= not(layer4_outputs(5600)) or (layer4_outputs(6644));
    outputs(9754) <= not(layer4_outputs(3545));
    outputs(9755) <= not(layer4_outputs(3223));
    outputs(9756) <= not(layer4_outputs(3145));
    outputs(9757) <= not(layer4_outputs(4037));
    outputs(9758) <= layer4_outputs(6095);
    outputs(9759) <= layer4_outputs(1895);
    outputs(9760) <= not((layer4_outputs(3767)) xor (layer4_outputs(6617)));
    outputs(9761) <= not(layer4_outputs(5149));
    outputs(9762) <= not(layer4_outputs(7909));
    outputs(9763) <= not(layer4_outputs(8945));
    outputs(9764) <= layer4_outputs(2513);
    outputs(9765) <= not((layer4_outputs(8083)) xor (layer4_outputs(269)));
    outputs(9766) <= layer4_outputs(9040);
    outputs(9767) <= layer4_outputs(5403);
    outputs(9768) <= not((layer4_outputs(5364)) xor (layer4_outputs(4648)));
    outputs(9769) <= layer4_outputs(8861);
    outputs(9770) <= (layer4_outputs(2573)) xor (layer4_outputs(5432));
    outputs(9771) <= not(layer4_outputs(5353));
    outputs(9772) <= not(layer4_outputs(4818));
    outputs(9773) <= not(layer4_outputs(1331));
    outputs(9774) <= not(layer4_outputs(9644));
    outputs(9775) <= not((layer4_outputs(4284)) xor (layer4_outputs(3820)));
    outputs(9776) <= not((layer4_outputs(5985)) xor (layer4_outputs(788)));
    outputs(9777) <= not((layer4_outputs(3161)) xor (layer4_outputs(3164)));
    outputs(9778) <= not(layer4_outputs(1875));
    outputs(9779) <= not((layer4_outputs(8485)) xor (layer4_outputs(10074)));
    outputs(9780) <= not(layer4_outputs(5637));
    outputs(9781) <= not((layer4_outputs(7731)) xor (layer4_outputs(5617)));
    outputs(9782) <= (layer4_outputs(6267)) and not (layer4_outputs(6839));
    outputs(9783) <= not((layer4_outputs(1031)) or (layer4_outputs(5805)));
    outputs(9784) <= (layer4_outputs(7694)) xor (layer4_outputs(5302));
    outputs(9785) <= (layer4_outputs(841)) and not (layer4_outputs(9851));
    outputs(9786) <= layer4_outputs(4694);
    outputs(9787) <= not(layer4_outputs(9051));
    outputs(9788) <= layer4_outputs(4352);
    outputs(9789) <= (layer4_outputs(8398)) xor (layer4_outputs(7496));
    outputs(9790) <= layer4_outputs(7299);
    outputs(9791) <= (layer4_outputs(4471)) xor (layer4_outputs(10079));
    outputs(9792) <= layer4_outputs(333);
    outputs(9793) <= not((layer4_outputs(5283)) xor (layer4_outputs(8114)));
    outputs(9794) <= not((layer4_outputs(3945)) or (layer4_outputs(4700)));
    outputs(9795) <= (layer4_outputs(828)) or (layer4_outputs(3639));
    outputs(9796) <= layer4_outputs(1550);
    outputs(9797) <= not(layer4_outputs(2581));
    outputs(9798) <= not((layer4_outputs(7197)) xor (layer4_outputs(8863)));
    outputs(9799) <= (layer4_outputs(6503)) xor (layer4_outputs(8498));
    outputs(9800) <= layer4_outputs(5352);
    outputs(9801) <= (layer4_outputs(8665)) xor (layer4_outputs(6032));
    outputs(9802) <= not(layer4_outputs(1320));
    outputs(9803) <= layer4_outputs(1778);
    outputs(9804) <= (layer4_outputs(6239)) xor (layer4_outputs(5153));
    outputs(9805) <= not(layer4_outputs(1433)) or (layer4_outputs(9330));
    outputs(9806) <= not((layer4_outputs(3114)) or (layer4_outputs(7568)));
    outputs(9807) <= not(layer4_outputs(6153));
    outputs(9808) <= not(layer4_outputs(5104));
    outputs(9809) <= not(layer4_outputs(337));
    outputs(9810) <= not((layer4_outputs(2919)) xor (layer4_outputs(3699)));
    outputs(9811) <= (layer4_outputs(10231)) or (layer4_outputs(2392));
    outputs(9812) <= not(layer4_outputs(6562));
    outputs(9813) <= layer4_outputs(5330);
    outputs(9814) <= not(layer4_outputs(10205));
    outputs(9815) <= '1';
    outputs(9816) <= not(layer4_outputs(3052));
    outputs(9817) <= (layer4_outputs(7530)) xor (layer4_outputs(10139));
    outputs(9818) <= layer4_outputs(6300);
    outputs(9819) <= not(layer4_outputs(1624));
    outputs(9820) <= not(layer4_outputs(1882));
    outputs(9821) <= layer4_outputs(8764);
    outputs(9822) <= layer4_outputs(8019);
    outputs(9823) <= not(layer4_outputs(7539));
    outputs(9824) <= not(layer4_outputs(1933));
    outputs(9825) <= layer4_outputs(6567);
    outputs(9826) <= not((layer4_outputs(6070)) xor (layer4_outputs(1083)));
    outputs(9827) <= (layer4_outputs(6637)) and not (layer4_outputs(4115));
    outputs(9828) <= (layer4_outputs(10223)) xor (layer4_outputs(3679));
    outputs(9829) <= (layer4_outputs(4076)) or (layer4_outputs(9924));
    outputs(9830) <= (layer4_outputs(3510)) or (layer4_outputs(1093));
    outputs(9831) <= layer4_outputs(1899);
    outputs(9832) <= layer4_outputs(9466);
    outputs(9833) <= not((layer4_outputs(881)) xor (layer4_outputs(3043)));
    outputs(9834) <= (layer4_outputs(6234)) xor (layer4_outputs(8213));
    outputs(9835) <= not((layer4_outputs(7572)) xor (layer4_outputs(4632)));
    outputs(9836) <= not(layer4_outputs(9699));
    outputs(9837) <= layer4_outputs(8669);
    outputs(9838) <= (layer4_outputs(8369)) and (layer4_outputs(3648));
    outputs(9839) <= not(layer4_outputs(4531));
    outputs(9840) <= not(layer4_outputs(4545));
    outputs(9841) <= (layer4_outputs(2107)) xor (layer4_outputs(5566));
    outputs(9842) <= layer4_outputs(5728);
    outputs(9843) <= not(layer4_outputs(7721)) or (layer4_outputs(2789));
    outputs(9844) <= layer4_outputs(1534);
    outputs(9845) <= not(layer4_outputs(1147));
    outputs(9846) <= (layer4_outputs(20)) xor (layer4_outputs(3915));
    outputs(9847) <= not((layer4_outputs(8027)) xor (layer4_outputs(4651)));
    outputs(9848) <= layer4_outputs(5728);
    outputs(9849) <= not(layer4_outputs(7769));
    outputs(9850) <= layer4_outputs(4223);
    outputs(9851) <= not(layer4_outputs(3935));
    outputs(9852) <= not((layer4_outputs(9245)) or (layer4_outputs(8602)));
    outputs(9853) <= layer4_outputs(1047);
    outputs(9854) <= not(layer4_outputs(6108));
    outputs(9855) <= not(layer4_outputs(5921));
    outputs(9856) <= not((layer4_outputs(4190)) xor (layer4_outputs(3971)));
    outputs(9857) <= not((layer4_outputs(4000)) xor (layer4_outputs(8300)));
    outputs(9858) <= layer4_outputs(9052);
    outputs(9859) <= not(layer4_outputs(2593));
    outputs(9860) <= not(layer4_outputs(5275));
    outputs(9861) <= (layer4_outputs(168)) xor (layer4_outputs(1025));
    outputs(9862) <= layer4_outputs(7112);
    outputs(9863) <= layer4_outputs(6281);
    outputs(9864) <= not((layer4_outputs(4730)) xor (layer4_outputs(5777)));
    outputs(9865) <= (layer4_outputs(9676)) and not (layer4_outputs(3978));
    outputs(9866) <= not(layer4_outputs(8770));
    outputs(9867) <= layer4_outputs(8450);
    outputs(9868) <= (layer4_outputs(5331)) xor (layer4_outputs(6822));
    outputs(9869) <= (layer4_outputs(4895)) and not (layer4_outputs(1099));
    outputs(9870) <= not(layer4_outputs(7412));
    outputs(9871) <= not(layer4_outputs(3301));
    outputs(9872) <= not((layer4_outputs(4536)) or (layer4_outputs(8082)));
    outputs(9873) <= not(layer4_outputs(9496));
    outputs(9874) <= layer4_outputs(7979);
    outputs(9875) <= layer4_outputs(4575);
    outputs(9876) <= (layer4_outputs(3156)) xor (layer4_outputs(5112));
    outputs(9877) <= not(layer4_outputs(8759));
    outputs(9878) <= (layer4_outputs(1290)) xor (layer4_outputs(1401));
    outputs(9879) <= not(layer4_outputs(2102));
    outputs(9880) <= not(layer4_outputs(1642));
    outputs(9881) <= (layer4_outputs(2728)) and not (layer4_outputs(5046));
    outputs(9882) <= not(layer4_outputs(8850));
    outputs(9883) <= not(layer4_outputs(8129));
    outputs(9884) <= not(layer4_outputs(5720));
    outputs(9885) <= (layer4_outputs(4529)) or (layer4_outputs(10165));
    outputs(9886) <= layer4_outputs(8738);
    outputs(9887) <= (layer4_outputs(2304)) and (layer4_outputs(3417));
    outputs(9888) <= (layer4_outputs(4033)) xor (layer4_outputs(512));
    outputs(9889) <= not((layer4_outputs(3417)) xor (layer4_outputs(2734)));
    outputs(9890) <= not(layer4_outputs(10134));
    outputs(9891) <= not(layer4_outputs(7080));
    outputs(9892) <= (layer4_outputs(664)) xor (layer4_outputs(9886));
    outputs(9893) <= layer4_outputs(1209);
    outputs(9894) <= not(layer4_outputs(7501));
    outputs(9895) <= layer4_outputs(4868);
    outputs(9896) <= not((layer4_outputs(9145)) xor (layer4_outputs(2738)));
    outputs(9897) <= layer4_outputs(6673);
    outputs(9898) <= not(layer4_outputs(6903));
    outputs(9899) <= (layer4_outputs(3514)) xor (layer4_outputs(7383));
    outputs(9900) <= (layer4_outputs(9796)) xor (layer4_outputs(978));
    outputs(9901) <= (layer4_outputs(4479)) xor (layer4_outputs(4631));
    outputs(9902) <= not(layer4_outputs(1668));
    outputs(9903) <= not((layer4_outputs(3599)) xor (layer4_outputs(9474)));
    outputs(9904) <= not((layer4_outputs(4264)) and (layer4_outputs(8204)));
    outputs(9905) <= layer4_outputs(2744);
    outputs(9906) <= layer4_outputs(4729);
    outputs(9907) <= (layer4_outputs(5857)) or (layer4_outputs(338));
    outputs(9908) <= not((layer4_outputs(1990)) xor (layer4_outputs(637)));
    outputs(9909) <= not(layer4_outputs(6378));
    outputs(9910) <= layer4_outputs(3058);
    outputs(9911) <= (layer4_outputs(6055)) xor (layer4_outputs(1862));
    outputs(9912) <= not(layer4_outputs(3439));
    outputs(9913) <= not(layer4_outputs(9185));
    outputs(9914) <= not((layer4_outputs(4600)) and (layer4_outputs(5505)));
    outputs(9915) <= not(layer4_outputs(7185));
    outputs(9916) <= not((layer4_outputs(1500)) xor (layer4_outputs(4828)));
    outputs(9917) <= not((layer4_outputs(2310)) xor (layer4_outputs(9225)));
    outputs(9918) <= layer4_outputs(8541);
    outputs(9919) <= not(layer4_outputs(7412));
    outputs(9920) <= (layer4_outputs(6011)) xor (layer4_outputs(10049));
    outputs(9921) <= layer4_outputs(5775);
    outputs(9922) <= not(layer4_outputs(4465));
    outputs(9923) <= (layer4_outputs(1247)) and (layer4_outputs(5523));
    outputs(9924) <= (layer4_outputs(8032)) xor (layer4_outputs(2508));
    outputs(9925) <= not(layer4_outputs(768)) or (layer4_outputs(7561));
    outputs(9926) <= not((layer4_outputs(1741)) or (layer4_outputs(7856)));
    outputs(9927) <= (layer4_outputs(8025)) xor (layer4_outputs(4877));
    outputs(9928) <= layer4_outputs(8081);
    outputs(9929) <= (layer4_outputs(673)) xor (layer4_outputs(5410));
    outputs(9930) <= not(layer4_outputs(3382));
    outputs(9931) <= not((layer4_outputs(4331)) xor (layer4_outputs(3528)));
    outputs(9932) <= layer4_outputs(4859);
    outputs(9933) <= (layer4_outputs(2195)) xor (layer4_outputs(8354));
    outputs(9934) <= not(layer4_outputs(482));
    outputs(9935) <= not(layer4_outputs(203));
    outputs(9936) <= not((layer4_outputs(5445)) xor (layer4_outputs(7415)));
    outputs(9937) <= (layer4_outputs(6045)) xor (layer4_outputs(479));
    outputs(9938) <= not((layer4_outputs(9085)) xor (layer4_outputs(8679)));
    outputs(9939) <= (layer4_outputs(4866)) and not (layer4_outputs(50));
    outputs(9940) <= '0';
    outputs(9941) <= (layer4_outputs(5749)) and (layer4_outputs(1529));
    outputs(9942) <= not(layer4_outputs(1692));
    outputs(9943) <= not(layer4_outputs(3066));
    outputs(9944) <= layer4_outputs(6191);
    outputs(9945) <= not((layer4_outputs(4122)) and (layer4_outputs(2477)));
    outputs(9946) <= not((layer4_outputs(963)) xor (layer4_outputs(6874)));
    outputs(9947) <= not(layer4_outputs(1627));
    outputs(9948) <= not((layer4_outputs(9662)) xor (layer4_outputs(8556)));
    outputs(9949) <= not((layer4_outputs(1826)) or (layer4_outputs(7382)));
    outputs(9950) <= not(layer4_outputs(7843));
    outputs(9951) <= not(layer4_outputs(190)) or (layer4_outputs(7257));
    outputs(9952) <= not((layer4_outputs(684)) or (layer4_outputs(206)));
    outputs(9953) <= (layer4_outputs(5195)) and (layer4_outputs(4343));
    outputs(9954) <= layer4_outputs(5282);
    outputs(9955) <= not(layer4_outputs(8101));
    outputs(9956) <= not(layer4_outputs(6696));
    outputs(9957) <= layer4_outputs(8343);
    outputs(9958) <= not((layer4_outputs(3046)) xor (layer4_outputs(4047)));
    outputs(9959) <= not(layer4_outputs(7061));
    outputs(9960) <= not(layer4_outputs(8723)) or (layer4_outputs(2936));
    outputs(9961) <= (layer4_outputs(3889)) xor (layer4_outputs(7318));
    outputs(9962) <= not(layer4_outputs(5896));
    outputs(9963) <= layer4_outputs(2216);
    outputs(9964) <= not((layer4_outputs(10164)) or (layer4_outputs(1913)));
    outputs(9965) <= not(layer4_outputs(5407));
    outputs(9966) <= (layer4_outputs(611)) xor (layer4_outputs(5441));
    outputs(9967) <= (layer4_outputs(591)) xor (layer4_outputs(7541));
    outputs(9968) <= not(layer4_outputs(890));
    outputs(9969) <= layer4_outputs(9711);
    outputs(9970) <= not((layer4_outputs(2735)) xor (layer4_outputs(1891)));
    outputs(9971) <= not(layer4_outputs(81));
    outputs(9972) <= (layer4_outputs(1612)) or (layer4_outputs(10133));
    outputs(9973) <= (layer4_outputs(6432)) xor (layer4_outputs(9290));
    outputs(9974) <= layer4_outputs(8716);
    outputs(9975) <= layer4_outputs(9497);
    outputs(9976) <= not((layer4_outputs(9641)) xor (layer4_outputs(1655)));
    outputs(9977) <= not((layer4_outputs(4063)) and (layer4_outputs(6196)));
    outputs(9978) <= layer4_outputs(4383);
    outputs(9979) <= not((layer4_outputs(3641)) xor (layer4_outputs(8931)));
    outputs(9980) <= layer4_outputs(9147);
    outputs(9981) <= not((layer4_outputs(2708)) or (layer4_outputs(8519)));
    outputs(9982) <= not(layer4_outputs(9060));
    outputs(9983) <= not(layer4_outputs(7281)) or (layer4_outputs(1822));
    outputs(9984) <= (layer4_outputs(5564)) xor (layer4_outputs(1022));
    outputs(9985) <= not(layer4_outputs(1038));
    outputs(9986) <= not(layer4_outputs(2630));
    outputs(9987) <= layer4_outputs(448);
    outputs(9988) <= (layer4_outputs(7304)) xor (layer4_outputs(5852));
    outputs(9989) <= not((layer4_outputs(8600)) xor (layer4_outputs(4001)));
    outputs(9990) <= (layer4_outputs(8688)) xor (layer4_outputs(427));
    outputs(9991) <= (layer4_outputs(113)) and not (layer4_outputs(8515));
    outputs(9992) <= layer4_outputs(8788);
    outputs(9993) <= not(layer4_outputs(591));
    outputs(9994) <= not(layer4_outputs(186)) or (layer4_outputs(7991));
    outputs(9995) <= not((layer4_outputs(6861)) xor (layer4_outputs(5674)));
    outputs(9996) <= not(layer4_outputs(2057));
    outputs(9997) <= layer4_outputs(3375);
    outputs(9998) <= not(layer4_outputs(2583));
    outputs(9999) <= (layer4_outputs(10008)) and (layer4_outputs(1247));
    outputs(10000) <= (layer4_outputs(1183)) and not (layer4_outputs(582));
    outputs(10001) <= not(layer4_outputs(1959));
    outputs(10002) <= layer4_outputs(2703);
    outputs(10003) <= not((layer4_outputs(10202)) xor (layer4_outputs(4769)));
    outputs(10004) <= (layer4_outputs(9217)) xor (layer4_outputs(9867));
    outputs(10005) <= layer4_outputs(3239);
    outputs(10006) <= (layer4_outputs(7800)) xor (layer4_outputs(9098));
    outputs(10007) <= not(layer4_outputs(2174));
    outputs(10008) <= not(layer4_outputs(8053));
    outputs(10009) <= layer4_outputs(659);
    outputs(10010) <= layer4_outputs(7225);
    outputs(10011) <= not(layer4_outputs(149));
    outputs(10012) <= not(layer4_outputs(6236)) or (layer4_outputs(4308));
    outputs(10013) <= not((layer4_outputs(9021)) xor (layer4_outputs(5126)));
    outputs(10014) <= not(layer4_outputs(3393));
    outputs(10015) <= layer4_outputs(3157);
    outputs(10016) <= not(layer4_outputs(2251));
    outputs(10017) <= layer4_outputs(6132);
    outputs(10018) <= not((layer4_outputs(8873)) xor (layer4_outputs(5359)));
    outputs(10019) <= (layer4_outputs(8872)) and (layer4_outputs(675));
    outputs(10020) <= not(layer4_outputs(9490));
    outputs(10021) <= not(layer4_outputs(6516));
    outputs(10022) <= not(layer4_outputs(2537));
    outputs(10023) <= not(layer4_outputs(7672));
    outputs(10024) <= not((layer4_outputs(6813)) or (layer4_outputs(7369)));
    outputs(10025) <= not(layer4_outputs(5975));
    outputs(10026) <= not((layer4_outputs(7586)) xor (layer4_outputs(4588)));
    outputs(10027) <= not(layer4_outputs(4584));
    outputs(10028) <= not(layer4_outputs(4477));
    outputs(10029) <= (layer4_outputs(6684)) or (layer4_outputs(415));
    outputs(10030) <= layer4_outputs(6011);
    outputs(10031) <= not(layer4_outputs(5124));
    outputs(10032) <= layer4_outputs(298);
    outputs(10033) <= not(layer4_outputs(7903));
    outputs(10034) <= not(layer4_outputs(5424));
    outputs(10035) <= not(layer4_outputs(10150)) or (layer4_outputs(5396));
    outputs(10036) <= not((layer4_outputs(3551)) xor (layer4_outputs(7742)));
    outputs(10037) <= (layer4_outputs(9444)) xor (layer4_outputs(4821));
    outputs(10038) <= (layer4_outputs(555)) and not (layer4_outputs(4030));
    outputs(10039) <= not((layer4_outputs(1067)) xor (layer4_outputs(1508)));
    outputs(10040) <= (layer4_outputs(9727)) xor (layer4_outputs(5702));
    outputs(10041) <= not(layer4_outputs(1941));
    outputs(10042) <= not(layer4_outputs(7133)) or (layer4_outputs(5910));
    outputs(10043) <= not((layer4_outputs(2479)) xor (layer4_outputs(1456)));
    outputs(10044) <= (layer4_outputs(3781)) xor (layer4_outputs(4509));
    outputs(10045) <= not((layer4_outputs(3657)) xor (layer4_outputs(7222)));
    outputs(10046) <= not((layer4_outputs(4387)) xor (layer4_outputs(3020)));
    outputs(10047) <= not(layer4_outputs(3884));
    outputs(10048) <= (layer4_outputs(6708)) xor (layer4_outputs(7515));
    outputs(10049) <= (layer4_outputs(6564)) xor (layer4_outputs(7211));
    outputs(10050) <= layer4_outputs(1044);
    outputs(10051) <= not(layer4_outputs(2615)) or (layer4_outputs(4966));
    outputs(10052) <= not(layer4_outputs(7882)) or (layer4_outputs(6283));
    outputs(10053) <= (layer4_outputs(5361)) or (layer4_outputs(4605));
    outputs(10054) <= not(layer4_outputs(129));
    outputs(10055) <= not(layer4_outputs(1076));
    outputs(10056) <= not(layer4_outputs(1791));
    outputs(10057) <= not((layer4_outputs(9033)) xor (layer4_outputs(8228)));
    outputs(10058) <= (layer4_outputs(6904)) xor (layer4_outputs(7882));
    outputs(10059) <= not(layer4_outputs(121));
    outputs(10060) <= layer4_outputs(9868);
    outputs(10061) <= layer4_outputs(2802);
    outputs(10062) <= not((layer4_outputs(10088)) xor (layer4_outputs(228)));
    outputs(10063) <= layer4_outputs(4414);
    outputs(10064) <= (layer4_outputs(1555)) and not (layer4_outputs(3480));
    outputs(10065) <= (layer4_outputs(4555)) xor (layer4_outputs(6334));
    outputs(10066) <= (layer4_outputs(3974)) and not (layer4_outputs(8087));
    outputs(10067) <= not(layer4_outputs(8036));
    outputs(10068) <= not(layer4_outputs(255));
    outputs(10069) <= not(layer4_outputs(6101));
    outputs(10070) <= not((layer4_outputs(9171)) xor (layer4_outputs(4586)));
    outputs(10071) <= not((layer4_outputs(9954)) xor (layer4_outputs(9350)));
    outputs(10072) <= (layer4_outputs(4665)) xor (layer4_outputs(6212));
    outputs(10073) <= not(layer4_outputs(1338));
    outputs(10074) <= (layer4_outputs(2561)) xor (layer4_outputs(2408));
    outputs(10075) <= not(layer4_outputs(9456));
    outputs(10076) <= not((layer4_outputs(4132)) xor (layer4_outputs(3489)));
    outputs(10077) <= layer4_outputs(9944);
    outputs(10078) <= not(layer4_outputs(2521));
    outputs(10079) <= layer4_outputs(10197);
    outputs(10080) <= not(layer4_outputs(291));
    outputs(10081) <= not((layer4_outputs(3448)) xor (layer4_outputs(2043)));
    outputs(10082) <= layer4_outputs(3947);
    outputs(10083) <= not(layer4_outputs(9394));
    outputs(10084) <= not(layer4_outputs(9383));
    outputs(10085) <= not(layer4_outputs(6957)) or (layer4_outputs(5623));
    outputs(10086) <= not((layer4_outputs(2638)) xor (layer4_outputs(3719)));
    outputs(10087) <= not((layer4_outputs(5200)) xor (layer4_outputs(3041)));
    outputs(10088) <= not(layer4_outputs(268));
    outputs(10089) <= not(layer4_outputs(9020)) or (layer4_outputs(8586));
    outputs(10090) <= not(layer4_outputs(6188));
    outputs(10091) <= layer4_outputs(2471);
    outputs(10092) <= (layer4_outputs(5820)) xor (layer4_outputs(3687));
    outputs(10093) <= layer4_outputs(2449);
    outputs(10094) <= not(layer4_outputs(222));
    outputs(10095) <= (layer4_outputs(7174)) xor (layer4_outputs(4117));
    outputs(10096) <= layer4_outputs(8049);
    outputs(10097) <= (layer4_outputs(8980)) xor (layer4_outputs(1138));
    outputs(10098) <= (layer4_outputs(501)) xor (layer4_outputs(4294));
    outputs(10099) <= not(layer4_outputs(7869));
    outputs(10100) <= layer4_outputs(5074);
    outputs(10101) <= (layer4_outputs(9141)) xor (layer4_outputs(7479));
    outputs(10102) <= not(layer4_outputs(3288));
    outputs(10103) <= not(layer4_outputs(299));
    outputs(10104) <= not((layer4_outputs(2205)) xor (layer4_outputs(287)));
    outputs(10105) <= not(layer4_outputs(373));
    outputs(10106) <= not(layer4_outputs(9192));
    outputs(10107) <= not(layer4_outputs(7876));
    outputs(10108) <= not(layer4_outputs(6389)) or (layer4_outputs(1776));
    outputs(10109) <= not((layer4_outputs(208)) xor (layer4_outputs(5474)));
    outputs(10110) <= not((layer4_outputs(4961)) xor (layer4_outputs(3534)));
    outputs(10111) <= (layer4_outputs(1773)) xor (layer4_outputs(7337));
    outputs(10112) <= layer4_outputs(9554);
    outputs(10113) <= layer4_outputs(3305);
    outputs(10114) <= not(layer4_outputs(1242));
    outputs(10115) <= layer4_outputs(1057);
    outputs(10116) <= (layer4_outputs(9008)) xor (layer4_outputs(5538));
    outputs(10117) <= layer4_outputs(7808);
    outputs(10118) <= not(layer4_outputs(7016));
    outputs(10119) <= not(layer4_outputs(1194));
    outputs(10120) <= layer4_outputs(7783);
    outputs(10121) <= layer4_outputs(1850);
    outputs(10122) <= (layer4_outputs(6129)) xor (layer4_outputs(6442));
    outputs(10123) <= layer4_outputs(5129);
    outputs(10124) <= layer4_outputs(1872);
    outputs(10125) <= layer4_outputs(4989);
    outputs(10126) <= not(layer4_outputs(2254));
    outputs(10127) <= not(layer4_outputs(7074));
    outputs(10128) <= not(layer4_outputs(8164));
    outputs(10129) <= layer4_outputs(7509);
    outputs(10130) <= not((layer4_outputs(6192)) xor (layer4_outputs(1877)));
    outputs(10131) <= (layer4_outputs(9949)) xor (layer4_outputs(5157));
    outputs(10132) <= not(layer4_outputs(2323));
    outputs(10133) <= (layer4_outputs(2601)) and (layer4_outputs(519));
    outputs(10134) <= layer4_outputs(3922);
    outputs(10135) <= layer4_outputs(5853);
    outputs(10136) <= (layer4_outputs(4397)) xor (layer4_outputs(6583));
    outputs(10137) <= layer4_outputs(3774);
    outputs(10138) <= layer4_outputs(4094);
    outputs(10139) <= layer4_outputs(5960);
    outputs(10140) <= (layer4_outputs(8698)) xor (layer4_outputs(5543));
    outputs(10141) <= not(layer4_outputs(10224));
    outputs(10142) <= not(layer4_outputs(3242));
    outputs(10143) <= not((layer4_outputs(2462)) xor (layer4_outputs(988)));
    outputs(10144) <= (layer4_outputs(7733)) xor (layer4_outputs(6467));
    outputs(10145) <= layer4_outputs(8992);
    outputs(10146) <= not(layer4_outputs(49));
    outputs(10147) <= not(layer4_outputs(7417));
    outputs(10148) <= (layer4_outputs(2364)) xor (layer4_outputs(7464));
    outputs(10149) <= not(layer4_outputs(4312)) or (layer4_outputs(1115));
    outputs(10150) <= not((layer4_outputs(3297)) or (layer4_outputs(8314)));
    outputs(10151) <= not((layer4_outputs(7264)) and (layer4_outputs(7124)));
    outputs(10152) <= layer4_outputs(1705);
    outputs(10153) <= not(layer4_outputs(4341));
    outputs(10154) <= layer4_outputs(5287);
    outputs(10155) <= not((layer4_outputs(2689)) or (layer4_outputs(5147)));
    outputs(10156) <= not(layer4_outputs(4246));
    outputs(10157) <= '1';
    outputs(10158) <= not(layer4_outputs(5909));
    outputs(10159) <= layer4_outputs(6526);
    outputs(10160) <= (layer4_outputs(7677)) xor (layer4_outputs(747));
    outputs(10161) <= layer4_outputs(2329);
    outputs(10162) <= (layer4_outputs(999)) and not (layer4_outputs(3557));
    outputs(10163) <= (layer4_outputs(9966)) xor (layer4_outputs(4688));
    outputs(10164) <= not(layer4_outputs(1003));
    outputs(10165) <= layer4_outputs(2664);
    outputs(10166) <= layer4_outputs(8941);
    outputs(10167) <= layer4_outputs(5072);
    outputs(10168) <= (layer4_outputs(6800)) xor (layer4_outputs(5107));
    outputs(10169) <= not(layer4_outputs(2148));
    outputs(10170) <= not((layer4_outputs(3878)) xor (layer4_outputs(5474)));
    outputs(10171) <= layer4_outputs(334);
    outputs(10172) <= not(layer4_outputs(9916));
    outputs(10173) <= layer4_outputs(56);
    outputs(10174) <= not(layer4_outputs(1958));
    outputs(10175) <= (layer4_outputs(3852)) and (layer4_outputs(5232));
    outputs(10176) <= not(layer4_outputs(4270));
    outputs(10177) <= (layer4_outputs(2127)) and (layer4_outputs(2058));
    outputs(10178) <= layer4_outputs(9091);
    outputs(10179) <= layer4_outputs(1084);
    outputs(10180) <= not((layer4_outputs(543)) xor (layer4_outputs(8030)));
    outputs(10181) <= (layer4_outputs(4642)) xor (layer4_outputs(5578));
    outputs(10182) <= not((layer4_outputs(8004)) xor (layer4_outputs(2645)));
    outputs(10183) <= not((layer4_outputs(9980)) xor (layer4_outputs(8654)));
    outputs(10184) <= (layer4_outputs(2215)) and not (layer4_outputs(8350));
    outputs(10185) <= not(layer4_outputs(6042));
    outputs(10186) <= not(layer4_outputs(4469)) or (layer4_outputs(3019));
    outputs(10187) <= (layer4_outputs(9865)) xor (layer4_outputs(2447));
    outputs(10188) <= not(layer4_outputs(942)) or (layer4_outputs(654));
    outputs(10189) <= not(layer4_outputs(936));
    outputs(10190) <= not(layer4_outputs(1639));
    outputs(10191) <= layer4_outputs(3247);
    outputs(10192) <= layer4_outputs(5450);
    outputs(10193) <= layer4_outputs(6540);
    outputs(10194) <= layer4_outputs(324);
    outputs(10195) <= layer4_outputs(774);
    outputs(10196) <= (layer4_outputs(6872)) xor (layer4_outputs(8847));
    outputs(10197) <= not(layer4_outputs(2073));
    outputs(10198) <= layer4_outputs(1140);
    outputs(10199) <= not((layer4_outputs(5991)) or (layer4_outputs(2137)));
    outputs(10200) <= layer4_outputs(296);
    outputs(10201) <= not(layer4_outputs(7072));
    outputs(10202) <= not(layer4_outputs(1463));
    outputs(10203) <= layer4_outputs(3629);
    outputs(10204) <= (layer4_outputs(4727)) xor (layer4_outputs(467));
    outputs(10205) <= (layer4_outputs(3414)) and (layer4_outputs(2848));
    outputs(10206) <= layer4_outputs(1086);
    outputs(10207) <= not(layer4_outputs(369));
    outputs(10208) <= not(layer4_outputs(2163)) or (layer4_outputs(5795));
    outputs(10209) <= not(layer4_outputs(5322));
    outputs(10210) <= layer4_outputs(9384);
    outputs(10211) <= (layer4_outputs(7358)) and (layer4_outputs(2984));
    outputs(10212) <= (layer4_outputs(1528)) and not (layer4_outputs(665));
    outputs(10213) <= layer4_outputs(8016);
    outputs(10214) <= layer4_outputs(4205);
    outputs(10215) <= (layer4_outputs(1336)) xor (layer4_outputs(5101));
    outputs(10216) <= not(layer4_outputs(1307));
    outputs(10217) <= layer4_outputs(4470);
    outputs(10218) <= (layer4_outputs(4582)) xor (layer4_outputs(6504));
    outputs(10219) <= not(layer4_outputs(5836));
    outputs(10220) <= layer4_outputs(1150);
    outputs(10221) <= not((layer4_outputs(2853)) xor (layer4_outputs(9922)));
    outputs(10222) <= layer4_outputs(5704);
    outputs(10223) <= not((layer4_outputs(2239)) xor (layer4_outputs(10136)));
    outputs(10224) <= layer4_outputs(5744);
    outputs(10225) <= (layer4_outputs(7516)) xor (layer4_outputs(9154));
    outputs(10226) <= not(layer4_outputs(6423));
    outputs(10227) <= layer4_outputs(8127);
    outputs(10228) <= not((layer4_outputs(4981)) xor (layer4_outputs(4215)));
    outputs(10229) <= (layer4_outputs(6035)) and not (layer4_outputs(5180));
    outputs(10230) <= (layer4_outputs(183)) xor (layer4_outputs(7265));
    outputs(10231) <= (layer4_outputs(3953)) xor (layer4_outputs(7566));
    outputs(10232) <= not(layer4_outputs(8796));
    outputs(10233) <= (layer4_outputs(8436)) xor (layer4_outputs(8970));
    outputs(10234) <= not(layer4_outputs(2096));
    outputs(10235) <= not((layer4_outputs(9452)) or (layer4_outputs(5559)));
    outputs(10236) <= not((layer4_outputs(8684)) or (layer4_outputs(7827)));
    outputs(10237) <= not(layer4_outputs(9900));
    outputs(10238) <= (layer4_outputs(7550)) xor (layer4_outputs(9844));
    outputs(10239) <= not(layer4_outputs(3162));

end Behavioral;
