library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(2559 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);
    signal layer1_outputs : std_logic_vector(2559 downto 0);
    signal layer2_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not(inputs(241)) or (inputs(119));
    layer0_outputs(1) <= inputs(146);
    layer0_outputs(2) <= (inputs(51)) or (inputs(138));
    layer0_outputs(3) <= '1';
    layer0_outputs(4) <= not((inputs(186)) or (inputs(5)));
    layer0_outputs(5) <= inputs(138);
    layer0_outputs(6) <= not(inputs(66));
    layer0_outputs(7) <= not(inputs(240));
    layer0_outputs(8) <= '1';
    layer0_outputs(9) <= not(inputs(27));
    layer0_outputs(10) <= (inputs(173)) and (inputs(218));
    layer0_outputs(11) <= (inputs(61)) or (inputs(43));
    layer0_outputs(12) <= (inputs(49)) and (inputs(250));
    layer0_outputs(13) <= (inputs(20)) and not (inputs(7));
    layer0_outputs(14) <= not(inputs(78));
    layer0_outputs(15) <= not(inputs(57)) or (inputs(168));
    layer0_outputs(16) <= not(inputs(187));
    layer0_outputs(17) <= (inputs(84)) and not (inputs(160));
    layer0_outputs(18) <= (inputs(195)) and not (inputs(57));
    layer0_outputs(19) <= '1';
    layer0_outputs(20) <= (inputs(230)) or (inputs(175));
    layer0_outputs(21) <= not(inputs(50)) or (inputs(138));
    layer0_outputs(22) <= '0';
    layer0_outputs(23) <= not(inputs(23));
    layer0_outputs(24) <= not(inputs(195));
    layer0_outputs(25) <= '0';
    layer0_outputs(26) <= (inputs(48)) or (inputs(1));
    layer0_outputs(27) <= not((inputs(230)) or (inputs(247)));
    layer0_outputs(28) <= inputs(178);
    layer0_outputs(29) <= inputs(246);
    layer0_outputs(30) <= not(inputs(126));
    layer0_outputs(31) <= (inputs(23)) and not (inputs(216));
    layer0_outputs(32) <= not((inputs(168)) xor (inputs(170)));
    layer0_outputs(33) <= inputs(232);
    layer0_outputs(34) <= (inputs(181)) and (inputs(161));
    layer0_outputs(35) <= (inputs(101)) and not (inputs(65));
    layer0_outputs(36) <= inputs(12);
    layer0_outputs(37) <= '1';
    layer0_outputs(38) <= not((inputs(55)) and (inputs(155)));
    layer0_outputs(39) <= not(inputs(4));
    layer0_outputs(40) <= inputs(198);
    layer0_outputs(41) <= '1';
    layer0_outputs(42) <= (inputs(216)) or (inputs(3));
    layer0_outputs(43) <= not(inputs(173)) or (inputs(153));
    layer0_outputs(44) <= not((inputs(225)) or (inputs(119)));
    layer0_outputs(45) <= not(inputs(105));
    layer0_outputs(46) <= inputs(40);
    layer0_outputs(47) <= inputs(103);
    layer0_outputs(48) <= not(inputs(25)) or (inputs(182));
    layer0_outputs(49) <= not(inputs(255));
    layer0_outputs(50) <= (inputs(33)) and not (inputs(78));
    layer0_outputs(51) <= inputs(85);
    layer0_outputs(52) <= not(inputs(131));
    layer0_outputs(53) <= inputs(68);
    layer0_outputs(54) <= inputs(169);
    layer0_outputs(55) <= not(inputs(199)) or (inputs(9));
    layer0_outputs(56) <= not(inputs(180));
    layer0_outputs(57) <= not(inputs(250)) or (inputs(148));
    layer0_outputs(58) <= '0';
    layer0_outputs(59) <= (inputs(60)) and not (inputs(149));
    layer0_outputs(60) <= (inputs(164)) or (inputs(139));
    layer0_outputs(61) <= (inputs(6)) or (inputs(126));
    layer0_outputs(62) <= (inputs(44)) xor (inputs(12));
    layer0_outputs(63) <= not(inputs(90));
    layer0_outputs(64) <= (inputs(229)) or (inputs(208));
    layer0_outputs(65) <= (inputs(33)) and (inputs(54));
    layer0_outputs(66) <= '0';
    layer0_outputs(67) <= inputs(211);
    layer0_outputs(68) <= (inputs(86)) and not (inputs(17));
    layer0_outputs(69) <= not(inputs(60));
    layer0_outputs(70) <= not((inputs(159)) or (inputs(115)));
    layer0_outputs(71) <= not(inputs(54));
    layer0_outputs(72) <= not(inputs(247));
    layer0_outputs(73) <= (inputs(221)) or (inputs(175));
    layer0_outputs(74) <= inputs(100);
    layer0_outputs(75) <= (inputs(112)) or (inputs(187));
    layer0_outputs(76) <= not(inputs(197));
    layer0_outputs(77) <= '1';
    layer0_outputs(78) <= not((inputs(155)) xor (inputs(104)));
    layer0_outputs(79) <= not(inputs(99));
    layer0_outputs(80) <= inputs(213);
    layer0_outputs(81) <= '1';
    layer0_outputs(82) <= inputs(42);
    layer0_outputs(83) <= inputs(21);
    layer0_outputs(84) <= '0';
    layer0_outputs(85) <= not((inputs(197)) or (inputs(140)));
    layer0_outputs(86) <= not((inputs(234)) or (inputs(186)));
    layer0_outputs(87) <= not((inputs(18)) or (inputs(6)));
    layer0_outputs(88) <= (inputs(112)) or (inputs(4));
    layer0_outputs(89) <= (inputs(64)) or (inputs(51));
    layer0_outputs(90) <= '0';
    layer0_outputs(91) <= inputs(233);
    layer0_outputs(92) <= inputs(151);
    layer0_outputs(93) <= (inputs(52)) or (inputs(108));
    layer0_outputs(94) <= not(inputs(156));
    layer0_outputs(95) <= not(inputs(218));
    layer0_outputs(96) <= not((inputs(30)) or (inputs(98)));
    layer0_outputs(97) <= not((inputs(198)) or (inputs(33)));
    layer0_outputs(98) <= inputs(221);
    layer0_outputs(99) <= not(inputs(231));
    layer0_outputs(100) <= (inputs(78)) or (inputs(131));
    layer0_outputs(101) <= not((inputs(207)) or (inputs(224)));
    layer0_outputs(102) <= not(inputs(111)) or (inputs(114));
    layer0_outputs(103) <= (inputs(65)) xor (inputs(79));
    layer0_outputs(104) <= not(inputs(231)) or (inputs(15));
    layer0_outputs(105) <= not((inputs(223)) and (inputs(193)));
    layer0_outputs(106) <= not(inputs(35)) or (inputs(29));
    layer0_outputs(107) <= inputs(85);
    layer0_outputs(108) <= not((inputs(49)) or (inputs(27)));
    layer0_outputs(109) <= not((inputs(226)) or (inputs(224)));
    layer0_outputs(110) <= not(inputs(148));
    layer0_outputs(111) <= not(inputs(142));
    layer0_outputs(112) <= not(inputs(205)) or (inputs(110));
    layer0_outputs(113) <= (inputs(18)) or (inputs(16));
    layer0_outputs(114) <= (inputs(117)) xor (inputs(255));
    layer0_outputs(115) <= not(inputs(219)) or (inputs(14));
    layer0_outputs(116) <= '1';
    layer0_outputs(117) <= not(inputs(191)) or (inputs(174));
    layer0_outputs(118) <= not(inputs(227));
    layer0_outputs(119) <= not(inputs(43));
    layer0_outputs(120) <= not(inputs(115));
    layer0_outputs(121) <= (inputs(170)) or (inputs(160));
    layer0_outputs(122) <= not((inputs(247)) or (inputs(50)));
    layer0_outputs(123) <= (inputs(229)) and (inputs(251));
    layer0_outputs(124) <= (inputs(155)) and not (inputs(177));
    layer0_outputs(125) <= not((inputs(241)) or (inputs(156)));
    layer0_outputs(126) <= (inputs(139)) and not (inputs(47));
    layer0_outputs(127) <= inputs(22);
    layer0_outputs(128) <= (inputs(71)) and (inputs(45));
    layer0_outputs(129) <= inputs(71);
    layer0_outputs(130) <= inputs(119);
    layer0_outputs(131) <= '0';
    layer0_outputs(132) <= not((inputs(11)) or (inputs(171)));
    layer0_outputs(133) <= not(inputs(69)) or (inputs(32));
    layer0_outputs(134) <= (inputs(52)) and not (inputs(159));
    layer0_outputs(135) <= (inputs(6)) and (inputs(88));
    layer0_outputs(136) <= not(inputs(90));
    layer0_outputs(137) <= not((inputs(104)) or (inputs(63)));
    layer0_outputs(138) <= not((inputs(125)) or (inputs(22)));
    layer0_outputs(139) <= '0';
    layer0_outputs(140) <= inputs(82);
    layer0_outputs(141) <= (inputs(153)) and (inputs(219));
    layer0_outputs(142) <= (inputs(178)) or (inputs(201));
    layer0_outputs(143) <= '0';
    layer0_outputs(144) <= (inputs(216)) or (inputs(144));
    layer0_outputs(145) <= (inputs(163)) or (inputs(165));
    layer0_outputs(146) <= not(inputs(204)) or (inputs(154));
    layer0_outputs(147) <= inputs(221);
    layer0_outputs(148) <= (inputs(46)) or (inputs(212));
    layer0_outputs(149) <= '1';
    layer0_outputs(150) <= (inputs(210)) or (inputs(241));
    layer0_outputs(151) <= inputs(85);
    layer0_outputs(152) <= (inputs(122)) and not (inputs(228));
    layer0_outputs(153) <= (inputs(233)) and (inputs(231));
    layer0_outputs(154) <= (inputs(146)) or (inputs(116));
    layer0_outputs(155) <= not(inputs(122)) or (inputs(28));
    layer0_outputs(156) <= (inputs(228)) and (inputs(162));
    layer0_outputs(157) <= '0';
    layer0_outputs(158) <= (inputs(219)) or (inputs(250));
    layer0_outputs(159) <= not(inputs(243));
    layer0_outputs(160) <= (inputs(133)) and (inputs(67));
    layer0_outputs(161) <= inputs(93);
    layer0_outputs(162) <= not(inputs(65));
    layer0_outputs(163) <= not(inputs(177)) or (inputs(15));
    layer0_outputs(164) <= (inputs(61)) or (inputs(76));
    layer0_outputs(165) <= not((inputs(71)) xor (inputs(98)));
    layer0_outputs(166) <= not(inputs(3)) or (inputs(220));
    layer0_outputs(167) <= not(inputs(34));
    layer0_outputs(168) <= not((inputs(73)) or (inputs(226)));
    layer0_outputs(169) <= not(inputs(178));
    layer0_outputs(170) <= '0';
    layer0_outputs(171) <= (inputs(64)) or (inputs(182));
    layer0_outputs(172) <= inputs(162);
    layer0_outputs(173) <= not(inputs(251)) or (inputs(214));
    layer0_outputs(174) <= (inputs(118)) and not (inputs(229));
    layer0_outputs(175) <= not((inputs(227)) or (inputs(18)));
    layer0_outputs(176) <= inputs(133);
    layer0_outputs(177) <= not(inputs(117));
    layer0_outputs(178) <= inputs(72);
    layer0_outputs(179) <= (inputs(184)) and not (inputs(127));
    layer0_outputs(180) <= inputs(255);
    layer0_outputs(181) <= (inputs(150)) and not (inputs(15));
    layer0_outputs(182) <= not((inputs(202)) and (inputs(41)));
    layer0_outputs(183) <= (inputs(8)) or (inputs(70));
    layer0_outputs(184) <= not(inputs(172));
    layer0_outputs(185) <= not((inputs(242)) and (inputs(215)));
    layer0_outputs(186) <= not(inputs(41));
    layer0_outputs(187) <= not(inputs(133));
    layer0_outputs(188) <= inputs(244);
    layer0_outputs(189) <= not(inputs(137));
    layer0_outputs(190) <= not((inputs(17)) or (inputs(229)));
    layer0_outputs(191) <= not((inputs(207)) or (inputs(212)));
    layer0_outputs(192) <= inputs(75);
    layer0_outputs(193) <= inputs(226);
    layer0_outputs(194) <= (inputs(81)) or (inputs(63));
    layer0_outputs(195) <= '1';
    layer0_outputs(196) <= not(inputs(165)) or (inputs(92));
    layer0_outputs(197) <= inputs(80);
    layer0_outputs(198) <= inputs(17);
    layer0_outputs(199) <= not(inputs(57)) or (inputs(3));
    layer0_outputs(200) <= inputs(164);
    layer0_outputs(201) <= (inputs(20)) and not (inputs(72));
    layer0_outputs(202) <= not((inputs(52)) or (inputs(218)));
    layer0_outputs(203) <= not(inputs(138));
    layer0_outputs(204) <= '0';
    layer0_outputs(205) <= not(inputs(230));
    layer0_outputs(206) <= (inputs(171)) or (inputs(218));
    layer0_outputs(207) <= inputs(126);
    layer0_outputs(208) <= (inputs(29)) and not (inputs(121));
    layer0_outputs(209) <= inputs(93);
    layer0_outputs(210) <= (inputs(44)) or (inputs(239));
    layer0_outputs(211) <= '1';
    layer0_outputs(212) <= (inputs(110)) and not (inputs(66));
    layer0_outputs(213) <= inputs(181);
    layer0_outputs(214) <= not(inputs(160));
    layer0_outputs(215) <= (inputs(38)) and not (inputs(175));
    layer0_outputs(216) <= not(inputs(46));
    layer0_outputs(217) <= not((inputs(89)) or (inputs(122)));
    layer0_outputs(218) <= not((inputs(163)) or (inputs(23)));
    layer0_outputs(219) <= not((inputs(109)) xor (inputs(178)));
    layer0_outputs(220) <= not(inputs(136));
    layer0_outputs(221) <= '1';
    layer0_outputs(222) <= (inputs(199)) and not (inputs(19));
    layer0_outputs(223) <= (inputs(108)) and (inputs(232));
    layer0_outputs(224) <= (inputs(134)) and (inputs(242));
    layer0_outputs(225) <= not(inputs(48));
    layer0_outputs(226) <= (inputs(49)) and not (inputs(113));
    layer0_outputs(227) <= '0';
    layer0_outputs(228) <= (inputs(39)) or (inputs(24));
    layer0_outputs(229) <= not(inputs(116));
    layer0_outputs(230) <= (inputs(239)) or (inputs(114));
    layer0_outputs(231) <= not(inputs(8));
    layer0_outputs(232) <= (inputs(24)) and (inputs(26));
    layer0_outputs(233) <= not(inputs(121)) or (inputs(210));
    layer0_outputs(234) <= not(inputs(217)) or (inputs(124));
    layer0_outputs(235) <= '0';
    layer0_outputs(236) <= inputs(165);
    layer0_outputs(237) <= not(inputs(180));
    layer0_outputs(238) <= (inputs(78)) or (inputs(92));
    layer0_outputs(239) <= not(inputs(194));
    layer0_outputs(240) <= (inputs(120)) xor (inputs(188));
    layer0_outputs(241) <= not(inputs(114));
    layer0_outputs(242) <= (inputs(179)) or (inputs(142));
    layer0_outputs(243) <= not(inputs(50));
    layer0_outputs(244) <= (inputs(131)) or (inputs(162));
    layer0_outputs(245) <= not(inputs(46)) or (inputs(146));
    layer0_outputs(246) <= inputs(24);
    layer0_outputs(247) <= (inputs(198)) and not (inputs(191));
    layer0_outputs(248) <= not(inputs(211));
    layer0_outputs(249) <= not(inputs(35));
    layer0_outputs(250) <= '0';
    layer0_outputs(251) <= not((inputs(134)) or (inputs(31)));
    layer0_outputs(252) <= '0';
    layer0_outputs(253) <= (inputs(179)) and not (inputs(172));
    layer0_outputs(254) <= not(inputs(186));
    layer0_outputs(255) <= inputs(182);
    layer0_outputs(256) <= not(inputs(182));
    layer0_outputs(257) <= '1';
    layer0_outputs(258) <= not(inputs(168));
    layer0_outputs(259) <= not(inputs(2)) or (inputs(123));
    layer0_outputs(260) <= not((inputs(157)) or (inputs(61)));
    layer0_outputs(261) <= inputs(166);
    layer0_outputs(262) <= inputs(181);
    layer0_outputs(263) <= '0';
    layer0_outputs(264) <= not(inputs(26)) or (inputs(154));
    layer0_outputs(265) <= not(inputs(132));
    layer0_outputs(266) <= not((inputs(7)) or (inputs(33)));
    layer0_outputs(267) <= (inputs(126)) and not (inputs(15));
    layer0_outputs(268) <= not((inputs(171)) or (inputs(149)));
    layer0_outputs(269) <= not((inputs(209)) or (inputs(104)));
    layer0_outputs(270) <= not(inputs(130));
    layer0_outputs(271) <= (inputs(40)) or (inputs(6));
    layer0_outputs(272) <= (inputs(75)) or (inputs(60));
    layer0_outputs(273) <= (inputs(229)) and not (inputs(223));
    layer0_outputs(274) <= not((inputs(69)) or (inputs(98)));
    layer0_outputs(275) <= not(inputs(230));
    layer0_outputs(276) <= not((inputs(144)) xor (inputs(179)));
    layer0_outputs(277) <= (inputs(210)) or (inputs(212));
    layer0_outputs(278) <= not(inputs(209));
    layer0_outputs(279) <= (inputs(180)) and not (inputs(73));
    layer0_outputs(280) <= inputs(154);
    layer0_outputs(281) <= not((inputs(255)) or (inputs(57)));
    layer0_outputs(282) <= (inputs(163)) or (inputs(149));
    layer0_outputs(283) <= inputs(229);
    layer0_outputs(284) <= not(inputs(84));
    layer0_outputs(285) <= (inputs(237)) and (inputs(242));
    layer0_outputs(286) <= not(inputs(236)) or (inputs(132));
    layer0_outputs(287) <= not(inputs(71));
    layer0_outputs(288) <= (inputs(136)) and not (inputs(128));
    layer0_outputs(289) <= '0';
    layer0_outputs(290) <= (inputs(225)) or (inputs(207));
    layer0_outputs(291) <= (inputs(184)) and (inputs(133));
    layer0_outputs(292) <= not(inputs(25)) or (inputs(127));
    layer0_outputs(293) <= '0';
    layer0_outputs(294) <= (inputs(88)) or (inputs(25));
    layer0_outputs(295) <= not(inputs(236)) or (inputs(113));
    layer0_outputs(296) <= not((inputs(118)) or (inputs(85)));
    layer0_outputs(297) <= not(inputs(10));
    layer0_outputs(298) <= (inputs(180)) and not (inputs(227));
    layer0_outputs(299) <= inputs(118);
    layer0_outputs(300) <= not(inputs(109)) or (inputs(246));
    layer0_outputs(301) <= not(inputs(53)) or (inputs(225));
    layer0_outputs(302) <= inputs(29);
    layer0_outputs(303) <= not((inputs(254)) or (inputs(94)));
    layer0_outputs(304) <= inputs(78);
    layer0_outputs(305) <= not(inputs(158)) or (inputs(181));
    layer0_outputs(306) <= inputs(198);
    layer0_outputs(307) <= '1';
    layer0_outputs(308) <= '0';
    layer0_outputs(309) <= not((inputs(182)) xor (inputs(12)));
    layer0_outputs(310) <= not((inputs(13)) and (inputs(66)));
    layer0_outputs(311) <= not(inputs(204)) or (inputs(128));
    layer0_outputs(312) <= not((inputs(224)) xor (inputs(188)));
    layer0_outputs(313) <= '0';
    layer0_outputs(314) <= inputs(14);
    layer0_outputs(315) <= not(inputs(97));
    layer0_outputs(316) <= not(inputs(119));
    layer0_outputs(317) <= not(inputs(118)) or (inputs(124));
    layer0_outputs(318) <= (inputs(52)) and not (inputs(33));
    layer0_outputs(319) <= (inputs(25)) or (inputs(63));
    layer0_outputs(320) <= not(inputs(112)) or (inputs(31));
    layer0_outputs(321) <= not(inputs(229)) or (inputs(255));
    layer0_outputs(322) <= inputs(158);
    layer0_outputs(323) <= '1';
    layer0_outputs(324) <= not(inputs(53));
    layer0_outputs(325) <= not((inputs(35)) or (inputs(108)));
    layer0_outputs(326) <= not(inputs(92));
    layer0_outputs(327) <= inputs(82);
    layer0_outputs(328) <= not(inputs(79));
    layer0_outputs(329) <= not(inputs(35));
    layer0_outputs(330) <= not(inputs(200)) or (inputs(81));
    layer0_outputs(331) <= not((inputs(129)) or (inputs(253)));
    layer0_outputs(332) <= (inputs(39)) and (inputs(103));
    layer0_outputs(333) <= not(inputs(125));
    layer0_outputs(334) <= not(inputs(130));
    layer0_outputs(335) <= (inputs(254)) and not (inputs(224));
    layer0_outputs(336) <= not((inputs(181)) xor (inputs(62)));
    layer0_outputs(337) <= inputs(116);
    layer0_outputs(338) <= '0';
    layer0_outputs(339) <= (inputs(2)) or (inputs(222));
    layer0_outputs(340) <= not(inputs(20));
    layer0_outputs(341) <= inputs(69);
    layer0_outputs(342) <= inputs(29);
    layer0_outputs(343) <= (inputs(211)) or (inputs(22));
    layer0_outputs(344) <= not(inputs(135));
    layer0_outputs(345) <= not(inputs(31));
    layer0_outputs(346) <= (inputs(12)) or (inputs(54));
    layer0_outputs(347) <= not(inputs(89));
    layer0_outputs(348) <= (inputs(238)) and not (inputs(71));
    layer0_outputs(349) <= inputs(90);
    layer0_outputs(350) <= not(inputs(117));
    layer0_outputs(351) <= inputs(196);
    layer0_outputs(352) <= inputs(99);
    layer0_outputs(353) <= (inputs(87)) and (inputs(31));
    layer0_outputs(354) <= not((inputs(128)) or (inputs(55)));
    layer0_outputs(355) <= inputs(76);
    layer0_outputs(356) <= not(inputs(121)) or (inputs(218));
    layer0_outputs(357) <= not(inputs(90));
    layer0_outputs(358) <= inputs(231);
    layer0_outputs(359) <= not((inputs(1)) and (inputs(192)));
    layer0_outputs(360) <= not(inputs(224));
    layer0_outputs(361) <= '0';
    layer0_outputs(362) <= not((inputs(254)) xor (inputs(104)));
    layer0_outputs(363) <= inputs(17);
    layer0_outputs(364) <= not(inputs(79));
    layer0_outputs(365) <= not((inputs(191)) or (inputs(35)));
    layer0_outputs(366) <= not((inputs(218)) xor (inputs(170)));
    layer0_outputs(367) <= inputs(153);
    layer0_outputs(368) <= inputs(113);
    layer0_outputs(369) <= not((inputs(244)) or (inputs(250)));
    layer0_outputs(370) <= not((inputs(47)) and (inputs(0)));
    layer0_outputs(371) <= not(inputs(127)) or (inputs(255));
    layer0_outputs(372) <= not(inputs(115));
    layer0_outputs(373) <= not(inputs(131));
    layer0_outputs(374) <= not(inputs(84));
    layer0_outputs(375) <= not(inputs(228));
    layer0_outputs(376) <= not(inputs(231)) or (inputs(48));
    layer0_outputs(377) <= inputs(130);
    layer0_outputs(378) <= not(inputs(185));
    layer0_outputs(379) <= not(inputs(150)) or (inputs(63));
    layer0_outputs(380) <= inputs(49);
    layer0_outputs(381) <= not(inputs(201)) or (inputs(215));
    layer0_outputs(382) <= inputs(170);
    layer0_outputs(383) <= (inputs(61)) and (inputs(183));
    layer0_outputs(384) <= inputs(97);
    layer0_outputs(385) <= '0';
    layer0_outputs(386) <= not((inputs(195)) or (inputs(53)));
    layer0_outputs(387) <= inputs(81);
    layer0_outputs(388) <= not((inputs(183)) and (inputs(234)));
    layer0_outputs(389) <= not(inputs(25)) or (inputs(40));
    layer0_outputs(390) <= (inputs(114)) or (inputs(115));
    layer0_outputs(391) <= not(inputs(94));
    layer0_outputs(392) <= (inputs(69)) or (inputs(204));
    layer0_outputs(393) <= not(inputs(55));
    layer0_outputs(394) <= inputs(180);
    layer0_outputs(395) <= inputs(62);
    layer0_outputs(396) <= (inputs(46)) or (inputs(37));
    layer0_outputs(397) <= not(inputs(88));
    layer0_outputs(398) <= not((inputs(149)) or (inputs(235)));
    layer0_outputs(399) <= inputs(217);
    layer0_outputs(400) <= not(inputs(199));
    layer0_outputs(401) <= (inputs(217)) xor (inputs(38));
    layer0_outputs(402) <= not((inputs(238)) or (inputs(53)));
    layer0_outputs(403) <= not(inputs(186)) or (inputs(27));
    layer0_outputs(404) <= '0';
    layer0_outputs(405) <= '0';
    layer0_outputs(406) <= inputs(183);
    layer0_outputs(407) <= (inputs(12)) and not (inputs(209));
    layer0_outputs(408) <= (inputs(31)) and not (inputs(181));
    layer0_outputs(409) <= not(inputs(104)) or (inputs(97));
    layer0_outputs(410) <= not((inputs(213)) or (inputs(141)));
    layer0_outputs(411) <= (inputs(108)) or (inputs(32));
    layer0_outputs(412) <= not((inputs(101)) or (inputs(145)));
    layer0_outputs(413) <= not((inputs(68)) or (inputs(108)));
    layer0_outputs(414) <= inputs(176);
    layer0_outputs(415) <= '0';
    layer0_outputs(416) <= (inputs(67)) or (inputs(122));
    layer0_outputs(417) <= inputs(146);
    layer0_outputs(418) <= inputs(239);
    layer0_outputs(419) <= '1';
    layer0_outputs(420) <= (inputs(97)) or (inputs(238));
    layer0_outputs(421) <= inputs(202);
    layer0_outputs(422) <= inputs(162);
    layer0_outputs(423) <= not(inputs(114)) or (inputs(156));
    layer0_outputs(424) <= inputs(93);
    layer0_outputs(425) <= not(inputs(198));
    layer0_outputs(426) <= (inputs(65)) or (inputs(153));
    layer0_outputs(427) <= not((inputs(181)) or (inputs(83)));
    layer0_outputs(428) <= not(inputs(14)) or (inputs(106));
    layer0_outputs(429) <= not(inputs(103));
    layer0_outputs(430) <= not((inputs(133)) xor (inputs(228)));
    layer0_outputs(431) <= not(inputs(162));
    layer0_outputs(432) <= (inputs(91)) and not (inputs(157));
    layer0_outputs(433) <= not(inputs(75));
    layer0_outputs(434) <= not((inputs(218)) or (inputs(158)));
    layer0_outputs(435) <= not((inputs(187)) xor (inputs(34)));
    layer0_outputs(436) <= (inputs(19)) or (inputs(122));
    layer0_outputs(437) <= (inputs(76)) and (inputs(9));
    layer0_outputs(438) <= not(inputs(122));
    layer0_outputs(439) <= (inputs(183)) and (inputs(42));
    layer0_outputs(440) <= not(inputs(194));
    layer0_outputs(441) <= (inputs(148)) and not (inputs(224));
    layer0_outputs(442) <= not(inputs(146));
    layer0_outputs(443) <= '0';
    layer0_outputs(444) <= not(inputs(182));
    layer0_outputs(445) <= not(inputs(255));
    layer0_outputs(446) <= not((inputs(83)) or (inputs(234)));
    layer0_outputs(447) <= not((inputs(173)) or (inputs(20)));
    layer0_outputs(448) <= not(inputs(119)) or (inputs(206));
    layer0_outputs(449) <= (inputs(170)) or (inputs(102));
    layer0_outputs(450) <= not((inputs(240)) and (inputs(170)));
    layer0_outputs(451) <= not(inputs(103)) or (inputs(163));
    layer0_outputs(452) <= not(inputs(7)) or (inputs(100));
    layer0_outputs(453) <= (inputs(146)) or (inputs(101));
    layer0_outputs(454) <= (inputs(88)) and not (inputs(108));
    layer0_outputs(455) <= inputs(118);
    layer0_outputs(456) <= not((inputs(54)) or (inputs(193)));
    layer0_outputs(457) <= not(inputs(204));
    layer0_outputs(458) <= not(inputs(34)) or (inputs(34));
    layer0_outputs(459) <= not(inputs(43));
    layer0_outputs(460) <= not((inputs(2)) or (inputs(7)));
    layer0_outputs(461) <= not(inputs(51)) or (inputs(54));
    layer0_outputs(462) <= (inputs(224)) or (inputs(81));
    layer0_outputs(463) <= not(inputs(99));
    layer0_outputs(464) <= not(inputs(155)) or (inputs(121));
    layer0_outputs(465) <= (inputs(21)) and not (inputs(66));
    layer0_outputs(466) <= inputs(227);
    layer0_outputs(467) <= '1';
    layer0_outputs(468) <= not(inputs(143));
    layer0_outputs(469) <= not((inputs(140)) or (inputs(84)));
    layer0_outputs(470) <= not(inputs(120)) or (inputs(146));
    layer0_outputs(471) <= (inputs(228)) and not (inputs(217));
    layer0_outputs(472) <= (inputs(244)) and (inputs(126));
    layer0_outputs(473) <= (inputs(208)) or (inputs(186));
    layer0_outputs(474) <= (inputs(71)) and not (inputs(66));
    layer0_outputs(475) <= not(inputs(175));
    layer0_outputs(476) <= inputs(37);
    layer0_outputs(477) <= not(inputs(178));
    layer0_outputs(478) <= not(inputs(114));
    layer0_outputs(479) <= not(inputs(223)) or (inputs(77));
    layer0_outputs(480) <= inputs(25);
    layer0_outputs(481) <= not(inputs(103));
    layer0_outputs(482) <= not(inputs(211));
    layer0_outputs(483) <= not(inputs(95));
    layer0_outputs(484) <= not(inputs(165)) or (inputs(89));
    layer0_outputs(485) <= not((inputs(53)) or (inputs(80)));
    layer0_outputs(486) <= not(inputs(153));
    layer0_outputs(487) <= not(inputs(106)) or (inputs(196));
    layer0_outputs(488) <= '0';
    layer0_outputs(489) <= (inputs(155)) and not (inputs(137));
    layer0_outputs(490) <= not(inputs(44));
    layer0_outputs(491) <= (inputs(199)) and not (inputs(134));
    layer0_outputs(492) <= '1';
    layer0_outputs(493) <= not((inputs(225)) or (inputs(31)));
    layer0_outputs(494) <= not(inputs(130));
    layer0_outputs(495) <= '0';
    layer0_outputs(496) <= not((inputs(111)) or (inputs(194)));
    layer0_outputs(497) <= not(inputs(121));
    layer0_outputs(498) <= not(inputs(232)) or (inputs(2));
    layer0_outputs(499) <= not(inputs(42));
    layer0_outputs(500) <= not(inputs(151));
    layer0_outputs(501) <= not(inputs(21)) or (inputs(85));
    layer0_outputs(502) <= not(inputs(68));
    layer0_outputs(503) <= not(inputs(157));
    layer0_outputs(504) <= inputs(77);
    layer0_outputs(505) <= inputs(195);
    layer0_outputs(506) <= not(inputs(125)) or (inputs(181));
    layer0_outputs(507) <= (inputs(18)) or (inputs(227));
    layer0_outputs(508) <= inputs(29);
    layer0_outputs(509) <= inputs(123);
    layer0_outputs(510) <= '1';
    layer0_outputs(511) <= (inputs(144)) or (inputs(130));
    layer0_outputs(512) <= not((inputs(234)) and (inputs(199)));
    layer0_outputs(513) <= (inputs(79)) or (inputs(202));
    layer0_outputs(514) <= inputs(112);
    layer0_outputs(515) <= '1';
    layer0_outputs(516) <= '0';
    layer0_outputs(517) <= inputs(15);
    layer0_outputs(518) <= (inputs(109)) and not (inputs(109));
    layer0_outputs(519) <= not((inputs(38)) xor (inputs(87)));
    layer0_outputs(520) <= not(inputs(83));
    layer0_outputs(521) <= not((inputs(190)) and (inputs(70)));
    layer0_outputs(522) <= (inputs(252)) or (inputs(98));
    layer0_outputs(523) <= not((inputs(34)) or (inputs(32)));
    layer0_outputs(524) <= not(inputs(94));
    layer0_outputs(525) <= not(inputs(121));
    layer0_outputs(526) <= (inputs(36)) or (inputs(60));
    layer0_outputs(527) <= '1';
    layer0_outputs(528) <= (inputs(215)) and not (inputs(39));
    layer0_outputs(529) <= (inputs(231)) and not (inputs(238));
    layer0_outputs(530) <= inputs(105);
    layer0_outputs(531) <= not(inputs(84));
    layer0_outputs(532) <= (inputs(6)) and not (inputs(221));
    layer0_outputs(533) <= inputs(228);
    layer0_outputs(534) <= inputs(26);
    layer0_outputs(535) <= inputs(59);
    layer0_outputs(536) <= not(inputs(26));
    layer0_outputs(537) <= (inputs(117)) and not (inputs(93));
    layer0_outputs(538) <= not((inputs(62)) xor (inputs(113)));
    layer0_outputs(539) <= inputs(131);
    layer0_outputs(540) <= (inputs(24)) and (inputs(149));
    layer0_outputs(541) <= inputs(56);
    layer0_outputs(542) <= (inputs(225)) or (inputs(195));
    layer0_outputs(543) <= (inputs(255)) and (inputs(70));
    layer0_outputs(544) <= (inputs(107)) xor (inputs(175));
    layer0_outputs(545) <= (inputs(120)) xor (inputs(133));
    layer0_outputs(546) <= (inputs(109)) and not (inputs(30));
    layer0_outputs(547) <= not((inputs(134)) or (inputs(3)));
    layer0_outputs(548) <= not((inputs(247)) and (inputs(88)));
    layer0_outputs(549) <= inputs(41);
    layer0_outputs(550) <= not(inputs(21)) or (inputs(99));
    layer0_outputs(551) <= not(inputs(23));
    layer0_outputs(552) <= not(inputs(146));
    layer0_outputs(553) <= (inputs(187)) xor (inputs(219));
    layer0_outputs(554) <= not(inputs(60));
    layer0_outputs(555) <= inputs(21);
    layer0_outputs(556) <= (inputs(189)) or (inputs(87));
    layer0_outputs(557) <= not(inputs(8));
    layer0_outputs(558) <= inputs(129);
    layer0_outputs(559) <= (inputs(103)) and not (inputs(8));
    layer0_outputs(560) <= inputs(177);
    layer0_outputs(561) <= (inputs(119)) or (inputs(88));
    layer0_outputs(562) <= not((inputs(175)) or (inputs(188)));
    layer0_outputs(563) <= (inputs(248)) and not (inputs(82));
    layer0_outputs(564) <= inputs(100);
    layer0_outputs(565) <= (inputs(46)) or (inputs(106));
    layer0_outputs(566) <= (inputs(211)) and (inputs(239));
    layer0_outputs(567) <= inputs(195);
    layer0_outputs(568) <= inputs(182);
    layer0_outputs(569) <= not((inputs(139)) or (inputs(204)));
    layer0_outputs(570) <= not(inputs(149)) or (inputs(36));
    layer0_outputs(571) <= not(inputs(81));
    layer0_outputs(572) <= inputs(224);
    layer0_outputs(573) <= not(inputs(226));
    layer0_outputs(574) <= inputs(22);
    layer0_outputs(575) <= '1';
    layer0_outputs(576) <= inputs(138);
    layer0_outputs(577) <= '1';
    layer0_outputs(578) <= '0';
    layer0_outputs(579) <= not(inputs(120));
    layer0_outputs(580) <= not(inputs(53));
    layer0_outputs(581) <= not(inputs(173)) or (inputs(14));
    layer0_outputs(582) <= '1';
    layer0_outputs(583) <= (inputs(241)) xor (inputs(11));
    layer0_outputs(584) <= not(inputs(104)) or (inputs(189));
    layer0_outputs(585) <= inputs(184);
    layer0_outputs(586) <= (inputs(211)) and not (inputs(103));
    layer0_outputs(587) <= not((inputs(172)) or (inputs(80)));
    layer0_outputs(588) <= not(inputs(220)) or (inputs(12));
    layer0_outputs(589) <= not(inputs(248)) or (inputs(29));
    layer0_outputs(590) <= not(inputs(223));
    layer0_outputs(591) <= inputs(17);
    layer0_outputs(592) <= not(inputs(221));
    layer0_outputs(593) <= not((inputs(98)) or (inputs(176)));
    layer0_outputs(594) <= not(inputs(174));
    layer0_outputs(595) <= not((inputs(148)) or (inputs(150)));
    layer0_outputs(596) <= (inputs(111)) xor (inputs(171));
    layer0_outputs(597) <= not(inputs(198));
    layer0_outputs(598) <= inputs(72);
    layer0_outputs(599) <= not((inputs(5)) or (inputs(253)));
    layer0_outputs(600) <= (inputs(126)) and not (inputs(153));
    layer0_outputs(601) <= inputs(123);
    layer0_outputs(602) <= (inputs(17)) and not (inputs(236));
    layer0_outputs(603) <= inputs(184);
    layer0_outputs(604) <= (inputs(15)) and not (inputs(47));
    layer0_outputs(605) <= not((inputs(36)) or (inputs(47)));
    layer0_outputs(606) <= (inputs(215)) and not (inputs(45));
    layer0_outputs(607) <= not((inputs(18)) xor (inputs(191)));
    layer0_outputs(608) <= (inputs(39)) or (inputs(107));
    layer0_outputs(609) <= not(inputs(128)) or (inputs(150));
    layer0_outputs(610) <= (inputs(148)) and not (inputs(95));
    layer0_outputs(611) <= not(inputs(84));
    layer0_outputs(612) <= not((inputs(39)) or (inputs(38)));
    layer0_outputs(613) <= not(inputs(122));
    layer0_outputs(614) <= not(inputs(142)) or (inputs(167));
    layer0_outputs(615) <= (inputs(117)) or (inputs(192));
    layer0_outputs(616) <= inputs(17);
    layer0_outputs(617) <= not(inputs(40));
    layer0_outputs(618) <= (inputs(39)) or (inputs(192));
    layer0_outputs(619) <= not((inputs(17)) or (inputs(111)));
    layer0_outputs(620) <= inputs(53);
    layer0_outputs(621) <= not((inputs(78)) and (inputs(232)));
    layer0_outputs(622) <= not(inputs(86));
    layer0_outputs(623) <= (inputs(28)) and not (inputs(248));
    layer0_outputs(624) <= not((inputs(170)) or (inputs(114)));
    layer0_outputs(625) <= (inputs(132)) and not (inputs(234));
    layer0_outputs(626) <= not((inputs(192)) xor (inputs(18)));
    layer0_outputs(627) <= not((inputs(144)) and (inputs(97)));
    layer0_outputs(628) <= inputs(237);
    layer0_outputs(629) <= not(inputs(232)) or (inputs(25));
    layer0_outputs(630) <= inputs(215);
    layer0_outputs(631) <= '0';
    layer0_outputs(632) <= inputs(167);
    layer0_outputs(633) <= (inputs(121)) and not (inputs(56));
    layer0_outputs(634) <= not(inputs(103)) or (inputs(111));
    layer0_outputs(635) <= inputs(169);
    layer0_outputs(636) <= not((inputs(203)) and (inputs(119)));
    layer0_outputs(637) <= not((inputs(206)) or (inputs(19)));
    layer0_outputs(638) <= not((inputs(172)) xor (inputs(205)));
    layer0_outputs(639) <= (inputs(147)) and not (inputs(166));
    layer0_outputs(640) <= '0';
    layer0_outputs(641) <= (inputs(12)) xor (inputs(56));
    layer0_outputs(642) <= not(inputs(168));
    layer0_outputs(643) <= not(inputs(38));
    layer0_outputs(644) <= (inputs(37)) and (inputs(210));
    layer0_outputs(645) <= not(inputs(149));
    layer0_outputs(646) <= (inputs(110)) or (inputs(157));
    layer0_outputs(647) <= inputs(42);
    layer0_outputs(648) <= (inputs(197)) and not (inputs(141));
    layer0_outputs(649) <= inputs(237);
    layer0_outputs(650) <= inputs(122);
    layer0_outputs(651) <= not((inputs(45)) and (inputs(17)));
    layer0_outputs(652) <= inputs(100);
    layer0_outputs(653) <= not(inputs(92)) or (inputs(210));
    layer0_outputs(654) <= (inputs(251)) xor (inputs(171));
    layer0_outputs(655) <= inputs(249);
    layer0_outputs(656) <= inputs(194);
    layer0_outputs(657) <= not((inputs(146)) or (inputs(170)));
    layer0_outputs(658) <= inputs(11);
    layer0_outputs(659) <= inputs(118);
    layer0_outputs(660) <= not(inputs(26)) or (inputs(208));
    layer0_outputs(661) <= not(inputs(49)) or (inputs(237));
    layer0_outputs(662) <= not(inputs(25)) or (inputs(132));
    layer0_outputs(663) <= (inputs(249)) and not (inputs(175));
    layer0_outputs(664) <= not(inputs(93));
    layer0_outputs(665) <= (inputs(160)) or (inputs(13));
    layer0_outputs(666) <= (inputs(134)) and not (inputs(16));
    layer0_outputs(667) <= (inputs(225)) and not (inputs(106));
    layer0_outputs(668) <= not((inputs(235)) or (inputs(79)));
    layer0_outputs(669) <= (inputs(219)) or (inputs(153));
    layer0_outputs(670) <= not((inputs(196)) and (inputs(187)));
    layer0_outputs(671) <= '1';
    layer0_outputs(672) <= not(inputs(237));
    layer0_outputs(673) <= '1';
    layer0_outputs(674) <= (inputs(7)) xor (inputs(42));
    layer0_outputs(675) <= '0';
    layer0_outputs(676) <= not((inputs(139)) and (inputs(135)));
    layer0_outputs(677) <= (inputs(104)) and not (inputs(126));
    layer0_outputs(678) <= (inputs(85)) or (inputs(145));
    layer0_outputs(679) <= '0';
    layer0_outputs(680) <= not(inputs(232)) or (inputs(110));
    layer0_outputs(681) <= (inputs(64)) or (inputs(60));
    layer0_outputs(682) <= '1';
    layer0_outputs(683) <= not(inputs(99));
    layer0_outputs(684) <= (inputs(206)) and not (inputs(7));
    layer0_outputs(685) <= inputs(39);
    layer0_outputs(686) <= not(inputs(102));
    layer0_outputs(687) <= not(inputs(4)) or (inputs(116));
    layer0_outputs(688) <= not(inputs(208)) or (inputs(0));
    layer0_outputs(689) <= inputs(208);
    layer0_outputs(690) <= not((inputs(146)) or (inputs(61)));
    layer0_outputs(691) <= not(inputs(78)) or (inputs(255));
    layer0_outputs(692) <= (inputs(99)) and (inputs(108));
    layer0_outputs(693) <= not(inputs(112));
    layer0_outputs(694) <= inputs(136);
    layer0_outputs(695) <= not((inputs(161)) or (inputs(144)));
    layer0_outputs(696) <= not((inputs(220)) or (inputs(238)));
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= (inputs(212)) and not (inputs(133));
    layer0_outputs(699) <= not(inputs(162));
    layer0_outputs(700) <= (inputs(211)) or (inputs(254));
    layer0_outputs(701) <= (inputs(95)) or (inputs(99));
    layer0_outputs(702) <= not((inputs(156)) or (inputs(9)));
    layer0_outputs(703) <= (inputs(185)) xor (inputs(217));
    layer0_outputs(704) <= not(inputs(110));
    layer0_outputs(705) <= not((inputs(185)) or (inputs(40)));
    layer0_outputs(706) <= (inputs(120)) and (inputs(140));
    layer0_outputs(707) <= (inputs(230)) or (inputs(101));
    layer0_outputs(708) <= '0';
    layer0_outputs(709) <= not((inputs(44)) or (inputs(247)));
    layer0_outputs(710) <= (inputs(191)) or (inputs(230));
    layer0_outputs(711) <= not(inputs(114));
    layer0_outputs(712) <= '0';
    layer0_outputs(713) <= (inputs(56)) and not (inputs(113));
    layer0_outputs(714) <= not(inputs(78)) or (inputs(171));
    layer0_outputs(715) <= (inputs(106)) and not (inputs(56));
    layer0_outputs(716) <= (inputs(85)) and not (inputs(175));
    layer0_outputs(717) <= not(inputs(188)) or (inputs(137));
    layer0_outputs(718) <= not(inputs(107)) or (inputs(190));
    layer0_outputs(719) <= (inputs(148)) or (inputs(89));
    layer0_outputs(720) <= (inputs(99)) and not (inputs(42));
    layer0_outputs(721) <= (inputs(116)) and not (inputs(125));
    layer0_outputs(722) <= not((inputs(191)) or (inputs(20)));
    layer0_outputs(723) <= '0';
    layer0_outputs(724) <= not((inputs(148)) or (inputs(110)));
    layer0_outputs(725) <= '1';
    layer0_outputs(726) <= not(inputs(28));
    layer0_outputs(727) <= inputs(120);
    layer0_outputs(728) <= not((inputs(159)) or (inputs(250)));
    layer0_outputs(729) <= (inputs(50)) and not (inputs(218));
    layer0_outputs(730) <= inputs(239);
    layer0_outputs(731) <= '0';
    layer0_outputs(732) <= inputs(100);
    layer0_outputs(733) <= inputs(196);
    layer0_outputs(734) <= '1';
    layer0_outputs(735) <= inputs(23);
    layer0_outputs(736) <= (inputs(11)) or (inputs(35));
    layer0_outputs(737) <= (inputs(235)) and not (inputs(49));
    layer0_outputs(738) <= (inputs(26)) and (inputs(29));
    layer0_outputs(739) <= inputs(228);
    layer0_outputs(740) <= (inputs(121)) or (inputs(151));
    layer0_outputs(741) <= not(inputs(71)) or (inputs(59));
    layer0_outputs(742) <= not(inputs(54));
    layer0_outputs(743) <= not((inputs(172)) xor (inputs(251)));
    layer0_outputs(744) <= not(inputs(110));
    layer0_outputs(745) <= not(inputs(166)) or (inputs(93));
    layer0_outputs(746) <= inputs(209);
    layer0_outputs(747) <= (inputs(107)) or (inputs(207));
    layer0_outputs(748) <= inputs(82);
    layer0_outputs(749) <= not(inputs(60));
    layer0_outputs(750) <= inputs(226);
    layer0_outputs(751) <= inputs(110);
    layer0_outputs(752) <= '1';
    layer0_outputs(753) <= (inputs(42)) or (inputs(48));
    layer0_outputs(754) <= not(inputs(123));
    layer0_outputs(755) <= not(inputs(211)) or (inputs(119));
    layer0_outputs(756) <= not((inputs(68)) or (inputs(94)));
    layer0_outputs(757) <= (inputs(138)) or (inputs(254));
    layer0_outputs(758) <= not(inputs(178));
    layer0_outputs(759) <= not((inputs(141)) and (inputs(104)));
    layer0_outputs(760) <= not(inputs(14)) or (inputs(87));
    layer0_outputs(761) <= inputs(10);
    layer0_outputs(762) <= not(inputs(169));
    layer0_outputs(763) <= not((inputs(135)) or (inputs(253)));
    layer0_outputs(764) <= not(inputs(189)) or (inputs(132));
    layer0_outputs(765) <= not((inputs(163)) or (inputs(21)));
    layer0_outputs(766) <= '1';
    layer0_outputs(767) <= not(inputs(102));
    layer0_outputs(768) <= not((inputs(58)) and (inputs(39)));
    layer0_outputs(769) <= (inputs(11)) xor (inputs(41));
    layer0_outputs(770) <= not(inputs(147));
    layer0_outputs(771) <= not(inputs(72));
    layer0_outputs(772) <= (inputs(216)) and not (inputs(47));
    layer0_outputs(773) <= (inputs(248)) or (inputs(142));
    layer0_outputs(774) <= inputs(113);
    layer0_outputs(775) <= not(inputs(211));
    layer0_outputs(776) <= (inputs(66)) xor (inputs(70));
    layer0_outputs(777) <= not(inputs(89)) or (inputs(163));
    layer0_outputs(778) <= (inputs(101)) xor (inputs(132));
    layer0_outputs(779) <= (inputs(119)) or (inputs(222));
    layer0_outputs(780) <= not(inputs(121));
    layer0_outputs(781) <= not(inputs(234));
    layer0_outputs(782) <= (inputs(128)) or (inputs(187));
    layer0_outputs(783) <= (inputs(147)) and not (inputs(18));
    layer0_outputs(784) <= not(inputs(9));
    layer0_outputs(785) <= inputs(95);
    layer0_outputs(786) <= not((inputs(242)) or (inputs(33)));
    layer0_outputs(787) <= inputs(188);
    layer0_outputs(788) <= inputs(28);
    layer0_outputs(789) <= inputs(135);
    layer0_outputs(790) <= not(inputs(168)) or (inputs(41));
    layer0_outputs(791) <= not((inputs(94)) xor (inputs(66)));
    layer0_outputs(792) <= '0';
    layer0_outputs(793) <= (inputs(142)) and not (inputs(240));
    layer0_outputs(794) <= '0';
    layer0_outputs(795) <= not(inputs(157));
    layer0_outputs(796) <= (inputs(255)) and not (inputs(241));
    layer0_outputs(797) <= '0';
    layer0_outputs(798) <= (inputs(153)) and not (inputs(9));
    layer0_outputs(799) <= not((inputs(65)) or (inputs(79)));
    layer0_outputs(800) <= not(inputs(189));
    layer0_outputs(801) <= (inputs(200)) or (inputs(208));
    layer0_outputs(802) <= inputs(228);
    layer0_outputs(803) <= not(inputs(147));
    layer0_outputs(804) <= not((inputs(215)) or (inputs(179)));
    layer0_outputs(805) <= (inputs(114)) or (inputs(37));
    layer0_outputs(806) <= (inputs(81)) and not (inputs(250));
    layer0_outputs(807) <= '1';
    layer0_outputs(808) <= not(inputs(226)) or (inputs(45));
    layer0_outputs(809) <= '0';
    layer0_outputs(810) <= (inputs(7)) or (inputs(208));
    layer0_outputs(811) <= (inputs(13)) and (inputs(1));
    layer0_outputs(812) <= (inputs(252)) and (inputs(9));
    layer0_outputs(813) <= not(inputs(127));
    layer0_outputs(814) <= not(inputs(181));
    layer0_outputs(815) <= not(inputs(109));
    layer0_outputs(816) <= inputs(231);
    layer0_outputs(817) <= not(inputs(175));
    layer0_outputs(818) <= not(inputs(204));
    layer0_outputs(819) <= (inputs(36)) or (inputs(111));
    layer0_outputs(820) <= inputs(105);
    layer0_outputs(821) <= (inputs(31)) and (inputs(202));
    layer0_outputs(822) <= not(inputs(74));
    layer0_outputs(823) <= inputs(187);
    layer0_outputs(824) <= not((inputs(35)) or (inputs(43)));
    layer0_outputs(825) <= not((inputs(249)) and (inputs(193)));
    layer0_outputs(826) <= inputs(248);
    layer0_outputs(827) <= (inputs(13)) and (inputs(35));
    layer0_outputs(828) <= (inputs(10)) and not (inputs(159));
    layer0_outputs(829) <= '0';
    layer0_outputs(830) <= (inputs(152)) and not (inputs(1));
    layer0_outputs(831) <= inputs(120);
    layer0_outputs(832) <= inputs(196);
    layer0_outputs(833) <= not((inputs(226)) or (inputs(233)));
    layer0_outputs(834) <= not((inputs(4)) or (inputs(38)));
    layer0_outputs(835) <= '1';
    layer0_outputs(836) <= (inputs(30)) or (inputs(219));
    layer0_outputs(837) <= not(inputs(253)) or (inputs(52));
    layer0_outputs(838) <= not((inputs(140)) or (inputs(158)));
    layer0_outputs(839) <= not(inputs(206));
    layer0_outputs(840) <= not((inputs(190)) or (inputs(217)));
    layer0_outputs(841) <= (inputs(10)) and not (inputs(144));
    layer0_outputs(842) <= '0';
    layer0_outputs(843) <= not(inputs(50));
    layer0_outputs(844) <= inputs(78);
    layer0_outputs(845) <= (inputs(227)) or (inputs(134));
    layer0_outputs(846) <= not(inputs(136));
    layer0_outputs(847) <= not(inputs(28));
    layer0_outputs(848) <= '1';
    layer0_outputs(849) <= (inputs(20)) or (inputs(191));
    layer0_outputs(850) <= not(inputs(230)) or (inputs(84));
    layer0_outputs(851) <= not(inputs(128));
    layer0_outputs(852) <= (inputs(105)) and not (inputs(193));
    layer0_outputs(853) <= '1';
    layer0_outputs(854) <= not((inputs(143)) or (inputs(156)));
    layer0_outputs(855) <= not(inputs(75)) or (inputs(103));
    layer0_outputs(856) <= not(inputs(167));
    layer0_outputs(857) <= (inputs(192)) or (inputs(241));
    layer0_outputs(858) <= not(inputs(91));
    layer0_outputs(859) <= (inputs(84)) and not (inputs(107));
    layer0_outputs(860) <= not(inputs(175));
    layer0_outputs(861) <= not(inputs(60));
    layer0_outputs(862) <= inputs(40);
    layer0_outputs(863) <= (inputs(187)) or (inputs(127));
    layer0_outputs(864) <= not((inputs(54)) or (inputs(98)));
    layer0_outputs(865) <= not((inputs(158)) or (inputs(208)));
    layer0_outputs(866) <= not(inputs(86)) or (inputs(34));
    layer0_outputs(867) <= not((inputs(15)) or (inputs(69)));
    layer0_outputs(868) <= not((inputs(99)) and (inputs(211)));
    layer0_outputs(869) <= '1';
    layer0_outputs(870) <= (inputs(85)) xor (inputs(189));
    layer0_outputs(871) <= not((inputs(194)) or (inputs(162)));
    layer0_outputs(872) <= not(inputs(193)) or (inputs(143));
    layer0_outputs(873) <= inputs(156);
    layer0_outputs(874) <= not((inputs(205)) or (inputs(215)));
    layer0_outputs(875) <= not(inputs(138));
    layer0_outputs(876) <= not(inputs(104)) or (inputs(110));
    layer0_outputs(877) <= inputs(230);
    layer0_outputs(878) <= not((inputs(129)) or (inputs(30)));
    layer0_outputs(879) <= not(inputs(148));
    layer0_outputs(880) <= not((inputs(209)) or (inputs(244)));
    layer0_outputs(881) <= not(inputs(91));
    layer0_outputs(882) <= inputs(2);
    layer0_outputs(883) <= inputs(239);
    layer0_outputs(884) <= (inputs(162)) and not (inputs(149));
    layer0_outputs(885) <= inputs(41);
    layer0_outputs(886) <= not(inputs(28));
    layer0_outputs(887) <= inputs(23);
    layer0_outputs(888) <= (inputs(49)) or (inputs(195));
    layer0_outputs(889) <= (inputs(229)) and not (inputs(60));
    layer0_outputs(890) <= '0';
    layer0_outputs(891) <= (inputs(109)) or (inputs(56));
    layer0_outputs(892) <= not((inputs(129)) xor (inputs(147)));
    layer0_outputs(893) <= '1';
    layer0_outputs(894) <= not(inputs(212));
    layer0_outputs(895) <= inputs(76);
    layer0_outputs(896) <= not((inputs(132)) or (inputs(114)));
    layer0_outputs(897) <= inputs(61);
    layer0_outputs(898) <= not(inputs(70)) or (inputs(125));
    layer0_outputs(899) <= (inputs(53)) and not (inputs(62));
    layer0_outputs(900) <= not((inputs(239)) or (inputs(164)));
    layer0_outputs(901) <= (inputs(234)) or (inputs(217));
    layer0_outputs(902) <= not(inputs(126)) or (inputs(222));
    layer0_outputs(903) <= not((inputs(210)) xor (inputs(126)));
    layer0_outputs(904) <= (inputs(228)) and not (inputs(95));
    layer0_outputs(905) <= (inputs(216)) xor (inputs(248));
    layer0_outputs(906) <= not((inputs(224)) or (inputs(12)));
    layer0_outputs(907) <= inputs(97);
    layer0_outputs(908) <= (inputs(33)) and not (inputs(131));
    layer0_outputs(909) <= not((inputs(123)) or (inputs(140)));
    layer0_outputs(910) <= inputs(70);
    layer0_outputs(911) <= not(inputs(163));
    layer0_outputs(912) <= not((inputs(83)) and (inputs(157)));
    layer0_outputs(913) <= not((inputs(238)) or (inputs(10)));
    layer0_outputs(914) <= (inputs(123)) and not (inputs(43));
    layer0_outputs(915) <= not((inputs(159)) or (inputs(54)));
    layer0_outputs(916) <= (inputs(144)) and not (inputs(105));
    layer0_outputs(917) <= inputs(7);
    layer0_outputs(918) <= not(inputs(21)) or (inputs(226));
    layer0_outputs(919) <= (inputs(248)) or (inputs(148));
    layer0_outputs(920) <= (inputs(227)) and not (inputs(192));
    layer0_outputs(921) <= (inputs(105)) and not (inputs(48));
    layer0_outputs(922) <= (inputs(82)) and not (inputs(140));
    layer0_outputs(923) <= not(inputs(248)) or (inputs(125));
    layer0_outputs(924) <= inputs(177);
    layer0_outputs(925) <= (inputs(112)) or (inputs(124));
    layer0_outputs(926) <= not((inputs(125)) or (inputs(6)));
    layer0_outputs(927) <= (inputs(65)) and not (inputs(169));
    layer0_outputs(928) <= not(inputs(7));
    layer0_outputs(929) <= (inputs(73)) and not (inputs(5));
    layer0_outputs(930) <= inputs(147);
    layer0_outputs(931) <= inputs(52);
    layer0_outputs(932) <= '0';
    layer0_outputs(933) <= '0';
    layer0_outputs(934) <= inputs(114);
    layer0_outputs(935) <= inputs(166);
    layer0_outputs(936) <= not((inputs(36)) or (inputs(3)));
    layer0_outputs(937) <= (inputs(100)) and not (inputs(77));
    layer0_outputs(938) <= not((inputs(236)) xor (inputs(80)));
    layer0_outputs(939) <= not((inputs(249)) or (inputs(12)));
    layer0_outputs(940) <= (inputs(17)) or (inputs(227));
    layer0_outputs(941) <= not(inputs(152)) or (inputs(123));
    layer0_outputs(942) <= inputs(119);
    layer0_outputs(943) <= '1';
    layer0_outputs(944) <= inputs(213);
    layer0_outputs(945) <= not(inputs(214)) or (inputs(183));
    layer0_outputs(946) <= (inputs(69)) and not (inputs(206));
    layer0_outputs(947) <= not((inputs(15)) or (inputs(53)));
    layer0_outputs(948) <= not(inputs(31));
    layer0_outputs(949) <= inputs(69);
    layer0_outputs(950) <= inputs(162);
    layer0_outputs(951) <= not((inputs(232)) and (inputs(71)));
    layer0_outputs(952) <= not((inputs(52)) or (inputs(33)));
    layer0_outputs(953) <= not((inputs(64)) and (inputs(124)));
    layer0_outputs(954) <= '1';
    layer0_outputs(955) <= not(inputs(146));
    layer0_outputs(956) <= not(inputs(43)) or (inputs(179));
    layer0_outputs(957) <= not(inputs(212));
    layer0_outputs(958) <= inputs(158);
    layer0_outputs(959) <= (inputs(137)) and not (inputs(120));
    layer0_outputs(960) <= '0';
    layer0_outputs(961) <= inputs(86);
    layer0_outputs(962) <= '0';
    layer0_outputs(963) <= '0';
    layer0_outputs(964) <= not(inputs(136));
    layer0_outputs(965) <= not(inputs(165));
    layer0_outputs(966) <= not((inputs(253)) or (inputs(11)));
    layer0_outputs(967) <= not(inputs(138));
    layer0_outputs(968) <= not(inputs(246));
    layer0_outputs(969) <= not((inputs(246)) or (inputs(110)));
    layer0_outputs(970) <= inputs(98);
    layer0_outputs(971) <= inputs(120);
    layer0_outputs(972) <= not(inputs(48)) or (inputs(101));
    layer0_outputs(973) <= not(inputs(231));
    layer0_outputs(974) <= (inputs(89)) or (inputs(92));
    layer0_outputs(975) <= not(inputs(54)) or (inputs(105));
    layer0_outputs(976) <= not(inputs(223));
    layer0_outputs(977) <= not(inputs(41));
    layer0_outputs(978) <= not((inputs(129)) or (inputs(124)));
    layer0_outputs(979) <= not(inputs(240));
    layer0_outputs(980) <= (inputs(195)) and (inputs(246));
    layer0_outputs(981) <= (inputs(50)) or (inputs(92));
    layer0_outputs(982) <= not(inputs(176)) or (inputs(176));
    layer0_outputs(983) <= not((inputs(113)) or (inputs(98)));
    layer0_outputs(984) <= not(inputs(83));
    layer0_outputs(985) <= '0';
    layer0_outputs(986) <= not(inputs(131));
    layer0_outputs(987) <= inputs(138);
    layer0_outputs(988) <= not((inputs(182)) or (inputs(101)));
    layer0_outputs(989) <= not(inputs(40));
    layer0_outputs(990) <= not(inputs(236));
    layer0_outputs(991) <= not(inputs(122));
    layer0_outputs(992) <= not((inputs(194)) or (inputs(193)));
    layer0_outputs(993) <= '1';
    layer0_outputs(994) <= inputs(177);
    layer0_outputs(995) <= not(inputs(132));
    layer0_outputs(996) <= not((inputs(235)) or (inputs(135)));
    layer0_outputs(997) <= '1';
    layer0_outputs(998) <= not(inputs(103));
    layer0_outputs(999) <= (inputs(233)) or (inputs(192));
    layer0_outputs(1000) <= (inputs(131)) and not (inputs(66));
    layer0_outputs(1001) <= not(inputs(116));
    layer0_outputs(1002) <= not(inputs(113));
    layer0_outputs(1003) <= not(inputs(145));
    layer0_outputs(1004) <= not((inputs(53)) and (inputs(244)));
    layer0_outputs(1005) <= not(inputs(3));
    layer0_outputs(1006) <= inputs(167);
    layer0_outputs(1007) <= not((inputs(96)) or (inputs(199)));
    layer0_outputs(1008) <= inputs(182);
    layer0_outputs(1009) <= not(inputs(97));
    layer0_outputs(1010) <= not(inputs(165));
    layer0_outputs(1011) <= not((inputs(173)) or (inputs(95)));
    layer0_outputs(1012) <= inputs(76);
    layer0_outputs(1013) <= (inputs(223)) or (inputs(150));
    layer0_outputs(1014) <= inputs(244);
    layer0_outputs(1015) <= inputs(73);
    layer0_outputs(1016) <= '1';
    layer0_outputs(1017) <= (inputs(91)) or (inputs(63));
    layer0_outputs(1018) <= inputs(154);
    layer0_outputs(1019) <= '1';
    layer0_outputs(1020) <= not(inputs(66));
    layer0_outputs(1021) <= not(inputs(229)) or (inputs(135));
    layer0_outputs(1022) <= inputs(147);
    layer0_outputs(1023) <= not((inputs(34)) or (inputs(40)));
    layer0_outputs(1024) <= inputs(119);
    layer0_outputs(1025) <= inputs(137);
    layer0_outputs(1026) <= (inputs(208)) or (inputs(9));
    layer0_outputs(1027) <= '0';
    layer0_outputs(1028) <= inputs(177);
    layer0_outputs(1029) <= (inputs(93)) or (inputs(156));
    layer0_outputs(1030) <= not(inputs(39)) or (inputs(56));
    layer0_outputs(1031) <= (inputs(160)) or (inputs(140));
    layer0_outputs(1032) <= inputs(169);
    layer0_outputs(1033) <= not((inputs(36)) or (inputs(94)));
    layer0_outputs(1034) <= not(inputs(27)) or (inputs(193));
    layer0_outputs(1035) <= not(inputs(200)) or (inputs(174));
    layer0_outputs(1036) <= inputs(85);
    layer0_outputs(1037) <= not(inputs(234));
    layer0_outputs(1038) <= not(inputs(209)) or (inputs(247));
    layer0_outputs(1039) <= (inputs(8)) or (inputs(57));
    layer0_outputs(1040) <= not((inputs(38)) or (inputs(75)));
    layer0_outputs(1041) <= (inputs(132)) or (inputs(18));
    layer0_outputs(1042) <= (inputs(45)) and not (inputs(255));
    layer0_outputs(1043) <= (inputs(13)) and not (inputs(254));
    layer0_outputs(1044) <= '0';
    layer0_outputs(1045) <= not(inputs(59));
    layer0_outputs(1046) <= not(inputs(187));
    layer0_outputs(1047) <= not(inputs(101)) or (inputs(1));
    layer0_outputs(1048) <= not(inputs(117)) or (inputs(254));
    layer0_outputs(1049) <= inputs(124);
    layer0_outputs(1050) <= inputs(83);
    layer0_outputs(1051) <= inputs(246);
    layer0_outputs(1052) <= not(inputs(92)) or (inputs(183));
    layer0_outputs(1053) <= (inputs(41)) and not (inputs(118));
    layer0_outputs(1054) <= '0';
    layer0_outputs(1055) <= not((inputs(225)) and (inputs(46)));
    layer0_outputs(1056) <= inputs(118);
    layer0_outputs(1057) <= not(inputs(163)) or (inputs(240));
    layer0_outputs(1058) <= inputs(107);
    layer0_outputs(1059) <= (inputs(160)) or (inputs(65));
    layer0_outputs(1060) <= not(inputs(108));
    layer0_outputs(1061) <= '0';
    layer0_outputs(1062) <= (inputs(192)) and not (inputs(82));
    layer0_outputs(1063) <= not((inputs(242)) and (inputs(250)));
    layer0_outputs(1064) <= (inputs(193)) xor (inputs(175));
    layer0_outputs(1065) <= inputs(84);
    layer0_outputs(1066) <= '1';
    layer0_outputs(1067) <= not((inputs(253)) or (inputs(167)));
    layer0_outputs(1068) <= (inputs(26)) and not (inputs(142));
    layer0_outputs(1069) <= inputs(233);
    layer0_outputs(1070) <= not((inputs(0)) or (inputs(202)));
    layer0_outputs(1071) <= not((inputs(29)) or (inputs(60)));
    layer0_outputs(1072) <= (inputs(117)) and not (inputs(222));
    layer0_outputs(1073) <= not(inputs(164));
    layer0_outputs(1074) <= (inputs(13)) or (inputs(74));
    layer0_outputs(1075) <= inputs(148);
    layer0_outputs(1076) <= not(inputs(103)) or (inputs(52));
    layer0_outputs(1077) <= not(inputs(7)) or (inputs(50));
    layer0_outputs(1078) <= not(inputs(41)) or (inputs(163));
    layer0_outputs(1079) <= (inputs(71)) and not (inputs(222));
    layer0_outputs(1080) <= inputs(11);
    layer0_outputs(1081) <= (inputs(189)) or (inputs(167));
    layer0_outputs(1082) <= not(inputs(203)) or (inputs(14));
    layer0_outputs(1083) <= not((inputs(126)) and (inputs(183)));
    layer0_outputs(1084) <= (inputs(165)) and not (inputs(96));
    layer0_outputs(1085) <= not((inputs(122)) or (inputs(17)));
    layer0_outputs(1086) <= inputs(172);
    layer0_outputs(1087) <= (inputs(5)) and not (inputs(239));
    layer0_outputs(1088) <= (inputs(110)) or (inputs(23));
    layer0_outputs(1089) <= '0';
    layer0_outputs(1090) <= not((inputs(222)) or (inputs(232)));
    layer0_outputs(1091) <= (inputs(87)) and not (inputs(157));
    layer0_outputs(1092) <= not(inputs(151)) or (inputs(80));
    layer0_outputs(1093) <= '0';
    layer0_outputs(1094) <= not(inputs(125)) or (inputs(3));
    layer0_outputs(1095) <= (inputs(220)) and not (inputs(227));
    layer0_outputs(1096) <= (inputs(112)) or (inputs(139));
    layer0_outputs(1097) <= '0';
    layer0_outputs(1098) <= not(inputs(160));
    layer0_outputs(1099) <= inputs(165);
    layer0_outputs(1100) <= inputs(101);
    layer0_outputs(1101) <= inputs(23);
    layer0_outputs(1102) <= not(inputs(96));
    layer0_outputs(1103) <= not((inputs(72)) or (inputs(239)));
    layer0_outputs(1104) <= '0';
    layer0_outputs(1105) <= inputs(88);
    layer0_outputs(1106) <= (inputs(209)) or (inputs(174));
    layer0_outputs(1107) <= (inputs(130)) and not (inputs(57));
    layer0_outputs(1108) <= not(inputs(158));
    layer0_outputs(1109) <= not(inputs(105));
    layer0_outputs(1110) <= not(inputs(68));
    layer0_outputs(1111) <= '0';
    layer0_outputs(1112) <= not(inputs(21));
    layer0_outputs(1113) <= (inputs(202)) and not (inputs(85));
    layer0_outputs(1114) <= (inputs(148)) and not (inputs(237));
    layer0_outputs(1115) <= (inputs(64)) or (inputs(225));
    layer0_outputs(1116) <= not((inputs(60)) or (inputs(170)));
    layer0_outputs(1117) <= inputs(72);
    layer0_outputs(1118) <= (inputs(24)) or (inputs(30));
    layer0_outputs(1119) <= not(inputs(162));
    layer0_outputs(1120) <= not((inputs(163)) or (inputs(180)));
    layer0_outputs(1121) <= inputs(178);
    layer0_outputs(1122) <= not(inputs(71));
    layer0_outputs(1123) <= not(inputs(143));
    layer0_outputs(1124) <= '0';
    layer0_outputs(1125) <= not((inputs(221)) or (inputs(192)));
    layer0_outputs(1126) <= not(inputs(235)) or (inputs(15));
    layer0_outputs(1127) <= '1';
    layer0_outputs(1128) <= (inputs(72)) and (inputs(154));
    layer0_outputs(1129) <= not((inputs(24)) or (inputs(158)));
    layer0_outputs(1130) <= not(inputs(90)) or (inputs(157));
    layer0_outputs(1131) <= not(inputs(66)) or (inputs(156));
    layer0_outputs(1132) <= not((inputs(207)) and (inputs(225)));
    layer0_outputs(1133) <= not(inputs(189)) or (inputs(101));
    layer0_outputs(1134) <= inputs(144);
    layer0_outputs(1135) <= not((inputs(245)) and (inputs(6)));
    layer0_outputs(1136) <= (inputs(206)) xor (inputs(139));
    layer0_outputs(1137) <= not(inputs(100));
    layer0_outputs(1138) <= (inputs(5)) or (inputs(59));
    layer0_outputs(1139) <= (inputs(209)) or (inputs(194));
    layer0_outputs(1140) <= inputs(188);
    layer0_outputs(1141) <= (inputs(40)) and not (inputs(162));
    layer0_outputs(1142) <= not((inputs(49)) or (inputs(67)));
    layer0_outputs(1143) <= (inputs(19)) or (inputs(61));
    layer0_outputs(1144) <= (inputs(32)) or (inputs(174));
    layer0_outputs(1145) <= not(inputs(26)) or (inputs(168));
    layer0_outputs(1146) <= inputs(174);
    layer0_outputs(1147) <= not(inputs(196));
    layer0_outputs(1148) <= (inputs(124)) and (inputs(35));
    layer0_outputs(1149) <= not(inputs(212)) or (inputs(52));
    layer0_outputs(1150) <= not((inputs(86)) or (inputs(176)));
    layer0_outputs(1151) <= inputs(136);
    layer0_outputs(1152) <= (inputs(27)) or (inputs(58));
    layer0_outputs(1153) <= (inputs(55)) and (inputs(187));
    layer0_outputs(1154) <= not(inputs(203)) or (inputs(34));
    layer0_outputs(1155) <= not(inputs(254));
    layer0_outputs(1156) <= not(inputs(59)) or (inputs(231));
    layer0_outputs(1157) <= not((inputs(95)) or (inputs(46)));
    layer0_outputs(1158) <= '1';
    layer0_outputs(1159) <= not(inputs(112)) or (inputs(27));
    layer0_outputs(1160) <= (inputs(91)) and not (inputs(59));
    layer0_outputs(1161) <= '1';
    layer0_outputs(1162) <= (inputs(93)) and not (inputs(251));
    layer0_outputs(1163) <= not((inputs(87)) or (inputs(132)));
    layer0_outputs(1164) <= not(inputs(62));
    layer0_outputs(1165) <= (inputs(173)) or (inputs(93));
    layer0_outputs(1166) <= not((inputs(240)) and (inputs(187)));
    layer0_outputs(1167) <= not(inputs(91));
    layer0_outputs(1168) <= not((inputs(237)) or (inputs(138)));
    layer0_outputs(1169) <= inputs(228);
    layer0_outputs(1170) <= not(inputs(217)) or (inputs(35));
    layer0_outputs(1171) <= '0';
    layer0_outputs(1172) <= inputs(7);
    layer0_outputs(1173) <= '1';
    layer0_outputs(1174) <= not(inputs(212));
    layer0_outputs(1175) <= inputs(101);
    layer0_outputs(1176) <= not(inputs(161));
    layer0_outputs(1177) <= '0';
    layer0_outputs(1178) <= inputs(226);
    layer0_outputs(1179) <= not(inputs(131)) or (inputs(205));
    layer0_outputs(1180) <= (inputs(36)) and not (inputs(98));
    layer0_outputs(1181) <= (inputs(124)) or (inputs(5));
    layer0_outputs(1182) <= inputs(31);
    layer0_outputs(1183) <= not((inputs(158)) or (inputs(76)));
    layer0_outputs(1184) <= inputs(181);
    layer0_outputs(1185) <= inputs(122);
    layer0_outputs(1186) <= not((inputs(236)) or (inputs(34)));
    layer0_outputs(1187) <= not(inputs(143));
    layer0_outputs(1188) <= inputs(176);
    layer0_outputs(1189) <= inputs(74);
    layer0_outputs(1190) <= not(inputs(36));
    layer0_outputs(1191) <= (inputs(140)) and (inputs(43));
    layer0_outputs(1192) <= inputs(100);
    layer0_outputs(1193) <= not(inputs(115));
    layer0_outputs(1194) <= not(inputs(90));
    layer0_outputs(1195) <= not(inputs(147)) or (inputs(63));
    layer0_outputs(1196) <= (inputs(46)) and not (inputs(241));
    layer0_outputs(1197) <= not(inputs(121));
    layer0_outputs(1198) <= (inputs(116)) or (inputs(133));
    layer0_outputs(1199) <= not((inputs(16)) or (inputs(33)));
    layer0_outputs(1200) <= not((inputs(111)) or (inputs(78)));
    layer0_outputs(1201) <= (inputs(16)) and not (inputs(96));
    layer0_outputs(1202) <= inputs(131);
    layer0_outputs(1203) <= (inputs(1)) or (inputs(199));
    layer0_outputs(1204) <= not(inputs(148));
    layer0_outputs(1205) <= (inputs(116)) and not (inputs(207));
    layer0_outputs(1206) <= inputs(194);
    layer0_outputs(1207) <= '1';
    layer0_outputs(1208) <= not(inputs(185)) or (inputs(248));
    layer0_outputs(1209) <= (inputs(11)) or (inputs(92));
    layer0_outputs(1210) <= (inputs(237)) and (inputs(185));
    layer0_outputs(1211) <= inputs(150);
    layer0_outputs(1212) <= not(inputs(145));
    layer0_outputs(1213) <= not(inputs(2));
    layer0_outputs(1214) <= (inputs(41)) and not (inputs(252));
    layer0_outputs(1215) <= inputs(97);
    layer0_outputs(1216) <= not(inputs(61));
    layer0_outputs(1217) <= not((inputs(247)) or (inputs(156)));
    layer0_outputs(1218) <= not(inputs(195));
    layer0_outputs(1219) <= inputs(58);
    layer0_outputs(1220) <= not(inputs(184));
    layer0_outputs(1221) <= not(inputs(80));
    layer0_outputs(1222) <= not(inputs(207));
    layer0_outputs(1223) <= not((inputs(117)) and (inputs(31)));
    layer0_outputs(1224) <= inputs(252);
    layer0_outputs(1225) <= not((inputs(207)) or (inputs(108)));
    layer0_outputs(1226) <= inputs(133);
    layer0_outputs(1227) <= not((inputs(93)) or (inputs(23)));
    layer0_outputs(1228) <= not((inputs(227)) or (inputs(224)));
    layer0_outputs(1229) <= not(inputs(216)) or (inputs(176));
    layer0_outputs(1230) <= (inputs(227)) xor (inputs(242));
    layer0_outputs(1231) <= not((inputs(189)) or (inputs(48)));
    layer0_outputs(1232) <= not(inputs(70));
    layer0_outputs(1233) <= '0';
    layer0_outputs(1234) <= not(inputs(90));
    layer0_outputs(1235) <= not((inputs(119)) or (inputs(162)));
    layer0_outputs(1236) <= (inputs(158)) xor (inputs(141));
    layer0_outputs(1237) <= not(inputs(233));
    layer0_outputs(1238) <= not(inputs(211));
    layer0_outputs(1239) <= (inputs(91)) and not (inputs(97));
    layer0_outputs(1240) <= (inputs(166)) or (inputs(163));
    layer0_outputs(1241) <= inputs(136);
    layer0_outputs(1242) <= (inputs(152)) and (inputs(189));
    layer0_outputs(1243) <= not(inputs(113));
    layer0_outputs(1244) <= not(inputs(203)) or (inputs(93));
    layer0_outputs(1245) <= '0';
    layer0_outputs(1246) <= (inputs(197)) and not (inputs(193));
    layer0_outputs(1247) <= not((inputs(9)) or (inputs(202)));
    layer0_outputs(1248) <= inputs(40);
    layer0_outputs(1249) <= (inputs(63)) and not (inputs(13));
    layer0_outputs(1250) <= not((inputs(190)) or (inputs(244)));
    layer0_outputs(1251) <= not(inputs(179));
    layer0_outputs(1252) <= inputs(62);
    layer0_outputs(1253) <= not(inputs(51)) or (inputs(225));
    layer0_outputs(1254) <= not((inputs(106)) or (inputs(208)));
    layer0_outputs(1255) <= (inputs(126)) and not (inputs(223));
    layer0_outputs(1256) <= inputs(203);
    layer0_outputs(1257) <= not(inputs(125));
    layer0_outputs(1258) <= (inputs(207)) or (inputs(16));
    layer0_outputs(1259) <= '0';
    layer0_outputs(1260) <= inputs(22);
    layer0_outputs(1261) <= '0';
    layer0_outputs(1262) <= (inputs(30)) or (inputs(44));
    layer0_outputs(1263) <= (inputs(36)) and not (inputs(217));
    layer0_outputs(1264) <= inputs(22);
    layer0_outputs(1265) <= not(inputs(51)) or (inputs(246));
    layer0_outputs(1266) <= '1';
    layer0_outputs(1267) <= not((inputs(168)) and (inputs(222)));
    layer0_outputs(1268) <= not((inputs(26)) or (inputs(218)));
    layer0_outputs(1269) <= (inputs(100)) or (inputs(70));
    layer0_outputs(1270) <= (inputs(34)) and not (inputs(34));
    layer0_outputs(1271) <= not(inputs(0));
    layer0_outputs(1272) <= (inputs(134)) or (inputs(218));
    layer0_outputs(1273) <= (inputs(171)) xor (inputs(219));
    layer0_outputs(1274) <= (inputs(241)) or (inputs(222));
    layer0_outputs(1275) <= not(inputs(98));
    layer0_outputs(1276) <= not(inputs(199));
    layer0_outputs(1277) <= (inputs(168)) or (inputs(48));
    layer0_outputs(1278) <= not(inputs(24));
    layer0_outputs(1279) <= (inputs(63)) and (inputs(154));
    layer0_outputs(1280) <= not((inputs(1)) or (inputs(219)));
    layer0_outputs(1281) <= not((inputs(219)) or (inputs(222)));
    layer0_outputs(1282) <= not(inputs(246)) or (inputs(74));
    layer0_outputs(1283) <= not(inputs(37));
    layer0_outputs(1284) <= not(inputs(232));
    layer0_outputs(1285) <= inputs(164);
    layer0_outputs(1286) <= not((inputs(61)) or (inputs(230)));
    layer0_outputs(1287) <= not(inputs(172));
    layer0_outputs(1288) <= not((inputs(232)) or (inputs(179)));
    layer0_outputs(1289) <= (inputs(39)) and not (inputs(19));
    layer0_outputs(1290) <= not((inputs(82)) or (inputs(183)));
    layer0_outputs(1291) <= (inputs(53)) or (inputs(108));
    layer0_outputs(1292) <= not((inputs(254)) or (inputs(132)));
    layer0_outputs(1293) <= not(inputs(21));
    layer0_outputs(1294) <= not(inputs(59)) or (inputs(145));
    layer0_outputs(1295) <= not(inputs(68));
    layer0_outputs(1296) <= inputs(24);
    layer0_outputs(1297) <= '0';
    layer0_outputs(1298) <= not((inputs(2)) or (inputs(220)));
    layer0_outputs(1299) <= not((inputs(211)) or (inputs(246)));
    layer0_outputs(1300) <= (inputs(157)) and not (inputs(67));
    layer0_outputs(1301) <= not((inputs(65)) or (inputs(84)));
    layer0_outputs(1302) <= (inputs(0)) or (inputs(127));
    layer0_outputs(1303) <= not(inputs(68)) or (inputs(242));
    layer0_outputs(1304) <= not((inputs(136)) and (inputs(132)));
    layer0_outputs(1305) <= not(inputs(230)) or (inputs(92));
    layer0_outputs(1306) <= not((inputs(66)) or (inputs(160)));
    layer0_outputs(1307) <= '1';
    layer0_outputs(1308) <= not(inputs(99));
    layer0_outputs(1309) <= not((inputs(158)) or (inputs(213)));
    layer0_outputs(1310) <= (inputs(166)) xor (inputs(164));
    layer0_outputs(1311) <= (inputs(128)) and (inputs(253));
    layer0_outputs(1312) <= '0';
    layer0_outputs(1313) <= (inputs(121)) and (inputs(172));
    layer0_outputs(1314) <= not(inputs(39));
    layer0_outputs(1315) <= not(inputs(75)) or (inputs(126));
    layer0_outputs(1316) <= not(inputs(230));
    layer0_outputs(1317) <= not((inputs(64)) and (inputs(127)));
    layer0_outputs(1318) <= inputs(147);
    layer0_outputs(1319) <= '0';
    layer0_outputs(1320) <= not((inputs(169)) or (inputs(198)));
    layer0_outputs(1321) <= not(inputs(74));
    layer0_outputs(1322) <= not((inputs(141)) or (inputs(193)));
    layer0_outputs(1323) <= '0';
    layer0_outputs(1324) <= inputs(217);
    layer0_outputs(1325) <= not((inputs(33)) or (inputs(128)));
    layer0_outputs(1326) <= not(inputs(87)) or (inputs(36));
    layer0_outputs(1327) <= '1';
    layer0_outputs(1328) <= inputs(88);
    layer0_outputs(1329) <= '1';
    layer0_outputs(1330) <= inputs(189);
    layer0_outputs(1331) <= not((inputs(141)) or (inputs(144)));
    layer0_outputs(1332) <= (inputs(195)) or (inputs(214));
    layer0_outputs(1333) <= not((inputs(4)) or (inputs(139)));
    layer0_outputs(1334) <= (inputs(71)) and not (inputs(85));
    layer0_outputs(1335) <= not((inputs(80)) and (inputs(150)));
    layer0_outputs(1336) <= not((inputs(73)) and (inputs(22)));
    layer0_outputs(1337) <= not(inputs(178));
    layer0_outputs(1338) <= not(inputs(34));
    layer0_outputs(1339) <= not(inputs(105));
    layer0_outputs(1340) <= inputs(83);
    layer0_outputs(1341) <= not(inputs(227));
    layer0_outputs(1342) <= inputs(125);
    layer0_outputs(1343) <= not((inputs(204)) or (inputs(220)));
    layer0_outputs(1344) <= not(inputs(66));
    layer0_outputs(1345) <= not((inputs(195)) or (inputs(27)));
    layer0_outputs(1346) <= (inputs(223)) or (inputs(241));
    layer0_outputs(1347) <= (inputs(28)) and not (inputs(186));
    layer0_outputs(1348) <= (inputs(145)) or (inputs(179));
    layer0_outputs(1349) <= inputs(251);
    layer0_outputs(1350) <= (inputs(145)) or (inputs(238));
    layer0_outputs(1351) <= inputs(252);
    layer0_outputs(1352) <= not(inputs(145));
    layer0_outputs(1353) <= not(inputs(244));
    layer0_outputs(1354) <= '0';
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= not(inputs(158)) or (inputs(241));
    layer0_outputs(1357) <= (inputs(88)) and not (inputs(221));
    layer0_outputs(1358) <= not((inputs(210)) or (inputs(24)));
    layer0_outputs(1359) <= inputs(180);
    layer0_outputs(1360) <= not((inputs(173)) or (inputs(22)));
    layer0_outputs(1361) <= (inputs(32)) or (inputs(218));
    layer0_outputs(1362) <= not(inputs(178));
    layer0_outputs(1363) <= inputs(35);
    layer0_outputs(1364) <= not((inputs(177)) or (inputs(221)));
    layer0_outputs(1365) <= (inputs(81)) or (inputs(146));
    layer0_outputs(1366) <= not(inputs(229));
    layer0_outputs(1367) <= not(inputs(2));
    layer0_outputs(1368) <= not((inputs(223)) or (inputs(224)));
    layer0_outputs(1369) <= inputs(102);
    layer0_outputs(1370) <= (inputs(10)) or (inputs(251));
    layer0_outputs(1371) <= not(inputs(199)) or (inputs(242));
    layer0_outputs(1372) <= not(inputs(100));
    layer0_outputs(1373) <= '1';
    layer0_outputs(1374) <= '1';
    layer0_outputs(1375) <= not(inputs(232));
    layer0_outputs(1376) <= inputs(84);
    layer0_outputs(1377) <= (inputs(151)) or (inputs(3));
    layer0_outputs(1378) <= not(inputs(161));
    layer0_outputs(1379) <= (inputs(44)) and not (inputs(163));
    layer0_outputs(1380) <= not((inputs(220)) or (inputs(148)));
    layer0_outputs(1381) <= (inputs(32)) or (inputs(142));
    layer0_outputs(1382) <= '0';
    layer0_outputs(1383) <= not(inputs(170)) or (inputs(147));
    layer0_outputs(1384) <= (inputs(59)) and (inputs(171));
    layer0_outputs(1385) <= not(inputs(163));
    layer0_outputs(1386) <= (inputs(203)) or (inputs(172));
    layer0_outputs(1387) <= (inputs(209)) or (inputs(72));
    layer0_outputs(1388) <= inputs(182);
    layer0_outputs(1389) <= '0';
    layer0_outputs(1390) <= not((inputs(8)) or (inputs(60)));
    layer0_outputs(1391) <= (inputs(151)) and (inputs(31));
    layer0_outputs(1392) <= (inputs(250)) and not (inputs(249));
    layer0_outputs(1393) <= inputs(71);
    layer0_outputs(1394) <= not((inputs(247)) and (inputs(132)));
    layer0_outputs(1395) <= (inputs(184)) and not (inputs(128));
    layer0_outputs(1396) <= not((inputs(53)) or (inputs(117)));
    layer0_outputs(1397) <= inputs(69);
    layer0_outputs(1398) <= (inputs(78)) or (inputs(35));
    layer0_outputs(1399) <= not(inputs(9)) or (inputs(213));
    layer0_outputs(1400) <= not((inputs(149)) or (inputs(68)));
    layer0_outputs(1401) <= inputs(245);
    layer0_outputs(1402) <= (inputs(17)) xor (inputs(48));
    layer0_outputs(1403) <= inputs(149);
    layer0_outputs(1404) <= not((inputs(54)) or (inputs(222)));
    layer0_outputs(1405) <= inputs(21);
    layer0_outputs(1406) <= (inputs(155)) or (inputs(254));
    layer0_outputs(1407) <= inputs(132);
    layer0_outputs(1408) <= not(inputs(118));
    layer0_outputs(1409) <= '1';
    layer0_outputs(1410) <= not(inputs(127));
    layer0_outputs(1411) <= inputs(71);
    layer0_outputs(1412) <= (inputs(192)) or (inputs(231));
    layer0_outputs(1413) <= (inputs(58)) and not (inputs(97));
    layer0_outputs(1414) <= not(inputs(83));
    layer0_outputs(1415) <= not((inputs(163)) or (inputs(99)));
    layer0_outputs(1416) <= inputs(75);
    layer0_outputs(1417) <= (inputs(142)) and not (inputs(31));
    layer0_outputs(1418) <= not((inputs(123)) or (inputs(149)));
    layer0_outputs(1419) <= (inputs(136)) and not (inputs(176));
    layer0_outputs(1420) <= inputs(84);
    layer0_outputs(1421) <= (inputs(129)) or (inputs(234));
    layer0_outputs(1422) <= not(inputs(188));
    layer0_outputs(1423) <= not(inputs(135)) or (inputs(254));
    layer0_outputs(1424) <= (inputs(35)) and not (inputs(233));
    layer0_outputs(1425) <= not(inputs(74));
    layer0_outputs(1426) <= inputs(151);
    layer0_outputs(1427) <= not(inputs(205));
    layer0_outputs(1428) <= not((inputs(178)) or (inputs(69)));
    layer0_outputs(1429) <= inputs(130);
    layer0_outputs(1430) <= (inputs(21)) or (inputs(92));
    layer0_outputs(1431) <= not(inputs(118)) or (inputs(159));
    layer0_outputs(1432) <= inputs(141);
    layer0_outputs(1433) <= inputs(13);
    layer0_outputs(1434) <= not(inputs(156)) or (inputs(1));
    layer0_outputs(1435) <= (inputs(52)) and not (inputs(35));
    layer0_outputs(1436) <= (inputs(7)) or (inputs(255));
    layer0_outputs(1437) <= inputs(166);
    layer0_outputs(1438) <= not((inputs(77)) or (inputs(192)));
    layer0_outputs(1439) <= inputs(233);
    layer0_outputs(1440) <= not(inputs(161));
    layer0_outputs(1441) <= '1';
    layer0_outputs(1442) <= (inputs(6)) or (inputs(55));
    layer0_outputs(1443) <= (inputs(127)) and (inputs(32));
    layer0_outputs(1444) <= (inputs(44)) and not (inputs(161));
    layer0_outputs(1445) <= not(inputs(150)) or (inputs(155));
    layer0_outputs(1446) <= inputs(118);
    layer0_outputs(1447) <= (inputs(115)) or (inputs(157));
    layer0_outputs(1448) <= not((inputs(242)) or (inputs(38)));
    layer0_outputs(1449) <= not(inputs(44)) or (inputs(147));
    layer0_outputs(1450) <= (inputs(87)) and not (inputs(151));
    layer0_outputs(1451) <= inputs(231);
    layer0_outputs(1452) <= not((inputs(28)) or (inputs(233)));
    layer0_outputs(1453) <= not(inputs(160));
    layer0_outputs(1454) <= not(inputs(60));
    layer0_outputs(1455) <= not(inputs(79)) or (inputs(64));
    layer0_outputs(1456) <= not((inputs(239)) or (inputs(183)));
    layer0_outputs(1457) <= not((inputs(140)) or (inputs(165)));
    layer0_outputs(1458) <= inputs(95);
    layer0_outputs(1459) <= (inputs(125)) or (inputs(3));
    layer0_outputs(1460) <= not(inputs(166));
    layer0_outputs(1461) <= inputs(23);
    layer0_outputs(1462) <= inputs(119);
    layer0_outputs(1463) <= inputs(92);
    layer0_outputs(1464) <= (inputs(214)) and not (inputs(14));
    layer0_outputs(1465) <= not(inputs(15));
    layer0_outputs(1466) <= not(inputs(41));
    layer0_outputs(1467) <= inputs(5);
    layer0_outputs(1468) <= not((inputs(196)) or (inputs(212)));
    layer0_outputs(1469) <= not(inputs(49));
    layer0_outputs(1470) <= not(inputs(82));
    layer0_outputs(1471) <= not(inputs(66));
    layer0_outputs(1472) <= inputs(9);
    layer0_outputs(1473) <= inputs(236);
    layer0_outputs(1474) <= (inputs(179)) or (inputs(247));
    layer0_outputs(1475) <= not(inputs(135));
    layer0_outputs(1476) <= not(inputs(7)) or (inputs(54));
    layer0_outputs(1477) <= inputs(255);
    layer0_outputs(1478) <= '1';
    layer0_outputs(1479) <= (inputs(183)) and not (inputs(102));
    layer0_outputs(1480) <= '0';
    layer0_outputs(1481) <= not(inputs(230));
    layer0_outputs(1482) <= (inputs(155)) and not (inputs(95));
    layer0_outputs(1483) <= not(inputs(71));
    layer0_outputs(1484) <= (inputs(70)) or (inputs(175));
    layer0_outputs(1485) <= inputs(194);
    layer0_outputs(1486) <= not(inputs(25));
    layer0_outputs(1487) <= inputs(128);
    layer0_outputs(1488) <= (inputs(91)) or (inputs(19));
    layer0_outputs(1489) <= (inputs(50)) or (inputs(237));
    layer0_outputs(1490) <= inputs(165);
    layer0_outputs(1491) <= not(inputs(57));
    layer0_outputs(1492) <= inputs(148);
    layer0_outputs(1493) <= not((inputs(185)) and (inputs(136)));
    layer0_outputs(1494) <= '1';
    layer0_outputs(1495) <= not((inputs(51)) or (inputs(203)));
    layer0_outputs(1496) <= (inputs(189)) or (inputs(79));
    layer0_outputs(1497) <= not((inputs(106)) or (inputs(89)));
    layer0_outputs(1498) <= (inputs(175)) or (inputs(252));
    layer0_outputs(1499) <= '1';
    layer0_outputs(1500) <= not((inputs(38)) or (inputs(62)));
    layer0_outputs(1501) <= (inputs(134)) and not (inputs(214));
    layer0_outputs(1502) <= '1';
    layer0_outputs(1503) <= not(inputs(20));
    layer0_outputs(1504) <= (inputs(159)) or (inputs(71));
    layer0_outputs(1505) <= (inputs(77)) or (inputs(135));
    layer0_outputs(1506) <= not(inputs(120));
    layer0_outputs(1507) <= (inputs(154)) and not (inputs(29));
    layer0_outputs(1508) <= not((inputs(250)) or (inputs(49)));
    layer0_outputs(1509) <= (inputs(64)) or (inputs(238));
    layer0_outputs(1510) <= not(inputs(114)) or (inputs(224));
    layer0_outputs(1511) <= not((inputs(83)) or (inputs(36)));
    layer0_outputs(1512) <= inputs(158);
    layer0_outputs(1513) <= not(inputs(228));
    layer0_outputs(1514) <= not(inputs(109));
    layer0_outputs(1515) <= '1';
    layer0_outputs(1516) <= not(inputs(25));
    layer0_outputs(1517) <= (inputs(115)) and not (inputs(209));
    layer0_outputs(1518) <= not(inputs(58));
    layer0_outputs(1519) <= '1';
    layer0_outputs(1520) <= '1';
    layer0_outputs(1521) <= not(inputs(25)) or (inputs(88));
    layer0_outputs(1522) <= not(inputs(237));
    layer0_outputs(1523) <= not(inputs(204)) or (inputs(43));
    layer0_outputs(1524) <= not(inputs(13));
    layer0_outputs(1525) <= not((inputs(16)) or (inputs(157)));
    layer0_outputs(1526) <= (inputs(119)) or (inputs(67));
    layer0_outputs(1527) <= (inputs(161)) and (inputs(249));
    layer0_outputs(1528) <= (inputs(216)) or (inputs(190));
    layer0_outputs(1529) <= not(inputs(123)) or (inputs(12));
    layer0_outputs(1530) <= not(inputs(95)) or (inputs(194));
    layer0_outputs(1531) <= (inputs(151)) or (inputs(32));
    layer0_outputs(1532) <= not(inputs(91));
    layer0_outputs(1533) <= not(inputs(172)) or (inputs(52));
    layer0_outputs(1534) <= not(inputs(236)) or (inputs(184));
    layer0_outputs(1535) <= not(inputs(61)) or (inputs(106));
    layer0_outputs(1536) <= '1';
    layer0_outputs(1537) <= (inputs(204)) and (inputs(102));
    layer0_outputs(1538) <= (inputs(234)) and not (inputs(26));
    layer0_outputs(1539) <= not(inputs(64));
    layer0_outputs(1540) <= (inputs(44)) and not (inputs(117));
    layer0_outputs(1541) <= not(inputs(73)) or (inputs(55));
    layer0_outputs(1542) <= inputs(40);
    layer0_outputs(1543) <= not(inputs(167)) or (inputs(77));
    layer0_outputs(1544) <= not(inputs(154));
    layer0_outputs(1545) <= (inputs(114)) and not (inputs(139));
    layer0_outputs(1546) <= not((inputs(14)) or (inputs(45)));
    layer0_outputs(1547) <= inputs(104);
    layer0_outputs(1548) <= not(inputs(177));
    layer0_outputs(1549) <= not(inputs(231));
    layer0_outputs(1550) <= not((inputs(102)) or (inputs(68)));
    layer0_outputs(1551) <= not(inputs(138));
    layer0_outputs(1552) <= (inputs(188)) and not (inputs(85));
    layer0_outputs(1553) <= inputs(92);
    layer0_outputs(1554) <= not(inputs(215)) or (inputs(93));
    layer0_outputs(1555) <= not(inputs(192)) or (inputs(138));
    layer0_outputs(1556) <= '0';
    layer0_outputs(1557) <= inputs(58);
    layer0_outputs(1558) <= not((inputs(165)) or (inputs(197)));
    layer0_outputs(1559) <= (inputs(2)) or (inputs(14));
    layer0_outputs(1560) <= '1';
    layer0_outputs(1561) <= inputs(159);
    layer0_outputs(1562) <= not((inputs(131)) or (inputs(119)));
    layer0_outputs(1563) <= (inputs(177)) xor (inputs(77));
    layer0_outputs(1564) <= not(inputs(24)) or (inputs(67));
    layer0_outputs(1565) <= inputs(62);
    layer0_outputs(1566) <= (inputs(184)) and not (inputs(176));
    layer0_outputs(1567) <= not((inputs(173)) or (inputs(142)));
    layer0_outputs(1568) <= not((inputs(183)) and (inputs(218)));
    layer0_outputs(1569) <= not(inputs(29)) or (inputs(170));
    layer0_outputs(1570) <= '0';
    layer0_outputs(1571) <= inputs(142);
    layer0_outputs(1572) <= inputs(96);
    layer0_outputs(1573) <= (inputs(122)) and not (inputs(245));
    layer0_outputs(1574) <= not(inputs(193)) or (inputs(46));
    layer0_outputs(1575) <= '1';
    layer0_outputs(1576) <= not((inputs(112)) and (inputs(139)));
    layer0_outputs(1577) <= inputs(22);
    layer0_outputs(1578) <= not(inputs(247));
    layer0_outputs(1579) <= '1';
    layer0_outputs(1580) <= not(inputs(192));
    layer0_outputs(1581) <= (inputs(80)) and (inputs(11));
    layer0_outputs(1582) <= not(inputs(153));
    layer0_outputs(1583) <= not(inputs(72)) or (inputs(30));
    layer0_outputs(1584) <= inputs(77);
    layer0_outputs(1585) <= not(inputs(154)) or (inputs(165));
    layer0_outputs(1586) <= not(inputs(164)) or (inputs(97));
    layer0_outputs(1587) <= not(inputs(248)) or (inputs(217));
    layer0_outputs(1588) <= not((inputs(223)) or (inputs(152)));
    layer0_outputs(1589) <= inputs(8);
    layer0_outputs(1590) <= inputs(247);
    layer0_outputs(1591) <= not((inputs(149)) and (inputs(67)));
    layer0_outputs(1592) <= not((inputs(99)) and (inputs(113)));
    layer0_outputs(1593) <= not(inputs(72)) or (inputs(174));
    layer0_outputs(1594) <= (inputs(167)) or (inputs(254));
    layer0_outputs(1595) <= '0';
    layer0_outputs(1596) <= (inputs(21)) and not (inputs(173));
    layer0_outputs(1597) <= not((inputs(54)) or (inputs(102)));
    layer0_outputs(1598) <= not(inputs(233));
    layer0_outputs(1599) <= not(inputs(176)) or (inputs(197));
    layer0_outputs(1600) <= inputs(115);
    layer0_outputs(1601) <= (inputs(104)) and not (inputs(94));
    layer0_outputs(1602) <= not((inputs(206)) or (inputs(169)));
    layer0_outputs(1603) <= not((inputs(3)) or (inputs(64)));
    layer0_outputs(1604) <= inputs(90);
    layer0_outputs(1605) <= (inputs(200)) and (inputs(220));
    layer0_outputs(1606) <= inputs(182);
    layer0_outputs(1607) <= (inputs(216)) or (inputs(94));
    layer0_outputs(1608) <= not(inputs(76));
    layer0_outputs(1609) <= (inputs(181)) or (inputs(237));
    layer0_outputs(1610) <= (inputs(84)) or (inputs(47));
    layer0_outputs(1611) <= not(inputs(100)) or (inputs(111));
    layer0_outputs(1612) <= (inputs(211)) or (inputs(234));
    layer0_outputs(1613) <= inputs(93);
    layer0_outputs(1614) <= not(inputs(120)) or (inputs(141));
    layer0_outputs(1615) <= not(inputs(26)) or (inputs(166));
    layer0_outputs(1616) <= not(inputs(132)) or (inputs(35));
    layer0_outputs(1617) <= (inputs(8)) and not (inputs(194));
    layer0_outputs(1618) <= (inputs(85)) or (inputs(144));
    layer0_outputs(1619) <= (inputs(107)) and not (inputs(229));
    layer0_outputs(1620) <= not((inputs(164)) or (inputs(68)));
    layer0_outputs(1621) <= inputs(96);
    layer0_outputs(1622) <= '0';
    layer0_outputs(1623) <= (inputs(163)) xor (inputs(0));
    layer0_outputs(1624) <= (inputs(23)) or (inputs(39));
    layer0_outputs(1625) <= (inputs(9)) and not (inputs(54));
    layer0_outputs(1626) <= (inputs(77)) or (inputs(16));
    layer0_outputs(1627) <= (inputs(106)) or (inputs(167));
    layer0_outputs(1628) <= (inputs(223)) xor (inputs(228));
    layer0_outputs(1629) <= inputs(179);
    layer0_outputs(1630) <= (inputs(156)) or (inputs(69));
    layer0_outputs(1631) <= '1';
    layer0_outputs(1632) <= not((inputs(245)) or (inputs(195)));
    layer0_outputs(1633) <= inputs(94);
    layer0_outputs(1634) <= (inputs(11)) and (inputs(69));
    layer0_outputs(1635) <= inputs(74);
    layer0_outputs(1636) <= '0';
    layer0_outputs(1637) <= inputs(111);
    layer0_outputs(1638) <= not(inputs(220));
    layer0_outputs(1639) <= inputs(19);
    layer0_outputs(1640) <= (inputs(107)) or (inputs(203));
    layer0_outputs(1641) <= (inputs(57)) and not (inputs(6));
    layer0_outputs(1642) <= not(inputs(97)) or (inputs(85));
    layer0_outputs(1643) <= (inputs(167)) and not (inputs(187));
    layer0_outputs(1644) <= inputs(240);
    layer0_outputs(1645) <= inputs(150);
    layer0_outputs(1646) <= (inputs(151)) and not (inputs(140));
    layer0_outputs(1647) <= (inputs(92)) and not (inputs(1));
    layer0_outputs(1648) <= not((inputs(52)) or (inputs(24)));
    layer0_outputs(1649) <= not(inputs(19)) or (inputs(177));
    layer0_outputs(1650) <= (inputs(217)) and not (inputs(14));
    layer0_outputs(1651) <= not(inputs(199)) or (inputs(238));
    layer0_outputs(1652) <= not(inputs(14));
    layer0_outputs(1653) <= (inputs(43)) or (inputs(3));
    layer0_outputs(1654) <= not(inputs(214)) or (inputs(238));
    layer0_outputs(1655) <= (inputs(63)) and not (inputs(164));
    layer0_outputs(1656) <= not(inputs(80)) or (inputs(41));
    layer0_outputs(1657) <= inputs(130);
    layer0_outputs(1658) <= (inputs(196)) and not (inputs(239));
    layer0_outputs(1659) <= not((inputs(83)) or (inputs(129)));
    layer0_outputs(1660) <= (inputs(29)) or (inputs(186));
    layer0_outputs(1661) <= not((inputs(247)) or (inputs(221)));
    layer0_outputs(1662) <= not((inputs(94)) and (inputs(16)));
    layer0_outputs(1663) <= (inputs(37)) and not (inputs(134));
    layer0_outputs(1664) <= not(inputs(176));
    layer0_outputs(1665) <= not((inputs(140)) or (inputs(111)));
    layer0_outputs(1666) <= (inputs(245)) and (inputs(247));
    layer0_outputs(1667) <= not((inputs(102)) or (inputs(62)));
    layer0_outputs(1668) <= not(inputs(25));
    layer0_outputs(1669) <= (inputs(117)) and not (inputs(3));
    layer0_outputs(1670) <= (inputs(180)) and not (inputs(41));
    layer0_outputs(1671) <= not(inputs(222)) or (inputs(217));
    layer0_outputs(1672) <= '1';
    layer0_outputs(1673) <= (inputs(146)) and not (inputs(240));
    layer0_outputs(1674) <= not((inputs(77)) or (inputs(37)));
    layer0_outputs(1675) <= not((inputs(8)) or (inputs(178)));
    layer0_outputs(1676) <= not((inputs(110)) or (inputs(158)));
    layer0_outputs(1677) <= inputs(24);
    layer0_outputs(1678) <= not(inputs(222));
    layer0_outputs(1679) <= (inputs(177)) or (inputs(247));
    layer0_outputs(1680) <= not((inputs(172)) or (inputs(234)));
    layer0_outputs(1681) <= not(inputs(186)) or (inputs(47));
    layer0_outputs(1682) <= inputs(27);
    layer0_outputs(1683) <= not((inputs(161)) or (inputs(188)));
    layer0_outputs(1684) <= (inputs(244)) or (inputs(95));
    layer0_outputs(1685) <= not((inputs(36)) or (inputs(101)));
    layer0_outputs(1686) <= (inputs(146)) and not (inputs(46));
    layer0_outputs(1687) <= not(inputs(166));
    layer0_outputs(1688) <= inputs(45);
    layer0_outputs(1689) <= not(inputs(98));
    layer0_outputs(1690) <= not((inputs(199)) or (inputs(178)));
    layer0_outputs(1691) <= '1';
    layer0_outputs(1692) <= (inputs(72)) and not (inputs(16));
    layer0_outputs(1693) <= (inputs(207)) or (inputs(151));
    layer0_outputs(1694) <= not((inputs(221)) xor (inputs(156)));
    layer0_outputs(1695) <= (inputs(162)) or (inputs(190));
    layer0_outputs(1696) <= (inputs(196)) or (inputs(110));
    layer0_outputs(1697) <= '1';
    layer0_outputs(1698) <= not((inputs(253)) or (inputs(90)));
    layer0_outputs(1699) <= not(inputs(116));
    layer0_outputs(1700) <= not(inputs(104)) or (inputs(4));
    layer0_outputs(1701) <= not((inputs(113)) and (inputs(223)));
    layer0_outputs(1702) <= (inputs(127)) and not (inputs(13));
    layer0_outputs(1703) <= (inputs(198)) and not (inputs(22));
    layer0_outputs(1704) <= (inputs(145)) or (inputs(235));
    layer0_outputs(1705) <= inputs(92);
    layer0_outputs(1706) <= not(inputs(25));
    layer0_outputs(1707) <= not(inputs(151)) or (inputs(66));
    layer0_outputs(1708) <= not((inputs(194)) or (inputs(0)));
    layer0_outputs(1709) <= not(inputs(174)) or (inputs(99));
    layer0_outputs(1710) <= inputs(116);
    layer0_outputs(1711) <= not((inputs(138)) or (inputs(209)));
    layer0_outputs(1712) <= not(inputs(83));
    layer0_outputs(1713) <= inputs(90);
    layer0_outputs(1714) <= not(inputs(201));
    layer0_outputs(1715) <= inputs(76);
    layer0_outputs(1716) <= '0';
    layer0_outputs(1717) <= (inputs(143)) or (inputs(181));
    layer0_outputs(1718) <= not(inputs(180));
    layer0_outputs(1719) <= '0';
    layer0_outputs(1720) <= '0';
    layer0_outputs(1721) <= not(inputs(148));
    layer0_outputs(1722) <= not(inputs(238));
    layer0_outputs(1723) <= inputs(65);
    layer0_outputs(1724) <= inputs(232);
    layer0_outputs(1725) <= not((inputs(161)) or (inputs(218)));
    layer0_outputs(1726) <= (inputs(188)) and not (inputs(77));
    layer0_outputs(1727) <= (inputs(239)) or (inputs(181));
    layer0_outputs(1728) <= not((inputs(200)) and (inputs(222)));
    layer0_outputs(1729) <= not((inputs(40)) or (inputs(95)));
    layer0_outputs(1730) <= not((inputs(162)) or (inputs(161)));
    layer0_outputs(1731) <= inputs(215);
    layer0_outputs(1732) <= inputs(103);
    layer0_outputs(1733) <= not(inputs(100));
    layer0_outputs(1734) <= (inputs(218)) or (inputs(80));
    layer0_outputs(1735) <= not(inputs(210));
    layer0_outputs(1736) <= not((inputs(33)) or (inputs(178)));
    layer0_outputs(1737) <= (inputs(152)) and not (inputs(118));
    layer0_outputs(1738) <= inputs(227);
    layer0_outputs(1739) <= not((inputs(155)) or (inputs(172)));
    layer0_outputs(1740) <= (inputs(101)) and not (inputs(249));
    layer0_outputs(1741) <= inputs(102);
    layer0_outputs(1742) <= not((inputs(194)) or (inputs(235)));
    layer0_outputs(1743) <= not((inputs(2)) or (inputs(210)));
    layer0_outputs(1744) <= inputs(226);
    layer0_outputs(1745) <= '0';
    layer0_outputs(1746) <= (inputs(26)) and not (inputs(113));
    layer0_outputs(1747) <= inputs(56);
    layer0_outputs(1748) <= inputs(109);
    layer0_outputs(1749) <= not(inputs(24));
    layer0_outputs(1750) <= inputs(128);
    layer0_outputs(1751) <= not(inputs(254));
    layer0_outputs(1752) <= (inputs(5)) and not (inputs(177));
    layer0_outputs(1753) <= '0';
    layer0_outputs(1754) <= not((inputs(240)) or (inputs(22)));
    layer0_outputs(1755) <= not(inputs(103));
    layer0_outputs(1756) <= '1';
    layer0_outputs(1757) <= (inputs(96)) or (inputs(77));
    layer0_outputs(1758) <= inputs(125);
    layer0_outputs(1759) <= not(inputs(110));
    layer0_outputs(1760) <= inputs(105);
    layer0_outputs(1761) <= inputs(226);
    layer0_outputs(1762) <= not(inputs(100)) or (inputs(225));
    layer0_outputs(1763) <= inputs(151);
    layer0_outputs(1764) <= (inputs(106)) and not (inputs(56));
    layer0_outputs(1765) <= not((inputs(226)) or (inputs(244)));
    layer0_outputs(1766) <= not((inputs(96)) or (inputs(124)));
    layer0_outputs(1767) <= not((inputs(239)) and (inputs(238)));
    layer0_outputs(1768) <= (inputs(110)) or (inputs(171));
    layer0_outputs(1769) <= inputs(185);
    layer0_outputs(1770) <= not((inputs(25)) or (inputs(75)));
    layer0_outputs(1771) <= inputs(69);
    layer0_outputs(1772) <= (inputs(129)) and (inputs(140));
    layer0_outputs(1773) <= (inputs(48)) or (inputs(95));
    layer0_outputs(1774) <= not(inputs(138));
    layer0_outputs(1775) <= not(inputs(95));
    layer0_outputs(1776) <= not(inputs(52));
    layer0_outputs(1777) <= (inputs(255)) or (inputs(167));
    layer0_outputs(1778) <= (inputs(99)) or (inputs(69));
    layer0_outputs(1779) <= inputs(98);
    layer0_outputs(1780) <= (inputs(49)) and not (inputs(125));
    layer0_outputs(1781) <= not(inputs(195));
    layer0_outputs(1782) <= not(inputs(162));
    layer0_outputs(1783) <= inputs(230);
    layer0_outputs(1784) <= not((inputs(70)) or (inputs(65)));
    layer0_outputs(1785) <= (inputs(176)) or (inputs(178));
    layer0_outputs(1786) <= not((inputs(128)) or (inputs(180)));
    layer0_outputs(1787) <= not(inputs(50));
    layer0_outputs(1788) <= not(inputs(145));
    layer0_outputs(1789) <= inputs(218);
    layer0_outputs(1790) <= not((inputs(107)) and (inputs(131)));
    layer0_outputs(1791) <= (inputs(112)) or (inputs(202));
    layer0_outputs(1792) <= not(inputs(209));
    layer0_outputs(1793) <= (inputs(154)) and not (inputs(10));
    layer0_outputs(1794) <= not(inputs(145)) or (inputs(240));
    layer0_outputs(1795) <= not(inputs(117));
    layer0_outputs(1796) <= (inputs(78)) or (inputs(61));
    layer0_outputs(1797) <= not(inputs(28));
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= (inputs(34)) or (inputs(90));
    layer0_outputs(1800) <= (inputs(160)) or (inputs(131));
    layer0_outputs(1801) <= not(inputs(140));
    layer0_outputs(1802) <= (inputs(245)) or (inputs(214));
    layer0_outputs(1803) <= not((inputs(78)) and (inputs(77)));
    layer0_outputs(1804) <= (inputs(96)) or (inputs(246));
    layer0_outputs(1805) <= (inputs(241)) or (inputs(7));
    layer0_outputs(1806) <= '1';
    layer0_outputs(1807) <= (inputs(164)) and not (inputs(43));
    layer0_outputs(1808) <= not((inputs(93)) or (inputs(169)));
    layer0_outputs(1809) <= not(inputs(53));
    layer0_outputs(1810) <= inputs(237);
    layer0_outputs(1811) <= inputs(14);
    layer0_outputs(1812) <= inputs(219);
    layer0_outputs(1813) <= not(inputs(192));
    layer0_outputs(1814) <= not(inputs(101));
    layer0_outputs(1815) <= (inputs(107)) or (inputs(108));
    layer0_outputs(1816) <= inputs(197);
    layer0_outputs(1817) <= inputs(120);
    layer0_outputs(1818) <= not((inputs(194)) or (inputs(179)));
    layer0_outputs(1819) <= not(inputs(226));
    layer0_outputs(1820) <= '1';
    layer0_outputs(1821) <= (inputs(106)) and not (inputs(219));
    layer0_outputs(1822) <= (inputs(11)) and not (inputs(165));
    layer0_outputs(1823) <= (inputs(230)) or (inputs(177));
    layer0_outputs(1824) <= inputs(1);
    layer0_outputs(1825) <= (inputs(70)) and not (inputs(42));
    layer0_outputs(1826) <= not(inputs(112));
    layer0_outputs(1827) <= inputs(128);
    layer0_outputs(1828) <= not((inputs(227)) or (inputs(229)));
    layer0_outputs(1829) <= not((inputs(20)) or (inputs(153)));
    layer0_outputs(1830) <= not((inputs(233)) or (inputs(157)));
    layer0_outputs(1831) <= not((inputs(58)) and (inputs(5)));
    layer0_outputs(1832) <= inputs(217);
    layer0_outputs(1833) <= not(inputs(130)) or (inputs(189));
    layer0_outputs(1834) <= inputs(24);
    layer0_outputs(1835) <= not((inputs(32)) or (inputs(224)));
    layer0_outputs(1836) <= not(inputs(26)) or (inputs(132));
    layer0_outputs(1837) <= not((inputs(206)) xor (inputs(3)));
    layer0_outputs(1838) <= '1';
    layer0_outputs(1839) <= (inputs(64)) and not (inputs(194));
    layer0_outputs(1840) <= inputs(147);
    layer0_outputs(1841) <= not((inputs(252)) or (inputs(169)));
    layer0_outputs(1842) <= '1';
    layer0_outputs(1843) <= inputs(0);
    layer0_outputs(1844) <= not(inputs(215));
    layer0_outputs(1845) <= (inputs(246)) or (inputs(64));
    layer0_outputs(1846) <= not((inputs(51)) or (inputs(36)));
    layer0_outputs(1847) <= not((inputs(218)) xor (inputs(236)));
    layer0_outputs(1848) <= not(inputs(136));
    layer0_outputs(1849) <= not((inputs(240)) or (inputs(127)));
    layer0_outputs(1850) <= not((inputs(174)) xor (inputs(127)));
    layer0_outputs(1851) <= not(inputs(214)) or (inputs(32));
    layer0_outputs(1852) <= not(inputs(219));
    layer0_outputs(1853) <= not(inputs(22));
    layer0_outputs(1854) <= not(inputs(180));
    layer0_outputs(1855) <= '1';
    layer0_outputs(1856) <= (inputs(104)) and not (inputs(114));
    layer0_outputs(1857) <= (inputs(106)) and not (inputs(205));
    layer0_outputs(1858) <= not((inputs(88)) xor (inputs(31)));
    layer0_outputs(1859) <= not(inputs(213));
    layer0_outputs(1860) <= not((inputs(148)) or (inputs(68)));
    layer0_outputs(1861) <= not(inputs(75));
    layer0_outputs(1862) <= (inputs(133)) or (inputs(28));
    layer0_outputs(1863) <= not(inputs(121));
    layer0_outputs(1864) <= not(inputs(40));
    layer0_outputs(1865) <= not(inputs(40));
    layer0_outputs(1866) <= (inputs(68)) or (inputs(35));
    layer0_outputs(1867) <= not((inputs(116)) or (inputs(162)));
    layer0_outputs(1868) <= not((inputs(228)) or (inputs(175)));
    layer0_outputs(1869) <= not(inputs(34));
    layer0_outputs(1870) <= inputs(23);
    layer0_outputs(1871) <= (inputs(208)) or (inputs(143));
    layer0_outputs(1872) <= '1';
    layer0_outputs(1873) <= not(inputs(55));
    layer0_outputs(1874) <= '0';
    layer0_outputs(1875) <= not(inputs(48));
    layer0_outputs(1876) <= '1';
    layer0_outputs(1877) <= inputs(227);
    layer0_outputs(1878) <= inputs(233);
    layer0_outputs(1879) <= not(inputs(19));
    layer0_outputs(1880) <= (inputs(99)) or (inputs(165));
    layer0_outputs(1881) <= (inputs(188)) or (inputs(222));
    layer0_outputs(1882) <= not(inputs(103));
    layer0_outputs(1883) <= not(inputs(180)) or (inputs(45));
    layer0_outputs(1884) <= not((inputs(156)) or (inputs(20)));
    layer0_outputs(1885) <= not(inputs(181));
    layer0_outputs(1886) <= (inputs(215)) or (inputs(105));
    layer0_outputs(1887) <= not(inputs(109));
    layer0_outputs(1888) <= inputs(168);
    layer0_outputs(1889) <= inputs(101);
    layer0_outputs(1890) <= (inputs(180)) and not (inputs(15));
    layer0_outputs(1891) <= not(inputs(179));
    layer0_outputs(1892) <= (inputs(126)) and not (inputs(63));
    layer0_outputs(1893) <= (inputs(218)) or (inputs(77));
    layer0_outputs(1894) <= not(inputs(24));
    layer0_outputs(1895) <= not(inputs(75)) or (inputs(146));
    layer0_outputs(1896) <= (inputs(182)) and not (inputs(157));
    layer0_outputs(1897) <= not((inputs(233)) or (inputs(242)));
    layer0_outputs(1898) <= inputs(202);
    layer0_outputs(1899) <= not(inputs(157));
    layer0_outputs(1900) <= '0';
    layer0_outputs(1901) <= not(inputs(229));
    layer0_outputs(1902) <= not(inputs(91));
    layer0_outputs(1903) <= not(inputs(178)) or (inputs(190));
    layer0_outputs(1904) <= not(inputs(106));
    layer0_outputs(1905) <= inputs(79);
    layer0_outputs(1906) <= (inputs(88)) and not (inputs(162));
    layer0_outputs(1907) <= not(inputs(72)) or (inputs(37));
    layer0_outputs(1908) <= (inputs(248)) or (inputs(246));
    layer0_outputs(1909) <= not(inputs(116));
    layer0_outputs(1910) <= '0';
    layer0_outputs(1911) <= inputs(5);
    layer0_outputs(1912) <= not(inputs(142)) or (inputs(239));
    layer0_outputs(1913) <= not((inputs(13)) or (inputs(135)));
    layer0_outputs(1914) <= inputs(180);
    layer0_outputs(1915) <= not(inputs(136)) or (inputs(68));
    layer0_outputs(1916) <= '0';
    layer0_outputs(1917) <= '0';
    layer0_outputs(1918) <= '1';
    layer0_outputs(1919) <= (inputs(235)) and not (inputs(162));
    layer0_outputs(1920) <= inputs(33);
    layer0_outputs(1921) <= inputs(183);
    layer0_outputs(1922) <= (inputs(130)) xor (inputs(180));
    layer0_outputs(1923) <= not(inputs(152)) or (inputs(159));
    layer0_outputs(1924) <= inputs(37);
    layer0_outputs(1925) <= not(inputs(127));
    layer0_outputs(1926) <= (inputs(21)) or (inputs(170));
    layer0_outputs(1927) <= not(inputs(106));
    layer0_outputs(1928) <= inputs(221);
    layer0_outputs(1929) <= not((inputs(206)) or (inputs(171)));
    layer0_outputs(1930) <= (inputs(225)) and not (inputs(216));
    layer0_outputs(1931) <= not(inputs(193)) or (inputs(239));
    layer0_outputs(1932) <= not((inputs(159)) or (inputs(124)));
    layer0_outputs(1933) <= not(inputs(204));
    layer0_outputs(1934) <= (inputs(243)) and (inputs(15));
    layer0_outputs(1935) <= (inputs(134)) and not (inputs(113));
    layer0_outputs(1936) <= not(inputs(173)) or (inputs(63));
    layer0_outputs(1937) <= not((inputs(206)) or (inputs(237)));
    layer0_outputs(1938) <= not(inputs(70)) or (inputs(31));
    layer0_outputs(1939) <= not(inputs(1));
    layer0_outputs(1940) <= inputs(110);
    layer0_outputs(1941) <= inputs(119);
    layer0_outputs(1942) <= (inputs(210)) and not (inputs(114));
    layer0_outputs(1943) <= (inputs(231)) or (inputs(174));
    layer0_outputs(1944) <= not(inputs(56));
    layer0_outputs(1945) <= (inputs(16)) and not (inputs(0));
    layer0_outputs(1946) <= not(inputs(67)) or (inputs(111));
    layer0_outputs(1947) <= (inputs(243)) and not (inputs(143));
    layer0_outputs(1948) <= not(inputs(213));
    layer0_outputs(1949) <= not(inputs(207));
    layer0_outputs(1950) <= not(inputs(41)) or (inputs(131));
    layer0_outputs(1951) <= (inputs(118)) or (inputs(159));
    layer0_outputs(1952) <= inputs(83);
    layer0_outputs(1953) <= (inputs(197)) or (inputs(17));
    layer0_outputs(1954) <= not((inputs(80)) and (inputs(133)));
    layer0_outputs(1955) <= inputs(104);
    layer0_outputs(1956) <= inputs(62);
    layer0_outputs(1957) <= not(inputs(212));
    layer0_outputs(1958) <= not((inputs(34)) xor (inputs(76)));
    layer0_outputs(1959) <= not((inputs(110)) or (inputs(198)));
    layer0_outputs(1960) <= not(inputs(144));
    layer0_outputs(1961) <= (inputs(225)) and not (inputs(45));
    layer0_outputs(1962) <= not(inputs(21)) or (inputs(190));
    layer0_outputs(1963) <= not((inputs(171)) and (inputs(221)));
    layer0_outputs(1964) <= not((inputs(80)) or (inputs(179)));
    layer0_outputs(1965) <= inputs(116);
    layer0_outputs(1966) <= not(inputs(231));
    layer0_outputs(1967) <= '1';
    layer0_outputs(1968) <= not((inputs(39)) or (inputs(245)));
    layer0_outputs(1969) <= '1';
    layer0_outputs(1970) <= not(inputs(87)) or (inputs(129));
    layer0_outputs(1971) <= (inputs(75)) and not (inputs(208));
    layer0_outputs(1972) <= inputs(229);
    layer0_outputs(1973) <= not(inputs(75));
    layer0_outputs(1974) <= not(inputs(100));
    layer0_outputs(1975) <= '1';
    layer0_outputs(1976) <= inputs(18);
    layer0_outputs(1977) <= not(inputs(107)) or (inputs(245));
    layer0_outputs(1978) <= not(inputs(125));
    layer0_outputs(1979) <= not((inputs(166)) and (inputs(137)));
    layer0_outputs(1980) <= (inputs(12)) or (inputs(21));
    layer0_outputs(1981) <= not(inputs(96)) or (inputs(207));
    layer0_outputs(1982) <= not(inputs(195)) or (inputs(112));
    layer0_outputs(1983) <= not(inputs(101));
    layer0_outputs(1984) <= '0';
    layer0_outputs(1985) <= not((inputs(22)) or (inputs(216)));
    layer0_outputs(1986) <= inputs(87);
    layer0_outputs(1987) <= '1';
    layer0_outputs(1988) <= not(inputs(125));
    layer0_outputs(1989) <= not(inputs(239));
    layer0_outputs(1990) <= inputs(211);
    layer0_outputs(1991) <= not(inputs(166));
    layer0_outputs(1992) <= not(inputs(185)) or (inputs(170));
    layer0_outputs(1993) <= (inputs(7)) and not (inputs(251));
    layer0_outputs(1994) <= inputs(134);
    layer0_outputs(1995) <= not(inputs(203)) or (inputs(37));
    layer0_outputs(1996) <= inputs(210);
    layer0_outputs(1997) <= (inputs(166)) or (inputs(230));
    layer0_outputs(1998) <= not(inputs(98)) or (inputs(243));
    layer0_outputs(1999) <= inputs(69);
    layer0_outputs(2000) <= not(inputs(179));
    layer0_outputs(2001) <= not((inputs(52)) and (inputs(42)));
    layer0_outputs(2002) <= not((inputs(22)) and (inputs(67)));
    layer0_outputs(2003) <= not(inputs(230));
    layer0_outputs(2004) <= (inputs(247)) and not (inputs(16));
    layer0_outputs(2005) <= not((inputs(249)) and (inputs(243)));
    layer0_outputs(2006) <= inputs(240);
    layer0_outputs(2007) <= inputs(36);
    layer0_outputs(2008) <= inputs(135);
    layer0_outputs(2009) <= not(inputs(204));
    layer0_outputs(2010) <= not(inputs(85));
    layer0_outputs(2011) <= (inputs(130)) or (inputs(161));
    layer0_outputs(2012) <= inputs(73);
    layer0_outputs(2013) <= inputs(167);
    layer0_outputs(2014) <= not((inputs(74)) or (inputs(171)));
    layer0_outputs(2015) <= '1';
    layer0_outputs(2016) <= inputs(220);
    layer0_outputs(2017) <= not(inputs(153)) or (inputs(241));
    layer0_outputs(2018) <= not(inputs(201));
    layer0_outputs(2019) <= (inputs(129)) or (inputs(6));
    layer0_outputs(2020) <= not(inputs(167)) or (inputs(85));
    layer0_outputs(2021) <= (inputs(8)) or (inputs(208));
    layer0_outputs(2022) <= (inputs(66)) or (inputs(198));
    layer0_outputs(2023) <= (inputs(128)) and not (inputs(152));
    layer0_outputs(2024) <= not((inputs(148)) or (inputs(172)));
    layer0_outputs(2025) <= (inputs(231)) and not (inputs(73));
    layer0_outputs(2026) <= not((inputs(20)) and (inputs(207)));
    layer0_outputs(2027) <= (inputs(190)) and not (inputs(239));
    layer0_outputs(2028) <= (inputs(11)) and not (inputs(190));
    layer0_outputs(2029) <= inputs(224);
    layer0_outputs(2030) <= (inputs(201)) and (inputs(196));
    layer0_outputs(2031) <= (inputs(46)) or (inputs(181));
    layer0_outputs(2032) <= '1';
    layer0_outputs(2033) <= (inputs(81)) and (inputs(175));
    layer0_outputs(2034) <= (inputs(253)) or (inputs(6));
    layer0_outputs(2035) <= not(inputs(165));
    layer0_outputs(2036) <= '0';
    layer0_outputs(2037) <= (inputs(252)) xor (inputs(243));
    layer0_outputs(2038) <= not((inputs(195)) xor (inputs(51)));
    layer0_outputs(2039) <= not(inputs(91)) or (inputs(178));
    layer0_outputs(2040) <= '1';
    layer0_outputs(2041) <= not((inputs(130)) xor (inputs(19)));
    layer0_outputs(2042) <= inputs(8);
    layer0_outputs(2043) <= not(inputs(118));
    layer0_outputs(2044) <= inputs(244);
    layer0_outputs(2045) <= (inputs(8)) and not (inputs(224));
    layer0_outputs(2046) <= inputs(64);
    layer0_outputs(2047) <= not(inputs(143));
    layer0_outputs(2048) <= inputs(134);
    layer0_outputs(2049) <= inputs(127);
    layer0_outputs(2050) <= not(inputs(150)) or (inputs(236));
    layer0_outputs(2051) <= (inputs(103)) and (inputs(17));
    layer0_outputs(2052) <= not(inputs(220)) or (inputs(113));
    layer0_outputs(2053) <= not(inputs(141));
    layer0_outputs(2054) <= '0';
    layer0_outputs(2055) <= not(inputs(133));
    layer0_outputs(2056) <= '0';
    layer0_outputs(2057) <= inputs(83);
    layer0_outputs(2058) <= not(inputs(61));
    layer0_outputs(2059) <= not(inputs(94));
    layer0_outputs(2060) <= not(inputs(124)) or (inputs(227));
    layer0_outputs(2061) <= not(inputs(46)) or (inputs(176));
    layer0_outputs(2062) <= (inputs(216)) or (inputs(112));
    layer0_outputs(2063) <= not(inputs(119)) or (inputs(2));
    layer0_outputs(2064) <= (inputs(100)) and not (inputs(141));
    layer0_outputs(2065) <= (inputs(205)) or (inputs(85));
    layer0_outputs(2066) <= not(inputs(106)) or (inputs(84));
    layer0_outputs(2067) <= (inputs(102)) or (inputs(88));
    layer0_outputs(2068) <= not((inputs(203)) or (inputs(39)));
    layer0_outputs(2069) <= not((inputs(104)) and (inputs(238)));
    layer0_outputs(2070) <= not((inputs(228)) or (inputs(189)));
    layer0_outputs(2071) <= inputs(8);
    layer0_outputs(2072) <= inputs(135);
    layer0_outputs(2073) <= not(inputs(135)) or (inputs(60));
    layer0_outputs(2074) <= (inputs(202)) or (inputs(4));
    layer0_outputs(2075) <= inputs(21);
    layer0_outputs(2076) <= not(inputs(14));
    layer0_outputs(2077) <= (inputs(121)) and not (inputs(177));
    layer0_outputs(2078) <= not((inputs(70)) or (inputs(86)));
    layer0_outputs(2079) <= inputs(97);
    layer0_outputs(2080) <= inputs(102);
    layer0_outputs(2081) <= (inputs(234)) or (inputs(210));
    layer0_outputs(2082) <= (inputs(205)) or (inputs(84));
    layer0_outputs(2083) <= '0';
    layer0_outputs(2084) <= not(inputs(89)) or (inputs(129));
    layer0_outputs(2085) <= not(inputs(177));
    layer0_outputs(2086) <= not(inputs(118));
    layer0_outputs(2087) <= (inputs(210)) or (inputs(89));
    layer0_outputs(2088) <= not(inputs(108));
    layer0_outputs(2089) <= (inputs(13)) xor (inputs(50));
    layer0_outputs(2090) <= (inputs(89)) xor (inputs(194));
    layer0_outputs(2091) <= not(inputs(58));
    layer0_outputs(2092) <= not(inputs(164));
    layer0_outputs(2093) <= (inputs(198)) or (inputs(254));
    layer0_outputs(2094) <= '0';
    layer0_outputs(2095) <= inputs(253);
    layer0_outputs(2096) <= not(inputs(199)) or (inputs(103));
    layer0_outputs(2097) <= '0';
    layer0_outputs(2098) <= not((inputs(8)) and (inputs(118)));
    layer0_outputs(2099) <= (inputs(200)) xor (inputs(214));
    layer0_outputs(2100) <= not(inputs(179)) or (inputs(3));
    layer0_outputs(2101) <= inputs(180);
    layer0_outputs(2102) <= (inputs(205)) and not (inputs(10));
    layer0_outputs(2103) <= (inputs(105)) and not (inputs(146));
    layer0_outputs(2104) <= not(inputs(136));
    layer0_outputs(2105) <= not((inputs(111)) or (inputs(121)));
    layer0_outputs(2106) <= not(inputs(168));
    layer0_outputs(2107) <= '1';
    layer0_outputs(2108) <= inputs(176);
    layer0_outputs(2109) <= (inputs(9)) or (inputs(254));
    layer0_outputs(2110) <= not((inputs(189)) or (inputs(70)));
    layer0_outputs(2111) <= not((inputs(31)) or (inputs(166)));
    layer0_outputs(2112) <= inputs(126);
    layer0_outputs(2113) <= not(inputs(57));
    layer0_outputs(2114) <= (inputs(38)) and not (inputs(205));
    layer0_outputs(2115) <= (inputs(15)) or (inputs(140));
    layer0_outputs(2116) <= (inputs(207)) or (inputs(150));
    layer0_outputs(2117) <= '0';
    layer0_outputs(2118) <= inputs(33);
    layer0_outputs(2119) <= not(inputs(233));
    layer0_outputs(2120) <= (inputs(150)) or (inputs(198));
    layer0_outputs(2121) <= not((inputs(70)) or (inputs(67)));
    layer0_outputs(2122) <= (inputs(206)) or (inputs(212));
    layer0_outputs(2123) <= not(inputs(120));
    layer0_outputs(2124) <= not(inputs(246));
    layer0_outputs(2125) <= inputs(100);
    layer0_outputs(2126) <= (inputs(106)) and not (inputs(176));
    layer0_outputs(2127) <= '0';
    layer0_outputs(2128) <= not(inputs(30));
    layer0_outputs(2129) <= (inputs(226)) or (inputs(59));
    layer0_outputs(2130) <= (inputs(181)) and not (inputs(211));
    layer0_outputs(2131) <= not((inputs(46)) or (inputs(55)));
    layer0_outputs(2132) <= (inputs(203)) or (inputs(223));
    layer0_outputs(2133) <= (inputs(166)) or (inputs(219));
    layer0_outputs(2134) <= inputs(159);
    layer0_outputs(2135) <= '1';
    layer0_outputs(2136) <= not(inputs(46));
    layer0_outputs(2137) <= not((inputs(205)) or (inputs(20)));
    layer0_outputs(2138) <= inputs(116);
    layer0_outputs(2139) <= not((inputs(0)) xor (inputs(10)));
    layer0_outputs(2140) <= not((inputs(204)) or (inputs(165)));
    layer0_outputs(2141) <= not((inputs(193)) xor (inputs(240)));
    layer0_outputs(2142) <= (inputs(55)) and not (inputs(121));
    layer0_outputs(2143) <= not((inputs(248)) or (inputs(246)));
    layer0_outputs(2144) <= (inputs(47)) and not (inputs(124));
    layer0_outputs(2145) <= not(inputs(86)) or (inputs(1));
    layer0_outputs(2146) <= inputs(115);
    layer0_outputs(2147) <= '0';
    layer0_outputs(2148) <= '1';
    layer0_outputs(2149) <= '1';
    layer0_outputs(2150) <= not((inputs(176)) or (inputs(84)));
    layer0_outputs(2151) <= not(inputs(247));
    layer0_outputs(2152) <= '0';
    layer0_outputs(2153) <= not((inputs(238)) or (inputs(76)));
    layer0_outputs(2154) <= not(inputs(150));
    layer0_outputs(2155) <= (inputs(235)) and not (inputs(86));
    layer0_outputs(2156) <= (inputs(117)) or (inputs(104));
    layer0_outputs(2157) <= not((inputs(201)) and (inputs(29)));
    layer0_outputs(2158) <= inputs(124);
    layer0_outputs(2159) <= (inputs(28)) or (inputs(196));
    layer0_outputs(2160) <= inputs(75);
    layer0_outputs(2161) <= (inputs(86)) and not (inputs(253));
    layer0_outputs(2162) <= not(inputs(30));
    layer0_outputs(2163) <= (inputs(113)) or (inputs(87));
    layer0_outputs(2164) <= not((inputs(38)) and (inputs(0)));
    layer0_outputs(2165) <= (inputs(191)) and not (inputs(42));
    layer0_outputs(2166) <= not(inputs(191));
    layer0_outputs(2167) <= (inputs(251)) and (inputs(225));
    layer0_outputs(2168) <= '1';
    layer0_outputs(2169) <= not(inputs(37));
    layer0_outputs(2170) <= not(inputs(106)) or (inputs(196));
    layer0_outputs(2171) <= (inputs(136)) and (inputs(101));
    layer0_outputs(2172) <= (inputs(36)) and not (inputs(137));
    layer0_outputs(2173) <= (inputs(3)) or (inputs(78));
    layer0_outputs(2174) <= inputs(32);
    layer0_outputs(2175) <= (inputs(186)) and (inputs(191));
    layer0_outputs(2176) <= not((inputs(27)) or (inputs(232)));
    layer0_outputs(2177) <= not(inputs(67));
    layer0_outputs(2178) <= not((inputs(232)) xor (inputs(200)));
    layer0_outputs(2179) <= inputs(149);
    layer0_outputs(2180) <= not(inputs(171)) or (inputs(67));
    layer0_outputs(2181) <= not(inputs(83));
    layer0_outputs(2182) <= inputs(114);
    layer0_outputs(2183) <= not(inputs(130));
    layer0_outputs(2184) <= (inputs(244)) or (inputs(130));
    layer0_outputs(2185) <= not((inputs(56)) or (inputs(161)));
    layer0_outputs(2186) <= not(inputs(164));
    layer0_outputs(2187) <= not(inputs(72));
    layer0_outputs(2188) <= inputs(74);
    layer0_outputs(2189) <= inputs(186);
    layer0_outputs(2190) <= not(inputs(137));
    layer0_outputs(2191) <= not(inputs(58));
    layer0_outputs(2192) <= not((inputs(160)) or (inputs(143)));
    layer0_outputs(2193) <= not(inputs(103));
    layer0_outputs(2194) <= (inputs(69)) or (inputs(209));
    layer0_outputs(2195) <= '0';
    layer0_outputs(2196) <= '1';
    layer0_outputs(2197) <= inputs(139);
    layer0_outputs(2198) <= inputs(127);
    layer0_outputs(2199) <= inputs(75);
    layer0_outputs(2200) <= not((inputs(226)) or (inputs(171)));
    layer0_outputs(2201) <= (inputs(117)) or (inputs(67));
    layer0_outputs(2202) <= not((inputs(87)) and (inputs(103)));
    layer0_outputs(2203) <= not(inputs(69)) or (inputs(105));
    layer0_outputs(2204) <= not(inputs(46)) or (inputs(209));
    layer0_outputs(2205) <= '0';
    layer0_outputs(2206) <= (inputs(37)) or (inputs(201));
    layer0_outputs(2207) <= inputs(172);
    layer0_outputs(2208) <= (inputs(183)) xor (inputs(213));
    layer0_outputs(2209) <= not(inputs(118));
    layer0_outputs(2210) <= inputs(19);
    layer0_outputs(2211) <= not(inputs(24));
    layer0_outputs(2212) <= (inputs(0)) and not (inputs(51));
    layer0_outputs(2213) <= not(inputs(231));
    layer0_outputs(2214) <= inputs(67);
    layer0_outputs(2215) <= (inputs(131)) and not (inputs(210));
    layer0_outputs(2216) <= not(inputs(22));
    layer0_outputs(2217) <= not((inputs(236)) or (inputs(208)));
    layer0_outputs(2218) <= not(inputs(228));
    layer0_outputs(2219) <= not(inputs(150));
    layer0_outputs(2220) <= not(inputs(195));
    layer0_outputs(2221) <= not(inputs(233));
    layer0_outputs(2222) <= not(inputs(203));
    layer0_outputs(2223) <= not(inputs(165)) or (inputs(239));
    layer0_outputs(2224) <= inputs(19);
    layer0_outputs(2225) <= inputs(144);
    layer0_outputs(2226) <= '0';
    layer0_outputs(2227) <= inputs(19);
    layer0_outputs(2228) <= not((inputs(89)) and (inputs(68)));
    layer0_outputs(2229) <= inputs(177);
    layer0_outputs(2230) <= inputs(98);
    layer0_outputs(2231) <= '1';
    layer0_outputs(2232) <= inputs(23);
    layer0_outputs(2233) <= '0';
    layer0_outputs(2234) <= not(inputs(248));
    layer0_outputs(2235) <= inputs(197);
    layer0_outputs(2236) <= (inputs(142)) and not (inputs(255));
    layer0_outputs(2237) <= not((inputs(207)) or (inputs(178)));
    layer0_outputs(2238) <= inputs(224);
    layer0_outputs(2239) <= not((inputs(33)) or (inputs(5)));
    layer0_outputs(2240) <= (inputs(170)) and not (inputs(127));
    layer0_outputs(2241) <= not(inputs(209));
    layer0_outputs(2242) <= not((inputs(175)) or (inputs(211)));
    layer0_outputs(2243) <= (inputs(174)) and (inputs(13));
    layer0_outputs(2244) <= (inputs(50)) or (inputs(154));
    layer0_outputs(2245) <= not((inputs(45)) or (inputs(52)));
    layer0_outputs(2246) <= not((inputs(207)) or (inputs(210)));
    layer0_outputs(2247) <= not(inputs(231)) or (inputs(115));
    layer0_outputs(2248) <= not(inputs(120)) or (inputs(143));
    layer0_outputs(2249) <= (inputs(26)) and not (inputs(243));
    layer0_outputs(2250) <= '0';
    layer0_outputs(2251) <= not(inputs(121));
    layer0_outputs(2252) <= '1';
    layer0_outputs(2253) <= (inputs(132)) and (inputs(101));
    layer0_outputs(2254) <= (inputs(96)) or (inputs(245));
    layer0_outputs(2255) <= inputs(89);
    layer0_outputs(2256) <= not(inputs(212));
    layer0_outputs(2257) <= (inputs(55)) and not (inputs(155));
    layer0_outputs(2258) <= (inputs(32)) or (inputs(95));
    layer0_outputs(2259) <= not(inputs(188)) or (inputs(3));
    layer0_outputs(2260) <= (inputs(177)) and not (inputs(205));
    layer0_outputs(2261) <= inputs(102);
    layer0_outputs(2262) <= inputs(209);
    layer0_outputs(2263) <= '1';
    layer0_outputs(2264) <= not((inputs(9)) or (inputs(246)));
    layer0_outputs(2265) <= not(inputs(112));
    layer0_outputs(2266) <= not((inputs(164)) or (inputs(255)));
    layer0_outputs(2267) <= not(inputs(59)) or (inputs(168));
    layer0_outputs(2268) <= not(inputs(246)) or (inputs(89));
    layer0_outputs(2269) <= (inputs(161)) or (inputs(164));
    layer0_outputs(2270) <= inputs(43);
    layer0_outputs(2271) <= not(inputs(10));
    layer0_outputs(2272) <= not(inputs(25));
    layer0_outputs(2273) <= '0';
    layer0_outputs(2274) <= not(inputs(109)) or (inputs(67));
    layer0_outputs(2275) <= inputs(191);
    layer0_outputs(2276) <= inputs(98);
    layer0_outputs(2277) <= not((inputs(159)) or (inputs(233)));
    layer0_outputs(2278) <= not(inputs(140));
    layer0_outputs(2279) <= not(inputs(121));
    layer0_outputs(2280) <= (inputs(179)) or (inputs(167));
    layer0_outputs(2281) <= not((inputs(107)) xor (inputs(182)));
    layer0_outputs(2282) <= not(inputs(179));
    layer0_outputs(2283) <= not(inputs(72));
    layer0_outputs(2284) <= inputs(160);
    layer0_outputs(2285) <= not(inputs(226));
    layer0_outputs(2286) <= not((inputs(142)) or (inputs(173)));
    layer0_outputs(2287) <= not(inputs(141));
    layer0_outputs(2288) <= inputs(76);
    layer0_outputs(2289) <= inputs(105);
    layer0_outputs(2290) <= (inputs(78)) xor (inputs(89));
    layer0_outputs(2291) <= (inputs(22)) and not (inputs(101));
    layer0_outputs(2292) <= (inputs(123)) and (inputs(41));
    layer0_outputs(2293) <= (inputs(199)) and (inputs(46));
    layer0_outputs(2294) <= (inputs(110)) and not (inputs(2));
    layer0_outputs(2295) <= (inputs(158)) or (inputs(203));
    layer0_outputs(2296) <= inputs(153);
    layer0_outputs(2297) <= '1';
    layer0_outputs(2298) <= not(inputs(254)) or (inputs(1));
    layer0_outputs(2299) <= '0';
    layer0_outputs(2300) <= '0';
    layer0_outputs(2301) <= not(inputs(64)) or (inputs(14));
    layer0_outputs(2302) <= '1';
    layer0_outputs(2303) <= (inputs(190)) or (inputs(214));
    layer0_outputs(2304) <= inputs(68);
    layer0_outputs(2305) <= (inputs(217)) and not (inputs(233));
    layer0_outputs(2306) <= (inputs(168)) or (inputs(183));
    layer0_outputs(2307) <= inputs(112);
    layer0_outputs(2308) <= inputs(168);
    layer0_outputs(2309) <= inputs(173);
    layer0_outputs(2310) <= not(inputs(107)) or (inputs(90));
    layer0_outputs(2311) <= not(inputs(25));
    layer0_outputs(2312) <= inputs(14);
    layer0_outputs(2313) <= not(inputs(26));
    layer0_outputs(2314) <= inputs(152);
    layer0_outputs(2315) <= not((inputs(97)) or (inputs(116)));
    layer0_outputs(2316) <= inputs(30);
    layer0_outputs(2317) <= not((inputs(27)) or (inputs(144)));
    layer0_outputs(2318) <= (inputs(34)) and not (inputs(65));
    layer0_outputs(2319) <= not(inputs(102)) or (inputs(32));
    layer0_outputs(2320) <= not(inputs(219));
    layer0_outputs(2321) <= not(inputs(180));
    layer0_outputs(2322) <= '0';
    layer0_outputs(2323) <= (inputs(120)) and (inputs(23));
    layer0_outputs(2324) <= not(inputs(72));
    layer0_outputs(2325) <= inputs(213);
    layer0_outputs(2326) <= inputs(167);
    layer0_outputs(2327) <= not(inputs(13));
    layer0_outputs(2328) <= (inputs(21)) and not (inputs(124));
    layer0_outputs(2329) <= inputs(98);
    layer0_outputs(2330) <= (inputs(211)) and not (inputs(105));
    layer0_outputs(2331) <= (inputs(51)) xor (inputs(242));
    layer0_outputs(2332) <= '0';
    layer0_outputs(2333) <= (inputs(59)) or (inputs(182));
    layer0_outputs(2334) <= (inputs(35)) and not (inputs(245));
    layer0_outputs(2335) <= not(inputs(225));
    layer0_outputs(2336) <= inputs(25);
    layer0_outputs(2337) <= (inputs(197)) and not (inputs(54));
    layer0_outputs(2338) <= inputs(25);
    layer0_outputs(2339) <= not((inputs(50)) and (inputs(40)));
    layer0_outputs(2340) <= (inputs(29)) and not (inputs(214));
    layer0_outputs(2341) <= not(inputs(154)) or (inputs(207));
    layer0_outputs(2342) <= (inputs(161)) or (inputs(39));
    layer0_outputs(2343) <= not((inputs(192)) or (inputs(159)));
    layer0_outputs(2344) <= not(inputs(37)) or (inputs(204));
    layer0_outputs(2345) <= (inputs(237)) and not (inputs(81));
    layer0_outputs(2346) <= (inputs(253)) or (inputs(164));
    layer0_outputs(2347) <= not((inputs(174)) or (inputs(102)));
    layer0_outputs(2348) <= (inputs(243)) and not (inputs(50));
    layer0_outputs(2349) <= inputs(74);
    layer0_outputs(2350) <= (inputs(138)) or (inputs(15));
    layer0_outputs(2351) <= inputs(60);
    layer0_outputs(2352) <= '1';
    layer0_outputs(2353) <= not(inputs(56));
    layer0_outputs(2354) <= not((inputs(81)) xor (inputs(76)));
    layer0_outputs(2355) <= not((inputs(177)) and (inputs(7)));
    layer0_outputs(2356) <= not((inputs(82)) xor (inputs(198)));
    layer0_outputs(2357) <= not(inputs(20));
    layer0_outputs(2358) <= '0';
    layer0_outputs(2359) <= not(inputs(142));
    layer0_outputs(2360) <= (inputs(18)) and not (inputs(33));
    layer0_outputs(2361) <= (inputs(60)) and not (inputs(243));
    layer0_outputs(2362) <= inputs(150);
    layer0_outputs(2363) <= not((inputs(122)) or (inputs(109)));
    layer0_outputs(2364) <= not((inputs(62)) or (inputs(238)));
    layer0_outputs(2365) <= not(inputs(245)) or (inputs(126));
    layer0_outputs(2366) <= not((inputs(107)) and (inputs(40)));
    layer0_outputs(2367) <= not(inputs(99));
    layer0_outputs(2368) <= (inputs(149)) or (inputs(151));
    layer0_outputs(2369) <= (inputs(37)) and not (inputs(113));
    layer0_outputs(2370) <= inputs(17);
    layer0_outputs(2371) <= not(inputs(92));
    layer0_outputs(2372) <= not(inputs(26)) or (inputs(153));
    layer0_outputs(2373) <= not((inputs(87)) and (inputs(5)));
    layer0_outputs(2374) <= not((inputs(5)) xor (inputs(97)));
    layer0_outputs(2375) <= not((inputs(61)) xor (inputs(127)));
    layer0_outputs(2376) <= (inputs(120)) and not (inputs(129));
    layer0_outputs(2377) <= not(inputs(138)) or (inputs(115));
    layer0_outputs(2378) <= (inputs(145)) and not (inputs(31));
    layer0_outputs(2379) <= (inputs(98)) and not (inputs(107));
    layer0_outputs(2380) <= not(inputs(189));
    layer0_outputs(2381) <= inputs(130);
    layer0_outputs(2382) <= not(inputs(143));
    layer0_outputs(2383) <= not((inputs(82)) and (inputs(95)));
    layer0_outputs(2384) <= (inputs(202)) or (inputs(172));
    layer0_outputs(2385) <= not((inputs(211)) or (inputs(238)));
    layer0_outputs(2386) <= not(inputs(117));
    layer0_outputs(2387) <= not((inputs(108)) or (inputs(131)));
    layer0_outputs(2388) <= inputs(205);
    layer0_outputs(2389) <= inputs(65);
    layer0_outputs(2390) <= not(inputs(230)) or (inputs(157));
    layer0_outputs(2391) <= (inputs(173)) xor (inputs(194));
    layer0_outputs(2392) <= inputs(29);
    layer0_outputs(2393) <= not(inputs(104)) or (inputs(186));
    layer0_outputs(2394) <= '0';
    layer0_outputs(2395) <= inputs(105);
    layer0_outputs(2396) <= (inputs(33)) and (inputs(86));
    layer0_outputs(2397) <= not(inputs(228)) or (inputs(67));
    layer0_outputs(2398) <= not((inputs(115)) and (inputs(250)));
    layer0_outputs(2399) <= inputs(228);
    layer0_outputs(2400) <= not((inputs(32)) or (inputs(8)));
    layer0_outputs(2401) <= '1';
    layer0_outputs(2402) <= (inputs(114)) xor (inputs(210));
    layer0_outputs(2403) <= (inputs(118)) and not (inputs(45));
    layer0_outputs(2404) <= inputs(68);
    layer0_outputs(2405) <= (inputs(38)) or (inputs(191));
    layer0_outputs(2406) <= (inputs(1)) or (inputs(32));
    layer0_outputs(2407) <= not(inputs(115)) or (inputs(236));
    layer0_outputs(2408) <= not(inputs(213));
    layer0_outputs(2409) <= '1';
    layer0_outputs(2410) <= not((inputs(187)) or (inputs(237)));
    layer0_outputs(2411) <= (inputs(14)) or (inputs(160));
    layer0_outputs(2412) <= inputs(208);
    layer0_outputs(2413) <= (inputs(93)) and not (inputs(120));
    layer0_outputs(2414) <= not(inputs(190)) or (inputs(94));
    layer0_outputs(2415) <= inputs(135);
    layer0_outputs(2416) <= (inputs(80)) or (inputs(170));
    layer0_outputs(2417) <= not((inputs(183)) or (inputs(68)));
    layer0_outputs(2418) <= not((inputs(98)) or (inputs(180)));
    layer0_outputs(2419) <= not((inputs(215)) or (inputs(190)));
    layer0_outputs(2420) <= inputs(82);
    layer0_outputs(2421) <= not((inputs(83)) or (inputs(145)));
    layer0_outputs(2422) <= '1';
    layer0_outputs(2423) <= not((inputs(70)) or (inputs(117)));
    layer0_outputs(2424) <= not(inputs(82));
    layer0_outputs(2425) <= inputs(8);
    layer0_outputs(2426) <= inputs(75);
    layer0_outputs(2427) <= not((inputs(85)) or (inputs(152)));
    layer0_outputs(2428) <= not(inputs(168));
    layer0_outputs(2429) <= (inputs(152)) or (inputs(99));
    layer0_outputs(2430) <= inputs(35);
    layer0_outputs(2431) <= not(inputs(85));
    layer0_outputs(2432) <= not((inputs(44)) xor (inputs(91)));
    layer0_outputs(2433) <= inputs(82);
    layer0_outputs(2434) <= not(inputs(206)) or (inputs(143));
    layer0_outputs(2435) <= not(inputs(54)) or (inputs(231));
    layer0_outputs(2436) <= inputs(148);
    layer0_outputs(2437) <= not(inputs(116));
    layer0_outputs(2438) <= not(inputs(45)) or (inputs(106));
    layer0_outputs(2439) <= not(inputs(151));
    layer0_outputs(2440) <= not(inputs(24));
    layer0_outputs(2441) <= '0';
    layer0_outputs(2442) <= not(inputs(37)) or (inputs(174));
    layer0_outputs(2443) <= not(inputs(105));
    layer0_outputs(2444) <= (inputs(255)) and not (inputs(56));
    layer0_outputs(2445) <= (inputs(82)) or (inputs(100));
    layer0_outputs(2446) <= (inputs(173)) and not (inputs(46));
    layer0_outputs(2447) <= (inputs(74)) or (inputs(43));
    layer0_outputs(2448) <= not(inputs(20));
    layer0_outputs(2449) <= not(inputs(66));
    layer0_outputs(2450) <= (inputs(133)) and not (inputs(55));
    layer0_outputs(2451) <= not(inputs(91));
    layer0_outputs(2452) <= not(inputs(203)) or (inputs(96));
    layer0_outputs(2453) <= (inputs(126)) and not (inputs(31));
    layer0_outputs(2454) <= not((inputs(161)) and (inputs(77)));
    layer0_outputs(2455) <= (inputs(234)) or (inputs(122));
    layer0_outputs(2456) <= not(inputs(123));
    layer0_outputs(2457) <= not(inputs(104));
    layer0_outputs(2458) <= (inputs(11)) and not (inputs(28));
    layer0_outputs(2459) <= not(inputs(130)) or (inputs(47));
    layer0_outputs(2460) <= (inputs(51)) or (inputs(79));
    layer0_outputs(2461) <= (inputs(96)) or (inputs(51));
    layer0_outputs(2462) <= (inputs(129)) or (inputs(70));
    layer0_outputs(2463) <= inputs(182);
    layer0_outputs(2464) <= not((inputs(94)) and (inputs(111)));
    layer0_outputs(2465) <= not(inputs(101));
    layer0_outputs(2466) <= not(inputs(114));
    layer0_outputs(2467) <= inputs(102);
    layer0_outputs(2468) <= not((inputs(139)) or (inputs(139)));
    layer0_outputs(2469) <= not(inputs(74));
    layer0_outputs(2470) <= inputs(90);
    layer0_outputs(2471) <= not((inputs(58)) and (inputs(249)));
    layer0_outputs(2472) <= not((inputs(142)) or (inputs(86)));
    layer0_outputs(2473) <= not(inputs(104));
    layer0_outputs(2474) <= (inputs(220)) and (inputs(208));
    layer0_outputs(2475) <= not(inputs(87));
    layer0_outputs(2476) <= '0';
    layer0_outputs(2477) <= (inputs(192)) and not (inputs(58));
    layer0_outputs(2478) <= not((inputs(183)) or (inputs(255)));
    layer0_outputs(2479) <= (inputs(201)) and not (inputs(122));
    layer0_outputs(2480) <= not(inputs(63));
    layer0_outputs(2481) <= (inputs(72)) and not (inputs(222));
    layer0_outputs(2482) <= (inputs(191)) or (inputs(175));
    layer0_outputs(2483) <= not(inputs(87));
    layer0_outputs(2484) <= inputs(24);
    layer0_outputs(2485) <= inputs(120);
    layer0_outputs(2486) <= not((inputs(135)) or (inputs(76)));
    layer0_outputs(2487) <= inputs(197);
    layer0_outputs(2488) <= not((inputs(27)) or (inputs(221)));
    layer0_outputs(2489) <= not(inputs(210));
    layer0_outputs(2490) <= not(inputs(205)) or (inputs(63));
    layer0_outputs(2491) <= not((inputs(15)) or (inputs(55)));
    layer0_outputs(2492) <= not(inputs(184));
    layer0_outputs(2493) <= (inputs(25)) or (inputs(48));
    layer0_outputs(2494) <= '0';
    layer0_outputs(2495) <= inputs(76);
    layer0_outputs(2496) <= not((inputs(100)) and (inputs(252)));
    layer0_outputs(2497) <= not((inputs(131)) and (inputs(86)));
    layer0_outputs(2498) <= not(inputs(236)) or (inputs(252));
    layer0_outputs(2499) <= inputs(190);
    layer0_outputs(2500) <= (inputs(130)) xor (inputs(164));
    layer0_outputs(2501) <= inputs(140);
    layer0_outputs(2502) <= inputs(116);
    layer0_outputs(2503) <= not((inputs(163)) xor (inputs(191)));
    layer0_outputs(2504) <= '0';
    layer0_outputs(2505) <= inputs(2);
    layer0_outputs(2506) <= inputs(240);
    layer0_outputs(2507) <= not((inputs(6)) xor (inputs(174)));
    layer0_outputs(2508) <= not((inputs(193)) or (inputs(64)));
    layer0_outputs(2509) <= not((inputs(166)) and (inputs(128)));
    layer0_outputs(2510) <= (inputs(201)) and not (inputs(5));
    layer0_outputs(2511) <= not(inputs(68)) or (inputs(10));
    layer0_outputs(2512) <= (inputs(5)) and not (inputs(147));
    layer0_outputs(2513) <= inputs(235);
    layer0_outputs(2514) <= (inputs(143)) or (inputs(158));
    layer0_outputs(2515) <= not((inputs(94)) or (inputs(58)));
    layer0_outputs(2516) <= not(inputs(196));
    layer0_outputs(2517) <= '1';
    layer0_outputs(2518) <= not(inputs(184)) or (inputs(47));
    layer0_outputs(2519) <= not((inputs(163)) or (inputs(142)));
    layer0_outputs(2520) <= not(inputs(167));
    layer0_outputs(2521) <= not((inputs(172)) and (inputs(215)));
    layer0_outputs(2522) <= not((inputs(196)) or (inputs(161)));
    layer0_outputs(2523) <= not((inputs(203)) and (inputs(126)));
    layer0_outputs(2524) <= (inputs(253)) and not (inputs(251));
    layer0_outputs(2525) <= inputs(133);
    layer0_outputs(2526) <= not((inputs(89)) or (inputs(28)));
    layer0_outputs(2527) <= not(inputs(80));
    layer0_outputs(2528) <= (inputs(133)) and not (inputs(16));
    layer0_outputs(2529) <= not(inputs(231));
    layer0_outputs(2530) <= not(inputs(238)) or (inputs(18));
    layer0_outputs(2531) <= not(inputs(152));
    layer0_outputs(2532) <= '1';
    layer0_outputs(2533) <= (inputs(229)) and (inputs(240));
    layer0_outputs(2534) <= inputs(208);
    layer0_outputs(2535) <= not(inputs(125)) or (inputs(233));
    layer0_outputs(2536) <= (inputs(71)) and not (inputs(147));
    layer0_outputs(2537) <= not(inputs(252)) or (inputs(236));
    layer0_outputs(2538) <= not((inputs(82)) or (inputs(102)));
    layer0_outputs(2539) <= (inputs(147)) and not (inputs(131));
    layer0_outputs(2540) <= not(inputs(28)) or (inputs(118));
    layer0_outputs(2541) <= not((inputs(248)) xor (inputs(200)));
    layer0_outputs(2542) <= '0';
    layer0_outputs(2543) <= '0';
    layer0_outputs(2544) <= not(inputs(115));
    layer0_outputs(2545) <= not(inputs(91));
    layer0_outputs(2546) <= not((inputs(7)) or (inputs(107)));
    layer0_outputs(2547) <= not(inputs(73));
    layer0_outputs(2548) <= inputs(109);
    layer0_outputs(2549) <= not((inputs(197)) and (inputs(189)));
    layer0_outputs(2550) <= inputs(148);
    layer0_outputs(2551) <= inputs(83);
    layer0_outputs(2552) <= not((inputs(111)) or (inputs(181)));
    layer0_outputs(2553) <= inputs(83);
    layer0_outputs(2554) <= not(inputs(135)) or (inputs(191));
    layer0_outputs(2555) <= inputs(165);
    layer0_outputs(2556) <= (inputs(49)) and not (inputs(81));
    layer0_outputs(2557) <= (inputs(180)) or (inputs(147));
    layer0_outputs(2558) <= not(inputs(90)) or (inputs(221));
    layer0_outputs(2559) <= inputs(166);
    layer1_outputs(0) <= layer0_outputs(1163);
    layer1_outputs(1) <= (layer0_outputs(1232)) and (layer0_outputs(1122));
    layer1_outputs(2) <= not((layer0_outputs(1064)) xor (layer0_outputs(2307)));
    layer1_outputs(3) <= layer0_outputs(1742);
    layer1_outputs(4) <= '1';
    layer1_outputs(5) <= (layer0_outputs(492)) or (layer0_outputs(510));
    layer1_outputs(6) <= not(layer0_outputs(769));
    layer1_outputs(7) <= (layer0_outputs(784)) and not (layer0_outputs(730));
    layer1_outputs(8) <= layer0_outputs(92);
    layer1_outputs(9) <= not(layer0_outputs(808));
    layer1_outputs(10) <= not(layer0_outputs(2219)) or (layer0_outputs(812));
    layer1_outputs(11) <= not((layer0_outputs(1853)) or (layer0_outputs(68)));
    layer1_outputs(12) <= not((layer0_outputs(2080)) or (layer0_outputs(597)));
    layer1_outputs(13) <= not(layer0_outputs(2381));
    layer1_outputs(14) <= not((layer0_outputs(2009)) and (layer0_outputs(696)));
    layer1_outputs(15) <= not(layer0_outputs(1455)) or (layer0_outputs(100));
    layer1_outputs(16) <= (layer0_outputs(1992)) and (layer0_outputs(2219));
    layer1_outputs(17) <= (layer0_outputs(946)) and not (layer0_outputs(1559));
    layer1_outputs(18) <= not(layer0_outputs(2122)) or (layer0_outputs(128));
    layer1_outputs(19) <= not(layer0_outputs(1837));
    layer1_outputs(20) <= not(layer0_outputs(7)) or (layer0_outputs(2104));
    layer1_outputs(21) <= layer0_outputs(722);
    layer1_outputs(22) <= (layer0_outputs(796)) or (layer0_outputs(720));
    layer1_outputs(23) <= (layer0_outputs(676)) and (layer0_outputs(395));
    layer1_outputs(24) <= not((layer0_outputs(458)) xor (layer0_outputs(1558)));
    layer1_outputs(25) <= layer0_outputs(641);
    layer1_outputs(26) <= (layer0_outputs(1482)) or (layer0_outputs(1224));
    layer1_outputs(27) <= (layer0_outputs(898)) and (layer0_outputs(711));
    layer1_outputs(28) <= not(layer0_outputs(2207));
    layer1_outputs(29) <= '0';
    layer1_outputs(30) <= (layer0_outputs(1163)) and not (layer0_outputs(919));
    layer1_outputs(31) <= (layer0_outputs(1920)) or (layer0_outputs(2248));
    layer1_outputs(32) <= (layer0_outputs(1081)) and not (layer0_outputs(1728));
    layer1_outputs(33) <= layer0_outputs(1616);
    layer1_outputs(34) <= layer0_outputs(2440);
    layer1_outputs(35) <= not(layer0_outputs(1051));
    layer1_outputs(36) <= not(layer0_outputs(1961));
    layer1_outputs(37) <= not(layer0_outputs(1735));
    layer1_outputs(38) <= not((layer0_outputs(1600)) or (layer0_outputs(1034)));
    layer1_outputs(39) <= not(layer0_outputs(158)) or (layer0_outputs(1757));
    layer1_outputs(40) <= not((layer0_outputs(1773)) and (layer0_outputs(2555)));
    layer1_outputs(41) <= (layer0_outputs(2335)) and (layer0_outputs(1784));
    layer1_outputs(42) <= not(layer0_outputs(314));
    layer1_outputs(43) <= '1';
    layer1_outputs(44) <= layer0_outputs(412);
    layer1_outputs(45) <= not(layer0_outputs(1393));
    layer1_outputs(46) <= layer0_outputs(1283);
    layer1_outputs(47) <= not(layer0_outputs(1703));
    layer1_outputs(48) <= (layer0_outputs(363)) and not (layer0_outputs(2331));
    layer1_outputs(49) <= '1';
    layer1_outputs(50) <= not(layer0_outputs(2320));
    layer1_outputs(51) <= (layer0_outputs(1659)) and (layer0_outputs(1912));
    layer1_outputs(52) <= (layer0_outputs(506)) or (layer0_outputs(1856));
    layer1_outputs(53) <= (layer0_outputs(239)) and not (layer0_outputs(119));
    layer1_outputs(54) <= not(layer0_outputs(1145));
    layer1_outputs(55) <= not((layer0_outputs(1460)) or (layer0_outputs(368)));
    layer1_outputs(56) <= (layer0_outputs(1845)) and not (layer0_outputs(1196));
    layer1_outputs(57) <= not((layer0_outputs(2038)) and (layer0_outputs(461)));
    layer1_outputs(58) <= layer0_outputs(1630);
    layer1_outputs(59) <= not(layer0_outputs(1635));
    layer1_outputs(60) <= '0';
    layer1_outputs(61) <= not((layer0_outputs(1784)) and (layer0_outputs(1306)));
    layer1_outputs(62) <= '0';
    layer1_outputs(63) <= layer0_outputs(2035);
    layer1_outputs(64) <= not((layer0_outputs(1359)) and (layer0_outputs(2398)));
    layer1_outputs(65) <= (layer0_outputs(1944)) and not (layer0_outputs(420));
    layer1_outputs(66) <= (layer0_outputs(285)) or (layer0_outputs(413));
    layer1_outputs(67) <= not(layer0_outputs(1274)) or (layer0_outputs(369));
    layer1_outputs(68) <= (layer0_outputs(584)) or (layer0_outputs(2212));
    layer1_outputs(69) <= layer0_outputs(1252);
    layer1_outputs(70) <= not(layer0_outputs(2514));
    layer1_outputs(71) <= layer0_outputs(2319);
    layer1_outputs(72) <= not(layer0_outputs(1487));
    layer1_outputs(73) <= not(layer0_outputs(906));
    layer1_outputs(74) <= (layer0_outputs(659)) and not (layer0_outputs(1459));
    layer1_outputs(75) <= (layer0_outputs(2124)) and not (layer0_outputs(802));
    layer1_outputs(76) <= layer0_outputs(2326);
    layer1_outputs(77) <= not((layer0_outputs(1523)) and (layer0_outputs(2490)));
    layer1_outputs(78) <= (layer0_outputs(1873)) and not (layer0_outputs(1113));
    layer1_outputs(79) <= not(layer0_outputs(795));
    layer1_outputs(80) <= not(layer0_outputs(585));
    layer1_outputs(81) <= (layer0_outputs(1901)) and (layer0_outputs(239));
    layer1_outputs(82) <= (layer0_outputs(390)) or (layer0_outputs(1893));
    layer1_outputs(83) <= not(layer0_outputs(1707));
    layer1_outputs(84) <= (layer0_outputs(264)) and not (layer0_outputs(790));
    layer1_outputs(85) <= layer0_outputs(273);
    layer1_outputs(86) <= (layer0_outputs(2406)) and not (layer0_outputs(2157));
    layer1_outputs(87) <= (layer0_outputs(1408)) and (layer0_outputs(1960));
    layer1_outputs(88) <= not(layer0_outputs(1240));
    layer1_outputs(89) <= layer0_outputs(33);
    layer1_outputs(90) <= (layer0_outputs(1466)) and not (layer0_outputs(2459));
    layer1_outputs(91) <= layer0_outputs(1438);
    layer1_outputs(92) <= (layer0_outputs(2277)) and (layer0_outputs(1548));
    layer1_outputs(93) <= not(layer0_outputs(1947));
    layer1_outputs(94) <= not(layer0_outputs(1018));
    layer1_outputs(95) <= layer0_outputs(2453);
    layer1_outputs(96) <= not((layer0_outputs(1599)) and (layer0_outputs(1976)));
    layer1_outputs(97) <= not((layer0_outputs(2179)) or (layer0_outputs(832)));
    layer1_outputs(98) <= not(layer0_outputs(1587)) or (layer0_outputs(605));
    layer1_outputs(99) <= not(layer0_outputs(999));
    layer1_outputs(100) <= (layer0_outputs(105)) or (layer0_outputs(1445));
    layer1_outputs(101) <= not((layer0_outputs(701)) and (layer0_outputs(1536)));
    layer1_outputs(102) <= (layer0_outputs(2507)) and not (layer0_outputs(355));
    layer1_outputs(103) <= not(layer0_outputs(1792)) or (layer0_outputs(358));
    layer1_outputs(104) <= layer0_outputs(1179);
    layer1_outputs(105) <= layer0_outputs(1794);
    layer1_outputs(106) <= (layer0_outputs(666)) and not (layer0_outputs(1589));
    layer1_outputs(107) <= layer0_outputs(2398);
    layer1_outputs(108) <= not((layer0_outputs(1956)) and (layer0_outputs(488)));
    layer1_outputs(109) <= not((layer0_outputs(1314)) and (layer0_outputs(2187)));
    layer1_outputs(110) <= not(layer0_outputs(2066));
    layer1_outputs(111) <= (layer0_outputs(1378)) and not (layer0_outputs(1285));
    layer1_outputs(112) <= not(layer0_outputs(2216));
    layer1_outputs(113) <= not(layer0_outputs(969)) or (layer0_outputs(659));
    layer1_outputs(114) <= layer0_outputs(2240);
    layer1_outputs(115) <= not((layer0_outputs(1226)) or (layer0_outputs(633)));
    layer1_outputs(116) <= layer0_outputs(1689);
    layer1_outputs(117) <= '1';
    layer1_outputs(118) <= (layer0_outputs(1174)) or (layer0_outputs(1192));
    layer1_outputs(119) <= not(layer0_outputs(462));
    layer1_outputs(120) <= (layer0_outputs(524)) and (layer0_outputs(72));
    layer1_outputs(121) <= not(layer0_outputs(152));
    layer1_outputs(122) <= layer0_outputs(1299);
    layer1_outputs(123) <= not(layer0_outputs(1793));
    layer1_outputs(124) <= not(layer0_outputs(1778));
    layer1_outputs(125) <= not(layer0_outputs(2339)) or (layer0_outputs(1081));
    layer1_outputs(126) <= layer0_outputs(377);
    layer1_outputs(127) <= not((layer0_outputs(2116)) xor (layer0_outputs(1957)));
    layer1_outputs(128) <= layer0_outputs(112);
    layer1_outputs(129) <= not((layer0_outputs(207)) or (layer0_outputs(1680)));
    layer1_outputs(130) <= not(layer0_outputs(2269));
    layer1_outputs(131) <= (layer0_outputs(1066)) and not (layer0_outputs(2465));
    layer1_outputs(132) <= layer0_outputs(755);
    layer1_outputs(133) <= layer0_outputs(1051);
    layer1_outputs(134) <= not((layer0_outputs(1618)) and (layer0_outputs(869)));
    layer1_outputs(135) <= not(layer0_outputs(388)) or (layer0_outputs(560));
    layer1_outputs(136) <= not(layer0_outputs(1940));
    layer1_outputs(137) <= not(layer0_outputs(2069)) or (layer0_outputs(691));
    layer1_outputs(138) <= layer0_outputs(2494);
    layer1_outputs(139) <= '1';
    layer1_outputs(140) <= not(layer0_outputs(27));
    layer1_outputs(141) <= not(layer0_outputs(1785)) or (layer0_outputs(1514));
    layer1_outputs(142) <= not(layer0_outputs(2341));
    layer1_outputs(143) <= not(layer0_outputs(1326)) or (layer0_outputs(1237));
    layer1_outputs(144) <= layer0_outputs(1508);
    layer1_outputs(145) <= layer0_outputs(624);
    layer1_outputs(146) <= not(layer0_outputs(1589)) or (layer0_outputs(348));
    layer1_outputs(147) <= not(layer0_outputs(2434)) or (layer0_outputs(1895));
    layer1_outputs(148) <= layer0_outputs(223);
    layer1_outputs(149) <= (layer0_outputs(1444)) and not (layer0_outputs(2134));
    layer1_outputs(150) <= (layer0_outputs(1911)) or (layer0_outputs(210));
    layer1_outputs(151) <= (layer0_outputs(1934)) or (layer0_outputs(1198));
    layer1_outputs(152) <= not(layer0_outputs(1815));
    layer1_outputs(153) <= not((layer0_outputs(192)) or (layer0_outputs(1626)));
    layer1_outputs(154) <= not(layer0_outputs(2434));
    layer1_outputs(155) <= (layer0_outputs(2086)) and (layer0_outputs(2038));
    layer1_outputs(156) <= layer0_outputs(1777);
    layer1_outputs(157) <= not(layer0_outputs(427));
    layer1_outputs(158) <= not(layer0_outputs(306));
    layer1_outputs(159) <= layer0_outputs(1204);
    layer1_outputs(160) <= not(layer0_outputs(279));
    layer1_outputs(161) <= (layer0_outputs(1882)) or (layer0_outputs(922));
    layer1_outputs(162) <= '1';
    layer1_outputs(163) <= '0';
    layer1_outputs(164) <= (layer0_outputs(1315)) and not (layer0_outputs(354));
    layer1_outputs(165) <= (layer0_outputs(2548)) and not (layer0_outputs(591));
    layer1_outputs(166) <= (layer0_outputs(1033)) and not (layer0_outputs(1748));
    layer1_outputs(167) <= layer0_outputs(357);
    layer1_outputs(168) <= not(layer0_outputs(594)) or (layer0_outputs(60));
    layer1_outputs(169) <= not(layer0_outputs(0)) or (layer0_outputs(1817));
    layer1_outputs(170) <= not((layer0_outputs(2538)) or (layer0_outputs(1459)));
    layer1_outputs(171) <= not(layer0_outputs(2410));
    layer1_outputs(172) <= (layer0_outputs(43)) and not (layer0_outputs(1043));
    layer1_outputs(173) <= (layer0_outputs(2222)) and not (layer0_outputs(2363));
    layer1_outputs(174) <= (layer0_outputs(1849)) and not (layer0_outputs(1867));
    layer1_outputs(175) <= (layer0_outputs(1280)) and (layer0_outputs(253));
    layer1_outputs(176) <= (layer0_outputs(1161)) and not (layer0_outputs(49));
    layer1_outputs(177) <= not((layer0_outputs(2463)) or (layer0_outputs(948)));
    layer1_outputs(178) <= '0';
    layer1_outputs(179) <= not(layer0_outputs(376));
    layer1_outputs(180) <= layer0_outputs(1606);
    layer1_outputs(181) <= layer0_outputs(92);
    layer1_outputs(182) <= (layer0_outputs(930)) xor (layer0_outputs(2065));
    layer1_outputs(183) <= (layer0_outputs(1980)) and (layer0_outputs(1700));
    layer1_outputs(184) <= not(layer0_outputs(2545));
    layer1_outputs(185) <= (layer0_outputs(2403)) and (layer0_outputs(188));
    layer1_outputs(186) <= not(layer0_outputs(1353)) or (layer0_outputs(772));
    layer1_outputs(187) <= layer0_outputs(69);
    layer1_outputs(188) <= layer0_outputs(1031);
    layer1_outputs(189) <= not(layer0_outputs(917)) or (layer0_outputs(680));
    layer1_outputs(190) <= not(layer0_outputs(2043));
    layer1_outputs(191) <= layer0_outputs(902);
    layer1_outputs(192) <= not(layer0_outputs(508)) or (layer0_outputs(2477));
    layer1_outputs(193) <= not((layer0_outputs(1203)) or (layer0_outputs(891)));
    layer1_outputs(194) <= not(layer0_outputs(1943));
    layer1_outputs(195) <= layer0_outputs(351);
    layer1_outputs(196) <= not(layer0_outputs(844)) or (layer0_outputs(545));
    layer1_outputs(197) <= layer0_outputs(1628);
    layer1_outputs(198) <= (layer0_outputs(1104)) and not (layer0_outputs(96));
    layer1_outputs(199) <= (layer0_outputs(1295)) or (layer0_outputs(193));
    layer1_outputs(200) <= layer0_outputs(1301);
    layer1_outputs(201) <= '1';
    layer1_outputs(202) <= not(layer0_outputs(2137));
    layer1_outputs(203) <= layer0_outputs(340);
    layer1_outputs(204) <= (layer0_outputs(1836)) or (layer0_outputs(923));
    layer1_outputs(205) <= (layer0_outputs(1851)) or (layer0_outputs(290));
    layer1_outputs(206) <= '0';
    layer1_outputs(207) <= not(layer0_outputs(1783));
    layer1_outputs(208) <= (layer0_outputs(1236)) and not (layer0_outputs(1910));
    layer1_outputs(209) <= not((layer0_outputs(170)) and (layer0_outputs(2300)));
    layer1_outputs(210) <= layer0_outputs(2296);
    layer1_outputs(211) <= (layer0_outputs(976)) or (layer0_outputs(1512));
    layer1_outputs(212) <= not(layer0_outputs(1003));
    layer1_outputs(213) <= '0';
    layer1_outputs(214) <= layer0_outputs(1687);
    layer1_outputs(215) <= layer0_outputs(1010);
    layer1_outputs(216) <= layer0_outputs(1386);
    layer1_outputs(217) <= (layer0_outputs(2100)) and not (layer0_outputs(246));
    layer1_outputs(218) <= layer0_outputs(657);
    layer1_outputs(219) <= layer0_outputs(453);
    layer1_outputs(220) <= (layer0_outputs(859)) or (layer0_outputs(1588));
    layer1_outputs(221) <= not(layer0_outputs(151));
    layer1_outputs(222) <= not(layer0_outputs(740)) or (layer0_outputs(1065));
    layer1_outputs(223) <= (layer0_outputs(1316)) and not (layer0_outputs(1311));
    layer1_outputs(224) <= layer0_outputs(1150);
    layer1_outputs(225) <= (layer0_outputs(787)) and not (layer0_outputs(1710));
    layer1_outputs(226) <= not(layer0_outputs(1208));
    layer1_outputs(227) <= (layer0_outputs(1947)) xor (layer0_outputs(1092));
    layer1_outputs(228) <= not(layer0_outputs(2287)) or (layer0_outputs(1402));
    layer1_outputs(229) <= not(layer0_outputs(157)) or (layer0_outputs(1441));
    layer1_outputs(230) <= (layer0_outputs(1621)) and not (layer0_outputs(823));
    layer1_outputs(231) <= not(layer0_outputs(2000)) or (layer0_outputs(478));
    layer1_outputs(232) <= (layer0_outputs(279)) or (layer0_outputs(2105));
    layer1_outputs(233) <= layer0_outputs(1292);
    layer1_outputs(234) <= not(layer0_outputs(1669)) or (layer0_outputs(2033));
    layer1_outputs(235) <= not(layer0_outputs(2325));
    layer1_outputs(236) <= (layer0_outputs(104)) or (layer0_outputs(125));
    layer1_outputs(237) <= layer0_outputs(1488);
    layer1_outputs(238) <= not(layer0_outputs(1786));
    layer1_outputs(239) <= layer0_outputs(1824);
    layer1_outputs(240) <= not(layer0_outputs(142));
    layer1_outputs(241) <= not((layer0_outputs(1613)) and (layer0_outputs(626)));
    layer1_outputs(242) <= not(layer0_outputs(114)) or (layer0_outputs(473));
    layer1_outputs(243) <= (layer0_outputs(1524)) and not (layer0_outputs(1619));
    layer1_outputs(244) <= (layer0_outputs(1396)) and not (layer0_outputs(1889));
    layer1_outputs(245) <= (layer0_outputs(1888)) and (layer0_outputs(406));
    layer1_outputs(246) <= layer0_outputs(820);
    layer1_outputs(247) <= (layer0_outputs(1210)) and not (layer0_outputs(1191));
    layer1_outputs(248) <= '1';
    layer1_outputs(249) <= not((layer0_outputs(1672)) xor (layer0_outputs(1061)));
    layer1_outputs(250) <= not((layer0_outputs(2338)) or (layer0_outputs(2188)));
    layer1_outputs(251) <= not(layer0_outputs(260));
    layer1_outputs(252) <= not(layer0_outputs(1662)) or (layer0_outputs(2304));
    layer1_outputs(253) <= not((layer0_outputs(430)) and (layer0_outputs(818)));
    layer1_outputs(254) <= layer0_outputs(1058);
    layer1_outputs(255) <= (layer0_outputs(590)) and not (layer0_outputs(2184));
    layer1_outputs(256) <= (layer0_outputs(763)) and not (layer0_outputs(1966));
    layer1_outputs(257) <= '1';
    layer1_outputs(258) <= not(layer0_outputs(1269)) or (layer0_outputs(1236));
    layer1_outputs(259) <= (layer0_outputs(248)) and not (layer0_outputs(2089));
    layer1_outputs(260) <= not(layer0_outputs(1102));
    layer1_outputs(261) <= not(layer0_outputs(765));
    layer1_outputs(262) <= not((layer0_outputs(1862)) and (layer0_outputs(1218)));
    layer1_outputs(263) <= not(layer0_outputs(752)) or (layer0_outputs(1038));
    layer1_outputs(264) <= not((layer0_outputs(270)) and (layer0_outputs(1008)));
    layer1_outputs(265) <= not((layer0_outputs(2476)) and (layer0_outputs(1573)));
    layer1_outputs(266) <= not(layer0_outputs(1177)) or (layer0_outputs(853));
    layer1_outputs(267) <= (layer0_outputs(1322)) and not (layer0_outputs(2379));
    layer1_outputs(268) <= not(layer0_outputs(1788)) or (layer0_outputs(1376));
    layer1_outputs(269) <= not((layer0_outputs(1190)) and (layer0_outputs(108)));
    layer1_outputs(270) <= (layer0_outputs(168)) and not (layer0_outputs(1465));
    layer1_outputs(271) <= not(layer0_outputs(2456));
    layer1_outputs(272) <= not(layer0_outputs(1301));
    layer1_outputs(273) <= not(layer0_outputs(1618));
    layer1_outputs(274) <= (layer0_outputs(2292)) or (layer0_outputs(229));
    layer1_outputs(275) <= not((layer0_outputs(2101)) or (layer0_outputs(810)));
    layer1_outputs(276) <= (layer0_outputs(153)) and (layer0_outputs(1580));
    layer1_outputs(277) <= layer0_outputs(1085);
    layer1_outputs(278) <= layer0_outputs(781);
    layer1_outputs(279) <= not((layer0_outputs(662)) or (layer0_outputs(1195)));
    layer1_outputs(280) <= not(layer0_outputs(600));
    layer1_outputs(281) <= not(layer0_outputs(1543)) or (layer0_outputs(2350));
    layer1_outputs(282) <= not(layer0_outputs(316)) or (layer0_outputs(2223));
    layer1_outputs(283) <= not((layer0_outputs(1303)) and (layer0_outputs(2317)));
    layer1_outputs(284) <= layer0_outputs(1121);
    layer1_outputs(285) <= layer0_outputs(52);
    layer1_outputs(286) <= not(layer0_outputs(687)) or (layer0_outputs(703));
    layer1_outputs(287) <= layer0_outputs(1870);
    layer1_outputs(288) <= layer0_outputs(1909);
    layer1_outputs(289) <= '0';
    layer1_outputs(290) <= (layer0_outputs(602)) xor (layer0_outputs(2304));
    layer1_outputs(291) <= not(layer0_outputs(2416));
    layer1_outputs(292) <= (layer0_outputs(1157)) and not (layer0_outputs(1379));
    layer1_outputs(293) <= (layer0_outputs(1840)) and not (layer0_outputs(1753));
    layer1_outputs(294) <= (layer0_outputs(364)) and (layer0_outputs(1062));
    layer1_outputs(295) <= not((layer0_outputs(1811)) or (layer0_outputs(657)));
    layer1_outputs(296) <= not(layer0_outputs(864)) or (layer0_outputs(566));
    layer1_outputs(297) <= not(layer0_outputs(318));
    layer1_outputs(298) <= not(layer0_outputs(758)) or (layer0_outputs(1451));
    layer1_outputs(299) <= layer0_outputs(384);
    layer1_outputs(300) <= layer0_outputs(695);
    layer1_outputs(301) <= not(layer0_outputs(2259));
    layer1_outputs(302) <= '1';
    layer1_outputs(303) <= '0';
    layer1_outputs(304) <= not(layer0_outputs(1484));
    layer1_outputs(305) <= layer0_outputs(1358);
    layer1_outputs(306) <= (layer0_outputs(1157)) and not (layer0_outputs(2031));
    layer1_outputs(307) <= not(layer0_outputs(529));
    layer1_outputs(308) <= not(layer0_outputs(711));
    layer1_outputs(309) <= not(layer0_outputs(1025));
    layer1_outputs(310) <= not((layer0_outputs(1223)) and (layer0_outputs(574)));
    layer1_outputs(311) <= not(layer0_outputs(251));
    layer1_outputs(312) <= (layer0_outputs(2108)) or (layer0_outputs(737));
    layer1_outputs(313) <= layer0_outputs(1841);
    layer1_outputs(314) <= (layer0_outputs(2518)) and (layer0_outputs(1456));
    layer1_outputs(315) <= '0';
    layer1_outputs(316) <= (layer0_outputs(1595)) and not (layer0_outputs(1603));
    layer1_outputs(317) <= not((layer0_outputs(2147)) or (layer0_outputs(1488)));
    layer1_outputs(318) <= (layer0_outputs(1512)) xor (layer0_outputs(411));
    layer1_outputs(319) <= layer0_outputs(276);
    layer1_outputs(320) <= not(layer0_outputs(2447));
    layer1_outputs(321) <= not(layer0_outputs(2549)) or (layer0_outputs(2344));
    layer1_outputs(322) <= layer0_outputs(1518);
    layer1_outputs(323) <= layer0_outputs(1251);
    layer1_outputs(324) <= not(layer0_outputs(137));
    layer1_outputs(325) <= not(layer0_outputs(1199)) or (layer0_outputs(535));
    layer1_outputs(326) <= (layer0_outputs(2385)) and (layer0_outputs(759));
    layer1_outputs(327) <= not(layer0_outputs(1793));
    layer1_outputs(328) <= (layer0_outputs(1063)) and (layer0_outputs(874));
    layer1_outputs(329) <= layer0_outputs(1788);
    layer1_outputs(330) <= '1';
    layer1_outputs(331) <= (layer0_outputs(2274)) and not (layer0_outputs(1540));
    layer1_outputs(332) <= (layer0_outputs(2512)) or (layer0_outputs(770));
    layer1_outputs(333) <= '1';
    layer1_outputs(334) <= not(layer0_outputs(830)) or (layer0_outputs(1272));
    layer1_outputs(335) <= not((layer0_outputs(1731)) or (layer0_outputs(798)));
    layer1_outputs(336) <= not((layer0_outputs(1565)) and (layer0_outputs(499)));
    layer1_outputs(337) <= not(layer0_outputs(1635)) or (layer0_outputs(497));
    layer1_outputs(338) <= (layer0_outputs(1569)) and not (layer0_outputs(996));
    layer1_outputs(339) <= not((layer0_outputs(519)) and (layer0_outputs(1826)));
    layer1_outputs(340) <= (layer0_outputs(1442)) or (layer0_outputs(1053));
    layer1_outputs(341) <= (layer0_outputs(1713)) xor (layer0_outputs(2547));
    layer1_outputs(342) <= not(layer0_outputs(410));
    layer1_outputs(343) <= not(layer0_outputs(1343));
    layer1_outputs(344) <= not(layer0_outputs(1065));
    layer1_outputs(345) <= not(layer0_outputs(1141));
    layer1_outputs(346) <= not((layer0_outputs(2529)) and (layer0_outputs(1368)));
    layer1_outputs(347) <= not(layer0_outputs(1137)) or (layer0_outputs(511));
    layer1_outputs(348) <= not(layer0_outputs(2241)) or (layer0_outputs(1056));
    layer1_outputs(349) <= not(layer0_outputs(101));
    layer1_outputs(350) <= not(layer0_outputs(838));
    layer1_outputs(351) <= layer0_outputs(1818);
    layer1_outputs(352) <= '0';
    layer1_outputs(353) <= '1';
    layer1_outputs(354) <= not((layer0_outputs(664)) and (layer0_outputs(550)));
    layer1_outputs(355) <= not((layer0_outputs(1425)) and (layer0_outputs(1465)));
    layer1_outputs(356) <= (layer0_outputs(1760)) and not (layer0_outputs(1278));
    layer1_outputs(357) <= not((layer0_outputs(1287)) and (layer0_outputs(1033)));
    layer1_outputs(358) <= (layer0_outputs(1908)) or (layer0_outputs(129));
    layer1_outputs(359) <= '0';
    layer1_outputs(360) <= (layer0_outputs(1808)) and not (layer0_outputs(1822));
    layer1_outputs(361) <= not(layer0_outputs(1802));
    layer1_outputs(362) <= not(layer0_outputs(592));
    layer1_outputs(363) <= '0';
    layer1_outputs(364) <= (layer0_outputs(338)) and (layer0_outputs(1097));
    layer1_outputs(365) <= layer0_outputs(1107);
    layer1_outputs(366) <= (layer0_outputs(2013)) or (layer0_outputs(824));
    layer1_outputs(367) <= layer0_outputs(242);
    layer1_outputs(368) <= (layer0_outputs(589)) and not (layer0_outputs(678));
    layer1_outputs(369) <= (layer0_outputs(2252)) or (layer0_outputs(1207));
    layer1_outputs(370) <= (layer0_outputs(2242)) and not (layer0_outputs(733));
    layer1_outputs(371) <= not(layer0_outputs(1202));
    layer1_outputs(372) <= '0';
    layer1_outputs(373) <= (layer0_outputs(621)) or (layer0_outputs(1705));
    layer1_outputs(374) <= not(layer0_outputs(449)) or (layer0_outputs(304));
    layer1_outputs(375) <= (layer0_outputs(894)) and (layer0_outputs(1133));
    layer1_outputs(376) <= not(layer0_outputs(1920));
    layer1_outputs(377) <= '0';
    layer1_outputs(378) <= (layer0_outputs(1835)) and not (layer0_outputs(466));
    layer1_outputs(379) <= (layer0_outputs(20)) or (layer0_outputs(2505));
    layer1_outputs(380) <= layer0_outputs(1965);
    layer1_outputs(381) <= layer0_outputs(371);
    layer1_outputs(382) <= not((layer0_outputs(400)) or (layer0_outputs(2357)));
    layer1_outputs(383) <= (layer0_outputs(1718)) or (layer0_outputs(1115));
    layer1_outputs(384) <= layer0_outputs(503);
    layer1_outputs(385) <= not(layer0_outputs(2276));
    layer1_outputs(386) <= (layer0_outputs(951)) and not (layer0_outputs(1962));
    layer1_outputs(387) <= (layer0_outputs(1481)) and not (layer0_outputs(792));
    layer1_outputs(388) <= (layer0_outputs(1164)) and not (layer0_outputs(2224));
    layer1_outputs(389) <= (layer0_outputs(1803)) and not (layer0_outputs(800));
    layer1_outputs(390) <= layer0_outputs(1190);
    layer1_outputs(391) <= layer0_outputs(2052);
    layer1_outputs(392) <= '0';
    layer1_outputs(393) <= layer0_outputs(99);
    layer1_outputs(394) <= not(layer0_outputs(457)) or (layer0_outputs(1490));
    layer1_outputs(395) <= '0';
    layer1_outputs(396) <= not((layer0_outputs(186)) and (layer0_outputs(2353)));
    layer1_outputs(397) <= (layer0_outputs(1134)) and (layer0_outputs(2469));
    layer1_outputs(398) <= layer0_outputs(1333);
    layer1_outputs(399) <= layer0_outputs(2008);
    layer1_outputs(400) <= not(layer0_outputs(1046));
    layer1_outputs(401) <= layer0_outputs(727);
    layer1_outputs(402) <= not(layer0_outputs(485));
    layer1_outputs(403) <= not(layer0_outputs(1216));
    layer1_outputs(404) <= (layer0_outputs(1894)) and not (layer0_outputs(1109));
    layer1_outputs(405) <= (layer0_outputs(876)) and not (layer0_outputs(623));
    layer1_outputs(406) <= layer0_outputs(1254);
    layer1_outputs(407) <= '1';
    layer1_outputs(408) <= (layer0_outputs(2391)) or (layer0_outputs(904));
    layer1_outputs(409) <= not((layer0_outputs(926)) or (layer0_outputs(1991)));
    layer1_outputs(410) <= (layer0_outputs(1929)) and not (layer0_outputs(269));
    layer1_outputs(411) <= (layer0_outputs(2389)) or (layer0_outputs(175));
    layer1_outputs(412) <= not((layer0_outputs(544)) or (layer0_outputs(1256)));
    layer1_outputs(413) <= not(layer0_outputs(930));
    layer1_outputs(414) <= not(layer0_outputs(2218));
    layer1_outputs(415) <= (layer0_outputs(1937)) and (layer0_outputs(498));
    layer1_outputs(416) <= layer0_outputs(836);
    layer1_outputs(417) <= not(layer0_outputs(2360)) or (layer0_outputs(619));
    layer1_outputs(418) <= layer0_outputs(826);
    layer1_outputs(419) <= not(layer0_outputs(542));
    layer1_outputs(420) <= layer0_outputs(378);
    layer1_outputs(421) <= (layer0_outputs(2124)) and (layer0_outputs(548));
    layer1_outputs(422) <= not((layer0_outputs(874)) and (layer0_outputs(2114)));
    layer1_outputs(423) <= not(layer0_outputs(2382));
    layer1_outputs(424) <= not((layer0_outputs(103)) and (layer0_outputs(938)));
    layer1_outputs(425) <= (layer0_outputs(703)) or (layer0_outputs(1768));
    layer1_outputs(426) <= (layer0_outputs(330)) or (layer0_outputs(1771));
    layer1_outputs(427) <= not(layer0_outputs(1136));
    layer1_outputs(428) <= not(layer0_outputs(866));
    layer1_outputs(429) <= (layer0_outputs(1400)) and not (layer0_outputs(2368));
    layer1_outputs(430) <= (layer0_outputs(1954)) and (layer0_outputs(1497));
    layer1_outputs(431) <= not((layer0_outputs(2210)) or (layer0_outputs(2253)));
    layer1_outputs(432) <= not(layer0_outputs(150));
    layer1_outputs(433) <= layer0_outputs(1152);
    layer1_outputs(434) <= not(layer0_outputs(1894));
    layer1_outputs(435) <= layer0_outputs(207);
    layer1_outputs(436) <= not(layer0_outputs(2002)) or (layer0_outputs(64));
    layer1_outputs(437) <= (layer0_outputs(1135)) and not (layer0_outputs(2039));
    layer1_outputs(438) <= layer0_outputs(1382);
    layer1_outputs(439) <= not(layer0_outputs(1930));
    layer1_outputs(440) <= not(layer0_outputs(1390));
    layer1_outputs(441) <= (layer0_outputs(1640)) or (layer0_outputs(1069));
    layer1_outputs(442) <= not(layer0_outputs(67));
    layer1_outputs(443) <= not(layer0_outputs(1056)) or (layer0_outputs(1227));
    layer1_outputs(444) <= '0';
    layer1_outputs(445) <= layer0_outputs(2256);
    layer1_outputs(446) <= not(layer0_outputs(1974)) or (layer0_outputs(1866));
    layer1_outputs(447) <= (layer0_outputs(50)) and not (layer0_outputs(2483));
    layer1_outputs(448) <= not(layer0_outputs(1276)) or (layer0_outputs(394));
    layer1_outputs(449) <= not(layer0_outputs(1834));
    layer1_outputs(450) <= not(layer0_outputs(1944));
    layer1_outputs(451) <= not((layer0_outputs(754)) or (layer0_outputs(2496)));
    layer1_outputs(452) <= (layer0_outputs(1966)) and (layer0_outputs(266));
    layer1_outputs(453) <= layer0_outputs(1746);
    layer1_outputs(454) <= (layer0_outputs(244)) or (layer0_outputs(1670));
    layer1_outputs(455) <= not(layer0_outputs(1935));
    layer1_outputs(456) <= layer0_outputs(1423);
    layer1_outputs(457) <= (layer0_outputs(1054)) or (layer0_outputs(1109));
    layer1_outputs(458) <= not((layer0_outputs(887)) or (layer0_outputs(2174)));
    layer1_outputs(459) <= not(layer0_outputs(2485));
    layer1_outputs(460) <= layer0_outputs(448);
    layer1_outputs(461) <= not(layer0_outputs(605));
    layer1_outputs(462) <= (layer0_outputs(1883)) and not (layer0_outputs(1789));
    layer1_outputs(463) <= layer0_outputs(754);
    layer1_outputs(464) <= not(layer0_outputs(1855)) or (layer0_outputs(183));
    layer1_outputs(465) <= layer0_outputs(1175);
    layer1_outputs(466) <= (layer0_outputs(1925)) and not (layer0_outputs(297));
    layer1_outputs(467) <= not(layer0_outputs(51));
    layer1_outputs(468) <= (layer0_outputs(2507)) and not (layer0_outputs(147));
    layer1_outputs(469) <= not(layer0_outputs(1036));
    layer1_outputs(470) <= (layer0_outputs(138)) and (layer0_outputs(2546));
    layer1_outputs(471) <= layer0_outputs(1000);
    layer1_outputs(472) <= layer0_outputs(2059);
    layer1_outputs(473) <= (layer0_outputs(2098)) and not (layer0_outputs(581));
    layer1_outputs(474) <= not((layer0_outputs(1620)) and (layer0_outputs(71)));
    layer1_outputs(475) <= (layer0_outputs(262)) and not (layer0_outputs(2342));
    layer1_outputs(476) <= not((layer0_outputs(2458)) and (layer0_outputs(2316)));
    layer1_outputs(477) <= '1';
    layer1_outputs(478) <= (layer0_outputs(1678)) and not (layer0_outputs(86));
    layer1_outputs(479) <= (layer0_outputs(1913)) and not (layer0_outputs(389));
    layer1_outputs(480) <= not(layer0_outputs(2235)) or (layer0_outputs(376));
    layer1_outputs(481) <= not(layer0_outputs(1782));
    layer1_outputs(482) <= not((layer0_outputs(1030)) and (layer0_outputs(1047)));
    layer1_outputs(483) <= layer0_outputs(1517);
    layer1_outputs(484) <= (layer0_outputs(841)) or (layer0_outputs(226));
    layer1_outputs(485) <= layer0_outputs(2008);
    layer1_outputs(486) <= not(layer0_outputs(2487)) or (layer0_outputs(774));
    layer1_outputs(487) <= not(layer0_outputs(148));
    layer1_outputs(488) <= not((layer0_outputs(2420)) or (layer0_outputs(2251)));
    layer1_outputs(489) <= (layer0_outputs(762)) and not (layer0_outputs(2556));
    layer1_outputs(490) <= (layer0_outputs(484)) and (layer0_outputs(1541));
    layer1_outputs(491) <= not(layer0_outputs(630));
    layer1_outputs(492) <= not(layer0_outputs(114));
    layer1_outputs(493) <= '0';
    layer1_outputs(494) <= layer0_outputs(246);
    layer1_outputs(495) <= not(layer0_outputs(1730)) or (layer0_outputs(883));
    layer1_outputs(496) <= layer0_outputs(145);
    layer1_outputs(497) <= (layer0_outputs(2365)) or (layer0_outputs(1202));
    layer1_outputs(498) <= (layer0_outputs(690)) and not (layer0_outputs(619));
    layer1_outputs(499) <= (layer0_outputs(430)) and (layer0_outputs(722));
    layer1_outputs(500) <= layer0_outputs(1289);
    layer1_outputs(501) <= not(layer0_outputs(790)) or (layer0_outputs(2333));
    layer1_outputs(502) <= layer0_outputs(63);
    layer1_outputs(503) <= '0';
    layer1_outputs(504) <= not(layer0_outputs(1235)) or (layer0_outputs(167));
    layer1_outputs(505) <= (layer0_outputs(1475)) and (layer0_outputs(1060));
    layer1_outputs(506) <= (layer0_outputs(2158)) and (layer0_outputs(68));
    layer1_outputs(507) <= '0';
    layer1_outputs(508) <= not(layer0_outputs(217));
    layer1_outputs(509) <= not(layer0_outputs(406));
    layer1_outputs(510) <= not((layer0_outputs(1530)) and (layer0_outputs(1738)));
    layer1_outputs(511) <= not(layer0_outputs(501));
    layer1_outputs(512) <= (layer0_outputs(159)) and not (layer0_outputs(810));
    layer1_outputs(513) <= (layer0_outputs(552)) and (layer0_outputs(2125));
    layer1_outputs(514) <= (layer0_outputs(1118)) and not (layer0_outputs(1686));
    layer1_outputs(515) <= (layer0_outputs(1862)) and (layer0_outputs(1586));
    layer1_outputs(516) <= not(layer0_outputs(1532));
    layer1_outputs(517) <= layer0_outputs(1333);
    layer1_outputs(518) <= (layer0_outputs(752)) or (layer0_outputs(767));
    layer1_outputs(519) <= (layer0_outputs(1602)) or (layer0_outputs(1120));
    layer1_outputs(520) <= '0';
    layer1_outputs(521) <= not(layer0_outputs(521)) or (layer0_outputs(1717));
    layer1_outputs(522) <= '0';
    layer1_outputs(523) <= (layer0_outputs(313)) and (layer0_outputs(1798));
    layer1_outputs(524) <= (layer0_outputs(1088)) and (layer0_outputs(1994));
    layer1_outputs(525) <= '0';
    layer1_outputs(526) <= layer0_outputs(339);
    layer1_outputs(527) <= not(layer0_outputs(508));
    layer1_outputs(528) <= not(layer0_outputs(772));
    layer1_outputs(529) <= (layer0_outputs(2520)) and not (layer0_outputs(261));
    layer1_outputs(530) <= not((layer0_outputs(843)) xor (layer0_outputs(151)));
    layer1_outputs(531) <= not(layer0_outputs(2014)) or (layer0_outputs(565));
    layer1_outputs(532) <= (layer0_outputs(653)) and not (layer0_outputs(2368));
    layer1_outputs(533) <= not(layer0_outputs(1246)) or (layer0_outputs(922));
    layer1_outputs(534) <= '1';
    layer1_outputs(535) <= layer0_outputs(1368);
    layer1_outputs(536) <= not(layer0_outputs(646));
    layer1_outputs(537) <= '1';
    layer1_outputs(538) <= layer0_outputs(78);
    layer1_outputs(539) <= not((layer0_outputs(1664)) and (layer0_outputs(1708)));
    layer1_outputs(540) <= layer0_outputs(1258);
    layer1_outputs(541) <= not((layer0_outputs(228)) and (layer0_outputs(1562)));
    layer1_outputs(542) <= not(layer0_outputs(1919));
    layer1_outputs(543) <= layer0_outputs(872);
    layer1_outputs(544) <= not(layer0_outputs(1951));
    layer1_outputs(545) <= (layer0_outputs(1850)) and (layer0_outputs(2341));
    layer1_outputs(546) <= (layer0_outputs(972)) and not (layer0_outputs(2030));
    layer1_outputs(547) <= layer0_outputs(1724);
    layer1_outputs(548) <= not(layer0_outputs(1902));
    layer1_outputs(549) <= layer0_outputs(814);
    layer1_outputs(550) <= '0';
    layer1_outputs(551) <= not(layer0_outputs(522));
    layer1_outputs(552) <= not((layer0_outputs(1761)) and (layer0_outputs(434)));
    layer1_outputs(553) <= layer0_outputs(1996);
    layer1_outputs(554) <= (layer0_outputs(1108)) and not (layer0_outputs(1458));
    layer1_outputs(555) <= '1';
    layer1_outputs(556) <= (layer0_outputs(446)) and (layer0_outputs(1649));
    layer1_outputs(557) <= not(layer0_outputs(1529));
    layer1_outputs(558) <= (layer0_outputs(2359)) and not (layer0_outputs(2205));
    layer1_outputs(559) <= (layer0_outputs(255)) or (layer0_outputs(1632));
    layer1_outputs(560) <= layer0_outputs(1015);
    layer1_outputs(561) <= not(layer0_outputs(1868));
    layer1_outputs(562) <= not(layer0_outputs(1344));
    layer1_outputs(563) <= not((layer0_outputs(2449)) or (layer0_outputs(949)));
    layer1_outputs(564) <= not((layer0_outputs(316)) and (layer0_outputs(2140)));
    layer1_outputs(565) <= not(layer0_outputs(1767)) or (layer0_outputs(2349));
    layer1_outputs(566) <= not(layer0_outputs(1864));
    layer1_outputs(567) <= not((layer0_outputs(1587)) and (layer0_outputs(1047)));
    layer1_outputs(568) <= layer0_outputs(215);
    layer1_outputs(569) <= (layer0_outputs(1740)) or (layer0_outputs(384));
    layer1_outputs(570) <= '1';
    layer1_outputs(571) <= (layer0_outputs(1102)) and not (layer0_outputs(1073));
    layer1_outputs(572) <= not(layer0_outputs(1915));
    layer1_outputs(573) <= (layer0_outputs(1519)) or (layer0_outputs(1392));
    layer1_outputs(574) <= not((layer0_outputs(1107)) or (layer0_outputs(2137)));
    layer1_outputs(575) <= not(layer0_outputs(82));
    layer1_outputs(576) <= not(layer0_outputs(2313));
    layer1_outputs(577) <= layer0_outputs(1252);
    layer1_outputs(578) <= layer0_outputs(918);
    layer1_outputs(579) <= layer0_outputs(311);
    layer1_outputs(580) <= layer0_outputs(214);
    layer1_outputs(581) <= (layer0_outputs(106)) xor (layer0_outputs(902));
    layer1_outputs(582) <= (layer0_outputs(539)) or (layer0_outputs(2254));
    layer1_outputs(583) <= (layer0_outputs(839)) and not (layer0_outputs(1726));
    layer1_outputs(584) <= '0';
    layer1_outputs(585) <= not(layer0_outputs(2178));
    layer1_outputs(586) <= (layer0_outputs(2428)) and not (layer0_outputs(1357));
    layer1_outputs(587) <= (layer0_outputs(2144)) or (layer0_outputs(1745));
    layer1_outputs(588) <= not(layer0_outputs(2511)) or (layer0_outputs(47));
    layer1_outputs(589) <= '1';
    layer1_outputs(590) <= not(layer0_outputs(2298)) or (layer0_outputs(191));
    layer1_outputs(591) <= layer0_outputs(1201);
    layer1_outputs(592) <= (layer0_outputs(953)) and (layer0_outputs(251));
    layer1_outputs(593) <= '1';
    layer1_outputs(594) <= not(layer0_outputs(2171));
    layer1_outputs(595) <= not(layer0_outputs(672));
    layer1_outputs(596) <= not((layer0_outputs(2519)) and (layer0_outputs(815)));
    layer1_outputs(597) <= not(layer0_outputs(2076)) or (layer0_outputs(15));
    layer1_outputs(598) <= layer0_outputs(1617);
    layer1_outputs(599) <= (layer0_outputs(52)) and not (layer0_outputs(133));
    layer1_outputs(600) <= not((layer0_outputs(751)) and (layer0_outputs(1828)));
    layer1_outputs(601) <= '0';
    layer1_outputs(602) <= not(layer0_outputs(1526)) or (layer0_outputs(1008));
    layer1_outputs(603) <= (layer0_outputs(1153)) or (layer0_outputs(1140));
    layer1_outputs(604) <= (layer0_outputs(514)) or (layer0_outputs(2052));
    layer1_outputs(605) <= layer0_outputs(637);
    layer1_outputs(606) <= not(layer0_outputs(1665)) or (layer0_outputs(1509));
    layer1_outputs(607) <= not(layer0_outputs(1785));
    layer1_outputs(608) <= layer0_outputs(551);
    layer1_outputs(609) <= not(layer0_outputs(1783)) or (layer0_outputs(383));
    layer1_outputs(610) <= not(layer0_outputs(295));
    layer1_outputs(611) <= layer0_outputs(617);
    layer1_outputs(612) <= not((layer0_outputs(1871)) or (layer0_outputs(1045)));
    layer1_outputs(613) <= (layer0_outputs(558)) or (layer0_outputs(1375));
    layer1_outputs(614) <= (layer0_outputs(2472)) and not (layer0_outputs(596));
    layer1_outputs(615) <= (layer0_outputs(127)) and (layer0_outputs(1510));
    layer1_outputs(616) <= not((layer0_outputs(678)) and (layer0_outputs(2106)));
    layer1_outputs(617) <= (layer0_outputs(1415)) and not (layer0_outputs(1964));
    layer1_outputs(618) <= (layer0_outputs(1076)) and not (layer0_outputs(1774));
    layer1_outputs(619) <= (layer0_outputs(399)) and not (layer0_outputs(1810));
    layer1_outputs(620) <= '1';
    layer1_outputs(621) <= layer0_outputs(1473);
    layer1_outputs(622) <= layer0_outputs(2448);
    layer1_outputs(623) <= (layer0_outputs(861)) and not (layer0_outputs(785));
    layer1_outputs(624) <= not(layer0_outputs(814)) or (layer0_outputs(1285));
    layer1_outputs(625) <= (layer0_outputs(364)) and not (layer0_outputs(586));
    layer1_outputs(626) <= layer0_outputs(824);
    layer1_outputs(627) <= not(layer0_outputs(778));
    layer1_outputs(628) <= (layer0_outputs(736)) and not (layer0_outputs(2536));
    layer1_outputs(629) <= (layer0_outputs(160)) or (layer0_outputs(1420));
    layer1_outputs(630) <= (layer0_outputs(2074)) or (layer0_outputs(1365));
    layer1_outputs(631) <= layer0_outputs(699);
    layer1_outputs(632) <= (layer0_outputs(1497)) or (layer0_outputs(785));
    layer1_outputs(633) <= layer0_outputs(2215);
    layer1_outputs(634) <= layer0_outputs(799);
    layer1_outputs(635) <= layer0_outputs(154);
    layer1_outputs(636) <= layer0_outputs(608);
    layer1_outputs(637) <= not(layer0_outputs(1547)) or (layer0_outputs(1113));
    layer1_outputs(638) <= (layer0_outputs(2233)) xor (layer0_outputs(17));
    layer1_outputs(639) <= layer0_outputs(331);
    layer1_outputs(640) <= not((layer0_outputs(2238)) or (layer0_outputs(2160)));
    layer1_outputs(641) <= layer0_outputs(2000);
    layer1_outputs(642) <= (layer0_outputs(2111)) and (layer0_outputs(878));
    layer1_outputs(643) <= not(layer0_outputs(1068));
    layer1_outputs(644) <= not((layer0_outputs(2439)) or (layer0_outputs(2175)));
    layer1_outputs(645) <= layer0_outputs(718);
    layer1_outputs(646) <= not((layer0_outputs(1667)) or (layer0_outputs(1945)));
    layer1_outputs(647) <= layer0_outputs(677);
    layer1_outputs(648) <= not(layer0_outputs(2559));
    layer1_outputs(649) <= not(layer0_outputs(2374)) or (layer0_outputs(2206));
    layer1_outputs(650) <= not((layer0_outputs(1356)) and (layer0_outputs(70)));
    layer1_outputs(651) <= not(layer0_outputs(2136)) or (layer0_outputs(2091));
    layer1_outputs(652) <= (layer0_outputs(2486)) and not (layer0_outputs(451));
    layer1_outputs(653) <= not((layer0_outputs(2390)) and (layer0_outputs(1170)));
    layer1_outputs(654) <= (layer0_outputs(2359)) and not (layer0_outputs(983));
    layer1_outputs(655) <= not(layer0_outputs(1796));
    layer1_outputs(656) <= (layer0_outputs(2094)) and not (layer0_outputs(89));
    layer1_outputs(657) <= layer0_outputs(98);
    layer1_outputs(658) <= (layer0_outputs(2074)) or (layer0_outputs(1069));
    layer1_outputs(659) <= not(layer0_outputs(1823));
    layer1_outputs(660) <= not(layer0_outputs(757));
    layer1_outputs(661) <= not(layer0_outputs(379));
    layer1_outputs(662) <= (layer0_outputs(1129)) and not (layer0_outputs(1164));
    layer1_outputs(663) <= not((layer0_outputs(2510)) xor (layer0_outputs(197)));
    layer1_outputs(664) <= (layer0_outputs(2003)) or (layer0_outputs(1006));
    layer1_outputs(665) <= not(layer0_outputs(791));
    layer1_outputs(666) <= (layer0_outputs(240)) and (layer0_outputs(2538));
    layer1_outputs(667) <= (layer0_outputs(359)) and not (layer0_outputs(2452));
    layer1_outputs(668) <= (layer0_outputs(1623)) or (layer0_outputs(640));
    layer1_outputs(669) <= layer0_outputs(2285);
    layer1_outputs(670) <= (layer0_outputs(173)) and not (layer0_outputs(1138));
    layer1_outputs(671) <= (layer0_outputs(947)) and (layer0_outputs(1591));
    layer1_outputs(672) <= not(layer0_outputs(1450));
    layer1_outputs(673) <= not(layer0_outputs(681));
    layer1_outputs(674) <= (layer0_outputs(134)) and not (layer0_outputs(1401));
    layer1_outputs(675) <= (layer0_outputs(1479)) or (layer0_outputs(1217));
    layer1_outputs(676) <= not((layer0_outputs(2192)) and (layer0_outputs(1715)));
    layer1_outputs(677) <= not(layer0_outputs(208)) or (layer0_outputs(2402));
    layer1_outputs(678) <= not((layer0_outputs(968)) or (layer0_outputs(1288)));
    layer1_outputs(679) <= (layer0_outputs(2213)) and not (layer0_outputs(1536));
    layer1_outputs(680) <= layer0_outputs(1032);
    layer1_outputs(681) <= (layer0_outputs(40)) and not (layer0_outputs(2023));
    layer1_outputs(682) <= (layer0_outputs(1060)) and (layer0_outputs(1525));
    layer1_outputs(683) <= not(layer0_outputs(1168));
    layer1_outputs(684) <= (layer0_outputs(1591)) and not (layer0_outputs(1257));
    layer1_outputs(685) <= not((layer0_outputs(2211)) or (layer0_outputs(682)));
    layer1_outputs(686) <= '0';
    layer1_outputs(687) <= not((layer0_outputs(79)) or (layer0_outputs(1637)));
    layer1_outputs(688) <= not(layer0_outputs(1402));
    layer1_outputs(689) <= (layer0_outputs(2386)) and not (layer0_outputs(1449));
    layer1_outputs(690) <= layer0_outputs(1068);
    layer1_outputs(691) <= '1';
    layer1_outputs(692) <= not(layer0_outputs(628));
    layer1_outputs(693) <= not(layer0_outputs(491)) or (layer0_outputs(1115));
    layer1_outputs(694) <= not(layer0_outputs(1503));
    layer1_outputs(695) <= not(layer0_outputs(980)) or (layer0_outputs(257));
    layer1_outputs(696) <= layer0_outputs(850);
    layer1_outputs(697) <= not((layer0_outputs(171)) or (layer0_outputs(1263)));
    layer1_outputs(698) <= not(layer0_outputs(660));
    layer1_outputs(699) <= layer0_outputs(1763);
    layer1_outputs(700) <= not(layer0_outputs(2306));
    layer1_outputs(701) <= (layer0_outputs(2557)) or (layer0_outputs(409));
    layer1_outputs(702) <= layer0_outputs(738);
    layer1_outputs(703) <= layer0_outputs(2343);
    layer1_outputs(704) <= not(layer0_outputs(1835));
    layer1_outputs(705) <= (layer0_outputs(887)) or (layer0_outputs(140));
    layer1_outputs(706) <= '1';
    layer1_outputs(707) <= not(layer0_outputs(2414)) or (layer0_outputs(2163));
    layer1_outputs(708) <= (layer0_outputs(570)) and (layer0_outputs(1119));
    layer1_outputs(709) <= not((layer0_outputs(397)) xor (layer0_outputs(1432)));
    layer1_outputs(710) <= not(layer0_outputs(1562));
    layer1_outputs(711) <= layer0_outputs(325);
    layer1_outputs(712) <= not((layer0_outputs(474)) xor (layer0_outputs(1279)));
    layer1_outputs(713) <= not(layer0_outputs(1744));
    layer1_outputs(714) <= not(layer0_outputs(1461)) or (layer0_outputs(451));
    layer1_outputs(715) <= '1';
    layer1_outputs(716) <= not((layer0_outputs(1998)) and (layer0_outputs(1189)));
    layer1_outputs(717) <= not(layer0_outputs(1091)) or (layer0_outputs(450));
    layer1_outputs(718) <= not((layer0_outputs(1417)) or (layer0_outputs(2280)));
    layer1_outputs(719) <= layer0_outputs(1258);
    layer1_outputs(720) <= (layer0_outputs(1310)) or (layer0_outputs(2319));
    layer1_outputs(721) <= not(layer0_outputs(225)) or (layer0_outputs(1761));
    layer1_outputs(722) <= layer0_outputs(702);
    layer1_outputs(723) <= layer0_outputs(650);
    layer1_outputs(724) <= not(layer0_outputs(1217));
    layer1_outputs(725) <= layer0_outputs(1486);
    layer1_outputs(726) <= (layer0_outputs(39)) or (layer0_outputs(414));
    layer1_outputs(727) <= not((layer0_outputs(1428)) and (layer0_outputs(370)));
    layer1_outputs(728) <= not(layer0_outputs(1870));
    layer1_outputs(729) <= layer0_outputs(399);
    layer1_outputs(730) <= not(layer0_outputs(1212)) or (layer0_outputs(700));
    layer1_outputs(731) <= (layer0_outputs(1755)) or (layer0_outputs(1334));
    layer1_outputs(732) <= (layer0_outputs(318)) and (layer0_outputs(55));
    layer1_outputs(733) <= not(layer0_outputs(1502)) or (layer0_outputs(2269));
    layer1_outputs(734) <= not(layer0_outputs(2466));
    layer1_outputs(735) <= layer0_outputs(2548);
    layer1_outputs(736) <= not(layer0_outputs(1832));
    layer1_outputs(737) <= '0';
    layer1_outputs(738) <= not(layer0_outputs(1194));
    layer1_outputs(739) <= not(layer0_outputs(580)) or (layer0_outputs(2075));
    layer1_outputs(740) <= (layer0_outputs(1633)) xor (layer0_outputs(1806));
    layer1_outputs(741) <= layer0_outputs(1430);
    layer1_outputs(742) <= not((layer0_outputs(534)) and (layer0_outputs(2079)));
    layer1_outputs(743) <= not(layer0_outputs(613)) or (layer0_outputs(2363));
    layer1_outputs(744) <= layer0_outputs(2355);
    layer1_outputs(745) <= layer0_outputs(1686);
    layer1_outputs(746) <= not(layer0_outputs(483)) or (layer0_outputs(2255));
    layer1_outputs(747) <= '1';
    layer1_outputs(748) <= (layer0_outputs(220)) and (layer0_outputs(903));
    layer1_outputs(749) <= not(layer0_outputs(1753)) or (layer0_outputs(1011));
    layer1_outputs(750) <= (layer0_outputs(515)) and not (layer0_outputs(1989));
    layer1_outputs(751) <= layer0_outputs(448);
    layer1_outputs(752) <= (layer0_outputs(229)) and not (layer0_outputs(93));
    layer1_outputs(753) <= not(layer0_outputs(444));
    layer1_outputs(754) <= (layer0_outputs(1071)) and (layer0_outputs(2135));
    layer1_outputs(755) <= not((layer0_outputs(1479)) or (layer0_outputs(418)));
    layer1_outputs(756) <= (layer0_outputs(1243)) and not (layer0_outputs(1887));
    layer1_outputs(757) <= (layer0_outputs(2451)) and not (layer0_outputs(1545));
    layer1_outputs(758) <= '0';
    layer1_outputs(759) <= not(layer0_outputs(1192)) or (layer0_outputs(1022));
    layer1_outputs(760) <= not(layer0_outputs(778));
    layer1_outputs(761) <= (layer0_outputs(1089)) and (layer0_outputs(1391));
    layer1_outputs(762) <= (layer0_outputs(2353)) or (layer0_outputs(236));
    layer1_outputs(763) <= not(layer0_outputs(1813));
    layer1_outputs(764) <= (layer0_outputs(2029)) or (layer0_outputs(1026));
    layer1_outputs(765) <= not(layer0_outputs(460));
    layer1_outputs(766) <= layer0_outputs(2199);
    layer1_outputs(767) <= not(layer0_outputs(2531));
    layer1_outputs(768) <= layer0_outputs(857);
    layer1_outputs(769) <= not((layer0_outputs(1711)) and (layer0_outputs(1656)));
    layer1_outputs(770) <= layer0_outputs(701);
    layer1_outputs(771) <= (layer0_outputs(773)) and (layer0_outputs(2131));
    layer1_outputs(772) <= not(layer0_outputs(1083)) or (layer0_outputs(786));
    layer1_outputs(773) <= layer0_outputs(18);
    layer1_outputs(774) <= (layer0_outputs(442)) and not (layer0_outputs(2375));
    layer1_outputs(775) <= (layer0_outputs(1906)) and not (layer0_outputs(291));
    layer1_outputs(776) <= layer0_outputs(1416);
    layer1_outputs(777) <= not((layer0_outputs(523)) and (layer0_outputs(337)));
    layer1_outputs(778) <= layer0_outputs(238);
    layer1_outputs(779) <= not((layer0_outputs(989)) or (layer0_outputs(689)));
    layer1_outputs(780) <= (layer0_outputs(1580)) and (layer0_outputs(973));
    layer1_outputs(781) <= layer0_outputs(2268);
    layer1_outputs(782) <= (layer0_outputs(1674)) and not (layer0_outputs(2506));
    layer1_outputs(783) <= (layer0_outputs(2519)) and (layer0_outputs(1597));
    layer1_outputs(784) <= not(layer0_outputs(1415));
    layer1_outputs(785) <= (layer0_outputs(2427)) and not (layer0_outputs(1940));
    layer1_outputs(786) <= layer0_outputs(1972);
    layer1_outputs(787) <= not((layer0_outputs(295)) and (layer0_outputs(1813)));
    layer1_outputs(788) <= not(layer0_outputs(28));
    layer1_outputs(789) <= not(layer0_outputs(2455)) or (layer0_outputs(2329));
    layer1_outputs(790) <= not(layer0_outputs(1214));
    layer1_outputs(791) <= '0';
    layer1_outputs(792) <= '1';
    layer1_outputs(793) <= not(layer0_outputs(417));
    layer1_outputs(794) <= layer0_outputs(72);
    layer1_outputs(795) <= layer0_outputs(610);
    layer1_outputs(796) <= not(layer0_outputs(863));
    layer1_outputs(797) <= '1';
    layer1_outputs(798) <= (layer0_outputs(1119)) or (layer0_outputs(210));
    layer1_outputs(799) <= not(layer0_outputs(1798)) or (layer0_outputs(825));
    layer1_outputs(800) <= not((layer0_outputs(267)) or (layer0_outputs(2232)));
    layer1_outputs(801) <= not(layer0_outputs(1064));
    layer1_outputs(802) <= not(layer0_outputs(1253));
    layer1_outputs(803) <= (layer0_outputs(1688)) and (layer0_outputs(837));
    layer1_outputs(804) <= (layer0_outputs(893)) and (layer0_outputs(482));
    layer1_outputs(805) <= not((layer0_outputs(858)) and (layer0_outputs(704)));
    layer1_outputs(806) <= (layer0_outputs(1879)) and not (layer0_outputs(827));
    layer1_outputs(807) <= not((layer0_outputs(2416)) or (layer0_outputs(113)));
    layer1_outputs(808) <= (layer0_outputs(904)) and (layer0_outputs(749));
    layer1_outputs(809) <= (layer0_outputs(1828)) and not (layer0_outputs(1896));
    layer1_outputs(810) <= (layer0_outputs(487)) and not (layer0_outputs(2072));
    layer1_outputs(811) <= '0';
    layer1_outputs(812) <= (layer0_outputs(2432)) and (layer0_outputs(1903));
    layer1_outputs(813) <= not(layer0_outputs(2244));
    layer1_outputs(814) <= not(layer0_outputs(1983));
    layer1_outputs(815) <= not((layer0_outputs(1489)) or (layer0_outputs(2305)));
    layer1_outputs(816) <= (layer0_outputs(1264)) and not (layer0_outputs(563));
    layer1_outputs(817) <= '1';
    layer1_outputs(818) <= not(layer0_outputs(1787));
    layer1_outputs(819) <= not(layer0_outputs(1993)) or (layer0_outputs(2342));
    layer1_outputs(820) <= not(layer0_outputs(1548)) or (layer0_outputs(2446));
    layer1_outputs(821) <= not(layer0_outputs(319));
    layer1_outputs(822) <= not(layer0_outputs(884));
    layer1_outputs(823) <= not(layer0_outputs(708)) or (layer0_outputs(840));
    layer1_outputs(824) <= (layer0_outputs(1719)) and (layer0_outputs(408));
    layer1_outputs(825) <= layer0_outputs(2288);
    layer1_outputs(826) <= (layer0_outputs(760)) and (layer0_outputs(1557));
    layer1_outputs(827) <= not((layer0_outputs(996)) or (layer0_outputs(574)));
    layer1_outputs(828) <= not((layer0_outputs(2006)) or (layer0_outputs(1116)));
    layer1_outputs(829) <= not((layer0_outputs(1082)) and (layer0_outputs(2522)));
    layer1_outputs(830) <= (layer0_outputs(309)) and not (layer0_outputs(1121));
    layer1_outputs(831) <= layer0_outputs(935);
    layer1_outputs(832) <= not(layer0_outputs(600));
    layer1_outputs(833) <= layer0_outputs(2017);
    layer1_outputs(834) <= not(layer0_outputs(721));
    layer1_outputs(835) <= (layer0_outputs(1344)) and not (layer0_outputs(2357));
    layer1_outputs(836) <= layer0_outputs(1262);
    layer1_outputs(837) <= not(layer0_outputs(2558)) or (layer0_outputs(1773));
    layer1_outputs(838) <= (layer0_outputs(1280)) and not (layer0_outputs(714));
    layer1_outputs(839) <= layer0_outputs(440);
    layer1_outputs(840) <= not((layer0_outputs(2243)) and (layer0_outputs(1967)));
    layer1_outputs(841) <= (layer0_outputs(750)) xor (layer0_outputs(1298));
    layer1_outputs(842) <= not((layer0_outputs(658)) or (layer0_outputs(2190)));
    layer1_outputs(843) <= layer0_outputs(505);
    layer1_outputs(844) <= not(layer0_outputs(477)) or (layer0_outputs(1227));
    layer1_outputs(845) <= not(layer0_outputs(206)) or (layer0_outputs(665));
    layer1_outputs(846) <= layer0_outputs(334);
    layer1_outputs(847) <= not(layer0_outputs(195)) or (layer0_outputs(315));
    layer1_outputs(848) <= not(layer0_outputs(1437));
    layer1_outputs(849) <= not(layer0_outputs(1225)) or (layer0_outputs(836));
    layer1_outputs(850) <= not((layer0_outputs(2371)) and (layer0_outputs(1775)));
    layer1_outputs(851) <= not(layer0_outputs(1211));
    layer1_outputs(852) <= (layer0_outputs(798)) and not (layer0_outputs(1582));
    layer1_outputs(853) <= not((layer0_outputs(907)) or (layer0_outputs(199)));
    layer1_outputs(854) <= layer0_outputs(2149);
    layer1_outputs(855) <= (layer0_outputs(2465)) and not (layer0_outputs(1340));
    layer1_outputs(856) <= layer0_outputs(474);
    layer1_outputs(857) <= not(layer0_outputs(2234));
    layer1_outputs(858) <= layer0_outputs(1126);
    layer1_outputs(859) <= layer0_outputs(1086);
    layer1_outputs(860) <= not((layer0_outputs(2013)) or (layer0_outputs(2179)));
    layer1_outputs(861) <= not((layer0_outputs(1077)) and (layer0_outputs(1237)));
    layer1_outputs(862) <= not(layer0_outputs(946));
    layer1_outputs(863) <= not(layer0_outputs(822));
    layer1_outputs(864) <= layer0_outputs(957);
    layer1_outputs(865) <= not((layer0_outputs(391)) and (layer0_outputs(615)));
    layer1_outputs(866) <= (layer0_outputs(2367)) and (layer0_outputs(317));
    layer1_outputs(867) <= not(layer0_outputs(2177)) or (layer0_outputs(1663));
    layer1_outputs(868) <= '1';
    layer1_outputs(869) <= layer0_outputs(1114);
    layer1_outputs(870) <= not(layer0_outputs(1361));
    layer1_outputs(871) <= layer0_outputs(1726);
    layer1_outputs(872) <= layer0_outputs(1801);
    layer1_outputs(873) <= layer0_outputs(889);
    layer1_outputs(874) <= not(layer0_outputs(2387));
    layer1_outputs(875) <= layer0_outputs(1308);
    layer1_outputs(876) <= (layer0_outputs(1040)) and not (layer0_outputs(1229));
    layer1_outputs(877) <= '1';
    layer1_outputs(878) <= not((layer0_outputs(827)) xor (layer0_outputs(2369)));
    layer1_outputs(879) <= layer0_outputs(341);
    layer1_outputs(880) <= (layer0_outputs(363)) or (layer0_outputs(2386));
    layer1_outputs(881) <= (layer0_outputs(2097)) or (layer0_outputs(2290));
    layer1_outputs(882) <= not((layer0_outputs(748)) and (layer0_outputs(1714)));
    layer1_outputs(883) <= (layer0_outputs(1585)) and not (layer0_outputs(418));
    layer1_outputs(884) <= layer0_outputs(1013);
    layer1_outputs(885) <= not(layer0_outputs(1440)) or (layer0_outputs(793));
    layer1_outputs(886) <= not((layer0_outputs(2404)) or (layer0_outputs(1952)));
    layer1_outputs(887) <= layer0_outputs(583);
    layer1_outputs(888) <= not(layer0_outputs(1439));
    layer1_outputs(889) <= not((layer0_outputs(576)) and (layer0_outputs(2092)));
    layer1_outputs(890) <= (layer0_outputs(190)) and (layer0_outputs(57));
    layer1_outputs(891) <= '1';
    layer1_outputs(892) <= not(layer0_outputs(1649)) or (layer0_outputs(2413));
    layer1_outputs(893) <= '0';
    layer1_outputs(894) <= (layer0_outputs(1105)) or (layer0_outputs(1313));
    layer1_outputs(895) <= layer0_outputs(1953);
    layer1_outputs(896) <= (layer0_outputs(564)) and not (layer0_outputs(1733));
    layer1_outputs(897) <= not(layer0_outputs(277));
    layer1_outputs(898) <= (layer0_outputs(1892)) and (layer0_outputs(320));
    layer1_outputs(899) <= (layer0_outputs(2090)) and not (layer0_outputs(1106));
    layer1_outputs(900) <= not(layer0_outputs(2176)) or (layer0_outputs(129));
    layer1_outputs(901) <= (layer0_outputs(402)) and not (layer0_outputs(1572));
    layer1_outputs(902) <= layer0_outputs(2119);
    layer1_outputs(903) <= layer0_outputs(490);
    layer1_outputs(904) <= not((layer0_outputs(1677)) and (layer0_outputs(1683)));
    layer1_outputs(905) <= not(layer0_outputs(1904));
    layer1_outputs(906) <= not(layer0_outputs(1574)) or (layer0_outputs(1559));
    layer1_outputs(907) <= not((layer0_outputs(1464)) and (layer0_outputs(1434)));
    layer1_outputs(908) <= layer0_outputs(1695);
    layer1_outputs(909) <= layer0_outputs(1926);
    layer1_outputs(910) <= not((layer0_outputs(1905)) and (layer0_outputs(1578)));
    layer1_outputs(911) <= not((layer0_outputs(846)) and (layer0_outputs(2017)));
    layer1_outputs(912) <= '0';
    layer1_outputs(913) <= not(layer0_outputs(24));
    layer1_outputs(914) <= layer0_outputs(999);
    layer1_outputs(915) <= '1';
    layer1_outputs(916) <= not(layer0_outputs(2048)) or (layer0_outputs(1861));
    layer1_outputs(917) <= (layer0_outputs(2462)) or (layer0_outputs(2132));
    layer1_outputs(918) <= (layer0_outputs(1005)) and (layer0_outputs(780));
    layer1_outputs(919) <= not(layer0_outputs(1550));
    layer1_outputs(920) <= layer0_outputs(2060);
    layer1_outputs(921) <= (layer0_outputs(2535)) and not (layer0_outputs(1903));
    layer1_outputs(922) <= layer0_outputs(2199);
    layer1_outputs(923) <= not(layer0_outputs(1977));
    layer1_outputs(924) <= not((layer0_outputs(462)) and (layer0_outputs(1650)));
    layer1_outputs(925) <= not(layer0_outputs(1445));
    layer1_outputs(926) <= (layer0_outputs(2513)) and not (layer0_outputs(1878));
    layer1_outputs(927) <= not(layer0_outputs(1188)) or (layer0_outputs(2433));
    layer1_outputs(928) <= not((layer0_outputs(869)) and (layer0_outputs(352)));
    layer1_outputs(929) <= not((layer0_outputs(1245)) or (layer0_outputs(2346)));
    layer1_outputs(930) <= layer0_outputs(1125);
    layer1_outputs(931) <= '1';
    layer1_outputs(932) <= (layer0_outputs(1105)) and (layer0_outputs(952));
    layer1_outputs(933) <= (layer0_outputs(1387)) or (layer0_outputs(74));
    layer1_outputs(934) <= (layer0_outputs(768)) and not (layer0_outputs(35));
    layer1_outputs(935) <= not((layer0_outputs(197)) or (layer0_outputs(1936)));
    layer1_outputs(936) <= not(layer0_outputs(1387));
    layer1_outputs(937) <= (layer0_outputs(2019)) or (layer0_outputs(1597));
    layer1_outputs(938) <= (layer0_outputs(501)) and not (layer0_outputs(747));
    layer1_outputs(939) <= not(layer0_outputs(719));
    layer1_outputs(940) <= not((layer0_outputs(1551)) and (layer0_outputs(1100)));
    layer1_outputs(941) <= not((layer0_outputs(734)) and (layer0_outputs(2215)));
    layer1_outputs(942) <= not(layer0_outputs(238));
    layer1_outputs(943) <= (layer0_outputs(1992)) xor (layer0_outputs(1528));
    layer1_outputs(944) <= layer0_outputs(1698);
    layer1_outputs(945) <= not(layer0_outputs(981));
    layer1_outputs(946) <= layer0_outputs(620);
    layer1_outputs(947) <= (layer0_outputs(2200)) and not (layer0_outputs(951));
    layer1_outputs(948) <= layer0_outputs(1496);
    layer1_outputs(949) <= layer0_outputs(1821);
    layer1_outputs(950) <= (layer0_outputs(1198)) and (layer0_outputs(756));
    layer1_outputs(951) <= (layer0_outputs(732)) and (layer0_outputs(590));
    layer1_outputs(952) <= (layer0_outputs(2394)) and not (layer0_outputs(1918));
    layer1_outputs(953) <= (layer0_outputs(2065)) and not (layer0_outputs(65));
    layer1_outputs(954) <= not((layer0_outputs(1228)) or (layer0_outputs(907)));
    layer1_outputs(955) <= not((layer0_outputs(1561)) or (layer0_outputs(1469)));
    layer1_outputs(956) <= not(layer0_outputs(2047)) or (layer0_outputs(107));
    layer1_outputs(957) <= not(layer0_outputs(1211));
    layer1_outputs(958) <= not(layer0_outputs(2503));
    layer1_outputs(959) <= not(layer0_outputs(661)) or (layer0_outputs(1426));
    layer1_outputs(960) <= not(layer0_outputs(2193));
    layer1_outputs(961) <= not(layer0_outputs(1325)) or (layer0_outputs(2207));
    layer1_outputs(962) <= (layer0_outputs(1324)) or (layer0_outputs(2081));
    layer1_outputs(963) <= not((layer0_outputs(1652)) and (layer0_outputs(1617)));
    layer1_outputs(964) <= (layer0_outputs(2189)) and (layer0_outputs(1670));
    layer1_outputs(965) <= not(layer0_outputs(70));
    layer1_outputs(966) <= not(layer0_outputs(29));
    layer1_outputs(967) <= not(layer0_outputs(450)) or (layer0_outputs(905));
    layer1_outputs(968) <= not(layer0_outputs(783));
    layer1_outputs(969) <= not((layer0_outputs(2534)) or (layer0_outputs(726)));
    layer1_outputs(970) <= (layer0_outputs(2504)) or (layer0_outputs(2197));
    layer1_outputs(971) <= not(layer0_outputs(372));
    layer1_outputs(972) <= not(layer0_outputs(299));
    layer1_outputs(973) <= layer0_outputs(730);
    layer1_outputs(974) <= (layer0_outputs(2380)) and not (layer0_outputs(1087));
    layer1_outputs(975) <= (layer0_outputs(1608)) and (layer0_outputs(271));
    layer1_outputs(976) <= not(layer0_outputs(1492));
    layer1_outputs(977) <= not((layer0_outputs(1491)) or (layer0_outputs(341)));
    layer1_outputs(978) <= not((layer0_outputs(917)) or (layer0_outputs(1684)));
    layer1_outputs(979) <= (layer0_outputs(2326)) and (layer0_outputs(2497));
    layer1_outputs(980) <= layer0_outputs(1024);
    layer1_outputs(981) <= not(layer0_outputs(2272));
    layer1_outputs(982) <= not((layer0_outputs(36)) xor (layer0_outputs(2015)));
    layer1_outputs(983) <= layer0_outputs(2555);
    layer1_outputs(984) <= (layer0_outputs(1308)) and not (layer0_outputs(1610));
    layer1_outputs(985) <= not(layer0_outputs(1403));
    layer1_outputs(986) <= (layer0_outputs(1750)) or (layer0_outputs(634));
    layer1_outputs(987) <= (layer0_outputs(746)) or (layer0_outputs(60));
    layer1_outputs(988) <= layer0_outputs(719);
    layer1_outputs(989) <= not((layer0_outputs(293)) xor (layer0_outputs(2229)));
    layer1_outputs(990) <= not((layer0_outputs(441)) or (layer0_outputs(1922)));
    layer1_outputs(991) <= not(layer0_outputs(1317)) or (layer0_outputs(901));
    layer1_outputs(992) <= (layer0_outputs(2369)) or (layer0_outputs(2085));
    layer1_outputs(993) <= not(layer0_outputs(1651)) or (layer0_outputs(864));
    layer1_outputs(994) <= not(layer0_outputs(1646));
    layer1_outputs(995) <= (layer0_outputs(1456)) or (layer0_outputs(741));
    layer1_outputs(996) <= '1';
    layer1_outputs(997) <= layer0_outputs(1727);
    layer1_outputs(998) <= not((layer0_outputs(1026)) and (layer0_outputs(2544)));
    layer1_outputs(999) <= (layer0_outputs(2216)) and (layer0_outputs(273));
    layer1_outputs(1000) <= not(layer0_outputs(1075));
    layer1_outputs(1001) <= (layer0_outputs(1342)) and not (layer0_outputs(1020));
    layer1_outputs(1002) <= (layer0_outputs(1547)) or (layer0_outputs(517));
    layer1_outputs(1003) <= (layer0_outputs(1147)) and (layer0_outputs(601));
    layer1_outputs(1004) <= (layer0_outputs(2202)) and (layer0_outputs(1583));
    layer1_outputs(1005) <= not((layer0_outputs(1765)) or (layer0_outputs(135)));
    layer1_outputs(1006) <= not(layer0_outputs(1791));
    layer1_outputs(1007) <= '1';
    layer1_outputs(1008) <= layer0_outputs(2125);
    layer1_outputs(1009) <= not(layer0_outputs(713));
    layer1_outputs(1010) <= not(layer0_outputs(2426));
    layer1_outputs(1011) <= not(layer0_outputs(612));
    layer1_outputs(1012) <= (layer0_outputs(280)) and not (layer0_outputs(1230));
    layer1_outputs(1013) <= not((layer0_outputs(2123)) or (layer0_outputs(1330)));
    layer1_outputs(1014) <= (layer0_outputs(296)) and not (layer0_outputs(2310));
    layer1_outputs(1015) <= layer0_outputs(163);
    layer1_outputs(1016) <= '1';
    layer1_outputs(1017) <= not(layer0_outputs(964));
    layer1_outputs(1018) <= not(layer0_outputs(1818));
    layer1_outputs(1019) <= (layer0_outputs(118)) and (layer0_outputs(1309));
    layer1_outputs(1020) <= layer0_outputs(345);
    layer1_outputs(1021) <= not(layer0_outputs(1858));
    layer1_outputs(1022) <= not((layer0_outputs(1039)) and (layer0_outputs(1343)));
    layer1_outputs(1023) <= not((layer0_outputs(578)) xor (layer0_outputs(2126)));
    layer1_outputs(1024) <= not((layer0_outputs(113)) or (layer0_outputs(494)));
    layer1_outputs(1025) <= (layer0_outputs(1406)) and not (layer0_outputs(2161));
    layer1_outputs(1026) <= (layer0_outputs(909)) and (layer0_outputs(2164));
    layer1_outputs(1027) <= (layer0_outputs(885)) and not (layer0_outputs(1337));
    layer1_outputs(1028) <= (layer0_outputs(1419)) and not (layer0_outputs(2028));
    layer1_outputs(1029) <= not(layer0_outputs(2097));
    layer1_outputs(1030) <= layer0_outputs(1890);
    layer1_outputs(1031) <= (layer0_outputs(1420)) and (layer0_outputs(354));
    layer1_outputs(1032) <= not(layer0_outputs(520));
    layer1_outputs(1033) <= not(layer0_outputs(193));
    layer1_outputs(1034) <= (layer0_outputs(533)) and not (layer0_outputs(1840));
    layer1_outputs(1035) <= layer0_outputs(541);
    layer1_outputs(1036) <= (layer0_outputs(2205)) and (layer0_outputs(382));
    layer1_outputs(1037) <= '1';
    layer1_outputs(1038) <= not(layer0_outputs(1367));
    layer1_outputs(1039) <= not((layer0_outputs(417)) and (layer0_outputs(2058)));
    layer1_outputs(1040) <= not(layer0_outputs(2112));
    layer1_outputs(1041) <= not(layer0_outputs(205)) or (layer0_outputs(402));
    layer1_outputs(1042) <= not(layer0_outputs(2310)) or (layer0_outputs(342));
    layer1_outputs(1043) <= (layer0_outputs(809)) and (layer0_outputs(2226));
    layer1_outputs(1044) <= (layer0_outputs(2352)) and (layer0_outputs(2003));
    layer1_outputs(1045) <= not(layer0_outputs(2043));
    layer1_outputs(1046) <= not(layer0_outputs(886)) or (layer0_outputs(1690));
    layer1_outputs(1047) <= not(layer0_outputs(1305));
    layer1_outputs(1048) <= not((layer0_outputs(1576)) and (layer0_outputs(424)));
    layer1_outputs(1049) <= layer0_outputs(1632);
    layer1_outputs(1050) <= not(layer0_outputs(2188));
    layer1_outputs(1051) <= not(layer0_outputs(966));
    layer1_outputs(1052) <= (layer0_outputs(106)) and not (layer0_outputs(35));
    layer1_outputs(1053) <= layer0_outputs(454);
    layer1_outputs(1054) <= (layer0_outputs(438)) and (layer0_outputs(941));
    layer1_outputs(1055) <= not((layer0_outputs(2502)) or (layer0_outputs(965)));
    layer1_outputs(1056) <= layer0_outputs(939);
    layer1_outputs(1057) <= '1';
    layer1_outputs(1058) <= not(layer0_outputs(324)) or (layer0_outputs(1366));
    layer1_outputs(1059) <= not(layer0_outputs(2133)) or (layer0_outputs(1588));
    layer1_outputs(1060) <= not(layer0_outputs(1853)) or (layer0_outputs(1657));
    layer1_outputs(1061) <= (layer0_outputs(1277)) and not (layer0_outputs(2438));
    layer1_outputs(1062) <= not(layer0_outputs(2110));
    layer1_outputs(1063) <= (layer0_outputs(1803)) and (layer0_outputs(585));
    layer1_outputs(1064) <= '0';
    layer1_outputs(1065) <= not((layer0_outputs(1720)) and (layer0_outputs(472)));
    layer1_outputs(1066) <= not(layer0_outputs(1123));
    layer1_outputs(1067) <= not((layer0_outputs(728)) or (layer0_outputs(160)));
    layer1_outputs(1068) <= not((layer0_outputs(1979)) and (layer0_outputs(326)));
    layer1_outputs(1069) <= not((layer0_outputs(2236)) and (layer0_outputs(310)));
    layer1_outputs(1070) <= layer0_outputs(950);
    layer1_outputs(1071) <= not((layer0_outputs(575)) or (layer0_outputs(1183)));
    layer1_outputs(1072) <= not(layer0_outputs(683));
    layer1_outputs(1073) <= (layer0_outputs(2198)) or (layer0_outputs(1680));
    layer1_outputs(1074) <= (layer0_outputs(1560)) and (layer0_outputs(360));
    layer1_outputs(1075) <= not((layer0_outputs(141)) xor (layer0_outputs(1515)));
    layer1_outputs(1076) <= (layer0_outputs(654)) and not (layer0_outputs(1766));
    layer1_outputs(1077) <= not((layer0_outputs(1137)) or (layer0_outputs(1914)));
    layer1_outputs(1078) <= not(layer0_outputs(373));
    layer1_outputs(1079) <= layer0_outputs(710);
    layer1_outputs(1080) <= not(layer0_outputs(478));
    layer1_outputs(1081) <= not(layer0_outputs(2433));
    layer1_outputs(1082) <= not((layer0_outputs(2414)) and (layer0_outputs(716)));
    layer1_outputs(1083) <= not(layer0_outputs(2103));
    layer1_outputs(1084) <= not(layer0_outputs(2547));
    layer1_outputs(1085) <= not(layer0_outputs(1011));
    layer1_outputs(1086) <= (layer0_outputs(1471)) and not (layer0_outputs(801));
    layer1_outputs(1087) <= layer0_outputs(1431);
    layer1_outputs(1088) <= layer0_outputs(1021);
    layer1_outputs(1089) <= not(layer0_outputs(1149));
    layer1_outputs(1090) <= not((layer0_outputs(1568)) or (layer0_outputs(2262)));
    layer1_outputs(1091) <= '1';
    layer1_outputs(1092) <= not(layer0_outputs(1960)) or (layer0_outputs(834));
    layer1_outputs(1093) <= not(layer0_outputs(2553)) or (layer0_outputs(77));
    layer1_outputs(1094) <= not((layer0_outputs(2445)) or (layer0_outputs(335)));
    layer1_outputs(1095) <= not((layer0_outputs(2239)) or (layer0_outputs(748)));
    layer1_outputs(1096) <= not(layer0_outputs(2260));
    layer1_outputs(1097) <= (layer0_outputs(2317)) and not (layer0_outputs(2542));
    layer1_outputs(1098) <= not(layer0_outputs(1461));
    layer1_outputs(1099) <= not(layer0_outputs(161));
    layer1_outputs(1100) <= not(layer0_outputs(461)) or (layer0_outputs(1800));
    layer1_outputs(1101) <= (layer0_outputs(938)) and not (layer0_outputs(805));
    layer1_outputs(1102) <= (layer0_outputs(595)) and (layer0_outputs(120));
    layer1_outputs(1103) <= (layer0_outputs(249)) and (layer0_outputs(1710));
    layer1_outputs(1104) <= not(layer0_outputs(1922));
    layer1_outputs(1105) <= not((layer0_outputs(1958)) or (layer0_outputs(1215)));
    layer1_outputs(1106) <= not(layer0_outputs(843)) or (layer0_outputs(401));
    layer1_outputs(1107) <= not(layer0_outputs(1339));
    layer1_outputs(1108) <= not(layer0_outputs(1749));
    layer1_outputs(1109) <= layer0_outputs(1206);
    layer1_outputs(1110) <= not(layer0_outputs(1925));
    layer1_outputs(1111) <= (layer0_outputs(707)) and not (layer0_outputs(1201));
    layer1_outputs(1112) <= not(layer0_outputs(2479));
    layer1_outputs(1113) <= (layer0_outputs(1538)) and not (layer0_outputs(755));
    layer1_outputs(1114) <= not(layer0_outputs(1199)) or (layer0_outputs(531));
    layer1_outputs(1115) <= layer0_outputs(2334);
    layer1_outputs(1116) <= layer0_outputs(2234);
    layer1_outputs(1117) <= not((layer0_outputs(875)) xor (layer0_outputs(1978)));
    layer1_outputs(1118) <= not(layer0_outputs(2265)) or (layer0_outputs(2393));
    layer1_outputs(1119) <= not(layer0_outputs(521)) or (layer0_outputs(2208));
    layer1_outputs(1120) <= not(layer0_outputs(923));
    layer1_outputs(1121) <= (layer0_outputs(31)) and not (layer0_outputs(994));
    layer1_outputs(1122) <= not(layer0_outputs(185)) or (layer0_outputs(642));
    layer1_outputs(1123) <= not(layer0_outputs(2395)) or (layer0_outputs(353));
    layer1_outputs(1124) <= not(layer0_outputs(732)) or (layer0_outputs(536));
    layer1_outputs(1125) <= layer0_outputs(686);
    layer1_outputs(1126) <= (layer0_outputs(381)) xor (layer0_outputs(662));
    layer1_outputs(1127) <= not((layer0_outputs(1200)) and (layer0_outputs(27)));
    layer1_outputs(1128) <= (layer0_outputs(2138)) and (layer0_outputs(872));
    layer1_outputs(1129) <= (layer0_outputs(225)) and not (layer0_outputs(1241));
    layer1_outputs(1130) <= '0';
    layer1_outputs(1131) <= not((layer0_outputs(802)) or (layer0_outputs(1084)));
    layer1_outputs(1132) <= not(layer0_outputs(1416));
    layer1_outputs(1133) <= not((layer0_outputs(1742)) and (layer0_outputs(447)));
    layer1_outputs(1134) <= (layer0_outputs(142)) xor (layer0_outputs(221));
    layer1_outputs(1135) <= (layer0_outputs(175)) and (layer0_outputs(1078));
    layer1_outputs(1136) <= not(layer0_outputs(2209)) or (layer0_outputs(1549));
    layer1_outputs(1137) <= not(layer0_outputs(118)) or (layer0_outputs(203));
    layer1_outputs(1138) <= not(layer0_outputs(820));
    layer1_outputs(1139) <= not(layer0_outputs(1610));
    layer1_outputs(1140) <= not(layer0_outputs(789));
    layer1_outputs(1141) <= not(layer0_outputs(1516));
    layer1_outputs(1142) <= layer0_outputs(738);
    layer1_outputs(1143) <= not((layer0_outputs(2392)) or (layer0_outputs(2227)));
    layer1_outputs(1144) <= '1';
    layer1_outputs(1145) <= not(layer0_outputs(952));
    layer1_outputs(1146) <= not(layer0_outputs(180));
    layer1_outputs(1147) <= not(layer0_outputs(879));
    layer1_outputs(1148) <= (layer0_outputs(140)) and not (layer0_outputs(2383));
    layer1_outputs(1149) <= '0';
    layer1_outputs(1150) <= (layer0_outputs(85)) or (layer0_outputs(191));
    layer1_outputs(1151) <= layer0_outputs(546);
    layer1_outputs(1152) <= (layer0_outputs(1352)) and not (layer0_outputs(500));
    layer1_outputs(1153) <= (layer0_outputs(775)) and (layer0_outputs(1874));
    layer1_outputs(1154) <= not(layer0_outputs(1755));
    layer1_outputs(1155) <= not(layer0_outputs(1672));
    layer1_outputs(1156) <= layer0_outputs(2267);
    layer1_outputs(1157) <= not(layer0_outputs(261));
    layer1_outputs(1158) <= layer0_outputs(1974);
    layer1_outputs(1159) <= not(layer0_outputs(455));
    layer1_outputs(1160) <= (layer0_outputs(1186)) and not (layer0_outputs(1912));
    layer1_outputs(1161) <= not((layer0_outputs(1699)) xor (layer0_outputs(803)));
    layer1_outputs(1162) <= '0';
    layer1_outputs(1163) <= layer0_outputs(2431);
    layer1_outputs(1164) <= not((layer0_outputs(1609)) or (layer0_outputs(181)));
    layer1_outputs(1165) <= (layer0_outputs(2383)) and not (layer0_outputs(1951));
    layer1_outputs(1166) <= (layer0_outputs(618)) and (layer0_outputs(2203));
    layer1_outputs(1167) <= not(layer0_outputs(695)) or (layer0_outputs(1467));
    layer1_outputs(1168) <= (layer0_outputs(1643)) or (layer0_outputs(1896));
    layer1_outputs(1169) <= not(layer0_outputs(1404));
    layer1_outputs(1170) <= not(layer0_outputs(1643));
    layer1_outputs(1171) <= (layer0_outputs(2259)) and (layer0_outputs(2484));
    layer1_outputs(1172) <= (layer0_outputs(1321)) and not (layer0_outputs(911));
    layer1_outputs(1173) <= not(layer0_outputs(1575)) or (layer0_outputs(1751));
    layer1_outputs(1174) <= layer0_outputs(557);
    layer1_outputs(1175) <= not(layer0_outputs(1037)) or (layer0_outputs(401));
    layer1_outputs(1176) <= not(layer0_outputs(773));
    layer1_outputs(1177) <= not(layer0_outputs(645)) or (layer0_outputs(54));
    layer1_outputs(1178) <= layer0_outputs(816);
    layer1_outputs(1179) <= (layer0_outputs(1225)) and not (layer0_outputs(1096));
    layer1_outputs(1180) <= (layer0_outputs(2202)) and (layer0_outputs(2356));
    layer1_outputs(1181) <= (layer0_outputs(1363)) and not (layer0_outputs(1517));
    layer1_outputs(1182) <= not(layer0_outputs(2035));
    layer1_outputs(1183) <= layer0_outputs(97);
    layer1_outputs(1184) <= not(layer0_outputs(2378)) or (layer0_outputs(124));
    layer1_outputs(1185) <= not((layer0_outputs(1370)) or (layer0_outputs(1924)));
    layer1_outputs(1186) <= layer0_outputs(671);
    layer1_outputs(1187) <= layer0_outputs(2280);
    layer1_outputs(1188) <= not(layer0_outputs(1380));
    layer1_outputs(1189) <= not((layer0_outputs(1270)) xor (layer0_outputs(629)));
    layer1_outputs(1190) <= layer0_outputs(2022);
    layer1_outputs(1191) <= not((layer0_outputs(1424)) or (layer0_outputs(1282)));
    layer1_outputs(1192) <= not(layer0_outputs(846)) or (layer0_outputs(950));
    layer1_outputs(1193) <= not(layer0_outputs(99));
    layer1_outputs(1194) <= (layer0_outputs(2473)) xor (layer0_outputs(2530));
    layer1_outputs(1195) <= not(layer0_outputs(569));
    layer1_outputs(1196) <= not(layer0_outputs(2128)) or (layer0_outputs(2105));
    layer1_outputs(1197) <= (layer0_outputs(713)) and not (layer0_outputs(2027));
    layer1_outputs(1198) <= layer0_outputs(274);
    layer1_outputs(1199) <= not((layer0_outputs(2055)) or (layer0_outputs(1471)));
    layer1_outputs(1200) <= not(layer0_outputs(1759)) or (layer0_outputs(1507));
    layer1_outputs(1201) <= not(layer0_outputs(1348));
    layer1_outputs(1202) <= layer0_outputs(1290);
    layer1_outputs(1203) <= layer0_outputs(165);
    layer1_outputs(1204) <= (layer0_outputs(328)) and not (layer0_outputs(608));
    layer1_outputs(1205) <= (layer0_outputs(1850)) and (layer0_outputs(2222));
    layer1_outputs(1206) <= (layer0_outputs(1453)) and (layer0_outputs(545));
    layer1_outputs(1207) <= not(layer0_outputs(1865));
    layer1_outputs(1208) <= layer0_outputs(753);
    layer1_outputs(1209) <= layer0_outputs(1935);
    layer1_outputs(1210) <= not((layer0_outputs(420)) or (layer0_outputs(102)));
    layer1_outputs(1211) <= (layer0_outputs(1624)) and not (layer0_outputs(1178));
    layer1_outputs(1212) <= (layer0_outputs(995)) and not (layer0_outputs(377));
    layer1_outputs(1213) <= not((layer0_outputs(386)) xor (layer0_outputs(1346)));
    layer1_outputs(1214) <= layer0_outputs(2400);
    layer1_outputs(1215) <= '0';
    layer1_outputs(1216) <= layer0_outputs(2527);
    layer1_outputs(1217) <= not(layer0_outputs(2101));
    layer1_outputs(1218) <= layer0_outputs(1747);
    layer1_outputs(1219) <= not((layer0_outputs(782)) or (layer0_outputs(1854)));
    layer1_outputs(1220) <= (layer0_outputs(599)) and not (layer0_outputs(1463));
    layer1_outputs(1221) <= not((layer0_outputs(910)) or (layer0_outputs(1418)));
    layer1_outputs(1222) <= (layer0_outputs(1242)) and not (layer0_outputs(2155));
    layer1_outputs(1223) <= layer0_outputs(881);
    layer1_outputs(1224) <= (layer0_outputs(538)) and (layer0_outputs(1676));
    layer1_outputs(1225) <= not(layer0_outputs(2020));
    layer1_outputs(1226) <= not(layer0_outputs(2169));
    layer1_outputs(1227) <= layer0_outputs(2330);
    layer1_outputs(1228) <= (layer0_outputs(332)) xor (layer0_outputs(2409));
    layer1_outputs(1229) <= layer0_outputs(2183);
    layer1_outputs(1230) <= layer0_outputs(656);
    layer1_outputs(1231) <= not((layer0_outputs(1897)) and (layer0_outputs(1886)));
    layer1_outputs(1232) <= not((layer0_outputs(746)) or (layer0_outputs(2412)));
    layer1_outputs(1233) <= not((layer0_outputs(1290)) and (layer0_outputs(1603)));
    layer1_outputs(1234) <= not(layer0_outputs(2374)) or (layer0_outputs(230));
    layer1_outputs(1235) <= not(layer0_outputs(2231));
    layer1_outputs(1236) <= not(layer0_outputs(1730)) or (layer0_outputs(816));
    layer1_outputs(1237) <= (layer0_outputs(373)) and (layer0_outputs(2045));
    layer1_outputs(1238) <= layer0_outputs(2053);
    layer1_outputs(1239) <= layer0_outputs(2413);
    layer1_outputs(1240) <= layer0_outputs(2349);
    layer1_outputs(1241) <= (layer0_outputs(130)) and not (layer0_outputs(2482));
    layer1_outputs(1242) <= layer0_outputs(1826);
    layer1_outputs(1243) <= (layer0_outputs(408)) and (layer0_outputs(2273));
    layer1_outputs(1244) <= not(layer0_outputs(1964));
    layer1_outputs(1245) <= layer0_outputs(497);
    layer1_outputs(1246) <= layer0_outputs(2356);
    layer1_outputs(1247) <= not(layer0_outputs(986)) or (layer0_outputs(269));
    layer1_outputs(1248) <= not((layer0_outputs(1668)) xor (layer0_outputs(178)));
    layer1_outputs(1249) <= '1';
    layer1_outputs(1250) <= '1';
    layer1_outputs(1251) <= (layer0_outputs(2464)) or (layer0_outputs(1816));
    layer1_outputs(1252) <= not(layer0_outputs(513)) or (layer0_outputs(1191));
    layer1_outputs(1253) <= (layer0_outputs(232)) and not (layer0_outputs(1483));
    layer1_outputs(1254) <= (layer0_outputs(927)) or (layer0_outputs(1533));
    layer1_outputs(1255) <= not(layer0_outputs(1833));
    layer1_outputs(1256) <= not((layer0_outputs(624)) and (layer0_outputs(1403)));
    layer1_outputs(1257) <= not(layer0_outputs(2005)) or (layer0_outputs(707));
    layer1_outputs(1258) <= not(layer0_outputs(332));
    layer1_outputs(1259) <= (layer0_outputs(2493)) and not (layer0_outputs(1015));
    layer1_outputs(1260) <= not(layer0_outputs(28));
    layer1_outputs(1261) <= '1';
    layer1_outputs(1262) <= layer0_outputs(1412);
    layer1_outputs(1263) <= not(layer0_outputs(914)) or (layer0_outputs(2274));
    layer1_outputs(1264) <= layer0_outputs(971);
    layer1_outputs(1265) <= (layer0_outputs(671)) xor (layer0_outputs(526));
    layer1_outputs(1266) <= (layer0_outputs(1277)) and not (layer0_outputs(407));
    layer1_outputs(1267) <= not(layer0_outputs(896)) or (layer0_outputs(2381));
    layer1_outputs(1268) <= (layer0_outputs(2376)) or (layer0_outputs(2048));
    layer1_outputs(1269) <= not(layer0_outputs(945));
    layer1_outputs(1270) <= (layer0_outputs(1126)) and (layer0_outputs(868));
    layer1_outputs(1271) <= layer0_outputs(219);
    layer1_outputs(1272) <= not(layer0_outputs(2181));
    layer1_outputs(1273) <= (layer0_outputs(1004)) and not (layer0_outputs(237));
    layer1_outputs(1274) <= (layer0_outputs(2499)) xor (layer0_outputs(1349));
    layer1_outputs(1275) <= layer0_outputs(2099);
    layer1_outputs(1276) <= '1';
    layer1_outputs(1277) <= not(layer0_outputs(645));
    layer1_outputs(1278) <= not((layer0_outputs(1184)) or (layer0_outputs(2170)));
    layer1_outputs(1279) <= not((layer0_outputs(914)) or (layer0_outputs(1489)));
    layer1_outputs(1280) <= (layer0_outputs(825)) and (layer0_outputs(1063));
    layer1_outputs(1281) <= (layer0_outputs(1736)) and not (layer0_outputs(1685));
    layer1_outputs(1282) <= layer0_outputs(67);
    layer1_outputs(1283) <= '1';
    layer1_outputs(1284) <= '1';
    layer1_outputs(1285) <= not(layer0_outputs(1764));
    layer1_outputs(1286) <= not(layer0_outputs(1421));
    layer1_outputs(1287) <= not((layer0_outputs(9)) and (layer0_outputs(80)));
    layer1_outputs(1288) <= not((layer0_outputs(966)) and (layer0_outputs(297)));
    layer1_outputs(1289) <= (layer0_outputs(2505)) or (layer0_outputs(1899));
    layer1_outputs(1290) <= '0';
    layer1_outputs(1291) <= not(layer0_outputs(1457));
    layer1_outputs(1292) <= not(layer0_outputs(1971));
    layer1_outputs(1293) <= layer0_outputs(398);
    layer1_outputs(1294) <= (layer0_outputs(312)) and (layer0_outputs(1009));
    layer1_outputs(1295) <= (layer0_outputs(1288)) and not (layer0_outputs(572));
    layer1_outputs(1296) <= not((layer0_outputs(1563)) or (layer0_outputs(2295)));
    layer1_outputs(1297) <= not((layer0_outputs(1668)) and (layer0_outputs(1271)));
    layer1_outputs(1298) <= not(layer0_outputs(1181));
    layer1_outputs(1299) <= not((layer0_outputs(1516)) or (layer0_outputs(1810)));
    layer1_outputs(1300) <= (layer0_outputs(599)) and not (layer0_outputs(1729));
    layer1_outputs(1301) <= not(layer0_outputs(1231)) or (layer0_outputs(988));
    layer1_outputs(1302) <= not(layer0_outputs(1269)) or (layer0_outputs(1117));
    layer1_outputs(1303) <= (layer0_outputs(1535)) and not (layer0_outputs(1429));
    layer1_outputs(1304) <= '0';
    layer1_outputs(1305) <= (layer0_outputs(683)) or (layer0_outputs(2467));
    layer1_outputs(1306) <= layer0_outputs(1463);
    layer1_outputs(1307) <= (layer0_outputs(1350)) and not (layer0_outputs(2447));
    layer1_outputs(1308) <= not((layer0_outputs(1637)) or (layer0_outputs(2362)));
    layer1_outputs(1309) <= (layer0_outputs(1804)) and not (layer0_outputs(692));
    layer1_outputs(1310) <= not((layer0_outputs(2501)) and (layer0_outputs(1963)));
    layer1_outputs(1311) <= '1';
    layer1_outputs(1312) <= not(layer0_outputs(839));
    layer1_outputs(1313) <= not(layer0_outputs(53));
    layer1_outputs(1314) <= '0';
    layer1_outputs(1315) <= not(layer0_outputs(1372));
    layer1_outputs(1316) <= not(layer0_outputs(299)) or (layer0_outputs(551));
    layer1_outputs(1317) <= layer0_outputs(920);
    layer1_outputs(1318) <= not(layer0_outputs(2153));
    layer1_outputs(1319) <= layer0_outputs(2493);
    layer1_outputs(1320) <= (layer0_outputs(492)) or (layer0_outputs(1787));
    layer1_outputs(1321) <= not(layer0_outputs(1082));
    layer1_outputs(1322) <= not((layer0_outputs(198)) or (layer0_outputs(1851)));
    layer1_outputs(1323) <= (layer0_outputs(1240)) and (layer0_outputs(1790));
    layer1_outputs(1324) <= layer0_outputs(2514);
    layer1_outputs(1325) <= layer0_outputs(1586);
    layer1_outputs(1326) <= layer0_outputs(739);
    layer1_outputs(1327) <= not(layer0_outputs(632)) or (layer0_outputs(2046));
    layer1_outputs(1328) <= layer0_outputs(900);
    layer1_outputs(1329) <= (layer0_outputs(1168)) and not (layer0_outputs(348));
    layer1_outputs(1330) <= not(layer0_outputs(2423)) or (layer0_outputs(604));
    layer1_outputs(1331) <= not((layer0_outputs(1307)) xor (layer0_outputs(156)));
    layer1_outputs(1332) <= (layer0_outputs(629)) and not (layer0_outputs(12));
    layer1_outputs(1333) <= not(layer0_outputs(350));
    layer1_outputs(1334) <= '1';
    layer1_outputs(1335) <= (layer0_outputs(1114)) and not (layer0_outputs(616));
    layer1_outputs(1336) <= layer0_outputs(1318);
    layer1_outputs(1337) <= (layer0_outputs(916)) or (layer0_outputs(1200));
    layer1_outputs(1338) <= '0';
    layer1_outputs(1339) <= layer0_outputs(642);
    layer1_outputs(1340) <= layer0_outputs(45);
    layer1_outputs(1341) <= not(layer0_outputs(2042));
    layer1_outputs(1342) <= not((layer0_outputs(580)) and (layer0_outputs(1607)));
    layer1_outputs(1343) <= not(layer0_outputs(1739)) or (layer0_outputs(2167));
    layer1_outputs(1344) <= not(layer0_outputs(234));
    layer1_outputs(1345) <= layer0_outputs(1740);
    layer1_outputs(1346) <= not(layer0_outputs(1972));
    layer1_outputs(1347) <= layer0_outputs(1596);
    layer1_outputs(1348) <= not(layer0_outputs(218));
    layer1_outputs(1349) <= not(layer0_outputs(2365));
    layer1_outputs(1350) <= not((layer0_outputs(1571)) and (layer0_outputs(1676)));
    layer1_outputs(1351) <= not(layer0_outputs(522));
    layer1_outputs(1352) <= layer0_outputs(993);
    layer1_outputs(1353) <= not((layer0_outputs(2522)) and (layer0_outputs(573)));
    layer1_outputs(1354) <= not((layer0_outputs(1694)) and (layer0_outputs(745)));
    layer1_outputs(1355) <= not(layer0_outputs(775));
    layer1_outputs(1356) <= not(layer0_outputs(1145));
    layer1_outputs(1357) <= not((layer0_outputs(1688)) or (layer0_outputs(1968)));
    layer1_outputs(1358) <= layer0_outputs(1658);
    layer1_outputs(1359) <= not((layer0_outputs(1130)) and (layer0_outputs(1990)));
    layer1_outputs(1360) <= layer0_outputs(187);
    layer1_outputs(1361) <= not((layer0_outputs(570)) or (layer0_outputs(465)));
    layer1_outputs(1362) <= not(layer0_outputs(1450));
    layer1_outputs(1363) <= (layer0_outputs(115)) and not (layer0_outputs(1507));
    layer1_outputs(1364) <= not((layer0_outputs(1928)) xor (layer0_outputs(110)));
    layer1_outputs(1365) <= (layer0_outputs(1294)) or (layer0_outputs(1889));
    layer1_outputs(1366) <= '0';
    layer1_outputs(1367) <= not(layer0_outputs(525));
    layer1_outputs(1368) <= (layer0_outputs(2474)) xor (layer0_outputs(1604));
    layer1_outputs(1369) <= not(layer0_outputs(1007));
    layer1_outputs(1370) <= layer0_outputs(669);
    layer1_outputs(1371) <= not(layer0_outputs(48));
    layer1_outputs(1372) <= (layer0_outputs(1472)) or (layer0_outputs(1274));
    layer1_outputs(1373) <= layer0_outputs(209);
    layer1_outputs(1374) <= (layer0_outputs(1701)) and not (layer0_outputs(1370));
    layer1_outputs(1375) <= not(layer0_outputs(892)) or (layer0_outputs(298));
    layer1_outputs(1376) <= (layer0_outputs(431)) and not (layer0_outputs(1474));
    layer1_outputs(1377) <= layer0_outputs(2041);
    layer1_outputs(1378) <= not(layer0_outputs(1219)) or (layer0_outputs(884));
    layer1_outputs(1379) <= layer0_outputs(1687);
    layer1_outputs(1380) <= not(layer0_outputs(2113));
    layer1_outputs(1381) <= not(layer0_outputs(1077));
    layer1_outputs(1382) <= not((layer0_outputs(505)) or (layer0_outputs(882)));
    layer1_outputs(1383) <= not((layer0_outputs(1392)) or (layer0_outputs(1410)));
    layer1_outputs(1384) <= layer0_outputs(1345);
    layer1_outputs(1385) <= (layer0_outputs(1473)) and not (layer0_outputs(516));
    layer1_outputs(1386) <= (layer0_outputs(654)) or (layer0_outputs(2318));
    layer1_outputs(1387) <= (layer0_outputs(1322)) and not (layer0_outputs(344));
    layer1_outputs(1388) <= layer0_outputs(1701);
    layer1_outputs(1389) <= layer0_outputs(2291);
    layer1_outputs(1390) <= not((layer0_outputs(2241)) and (layer0_outputs(2525)));
    layer1_outputs(1391) <= not(layer0_outputs(1572)) or (layer0_outputs(2079));
    layer1_outputs(1392) <= not(layer0_outputs(606));
    layer1_outputs(1393) <= (layer0_outputs(1244)) and (layer0_outputs(2373));
    layer1_outputs(1394) <= (layer0_outputs(1043)) xor (layer0_outputs(272));
    layer1_outputs(1395) <= not(layer0_outputs(982)) or (layer0_outputs(2189));
    layer1_outputs(1396) <= not(layer0_outputs(2329));
    layer1_outputs(1397) <= not(layer0_outputs(1611)) or (layer0_outputs(1000));
    layer1_outputs(1398) <= (layer0_outputs(303)) and not (layer0_outputs(83));
    layer1_outputs(1399) <= not((layer0_outputs(602)) xor (layer0_outputs(336)));
    layer1_outputs(1400) <= not((layer0_outputs(422)) or (layer0_outputs(961)));
    layer1_outputs(1401) <= layer0_outputs(172);
    layer1_outputs(1402) <= '0';
    layer1_outputs(1403) <= not(layer0_outputs(564));
    layer1_outputs(1404) <= layer0_outputs(1653);
    layer1_outputs(1405) <= not(layer0_outputs(2254));
    layer1_outputs(1406) <= not((layer0_outputs(1418)) or (layer0_outputs(2311)));
    layer1_outputs(1407) <= (layer0_outputs(2292)) and not (layer0_outputs(199));
    layer1_outputs(1408) <= layer0_outputs(539);
    layer1_outputs(1409) <= layer0_outputs(1466);
    layer1_outputs(1410) <= (layer0_outputs(1705)) or (layer0_outputs(1506));
    layer1_outputs(1411) <= not(layer0_outputs(686)) or (layer0_outputs(1276));
    layer1_outputs(1412) <= not(layer0_outputs(2186));
    layer1_outputs(1413) <= not(layer0_outputs(1679));
    layer1_outputs(1414) <= layer0_outputs(921);
    layer1_outputs(1415) <= (layer0_outputs(190)) and (layer0_outputs(1598));
    layer1_outputs(1416) <= not((layer0_outputs(669)) and (layer0_outputs(468)));
    layer1_outputs(1417) <= layer0_outputs(2529);
    layer1_outputs(1418) <= not(layer0_outputs(1123));
    layer1_outputs(1419) <= layer0_outputs(1485);
    layer1_outputs(1420) <= (layer0_outputs(1830)) and not (layer0_outputs(2227));
    layer1_outputs(1421) <= (layer0_outputs(1797)) and (layer0_outputs(1108));
    layer1_outputs(1422) <= (layer0_outputs(943)) and (layer0_outputs(2554));
    layer1_outputs(1423) <= layer0_outputs(1708);
    layer1_outputs(1424) <= layer0_outputs(636);
    layer1_outputs(1425) <= not(layer0_outputs(1176)) or (layer0_outputs(1626));
    layer1_outputs(1426) <= not((layer0_outputs(553)) and (layer0_outputs(2367)));
    layer1_outputs(1427) <= (layer0_outputs(1557)) and not (layer0_outputs(1545));
    layer1_outputs(1428) <= not(layer0_outputs(1034)) or (layer0_outputs(706));
    layer1_outputs(1429) <= not(layer0_outputs(2260)) or (layer0_outputs(10));
    layer1_outputs(1430) <= not((layer0_outputs(1918)) or (layer0_outputs(245)));
    layer1_outputs(1431) <= not(layer0_outputs(470));
    layer1_outputs(1432) <= not((layer0_outputs(817)) or (layer0_outputs(1007)));
    layer1_outputs(1433) <= (layer0_outputs(222)) or (layer0_outputs(635));
    layer1_outputs(1434) <= not((layer0_outputs(1012)) or (layer0_outputs(1405)));
    layer1_outputs(1435) <= not(layer0_outputs(1448));
    layer1_outputs(1436) <= not(layer0_outputs(584));
    layer1_outputs(1437) <= layer0_outputs(970);
    layer1_outputs(1438) <= (layer0_outputs(2308)) and (layer0_outputs(1425));
    layer1_outputs(1439) <= not(layer0_outputs(1189)) or (layer0_outputs(795));
    layer1_outputs(1440) <= not(layer0_outputs(2291)) or (layer0_outputs(189));
    layer1_outputs(1441) <= not(layer0_outputs(2265)) or (layer0_outputs(776));
    layer1_outputs(1442) <= '0';
    layer1_outputs(1443) <= layer0_outputs(710);
    layer1_outputs(1444) <= not(layer0_outputs(2010));
    layer1_outputs(1445) <= not(layer0_outputs(562)) or (layer0_outputs(1221));
    layer1_outputs(1446) <= '0';
    layer1_outputs(1447) <= (layer0_outputs(1249)) or (layer0_outputs(858));
    layer1_outputs(1448) <= not(layer0_outputs(320)) or (layer0_outputs(554));
    layer1_outputs(1449) <= not(layer0_outputs(2162));
    layer1_outputs(1450) <= not(layer0_outputs(1139));
    layer1_outputs(1451) <= (layer0_outputs(457)) or (layer0_outputs(2445));
    layer1_outputs(1452) <= not(layer0_outputs(2069)) or (layer0_outputs(1990));
    layer1_outputs(1453) <= not(layer0_outputs(1469)) or (layer0_outputs(302));
    layer1_outputs(1454) <= '0';
    layer1_outputs(1455) <= not(layer0_outputs(1215)) or (layer0_outputs(1965));
    layer1_outputs(1456) <= not((layer0_outputs(147)) and (layer0_outputs(953)));
    layer1_outputs(1457) <= not(layer0_outputs(1462));
    layer1_outputs(1458) <= not(layer0_outputs(2481)) or (layer0_outputs(2441));
    layer1_outputs(1459) <= (layer0_outputs(1825)) and not (layer0_outputs(1526));
    layer1_outputs(1460) <= not(layer0_outputs(1525));
    layer1_outputs(1461) <= not(layer0_outputs(1486));
    layer1_outputs(1462) <= not(layer0_outputs(2018)) or (layer0_outputs(1125));
    layer1_outputs(1463) <= '0';
    layer1_outputs(1464) <= layer0_outputs(983);
    layer1_outputs(1465) <= (layer0_outputs(237)) and not (layer0_outputs(1388));
    layer1_outputs(1466) <= (layer0_outputs(444)) or (layer0_outputs(2549));
    layer1_outputs(1467) <= '0';
    layer1_outputs(1468) <= not((layer0_outputs(1827)) or (layer0_outputs(172)));
    layer1_outputs(1469) <= (layer0_outputs(636)) and not (layer0_outputs(188));
    layer1_outputs(1470) <= not(layer0_outputs(1633)) or (layer0_outputs(1539));
    layer1_outputs(1471) <= '0';
    layer1_outputs(1472) <= (layer0_outputs(1558)) or (layer0_outputs(1985));
    layer1_outputs(1473) <= layer0_outputs(2191);
    layer1_outputs(1474) <= not(layer0_outputs(1203));
    layer1_outputs(1475) <= layer0_outputs(1041);
    layer1_outputs(1476) <= (layer0_outputs(2111)) or (layer0_outputs(1447));
    layer1_outputs(1477) <= (layer0_outputs(915)) or (layer0_outputs(1843));
    layer1_outputs(1478) <= (layer0_outputs(2047)) and not (layer0_outputs(1921));
    layer1_outputs(1479) <= layer0_outputs(2235);
    layer1_outputs(1480) <= layer0_outputs(1699);
    layer1_outputs(1481) <= not(layer0_outputs(881));
    layer1_outputs(1482) <= layer0_outputs(1521);
    layer1_outputs(1483) <= (layer0_outputs(1005)) and not (layer0_outputs(2));
    layer1_outputs(1484) <= layer0_outputs(1385);
    layer1_outputs(1485) <= (layer0_outputs(943)) and not (layer0_outputs(365));
    layer1_outputs(1486) <= layer0_outputs(2261);
    layer1_outputs(1487) <= not((layer0_outputs(2142)) or (layer0_outputs(150)));
    layer1_outputs(1488) <= not((layer0_outputs(2466)) xor (layer0_outputs(2010)));
    layer1_outputs(1489) <= not(layer0_outputs(426)) or (layer0_outputs(562));
    layer1_outputs(1490) <= (layer0_outputs(2247)) or (layer0_outputs(2086));
    layer1_outputs(1491) <= not(layer0_outputs(1671));
    layer1_outputs(1492) <= (layer0_outputs(1122)) or (layer0_outputs(2314));
    layer1_outputs(1493) <= not(layer0_outputs(518)) or (layer0_outputs(1353));
    layer1_outputs(1494) <= not(layer0_outputs(2380)) or (layer0_outputs(2061));
    layer1_outputs(1495) <= (layer0_outputs(105)) and (layer0_outputs(2277));
    layer1_outputs(1496) <= layer0_outputs(1971);
    layer1_outputs(1497) <= layer0_outputs(2004);
    layer1_outputs(1498) <= (layer0_outputs(865)) and (layer0_outputs(913));
    layer1_outputs(1499) <= not((layer0_outputs(1583)) and (layer0_outputs(286)));
    layer1_outputs(1500) <= layer0_outputs(2171);
    layer1_outputs(1501) <= (layer0_outputs(266)) and (layer0_outputs(1523));
    layer1_outputs(1502) <= not(layer0_outputs(1942));
    layer1_outputs(1503) <= (layer0_outputs(1662)) or (layer0_outputs(260));
    layer1_outputs(1504) <= not(layer0_outputs(2551));
    layer1_outputs(1505) <= not(layer0_outputs(2553));
    layer1_outputs(1506) <= '1';
    layer1_outputs(1507) <= layer0_outputs(1642);
    layer1_outputs(1508) <= not((layer0_outputs(672)) or (layer0_outputs(109)));
    layer1_outputs(1509) <= layer0_outputs(2544);
    layer1_outputs(1510) <= '0';
    layer1_outputs(1511) <= layer0_outputs(1991);
    layer1_outputs(1512) <= '1';
    layer1_outputs(1513) <= layer0_outputs(767);
    layer1_outputs(1514) <= (layer0_outputs(2478)) or (layer0_outputs(1641));
    layer1_outputs(1515) <= layer0_outputs(2497);
    layer1_outputs(1516) <= layer0_outputs(2346);
    layer1_outputs(1517) <= (layer0_outputs(1674)) and not (layer0_outputs(532));
    layer1_outputs(1518) <= not((layer0_outputs(2246)) and (layer0_outputs(1221)));
    layer1_outputs(1519) <= not(layer0_outputs(2120));
    layer1_outputs(1520) <= not(layer0_outputs(2245)) or (layer0_outputs(1757));
    layer1_outputs(1521) <= (layer0_outputs(1921)) and not (layer0_outputs(2351));
    layer1_outputs(1522) <= not(layer0_outputs(2004));
    layer1_outputs(1523) <= (layer0_outputs(1807)) or (layer0_outputs(280));
    layer1_outputs(1524) <= (layer0_outputs(2309)) or (layer0_outputs(903));
    layer1_outputs(1525) <= (layer0_outputs(1414)) and not (layer0_outputs(588));
    layer1_outputs(1526) <= not(layer0_outputs(531));
    layer1_outputs(1527) <= (layer0_outputs(2096)) or (layer0_outputs(829));
    layer1_outputs(1528) <= not(layer0_outputs(1638)) or (layer0_outputs(421));
    layer1_outputs(1529) <= (layer0_outputs(1426)) and not (layer0_outputs(88));
    layer1_outputs(1530) <= (layer0_outputs(1513)) and not (layer0_outputs(685));
    layer1_outputs(1531) <= not(layer0_outputs(1577)) or (layer0_outputs(655));
    layer1_outputs(1532) <= not((layer0_outputs(2095)) or (layer0_outputs(1098)));
    layer1_outputs(1533) <= (layer0_outputs(1973)) and (layer0_outputs(1474));
    layer1_outputs(1534) <= (layer0_outputs(693)) and not (layer0_outputs(1029));
    layer1_outputs(1535) <= not(layer0_outputs(209));
    layer1_outputs(1536) <= (layer0_outputs(1887)) and (layer0_outputs(1911));
    layer1_outputs(1537) <= (layer0_outputs(224)) and not (layer0_outputs(527));
    layer1_outputs(1538) <= not(layer0_outputs(1023)) or (layer0_outputs(771));
    layer1_outputs(1539) <= not(layer0_outputs(1414)) or (layer0_outputs(213));
    layer1_outputs(1540) <= layer0_outputs(1214);
    layer1_outputs(1541) <= not(layer0_outputs(2420));
    layer1_outputs(1542) <= '0';
    layer1_outputs(1543) <= layer0_outputs(1365);
    layer1_outputs(1544) <= '1';
    layer1_outputs(1545) <= not(layer0_outputs(1819));
    layer1_outputs(1546) <= not(layer0_outputs(2289));
    layer1_outputs(1547) <= layer0_outputs(1072);
    layer1_outputs(1548) <= (layer0_outputs(407)) or (layer0_outputs(2203));
    layer1_outputs(1549) <= layer0_outputs(1267);
    layer1_outputs(1550) <= (layer0_outputs(2249)) and not (layer0_outputs(649));
    layer1_outputs(1551) <= not(layer0_outputs(1522)) or (layer0_outputs(2344));
    layer1_outputs(1552) <= not(layer0_outputs(356));
    layer1_outputs(1553) <= layer0_outputs(2095);
    layer1_outputs(1554) <= (layer0_outputs(614)) and not (layer0_outputs(1776));
    layer1_outputs(1555) <= not((layer0_outputs(2049)) or (layer0_outputs(1348)));
    layer1_outputs(1556) <= layer0_outputs(2088);
    layer1_outputs(1557) <= not((layer0_outputs(2312)) or (layer0_outputs(2175)));
    layer1_outputs(1558) <= not((layer0_outputs(1411)) xor (layer0_outputs(1741)));
    layer1_outputs(1559) <= not(layer0_outputs(1723));
    layer1_outputs(1560) <= layer0_outputs(441);
    layer1_outputs(1561) <= not(layer0_outputs(1901));
    layer1_outputs(1562) <= '1';
    layer1_outputs(1563) <= layer0_outputs(2161);
    layer1_outputs(1564) <= not((layer0_outputs(1042)) xor (layer0_outputs(1973)));
    layer1_outputs(1565) <= not(layer0_outputs(2552));
    layer1_outputs(1566) <= (layer0_outputs(11)) xor (layer0_outputs(2340));
    layer1_outputs(1567) <= (layer0_outputs(1946)) and not (layer0_outputs(94));
    layer1_outputs(1568) <= not(layer0_outputs(751));
    layer1_outputs(1569) <= layer0_outputs(606);
    layer1_outputs(1570) <= not(layer0_outputs(1446)) or (layer0_outputs(1162));
    layer1_outputs(1571) <= '0';
    layer1_outputs(1572) <= not(layer0_outputs(2109));
    layer1_outputs(1573) <= layer0_outputs(455);
    layer1_outputs(1574) <= (layer0_outputs(1948)) and not (layer0_outputs(2557));
    layer1_outputs(1575) <= not(layer0_outputs(2178));
    layer1_outputs(1576) <= (layer0_outputs(1848)) and not (layer0_outputs(1888));
    layer1_outputs(1577) <= (layer0_outputs(2278)) and not (layer0_outputs(1165));
    layer1_outputs(1578) <= not((layer0_outputs(852)) or (layer0_outputs(176)));
    layer1_outputs(1579) <= not(layer0_outputs(866)) or (layer0_outputs(337));
    layer1_outputs(1580) <= layer0_outputs(1638);
    layer1_outputs(1581) <= '0';
    layer1_outputs(1582) <= (layer0_outputs(201)) and not (layer0_outputs(1319));
    layer1_outputs(1583) <= layer0_outputs(1305);
    layer1_outputs(1584) <= '1';
    layer1_outputs(1585) <= layer0_outputs(493);
    layer1_outputs(1586) <= not(layer0_outputs(632));
    layer1_outputs(1587) <= (layer0_outputs(416)) and not (layer0_outputs(1490));
    layer1_outputs(1588) <= layer0_outputs(1025);
    layer1_outputs(1589) <= (layer0_outputs(1891)) and not (layer0_outputs(2143));
    layer1_outputs(1590) <= not(layer0_outputs(303));
    layer1_outputs(1591) <= layer0_outputs(2072);
    layer1_outputs(1592) <= (layer0_outputs(2391)) and not (layer0_outputs(1449));
    layer1_outputs(1593) <= not((layer0_outputs(679)) and (layer0_outputs(1044)));
    layer1_outputs(1594) <= not(layer0_outputs(1101)) or (layer0_outputs(1696));
    layer1_outputs(1595) <= not(layer0_outputs(355));
    layer1_outputs(1596) <= '0';
    layer1_outputs(1597) <= (layer0_outputs(1898)) or (layer0_outputs(315));
    layer1_outputs(1598) <= not((layer0_outputs(1111)) and (layer0_outputs(2448)));
    layer1_outputs(1599) <= not(layer0_outputs(1366)) or (layer0_outputs(967));
    layer1_outputs(1600) <= not(layer0_outputs(1599));
    layer1_outputs(1601) <= layer0_outputs(89);
    layer1_outputs(1602) <= not(layer0_outputs(2281));
    layer1_outputs(1603) <= not((layer0_outputs(1048)) and (layer0_outputs(1884)));
    layer1_outputs(1604) <= not(layer0_outputs(91)) or (layer0_outputs(1542));
    layer1_outputs(1605) <= (layer0_outputs(591)) and not (layer0_outputs(2411));
    layer1_outputs(1606) <= '1';
    layer1_outputs(1607) <= not(layer0_outputs(275));
    layer1_outputs(1608) <= layer0_outputs(637);
    layer1_outputs(1609) <= not(layer0_outputs(126)) or (layer0_outputs(2536));
    layer1_outputs(1610) <= layer0_outputs(458);
    layer1_outputs(1611) <= not((layer0_outputs(133)) and (layer0_outputs(1001)));
    layer1_outputs(1612) <= layer0_outputs(1023);
    layer1_outputs(1613) <= not(layer0_outputs(1795)) or (layer0_outputs(1468));
    layer1_outputs(1614) <= layer0_outputs(750);
    layer1_outputs(1615) <= not(layer0_outputs(1291));
    layer1_outputs(1616) <= layer0_outputs(899);
    layer1_outputs(1617) <= not(layer0_outputs(737));
    layer1_outputs(1618) <= not((layer0_outputs(1644)) xor (layer0_outputs(895)));
    layer1_outputs(1619) <= layer0_outputs(1212);
    layer1_outputs(1620) <= not(layer0_outputs(911));
    layer1_outputs(1621) <= (layer0_outputs(1777)) and not (layer0_outputs(968));
    layer1_outputs(1622) <= (layer0_outputs(1028)) xor (layer0_outputs(594));
    layer1_outputs(1623) <= (layer0_outputs(2119)) or (layer0_outputs(1197));
    layer1_outputs(1624) <= not(layer0_outputs(2130)) or (layer0_outputs(1505));
    layer1_outputs(1625) <= layer0_outputs(756);
    layer1_outputs(1626) <= not(layer0_outputs(2421));
    layer1_outputs(1627) <= (layer0_outputs(136)) and (layer0_outputs(1681));
    layer1_outputs(1628) <= not(layer0_outputs(1985));
    layer1_outputs(1629) <= '0';
    layer1_outputs(1630) <= (layer0_outputs(2481)) and (layer0_outputs(2423));
    layer1_outputs(1631) <= layer0_outputs(1253);
    layer1_outputs(1632) <= not(layer0_outputs(880));
    layer1_outputs(1633) <= (layer0_outputs(296)) and not (layer0_outputs(2307));
    layer1_outputs(1634) <= not(layer0_outputs(2264));
    layer1_outputs(1635) <= (layer0_outputs(771)) or (layer0_outputs(1634));
    layer1_outputs(1636) <= layer0_outputs(833);
    layer1_outputs(1637) <= layer0_outputs(43);
    layer1_outputs(1638) <= (layer0_outputs(652)) and not (layer0_outputs(2068));
    layer1_outputs(1639) <= not(layer0_outputs(91));
    layer1_outputs(1640) <= not(layer0_outputs(2323));
    layer1_outputs(1641) <= (layer0_outputs(1952)) and not (layer0_outputs(1715));
    layer1_outputs(1642) <= not(layer0_outputs(647));
    layer1_outputs(1643) <= (layer0_outputs(2266)) and not (layer0_outputs(2093));
    layer1_outputs(1644) <= '1';
    layer1_outputs(1645) <= layer0_outputs(1430);
    layer1_outputs(1646) <= not(layer0_outputs(598));
    layer1_outputs(1647) <= not((layer0_outputs(994)) or (layer0_outputs(1508)));
    layer1_outputs(1648) <= layer0_outputs(1654);
    layer1_outputs(1649) <= not(layer0_outputs(882));
    layer1_outputs(1650) <= (layer0_outputs(2328)) and not (layer0_outputs(1875));
    layer1_outputs(1651) <= not((layer0_outputs(1331)) and (layer0_outputs(1476)));
    layer1_outputs(1652) <= not(layer0_outputs(476)) or (layer0_outputs(1500));
    layer1_outputs(1653) <= (layer0_outputs(1737)) and not (layer0_outputs(134));
    layer1_outputs(1654) <= not(layer0_outputs(1296)) or (layer0_outputs(2556));
    layer1_outputs(1655) <= (layer0_outputs(1265)) and not (layer0_outputs(436));
    layer1_outputs(1656) <= layer0_outputs(1567);
    layer1_outputs(1657) <= (layer0_outputs(247)) and not (layer0_outputs(25));
    layer1_outputs(1658) <= (layer0_outputs(1395)) and not (layer0_outputs(1582));
    layer1_outputs(1659) <= (layer0_outputs(2154)) and (layer0_outputs(2530));
    layer1_outputs(1660) <= layer0_outputs(74);
    layer1_outputs(1661) <= not((layer0_outputs(502)) or (layer0_outputs(1780)));
    layer1_outputs(1662) <= (layer0_outputs(1234)) or (layer0_outputs(2236));
    layer1_outputs(1663) <= not(layer0_outputs(1303));
    layer1_outputs(1664) <= layer0_outputs(2352);
    layer1_outputs(1665) <= (layer0_outputs(1156)) and not (layer0_outputs(1345));
    layer1_outputs(1666) <= layer0_outputs(292);
    layer1_outputs(1667) <= not((layer0_outputs(1187)) and (layer0_outputs(514)));
    layer1_outputs(1668) <= (layer0_outputs(446)) and not (layer0_outputs(232));
    layer1_outputs(1669) <= not(layer0_outputs(507));
    layer1_outputs(1670) <= not(layer0_outputs(1169));
    layer1_outputs(1671) <= layer0_outputs(1542);
    layer1_outputs(1672) <= layer0_outputs(1606);
    layer1_outputs(1673) <= (layer0_outputs(1750)) or (layer0_outputs(34));
    layer1_outputs(1674) <= (layer0_outputs(2495)) and not (layer0_outputs(2293));
    layer1_outputs(1675) <= (layer0_outputs(668)) and not (layer0_outputs(1625));
    layer1_outputs(1676) <= not(layer0_outputs(2407)) or (layer0_outputs(1302));
    layer1_outputs(1677) <= (layer0_outputs(819)) and not (layer0_outputs(2284));
    layer1_outputs(1678) <= (layer0_outputs(1734)) or (layer0_outputs(940));
    layer1_outputs(1679) <= layer0_outputs(1328);
    layer1_outputs(1680) <= layer0_outputs(2201);
    layer1_outputs(1681) <= not(layer0_outputs(507));
    layer1_outputs(1682) <= not((layer0_outputs(2173)) or (layer0_outputs(849)));
    layer1_outputs(1683) <= not(layer0_outputs(189));
    layer1_outputs(1684) <= (layer0_outputs(288)) and not (layer0_outputs(2016));
    layer1_outputs(1685) <= not(layer0_outputs(42));
    layer1_outputs(1686) <= (layer0_outputs(241)) and not (layer0_outputs(1437));
    layer1_outputs(1687) <= not(layer0_outputs(2537)) or (layer0_outputs(1677));
    layer1_outputs(1688) <= (layer0_outputs(2242)) and (layer0_outputs(2402));
    layer1_outputs(1689) <= not(layer0_outputs(2516));
    layer1_outputs(1690) <= not(layer0_outputs(1079)) or (layer0_outputs(1601));
    layer1_outputs(1691) <= (layer0_outputs(610)) and not (layer0_outputs(1059));
    layer1_outputs(1692) <= not((layer0_outputs(908)) or (layer0_outputs(2495)));
    layer1_outputs(1693) <= not(layer0_outputs(281)) or (layer0_outputs(1130));
    layer1_outputs(1694) <= not(layer0_outputs(1057));
    layer1_outputs(1695) <= (layer0_outputs(1035)) or (layer0_outputs(744));
    layer1_outputs(1696) <= not(layer0_outputs(1267)) or (layer0_outputs(2467));
    layer1_outputs(1697) <= not(layer0_outputs(390));
    layer1_outputs(1698) <= not((layer0_outputs(1666)) and (layer0_outputs(192)));
    layer1_outputs(1699) <= not(layer0_outputs(944)) or (layer0_outputs(2272));
    layer1_outputs(1700) <= layer0_outputs(29);
    layer1_outputs(1701) <= layer0_outputs(64);
    layer1_outputs(1702) <= not(layer0_outputs(2324)) or (layer0_outputs(2485));
    layer1_outputs(1703) <= not((layer0_outputs(897)) or (layer0_outputs(122)));
    layer1_outputs(1704) <= not(layer0_outputs(724));
    layer1_outputs(1705) <= not((layer0_outputs(323)) and (layer0_outputs(1298)));
    layer1_outputs(1706) <= layer0_outputs(935);
    layer1_outputs(1707) <= not(layer0_outputs(1937)) or (layer0_outputs(1941));
    layer1_outputs(1708) <= layer0_outputs(2099);
    layer1_outputs(1709) <= '1';
    layer1_outputs(1710) <= not(layer0_outputs(1142)) or (layer0_outputs(1213));
    layer1_outputs(1711) <= not((layer0_outputs(1364)) and (layer0_outputs(445)));
    layer1_outputs(1712) <= (layer0_outputs(614)) and (layer0_outputs(888));
    layer1_outputs(1713) <= layer0_outputs(1880);
    layer1_outputs(1714) <= (layer0_outputs(2059)) and not (layer0_outputs(1744));
    layer1_outputs(1715) <= not(layer0_outputs(769));
    layer1_outputs(1716) <= not(layer0_outputs(1948));
    layer1_outputs(1717) <= (layer0_outputs(1148)) or (layer0_outputs(1457));
    layer1_outputs(1718) <= not(layer0_outputs(597));
    layer1_outputs(1719) <= not(layer0_outputs(1845)) or (layer0_outputs(304));
    layer1_outputs(1720) <= not(layer0_outputs(860)) or (layer0_outputs(794));
    layer1_outputs(1721) <= (layer0_outputs(486)) and not (layer0_outputs(1725));
    layer1_outputs(1722) <= not(layer0_outputs(155));
    layer1_outputs(1723) <= not(layer0_outputs(76));
    layer1_outputs(1724) <= (layer0_outputs(144)) and (layer0_outputs(1704));
    layer1_outputs(1725) <= not((layer0_outputs(319)) or (layer0_outputs(1629)));
    layer1_outputs(1726) <= not(layer0_outputs(1621));
    layer1_outputs(1727) <= (layer0_outputs(1383)) and not (layer0_outputs(1975));
    layer1_outputs(1728) <= (layer0_outputs(431)) or (layer0_outputs(715));
    layer1_outputs(1729) <= not((layer0_outputs(931)) or (layer0_outputs(965)));
    layer1_outputs(1730) <= not((layer0_outputs(1436)) and (layer0_outputs(270)));
    layer1_outputs(1731) <= layer0_outputs(276);
    layer1_outputs(1732) <= (layer0_outputs(2508)) or (layer0_outputs(2392));
    layer1_outputs(1733) <= (layer0_outputs(2309)) and not (layer0_outputs(1702));
    layer1_outputs(1734) <= (layer0_outputs(563)) and not (layer0_outputs(2533));
    layer1_outputs(1735) <= (layer0_outputs(1330)) xor (layer0_outputs(1928));
    layer1_outputs(1736) <= not((layer0_outputs(284)) or (layer0_outputs(660)));
    layer1_outputs(1737) <= not(layer0_outputs(1231));
    layer1_outputs(1738) <= '0';
    layer1_outputs(1739) <= layer0_outputs(23);
    layer1_outputs(1740) <= (layer0_outputs(1241)) and not (layer0_outputs(910));
    layer1_outputs(1741) <= (layer0_outputs(435)) and (layer0_outputs(694));
    layer1_outputs(1742) <= layer0_outputs(936);
    layer1_outputs(1743) <= layer0_outputs(1794);
    layer1_outputs(1744) <= not(layer0_outputs(838)) or (layer0_outputs(154));
    layer1_outputs(1745) <= not((layer0_outputs(2077)) and (layer0_outputs(1721)));
    layer1_outputs(1746) <= not(layer0_outputs(1084));
    layer1_outputs(1747) <= layer0_outputs(2454);
    layer1_outputs(1748) <= not(layer0_outputs(2469));
    layer1_outputs(1749) <= not((layer0_outputs(1584)) xor (layer0_outputs(1321)));
    layer1_outputs(1750) <= not(layer0_outputs(973));
    layer1_outputs(1751) <= not(layer0_outputs(124));
    layer1_outputs(1752) <= not(layer0_outputs(2301)) or (layer0_outputs(182));
    layer1_outputs(1753) <= not(layer0_outputs(1220));
    layer1_outputs(1754) <= '1';
    layer1_outputs(1755) <= layer0_outputs(1909);
    layer1_outputs(1756) <= not((layer0_outputs(272)) or (layer0_outputs(2461)));
    layer1_outputs(1757) <= not(layer0_outputs(1350));
    layer1_outputs(1758) <= (layer0_outputs(2046)) and not (layer0_outputs(1499));
    layer1_outputs(1759) <= not(layer0_outputs(2085)) or (layer0_outputs(123));
    layer1_outputs(1760) <= '0';
    layer1_outputs(1761) <= (layer0_outputs(2164)) and not (layer0_outputs(155));
    layer1_outputs(1762) <= layer0_outputs(1419);
    layer1_outputs(1763) <= not(layer0_outputs(766)) or (layer0_outputs(87));
    layer1_outputs(1764) <= not((layer0_outputs(1304)) and (layer0_outputs(1412)));
    layer1_outputs(1765) <= not((layer0_outputs(863)) and (layer0_outputs(1139)));
    layer1_outputs(1766) <= (layer0_outputs(1149)) and not (layer0_outputs(586));
    layer1_outputs(1767) <= (layer0_outputs(805)) xor (layer0_outputs(1409));
    layer1_outputs(1768) <= not(layer0_outputs(1377));
    layer1_outputs(1769) <= not(layer0_outputs(1421)) or (layer0_outputs(1661));
    layer1_outputs(1770) <= layer0_outputs(791);
    layer1_outputs(1771) <= (layer0_outputs(2406)) and not (layer0_outputs(1050));
    layer1_outputs(1772) <= (layer0_outputs(729)) or (layer0_outputs(2306));
    layer1_outputs(1773) <= not(layer0_outputs(2193));
    layer1_outputs(1774) <= (layer0_outputs(1982)) and not (layer0_outputs(1002));
    layer1_outputs(1775) <= not(layer0_outputs(1713));
    layer1_outputs(1776) <= '0';
    layer1_outputs(1777) <= (layer0_outputs(511)) or (layer0_outputs(1369));
    layer1_outputs(1778) <= (layer0_outputs(200)) and not (layer0_outputs(268));
    layer1_outputs(1779) <= (layer0_outputs(1915)) and not (layer0_outputs(1902));
    layer1_outputs(1780) <= not(layer0_outputs(978)) or (layer0_outputs(329));
    layer1_outputs(1781) <= '1';
    layer1_outputs(1782) <= not(layer0_outputs(530)) or (layer0_outputs(2115));
    layer1_outputs(1783) <= '0';
    layer1_outputs(1784) <= (layer0_outputs(1847)) and not (layer0_outputs(1607));
    layer1_outputs(1785) <= (layer0_outputs(879)) and (layer0_outputs(244));
    layer1_outputs(1786) <= not((layer0_outputs(1594)) or (layer0_outputs(391)));
    layer1_outputs(1787) <= not((layer0_outputs(622)) and (layer0_outputs(955)));
    layer1_outputs(1788) <= not(layer0_outputs(1846));
    layer1_outputs(1789) <= not(layer0_outputs(259)) or (layer0_outputs(2154));
    layer1_outputs(1790) <= layer0_outputs(2502);
    layer1_outputs(1791) <= (layer0_outputs(1235)) and not (layer0_outputs(1808));
    layer1_outputs(1792) <= (layer0_outputs(277)) or (layer0_outputs(1953));
    layer1_outputs(1793) <= '0';
    layer1_outputs(1794) <= layer0_outputs(1914);
    layer1_outputs(1795) <= not((layer0_outputs(552)) and (layer0_outputs(1293)));
    layer1_outputs(1796) <= (layer0_outputs(579)) or (layer0_outputs(1381));
    layer1_outputs(1797) <= not(layer0_outputs(593)) or (layer0_outputs(899));
    layer1_outputs(1798) <= not(layer0_outputs(1805)) or (layer0_outputs(2022));
    layer1_outputs(1799) <= layer0_outputs(2287);
    layer1_outputs(1800) <= not(layer0_outputs(137));
    layer1_outputs(1801) <= not(layer0_outputs(2145)) or (layer0_outputs(1210));
    layer1_outputs(1802) <= not(layer0_outputs(804)) or (layer0_outputs(2173));
    layer1_outputs(1803) <= layer0_outputs(1598);
    layer1_outputs(1804) <= layer0_outputs(969);
    layer1_outputs(1805) <= (layer0_outputs(1577)) or (layer0_outputs(806));
    layer1_outputs(1806) <= not(layer0_outputs(1737)) or (layer0_outputs(1986));
    layer1_outputs(1807) <= not((layer0_outputs(1433)) or (layer0_outputs(1196)));
    layer1_outputs(1808) <= not(layer0_outputs(665));
    layer1_outputs(1809) <= not(layer0_outputs(978));
    layer1_outputs(1810) <= not(layer0_outputs(649));
    layer1_outputs(1811) <= '0';
    layer1_outputs(1812) <= not(layer0_outputs(31));
    layer1_outputs(1813) <= layer0_outputs(1624);
    layer1_outputs(1814) <= '0';
    layer1_outputs(1815) <= (layer0_outputs(967)) and (layer0_outputs(1166));
    layer1_outputs(1816) <= not((layer0_outputs(380)) or (layer0_outputs(569)));
    layer1_outputs(1817) <= (layer0_outputs(1399)) and not (layer0_outputs(2268));
    layer1_outputs(1818) <= (layer0_outputs(2106)) or (layer0_outputs(2298));
    layer1_outputs(1819) <= not(layer0_outputs(1856)) or (layer0_outputs(1144));
    layer1_outputs(1820) <= (layer0_outputs(2373)) and not (layer0_outputs(895));
    layer1_outputs(1821) <= '0';
    layer1_outputs(1822) <= not(layer0_outputs(282));
    layer1_outputs(1823) <= not((layer0_outputs(435)) and (layer0_outputs(1831)));
    layer1_outputs(1824) <= '0';
    layer1_outputs(1825) <= (layer0_outputs(990)) and (layer0_outputs(1681));
    layer1_outputs(1826) <= not(layer0_outputs(975)) or (layer0_outputs(934));
    layer1_outputs(1827) <= layer0_outputs(499);
    layer1_outputs(1828) <= not((layer0_outputs(1982)) and (layer0_outputs(2480)));
    layer1_outputs(1829) <= (layer0_outputs(2071)) or (layer0_outputs(121));
    layer1_outputs(1830) <= layer0_outputs(2120);
    layer1_outputs(1831) <= (layer0_outputs(95)) or (layer0_outputs(2472));
    layer1_outputs(1832) <= (layer0_outputs(1605)) and not (layer0_outputs(852));
    layer1_outputs(1833) <= not(layer0_outputs(220));
    layer1_outputs(1834) <= '0';
    layer1_outputs(1835) <= (layer0_outputs(369)) and not (layer0_outputs(2501));
    layer1_outputs(1836) <= not(layer0_outputs(205));
    layer1_outputs(1837) <= (layer0_outputs(1743)) and not (layer0_outputs(2170));
    layer1_outputs(1838) <= (layer0_outputs(2302)) and (layer0_outputs(2458));
    layer1_outputs(1839) <= (layer0_outputs(506)) xor (layer0_outputs(432));
    layer1_outputs(1840) <= (layer0_outputs(1364)) and not (layer0_outputs(2337));
    layer1_outputs(1841) <= (layer0_outputs(1083)) or (layer0_outputs(558));
    layer1_outputs(1842) <= (layer0_outputs(503)) or (layer0_outputs(1289));
    layer1_outputs(1843) <= not(layer0_outputs(1088));
    layer1_outputs(1844) <= (layer0_outputs(1854)) and (layer0_outputs(258));
    layer1_outputs(1845) <= (layer0_outputs(871)) and (layer0_outputs(496));
    layer1_outputs(1846) <= (layer0_outputs(1379)) or (layer0_outputs(1443));
    layer1_outputs(1847) <= (layer0_outputs(908)) or (layer0_outputs(873));
    layer1_outputs(1848) <= '0';
    layer1_outputs(1849) <= not(layer0_outputs(627)) or (layer0_outputs(740));
    layer1_outputs(1850) <= layer0_outputs(568);
    layer1_outputs(1851) <= not(layer0_outputs(945)) or (layer0_outputs(1871));
    layer1_outputs(1852) <= layer0_outputs(826);
    layer1_outputs(1853) <= layer0_outputs(1678);
    layer1_outputs(1854) <= not(layer0_outputs(777));
    layer1_outputs(1855) <= not(layer0_outputs(2026)) or (layer0_outputs(39));
    layer1_outputs(1856) <= layer0_outputs(528);
    layer1_outputs(1857) <= layer0_outputs(1859);
    layer1_outputs(1858) <= '0';
    layer1_outputs(1859) <= layer0_outputs(2230);
    layer1_outputs(1860) <= not((layer0_outputs(1159)) and (layer0_outputs(2156)));
    layer1_outputs(1861) <= not(layer0_outputs(788)) or (layer0_outputs(635));
    layer1_outputs(1862) <= '0';
    layer1_outputs(1863) <= not(layer0_outputs(425));
    layer1_outputs(1864) <= not(layer0_outputs(437));
    layer1_outputs(1865) <= layer0_outputs(459);
    layer1_outputs(1866) <= not(layer0_outputs(115));
    layer1_outputs(1867) <= not(layer0_outputs(1568));
    layer1_outputs(1868) <= not(layer0_outputs(1746));
    layer1_outputs(1869) <= (layer0_outputs(568)) or (layer0_outputs(1170));
    layer1_outputs(1870) <= not(layer0_outputs(2426));
    layer1_outputs(1871) <= not(layer0_outputs(1057));
    layer1_outputs(1872) <= not(layer0_outputs(1030)) or (layer0_outputs(2457));
    layer1_outputs(1873) <= (layer0_outputs(868)) and not (layer0_outputs(2294));
    layer1_outputs(1874) <= layer0_outputs(2443);
    layer1_outputs(1875) <= not((layer0_outputs(2432)) or (layer0_outputs(2316)));
    layer1_outputs(1876) <= (layer0_outputs(85)) and not (layer0_outputs(875));
    layer1_outputs(1877) <= not(layer0_outputs(2128)) or (layer0_outputs(2411));
    layer1_outputs(1878) <= not((layer0_outputs(877)) or (layer0_outputs(1294)));
    layer1_outputs(1879) <= (layer0_outputs(194)) or (layer0_outputs(2194));
    layer1_outputs(1880) <= not((layer0_outputs(927)) or (layer0_outputs(2172)));
    layer1_outputs(1881) <= layer0_outputs(2376);
    layer1_outputs(1882) <= layer0_outputs(1205);
    layer1_outputs(1883) <= not(layer0_outputs(2303));
    layer1_outputs(1884) <= not(layer0_outputs(1775)) or (layer0_outputs(540));
    layer1_outputs(1885) <= not((layer0_outputs(1389)) and (layer0_outputs(1812)));
    layer1_outputs(1886) <= not(layer0_outputs(977));
    layer1_outputs(1887) <= layer0_outputs(321);
    layer1_outputs(1888) <= (layer0_outputs(1477)) and (layer0_outputs(1094));
    layer1_outputs(1889) <= layer0_outputs(880);
    layer1_outputs(1890) <= not(layer0_outputs(2279));
    layer1_outputs(1891) <= layer0_outputs(1096);
    layer1_outputs(1892) <= not(layer0_outputs(1440)) or (layer0_outputs(1359));
    layer1_outputs(1893) <= not(layer0_outputs(325));
    layer1_outputs(1894) <= not(layer0_outputs(1938)) or (layer0_outputs(643));
    layer1_outputs(1895) <= layer0_outputs(248);
    layer1_outputs(1896) <= not(layer0_outputs(2470)) or (layer0_outputs(1842));
    layer1_outputs(1897) <= not(layer0_outputs(854));
    layer1_outputs(1898) <= not((layer0_outputs(305)) and (layer0_outputs(1751)));
    layer1_outputs(1899) <= not(layer0_outputs(2451));
    layer1_outputs(1900) <= (layer0_outputs(1647)) and not (layer0_outputs(2371));
    layer1_outputs(1901) <= layer0_outputs(1645);
    layer1_outputs(1902) <= not(layer0_outputs(1797)) or (layer0_outputs(504));
    layer1_outputs(1903) <= not(layer0_outputs(813));
    layer1_outputs(1904) <= layer0_outputs(828);
    layer1_outputs(1905) <= not(layer0_outputs(498));
    layer1_outputs(1906) <= not(layer0_outputs(540));
    layer1_outputs(1907) <= layer0_outputs(1275);
    layer1_outputs(1908) <= (layer0_outputs(2275)) and (layer0_outputs(1035));
    layer1_outputs(1909) <= (layer0_outputs(356)) and not (layer0_outputs(327));
    layer1_outputs(1910) <= layer0_outputs(2096);
    layer1_outputs(1911) <= not((layer0_outputs(344)) and (layer0_outputs(466)));
    layer1_outputs(1912) <= layer0_outputs(1417);
    layer1_outputs(1913) <= not((layer0_outputs(648)) xor (layer0_outputs(1868)));
    layer1_outputs(1914) <= (layer0_outputs(1226)) or (layer0_outputs(1510));
    layer1_outputs(1915) <= (layer0_outputs(1671)) and not (layer0_outputs(1156));
    layer1_outputs(1916) <= layer0_outputs(876);
    layer1_outputs(1917) <= (layer0_outputs(30)) and not (layer0_outputs(311));
    layer1_outputs(1918) <= layer0_outputs(1942);
    layer1_outputs(1919) <= '1';
    layer1_outputs(1920) <= layer0_outputs(482);
    layer1_outputs(1921) <= not(layer0_outputs(2042)) or (layer0_outputs(2370));
    layer1_outputs(1922) <= layer0_outputs(256);
    layer1_outputs(1923) <= '0';
    layer1_outputs(1924) <= (layer0_outputs(2345)) and (layer0_outputs(1249));
    layer1_outputs(1925) <= layer0_outputs(980);
    layer1_outputs(1926) <= (layer0_outputs(1054)) xor (layer0_outputs(2488));
    layer1_outputs(1927) <= (layer0_outputs(850)) and not (layer0_outputs(2295));
    layer1_outputs(1928) <= not(layer0_outputs(1867));
    layer1_outputs(1929) <= (layer0_outputs(2552)) and (layer0_outputs(1741));
    layer1_outputs(1930) <= layer0_outputs(427);
    layer1_outputs(1931) <= not(layer0_outputs(1017)) or (layer0_outputs(2521));
    layer1_outputs(1932) <= '1';
    layer1_outputs(1933) <= (layer0_outputs(259)) and not (layer0_outputs(104));
    layer1_outputs(1934) <= (layer0_outputs(928)) and not (layer0_outputs(905));
    layer1_outputs(1935) <= (layer0_outputs(42)) or (layer0_outputs(959));
    layer1_outputs(1936) <= (layer0_outputs(2240)) or (layer0_outputs(1300));
    layer1_outputs(1937) <= layer0_outputs(416);
    layer1_outputs(1938) <= not(layer0_outputs(523)) or (layer0_outputs(2070));
    layer1_outputs(1939) <= (layer0_outputs(1608)) xor (layer0_outputs(2256));
    layer1_outputs(1940) <= layer0_outputs(1923);
    layer1_outputs(1941) <= not((layer0_outputs(1816)) and (layer0_outputs(1358)));
    layer1_outputs(1942) <= layer0_outputs(1046);
    layer1_outputs(1943) <= not(layer0_outputs(2509)) or (layer0_outputs(2129));
    layer1_outputs(1944) <= layer0_outputs(1596);
    layer1_outputs(1945) <= (layer0_outputs(860)) or (layer0_outputs(2057));
    layer1_outputs(1946) <= (layer0_outputs(7)) and not (layer0_outputs(2384));
    layer1_outputs(1947) <= (layer0_outputs(2005)) and (layer0_outputs(780));
    layer1_outputs(1948) <= layer0_outputs(1815);
    layer1_outputs(1949) <= not(layer0_outputs(162)) or (layer0_outputs(1550));
    layer1_outputs(1950) <= not(layer0_outputs(1844)) or (layer0_outputs(2311));
    layer1_outputs(1951) <= layer0_outputs(1250);
    layer1_outputs(1952) <= not(layer0_outputs(1042));
    layer1_outputs(1953) <= (layer0_outputs(1655)) or (layer0_outputs(1304));
    layer1_outputs(1954) <= (layer0_outputs(684)) xor (layer0_outputs(2058));
    layer1_outputs(1955) <= not(layer0_outputs(231)) or (layer0_outputs(164));
    layer1_outputs(1956) <= layer0_outputs(955);
    layer1_outputs(1957) <= layer0_outputs(1281);
    layer1_outputs(1958) <= not(layer0_outputs(1981)) or (layer0_outputs(2009));
    layer1_outputs(1959) <= not(layer0_outputs(878));
    layer1_outputs(1960) <= layer0_outputs(178);
    layer1_outputs(1961) <= (layer0_outputs(2364)) and not (layer0_outputs(1905));
    layer1_outputs(1962) <= layer0_outputs(1099);
    layer1_outputs(1963) <= not(layer0_outputs(2436));
    layer1_outputs(1964) <= not(layer0_outputs(2114));
    layer1_outputs(1965) <= not((layer0_outputs(398)) and (layer0_outputs(278)));
    layer1_outputs(1966) <= not(layer0_outputs(1094));
    layer1_outputs(1967) <= layer0_outputs(2286);
    layer1_outputs(1968) <= not((layer0_outputs(14)) and (layer0_outputs(2255)));
    layer1_outputs(1969) <= (layer0_outputs(1372)) and not (layer0_outputs(2062));
    layer1_outputs(1970) <= not(layer0_outputs(781)) or (layer0_outputs(1593));
    layer1_outputs(1971) <= not(layer0_outputs(350));
    layer1_outputs(1972) <= not(layer0_outputs(1427));
    layer1_outputs(1973) <= layer0_outputs(138);
    layer1_outputs(1974) <= layer0_outputs(1733);
    layer1_outputs(1975) <= not((layer0_outputs(942)) and (layer0_outputs(1849)));
    layer1_outputs(1976) <= not(layer0_outputs(111)) or (layer0_outputs(1443));
    layer1_outputs(1977) <= '0';
    layer1_outputs(1978) <= (layer0_outputs(2152)) or (layer0_outputs(1012));
    layer1_outputs(1979) <= not(layer0_outputs(2023));
    layer1_outputs(1980) <= not((layer0_outputs(381)) and (layer0_outputs(1555)));
    layer1_outputs(1981) <= '1';
    layer1_outputs(1982) <= layer0_outputs(1244);
    layer1_outputs(1983) <= (layer0_outputs(575)) or (layer0_outputs(1373));
    layer1_outputs(1984) <= not(layer0_outputs(2500));
    layer1_outputs(1985) <= not(layer0_outputs(1627));
    layer1_outputs(1986) <= not(layer0_outputs(1735));
    layer1_outputs(1987) <= not(layer0_outputs(20));
    layer1_outputs(1988) <= not(layer0_outputs(2070));
    layer1_outputs(1989) <= not(layer0_outputs(362)) or (layer0_outputs(1859));
    layer1_outputs(1990) <= '1';
    layer1_outputs(1991) <= '0';
    layer1_outputs(1992) <= not(layer0_outputs(1527)) or (layer0_outputs(1174));
    layer1_outputs(1993) <= not((layer0_outputs(2102)) or (layer0_outputs(1300)));
    layer1_outputs(1994) <= layer0_outputs(1615);
    layer1_outputs(1995) <= layer0_outputs(1722);
    layer1_outputs(1996) <= not(layer0_outputs(2418));
    layer1_outputs(1997) <= not(layer0_outputs(998)) or (layer0_outputs(1657));
    layer1_outputs(1998) <= (layer0_outputs(2102)) or (layer0_outputs(2436));
    layer1_outputs(1999) <= not(layer0_outputs(1080)) or (layer0_outputs(940));
    layer1_outputs(2000) <= (layer0_outputs(1172)) and (layer0_outputs(768));
    layer1_outputs(2001) <= not(layer0_outputs(1313));
    layer1_outputs(2002) <= not(layer0_outputs(30)) or (layer0_outputs(123));
    layer1_outputs(2003) <= layer0_outputs(1679);
    layer1_outputs(2004) <= (layer0_outputs(228)) and (layer0_outputs(1869));
    layer1_outputs(2005) <= not(layer0_outputs(1120));
    layer1_outputs(2006) <= not((layer0_outputs(2039)) xor (layer0_outputs(1652)));
    layer1_outputs(2007) <= (layer0_outputs(2266)) and not (layer0_outputs(765));
    layer1_outputs(2008) <= layer0_outputs(265);
    layer1_outputs(2009) <= not(layer0_outputs(2024));
    layer1_outputs(2010) <= layer0_outputs(177);
    layer1_outputs(2011) <= not(layer0_outputs(541)) or (layer0_outputs(117));
    layer1_outputs(2012) <= not((layer0_outputs(1722)) and (layer0_outputs(2073)));
    layer1_outputs(2013) <= not(layer0_outputs(1336));
    layer1_outputs(2014) <= '1';
    layer1_outputs(2015) <= not(layer0_outputs(80)) or (layer0_outputs(226));
    layer1_outputs(2016) <= layer0_outputs(2146);
    layer1_outputs(2017) <= layer0_outputs(670);
    layer1_outputs(2018) <= layer0_outputs(2276);
    layer1_outputs(2019) <= (layer0_outputs(1476)) xor (layer0_outputs(424));
    layer1_outputs(2020) <= not(layer0_outputs(1435));
    layer1_outputs(2021) <= layer0_outputs(770);
    layer1_outputs(2022) <= layer0_outputs(544);
    layer1_outputs(2023) <= (layer0_outputs(1326)) and (layer0_outputs(2230));
    layer1_outputs(2024) <= not(layer0_outputs(2275));
    layer1_outputs(2025) <= (layer0_outputs(2267)) or (layer0_outputs(1332));
    layer1_outputs(2026) <= not((layer0_outputs(1736)) and (layer0_outputs(1817)));
    layer1_outputs(2027) <= not((layer0_outputs(761)) and (layer0_outputs(410)));
    layer1_outputs(2028) <= layer0_outputs(2185);
    layer1_outputs(2029) <= layer0_outputs(721);
    layer1_outputs(2030) <= (layer0_outputs(971)) and not (layer0_outputs(1268));
    layer1_outputs(2031) <= layer0_outputs(1136);
    layer1_outputs(2032) <= layer0_outputs(2437);
    layer1_outputs(2033) <= '1';
    layer1_outputs(2034) <= not(layer0_outputs(1339)) or (layer0_outputs(1770));
    layer1_outputs(2035) <= layer0_outputs(1908);
    layer1_outputs(2036) <= not(layer0_outputs(926)) or (layer0_outputs(849));
    layer1_outputs(2037) <= not(layer0_outputs(98)) or (layer0_outputs(13));
    layer1_outputs(2038) <= not((layer0_outputs(1780)) or (layer0_outputs(656)));
    layer1_outputs(2039) <= not((layer0_outputs(867)) and (layer0_outputs(1837)));
    layer1_outputs(2040) <= not((layer0_outputs(1765)) or (layer0_outputs(2550)));
    layer1_outputs(2041) <= not(layer0_outputs(82));
    layer1_outputs(2042) <= (layer0_outputs(867)) and not (layer0_outputs(1897));
    layer1_outputs(2043) <= (layer0_outputs(12)) or (layer0_outputs(1628));
    layer1_outputs(2044) <= (layer0_outputs(1551)) and (layer0_outputs(1823));
    layer1_outputs(2045) <= layer0_outputs(639);
    layer1_outputs(2046) <= (layer0_outputs(2057)) and not (layer0_outputs(1504));
    layer1_outputs(2047) <= layer0_outputs(611);
    layer1_outputs(2048) <= layer0_outputs(2331);
    layer1_outputs(2049) <= (layer0_outputs(2073)) and (layer0_outputs(762));
    layer1_outputs(2050) <= not(layer0_outputs(1090));
    layer1_outputs(2051) <= (layer0_outputs(1213)) and not (layer0_outputs(333));
    layer1_outputs(2052) <= '1';
    layer1_outputs(2053) <= not(layer0_outputs(1762)) or (layer0_outputs(1863));
    layer1_outputs(2054) <= not((layer0_outputs(1371)) or (layer0_outputs(83)));
    layer1_outputs(2055) <= (layer0_outputs(1552)) or (layer0_outputs(1049));
    layer1_outputs(2056) <= not(layer0_outputs(6));
    layer1_outputs(2057) <= (layer0_outputs(1052)) and not (layer0_outputs(1781));
    layer1_outputs(2058) <= not(layer0_outputs(2232)) or (layer0_outputs(1270));
    layer1_outputs(2059) <= (layer0_outputs(607)) and not (layer0_outputs(2533));
    layer1_outputs(2060) <= not(layer0_outputs(1877)) or (layer0_outputs(929));
    layer1_outputs(2061) <= not(layer0_outputs(2112)) or (layer0_outputs(1182));
    layer1_outputs(2062) <= (layer0_outputs(1408)) or (layer0_outputs(1406));
    layer1_outputs(2063) <= layer0_outputs(1436);
    layer1_outputs(2064) <= not(layer0_outputs(1873));
    layer1_outputs(2065) <= layer0_outputs(991);
    layer1_outputs(2066) <= not(layer0_outputs(15)) or (layer0_outputs(476));
    layer1_outputs(2067) <= (layer0_outputs(1501)) or (layer0_outputs(1825));
    layer1_outputs(2068) <= not((layer0_outputs(982)) xor (layer0_outputs(779)));
    layer1_outputs(2069) <= '0';
    layer1_outputs(2070) <= not(layer0_outputs(990)) or (layer0_outputs(2034));
    layer1_outputs(2071) <= not(layer0_outputs(847)) or (layer0_outputs(1552));
    layer1_outputs(2072) <= layer0_outputs(1796);
    layer1_outputs(2073) <= not(layer0_outputs(380));
    layer1_outputs(2074) <= not(layer0_outputs(2415));
    layer1_outputs(2075) <= not(layer0_outputs(2122));
    layer1_outputs(2076) <= not(layer0_outputs(2044)) or (layer0_outputs(674));
    layer1_outputs(2077) <= not((layer0_outputs(389)) or (layer0_outputs(2228)));
    layer1_outputs(2078) <= not((layer0_outputs(146)) and (layer0_outputs(2257)));
    layer1_outputs(2079) <= not((layer0_outputs(1099)) or (layer0_outputs(1095)));
    layer1_outputs(2080) <= not(layer0_outputs(1347));
    layer1_outputs(2081) <= not(layer0_outputs(2498)) or (layer0_outputs(550));
    layer1_outputs(2082) <= not(layer0_outputs(2503));
    layer1_outputs(2083) <= not((layer0_outputs(1503)) xor (layer0_outputs(1160)));
    layer1_outputs(2084) <= not(layer0_outputs(120));
    layer1_outputs(2085) <= (layer0_outputs(2478)) and not (layer0_outputs(1481));
    layer1_outputs(2086) <= layer0_outputs(1531);
    layer1_outputs(2087) <= not(layer0_outputs(700));
    layer1_outputs(2088) <= layer0_outputs(1847);
    layer1_outputs(2089) <= not((layer0_outputs(2273)) and (layer0_outputs(414)));
    layer1_outputs(2090) <= not(layer0_outputs(439));
    layer1_outputs(2091) <= (layer0_outputs(403)) and not (layer0_outputs(1188));
    layer1_outputs(2092) <= not(layer0_outputs(2471));
    layer1_outputs(2093) <= not((layer0_outputs(900)) and (layer0_outputs(2320)));
    layer1_outputs(2094) <= not(layer0_outputs(1080));
    layer1_outputs(2095) <= layer0_outputs(862);
    layer1_outputs(2096) <= layer0_outputs(2180);
    layer1_outputs(2097) <= layer0_outputs(1433);
    layer1_outputs(2098) <= not(layer0_outputs(1498)) or (layer0_outputs(333));
    layer1_outputs(2099) <= (layer0_outputs(741)) and not (layer0_outputs(912));
    layer1_outputs(2100) <= not((layer0_outputs(375)) or (layer0_outputs(648)));
    layer1_outputs(2101) <= (layer0_outputs(265)) and not (layer0_outputs(2050));
    layer1_outputs(2102) <= layer0_outputs(486);
    layer1_outputs(2103) <= (layer0_outputs(2089)) and (layer0_outputs(493));
    layer1_outputs(2104) <= layer0_outputs(393);
    layer1_outputs(2105) <= layer0_outputs(1238);
    layer1_outputs(2106) <= (layer0_outputs(1337)) and not (layer0_outputs(1537));
    layer1_outputs(2107) <= (layer0_outputs(1501)) or (layer0_outputs(934));
    layer1_outputs(2108) <= not((layer0_outputs(2337)) or (layer0_outputs(9)));
    layer1_outputs(2109) <= (layer0_outputs(958)) xor (layer0_outputs(264));
    layer1_outputs(2110) <= layer0_outputs(1706);
    layer1_outputs(2111) <= not((layer0_outputs(2527)) and (layer0_outputs(1648)));
    layer1_outputs(2112) <= not(layer0_outputs(2025)) or (layer0_outputs(2332));
    layer1_outputs(2113) <= layer0_outputs(2475);
    layer1_outputs(2114) <= not(layer0_outputs(1183));
    layer1_outputs(2115) <= (layer0_outputs(485)) or (layer0_outputs(1716));
    layer1_outputs(2116) <= (layer0_outputs(2100)) and not (layer0_outputs(1754));
    layer1_outputs(2117) <= (layer0_outputs(1721)) or (layer0_outputs(2133));
    layer1_outputs(2118) <= not(layer0_outputs(1505));
    layer1_outputs(2119) <= not(layer0_outputs(2475));
    layer1_outputs(2120) <= (layer0_outputs(1405)) or (layer0_outputs(1931));
    layer1_outputs(2121) <= (layer0_outputs(538)) and (layer0_outputs(483));
    layer1_outputs(2122) <= (layer0_outputs(519)) and not (layer0_outputs(1811));
    layer1_outputs(2123) <= not(layer0_outputs(312));
    layer1_outputs(2124) <= layer0_outputs(1310);
    layer1_outputs(2125) <= not(layer0_outputs(1669));
    layer1_outputs(2126) <= '0';
    layer1_outputs(2127) <= layer0_outputs(217);
    layer1_outputs(2128) <= (layer0_outputs(1574)) and (layer0_outputs(2158));
    layer1_outputs(2129) <= not(layer0_outputs(963));
    layer1_outputs(2130) <= (layer0_outputs(735)) and not (layer0_outputs(1961));
    layer1_outputs(2131) <= not(layer0_outputs(346));
    layer1_outputs(2132) <= layer0_outputs(1881);
    layer1_outputs(2133) <= layer0_outputs(1320);
    layer1_outputs(2134) <= (layer0_outputs(305)) and (layer0_outputs(2183));
    layer1_outputs(2135) <= layer0_outputs(1696);
    layer1_outputs(2136) <= not(layer0_outputs(1278));
    layer1_outputs(2137) <= (layer0_outputs(2404)) and not (layer0_outputs(2006));
    layer1_outputs(2138) <= not(layer0_outputs(892));
    layer1_outputs(2139) <= '1';
    layer1_outputs(2140) <= (layer0_outputs(79)) or (layer0_outputs(2037));
    layer1_outputs(2141) <= layer0_outputs(652);
    layer1_outputs(2142) <= (layer0_outputs(2082)) or (layer0_outputs(1146));
    layer1_outputs(2143) <= not((layer0_outputs(1439)) or (layer0_outputs(1927)));
    layer1_outputs(2144) <= not((layer0_outputs(2397)) or (layer0_outputs(387)));
    layer1_outputs(2145) <= (layer0_outputs(800)) and not (layer0_outputs(1));
    layer1_outputs(2146) <= not(layer0_outputs(851));
    layer1_outputs(2147) <= not((layer0_outputs(1338)) and (layer0_outputs(554)));
    layer1_outputs(2148) <= not((layer0_outputs(1383)) and (layer0_outputs(1195)));
    layer1_outputs(2149) <= not(layer0_outputs(1247)) or (layer0_outputs(1067));
    layer1_outputs(2150) <= not(layer0_outputs(1017));
    layer1_outputs(2151) <= layer0_outputs(487);
    layer1_outputs(2152) <= not((layer0_outputs(2078)) and (layer0_outputs(1977)));
    layer1_outputs(2153) <= (layer0_outputs(2018)) and not (layer0_outputs(2294));
    layer1_outputs(2154) <= not(layer0_outputs(692));
    layer1_outputs(2155) <= not((layer0_outputs(718)) and (layer0_outputs(1511)));
    layer1_outputs(2156) <= (layer0_outputs(1754)) or (layer0_outputs(2151));
    layer1_outputs(2157) <= not(layer0_outputs(494)) or (layer0_outputs(1629));
    layer1_outputs(2158) <= not(layer0_outputs(1098));
    layer1_outputs(2159) <= not(layer0_outputs(1872)) or (layer0_outputs(885));
    layer1_outputs(2160) <= (layer0_outputs(479)) and not (layer0_outputs(1814));
    layer1_outputs(2161) <= not(layer0_outputs(1110)) or (layer0_outputs(73));
    layer1_outputs(2162) <= (layer0_outputs(1397)) or (layer0_outputs(127));
    layer1_outputs(2163) <= not(layer0_outputs(2322)) or (layer0_outputs(2358));
    layer1_outputs(2164) <= '0';
    layer1_outputs(2165) <= '0';
    layer1_outputs(2166) <= '1';
    layer1_outputs(2167) <= not(layer0_outputs(2163));
    layer1_outputs(2168) <= (layer0_outputs(2297)) or (layer0_outputs(200));
    layer1_outputs(2169) <= '0';
    layer1_outputs(2170) <= not(layer0_outputs(268));
    layer1_outputs(2171) <= not((layer0_outputs(11)) and (layer0_outputs(366)));
    layer1_outputs(2172) <= (layer0_outputs(2211)) or (layer0_outputs(1153));
    layer1_outputs(2173) <= not(layer0_outputs(1555)) or (layer0_outputs(833));
    layer1_outputs(2174) <= not((layer0_outputs(764)) or (layer0_outputs(242)));
    layer1_outputs(2175) <= (layer0_outputs(2540)) and (layer0_outputs(300));
    layer1_outputs(2176) <= (layer0_outputs(202)) and not (layer0_outputs(2401));
    layer1_outputs(2177) <= not((layer0_outputs(1193)) or (layer0_outputs(284)));
    layer1_outputs(2178) <= (layer0_outputs(1019)) or (layer0_outputs(1967));
    layer1_outputs(2179) <= '1';
    layer1_outputs(2180) <= not(layer0_outputs(1239)) or (layer0_outputs(1429));
    layer1_outputs(2181) <= not(layer0_outputs(1933)) or (layer0_outputs(601));
    layer1_outputs(2182) <= not(layer0_outputs(877));
    layer1_outputs(2183) <= not((layer0_outputs(1341)) and (layer0_outputs(440)));
    layer1_outputs(2184) <= not(layer0_outputs(2063));
    layer1_outputs(2185) <= not(layer0_outputs(862)) or (layer0_outputs(1957));
    layer1_outputs(2186) <= not(layer0_outputs(704)) or (layer0_outputs(1422));
    layer1_outputs(2187) <= (layer0_outputs(1254)) and not (layer0_outputs(135));
    layer1_outputs(2188) <= layer0_outputs(343);
    layer1_outputs(2189) <= (layer0_outputs(479)) and (layer0_outputs(2223));
    layer1_outputs(2190) <= (layer0_outputs(385)) and not (layer0_outputs(1520));
    layer1_outputs(2191) <= layer0_outputs(855);
    layer1_outputs(2192) <= (layer0_outputs(2033)) and (layer0_outputs(1220));
    layer1_outputs(2193) <= (layer0_outputs(452)) and not (layer0_outputs(526));
    layer1_outputs(2194) <= '1';
    layer1_outputs(2195) <= layer0_outputs(96);
    layer1_outputs(2196) <= (layer0_outputs(2093)) and not (layer0_outputs(1444));
    layer1_outputs(2197) <= not(layer0_outputs(2011));
    layer1_outputs(2198) <= (layer0_outputs(2107)) or (layer0_outputs(347));
    layer1_outputs(2199) <= (layer0_outputs(2491)) and not (layer0_outputs(283));
    layer1_outputs(2200) <= layer0_outputs(694);
    layer1_outputs(2201) <= not(layer0_outputs(2246));
    layer1_outputs(2202) <= not(layer0_outputs(1));
    layer1_outputs(2203) <= layer0_outputs(831);
    layer1_outputs(2204) <= (layer0_outputs(301)) and (layer0_outputs(1260));
    layer1_outputs(2205) <= not((layer0_outputs(1385)) and (layer0_outputs(2511)));
    layer1_outputs(2206) <= not(layer0_outputs(2166)) or (layer0_outputs(1898));
    layer1_outputs(2207) <= layer0_outputs(1085);
    layer1_outputs(2208) <= not(layer0_outputs(469));
    layer1_outputs(2209) <= not((layer0_outputs(2347)) and (layer0_outputs(323)));
    layer1_outputs(2210) <= not(layer0_outputs(1075)) or (layer0_outputs(378));
    layer1_outputs(2211) <= not(layer0_outputs(177)) or (layer0_outputs(883));
    layer1_outputs(2212) <= not(layer0_outputs(1087));
    layer1_outputs(2213) <= layer0_outputs(1955);
    layer1_outputs(2214) <= not(layer0_outputs(1155)) or (layer0_outputs(680));
    layer1_outputs(2215) <= layer0_outputs(1927);
    layer1_outputs(2216) <= layer0_outputs(720);
    layer1_outputs(2217) <= layer0_outputs(322);
    layer1_outputs(2218) <= '1';
    layer1_outputs(2219) <= (layer0_outputs(1024)) or (layer0_outputs(10));
    layer1_outputs(2220) <= layer0_outputs(358);
    layer1_outputs(2221) <= '1';
    layer1_outputs(2222) <= '1';
    layer1_outputs(2223) <= not(layer0_outputs(302));
    layer1_outputs(2224) <= layer0_outputs(2460);
    layer1_outputs(2225) <= layer0_outputs(1778);
    layer1_outputs(2226) <= layer0_outputs(1553);
    layer1_outputs(2227) <= layer0_outputs(747);
    layer1_outputs(2228) <= (layer0_outputs(1533)) and (layer0_outputs(1683));
    layer1_outputs(2229) <= layer0_outputs(1891);
    layer1_outputs(2230) <= not(layer0_outputs(145));
    layer1_outputs(2231) <= (layer0_outputs(2150)) and (layer0_outputs(224));
    layer1_outputs(2232) <= not((layer0_outputs(1223)) and (layer0_outputs(1186)));
    layer1_outputs(2233) <= layer0_outputs(2204);
    layer1_outputs(2234) <= '1';
    layer1_outputs(2235) <= layer0_outputs(1829);
    layer1_outputs(2236) <= not((layer0_outputs(1612)) or (layer0_outputs(1758)));
    layer1_outputs(2237) <= layer0_outputs(459);
    layer1_outputs(2238) <= not(layer0_outputs(1511)) or (layer0_outputs(1769));
    layer1_outputs(2239) <= layer0_outputs(174);
    layer1_outputs(2240) <= layer0_outputs(2425);
    layer1_outputs(2241) <= (layer0_outputs(428)) and not (layer0_outputs(776));
    layer1_outputs(2242) <= (layer0_outputs(2080)) and not (layer0_outputs(764));
    layer1_outputs(2243) <= not(layer0_outputs(374));
    layer1_outputs(2244) <= (layer0_outputs(2147)) or (layer0_outputs(2145));
    layer1_outputs(2245) <= not(layer0_outputs(2315)) or (layer0_outputs(1482));
    layer1_outputs(2246) <= not(layer0_outputs(942)) or (layer0_outputs(1869));
    layer1_outputs(2247) <= not(layer0_outputs(2345));
    layer1_outputs(2248) <= layer0_outputs(2150);
    layer1_outputs(2249) <= (layer0_outputs(2296)) and (layer0_outputs(1074));
    layer1_outputs(2250) <= not(layer0_outputs(1834)) or (layer0_outputs(688));
    layer1_outputs(2251) <= not(layer0_outputs(1955)) or (layer0_outputs(1907));
    layer1_outputs(2252) <= (layer0_outputs(2141)) or (layer0_outputs(1242));
    layer1_outputs(2253) <= layer0_outputs(2500);
    layer1_outputs(2254) <= (layer0_outputs(470)) and not (layer0_outputs(689));
    layer1_outputs(2255) <= not(layer0_outputs(477)) or (layer0_outputs(2045));
    layer1_outputs(2256) <= not(layer0_outputs(1932)) or (layer0_outputs(411));
    layer1_outputs(2257) <= layer0_outputs(2021);
    layer1_outputs(2258) <= (layer0_outputs(1470)) and not (layer0_outputs(2270));
    layer1_outputs(2259) <= not((layer0_outputs(2213)) and (layer0_outputs(817)));
    layer1_outputs(2260) <= layer0_outputs(2220);
    layer1_outputs(2261) <= not(layer0_outputs(111)) or (layer0_outputs(2));
    layer1_outputs(2262) <= not(layer0_outputs(2459)) or (layer0_outputs(567));
    layer1_outputs(2263) <= (layer0_outputs(1468)) xor (layer0_outputs(2388));
    layer1_outputs(2264) <= '0';
    layer1_outputs(2265) <= not(layer0_outputs(4)) or (layer0_outputs(18));
    layer1_outputs(2266) <= '1';
    layer1_outputs(2267) <= not((layer0_outputs(1208)) xor (layer0_outputs(1357)));
    layer1_outputs(2268) <= (layer0_outputs(2394)) and (layer0_outputs(4));
    layer1_outputs(2269) <= layer0_outputs(2397);
    layer1_outputs(2270) <= '0';
    layer1_outputs(2271) <= (layer0_outputs(2443)) and (layer0_outputs(1812));
    layer1_outputs(2272) <= not(layer0_outputs(255)) or (layer0_outputs(705));
    layer1_outputs(2273) <= (layer0_outputs(1275)) and (layer0_outputs(647));
    layer1_outputs(2274) <= '1';
    layer1_outputs(2275) <= not((layer0_outputs(2315)) and (layer0_outputs(1712)));
    layer1_outputs(2276) <= (layer0_outputs(100)) or (layer0_outputs(620));
    layer1_outputs(2277) <= (layer0_outputs(2165)) or (layer0_outputs(1066));
    layer1_outputs(2278) <= not((layer0_outputs(2165)) xor (layer0_outputs(787)));
    layer1_outputs(2279) <= layer0_outputs(1205);
    layer1_outputs(2280) <= layer0_outputs(245);
    layer1_outputs(2281) <= (layer0_outputs(2283)) and not (layer0_outputs(2534));
    layer1_outputs(2282) <= (layer0_outputs(2490)) and (layer0_outputs(432));
    layer1_outputs(2283) <= (layer0_outputs(1257)) and (layer0_outputs(670));
    layer1_outputs(2284) <= (layer0_outputs(44)) or (layer0_outputs(368));
    layer1_outputs(2285) <= (layer0_outputs(2237)) xor (layer0_outputs(433));
    layer1_outputs(2286) <= not(layer0_outputs(122)) or (layer0_outputs(75));
    layer1_outputs(2287) <= layer0_outputs(831);
    layer1_outputs(2288) <= not(layer0_outputs(1495));
    layer1_outputs(2289) <= layer0_outputs(643);
    layer1_outputs(2290) <= not(layer0_outputs(169));
    layer1_outputs(2291) <= '0';
    layer1_outputs(2292) <= not((layer0_outputs(475)) and (layer0_outputs(1185)));
    layer1_outputs(2293) <= not((layer0_outputs(530)) or (layer0_outputs(1462)));
    layer1_outputs(2294) <= not(layer0_outputs(2217)) or (layer0_outputs(646));
    layer1_outputs(2295) <= layer0_outputs(1036);
    layer1_outputs(2296) <= not((layer0_outputs(625)) xor (layer0_outputs(1103)));
    layer1_outputs(2297) <= not((layer0_outputs(593)) and (layer0_outputs(804)));
    layer1_outputs(2298) <= not(layer0_outputs(979)) or (layer0_outputs(528));
    layer1_outputs(2299) <= not((layer0_outputs(576)) and (layer0_outputs(992)));
    layer1_outputs(2300) <= not(layer0_outputs(2166)) or (layer0_outputs(561));
    layer1_outputs(2301) <= not((layer0_outputs(1380)) or (layer0_outputs(2524)));
    layer1_outputs(2302) <= not(layer0_outputs(1133));
    layer1_outputs(2303) <= not((layer0_outputs(993)) or (layer0_outputs(37)));
    layer1_outputs(2304) <= not(layer0_outputs(2489));
    layer1_outputs(2305) <= '0';
    layer1_outputs(2306) <= not((layer0_outputs(310)) and (layer0_outputs(164)));
    layer1_outputs(2307) <= not(layer0_outputs(1493));
    layer1_outputs(2308) <= '1';
    layer1_outputs(2309) <= (layer0_outputs(1143)) and not (layer0_outputs(1177));
    layer1_outputs(2310) <= (layer0_outputs(1169)) or (layer0_outputs(1943));
    layer1_outputs(2311) <= (layer0_outputs(77)) and not (layer0_outputs(1792));
    layer1_outputs(2312) <= not(layer0_outputs(837)) or (layer0_outputs(2067));
    layer1_outputs(2313) <= layer0_outputs(1619);
    layer1_outputs(2314) <= (layer0_outputs(1666)) and (layer0_outputs(1691));
    layer1_outputs(2315) <= (layer0_outputs(1571)) or (layer0_outputs(156));
    layer1_outputs(2316) <= layer0_outputs(690);
    layer1_outputs(2317) <= not(layer0_outputs(1768)) or (layer0_outputs(663));
    layer1_outputs(2318) <= layer0_outputs(921);
    layer1_outputs(2319) <= layer0_outputs(556);
    layer1_outputs(2320) <= not((layer0_outputs(2155)) or (layer0_outputs(437)));
    layer1_outputs(2321) <= not(layer0_outputs(347));
    layer1_outputs(2322) <= (layer0_outputs(1224)) and (layer0_outputs(615));
    layer1_outputs(2323) <= not((layer0_outputs(1287)) and (layer0_outputs(1534)));
    layer1_outputs(2324) <= (layer0_outputs(103)) and not (layer0_outputs(2396));
    layer1_outputs(2325) <= not(layer0_outputs(1393)) or (layer0_outputs(339));
    layer1_outputs(2326) <= not((layer0_outputs(206)) or (layer0_outputs(1049)));
    layer1_outputs(2327) <= not(layer0_outputs(856));
    layer1_outputs(2328) <= not(layer0_outputs(2103)) or (layer0_outputs(396));
    layer1_outputs(2329) <= not((layer0_outputs(1786)) xor (layer0_outputs(1566)));
    layer1_outputs(2330) <= (layer0_outputs(2146)) or (layer0_outputs(1351));
    layer1_outputs(2331) <= layer0_outputs(699);
    layer1_outputs(2332) <= layer0_outputs(271);
    layer1_outputs(2333) <= (layer0_outputs(1804)) and not (layer0_outputs(1171));
    layer1_outputs(2334) <= not(layer0_outputs(512)) or (layer0_outputs(2245));
    layer1_outputs(2335) <= not((layer0_outputs(644)) or (layer0_outputs(2321)));
    layer1_outputs(2336) <= (layer0_outputs(2001)) and not (layer0_outputs(1760));
    layer1_outputs(2337) <= (layer0_outputs(187)) and not (layer0_outputs(2020));
    layer1_outputs(2338) <= layer0_outputs(1243);
    layer1_outputs(2339) <= layer0_outputs(2092);
    layer1_outputs(2340) <= '0';
    layer1_outputs(2341) <= '0';
    layer1_outputs(2342) <= not(layer0_outputs(2486));
    layer1_outputs(2343) <= not(layer0_outputs(2334));
    layer1_outputs(2344) <= '0';
    layer1_outputs(2345) <= layer0_outputs(17);
    layer1_outputs(2346) <= not((layer0_outputs(1821)) and (layer0_outputs(581)));
    layer1_outputs(2347) <= '0';
    layer1_outputs(2348) <= layer0_outputs(236);
    layer1_outputs(2349) <= not(layer0_outputs(2541)) or (layer0_outputs(1956));
    layer1_outputs(2350) <= not(layer0_outputs(1799));
    layer1_outputs(2351) <= (layer0_outputs(423)) and not (layer0_outputs(2515));
    layer1_outputs(2352) <= not(layer0_outputs(2473));
    layer1_outputs(2353) <= layer0_outputs(1999);
    layer1_outputs(2354) <= (layer0_outputs(1331)) and not (layer0_outputs(1614));
    layer1_outputs(2355) <= (layer0_outputs(453)) and (layer0_outputs(664));
    layer1_outputs(2356) <= layer0_outputs(481);
    layer1_outputs(2357) <= not((layer0_outputs(392)) or (layer0_outputs(1660)));
    layer1_outputs(2358) <= layer0_outputs(2129);
    layer1_outputs(2359) <= '0';
    layer1_outputs(2360) <= (layer0_outputs(2174)) or (layer0_outputs(456));
    layer1_outputs(2361) <= '0';
    layer1_outputs(2362) <= (layer0_outputs(1002)) xor (layer0_outputs(1820));
    layer1_outputs(2363) <= layer0_outputs(2361);
    layer1_outputs(2364) <= not((layer0_outputs(2484)) and (layer0_outputs(1987)));
    layer1_outputs(2365) <= not(layer0_outputs(395));
    layer1_outputs(2366) <= layer0_outputs(212);
    layer1_outputs(2367) <= (layer0_outputs(889)) and (layer0_outputs(972));
    layer1_outputs(2368) <= (layer0_outputs(2460)) and not (layer0_outputs(571));
    layer1_outputs(2369) <= not(layer0_outputs(744)) or (layer0_outputs(1673));
    layer1_outputs(2370) <= layer0_outputs(2408);
    layer1_outputs(2371) <= layer0_outputs(262);
    layer1_outputs(2372) <= layer0_outputs(2417);
    layer1_outputs(2373) <= not((layer0_outputs(63)) or (layer0_outputs(821)));
    layer1_outputs(2374) <= not(layer0_outputs(1609));
    layer1_outputs(2375) <= layer0_outputs(1238);
    layer1_outputs(2376) <= not(layer0_outputs(2084));
    layer1_outputs(2377) <= '0';
    layer1_outputs(2378) <= not(layer0_outputs(425)) or (layer0_outputs(548));
    layer1_outputs(2379) <= layer0_outputs(1880);
    layer1_outputs(2380) <= not(layer0_outputs(463)) or (layer0_outputs(128));
    layer1_outputs(2381) <= not((layer0_outputs(1347)) or (layer0_outputs(198)));
    layer1_outputs(2382) <= (layer0_outputs(958)) or (layer0_outputs(2528));
    layer1_outputs(2383) <= layer0_outputs(136);
    layer1_outputs(2384) <= (layer0_outputs(1396)) or (layer0_outputs(1438));
    layer1_outputs(2385) <= not(layer0_outputs(274));
    layer1_outputs(2386) <= not(layer0_outputs(1132)) or (layer0_outputs(464));
    layer1_outputs(2387) <= not(layer0_outputs(561));
    layer1_outputs(2388) <= not(layer0_outputs(196));
    layer1_outputs(2389) <= not(layer0_outputs(592));
    layer1_outputs(2390) <= layer0_outputs(1071);
    layer1_outputs(2391) <= (layer0_outputs(1634)) and (layer0_outputs(2360));
    layer1_outputs(2392) <= (layer0_outputs(717)) and not (layer0_outputs(2184));
    layer1_outputs(2393) <= layer0_outputs(2424);
    layer1_outputs(2394) <= layer0_outputs(394);
    layer1_outputs(2395) <= not((layer0_outputs(2424)) and (layer0_outputs(1362)));
    layer1_outputs(2396) <= (layer0_outputs(2221)) and (layer0_outputs(2282));
    layer1_outputs(2397) <= layer0_outputs(180);
    layer1_outputs(2398) <= (layer0_outputs(2162)) and not (layer0_outputs(56));
    layer1_outputs(2399) <= layer0_outputs(496);
    layer1_outputs(2400) <= '0';
    layer1_outputs(2401) <= not(layer0_outputs(1143)) or (layer0_outputs(2289));
    layer1_outputs(2402) <= layer0_outputs(1273);
    layer1_outputs(2403) <= '1';
    layer1_outputs(2404) <= (layer0_outputs(1732)) xor (layer0_outputs(481));
    layer1_outputs(2405) <= not((layer0_outputs(1564)) or (layer0_outputs(1702)));
    layer1_outputs(2406) <= (layer0_outputs(1336)) and (layer0_outputs(1884));
    layer1_outputs(2407) <= (layer0_outputs(609)) and not (layer0_outputs(2479));
    layer1_outputs(2408) <= not(layer0_outputs(1800));
    layer1_outputs(2409) <= layer0_outputs(349);
    layer1_outputs(2410) <= (layer0_outputs(2455)) or (layer0_outputs(1230));
    layer1_outputs(2411) <= not(layer0_outputs(1852));
    layer1_outputs(2412) <= (layer0_outputs(1883)) and (layer0_outputs(1329));
    layer1_outputs(2413) <= (layer0_outputs(2077)) and not (layer0_outputs(298));
    layer1_outputs(2414) <= layer0_outputs(1546);
    layer1_outputs(2415) <= '1';
    layer1_outputs(2416) <= (layer0_outputs(1988)) and not (layer0_outputs(489));
    layer1_outputs(2417) <= not(layer0_outputs(1341));
    layer1_outputs(2418) <= not(layer0_outputs(661)) or (layer0_outputs(1544));
    layer1_outputs(2419) <= (layer0_outputs(684)) or (layer0_outputs(233));
    layer1_outputs(2420) <= (layer0_outputs(1795)) and not (layer0_outputs(2063));
    layer1_outputs(2421) <= not(layer0_outputs(603)) or (layer0_outputs(1281));
    layer1_outputs(2422) <= not(layer0_outputs(202)) or (layer0_outputs(1050));
    layer1_outputs(2423) <= layer0_outputs(56);
    layer1_outputs(2424) <= not(layer0_outputs(509)) or (layer0_outputs(970));
    layer1_outputs(2425) <= (layer0_outputs(423)) and (layer0_outputs(549));
    layer1_outputs(2426) <= (layer0_outputs(2483)) and not (layer0_outputs(51));
    layer1_outputs(2427) <= (layer0_outputs(2509)) and (layer0_outputs(2209));
    layer1_outputs(2428) <= not(layer0_outputs(2419)) or (layer0_outputs(631));
    layer1_outputs(2429) <= not((layer0_outputs(2060)) or (layer0_outputs(26)));
    layer1_outputs(2430) <= '1';
    layer1_outputs(2431) <= layer0_outputs(1112);
    layer1_outputs(2432) <= (layer0_outputs(434)) and (layer0_outputs(1222));
    layer1_outputs(2433) <= (layer0_outputs(469)) and not (layer0_outputs(1101));
    layer1_outputs(2434) <= not((layer0_outputs(329)) and (layer0_outputs(749)));
    layer1_outputs(2435) <= layer0_outputs(2422);
    layer1_outputs(2436) <= layer0_outputs(1605);
    layer1_outputs(2437) <= (layer0_outputs(2088)) and (layer0_outputs(2036));
    layer1_outputs(2438) <= layer0_outputs(987);
    layer1_outputs(2439) <= '1';
    layer1_outputs(2440) <= not(layer0_outputs(555));
    layer1_outputs(2441) <= (layer0_outputs(974)) and (layer0_outputs(165));
    layer1_outputs(2442) <= (layer0_outputs(1963)) and (layer0_outputs(641));
    layer1_outputs(2443) <= not((layer0_outputs(1900)) or (layer0_outputs(1881)));
    layer1_outputs(2444) <= (layer0_outputs(1893)) or (layer0_outputs(65));
    layer1_outputs(2445) <= (layer0_outputs(587)) and not (layer0_outputs(1692));
    layer1_outputs(2446) <= not((layer0_outputs(1306)) and (layer0_outputs(742)));
    layer1_outputs(2447) <= not(layer0_outputs(322)) or (layer0_outputs(543));
    layer1_outputs(2448) <= not(layer0_outputs(1259)) or (layer0_outputs(2026));
    layer1_outputs(2449) <= not(layer0_outputs(2323));
    layer1_outputs(2450) <= not((layer0_outputs(2350)) or (layer0_outputs(2126)));
    layer1_outputs(2451) <= (layer0_outputs(627)) and (layer0_outputs(1454));
    layer1_outputs(2452) <= not(layer0_outputs(742));
    layer1_outputs(2453) <= layer0_outputs(2187);
    layer1_outputs(2454) <= not(layer0_outputs(1411));
    layer1_outputs(2455) <= not(layer0_outputs(1860));
    layer1_outputs(2456) <= (layer0_outputs(1142)) or (layer0_outputs(549));
    layer1_outputs(2457) <= not(layer0_outputs(638));
    layer1_outputs(2458) <= layer0_outputs(352);
    layer1_outputs(2459) <= (layer0_outputs(1857)) or (layer0_outputs(1509));
    layer1_outputs(2460) <= layer0_outputs(1028);
    layer1_outputs(2461) <= not(layer0_outputs(1332));
    layer1_outputs(2462) <= (layer0_outputs(529)) and not (layer0_outputs(1061));
    layer1_outputs(2463) <= '1';
    layer1_outputs(2464) <= layer0_outputs(231);
    layer1_outputs(2465) <= layer0_outputs(618);
    layer1_outputs(2466) <= (layer0_outputs(2136)) and not (layer0_outputs(1147));
    layer1_outputs(2467) <= not(layer0_outputs(1581)) or (layer0_outputs(667));
    layer1_outputs(2468) <= not(layer0_outputs(1531));
    layer1_outputs(2469) <= not((layer0_outputs(69)) and (layer0_outputs(1913)));
    layer1_outputs(2470) <= '1';
    layer1_outputs(2471) <= not(layer0_outputs(851));
    layer1_outputs(2472) <= layer0_outputs(1779);
    layer1_outputs(2473) <= layer0_outputs(1078);
    layer1_outputs(2474) <= (layer0_outputs(2253)) or (layer0_outputs(360));
    layer1_outputs(2475) <= not(layer0_outputs(1664));
    layer1_outputs(2476) <= layer0_outputs(2439);
    layer1_outputs(2477) <= (layer0_outputs(168)) and not (layer0_outputs(0));
    layer1_outputs(2478) <= (layer0_outputs(1675)) or (layer0_outputs(915));
    layer1_outputs(2479) <= not(layer0_outputs(1996));
    layer1_outputs(2480) <= not(layer0_outputs(1916)) or (layer0_outputs(2040));
    layer1_outputs(2481) <= (layer0_outputs(1941)) or (layer0_outputs(625));
    layer1_outputs(2482) <= layer0_outputs(314);
    layer1_outputs(2483) <= not(layer0_outputs(1860)) or (layer0_outputs(1999));
    layer1_outputs(2484) <= not((layer0_outputs(2462)) and (layer0_outputs(2435)));
    layer1_outputs(2485) <= not((layer0_outputs(918)) and (layer0_outputs(524)));
    layer1_outputs(2486) <= not((layer0_outputs(1041)) or (layer0_outputs(1541)));
    layer1_outputs(2487) <= layer0_outputs(287);
    layer1_outputs(2488) <= not(layer0_outputs(1302));
    layer1_outputs(2489) <= layer0_outputs(1172);
    layer1_outputs(2490) <= (layer0_outputs(2318)) or (layer0_outputs(1567));
    layer1_outputs(2491) <= not(layer0_outputs(1799));
    layer1_outputs(2492) <= layer0_outputs(2336);
    layer1_outputs(2493) <= (layer0_outputs(1058)) and (layer0_outputs(2395));
    layer1_outputs(2494) <= (layer0_outputs(1073)) and not (layer0_outputs(2032));
    layer1_outputs(2495) <= not(layer0_outputs(709));
    layer1_outputs(2496) <= (layer0_outputs(1809)) and not (layer0_outputs(1543));
    layer1_outputs(2497) <= (layer0_outputs(181)) and not (layer0_outputs(2442));
    layer1_outputs(2498) <= layer0_outputs(153);
    layer1_outputs(2499) <= not(layer0_outputs(533));
    layer1_outputs(2500) <= not(layer0_outputs(442)) or (layer0_outputs(1272));
    layer1_outputs(2501) <= '0';
    layer1_outputs(2502) <= layer0_outputs(2399);
    layer1_outputs(2503) <= '0';
    layer1_outputs(2504) <= not(layer0_outputs(1360));
    layer1_outputs(2505) <= layer0_outputs(2437);
    layer1_outputs(2506) <= layer0_outputs(480);
    layer1_outputs(2507) <= not(layer0_outputs(1600));
    layer1_outputs(2508) <= not(layer0_outputs(870)) or (layer0_outputs(1916));
    layer1_outputs(2509) <= layer0_outputs(1614);
    layer1_outputs(2510) <= not((layer0_outputs(1875)) and (layer0_outputs(1978)));
    layer1_outputs(2511) <= not(layer0_outputs(254)) or (layer0_outputs(2428));
    layer1_outputs(2512) <= layer0_outputs(1165);
    layer1_outputs(2513) <= (layer0_outputs(1360)) and (layer0_outputs(2540));
    layer1_outputs(2514) <= not((layer0_outputs(2221)) xor (layer0_outputs(1003)));
    layer1_outputs(2515) <= layer0_outputs(1885);
    layer1_outputs(2516) <= (layer0_outputs(2524)) or (layer0_outputs(937));
    layer1_outputs(2517) <= layer0_outputs(33);
    layer1_outputs(2518) <= (layer0_outputs(547)) and not (layer0_outputs(26));
    layer1_outputs(2519) <= not((layer0_outputs(2262)) or (layer0_outputs(1639)));
    layer1_outputs(2520) <= not(layer0_outputs(1167));
    layer1_outputs(2521) <= not(layer0_outputs(537));
    layer1_outputs(2522) <= not((layer0_outputs(928)) or (layer0_outputs(454)));
    layer1_outputs(2523) <= (layer0_outputs(117)) and not (layer0_outputs(1264));
    layer1_outputs(2524) <= not(layer0_outputs(2190));
    layer1_outputs(2525) <= (layer0_outputs(1492)) and not (layer0_outputs(409));
    layer1_outputs(2526) <= not((layer0_outputs(1204)) or (layer0_outputs(2457)));
    layer1_outputs(2527) <= (layer0_outputs(1807)) and not (layer0_outputs(1407));
    layer1_outputs(2528) <= not(layer0_outputs(463));
    layer1_outputs(2529) <= not(layer0_outputs(546));
    layer1_outputs(2530) <= not(layer0_outputs(2011)) or (layer0_outputs(698));
    layer1_outputs(2531) <= layer0_outputs(1646);
    layer1_outputs(2532) <= (layer0_outputs(204)) and not (layer0_outputs(2537));
    layer1_outputs(2533) <= (layer0_outputs(1861)) and not (layer0_outputs(897));
    layer1_outputs(2534) <= not((layer0_outputs(855)) and (layer0_outputs(1151)));
    layer1_outputs(2535) <= (layer0_outputs(1067)) and not (layer0_outputs(334));
    layer1_outputs(2536) <= layer0_outputs(658);
    layer1_outputs(2537) <= (layer0_outputs(2446)) and not (layer0_outputs(502));
    layer1_outputs(2538) <= (layer0_outputs(445)) and (layer0_outputs(2104));
    layer1_outputs(2539) <= layer0_outputs(2012);
    layer1_outputs(2540) <= not(layer0_outputs(2301)) or (layer0_outputs(1766));
    layer1_outputs(2541) <= (layer0_outputs(2364)) and not (layer0_outputs(1180));
    layer1_outputs(2542) <= layer0_outputs(565);
    layer1_outputs(2543) <= not(layer0_outputs(2214)) or (layer0_outputs(215));
    layer1_outputs(2544) <= not((layer0_outputs(2489)) or (layer0_outputs(2518)));
    layer1_outputs(2545) <= (layer0_outputs(2201)) and not (layer0_outputs(2108));
    layer1_outputs(2546) <= not((layer0_outputs(1998)) or (layer0_outputs(2206)));
    layer1_outputs(2547) <= not(layer0_outputs(803));
    layer1_outputs(2548) <= (layer0_outputs(1400)) or (layer0_outputs(46));
    layer1_outputs(2549) <= layer0_outputs(2410);
    layer1_outputs(2550) <= (layer0_outputs(152)) and (layer0_outputs(2151));
    layer1_outputs(2551) <= not(layer0_outputs(801));
    layer1_outputs(2552) <= not(layer0_outputs(894));
    layer1_outputs(2553) <= not(layer0_outputs(1284));
    layer1_outputs(2554) <= not((layer0_outputs(1381)) or (layer0_outputs(2087)));
    layer1_outputs(2555) <= not(layer0_outputs(2148)) or (layer0_outputs(2132));
    layer1_outputs(2556) <= not(layer0_outputs(2405));
    layer1_outputs(2557) <= not(layer0_outputs(2290));
    layer1_outputs(2558) <= not(layer0_outputs(793));
    layer1_outputs(2559) <= (layer0_outputs(2340)) or (layer0_outputs(743));
    layer2_outputs(0) <= not(layer1_outputs(221));
    layer2_outputs(1) <= layer1_outputs(2093);
    layer2_outputs(2) <= not(layer1_outputs(2337));
    layer2_outputs(3) <= not(layer1_outputs(805));
    layer2_outputs(4) <= (layer1_outputs(1197)) and (layer1_outputs(963));
    layer2_outputs(5) <= not(layer1_outputs(1982)) or (layer1_outputs(1269));
    layer2_outputs(6) <= not((layer1_outputs(1780)) and (layer1_outputs(873)));
    layer2_outputs(7) <= '1';
    layer2_outputs(8) <= not(layer1_outputs(1169)) or (layer1_outputs(149));
    layer2_outputs(9) <= not(layer1_outputs(1581)) or (layer1_outputs(1614));
    layer2_outputs(10) <= not(layer1_outputs(859));
    layer2_outputs(11) <= layer1_outputs(438);
    layer2_outputs(12) <= not(layer1_outputs(929));
    layer2_outputs(13) <= (layer1_outputs(531)) or (layer1_outputs(2183));
    layer2_outputs(14) <= layer1_outputs(933);
    layer2_outputs(15) <= (layer1_outputs(430)) and not (layer1_outputs(1647));
    layer2_outputs(16) <= not(layer1_outputs(0)) or (layer1_outputs(1997));
    layer2_outputs(17) <= not((layer1_outputs(2341)) and (layer1_outputs(715)));
    layer2_outputs(18) <= (layer1_outputs(1645)) and not (layer1_outputs(1553));
    layer2_outputs(19) <= (layer1_outputs(50)) and (layer1_outputs(2233));
    layer2_outputs(20) <= not(layer1_outputs(1042));
    layer2_outputs(21) <= layer1_outputs(1176);
    layer2_outputs(22) <= layer1_outputs(1213);
    layer2_outputs(23) <= not(layer1_outputs(1451)) or (layer1_outputs(2420));
    layer2_outputs(24) <= layer1_outputs(669);
    layer2_outputs(25) <= (layer1_outputs(802)) or (layer1_outputs(2295));
    layer2_outputs(26) <= '1';
    layer2_outputs(27) <= (layer1_outputs(2299)) and not (layer1_outputs(569));
    layer2_outputs(28) <= (layer1_outputs(888)) or (layer1_outputs(890));
    layer2_outputs(29) <= (layer1_outputs(1737)) and (layer1_outputs(951));
    layer2_outputs(30) <= not(layer1_outputs(886));
    layer2_outputs(31) <= not(layer1_outputs(2255)) or (layer1_outputs(1774));
    layer2_outputs(32) <= layer1_outputs(558);
    layer2_outputs(33) <= '0';
    layer2_outputs(34) <= (layer1_outputs(2400)) and not (layer1_outputs(2234));
    layer2_outputs(35) <= not(layer1_outputs(1277)) or (layer1_outputs(2046));
    layer2_outputs(36) <= layer1_outputs(173);
    layer2_outputs(37) <= not(layer1_outputs(1594));
    layer2_outputs(38) <= not(layer1_outputs(1056));
    layer2_outputs(39) <= layer1_outputs(2548);
    layer2_outputs(40) <= (layer1_outputs(1304)) and not (layer1_outputs(849));
    layer2_outputs(41) <= (layer1_outputs(1108)) or (layer1_outputs(2425));
    layer2_outputs(42) <= (layer1_outputs(1968)) and (layer1_outputs(962));
    layer2_outputs(43) <= not(layer1_outputs(1690));
    layer2_outputs(44) <= not(layer1_outputs(495)) or (layer1_outputs(770));
    layer2_outputs(45) <= not(layer1_outputs(1622));
    layer2_outputs(46) <= not(layer1_outputs(1350)) or (layer1_outputs(2141));
    layer2_outputs(47) <= (layer1_outputs(2297)) and not (layer1_outputs(825));
    layer2_outputs(48) <= (layer1_outputs(172)) and not (layer1_outputs(294));
    layer2_outputs(49) <= (layer1_outputs(1917)) or (layer1_outputs(2144));
    layer2_outputs(50) <= (layer1_outputs(637)) and (layer1_outputs(1358));
    layer2_outputs(51) <= (layer1_outputs(107)) and not (layer1_outputs(2295));
    layer2_outputs(52) <= (layer1_outputs(2387)) or (layer1_outputs(1252));
    layer2_outputs(53) <= layer1_outputs(2453);
    layer2_outputs(54) <= not(layer1_outputs(882)) or (layer1_outputs(628));
    layer2_outputs(55) <= not(layer1_outputs(598));
    layer2_outputs(56) <= (layer1_outputs(2294)) and not (layer1_outputs(491));
    layer2_outputs(57) <= layer1_outputs(1079);
    layer2_outputs(58) <= (layer1_outputs(1623)) and not (layer1_outputs(2172));
    layer2_outputs(59) <= layer1_outputs(2187);
    layer2_outputs(60) <= not(layer1_outputs(124));
    layer2_outputs(61) <= layer1_outputs(97);
    layer2_outputs(62) <= (layer1_outputs(2420)) and not (layer1_outputs(795));
    layer2_outputs(63) <= layer1_outputs(2257);
    layer2_outputs(64) <= (layer1_outputs(1342)) and (layer1_outputs(1178));
    layer2_outputs(65) <= (layer1_outputs(63)) or (layer1_outputs(1736));
    layer2_outputs(66) <= layer1_outputs(2481);
    layer2_outputs(67) <= not((layer1_outputs(926)) xor (layer1_outputs(813)));
    layer2_outputs(68) <= not(layer1_outputs(1157));
    layer2_outputs(69) <= not(layer1_outputs(860));
    layer2_outputs(70) <= not((layer1_outputs(703)) and (layer1_outputs(366)));
    layer2_outputs(71) <= not(layer1_outputs(80));
    layer2_outputs(72) <= (layer1_outputs(377)) xor (layer1_outputs(1938));
    layer2_outputs(73) <= not(layer1_outputs(1780)) or (layer1_outputs(93));
    layer2_outputs(74) <= (layer1_outputs(1407)) or (layer1_outputs(2315));
    layer2_outputs(75) <= not((layer1_outputs(81)) and (layer1_outputs(2178)));
    layer2_outputs(76) <= not(layer1_outputs(1192)) or (layer1_outputs(1479));
    layer2_outputs(77) <= not(layer1_outputs(446)) or (layer1_outputs(2248));
    layer2_outputs(78) <= not(layer1_outputs(194)) or (layer1_outputs(547));
    layer2_outputs(79) <= not(layer1_outputs(2406)) or (layer1_outputs(586));
    layer2_outputs(80) <= layer1_outputs(2379);
    layer2_outputs(81) <= not(layer1_outputs(1073));
    layer2_outputs(82) <= not(layer1_outputs(1690)) or (layer1_outputs(914));
    layer2_outputs(83) <= (layer1_outputs(1417)) and (layer1_outputs(1319));
    layer2_outputs(84) <= layer1_outputs(1374);
    layer2_outputs(85) <= (layer1_outputs(944)) and (layer1_outputs(102));
    layer2_outputs(86) <= layer1_outputs(857);
    layer2_outputs(87) <= not(layer1_outputs(1612));
    layer2_outputs(88) <= (layer1_outputs(1466)) and not (layer1_outputs(1978));
    layer2_outputs(89) <= layer1_outputs(1922);
    layer2_outputs(90) <= (layer1_outputs(260)) and (layer1_outputs(1289));
    layer2_outputs(91) <= layer1_outputs(424);
    layer2_outputs(92) <= (layer1_outputs(1959)) or (layer1_outputs(1315));
    layer2_outputs(93) <= not(layer1_outputs(122));
    layer2_outputs(94) <= not(layer1_outputs(2196));
    layer2_outputs(95) <= not((layer1_outputs(2036)) and (layer1_outputs(1362)));
    layer2_outputs(96) <= '1';
    layer2_outputs(97) <= (layer1_outputs(2268)) or (layer1_outputs(2070));
    layer2_outputs(98) <= (layer1_outputs(387)) and not (layer1_outputs(89));
    layer2_outputs(99) <= layer1_outputs(1482);
    layer2_outputs(100) <= not(layer1_outputs(2143));
    layer2_outputs(101) <= not(layer1_outputs(632));
    layer2_outputs(102) <= not(layer1_outputs(111));
    layer2_outputs(103) <= (layer1_outputs(957)) and not (layer1_outputs(610));
    layer2_outputs(104) <= (layer1_outputs(343)) or (layer1_outputs(208));
    layer2_outputs(105) <= not(layer1_outputs(1093)) or (layer1_outputs(1503));
    layer2_outputs(106) <= layer1_outputs(2328);
    layer2_outputs(107) <= not(layer1_outputs(1812)) or (layer1_outputs(1905));
    layer2_outputs(108) <= not(layer1_outputs(1704));
    layer2_outputs(109) <= (layer1_outputs(179)) and (layer1_outputs(1263));
    layer2_outputs(110) <= not(layer1_outputs(2343));
    layer2_outputs(111) <= layer1_outputs(2547);
    layer2_outputs(112) <= not((layer1_outputs(539)) or (layer1_outputs(521)));
    layer2_outputs(113) <= layer1_outputs(990);
    layer2_outputs(114) <= '1';
    layer2_outputs(115) <= not(layer1_outputs(501)) or (layer1_outputs(1245));
    layer2_outputs(116) <= (layer1_outputs(1913)) and not (layer1_outputs(1890));
    layer2_outputs(117) <= not((layer1_outputs(425)) and (layer1_outputs(754)));
    layer2_outputs(118) <= not(layer1_outputs(1797));
    layer2_outputs(119) <= (layer1_outputs(287)) and not (layer1_outputs(1083));
    layer2_outputs(120) <= not(layer1_outputs(2256));
    layer2_outputs(121) <= not(layer1_outputs(905));
    layer2_outputs(122) <= layer1_outputs(1589);
    layer2_outputs(123) <= not(layer1_outputs(884));
    layer2_outputs(124) <= not(layer1_outputs(585));
    layer2_outputs(125) <= not(layer1_outputs(671)) or (layer1_outputs(1645));
    layer2_outputs(126) <= not(layer1_outputs(897)) or (layer1_outputs(2057));
    layer2_outputs(127) <= not((layer1_outputs(453)) or (layer1_outputs(185)));
    layer2_outputs(128) <= layer1_outputs(2051);
    layer2_outputs(129) <= layer1_outputs(1843);
    layer2_outputs(130) <= not((layer1_outputs(809)) and (layer1_outputs(1732)));
    layer2_outputs(131) <= not((layer1_outputs(1187)) or (layer1_outputs(794)));
    layer2_outputs(132) <= layer1_outputs(1276);
    layer2_outputs(133) <= not((layer1_outputs(234)) and (layer1_outputs(846)));
    layer2_outputs(134) <= (layer1_outputs(1668)) and (layer1_outputs(519));
    layer2_outputs(135) <= layer1_outputs(2472);
    layer2_outputs(136) <= not(layer1_outputs(267));
    layer2_outputs(137) <= not(layer1_outputs(2552));
    layer2_outputs(138) <= not(layer1_outputs(738));
    layer2_outputs(139) <= not(layer1_outputs(2465));
    layer2_outputs(140) <= layer1_outputs(2411);
    layer2_outputs(141) <= not((layer1_outputs(1786)) or (layer1_outputs(1080)));
    layer2_outputs(142) <= '1';
    layer2_outputs(143) <= layer1_outputs(971);
    layer2_outputs(144) <= not(layer1_outputs(282));
    layer2_outputs(145) <= layer1_outputs(773);
    layer2_outputs(146) <= not(layer1_outputs(2350));
    layer2_outputs(147) <= not(layer1_outputs(92));
    layer2_outputs(148) <= (layer1_outputs(1335)) or (layer1_outputs(844));
    layer2_outputs(149) <= '1';
    layer2_outputs(150) <= layer1_outputs(2127);
    layer2_outputs(151) <= (layer1_outputs(1979)) and not (layer1_outputs(496));
    layer2_outputs(152) <= (layer1_outputs(2275)) and not (layer1_outputs(1449));
    layer2_outputs(153) <= '0';
    layer2_outputs(154) <= not(layer1_outputs(566));
    layer2_outputs(155) <= not((layer1_outputs(721)) and (layer1_outputs(1811)));
    layer2_outputs(156) <= layer1_outputs(1746);
    layer2_outputs(157) <= (layer1_outputs(793)) and not (layer1_outputs(2079));
    layer2_outputs(158) <= layer1_outputs(1393);
    layer2_outputs(159) <= not(layer1_outputs(27));
    layer2_outputs(160) <= layer1_outputs(1846);
    layer2_outputs(161) <= not(layer1_outputs(2253));
    layer2_outputs(162) <= not((layer1_outputs(2207)) and (layer1_outputs(1010)));
    layer2_outputs(163) <= layer1_outputs(1430);
    layer2_outputs(164) <= not(layer1_outputs(1026));
    layer2_outputs(165) <= not(layer1_outputs(2351));
    layer2_outputs(166) <= '0';
    layer2_outputs(167) <= layer1_outputs(576);
    layer2_outputs(168) <= layer1_outputs(1762);
    layer2_outputs(169) <= not(layer1_outputs(918));
    layer2_outputs(170) <= not(layer1_outputs(572));
    layer2_outputs(171) <= layer1_outputs(606);
    layer2_outputs(172) <= not(layer1_outputs(548));
    layer2_outputs(173) <= (layer1_outputs(1534)) and not (layer1_outputs(1392));
    layer2_outputs(174) <= (layer1_outputs(2182)) or (layer1_outputs(126));
    layer2_outputs(175) <= not((layer1_outputs(2493)) or (layer1_outputs(2283)));
    layer2_outputs(176) <= '0';
    layer2_outputs(177) <= (layer1_outputs(39)) and not (layer1_outputs(1326));
    layer2_outputs(178) <= layer1_outputs(2539);
    layer2_outputs(179) <= layer1_outputs(1919);
    layer2_outputs(180) <= (layer1_outputs(452)) and not (layer1_outputs(48));
    layer2_outputs(181) <= not(layer1_outputs(1518));
    layer2_outputs(182) <= layer1_outputs(1330);
    layer2_outputs(183) <= '1';
    layer2_outputs(184) <= not((layer1_outputs(885)) xor (layer1_outputs(800)));
    layer2_outputs(185) <= layer1_outputs(1375);
    layer2_outputs(186) <= not(layer1_outputs(2375)) or (layer1_outputs(484));
    layer2_outputs(187) <= not(layer1_outputs(1551));
    layer2_outputs(188) <= not(layer1_outputs(1152)) or (layer1_outputs(58));
    layer2_outputs(189) <= not(layer1_outputs(123));
    layer2_outputs(190) <= (layer1_outputs(396)) and (layer1_outputs(1364));
    layer2_outputs(191) <= not((layer1_outputs(864)) and (layer1_outputs(1019)));
    layer2_outputs(192) <= layer1_outputs(900);
    layer2_outputs(193) <= not((layer1_outputs(497)) and (layer1_outputs(701)));
    layer2_outputs(194) <= (layer1_outputs(722)) and (layer1_outputs(233));
    layer2_outputs(195) <= (layer1_outputs(2353)) xor (layer1_outputs(706));
    layer2_outputs(196) <= not(layer1_outputs(1439)) or (layer1_outputs(2007));
    layer2_outputs(197) <= (layer1_outputs(327)) and not (layer1_outputs(2013));
    layer2_outputs(198) <= (layer1_outputs(2544)) or (layer1_outputs(1982));
    layer2_outputs(199) <= '1';
    layer2_outputs(200) <= (layer1_outputs(716)) and (layer1_outputs(390));
    layer2_outputs(201) <= not(layer1_outputs(1498)) or (layer1_outputs(2270));
    layer2_outputs(202) <= not((layer1_outputs(1693)) or (layer1_outputs(564)));
    layer2_outputs(203) <= (layer1_outputs(2128)) xor (layer1_outputs(1751));
    layer2_outputs(204) <= not((layer1_outputs(1579)) or (layer1_outputs(2084)));
    layer2_outputs(205) <= layer1_outputs(1702);
    layer2_outputs(206) <= not(layer1_outputs(1801));
    layer2_outputs(207) <= not(layer1_outputs(1714)) or (layer1_outputs(2504));
    layer2_outputs(208) <= not((layer1_outputs(2203)) or (layer1_outputs(1275)));
    layer2_outputs(209) <= not(layer1_outputs(1980)) or (layer1_outputs(1929));
    layer2_outputs(210) <= (layer1_outputs(40)) and not (layer1_outputs(1573));
    layer2_outputs(211) <= not(layer1_outputs(553));
    layer2_outputs(212) <= not((layer1_outputs(2510)) and (layer1_outputs(1064)));
    layer2_outputs(213) <= not(layer1_outputs(1604));
    layer2_outputs(214) <= not(layer1_outputs(2259));
    layer2_outputs(215) <= not((layer1_outputs(925)) or (layer1_outputs(1437)));
    layer2_outputs(216) <= layer1_outputs(901);
    layer2_outputs(217) <= layer1_outputs(256);
    layer2_outputs(218) <= (layer1_outputs(134)) and (layer1_outputs(136));
    layer2_outputs(219) <= not(layer1_outputs(1214));
    layer2_outputs(220) <= '0';
    layer2_outputs(221) <= not((layer1_outputs(108)) or (layer1_outputs(1562)));
    layer2_outputs(222) <= layer1_outputs(1302);
    layer2_outputs(223) <= layer1_outputs(2096);
    layer2_outputs(224) <= (layer1_outputs(1904)) and (layer1_outputs(1831));
    layer2_outputs(225) <= not((layer1_outputs(1775)) or (layer1_outputs(2555)));
    layer2_outputs(226) <= layer1_outputs(440);
    layer2_outputs(227) <= layer1_outputs(1921);
    layer2_outputs(228) <= (layer1_outputs(67)) and not (layer1_outputs(1892));
    layer2_outputs(229) <= not(layer1_outputs(2044)) or (layer1_outputs(2034));
    layer2_outputs(230) <= (layer1_outputs(1270)) and (layer1_outputs(1181));
    layer2_outputs(231) <= not(layer1_outputs(1957)) or (layer1_outputs(1321));
    layer2_outputs(232) <= layer1_outputs(292);
    layer2_outputs(233) <= not(layer1_outputs(34));
    layer2_outputs(234) <= not(layer1_outputs(673));
    layer2_outputs(235) <= not(layer1_outputs(2243));
    layer2_outputs(236) <= layer1_outputs(192);
    layer2_outputs(237) <= not(layer1_outputs(1248)) or (layer1_outputs(1790));
    layer2_outputs(238) <= (layer1_outputs(415)) and (layer1_outputs(2373));
    layer2_outputs(239) <= layer1_outputs(1101);
    layer2_outputs(240) <= (layer1_outputs(865)) and (layer1_outputs(2433));
    layer2_outputs(241) <= not((layer1_outputs(1234)) or (layer1_outputs(2288)));
    layer2_outputs(242) <= layer1_outputs(1601);
    layer2_outputs(243) <= not((layer1_outputs(1896)) or (layer1_outputs(2178)));
    layer2_outputs(244) <= not(layer1_outputs(2191));
    layer2_outputs(245) <= not(layer1_outputs(832)) or (layer1_outputs(237));
    layer2_outputs(246) <= not((layer1_outputs(1251)) and (layer1_outputs(2055)));
    layer2_outputs(247) <= not(layer1_outputs(1535)) or (layer1_outputs(1679));
    layer2_outputs(248) <= layer1_outputs(1677);
    layer2_outputs(249) <= '0';
    layer2_outputs(250) <= not(layer1_outputs(1183)) or (layer1_outputs(1776));
    layer2_outputs(251) <= not(layer1_outputs(392));
    layer2_outputs(252) <= not(layer1_outputs(1569)) or (layer1_outputs(1702));
    layer2_outputs(253) <= (layer1_outputs(1085)) xor (layer1_outputs(917));
    layer2_outputs(254) <= (layer1_outputs(1254)) or (layer1_outputs(2508));
    layer2_outputs(255) <= (layer1_outputs(1002)) or (layer1_outputs(1642));
    layer2_outputs(256) <= not(layer1_outputs(1069));
    layer2_outputs(257) <= (layer1_outputs(1593)) and (layer1_outputs(2278));
    layer2_outputs(258) <= not(layer1_outputs(366));
    layer2_outputs(259) <= (layer1_outputs(638)) or (layer1_outputs(1028));
    layer2_outputs(260) <= layer1_outputs(1536);
    layer2_outputs(261) <= not((layer1_outputs(1305)) and (layer1_outputs(2407)));
    layer2_outputs(262) <= not(layer1_outputs(1216)) or (layer1_outputs(946));
    layer2_outputs(263) <= not((layer1_outputs(2168)) or (layer1_outputs(805)));
    layer2_outputs(264) <= (layer1_outputs(2050)) and not (layer1_outputs(947));
    layer2_outputs(265) <= layer1_outputs(2070);
    layer2_outputs(266) <= not(layer1_outputs(1490));
    layer2_outputs(267) <= layer1_outputs(2124);
    layer2_outputs(268) <= (layer1_outputs(70)) and not (layer1_outputs(1817));
    layer2_outputs(269) <= layer1_outputs(1088);
    layer2_outputs(270) <= not(layer1_outputs(2398));
    layer2_outputs(271) <= not(layer1_outputs(1416));
    layer2_outputs(272) <= layer1_outputs(574);
    layer2_outputs(273) <= (layer1_outputs(626)) xor (layer1_outputs(1050));
    layer2_outputs(274) <= (layer1_outputs(2467)) and not (layer1_outputs(2160));
    layer2_outputs(275) <= not(layer1_outputs(196)) or (layer1_outputs(1683));
    layer2_outputs(276) <= not(layer1_outputs(1814)) or (layer1_outputs(1435));
    layer2_outputs(277) <= (layer1_outputs(302)) and not (layer1_outputs(720));
    layer2_outputs(278) <= layer1_outputs(2157);
    layer2_outputs(279) <= (layer1_outputs(2477)) and not (layer1_outputs(1592));
    layer2_outputs(280) <= not((layer1_outputs(884)) and (layer1_outputs(297)));
    layer2_outputs(281) <= (layer1_outputs(2027)) and not (layer1_outputs(511));
    layer2_outputs(282) <= not(layer1_outputs(1492)) or (layer1_outputs(371));
    layer2_outputs(283) <= not(layer1_outputs(1522)) or (layer1_outputs(771));
    layer2_outputs(284) <= layer1_outputs(1208);
    layer2_outputs(285) <= (layer1_outputs(1061)) or (layer1_outputs(1666));
    layer2_outputs(286) <= layer1_outputs(1728);
    layer2_outputs(287) <= layer1_outputs(1590);
    layer2_outputs(288) <= not((layer1_outputs(46)) and (layer1_outputs(380)));
    layer2_outputs(289) <= (layer1_outputs(2519)) and not (layer1_outputs(1980));
    layer2_outputs(290) <= not(layer1_outputs(140));
    layer2_outputs(291) <= not((layer1_outputs(422)) and (layer1_outputs(187)));
    layer2_outputs(292) <= (layer1_outputs(2466)) and not (layer1_outputs(2128));
    layer2_outputs(293) <= layer1_outputs(1781);
    layer2_outputs(294) <= layer1_outputs(1236);
    layer2_outputs(295) <= '1';
    layer2_outputs(296) <= (layer1_outputs(1591)) and not (layer1_outputs(113));
    layer2_outputs(297) <= not((layer1_outputs(2354)) or (layer1_outputs(2429)));
    layer2_outputs(298) <= layer1_outputs(2346);
    layer2_outputs(299) <= not((layer1_outputs(2449)) or (layer1_outputs(2271)));
    layer2_outputs(300) <= layer1_outputs(1239);
    layer2_outputs(301) <= not((layer1_outputs(347)) or (layer1_outputs(529)));
    layer2_outputs(302) <= not(layer1_outputs(1877));
    layer2_outputs(303) <= layer1_outputs(1379);
    layer2_outputs(304) <= not(layer1_outputs(217)) or (layer1_outputs(2192));
    layer2_outputs(305) <= (layer1_outputs(1000)) and not (layer1_outputs(2481));
    layer2_outputs(306) <= (layer1_outputs(2445)) and not (layer1_outputs(2533));
    layer2_outputs(307) <= not(layer1_outputs(47)) or (layer1_outputs(250));
    layer2_outputs(308) <= not((layer1_outputs(1145)) or (layer1_outputs(1363)));
    layer2_outputs(309) <= not(layer1_outputs(1809)) or (layer1_outputs(401));
    layer2_outputs(310) <= '0';
    layer2_outputs(311) <= not(layer1_outputs(1671));
    layer2_outputs(312) <= not(layer1_outputs(755));
    layer2_outputs(313) <= (layer1_outputs(65)) and not (layer1_outputs(2387));
    layer2_outputs(314) <= (layer1_outputs(482)) and not (layer1_outputs(596));
    layer2_outputs(315) <= (layer1_outputs(2139)) and not (layer1_outputs(1271));
    layer2_outputs(316) <= not(layer1_outputs(145)) or (layer1_outputs(350));
    layer2_outputs(317) <= (layer1_outputs(2141)) or (layer1_outputs(1092));
    layer2_outputs(318) <= layer1_outputs(2484);
    layer2_outputs(319) <= not(layer1_outputs(1734));
    layer2_outputs(320) <= layer1_outputs(1755);
    layer2_outputs(321) <= not((layer1_outputs(309)) or (layer1_outputs(1536)));
    layer2_outputs(322) <= not(layer1_outputs(1288));
    layer2_outputs(323) <= (layer1_outputs(725)) and not (layer1_outputs(202));
    layer2_outputs(324) <= not(layer1_outputs(1875));
    layer2_outputs(325) <= (layer1_outputs(787)) or (layer1_outputs(1735));
    layer2_outputs(326) <= (layer1_outputs(1078)) or (layer1_outputs(885));
    layer2_outputs(327) <= not((layer1_outputs(204)) or (layer1_outputs(2439)));
    layer2_outputs(328) <= not(layer1_outputs(1177));
    layer2_outputs(329) <= not(layer1_outputs(1268));
    layer2_outputs(330) <= not(layer1_outputs(1214)) or (layer1_outputs(2057));
    layer2_outputs(331) <= (layer1_outputs(1275)) and (layer1_outputs(1745));
    layer2_outputs(332) <= not(layer1_outputs(940));
    layer2_outputs(333) <= not(layer1_outputs(1448));
    layer2_outputs(334) <= layer1_outputs(863);
    layer2_outputs(335) <= not(layer1_outputs(1902));
    layer2_outputs(336) <= not(layer1_outputs(2300)) or (layer1_outputs(649));
    layer2_outputs(337) <= layer1_outputs(338);
    layer2_outputs(338) <= not((layer1_outputs(667)) or (layer1_outputs(404)));
    layer2_outputs(339) <= (layer1_outputs(1130)) and not (layer1_outputs(1042));
    layer2_outputs(340) <= (layer1_outputs(1894)) and not (layer1_outputs(2443));
    layer2_outputs(341) <= (layer1_outputs(2119)) or (layer1_outputs(1627));
    layer2_outputs(342) <= layer1_outputs(2044);
    layer2_outputs(343) <= not(layer1_outputs(1881)) or (layer1_outputs(1516));
    layer2_outputs(344) <= (layer1_outputs(1988)) or (layer1_outputs(1986));
    layer2_outputs(345) <= layer1_outputs(7);
    layer2_outputs(346) <= not(layer1_outputs(1833));
    layer2_outputs(347) <= not(layer1_outputs(5)) or (layer1_outputs(2016));
    layer2_outputs(348) <= layer1_outputs(675);
    layer2_outputs(349) <= layer1_outputs(1131);
    layer2_outputs(350) <= (layer1_outputs(986)) and not (layer1_outputs(657));
    layer2_outputs(351) <= (layer1_outputs(205)) or (layer1_outputs(840));
    layer2_outputs(352) <= (layer1_outputs(1749)) xor (layer1_outputs(1043));
    layer2_outputs(353) <= not(layer1_outputs(2343));
    layer2_outputs(354) <= (layer1_outputs(1463)) or (layer1_outputs(1054));
    layer2_outputs(355) <= layer1_outputs(1005);
    layer2_outputs(356) <= not(layer1_outputs(2261));
    layer2_outputs(357) <= not(layer1_outputs(1242));
    layer2_outputs(358) <= not(layer1_outputs(1671));
    layer2_outputs(359) <= not((layer1_outputs(559)) and (layer1_outputs(445)));
    layer2_outputs(360) <= not((layer1_outputs(2521)) and (layer1_outputs(636)));
    layer2_outputs(361) <= (layer1_outputs(839)) and not (layer1_outputs(1866));
    layer2_outputs(362) <= not(layer1_outputs(322));
    layer2_outputs(363) <= (layer1_outputs(1454)) xor (layer1_outputs(872));
    layer2_outputs(364) <= layer1_outputs(2276);
    layer2_outputs(365) <= layer1_outputs(9);
    layer2_outputs(366) <= not((layer1_outputs(178)) xor (layer1_outputs(1856)));
    layer2_outputs(367) <= (layer1_outputs(491)) or (layer1_outputs(1154));
    layer2_outputs(368) <= layer1_outputs(2197);
    layer2_outputs(369) <= '1';
    layer2_outputs(370) <= not((layer1_outputs(2202)) and (layer1_outputs(1377)));
    layer2_outputs(371) <= not(layer1_outputs(1667)) or (layer1_outputs(2039));
    layer2_outputs(372) <= (layer1_outputs(2461)) and (layer1_outputs(1369));
    layer2_outputs(373) <= layer1_outputs(2087);
    layer2_outputs(374) <= layer1_outputs(1240);
    layer2_outputs(375) <= not(layer1_outputs(2073)) or (layer1_outputs(749));
    layer2_outputs(376) <= (layer1_outputs(2357)) and not (layer1_outputs(1278));
    layer2_outputs(377) <= not(layer1_outputs(1187));
    layer2_outputs(378) <= layer1_outputs(1804);
    layer2_outputs(379) <= not((layer1_outputs(642)) or (layer1_outputs(1668)));
    layer2_outputs(380) <= layer1_outputs(2061);
    layer2_outputs(381) <= (layer1_outputs(1661)) or (layer1_outputs(1674));
    layer2_outputs(382) <= not(layer1_outputs(173));
    layer2_outputs(383) <= not((layer1_outputs(1176)) and (layer1_outputs(1889)));
    layer2_outputs(384) <= layer1_outputs(1826);
    layer2_outputs(385) <= not(layer1_outputs(2340));
    layer2_outputs(386) <= (layer1_outputs(1457)) and (layer1_outputs(1557));
    layer2_outputs(387) <= layer1_outputs(2068);
    layer2_outputs(388) <= not(layer1_outputs(555));
    layer2_outputs(389) <= layer1_outputs(950);
    layer2_outputs(390) <= not(layer1_outputs(1310)) or (layer1_outputs(528));
    layer2_outputs(391) <= not(layer1_outputs(2312));
    layer2_outputs(392) <= layer1_outputs(118);
    layer2_outputs(393) <= not(layer1_outputs(1756));
    layer2_outputs(394) <= not((layer1_outputs(358)) and (layer1_outputs(1138)));
    layer2_outputs(395) <= not(layer1_outputs(819)) or (layer1_outputs(1960));
    layer2_outputs(396) <= layer1_outputs(2152);
    layer2_outputs(397) <= layer1_outputs(922);
    layer2_outputs(398) <= not(layer1_outputs(21)) or (layer1_outputs(271));
    layer2_outputs(399) <= layer1_outputs(972);
    layer2_outputs(400) <= (layer1_outputs(2303)) xor (layer1_outputs(674));
    layer2_outputs(401) <= not(layer1_outputs(1256));
    layer2_outputs(402) <= not(layer1_outputs(1994)) or (layer1_outputs(194));
    layer2_outputs(403) <= not((layer1_outputs(1643)) and (layer1_outputs(2448)));
    layer2_outputs(404) <= layer1_outputs(1019);
    layer2_outputs(405) <= not((layer1_outputs(2421)) xor (layer1_outputs(1146)));
    layer2_outputs(406) <= layer1_outputs(311);
    layer2_outputs(407) <= layer1_outputs(1047);
    layer2_outputs(408) <= (layer1_outputs(1076)) xor (layer1_outputs(100));
    layer2_outputs(409) <= layer1_outputs(718);
    layer2_outputs(410) <= layer1_outputs(1268);
    layer2_outputs(411) <= not((layer1_outputs(2525)) or (layer1_outputs(2377)));
    layer2_outputs(412) <= not((layer1_outputs(1595)) and (layer1_outputs(1008)));
    layer2_outputs(413) <= layer1_outputs(1496);
    layer2_outputs(414) <= layer1_outputs(2066);
    layer2_outputs(415) <= layer1_outputs(1746);
    layer2_outputs(416) <= not(layer1_outputs(361));
    layer2_outputs(417) <= (layer1_outputs(1575)) and not (layer1_outputs(2550));
    layer2_outputs(418) <= layer1_outputs(1068);
    layer2_outputs(419) <= (layer1_outputs(1029)) xor (layer1_outputs(689));
    layer2_outputs(420) <= (layer1_outputs(1765)) and (layer1_outputs(169));
    layer2_outputs(421) <= not((layer1_outputs(2488)) and (layer1_outputs(646)));
    layer2_outputs(422) <= layer1_outputs(1808);
    layer2_outputs(423) <= not(layer1_outputs(2281)) or (layer1_outputs(393));
    layer2_outputs(424) <= (layer1_outputs(80)) and not (layer1_outputs(2433));
    layer2_outputs(425) <= (layer1_outputs(2248)) xor (layer1_outputs(392));
    layer2_outputs(426) <= not(layer1_outputs(1269));
    layer2_outputs(427) <= (layer1_outputs(2324)) and (layer1_outputs(1639));
    layer2_outputs(428) <= '1';
    layer2_outputs(429) <= (layer1_outputs(363)) or (layer1_outputs(1872));
    layer2_outputs(430) <= layer1_outputs(1686);
    layer2_outputs(431) <= '1';
    layer2_outputs(432) <= not(layer1_outputs(2227));
    layer2_outputs(433) <= not(layer1_outputs(426)) or (layer1_outputs(1918));
    layer2_outputs(434) <= layer1_outputs(1328);
    layer2_outputs(435) <= not(layer1_outputs(680));
    layer2_outputs(436) <= layer1_outputs(1477);
    layer2_outputs(437) <= layer1_outputs(1301);
    layer2_outputs(438) <= not((layer1_outputs(1921)) or (layer1_outputs(2175)));
    layer2_outputs(439) <= (layer1_outputs(1958)) and not (layer1_outputs(706));
    layer2_outputs(440) <= (layer1_outputs(806)) and not (layer1_outputs(1009));
    layer2_outputs(441) <= not(layer1_outputs(2169)) or (layer1_outputs(982));
    layer2_outputs(442) <= layer1_outputs(2137);
    layer2_outputs(443) <= not(layer1_outputs(464));
    layer2_outputs(444) <= not(layer1_outputs(1599)) or (layer1_outputs(1893));
    layer2_outputs(445) <= not(layer1_outputs(2331));
    layer2_outputs(446) <= not(layer1_outputs(13)) or (layer1_outputs(687));
    layer2_outputs(447) <= not((layer1_outputs(1539)) xor (layer1_outputs(1811)));
    layer2_outputs(448) <= layer1_outputs(782);
    layer2_outputs(449) <= not(layer1_outputs(156));
    layer2_outputs(450) <= layer1_outputs(31);
    layer2_outputs(451) <= (layer1_outputs(57)) and not (layer1_outputs(554));
    layer2_outputs(452) <= (layer1_outputs(1860)) xor (layer1_outputs(2021));
    layer2_outputs(453) <= not((layer1_outputs(24)) and (layer1_outputs(1332)));
    layer2_outputs(454) <= not(layer1_outputs(2474)) or (layer1_outputs(942));
    layer2_outputs(455) <= not(layer1_outputs(1212));
    layer2_outputs(456) <= (layer1_outputs(594)) or (layer1_outputs(1066));
    layer2_outputs(457) <= not(layer1_outputs(816));
    layer2_outputs(458) <= (layer1_outputs(356)) or (layer1_outputs(634));
    layer2_outputs(459) <= layer1_outputs(212);
    layer2_outputs(460) <= layer1_outputs(1360);
    layer2_outputs(461) <= not(layer1_outputs(1815)) or (layer1_outputs(1800));
    layer2_outputs(462) <= not(layer1_outputs(1273));
    layer2_outputs(463) <= layer1_outputs(391);
    layer2_outputs(464) <= not(layer1_outputs(1460)) or (layer1_outputs(2339));
    layer2_outputs(465) <= not(layer1_outputs(443));
    layer2_outputs(466) <= not((layer1_outputs(1716)) or (layer1_outputs(667)));
    layer2_outputs(467) <= (layer1_outputs(2091)) and not (layer1_outputs(1118));
    layer2_outputs(468) <= not((layer1_outputs(1893)) or (layer1_outputs(1145)));
    layer2_outputs(469) <= layer1_outputs(2184);
    layer2_outputs(470) <= (layer1_outputs(589)) and (layer1_outputs(77));
    layer2_outputs(471) <= layer1_outputs(1292);
    layer2_outputs(472) <= not(layer1_outputs(643));
    layer2_outputs(473) <= not(layer1_outputs(577));
    layer2_outputs(474) <= layer1_outputs(539);
    layer2_outputs(475) <= layer1_outputs(1370);
    layer2_outputs(476) <= (layer1_outputs(1502)) and not (layer1_outputs(1651));
    layer2_outputs(477) <= (layer1_outputs(1718)) and (layer1_outputs(655));
    layer2_outputs(478) <= not(layer1_outputs(923)) or (layer1_outputs(1839));
    layer2_outputs(479) <= not((layer1_outputs(430)) and (layer1_outputs(2475)));
    layer2_outputs(480) <= not(layer1_outputs(1450)) or (layer1_outputs(1327));
    layer2_outputs(481) <= not(layer1_outputs(1549)) or (layer1_outputs(894));
    layer2_outputs(482) <= not(layer1_outputs(132));
    layer2_outputs(483) <= not(layer1_outputs(1223));
    layer2_outputs(484) <= layer1_outputs(18);
    layer2_outputs(485) <= layer1_outputs(144);
    layer2_outputs(486) <= layer1_outputs(2367);
    layer2_outputs(487) <= not(layer1_outputs(1555)) or (layer1_outputs(312));
    layer2_outputs(488) <= not((layer1_outputs(652)) or (layer1_outputs(2349)));
    layer2_outputs(489) <= layer1_outputs(613);
    layer2_outputs(490) <= not(layer1_outputs(1964)) or (layer1_outputs(1543));
    layer2_outputs(491) <= layer1_outputs(2358);
    layer2_outputs(492) <= not((layer1_outputs(948)) xor (layer1_outputs(1291)));
    layer2_outputs(493) <= layer1_outputs(1902);
    layer2_outputs(494) <= layer1_outputs(1656);
    layer2_outputs(495) <= not(layer1_outputs(1527)) or (layer1_outputs(167));
    layer2_outputs(496) <= not(layer1_outputs(811)) or (layer1_outputs(758));
    layer2_outputs(497) <= not(layer1_outputs(1038));
    layer2_outputs(498) <= not(layer1_outputs(308));
    layer2_outputs(499) <= not(layer1_outputs(432)) or (layer1_outputs(250));
    layer2_outputs(500) <= not(layer1_outputs(414)) or (layer1_outputs(230));
    layer2_outputs(501) <= '0';
    layer2_outputs(502) <= layer1_outputs(768);
    layer2_outputs(503) <= (layer1_outputs(1549)) and (layer1_outputs(1912));
    layer2_outputs(504) <= (layer1_outputs(1202)) and not (layer1_outputs(1850));
    layer2_outputs(505) <= not(layer1_outputs(1538));
    layer2_outputs(506) <= not(layer1_outputs(2432));
    layer2_outputs(507) <= not((layer1_outputs(2002)) or (layer1_outputs(2522)));
    layer2_outputs(508) <= layer1_outputs(313);
    layer2_outputs(509) <= not(layer1_outputs(231));
    layer2_outputs(510) <= layer1_outputs(1681);
    layer2_outputs(511) <= (layer1_outputs(1629)) and not (layer1_outputs(2083));
    layer2_outputs(512) <= (layer1_outputs(2208)) and not (layer1_outputs(1030));
    layer2_outputs(513) <= not(layer1_outputs(2381));
    layer2_outputs(514) <= not(layer1_outputs(777));
    layer2_outputs(515) <= layer1_outputs(55);
    layer2_outputs(516) <= (layer1_outputs(1747)) and not (layer1_outputs(1234));
    layer2_outputs(517) <= not(layer1_outputs(1129));
    layer2_outputs(518) <= layer1_outputs(2335);
    layer2_outputs(519) <= layer1_outputs(451);
    layer2_outputs(520) <= (layer1_outputs(23)) or (layer1_outputs(687));
    layer2_outputs(521) <= (layer1_outputs(83)) and not (layer1_outputs(212));
    layer2_outputs(522) <= not(layer1_outputs(76));
    layer2_outputs(523) <= not(layer1_outputs(2318));
    layer2_outputs(524) <= not(layer1_outputs(1178)) or (layer1_outputs(2229));
    layer2_outputs(525) <= layer1_outputs(511);
    layer2_outputs(526) <= not(layer1_outputs(2140)) or (layer1_outputs(2212));
    layer2_outputs(527) <= not(layer1_outputs(314));
    layer2_outputs(528) <= not(layer1_outputs(2356));
    layer2_outputs(529) <= not(layer1_outputs(508));
    layer2_outputs(530) <= layer1_outputs(623);
    layer2_outputs(531) <= (layer1_outputs(130)) and (layer1_outputs(467));
    layer2_outputs(532) <= not((layer1_outputs(2234)) and (layer1_outputs(1333)));
    layer2_outputs(533) <= layer1_outputs(472);
    layer2_outputs(534) <= not((layer1_outputs(2317)) and (layer1_outputs(2025)));
    layer2_outputs(535) <= not(layer1_outputs(24));
    layer2_outputs(536) <= not(layer1_outputs(456));
    layer2_outputs(537) <= not(layer1_outputs(2346));
    layer2_outputs(538) <= not((layer1_outputs(1264)) and (layer1_outputs(1104)));
    layer2_outputs(539) <= not(layer1_outputs(1864));
    layer2_outputs(540) <= not(layer1_outputs(1583)) or (layer1_outputs(1193));
    layer2_outputs(541) <= not(layer1_outputs(2521));
    layer2_outputs(542) <= not(layer1_outputs(96)) or (layer1_outputs(1121));
    layer2_outputs(543) <= not((layer1_outputs(1210)) xor (layer1_outputs(1800)));
    layer2_outputs(544) <= layer1_outputs(899);
    layer2_outputs(545) <= not((layer1_outputs(2428)) and (layer1_outputs(390)));
    layer2_outputs(546) <= not((layer1_outputs(2370)) or (layer1_outputs(1784)));
    layer2_outputs(547) <= not(layer1_outputs(1620));
    layer2_outputs(548) <= (layer1_outputs(1307)) or (layer1_outputs(1698));
    layer2_outputs(549) <= not((layer1_outputs(625)) and (layer1_outputs(1635)));
    layer2_outputs(550) <= not((layer1_outputs(1179)) and (layer1_outputs(1216)));
    layer2_outputs(551) <= layer1_outputs(2299);
    layer2_outputs(552) <= not((layer1_outputs(1927)) and (layer1_outputs(692)));
    layer2_outputs(553) <= (layer1_outputs(599)) and (layer1_outputs(858));
    layer2_outputs(554) <= '0';
    layer2_outputs(555) <= layer1_outputs(2029);
    layer2_outputs(556) <= layer1_outputs(1768);
    layer2_outputs(557) <= (layer1_outputs(126)) xor (layer1_outputs(580));
    layer2_outputs(558) <= (layer1_outputs(883)) and (layer1_outputs(180));
    layer2_outputs(559) <= not(layer1_outputs(1626));
    layer2_outputs(560) <= not((layer1_outputs(1210)) xor (layer1_outputs(2247)));
    layer2_outputs(561) <= not(layer1_outputs(1413));
    layer2_outputs(562) <= (layer1_outputs(100)) or (layer1_outputs(1263));
    layer2_outputs(563) <= not(layer1_outputs(2255)) or (layer1_outputs(1745));
    layer2_outputs(564) <= not(layer1_outputs(2078)) or (layer1_outputs(307));
    layer2_outputs(565) <= not(layer1_outputs(989));
    layer2_outputs(566) <= (layer1_outputs(1585)) and (layer1_outputs(1469));
    layer2_outputs(567) <= (layer1_outputs(105)) and not (layer1_outputs(580));
    layer2_outputs(568) <= not(layer1_outputs(1964));
    layer2_outputs(569) <= not(layer1_outputs(1287));
    layer2_outputs(570) <= not(layer1_outputs(1310)) or (layer1_outputs(1220));
    layer2_outputs(571) <= layer1_outputs(741);
    layer2_outputs(572) <= layer1_outputs(122);
    layer2_outputs(573) <= (layer1_outputs(1306)) or (layer1_outputs(1371));
    layer2_outputs(574) <= not(layer1_outputs(1260)) or (layer1_outputs(203));
    layer2_outputs(575) <= layer1_outputs(1625);
    layer2_outputs(576) <= (layer1_outputs(1451)) and (layer1_outputs(236));
    layer2_outputs(577) <= not(layer1_outputs(2517));
    layer2_outputs(578) <= not((layer1_outputs(612)) and (layer1_outputs(1822)));
    layer2_outputs(579) <= layer1_outputs(2510);
    layer2_outputs(580) <= not((layer1_outputs(2298)) and (layer1_outputs(1697)));
    layer2_outputs(581) <= (layer1_outputs(1126)) xor (layer1_outputs(1812));
    layer2_outputs(582) <= not(layer1_outputs(1292)) or (layer1_outputs(349));
    layer2_outputs(583) <= not((layer1_outputs(895)) and (layer1_outputs(1935)));
    layer2_outputs(584) <= not(layer1_outputs(147)) or (layer1_outputs(807));
    layer2_outputs(585) <= layer1_outputs(953);
    layer2_outputs(586) <= not((layer1_outputs(1949)) xor (layer1_outputs(2179)));
    layer2_outputs(587) <= not((layer1_outputs(2529)) or (layer1_outputs(1337)));
    layer2_outputs(588) <= (layer1_outputs(617)) and (layer1_outputs(1014));
    layer2_outputs(589) <= layer1_outputs(1949);
    layer2_outputs(590) <= (layer1_outputs(215)) xor (layer1_outputs(868));
    layer2_outputs(591) <= layer1_outputs(2184);
    layer2_outputs(592) <= not(layer1_outputs(1382)) or (layer1_outputs(1739));
    layer2_outputs(593) <= not((layer1_outputs(505)) or (layer1_outputs(2380)));
    layer2_outputs(594) <= not((layer1_outputs(195)) or (layer1_outputs(2446)));
    layer2_outputs(595) <= layer1_outputs(947);
    layer2_outputs(596) <= layer1_outputs(1319);
    layer2_outputs(597) <= not(layer1_outputs(90)) or (layer1_outputs(1586));
    layer2_outputs(598) <= layer1_outputs(59);
    layer2_outputs(599) <= layer1_outputs(351);
    layer2_outputs(600) <= not(layer1_outputs(633));
    layer2_outputs(601) <= (layer1_outputs(2520)) or (layer1_outputs(435));
    layer2_outputs(602) <= not(layer1_outputs(2518));
    layer2_outputs(603) <= not(layer1_outputs(1271));
    layer2_outputs(604) <= not(layer1_outputs(745));
    layer2_outputs(605) <= (layer1_outputs(1403)) xor (layer1_outputs(359));
    layer2_outputs(606) <= not(layer1_outputs(1103));
    layer2_outputs(607) <= (layer1_outputs(2223)) and not (layer1_outputs(2260));
    layer2_outputs(608) <= (layer1_outputs(1682)) and not (layer1_outputs(1955));
    layer2_outputs(609) <= layer1_outputs(1986);
    layer2_outputs(610) <= not(layer1_outputs(954));
    layer2_outputs(611) <= layer1_outputs(427);
    layer2_outputs(612) <= not((layer1_outputs(2160)) or (layer1_outputs(1661)));
    layer2_outputs(613) <= (layer1_outputs(527)) and (layer1_outputs(2558));
    layer2_outputs(614) <= (layer1_outputs(1122)) and not (layer1_outputs(1024));
    layer2_outputs(615) <= not(layer1_outputs(1424)) or (layer1_outputs(1344));
    layer2_outputs(616) <= (layer1_outputs(1930)) and (layer1_outputs(1325));
    layer2_outputs(617) <= (layer1_outputs(1491)) or (layer1_outputs(1909));
    layer2_outputs(618) <= not((layer1_outputs(319)) and (layer1_outputs(779)));
    layer2_outputs(619) <= (layer1_outputs(579)) and not (layer1_outputs(2244));
    layer2_outputs(620) <= not(layer1_outputs(1315));
    layer2_outputs(621) <= not(layer1_outputs(1630)) or (layer1_outputs(388));
    layer2_outputs(622) <= not((layer1_outputs(633)) and (layer1_outputs(2559)));
    layer2_outputs(623) <= '1';
    layer2_outputs(624) <= layer1_outputs(2062);
    layer2_outputs(625) <= (layer1_outputs(2076)) and not (layer1_outputs(2286));
    layer2_outputs(626) <= layer1_outputs(99);
    layer2_outputs(627) <= layer1_outputs(1244);
    layer2_outputs(628) <= layer1_outputs(2530);
    layer2_outputs(629) <= layer1_outputs(8);
    layer2_outputs(630) <= not((layer1_outputs(1207)) or (layer1_outputs(2007)));
    layer2_outputs(631) <= (layer1_outputs(284)) or (layer1_outputs(843));
    layer2_outputs(632) <= not((layer1_outputs(1601)) or (layer1_outputs(617)));
    layer2_outputs(633) <= not(layer1_outputs(2151));
    layer2_outputs(634) <= not((layer1_outputs(995)) or (layer1_outputs(2434)));
    layer2_outputs(635) <= (layer1_outputs(622)) and not (layer1_outputs(2221));
    layer2_outputs(636) <= not(layer1_outputs(379));
    layer2_outputs(637) <= layer1_outputs(2554);
    layer2_outputs(638) <= not((layer1_outputs(740)) and (layer1_outputs(58)));
    layer2_outputs(639) <= (layer1_outputs(1316)) and not (layer1_outputs(500));
    layer2_outputs(640) <= (layer1_outputs(834)) or (layer1_outputs(1761));
    layer2_outputs(641) <= not(layer1_outputs(640));
    layer2_outputs(642) <= layer1_outputs(2390);
    layer2_outputs(643) <= (layer1_outputs(2037)) and (layer1_outputs(806));
    layer2_outputs(644) <= not((layer1_outputs(1813)) and (layer1_outputs(2373)));
    layer2_outputs(645) <= layer1_outputs(2045);
    layer2_outputs(646) <= not(layer1_outputs(1436));
    layer2_outputs(647) <= not(layer1_outputs(1528));
    layer2_outputs(648) <= (layer1_outputs(1161)) and not (layer1_outputs(2132));
    layer2_outputs(649) <= not(layer1_outputs(2175));
    layer2_outputs(650) <= (layer1_outputs(170)) and not (layer1_outputs(164));
    layer2_outputs(651) <= not((layer1_outputs(277)) and (layer1_outputs(727)));
    layer2_outputs(652) <= '0';
    layer2_outputs(653) <= layer1_outputs(2523);
    layer2_outputs(654) <= layer1_outputs(1442);
    layer2_outputs(655) <= layer1_outputs(1685);
    layer2_outputs(656) <= (layer1_outputs(396)) and (layer1_outputs(1751));
    layer2_outputs(657) <= not(layer1_outputs(697));
    layer2_outputs(658) <= layer1_outputs(367);
    layer2_outputs(659) <= not(layer1_outputs(1423));
    layer2_outputs(660) <= not(layer1_outputs(2254));
    layer2_outputs(661) <= layer1_outputs(2554);
    layer2_outputs(662) <= not(layer1_outputs(1511)) or (layer1_outputs(10));
    layer2_outputs(663) <= layer1_outputs(1128);
    layer2_outputs(664) <= layer1_outputs(425);
    layer2_outputs(665) <= not(layer1_outputs(2312));
    layer2_outputs(666) <= (layer1_outputs(413)) and not (layer1_outputs(74));
    layer2_outputs(667) <= not((layer1_outputs(1736)) or (layer1_outputs(473)));
    layer2_outputs(668) <= not(layer1_outputs(558)) or (layer1_outputs(814));
    layer2_outputs(669) <= (layer1_outputs(2101)) and not (layer1_outputs(1524));
    layer2_outputs(670) <= not((layer1_outputs(101)) xor (layer1_outputs(2484)));
    layer2_outputs(671) <= layer1_outputs(873);
    layer2_outputs(672) <= not((layer1_outputs(1385)) or (layer1_outputs(1119)));
    layer2_outputs(673) <= (layer1_outputs(154)) or (layer1_outputs(1034));
    layer2_outputs(674) <= not(layer1_outputs(2495));
    layer2_outputs(675) <= not((layer1_outputs(83)) or (layer1_outputs(743)));
    layer2_outputs(676) <= not(layer1_outputs(1191)) or (layer1_outputs(514));
    layer2_outputs(677) <= not(layer1_outputs(453));
    layer2_outputs(678) <= not((layer1_outputs(1188)) or (layer1_outputs(964)));
    layer2_outputs(679) <= not(layer1_outputs(402)) or (layer1_outputs(820));
    layer2_outputs(680) <= not(layer1_outputs(361));
    layer2_outputs(681) <= (layer1_outputs(484)) or (layer1_outputs(382));
    layer2_outputs(682) <= not((layer1_outputs(1968)) or (layer1_outputs(1600)));
    layer2_outputs(683) <= (layer1_outputs(1250)) and (layer1_outputs(2320));
    layer2_outputs(684) <= not(layer1_outputs(1539)) or (layer1_outputs(1844));
    layer2_outputs(685) <= '1';
    layer2_outputs(686) <= (layer1_outputs(1293)) and not (layer1_outputs(1291));
    layer2_outputs(687) <= not((layer1_outputs(2280)) and (layer1_outputs(902)));
    layer2_outputs(688) <= not(layer1_outputs(463)) or (layer1_outputs(1478));
    layer2_outputs(689) <= (layer1_outputs(140)) and not (layer1_outputs(1615));
    layer2_outputs(690) <= not(layer1_outputs(127));
    layer2_outputs(691) <= layer1_outputs(1841);
    layer2_outputs(692) <= not(layer1_outputs(725));
    layer2_outputs(693) <= not(layer1_outputs(2383));
    layer2_outputs(694) <= not(layer1_outputs(2053));
    layer2_outputs(695) <= not(layer1_outputs(2556));
    layer2_outputs(696) <= (layer1_outputs(2421)) and (layer1_outputs(264));
    layer2_outputs(697) <= (layer1_outputs(1308)) and not (layer1_outputs(1155));
    layer2_outputs(698) <= not(layer1_outputs(2458)) or (layer1_outputs(2164));
    layer2_outputs(699) <= layer1_outputs(2483);
    layer2_outputs(700) <= not((layer1_outputs(1321)) and (layer1_outputs(2502)));
    layer2_outputs(701) <= (layer1_outputs(829)) and (layer1_outputs(1855));
    layer2_outputs(702) <= not((layer1_outputs(1783)) xor (layer1_outputs(31)));
    layer2_outputs(703) <= not((layer1_outputs(541)) or (layer1_outputs(1724)));
    layer2_outputs(704) <= layer1_outputs(2535);
    layer2_outputs(705) <= not(layer1_outputs(1217));
    layer2_outputs(706) <= (layer1_outputs(105)) and (layer1_outputs(2461));
    layer2_outputs(707) <= not(layer1_outputs(2059));
    layer2_outputs(708) <= layer1_outputs(1068);
    layer2_outputs(709) <= not(layer1_outputs(1970));
    layer2_outputs(710) <= (layer1_outputs(645)) and not (layer1_outputs(464));
    layer2_outputs(711) <= layer1_outputs(772);
    layer2_outputs(712) <= layer1_outputs(1686);
    layer2_outputs(713) <= (layer1_outputs(2174)) or (layer1_outputs(1035));
    layer2_outputs(714) <= (layer1_outputs(2372)) and not (layer1_outputs(1227));
    layer2_outputs(715) <= (layer1_outputs(1444)) or (layer1_outputs(1859));
    layer2_outputs(716) <= (layer1_outputs(103)) and not (layer1_outputs(2371));
    layer2_outputs(717) <= not((layer1_outputs(82)) or (layer1_outputs(1678)));
    layer2_outputs(718) <= (layer1_outputs(1152)) and (layer1_outputs(747));
    layer2_outputs(719) <= not(layer1_outputs(1418)) or (layer1_outputs(352));
    layer2_outputs(720) <= (layer1_outputs(1733)) or (layer1_outputs(1203));
    layer2_outputs(721) <= not(layer1_outputs(546));
    layer2_outputs(722) <= not(layer1_outputs(1876));
    layer2_outputs(723) <= (layer1_outputs(451)) and not (layer1_outputs(127));
    layer2_outputs(724) <= not(layer1_outputs(421));
    layer2_outputs(725) <= layer1_outputs(20);
    layer2_outputs(726) <= layer1_outputs(963);
    layer2_outputs(727) <= (layer1_outputs(132)) and not (layer1_outputs(454));
    layer2_outputs(728) <= not(layer1_outputs(210));
    layer2_outputs(729) <= layer1_outputs(603);
    layer2_outputs(730) <= not(layer1_outputs(1722));
    layer2_outputs(731) <= (layer1_outputs(971)) or (layer1_outputs(2493));
    layer2_outputs(732) <= '1';
    layer2_outputs(733) <= layer1_outputs(1908);
    layer2_outputs(734) <= not((layer1_outputs(1554)) or (layer1_outputs(701)));
    layer2_outputs(735) <= not(layer1_outputs(2460)) or (layer1_outputs(1111));
    layer2_outputs(736) <= (layer1_outputs(1362)) and (layer1_outputs(1558));
    layer2_outputs(737) <= not((layer1_outputs(1514)) and (layer1_outputs(1631)));
    layer2_outputs(738) <= '0';
    layer2_outputs(739) <= not(layer1_outputs(1962));
    layer2_outputs(740) <= not(layer1_outputs(649));
    layer2_outputs(741) <= not(layer1_outputs(1340)) or (layer1_outputs(181));
    layer2_outputs(742) <= layer1_outputs(2551);
    layer2_outputs(743) <= layer1_outputs(340);
    layer2_outputs(744) <= not(layer1_outputs(2526)) or (layer1_outputs(1307));
    layer2_outputs(745) <= layer1_outputs(437);
    layer2_outputs(746) <= not(layer1_outputs(1265)) or (layer1_outputs(2101));
    layer2_outputs(747) <= layer1_outputs(843);
    layer2_outputs(748) <= (layer1_outputs(1880)) and not (layer1_outputs(733));
    layer2_outputs(749) <= not((layer1_outputs(1164)) xor (layer1_outputs(601)));
    layer2_outputs(750) <= not(layer1_outputs(317));
    layer2_outputs(751) <= layer1_outputs(1465);
    layer2_outputs(752) <= not((layer1_outputs(61)) and (layer1_outputs(1820)));
    layer2_outputs(753) <= (layer1_outputs(467)) and not (layer1_outputs(2474));
    layer2_outputs(754) <= not((layer1_outputs(2095)) or (layer1_outputs(609)));
    layer2_outputs(755) <= (layer1_outputs(2393)) and not (layer1_outputs(1916));
    layer2_outputs(756) <= not(layer1_outputs(482));
    layer2_outputs(757) <= (layer1_outputs(1922)) and (layer1_outputs(2220));
    layer2_outputs(758) <= layer1_outputs(1488);
    layer2_outputs(759) <= (layer1_outputs(2430)) and not (layer1_outputs(765));
    layer2_outputs(760) <= (layer1_outputs(1139)) and not (layer1_outputs(652));
    layer2_outputs(761) <= layer1_outputs(1179);
    layer2_outputs(762) <= layer1_outputs(191);
    layer2_outputs(763) <= not(layer1_outputs(1579)) or (layer1_outputs(550));
    layer2_outputs(764) <= (layer1_outputs(2228)) and not (layer1_outputs(2314));
    layer2_outputs(765) <= not((layer1_outputs(416)) and (layer1_outputs(362)));
    layer2_outputs(766) <= not((layer1_outputs(68)) and (layer1_outputs(2098)));
    layer2_outputs(767) <= (layer1_outputs(576)) and not (layer1_outputs(1521));
    layer2_outputs(768) <= layer1_outputs(1731);
    layer2_outputs(769) <= layer1_outputs(1476);
    layer2_outputs(770) <= not(layer1_outputs(2336));
    layer2_outputs(771) <= not(layer1_outputs(29));
    layer2_outputs(772) <= not(layer1_outputs(593));
    layer2_outputs(773) <= (layer1_outputs(1901)) or (layer1_outputs(1874));
    layer2_outputs(774) <= not(layer1_outputs(354)) or (layer1_outputs(1001));
    layer2_outputs(775) <= not(layer1_outputs(2499));
    layer2_outputs(776) <= not(layer1_outputs(1006));
    layer2_outputs(777) <= not(layer1_outputs(1398)) or (layer1_outputs(2546));
    layer2_outputs(778) <= not(layer1_outputs(220));
    layer2_outputs(779) <= not(layer1_outputs(2080)) or (layer1_outputs(1423));
    layer2_outputs(780) <= not((layer1_outputs(150)) or (layer1_outputs(2031)));
    layer2_outputs(781) <= (layer1_outputs(2390)) and not (layer1_outputs(1663));
    layer2_outputs(782) <= not((layer1_outputs(562)) and (layer1_outputs(176)));
    layer2_outputs(783) <= not(layer1_outputs(1414));
    layer2_outputs(784) <= (layer1_outputs(2099)) or (layer1_outputs(2462));
    layer2_outputs(785) <= not(layer1_outputs(1880));
    layer2_outputs(786) <= layer1_outputs(1851);
    layer2_outputs(787) <= layer1_outputs(553);
    layer2_outputs(788) <= not(layer1_outputs(1974)) or (layer1_outputs(1859));
    layer2_outputs(789) <= not((layer1_outputs(1794)) or (layer1_outputs(252)));
    layer2_outputs(790) <= not(layer1_outputs(373)) or (layer1_outputs(1698));
    layer2_outputs(791) <= layer1_outputs(264);
    layer2_outputs(792) <= not(layer1_outputs(925));
    layer2_outputs(793) <= layer1_outputs(1497);
    layer2_outputs(794) <= not(layer1_outputs(2118));
    layer2_outputs(795) <= layer1_outputs(112);
    layer2_outputs(796) <= not((layer1_outputs(1883)) xor (layer1_outputs(1983)));
    layer2_outputs(797) <= layer1_outputs(1441);
    layer2_outputs(798) <= not(layer1_outputs(510)) or (layer1_outputs(32));
    layer2_outputs(799) <= layer1_outputs(1105);
    layer2_outputs(800) <= layer1_outputs(2384);
    layer2_outputs(801) <= not(layer1_outputs(1765)) or (layer1_outputs(2440));
    layer2_outputs(802) <= not(layer1_outputs(411)) or (layer1_outputs(1452));
    layer2_outputs(803) <= not(layer1_outputs(1910));
    layer2_outputs(804) <= not(layer1_outputs(2181));
    layer2_outputs(805) <= not(layer1_outputs(1967));
    layer2_outputs(806) <= (layer1_outputs(2269)) and not (layer1_outputs(808));
    layer2_outputs(807) <= (layer1_outputs(627)) and not (layer1_outputs(1100));
    layer2_outputs(808) <= not(layer1_outputs(1899));
    layer2_outputs(809) <= layer1_outputs(880);
    layer2_outputs(810) <= layer1_outputs(709);
    layer2_outputs(811) <= not(layer1_outputs(662));
    layer2_outputs(812) <= layer1_outputs(2549);
    layer2_outputs(813) <= not((layer1_outputs(273)) and (layer1_outputs(2011)));
    layer2_outputs(814) <= not((layer1_outputs(1973)) and (layer1_outputs(1381)));
    layer2_outputs(815) <= not(layer1_outputs(2524));
    layer2_outputs(816) <= (layer1_outputs(224)) and not (layer1_outputs(219));
    layer2_outputs(817) <= not(layer1_outputs(2095));
    layer2_outputs(818) <= not(layer1_outputs(2284)) or (layer1_outputs(1525));
    layer2_outputs(819) <= not((layer1_outputs(2286)) and (layer1_outputs(158)));
    layer2_outputs(820) <= not((layer1_outputs(84)) xor (layer1_outputs(671)));
    layer2_outputs(821) <= (layer1_outputs(323)) and (layer1_outputs(433));
    layer2_outputs(822) <= not((layer1_outputs(1803)) or (layer1_outputs(2313)));
    layer2_outputs(823) <= (layer1_outputs(1059)) and not (layer1_outputs(557));
    layer2_outputs(824) <= not(layer1_outputs(691));
    layer2_outputs(825) <= not(layer1_outputs(2283));
    layer2_outputs(826) <= not(layer1_outputs(1193)) or (layer1_outputs(1102));
    layer2_outputs(827) <= layer1_outputs(900);
    layer2_outputs(828) <= not(layer1_outputs(1296)) or (layer1_outputs(909));
    layer2_outputs(829) <= not(layer1_outputs(1598)) or (layer1_outputs(1655));
    layer2_outputs(830) <= not(layer1_outputs(2017)) or (layer1_outputs(2265));
    layer2_outputs(831) <= (layer1_outputs(2145)) and not (layer1_outputs(2498));
    layer2_outputs(832) <= layer1_outputs(2146);
    layer2_outputs(833) <= (layer1_outputs(2339)) and not (layer1_outputs(2443));
    layer2_outputs(834) <= layer1_outputs(2209);
    layer2_outputs(835) <= not(layer1_outputs(2058));
    layer2_outputs(836) <= not(layer1_outputs(1127));
    layer2_outputs(837) <= (layer1_outputs(2436)) or (layer1_outputs(526));
    layer2_outputs(838) <= not(layer1_outputs(414)) or (layer1_outputs(1453));
    layer2_outputs(839) <= not(layer1_outputs(1295)) or (layer1_outputs(2270));
    layer2_outputs(840) <= not(layer1_outputs(541)) or (layer1_outputs(1481));
    layer2_outputs(841) <= not(layer1_outputs(232));
    layer2_outputs(842) <= layer1_outputs(1660);
    layer2_outputs(843) <= not(layer1_outputs(936)) or (layer1_outputs(243));
    layer2_outputs(844) <= not(layer1_outputs(2082));
    layer2_outputs(845) <= (layer1_outputs(1899)) or (layer1_outputs(224));
    layer2_outputs(846) <= (layer1_outputs(1535)) and not (layer1_outputs(1748));
    layer2_outputs(847) <= (layer1_outputs(2116)) or (layer1_outputs(2189));
    layer2_outputs(848) <= not(layer1_outputs(315)) or (layer1_outputs(1261));
    layer2_outputs(849) <= layer1_outputs(1867);
    layer2_outputs(850) <= layer1_outputs(1361);
    layer2_outputs(851) <= not(layer1_outputs(1426)) or (layer1_outputs(1460));
    layer2_outputs(852) <= (layer1_outputs(1054)) or (layer1_outputs(719));
    layer2_outputs(853) <= (layer1_outputs(2527)) or (layer1_outputs(1323));
    layer2_outputs(854) <= not((layer1_outputs(2170)) and (layer1_outputs(2200)));
    layer2_outputs(855) <= layer1_outputs(1951);
    layer2_outputs(856) <= not((layer1_outputs(144)) and (layer1_outputs(1551)));
    layer2_outputs(857) <= not(layer1_outputs(1864)) or (layer1_outputs(2130));
    layer2_outputs(858) <= not(layer1_outputs(910));
    layer2_outputs(859) <= not(layer1_outputs(1772));
    layer2_outputs(860) <= not((layer1_outputs(139)) and (layer1_outputs(939)));
    layer2_outputs(861) <= layer1_outputs(1107);
    layer2_outputs(862) <= (layer1_outputs(395)) or (layer1_outputs(288));
    layer2_outputs(863) <= (layer1_outputs(1695)) and not (layer1_outputs(1868));
    layer2_outputs(864) <= not((layer1_outputs(6)) and (layer1_outputs(672)));
    layer2_outputs(865) <= layer1_outputs(2245);
    layer2_outputs(866) <= not(layer1_outputs(650));
    layer2_outputs(867) <= not(layer1_outputs(1208));
    layer2_outputs(868) <= not(layer1_outputs(6)) or (layer1_outputs(752));
    layer2_outputs(869) <= not(layer1_outputs(892));
    layer2_outputs(870) <= layer1_outputs(866);
    layer2_outputs(871) <= layer1_outputs(1072);
    layer2_outputs(872) <= not((layer1_outputs(785)) or (layer1_outputs(658)));
    layer2_outputs(873) <= layer1_outputs(93);
    layer2_outputs(874) <= (layer1_outputs(340)) and not (layer1_outputs(1680));
    layer2_outputs(875) <= layer1_outputs(2226);
    layer2_outputs(876) <= layer1_outputs(436);
    layer2_outputs(877) <= layer1_outputs(1936);
    layer2_outputs(878) <= not(layer1_outputs(431)) or (layer1_outputs(1399));
    layer2_outputs(879) <= (layer1_outputs(2304)) or (layer1_outputs(2118));
    layer2_outputs(880) <= layer1_outputs(485);
    layer2_outputs(881) <= (layer1_outputs(303)) and (layer1_outputs(1385));
    layer2_outputs(882) <= not(layer1_outputs(928)) or (layer1_outputs(982));
    layer2_outputs(883) <= not(layer1_outputs(1442));
    layer2_outputs(884) <= (layer1_outputs(231)) and not (layer1_outputs(2365));
    layer2_outputs(885) <= layer1_outputs(169);
    layer2_outputs(886) <= (layer1_outputs(2112)) and not (layer1_outputs(2505));
    layer2_outputs(887) <= not((layer1_outputs(2454)) and (layer1_outputs(1049)));
    layer2_outputs(888) <= not(layer1_outputs(123));
    layer2_outputs(889) <= not(layer1_outputs(1840));
    layer2_outputs(890) <= not((layer1_outputs(1996)) or (layer1_outputs(2138)));
    layer2_outputs(891) <= not(layer1_outputs(1897));
    layer2_outputs(892) <= not(layer1_outputs(1942));
    layer2_outputs(893) <= not(layer1_outputs(1086));
    layer2_outputs(894) <= not(layer1_outputs(167));
    layer2_outputs(895) <= not((layer1_outputs(15)) and (layer1_outputs(301)));
    layer2_outputs(896) <= (layer1_outputs(1820)) and not (layer1_outputs(2063));
    layer2_outputs(897) <= (layer1_outputs(1355)) and (layer1_outputs(1146));
    layer2_outputs(898) <= not(layer1_outputs(1289));
    layer2_outputs(899) <= not(layer1_outputs(400));
    layer2_outputs(900) <= not((layer1_outputs(2476)) and (layer1_outputs(1744)));
    layer2_outputs(901) <= not((layer1_outputs(2078)) xor (layer1_outputs(1473)));
    layer2_outputs(902) <= layer1_outputs(1550);
    layer2_outputs(903) <= not(layer1_outputs(810));
    layer2_outputs(904) <= layer1_outputs(1561);
    layer2_outputs(905) <= (layer1_outputs(2410)) or (layer1_outputs(137));
    layer2_outputs(906) <= not(layer1_outputs(847));
    layer2_outputs(907) <= not(layer1_outputs(1879));
    layer2_outputs(908) <= (layer1_outputs(2281)) and not (layer1_outputs(2159));
    layer2_outputs(909) <= layer1_outputs(2180);
    layer2_outputs(910) <= (layer1_outputs(2071)) and (layer1_outputs(2441));
    layer2_outputs(911) <= layer1_outputs(935);
    layer2_outputs(912) <= (layer1_outputs(2442)) and (layer1_outputs(1845));
    layer2_outputs(913) <= (layer1_outputs(244)) and (layer1_outputs(1041));
    layer2_outputs(914) <= not(layer1_outputs(1944));
    layer2_outputs(915) <= not(layer1_outputs(1749));
    layer2_outputs(916) <= layer1_outputs(682);
    layer2_outputs(917) <= (layer1_outputs(965)) or (layer1_outputs(487));
    layer2_outputs(918) <= (layer1_outputs(2511)) and not (layer1_outputs(255));
    layer2_outputs(919) <= not((layer1_outputs(786)) or (layer1_outputs(904)));
    layer2_outputs(920) <= (layer1_outputs(889)) and (layer1_outputs(417));
    layer2_outputs(921) <= (layer1_outputs(2053)) and not (layer1_outputs(516));
    layer2_outputs(922) <= (layer1_outputs(1313)) and (layer1_outputs(2543));
    layer2_outputs(923) <= layer1_outputs(1915);
    layer2_outputs(924) <= (layer1_outputs(276)) or (layer1_outputs(670));
    layer2_outputs(925) <= not((layer1_outputs(1040)) xor (layer1_outputs(1084)));
    layer2_outputs(926) <= not((layer1_outputs(1838)) or (layer1_outputs(1845)));
    layer2_outputs(927) <= (layer1_outputs(2440)) and not (layer1_outputs(318));
    layer2_outputs(928) <= (layer1_outputs(2545)) and (layer1_outputs(723));
    layer2_outputs(929) <= not((layer1_outputs(1718)) xor (layer1_outputs(2316)));
    layer2_outputs(930) <= (layer1_outputs(320)) or (layer1_outputs(2516));
    layer2_outputs(931) <= not(layer1_outputs(1496));
    layer2_outputs(932) <= not(layer1_outputs(1703));
    layer2_outputs(933) <= not(layer1_outputs(1548)) or (layer1_outputs(2319));
    layer2_outputs(934) <= layer1_outputs(2026);
    layer2_outputs(935) <= not((layer1_outputs(1462)) and (layer1_outputs(521)));
    layer2_outputs(936) <= (layer1_outputs(205)) or (layer1_outputs(1805));
    layer2_outputs(937) <= not(layer1_outputs(1392));
    layer2_outputs(938) <= (layer1_outputs(2202)) or (layer1_outputs(1903));
    layer2_outputs(939) <= (layer1_outputs(1045)) and (layer1_outputs(2040));
    layer2_outputs(940) <= layer1_outputs(1023);
    layer2_outputs(941) <= not(layer1_outputs(1530));
    layer2_outputs(942) <= not(layer1_outputs(1094));
    layer2_outputs(943) <= layer1_outputs(1171);
    layer2_outputs(944) <= not((layer1_outputs(1502)) and (layer1_outputs(1135)));
    layer2_outputs(945) <= (layer1_outputs(1165)) and not (layer1_outputs(2436));
    layer2_outputs(946) <= not((layer1_outputs(2154)) and (layer1_outputs(1221)));
    layer2_outputs(947) <= (layer1_outputs(2120)) and (layer1_outputs(501));
    layer2_outputs(948) <= (layer1_outputs(403)) xor (layer1_outputs(1259));
    layer2_outputs(949) <= (layer1_outputs(1628)) or (layer1_outputs(1011));
    layer2_outputs(950) <= not(layer1_outputs(570));
    layer2_outputs(951) <= not(layer1_outputs(239)) or (layer1_outputs(862));
    layer2_outputs(952) <= not((layer1_outputs(73)) and (layer1_outputs(631)));
    layer2_outputs(953) <= not((layer1_outputs(1687)) or (layer1_outputs(2149)));
    layer2_outputs(954) <= not(layer1_outputs(881));
    layer2_outputs(955) <= not(layer1_outputs(622));
    layer2_outputs(956) <= layer1_outputs(648);
    layer2_outputs(957) <= layer1_outputs(647);
    layer2_outputs(958) <= not(layer1_outputs(901));
    layer2_outputs(959) <= not((layer1_outputs(158)) or (layer1_outputs(1605)));
    layer2_outputs(960) <= not(layer1_outputs(1631));
    layer2_outputs(961) <= not((layer1_outputs(1499)) or (layer1_outputs(301)));
    layer2_outputs(962) <= layer1_outputs(855);
    layer2_outputs(963) <= (layer1_outputs(1999)) or (layer1_outputs(1284));
    layer2_outputs(964) <= (layer1_outputs(1956)) and (layer1_outputs(855));
    layer2_outputs(965) <= not(layer1_outputs(1616));
    layer2_outputs(966) <= layer1_outputs(1792);
    layer2_outputs(967) <= (layer1_outputs(336)) and not (layer1_outputs(513));
    layer2_outputs(968) <= not(layer1_outputs(1995));
    layer2_outputs(969) <= (layer1_outputs(1173)) and (layer1_outputs(921));
    layer2_outputs(970) <= not(layer1_outputs(372)) or (layer1_outputs(416));
    layer2_outputs(971) <= not((layer1_outputs(903)) and (layer1_outputs(1865)));
    layer2_outputs(972) <= layer1_outputs(48);
    layer2_outputs(973) <= not(layer1_outputs(1163));
    layer2_outputs(974) <= layer1_outputs(815);
    layer2_outputs(975) <= (layer1_outputs(1615)) and not (layer1_outputs(739));
    layer2_outputs(976) <= (layer1_outputs(1165)) and not (layer1_outputs(276));
    layer2_outputs(977) <= not(layer1_outputs(1281));
    layer2_outputs(978) <= '0';
    layer2_outputs(979) <= (layer1_outputs(1840)) or (layer1_outputs(1072));
    layer2_outputs(980) <= not(layer1_outputs(920));
    layer2_outputs(981) <= not((layer1_outputs(2464)) and (layer1_outputs(2545)));
    layer2_outputs(982) <= (layer1_outputs(2130)) or (layer1_outputs(1116));
    layer2_outputs(983) <= (layer1_outputs(756)) or (layer1_outputs(837));
    layer2_outputs(984) <= (layer1_outputs(1521)) or (layer1_outputs(1005));
    layer2_outputs(985) <= not(layer1_outputs(1788));
    layer2_outputs(986) <= layer1_outputs(2514);
    layer2_outputs(987) <= layer1_outputs(812);
    layer2_outputs(988) <= (layer1_outputs(360)) and not (layer1_outputs(1759));
    layer2_outputs(989) <= layer1_outputs(938);
    layer2_outputs(990) <= not(layer1_outputs(2108));
    layer2_outputs(991) <= layer1_outputs(2084);
    layer2_outputs(992) <= not(layer1_outputs(1501));
    layer2_outputs(993) <= not(layer1_outputs(174)) or (layer1_outputs(1884));
    layer2_outputs(994) <= not((layer1_outputs(332)) and (layer1_outputs(788)));
    layer2_outputs(995) <= not(layer1_outputs(2386));
    layer2_outputs(996) <= not(layer1_outputs(1132)) or (layer1_outputs(1467));
    layer2_outputs(997) <= not(layer1_outputs(2065));
    layer2_outputs(998) <= layer1_outputs(997);
    layer2_outputs(999) <= not(layer1_outputs(1459));
    layer2_outputs(1000) <= not(layer1_outputs(1928));
    layer2_outputs(1001) <= not(layer1_outputs(1419));
    layer2_outputs(1002) <= not(layer1_outputs(1061));
    layer2_outputs(1003) <= not(layer1_outputs(439));
    layer2_outputs(1004) <= '0';
    layer2_outputs(1005) <= (layer1_outputs(134)) and not (layer1_outputs(222));
    layer2_outputs(1006) <= layer1_outputs(1282);
    layer2_outputs(1007) <= (layer1_outputs(2364)) and (layer1_outputs(1139));
    layer2_outputs(1008) <= layer1_outputs(442);
    layer2_outputs(1009) <= layer1_outputs(460);
    layer2_outputs(1010) <= layer1_outputs(2086);
    layer2_outputs(1011) <= layer1_outputs(159);
    layer2_outputs(1012) <= not(layer1_outputs(2149));
    layer2_outputs(1013) <= layer1_outputs(2213);
    layer2_outputs(1014) <= not(layer1_outputs(241)) or (layer1_outputs(152));
    layer2_outputs(1015) <= not(layer1_outputs(1532));
    layer2_outputs(1016) <= not(layer1_outputs(1897)) or (layer1_outputs(1376));
    layer2_outputs(1017) <= (layer1_outputs(1033)) and (layer1_outputs(886));
    layer2_outputs(1018) <= not((layer1_outputs(1658)) or (layer1_outputs(202)));
    layer2_outputs(1019) <= not(layer1_outputs(211)) or (layer1_outputs(596));
    layer2_outputs(1020) <= (layer1_outputs(1556)) and not (layer1_outputs(650));
    layer2_outputs(1021) <= (layer1_outputs(2369)) or (layer1_outputs(1472));
    layer2_outputs(1022) <= not((layer1_outputs(245)) or (layer1_outputs(2438)));
    layer2_outputs(1023) <= (layer1_outputs(10)) and not (layer1_outputs(906));
    layer2_outputs(1024) <= layer1_outputs(88);
    layer2_outputs(1025) <= layer1_outputs(1901);
    layer2_outputs(1026) <= '0';
    layer2_outputs(1027) <= not((layer1_outputs(62)) xor (layer1_outputs(1824)));
    layer2_outputs(1028) <= not(layer1_outputs(1700)) or (layer1_outputs(1444));
    layer2_outputs(1029) <= layer1_outputs(1547);
    layer2_outputs(1030) <= layer1_outputs(2258);
    layer2_outputs(1031) <= not(layer1_outputs(2479)) or (layer1_outputs(1282));
    layer2_outputs(1032) <= not(layer1_outputs(1037));
    layer2_outputs(1033) <= (layer1_outputs(656)) and not (layer1_outputs(2216));
    layer2_outputs(1034) <= layer1_outputs(75);
    layer2_outputs(1035) <= not(layer1_outputs(19));
    layer2_outputs(1036) <= not((layer1_outputs(1675)) and (layer1_outputs(2235)));
    layer2_outputs(1037) <= (layer1_outputs(257)) and (layer1_outputs(299));
    layer2_outputs(1038) <= not(layer1_outputs(635));
    layer2_outputs(1039) <= '0';
    layer2_outputs(1040) <= not(layer1_outputs(956));
    layer2_outputs(1041) <= not((layer1_outputs(2009)) or (layer1_outputs(1410)));
    layer2_outputs(1042) <= not(layer1_outputs(2212)) or (layer1_outputs(1353));
    layer2_outputs(1043) <= not(layer1_outputs(513));
    layer2_outputs(1044) <= not(layer1_outputs(290)) or (layer1_outputs(2242));
    layer2_outputs(1045) <= not(layer1_outputs(1741));
    layer2_outputs(1046) <= not(layer1_outputs(2106)) or (layer1_outputs(238));
    layer2_outputs(1047) <= (layer1_outputs(45)) and not (layer1_outputs(2372));
    layer2_outputs(1048) <= (layer1_outputs(2025)) and not (layer1_outputs(1857));
    layer2_outputs(1049) <= (layer1_outputs(1704)) and not (layer1_outputs(95));
    layer2_outputs(1050) <= (layer1_outputs(600)) and not (layer1_outputs(1669));
    layer2_outputs(1051) <= (layer1_outputs(385)) and not (layer1_outputs(474));
    layer2_outputs(1052) <= not(layer1_outputs(1829));
    layer2_outputs(1053) <= layer1_outputs(1575);
    layer2_outputs(1054) <= not(layer1_outputs(1835)) or (layer1_outputs(1713));
    layer2_outputs(1055) <= not(layer1_outputs(713)) or (layer1_outputs(1479));
    layer2_outputs(1056) <= not(layer1_outputs(1946));
    layer2_outputs(1057) <= layer1_outputs(2127);
    layer2_outputs(1058) <= layer1_outputs(871);
    layer2_outputs(1059) <= layer1_outputs(1912);
    layer2_outputs(1060) <= not(layer1_outputs(532));
    layer2_outputs(1061) <= not(layer1_outputs(532)) or (layer1_outputs(761));
    layer2_outputs(1062) <= not(layer1_outputs(109));
    layer2_outputs(1063) <= not(layer1_outputs(1039));
    layer2_outputs(1064) <= (layer1_outputs(583)) and (layer1_outputs(1039));
    layer2_outputs(1065) <= (layer1_outputs(1655)) and not (layer1_outputs(1597));
    layer2_outputs(1066) <= (layer1_outputs(1092)) and not (layer1_outputs(1195));
    layer2_outputs(1067) <= not((layer1_outputs(2291)) xor (layer1_outputs(943)));
    layer2_outputs(1068) <= not((layer1_outputs(1790)) or (layer1_outputs(1879)));
    layer2_outputs(1069) <= (layer1_outputs(515)) and not (layer1_outputs(1491));
    layer2_outputs(1070) <= not(layer1_outputs(245));
    layer2_outputs(1071) <= (layer1_outputs(181)) and not (layer1_outputs(1821));
    layer2_outputs(1072) <= not(layer1_outputs(1060));
    layer2_outputs(1073) <= not((layer1_outputs(785)) xor (layer1_outputs(1783)));
    layer2_outputs(1074) <= layer1_outputs(1417);
    layer2_outputs(1075) <= not(layer1_outputs(2094)) or (layer1_outputs(803));
    layer2_outputs(1076) <= layer1_outputs(184);
    layer2_outputs(1077) <= not(layer1_outputs(1764)) or (layer1_outputs(1230));
    layer2_outputs(1078) <= layer1_outputs(237);
    layer2_outputs(1079) <= layer1_outputs(666);
    layer2_outputs(1080) <= layer1_outputs(223);
    layer2_outputs(1081) <= not(layer1_outputs(1810)) or (layer1_outputs(1048));
    layer2_outputs(1082) <= not(layer1_outputs(214));
    layer2_outputs(1083) <= (layer1_outputs(1488)) and not (layer1_outputs(2327));
    layer2_outputs(1084) <= (layer1_outputs(2087)) and not (layer1_outputs(827));
    layer2_outputs(1085) <= (layer1_outputs(2150)) and not (layer1_outputs(1650));
    layer2_outputs(1086) <= not((layer1_outputs(1648)) and (layer1_outputs(2075)));
    layer2_outputs(1087) <= not(layer1_outputs(1509));
    layer2_outputs(1088) <= not((layer1_outputs(2337)) and (layer1_outputs(2230)));
    layer2_outputs(1089) <= not(layer1_outputs(1934));
    layer2_outputs(1090) <= layer1_outputs(2382);
    layer2_outputs(1091) <= not(layer1_outputs(297));
    layer2_outputs(1092) <= layer1_outputs(1711);
    layer2_outputs(1093) <= layer1_outputs(814);
    layer2_outputs(1094) <= not((layer1_outputs(72)) and (layer1_outputs(1740)));
    layer2_outputs(1095) <= not(layer1_outputs(1358)) or (layer1_outputs(949));
    layer2_outputs(1096) <= not((layer1_outputs(120)) and (layer1_outputs(2125)));
    layer2_outputs(1097) <= layer1_outputs(1013);
    layer2_outputs(1098) <= not(layer1_outputs(1657));
    layer2_outputs(1099) <= not(layer1_outputs(253)) or (layer1_outputs(2307));
    layer2_outputs(1100) <= (layer1_outputs(1552)) and not (layer1_outputs(2475));
    layer2_outputs(1101) <= (layer1_outputs(2541)) and not (layer1_outputs(2359));
    layer2_outputs(1102) <= (layer1_outputs(1280)) xor (layer1_outputs(740));
    layer2_outputs(1103) <= '1';
    layer2_outputs(1104) <= not(layer1_outputs(1077));
    layer2_outputs(1105) <= layer1_outputs(924);
    layer2_outputs(1106) <= not(layer1_outputs(692)) or (layer1_outputs(1873));
    layer2_outputs(1107) <= not(layer1_outputs(189)) or (layer1_outputs(2214));
    layer2_outputs(1108) <= not(layer1_outputs(837));
    layer2_outputs(1109) <= not((layer1_outputs(223)) or (layer1_outputs(186)));
    layer2_outputs(1110) <= not((layer1_outputs(1563)) or (layer1_outputs(2142)));
    layer2_outputs(1111) <= (layer1_outputs(2379)) and not (layer1_outputs(1540));
    layer2_outputs(1112) <= layer1_outputs(1277);
    layer2_outputs(1113) <= not(layer1_outputs(2215));
    layer2_outputs(1114) <= (layer1_outputs(64)) and not (layer1_outputs(1966));
    layer2_outputs(1115) <= (layer1_outputs(1608)) and not (layer1_outputs(829));
    layer2_outputs(1116) <= (layer1_outputs(1150)) and not (layer1_outputs(226));
    layer2_outputs(1117) <= layer1_outputs(193);
    layer2_outputs(1118) <= not(layer1_outputs(419));
    layer2_outputs(1119) <= not(layer1_outputs(1137)) or (layer1_outputs(1115));
    layer2_outputs(1120) <= (layer1_outputs(441)) and (layer1_outputs(172));
    layer2_outputs(1121) <= not(layer1_outputs(1795));
    layer2_outputs(1122) <= layer1_outputs(417);
    layer2_outputs(1123) <= layer1_outputs(348);
    layer2_outputs(1124) <= (layer1_outputs(1931)) and not (layer1_outputs(2401));
    layer2_outputs(1125) <= not(layer1_outputs(595));
    layer2_outputs(1126) <= (layer1_outputs(2302)) or (layer1_outputs(1567));
    layer2_outputs(1127) <= (layer1_outputs(2097)) or (layer1_outputs(1920));
    layer2_outputs(1128) <= (layer1_outputs(1302)) and not (layer1_outputs(481));
    layer2_outputs(1129) <= not((layer1_outputs(448)) or (layer1_outputs(1173)));
    layer2_outputs(1130) <= layer1_outputs(902);
    layer2_outputs(1131) <= not((layer1_outputs(2559)) or (layer1_outputs(1189)));
    layer2_outputs(1132) <= not(layer1_outputs(46)) or (layer1_outputs(694));
    layer2_outputs(1133) <= not((layer1_outputs(1339)) and (layer1_outputs(1388)));
    layer2_outputs(1134) <= (layer1_outputs(370)) and (layer1_outputs(2235));
    layer2_outputs(1135) <= not(layer1_outputs(66)) or (layer1_outputs(1761));
    layer2_outputs(1136) <= not((layer1_outputs(119)) and (layer1_outputs(2285)));
    layer2_outputs(1137) <= not(layer1_outputs(87)) or (layer1_outputs(2500));
    layer2_outputs(1138) <= not(layer1_outputs(364));
    layer2_outputs(1139) <= not((layer1_outputs(42)) and (layer1_outputs(1729)));
    layer2_outputs(1140) <= (layer1_outputs(395)) xor (layer1_outputs(1529));
    layer2_outputs(1141) <= (layer1_outputs(1533)) and not (layer1_outputs(1688));
    layer2_outputs(1142) <= not(layer1_outputs(2523)) or (layer1_outputs(2512));
    layer2_outputs(1143) <= not(layer1_outputs(465));
    layer2_outputs(1144) <= not(layer1_outputs(614)) or (layer1_outputs(1677));
    layer2_outputs(1145) <= layer1_outputs(1109);
    layer2_outputs(1146) <= layer1_outputs(1815);
    layer2_outputs(1147) <= not(layer1_outputs(1799));
    layer2_outputs(1148) <= not(layer1_outputs(1640)) or (layer1_outputs(51));
    layer2_outputs(1149) <= '0';
    layer2_outputs(1150) <= not((layer1_outputs(1760)) xor (layer1_outputs(2195)));
    layer2_outputs(1151) <= not(layer1_outputs(802));
    layer2_outputs(1152) <= (layer1_outputs(1158)) and (layer1_outputs(751));
    layer2_outputs(1153) <= not(layer1_outputs(1066));
    layer2_outputs(1154) <= layer1_outputs(2466);
    layer2_outputs(1155) <= layer1_outputs(494);
    layer2_outputs(1156) <= (layer1_outputs(114)) and not (layer1_outputs(360));
    layer2_outputs(1157) <= layer1_outputs(1333);
    layer2_outputs(1158) <= not(layer1_outputs(1874));
    layer2_outputs(1159) <= layer1_outputs(734);
    layer2_outputs(1160) <= not(layer1_outputs(651));
    layer2_outputs(1161) <= layer1_outputs(1799);
    layer2_outputs(1162) <= not(layer1_outputs(2185)) or (layer1_outputs(357));
    layer2_outputs(1163) <= layer1_outputs(1882);
    layer2_outputs(1164) <= '1';
    layer2_outputs(1165) <= (layer1_outputs(227)) and not (layer1_outputs(1959));
    layer2_outputs(1166) <= not((layer1_outputs(2107)) or (layer1_outputs(1206)));
    layer2_outputs(1167) <= layer1_outputs(254);
    layer2_outputs(1168) <= not(layer1_outputs(2210));
    layer2_outputs(1169) <= not(layer1_outputs(1649)) or (layer1_outputs(180));
    layer2_outputs(1170) <= layer1_outputs(787);
    layer2_outputs(1171) <= layer1_outputs(1634);
    layer2_outputs(1172) <= not((layer1_outputs(2113)) xor (layer1_outputs(1886)));
    layer2_outputs(1173) <= not(layer1_outputs(2536));
    layer2_outputs(1174) <= layer1_outputs(1485);
    layer2_outputs(1175) <= not(layer1_outputs(216));
    layer2_outputs(1176) <= not(layer1_outputs(1796));
    layer2_outputs(1177) <= not(layer1_outputs(1952));
    layer2_outputs(1178) <= not(layer1_outputs(1070));
    layer2_outputs(1179) <= not(layer1_outputs(20));
    layer2_outputs(1180) <= not(layer1_outputs(613));
    layer2_outputs(1181) <= not(layer1_outputs(71));
    layer2_outputs(1182) <= layer1_outputs(405);
    layer2_outputs(1183) <= (layer1_outputs(1081)) and not (layer1_outputs(2455));
    layer2_outputs(1184) <= not(layer1_outputs(2432));
    layer2_outputs(1185) <= (layer1_outputs(1802)) and (layer1_outputs(1316));
    layer2_outputs(1186) <= (layer1_outputs(1185)) and (layer1_outputs(313));
    layer2_outputs(1187) <= not(layer1_outputs(211)) or (layer1_outputs(1785));
    layer2_outputs(1188) <= not(layer1_outputs(793)) or (layer1_outputs(1938));
    layer2_outputs(1189) <= (layer1_outputs(1976)) or (layer1_outputs(263));
    layer2_outputs(1190) <= not(layer1_outputs(1808));
    layer2_outputs(1191) <= not((layer1_outputs(673)) and (layer1_outputs(1652)));
    layer2_outputs(1192) <= not(layer1_outputs(1382));
    layer2_outputs(1193) <= not(layer1_outputs(489));
    layer2_outputs(1194) <= not((layer1_outputs(956)) xor (layer1_outputs(1508)));
    layer2_outputs(1195) <= layer1_outputs(375);
    layer2_outputs(1196) <= (layer1_outputs(304)) xor (layer1_outputs(1742));
    layer2_outputs(1197) <= not(layer1_outputs(143)) or (layer1_outputs(926));
    layer2_outputs(1198) <= not(layer1_outputs(1112));
    layer2_outputs(1199) <= not(layer1_outputs(1858)) or (layer1_outputs(2105));
    layer2_outputs(1200) <= not(layer1_outputs(2006)) or (layer1_outputs(769));
    layer2_outputs(1201) <= not(layer1_outputs(71));
    layer2_outputs(1202) <= not(layer1_outputs(822));
    layer2_outputs(1203) <= not(layer1_outputs(666));
    layer2_outputs(1204) <= not(layer1_outputs(283));
    layer2_outputs(1205) <= layer1_outputs(2309);
    layer2_outputs(1206) <= not(layer1_outputs(458));
    layer2_outputs(1207) <= layer1_outputs(195);
    layer2_outputs(1208) <= not(layer1_outputs(434));
    layer2_outputs(1209) <= not(layer1_outputs(2148));
    layer2_outputs(1210) <= layer1_outputs(78);
    layer2_outputs(1211) <= not(layer1_outputs(2457));
    layer2_outputs(1212) <= not(layer1_outputs(2003));
    layer2_outputs(1213) <= (layer1_outputs(592)) xor (layer1_outputs(1545));
    layer2_outputs(1214) <= not((layer1_outputs(578)) or (layer1_outputs(588)));
    layer2_outputs(1215) <= layer1_outputs(1468);
    layer2_outputs(1216) <= (layer1_outputs(754)) and not (layer1_outputs(38));
    layer2_outputs(1217) <= (layer1_outputs(1962)) and (layer1_outputs(1169));
    layer2_outputs(1218) <= (layer1_outputs(2389)) or (layer1_outputs(538));
    layer2_outputs(1219) <= (layer1_outputs(1774)) xor (layer1_outputs(377));
    layer2_outputs(1220) <= not(layer1_outputs(2307)) or (layer1_outputs(2321));
    layer2_outputs(1221) <= (layer1_outputs(2334)) and not (layer1_outputs(1413));
    layer2_outputs(1222) <= not(layer1_outputs(1884));
    layer2_outputs(1223) <= (layer1_outputs(1225)) or (layer1_outputs(2550));
    layer2_outputs(1224) <= not(layer1_outputs(2318));
    layer2_outputs(1225) <= layer1_outputs(637);
    layer2_outputs(1226) <= (layer1_outputs(1238)) and not (layer1_outputs(1517));
    layer2_outputs(1227) <= not(layer1_outputs(659));
    layer2_outputs(1228) <= not(layer1_outputs(1998));
    layer2_outputs(1229) <= layer1_outputs(300);
    layer2_outputs(1230) <= not(layer1_outputs(285));
    layer2_outputs(1231) <= (layer1_outputs(1858)) and not (layer1_outputs(2116));
    layer2_outputs(1232) <= (layer1_outputs(2397)) or (layer1_outputs(1773));
    layer2_outputs(1233) <= not(layer1_outputs(1241));
    layer2_outputs(1234) <= not(layer1_outputs(1770)) or (layer1_outputs(967));
    layer2_outputs(1235) <= not((layer1_outputs(876)) or (layer1_outputs(2553)));
    layer2_outputs(1236) <= not(layer1_outputs(845));
    layer2_outputs(1237) <= not(layer1_outputs(773));
    layer2_outputs(1238) <= not(layer1_outputs(1028)) or (layer1_outputs(733));
    layer2_outputs(1239) <= not(layer1_outputs(477)) or (layer1_outputs(678));
    layer2_outputs(1240) <= (layer1_outputs(1641)) or (layer1_outputs(1849));
    layer2_outputs(1241) <= layer1_outputs(269);
    layer2_outputs(1242) <= (layer1_outputs(1151)) and not (layer1_outputs(1126));
    layer2_outputs(1243) <= not((layer1_outputs(2504)) or (layer1_outputs(479)));
    layer2_outputs(1244) <= not((layer1_outputs(475)) or (layer1_outputs(767)));
    layer2_outputs(1245) <= layer1_outputs(28);
    layer2_outputs(1246) <= not(layer1_outputs(149)) or (layer1_outputs(1760));
    layer2_outputs(1247) <= (layer1_outputs(2121)) and not (layer1_outputs(828));
    layer2_outputs(1248) <= layer1_outputs(1630);
    layer2_outputs(1249) <= not(layer1_outputs(1837));
    layer2_outputs(1250) <= not(layer1_outputs(77));
    layer2_outputs(1251) <= not((layer1_outputs(1699)) and (layer1_outputs(1618)));
    layer2_outputs(1252) <= not((layer1_outputs(516)) xor (layer1_outputs(1151)));
    layer2_outputs(1253) <= (layer1_outputs(1684)) and not (layer1_outputs(1532));
    layer2_outputs(1254) <= (layer1_outputs(1270)) and not (layer1_outputs(958));
    layer2_outputs(1255) <= layer1_outputs(116);
    layer2_outputs(1256) <= layer1_outputs(1917);
    layer2_outputs(1257) <= not(layer1_outputs(153));
    layer2_outputs(1258) <= layer1_outputs(607);
    layer2_outputs(1259) <= layer1_outputs(1194);
    layer2_outputs(1260) <= (layer1_outputs(812)) or (layer1_outputs(2397));
    layer2_outputs(1261) <= not(layer1_outputs(2396));
    layer2_outputs(1262) <= not(layer1_outputs(975));
    layer2_outputs(1263) <= not((layer1_outputs(1888)) xor (layer1_outputs(2540)));
    layer2_outputs(1264) <= (layer1_outputs(1297)) and not (layer1_outputs(369));
    layer2_outputs(1265) <= (layer1_outputs(1031)) and (layer1_outputs(139));
    layer2_outputs(1266) <= not(layer1_outputs(602));
    layer2_outputs(1267) <= not(layer1_outputs(1805));
    layer2_outputs(1268) <= layer1_outputs(1082);
    layer2_outputs(1269) <= not(layer1_outputs(976)) or (layer1_outputs(2389));
    layer2_outputs(1270) <= not((layer1_outputs(1368)) or (layer1_outputs(1383)));
    layer2_outputs(1271) <= not(layer1_outputs(1667)) or (layer1_outputs(2111));
    layer2_outputs(1272) <= (layer1_outputs(664)) or (layer1_outputs(1154));
    layer2_outputs(1273) <= not((layer1_outputs(2430)) xor (layer1_outputs(1632)));
    layer2_outputs(1274) <= not(layer1_outputs(2268)) or (layer1_outputs(931));
    layer2_outputs(1275) <= not(layer1_outputs(1372));
    layer2_outputs(1276) <= not(layer1_outputs(981));
    layer2_outputs(1277) <= (layer1_outputs(1485)) or (layer1_outputs(2026));
    layer2_outputs(1278) <= not(layer1_outputs(1017)) or (layer1_outputs(1782));
    layer2_outputs(1279) <= not(layer1_outputs(1889));
    layer2_outputs(1280) <= not(layer1_outputs(1691));
    layer2_outputs(1281) <= (layer1_outputs(2056)) or (layer1_outputs(597));
    layer2_outputs(1282) <= not(layer1_outputs(815));
    layer2_outputs(1283) <= (layer1_outputs(2203)) and not (layer1_outputs(1160));
    layer2_outputs(1284) <= layer1_outputs(2047);
    layer2_outputs(1285) <= layer1_outputs(459);
    layer2_outputs(1286) <= not((layer1_outputs(1204)) or (layer1_outputs(1827)));
    layer2_outputs(1287) <= (layer1_outputs(367)) or (layer1_outputs(2263));
    layer2_outputs(1288) <= not(layer1_outputs(280)) or (layer1_outputs(1278));
    layer2_outputs(1289) <= not(layer1_outputs(866));
    layer2_outputs(1290) <= (layer1_outputs(305)) or (layer1_outputs(2231));
    layer2_outputs(1291) <= not(layer1_outputs(1356));
    layer2_outputs(1292) <= not(layer1_outputs(1796)) or (layer1_outputs(1450));
    layer2_outputs(1293) <= layer1_outputs(1374);
    layer2_outputs(1294) <= not(layer1_outputs(1614)) or (layer1_outputs(708));
    layer2_outputs(1295) <= not(layer1_outputs(1457));
    layer2_outputs(1296) <= not((layer1_outputs(1127)) and (layer1_outputs(1710)));
    layer2_outputs(1297) <= layer1_outputs(2022);
    layer2_outputs(1298) <= not(layer1_outputs(1202)) or (layer1_outputs(966));
    layer2_outputs(1299) <= not((layer1_outputs(435)) and (layer1_outputs(2271)));
    layer2_outputs(1300) <= not(layer1_outputs(1262));
    layer2_outputs(1301) <= not(layer1_outputs(1769));
    layer2_outputs(1302) <= (layer1_outputs(1400)) and not (layer1_outputs(1626));
    layer2_outputs(1303) <= (layer1_outputs(234)) and not (layer1_outputs(1164));
    layer2_outputs(1304) <= (layer1_outputs(1871)) or (layer1_outputs(1412));
    layer2_outputs(1305) <= (layer1_outputs(2531)) and not (layer1_outputs(1364));
    layer2_outputs(1306) <= not((layer1_outputs(2471)) xor (layer1_outputs(2252)));
    layer2_outputs(1307) <= (layer1_outputs(487)) and not (layer1_outputs(251));
    layer2_outputs(1308) <= not(layer1_outputs(512));
    layer2_outputs(1309) <= layer1_outputs(616);
    layer2_outputs(1310) <= not((layer1_outputs(2243)) and (layer1_outputs(992)));
    layer2_outputs(1311) <= layer1_outputs(310);
    layer2_outputs(1312) <= (layer1_outputs(1338)) or (layer1_outputs(468));
    layer2_outputs(1313) <= layer1_outputs(1106);
    layer2_outputs(1314) <= not(layer1_outputs(2072));
    layer2_outputs(1315) <= not(layer1_outputs(81));
    layer2_outputs(1316) <= (layer1_outputs(1226)) and (layer1_outputs(1393));
    layer2_outputs(1317) <= not(layer1_outputs(34)) or (layer1_outputs(2000));
    layer2_outputs(1318) <= not(layer1_outputs(324)) or (layer1_outputs(879));
    layer2_outputs(1319) <= layer1_outputs(780);
    layer2_outputs(1320) <= (layer1_outputs(1190)) or (layer1_outputs(1397));
    layer2_outputs(1321) <= layer1_outputs(1789);
    layer2_outputs(1322) <= layer1_outputs(1422);
    layer2_outputs(1323) <= layer1_outputs(2431);
    layer2_outputs(1324) <= layer1_outputs(1782);
    layer2_outputs(1325) <= (layer1_outputs(41)) and not (layer1_outputs(1657));
    layer2_outputs(1326) <= (layer1_outputs(179)) and (layer1_outputs(1349));
    layer2_outputs(1327) <= (layer1_outputs(2073)) and not (layer1_outputs(2261));
    layer2_outputs(1328) <= not(layer1_outputs(1134));
    layer2_outputs(1329) <= (layer1_outputs(810)) and not (layer1_outputs(442));
    layer2_outputs(1330) <= layer1_outputs(1777);
    layer2_outputs(1331) <= (layer1_outputs(92)) or (layer1_outputs(659));
    layer2_outputs(1332) <= not((layer1_outputs(1854)) and (layer1_outputs(236)));
    layer2_outputs(1333) <= (layer1_outputs(1098)) or (layer1_outputs(2099));
    layer2_outputs(1334) <= not((layer1_outputs(813)) and (layer1_outputs(1625)));
    layer2_outputs(1335) <= layer1_outputs(135);
    layer2_outputs(1336) <= not(layer1_outputs(1227));
    layer2_outputs(1337) <= not(layer1_outputs(406));
    layer2_outputs(1338) <= layer1_outputs(645);
    layer2_outputs(1339) <= (layer1_outputs(45)) and not (layer1_outputs(336));
    layer2_outputs(1340) <= not(layer1_outputs(2165));
    layer2_outputs(1341) <= (layer1_outputs(1973)) and not (layer1_outputs(1226));
    layer2_outputs(1342) <= (layer1_outputs(1728)) and (layer1_outputs(2199));
    layer2_outputs(1343) <= not((layer1_outputs(676)) and (layer1_outputs(1083)));
    layer2_outputs(1344) <= not((layer1_outputs(37)) and (layer1_outputs(1515)));
    layer2_outputs(1345) <= layer1_outputs(2041);
    layer2_outputs(1346) <= (layer1_outputs(1541)) and not (layer1_outputs(502));
    layer2_outputs(1347) <= layer1_outputs(98);
    layer2_outputs(1348) <= not((layer1_outputs(681)) or (layer1_outputs(1543)));
    layer2_outputs(1349) <= layer1_outputs(560);
    layer2_outputs(1350) <= '1';
    layer2_outputs(1351) <= layer1_outputs(1044);
    layer2_outputs(1352) <= not((layer1_outputs(2135)) and (layer1_outputs(883)));
    layer2_outputs(1353) <= (layer1_outputs(676)) and not (layer1_outputs(2396));
    layer2_outputs(1354) <= (layer1_outputs(63)) and (layer1_outputs(1140));
    layer2_outputs(1355) <= layer1_outputs(2068);
    layer2_outputs(1356) <= layer1_outputs(1750);
    layer2_outputs(1357) <= layer1_outputs(875);
    layer2_outputs(1358) <= not(layer1_outputs(2259)) or (layer1_outputs(1306));
    layer2_outputs(1359) <= (layer1_outputs(1232)) and (layer1_outputs(128));
    layer2_outputs(1360) <= not(layer1_outputs(2022)) or (layer1_outputs(698));
    layer2_outputs(1361) <= '0';
    layer2_outputs(1362) <= not(layer1_outputs(2289)) or (layer1_outputs(294));
    layer2_outputs(1363) <= not((layer1_outputs(1883)) or (layer1_outputs(736)));
    layer2_outputs(1364) <= '0';
    layer2_outputs(1365) <= layer1_outputs(309);
    layer2_outputs(1366) <= not((layer1_outputs(1091)) or (layer1_outputs(189)));
    layer2_outputs(1367) <= (layer1_outputs(1487)) xor (layer1_outputs(1317));
    layer2_outputs(1368) <= not(layer1_outputs(1694));
    layer2_outputs(1369) <= (layer1_outputs(2400)) and not (layer1_outputs(2463));
    layer2_outputs(1370) <= not(layer1_outputs(644)) or (layer1_outputs(1523));
    layer2_outputs(1371) <= '1';
    layer2_outputs(1372) <= (layer1_outputs(1357)) xor (layer1_outputs(1637));
    layer2_outputs(1373) <= not(layer1_outputs(1098)) or (layer1_outputs(702));
    layer2_outputs(1374) <= layer1_outputs(826);
    layer2_outputs(1375) <= not((layer1_outputs(1830)) xor (layer1_outputs(799)));
    layer2_outputs(1376) <= layer1_outputs(1225);
    layer2_outputs(1377) <= not((layer1_outputs(133)) xor (layer1_outputs(1366)));
    layer2_outputs(1378) <= layer1_outputs(254);
    layer2_outputs(1379) <= not((layer1_outputs(1082)) and (layer1_outputs(116)));
    layer2_outputs(1380) <= (layer1_outputs(1422)) or (layer1_outputs(540));
    layer2_outputs(1381) <= not(layer1_outputs(790));
    layer2_outputs(1382) <= not(layer1_outputs(53));
    layer2_outputs(1383) <= (layer1_outputs(538)) or (layer1_outputs(737));
    layer2_outputs(1384) <= not((layer1_outputs(1221)) and (layer1_outputs(311)));
    layer2_outputs(1385) <= not(layer1_outputs(1562)) or (layer1_outputs(1576));
    layer2_outputs(1386) <= layer1_outputs(235);
    layer2_outputs(1387) <= (layer1_outputs(1612)) xor (layer1_outputs(912));
    layer2_outputs(1388) <= not(layer1_outputs(1577));
    layer2_outputs(1389) <= not(layer1_outputs(1396));
    layer2_outputs(1390) <= (layer1_outputs(268)) and not (layer1_outputs(2174));
    layer2_outputs(1391) <= layer1_outputs(1188);
    layer2_outputs(1392) <= not(layer1_outputs(783));
    layer2_outputs(1393) <= '1';
    layer2_outputs(1394) <= (layer1_outputs(104)) and (layer1_outputs(847));
    layer2_outputs(1395) <= (layer1_outputs(2250)) and not (layer1_outputs(1022));
    layer2_outputs(1396) <= not((layer1_outputs(1809)) or (layer1_outputs(1486)));
    layer2_outputs(1397) <= not(layer1_outputs(998)) or (layer1_outputs(2405));
    layer2_outputs(1398) <= not(layer1_outputs(1398));
    layer2_outputs(1399) <= not(layer1_outputs(936)) or (layer1_outputs(2530));
    layer2_outputs(1400) <= layer1_outputs(1836);
    layer2_outputs(1401) <= '1';
    layer2_outputs(1402) <= not(layer1_outputs(373)) or (layer1_outputs(1218));
    layer2_outputs(1403) <= not((layer1_outputs(2279)) or (layer1_outputs(677)));
    layer2_outputs(1404) <= layer1_outputs(66);
    layer2_outputs(1405) <= '1';
    layer2_outputs(1406) <= not(layer1_outputs(2240));
    layer2_outputs(1407) <= not(layer1_outputs(2426));
    layer2_outputs(1408) <= not(layer1_outputs(1720));
    layer2_outputs(1409) <= (layer1_outputs(470)) or (layer1_outputs(2382));
    layer2_outputs(1410) <= not(layer1_outputs(130));
    layer2_outputs(1411) <= not(layer1_outputs(1478)) or (layer1_outputs(2163));
    layer2_outputs(1412) <= not(layer1_outputs(1096)) or (layer1_outputs(346));
    layer2_outputs(1413) <= (layer1_outputs(450)) or (layer1_outputs(447));
    layer2_outputs(1414) <= not(layer1_outputs(937));
    layer2_outputs(1415) <= layer1_outputs(1070);
    layer2_outputs(1416) <= (layer1_outputs(556)) and (layer1_outputs(2153));
    layer2_outputs(1417) <= (layer1_outputs(1717)) and not (layer1_outputs(762));
    layer2_outputs(1418) <= not((layer1_outputs(2478)) and (layer1_outputs(490)));
    layer2_outputs(1419) <= not(layer1_outputs(2402));
    layer2_outputs(1420) <= (layer1_outputs(1903)) or (layer1_outputs(1335));
    layer2_outputs(1421) <= not(layer1_outputs(399));
    layer2_outputs(1422) <= not(layer1_outputs(2506));
    layer2_outputs(1423) <= (layer1_outputs(2355)) and not (layer1_outputs(2497));
    layer2_outputs(1424) <= (layer1_outputs(995)) or (layer1_outputs(717));
    layer2_outputs(1425) <= (layer1_outputs(331)) and not (layer1_outputs(1415));
    layer2_outputs(1426) <= not(layer1_outputs(2315));
    layer2_outputs(1427) <= (layer1_outputs(639)) and not (layer1_outputs(766));
    layer2_outputs(1428) <= not((layer1_outputs(594)) and (layer1_outputs(1095)));
    layer2_outputs(1429) <= not(layer1_outputs(61));
    layer2_outputs(1430) <= not(layer1_outputs(1813)) or (layer1_outputs(1230));
    layer2_outputs(1431) <= (layer1_outputs(969)) and (layer1_outputs(1125));
    layer2_outputs(1432) <= (layer1_outputs(1900)) or (layer1_outputs(1969));
    layer2_outputs(1433) <= not(layer1_outputs(742));
    layer2_outputs(1434) <= layer1_outputs(735);
    layer2_outputs(1435) <= layer1_outputs(1947);
    layer2_outputs(1436) <= not((layer1_outputs(2215)) and (layer1_outputs(509)));
    layer2_outputs(1437) <= not(layer1_outputs(1766));
    layer2_outputs(1438) <= layer1_outputs(1159);
    layer2_outputs(1439) <= not((layer1_outputs(1239)) or (layer1_outputs(746)));
    layer2_outputs(1440) <= layer1_outputs(215);
    layer2_outputs(1441) <= (layer1_outputs(2469)) and (layer1_outputs(2001));
    layer2_outputs(1442) <= not(layer1_outputs(1236));
    layer2_outputs(1443) <= not(layer1_outputs(2138));
    layer2_outputs(1444) <= layer1_outputs(492);
    layer2_outputs(1445) <= not(layer1_outputs(151)) or (layer1_outputs(1222));
    layer2_outputs(1446) <= (layer1_outputs(190)) and (layer1_outputs(1107));
    layer2_outputs(1447) <= (layer1_outputs(1992)) and (layer1_outputs(314));
    layer2_outputs(1448) <= (layer1_outputs(2123)) xor (layer1_outputs(579));
    layer2_outputs(1449) <= (layer1_outputs(1090)) or (layer1_outputs(852));
    layer2_outputs(1450) <= not((layer1_outputs(290)) and (layer1_outputs(2060)));
    layer2_outputs(1451) <= layer1_outputs(51);
    layer2_outputs(1452) <= not(layer1_outputs(611));
    layer2_outputs(1453) <= not(layer1_outputs(945));
    layer2_outputs(1454) <= layer1_outputs(1020);
    layer2_outputs(1455) <= (layer1_outputs(835)) and not (layer1_outputs(2324));
    layer2_outputs(1456) <= (layer1_outputs(1941)) and (layer1_outputs(1046));
    layer2_outputs(1457) <= '0';
    layer2_outputs(1458) <= not(layer1_outputs(2001));
    layer2_outputs(1459) <= not(layer1_outputs(2131));
    layer2_outputs(1460) <= '0';
    layer2_outputs(1461) <= (layer1_outputs(410)) and not (layer1_outputs(977));
    layer2_outputs(1462) <= layer1_outputs(448);
    layer2_outputs(1463) <= layer1_outputs(862);
    layer2_outputs(1464) <= not((layer1_outputs(1590)) xor (layer1_outputs(2256)));
    layer2_outputs(1465) <= (layer1_outputs(199)) and (layer1_outputs(1963));
    layer2_outputs(1466) <= layer1_outputs(1365);
    layer2_outputs(1467) <= layer1_outputs(1433);
    layer2_outputs(1468) <= '0';
    layer2_outputs(1469) <= not(layer1_outputs(378)) or (layer1_outputs(32));
    layer2_outputs(1470) <= layer1_outputs(1787);
    layer2_outputs(1471) <= not(layer1_outputs(908));
    layer2_outputs(1472) <= layer1_outputs(152);
    layer2_outputs(1473) <= layer1_outputs(2029);
    layer2_outputs(1474) <= (layer1_outputs(2258)) or (layer1_outputs(2301));
    layer2_outputs(1475) <= '0';
    layer2_outputs(1476) <= layer1_outputs(851);
    layer2_outputs(1477) <= not(layer1_outputs(1011));
    layer2_outputs(1478) <= (layer1_outputs(1397)) and not (layer1_outputs(2217));
    layer2_outputs(1479) <= (layer1_outputs(542)) or (layer1_outputs(842));
    layer2_outputs(1480) <= not((layer1_outputs(1673)) or (layer1_outputs(2462)));
    layer2_outputs(1481) <= (layer1_outputs(1853)) and not (layer1_outputs(1365));
    layer2_outputs(1482) <= not((layer1_outputs(1935)) or (layer1_outputs(1222)));
    layer2_outputs(1483) <= '0';
    layer2_outputs(1484) <= (layer1_outputs(275)) or (layer1_outputs(2054));
    layer2_outputs(1485) <= not(layer1_outputs(1843));
    layer2_outputs(1486) <= not(layer1_outputs(776));
    layer2_outputs(1487) <= not(layer1_outputs(1950));
    layer2_outputs(1488) <= not(layer1_outputs(1856)) or (layer1_outputs(1351));
    layer2_outputs(1489) <= not(layer1_outputs(2134));
    layer2_outputs(1490) <= (layer1_outputs(1281)) and not (layer1_outputs(1167));
    layer2_outputs(1491) <= (layer1_outputs(1409)) and not (layer1_outputs(1390));
    layer2_outputs(1492) <= not(layer1_outputs(1628));
    layer2_outputs(1493) <= (layer1_outputs(624)) and (layer1_outputs(1818));
    layer2_outputs(1494) <= not(layer1_outputs(13)) or (layer1_outputs(2322));
    layer2_outputs(1495) <= not(layer1_outputs(1295));
    layer2_outputs(1496) <= layer1_outputs(780);
    layer2_outputs(1497) <= layer1_outputs(1258);
    layer2_outputs(1498) <= not(layer1_outputs(1576)) or (layer1_outputs(552));
    layer2_outputs(1499) <= (layer1_outputs(1609)) and not (layer1_outputs(365));
    layer2_outputs(1500) <= not(layer1_outputs(1429));
    layer2_outputs(1501) <= (layer1_outputs(2236)) or (layer1_outputs(1001));
    layer2_outputs(1502) <= layer1_outputs(2408);
    layer2_outputs(1503) <= not((layer1_outputs(1161)) xor (layer1_outputs(2532)));
    layer2_outputs(1504) <= layer1_outputs(1004);
    layer2_outputs(1505) <= not(layer1_outputs(2038));
    layer2_outputs(1506) <= (layer1_outputs(999)) or (layer1_outputs(1172));
    layer2_outputs(1507) <= (layer1_outputs(1049)) xor (layer1_outputs(117));
    layer2_outputs(1508) <= (layer1_outputs(850)) and not (layer1_outputs(1936));
    layer2_outputs(1509) <= not((layer1_outputs(230)) or (layer1_outputs(121)));
    layer2_outputs(1510) <= layer1_outputs(709);
    layer2_outputs(1511) <= not(layer1_outputs(1990));
    layer2_outputs(1512) <= not(layer1_outputs(1325)) or (layer1_outputs(1148));
    layer2_outputs(1513) <= layer1_outputs(850);
    layer2_outputs(1514) <= (layer1_outputs(631)) and not (layer1_outputs(983));
    layer2_outputs(1515) <= '1';
    layer2_outputs(1516) <= layer1_outputs(1396);
    layer2_outputs(1517) <= (layer1_outputs(976)) and (layer1_outputs(647));
    layer2_outputs(1518) <= layer1_outputs(207);
    layer2_outputs(1519) <= (layer1_outputs(1568)) and (layer1_outputs(985));
    layer2_outputs(1520) <= not(layer1_outputs(604)) or (layer1_outputs(1341));
    layer2_outputs(1521) <= layer1_outputs(959);
    layer2_outputs(1522) <= not((layer1_outputs(2275)) or (layer1_outputs(1147)));
    layer2_outputs(1523) <= (layer1_outputs(510)) and (layer1_outputs(183));
    layer2_outputs(1524) <= not(layer1_outputs(1979));
    layer2_outputs(1525) <= not(layer1_outputs(851)) or (layer1_outputs(1988));
    layer2_outputs(1526) <= not(layer1_outputs(959));
    layer2_outputs(1527) <= (layer1_outputs(4)) xor (layer1_outputs(919));
    layer2_outputs(1528) <= not((layer1_outputs(922)) or (layer1_outputs(2015)));
    layer2_outputs(1529) <= layer1_outputs(1069);
    layer2_outputs(1530) <= not(layer1_outputs(2297));
    layer2_outputs(1531) <= not(layer1_outputs(1701));
    layer2_outputs(1532) <= not((layer1_outputs(2399)) or (layer1_outputs(1924)));
    layer2_outputs(1533) <= (layer1_outputs(65)) and not (layer1_outputs(1554));
    layer2_outputs(1534) <= (layer1_outputs(439)) or (layer1_outputs(1378));
    layer2_outputs(1535) <= not(layer1_outputs(708));
    layer2_outputs(1536) <= not((layer1_outputs(1469)) and (layer1_outputs(2473)));
    layer2_outputs(1537) <= layer1_outputs(344);
    layer2_outputs(1538) <= (layer1_outputs(1624)) and (layer1_outputs(514));
    layer2_outputs(1539) <= layer1_outputs(1772);
    layer2_outputs(1540) <= (layer1_outputs(1467)) or (layer1_outputs(11));
    layer2_outputs(1541) <= not(layer1_outputs(1511));
    layer2_outputs(1542) <= (layer1_outputs(274)) and not (layer1_outputs(2311));
    layer2_outputs(1543) <= (layer1_outputs(1524)) and (layer1_outputs(1933));
    layer2_outputs(1544) <= (layer1_outputs(64)) and not (layer1_outputs(1689));
    layer2_outputs(1545) <= not(layer1_outputs(85)) or (layer1_outputs(955));
    layer2_outputs(1546) <= not(layer1_outputs(1895)) or (layer1_outputs(434));
    layer2_outputs(1547) <= layer1_outputs(165);
    layer2_outputs(1548) <= not(layer1_outputs(324)) or (layer1_outputs(164));
    layer2_outputs(1549) <= not(layer1_outputs(1644)) or (layer1_outputs(1725));
    layer2_outputs(1550) <= (layer1_outputs(999)) or (layer1_outputs(641));
    layer2_outputs(1551) <= layer1_outputs(35);
    layer2_outputs(1552) <= layer1_outputs(483);
    layer2_outputs(1553) <= not(layer1_outputs(1741));
    layer2_outputs(1554) <= not(layer1_outputs(2023));
    layer2_outputs(1555) <= not(layer1_outputs(1022));
    layer2_outputs(1556) <= (layer1_outputs(2459)) and not (layer1_outputs(1852));
    layer2_outputs(1557) <= not((layer1_outputs(2106)) and (layer1_outputs(698)));
    layer2_outputs(1558) <= not((layer1_outputs(114)) or (layer1_outputs(343)));
    layer2_outputs(1559) <= not(layer1_outputs(2456));
    layer2_outputs(1560) <= not(layer1_outputs(778)) or (layer1_outputs(750));
    layer2_outputs(1561) <= layer1_outputs(1965);
    layer2_outputs(1562) <= not(layer1_outputs(59)) or (layer1_outputs(1771));
    layer2_outputs(1563) <= layer1_outputs(2223);
    layer2_outputs(1564) <= not(layer1_outputs(2229));
    layer2_outputs(1565) <= (layer1_outputs(833)) or (layer1_outputs(1142));
    layer2_outputs(1566) <= not(layer1_outputs(1750));
    layer2_outputs(1567) <= not(layer1_outputs(1956)) or (layer1_outputs(2293));
    layer2_outputs(1568) <= not(layer1_outputs(1670));
    layer2_outputs(1569) <= not(layer1_outputs(1406));
    layer2_outputs(1570) <= layer1_outputs(2385);
    layer2_outputs(1571) <= (layer1_outputs(1224)) and not (layer1_outputs(2388));
    layer2_outputs(1572) <= layer1_outputs(1371);
    layer2_outputs(1573) <= (layer1_outputs(1190)) or (layer1_outputs(1691));
    layer2_outputs(1574) <= (layer1_outputs(1526)) and not (layer1_outputs(293));
    layer2_outputs(1575) <= not(layer1_outputs(1565));
    layer2_outputs(1576) <= not((layer1_outputs(1816)) or (layer1_outputs(498)));
    layer2_outputs(1577) <= (layer1_outputs(131)) and not (layer1_outputs(707));
    layer2_outputs(1578) <= not(layer1_outputs(721));
    layer2_outputs(1579) <= layer1_outputs(1837);
    layer2_outputs(1580) <= not(layer1_outputs(1473));
    layer2_outputs(1581) <= not((layer1_outputs(278)) and (layer1_outputs(2028)));
    layer2_outputs(1582) <= not(layer1_outputs(845)) or (layer1_outputs(1567));
    layer2_outputs(1583) <= (layer1_outputs(700)) and not (layer1_outputs(1555));
    layer2_outputs(1584) <= layer1_outputs(2241);
    layer2_outputs(1585) <= not(layer1_outputs(1134)) or (layer1_outputs(1545));
    layer2_outputs(1586) <= layer1_outputs(991);
    layer2_outputs(1587) <= layer1_outputs(2492);
    layer2_outputs(1588) <= (layer1_outputs(2310)) and not (layer1_outputs(2239));
    layer2_outputs(1589) <= (layer1_outputs(2296)) or (layer1_outputs(2290));
    layer2_outputs(1590) <= (layer1_outputs(1456)) and not (layer1_outputs(1419));
    layer2_outputs(1591) <= not((layer1_outputs(1405)) or (layer1_outputs(1658)));
    layer2_outputs(1592) <= not((layer1_outputs(1854)) and (layer1_outputs(1495)));
    layer2_outputs(1593) <= layer1_outputs(2369);
    layer2_outputs(1594) <= (layer1_outputs(1015)) and not (layer1_outputs(1798));
    layer2_outputs(1595) <= (layer1_outputs(686)) xor (layer1_outputs(2207));
    layer2_outputs(1596) <= not(layer1_outputs(629));
    layer2_outputs(1597) <= not(layer1_outputs(2018));
    layer2_outputs(1598) <= not(layer1_outputs(830)) or (layer1_outputs(1828));
    layer2_outputs(1599) <= not((layer1_outputs(1898)) or (layer1_outputs(658)));
    layer2_outputs(1600) <= not(layer1_outputs(1294)) or (layer1_outputs(295));
    layer2_outputs(1601) <= not(layer1_outputs(1196));
    layer2_outputs(1602) <= layer1_outputs(436);
    layer2_outputs(1603) <= not(layer1_outputs(2080)) or (layer1_outputs(1428));
    layer2_outputs(1604) <= not(layer1_outputs(1740));
    layer2_outputs(1605) <= (layer1_outputs(1500)) or (layer1_outputs(1742));
    layer2_outputs(1606) <= layer1_outputs(967);
    layer2_outputs(1607) <= (layer1_outputs(1916)) and not (layer1_outputs(1438));
    layer2_outputs(1608) <= not((layer1_outputs(1133)) or (layer1_outputs(1776)));
    layer2_outputs(1609) <= not((layer1_outputs(545)) and (layer1_outputs(1501)));
    layer2_outputs(1610) <= layer1_outputs(2502);
    layer2_outputs(1611) <= (layer1_outputs(2162)) and not (layer1_outputs(1167));
    layer2_outputs(1612) <= not(layer1_outputs(1886)) or (layer1_outputs(1754));
    layer2_outputs(1613) <= not((layer1_outputs(2287)) and (layer1_outputs(2105)));
    layer2_outputs(1614) <= layer1_outputs(1672);
    layer2_outputs(1615) <= '0';
    layer2_outputs(1616) <= (layer1_outputs(2451)) and (layer1_outputs(1138));
    layer2_outputs(1617) <= not(layer1_outputs(796));
    layer2_outputs(1618) <= (layer1_outputs(2487)) xor (layer1_outputs(1934));
    layer2_outputs(1619) <= layer1_outputs(188);
    layer2_outputs(1620) <= (layer1_outputs(1838)) or (layer1_outputs(1914));
    layer2_outputs(1621) <= (layer1_outputs(1421)) and (layer1_outputs(1710));
    layer2_outputs(1622) <= not((layer1_outputs(1388)) xor (layer1_outputs(2414)));
    layer2_outputs(1623) <= not((layer1_outputs(1000)) or (layer1_outputs(485)));
    layer2_outputs(1624) <= (layer1_outputs(661)) and not (layer1_outputs(1020));
    layer2_outputs(1625) <= not(layer1_outputs(1504)) or (layer1_outputs(1715));
    layer2_outputs(1626) <= (layer1_outputs(796)) and not (layer1_outputs(1237));
    layer2_outputs(1627) <= layer1_outputs(60);
    layer2_outputs(1628) <= layer1_outputs(1180);
    layer2_outputs(1629) <= not((layer1_outputs(243)) or (layer1_outputs(2330)));
    layer2_outputs(1630) <= layer1_outputs(781);
    layer2_outputs(1631) <= layer1_outputs(2211);
    layer2_outputs(1632) <= (layer1_outputs(282)) and (layer1_outputs(1887));
    layer2_outputs(1633) <= not(layer1_outputs(1329)) or (layer1_outputs(1274));
    layer2_outputs(1634) <= (layer1_outputs(300)) or (layer1_outputs(2110));
    layer2_outputs(1635) <= not((layer1_outputs(2334)) and (layer1_outputs(2093)));
    layer2_outputs(1636) <= not(layer1_outputs(28)) or (layer1_outputs(478));
    layer2_outputs(1637) <= (layer1_outputs(1571)) and not (layer1_outputs(2490));
    layer2_outputs(1638) <= not(layer1_outputs(552));
    layer2_outputs(1639) <= not(layer1_outputs(2058));
    layer2_outputs(1640) <= (layer1_outputs(1150)) and not (layer1_outputs(138));
    layer2_outputs(1641) <= not(layer1_outputs(2173));
    layer2_outputs(1642) <= (layer1_outputs(2122)) and not (layer1_outputs(1133));
    layer2_outputs(1643) <= (layer1_outputs(595)) xor (layer1_outputs(927));
    layer2_outputs(1644) <= not(layer1_outputs(2388)) or (layer1_outputs(387));
    layer2_outputs(1645) <= not(layer1_outputs(1937));
    layer2_outputs(1646) <= not(layer1_outputs(457)) or (layer1_outputs(852));
    layer2_outputs(1647) <= layer1_outputs(432);
    layer2_outputs(1648) <= (layer1_outputs(1359)) and (layer1_outputs(53));
    layer2_outputs(1649) <= layer1_outputs(408);
    layer2_outputs(1650) <= not(layer1_outputs(2323)) or (layer1_outputs(124));
    layer2_outputs(1651) <= not((layer1_outputs(329)) and (layer1_outputs(861)));
    layer2_outputs(1652) <= not(layer1_outputs(1171));
    layer2_outputs(1653) <= not(layer1_outputs(25)) or (layer1_outputs(443));
    layer2_outputs(1654) <= not(layer1_outputs(1472));
    layer2_outputs(1655) <= (layer1_outputs(456)) and not (layer1_outputs(575));
    layer2_outputs(1656) <= layer1_outputs(2460);
    layer2_outputs(1657) <= '0';
    layer2_outputs(1658) <= not(layer1_outputs(2322)) or (layer1_outputs(703));
    layer2_outputs(1659) <= layer1_outputs(1184);
    layer2_outputs(1660) <= (layer1_outputs(333)) and (layer1_outputs(1280));
    layer2_outputs(1661) <= not(layer1_outputs(339)) or (layer1_outputs(2241));
    layer2_outputs(1662) <= not(layer1_outputs(207));
    layer2_outputs(1663) <= (layer1_outputs(1946)) and not (layer1_outputs(2267));
    layer2_outputs(1664) <= (layer1_outputs(1233)) and not (layer1_outputs(374));
    layer2_outputs(1665) <= not(layer1_outputs(2458));
    layer2_outputs(1666) <= not(layer1_outputs(1573));
    layer2_outputs(1667) <= not(layer1_outputs(2360));
    layer2_outputs(1668) <= not((layer1_outputs(238)) and (layer1_outputs(742)));
    layer2_outputs(1669) <= (layer1_outputs(984)) and not (layer1_outputs(1253));
    layer2_outputs(1670) <= (layer1_outputs(1175)) and (layer1_outputs(1246));
    layer2_outputs(1671) <= layer1_outputs(536);
    layer2_outputs(1672) <= not(layer1_outputs(2012));
    layer2_outputs(1673) <= layer1_outputs(1569);
    layer2_outputs(1674) <= not(layer1_outputs(1907));
    layer2_outputs(1675) <= not(layer1_outputs(2326));
    layer2_outputs(1676) <= layer1_outputs(627);
    layer2_outputs(1677) <= (layer1_outputs(973)) or (layer1_outputs(1847));
    layer2_outputs(1678) <= layer1_outputs(478);
    layer2_outputs(1679) <= not((layer1_outputs(321)) and (layer1_outputs(2032)));
    layer2_outputs(1680) <= (layer1_outputs(2310)) and not (layer1_outputs(2345));
    layer2_outputs(1681) <= not(layer1_outputs(110));
    layer2_outputs(1682) <= (layer1_outputs(1483)) and not (layer1_outputs(1994));
    layer2_outputs(1683) <= not(layer1_outputs(1018)) or (layer1_outputs(1199));
    layer2_outputs(1684) <= not(layer1_outputs(714)) or (layer1_outputs(1642));
    layer2_outputs(1685) <= not(layer1_outputs(476)) or (layer1_outputs(272));
    layer2_outputs(1686) <= not(layer1_outputs(52)) or (layer1_outputs(1974));
    layer2_outputs(1687) <= not(layer1_outputs(2067)) or (layer1_outputs(608));
    layer2_outputs(1688) <= not(layer1_outputs(267));
    layer2_outputs(1689) <= layer1_outputs(1711);
    layer2_outputs(1690) <= (layer1_outputs(1322)) and not (layer1_outputs(2021));
    layer2_outputs(1691) <= (layer1_outputs(629)) and not (layer1_outputs(1114));
    layer2_outputs(1692) <= not(layer1_outputs(375));
    layer2_outputs(1693) <= not(layer1_outputs(996)) or (layer1_outputs(1870));
    layer2_outputs(1694) <= not(layer1_outputs(2468));
    layer2_outputs(1695) <= (layer1_outputs(2188)) and (layer1_outputs(2120));
    layer2_outputs(1696) <= layer1_outputs(1312);
    layer2_outputs(1697) <= not(layer1_outputs(156));
    layer2_outputs(1698) <= not(layer1_outputs(1474));
    layer2_outputs(1699) <= (layer1_outputs(2008)) and not (layer1_outputs(306));
    layer2_outputs(1700) <= layer1_outputs(935);
    layer2_outputs(1701) <= (layer1_outputs(517)) and not (layer1_outputs(898));
    layer2_outputs(1702) <= '0';
    layer2_outputs(1703) <= not(layer1_outputs(790));
    layer2_outputs(1704) <= not(layer1_outputs(383)) or (layer1_outputs(774));
    layer2_outputs(1705) <= layer1_outputs(952);
    layer2_outputs(1706) <= not((layer1_outputs(568)) and (layer1_outputs(2125)));
    layer2_outputs(1707) <= not(layer1_outputs(1170));
    layer2_outputs(1708) <= not(layer1_outputs(1137));
    layer2_outputs(1709) <= not(layer1_outputs(2201));
    layer2_outputs(1710) <= layer1_outputs(1706);
    layer2_outputs(1711) <= not(layer1_outputs(1708)) or (layer1_outputs(1331));
    layer2_outputs(1712) <= layer1_outputs(469);
    layer2_outputs(1713) <= not(layer1_outputs(1757));
    layer2_outputs(1714) <= not(layer1_outputs(1572));
    layer2_outputs(1715) <= not(layer1_outputs(2191)) or (layer1_outputs(2348));
    layer2_outputs(1716) <= not((layer1_outputs(298)) or (layer1_outputs(587)));
    layer2_outputs(1717) <= (layer1_outputs(2088)) and not (layer1_outputs(11));
    layer2_outputs(1718) <= not(layer1_outputs(480));
    layer2_outputs(1719) <= not(layer1_outputs(128)) or (layer1_outputs(2427));
    layer2_outputs(1720) <= not(layer1_outputs(602));
    layer2_outputs(1721) <= (layer1_outputs(1297)) and not (layer1_outputs(428));
    layer2_outputs(1722) <= not(layer1_outputs(2483));
    layer2_outputs(1723) <= layer1_outputs(2509);
    layer2_outputs(1724) <= '1';
    layer2_outputs(1725) <= not((layer1_outputs(1038)) and (layer1_outputs(1537)));
    layer2_outputs(1726) <= (layer1_outputs(287)) and not (layer1_outputs(917));
    layer2_outputs(1727) <= not(layer1_outputs(827));
    layer2_outputs(1728) <= (layer1_outputs(1224)) and not (layer1_outputs(168));
    layer2_outputs(1729) <= not(layer1_outputs(1759));
    layer2_outputs(1730) <= layer1_outputs(1972);
    layer2_outputs(1731) <= (layer1_outputs(2240)) and (layer1_outputs(2185));
    layer2_outputs(1732) <= layer1_outputs(338);
    layer2_outputs(1733) <= (layer1_outputs(582)) and not (layer1_outputs(2204));
    layer2_outputs(1734) <= (layer1_outputs(2522)) or (layer1_outputs(2170));
    layer2_outputs(1735) <= layer1_outputs(605);
    layer2_outputs(1736) <= (layer1_outputs(1260)) or (layer1_outputs(966));
    layer2_outputs(1737) <= not(layer1_outputs(121));
    layer2_outputs(1738) <= not(layer1_outputs(571)) or (layer1_outputs(1));
    layer2_outputs(1739) <= (layer1_outputs(1767)) and not (layer1_outputs(705));
    layer2_outputs(1740) <= (layer1_outputs(1367)) or (layer1_outputs(2392));
    layer2_outputs(1741) <= not(layer1_outputs(1143));
    layer2_outputs(1742) <= not(layer1_outputs(1503));
    layer2_outputs(1743) <= not(layer1_outputs(2371));
    layer2_outputs(1744) <= not(layer1_outputs(191)) or (layer1_outputs(661));
    layer2_outputs(1745) <= (layer1_outputs(741)) and not (layer1_outputs(1670));
    layer2_outputs(1746) <= not((layer1_outputs(306)) and (layer1_outputs(1663)));
    layer2_outputs(1747) <= not(layer1_outputs(949)) or (layer1_outputs(2232));
    layer2_outputs(1748) <= not(layer1_outputs(486));
    layer2_outputs(1749) <= not(layer1_outputs(1933));
    layer2_outputs(1750) <= (layer1_outputs(372)) and (layer1_outputs(1218));
    layer2_outputs(1751) <= not(layer1_outputs(2010));
    layer2_outputs(1752) <= not(layer1_outputs(1817));
    layer2_outputs(1753) <= layer1_outputs(690);
    layer2_outputs(1754) <= layer1_outputs(1232);
    layer2_outputs(1755) <= not(layer1_outputs(809));
    layer2_outputs(1756) <= not(layer1_outputs(376)) or (layer1_outputs(19));
    layer2_outputs(1757) <= (layer1_outputs(1071)) and (layer1_outputs(591));
    layer2_outputs(1758) <= not(layer1_outputs(1829));
    layer2_outputs(1759) <= (layer1_outputs(1926)) and (layer1_outputs(2117));
    layer2_outputs(1760) <= (layer1_outputs(2161)) and not (layer1_outputs(857));
    layer2_outputs(1761) <= (layer1_outputs(1633)) and (layer1_outputs(1507));
    layer2_outputs(1762) <= layer1_outputs(2409);
    layer2_outputs(1763) <= not((layer1_outputs(198)) and (layer1_outputs(1716)));
    layer2_outputs(1764) <= not(layer1_outputs(639));
    layer2_outputs(1765) <= not((layer1_outputs(1025)) or (layer1_outputs(155)));
    layer2_outputs(1766) <= not(layer1_outputs(422));
    layer2_outputs(1767) <= '0';
    layer2_outputs(1768) <= layer1_outputs(200);
    layer2_outputs(1769) <= not(layer1_outputs(16)) or (layer1_outputs(1616));
    layer2_outputs(1770) <= (layer1_outputs(1175)) or (layer1_outputs(1267));
    layer2_outputs(1771) <= layer1_outputs(327);
    layer2_outputs(1772) <= not(layer1_outputs(858)) or (layer1_outputs(2132));
    layer2_outputs(1773) <= (layer1_outputs(1705)) and not (layer1_outputs(2380));
    layer2_outputs(1774) <= (layer1_outputs(2518)) and (layer1_outputs(1410));
    layer2_outputs(1775) <= not((layer1_outputs(536)) or (layer1_outputs(1683)));
    layer2_outputs(1776) <= not(layer1_outputs(760));
    layer2_outputs(1777) <= not(layer1_outputs(1825)) or (layer1_outputs(1586));
    layer2_outputs(1778) <= not(layer1_outputs(1334)) or (layer1_outputs(2402));
    layer2_outputs(1779) <= not(layer1_outputs(1117)) or (layer1_outputs(26));
    layer2_outputs(1780) <= not((layer1_outputs(533)) and (layer1_outputs(1766)));
    layer2_outputs(1781) <= not(layer1_outputs(668));
    layer2_outputs(1782) <= layer1_outputs(1464);
    layer2_outputs(1783) <= layer1_outputs(2030);
    layer2_outputs(1784) <= (layer1_outputs(1871)) or (layer1_outputs(1722));
    layer2_outputs(1785) <= layer1_outputs(1659);
    layer2_outputs(1786) <= not(layer1_outputs(968));
    layer2_outputs(1787) <= not((layer1_outputs(2398)) or (layer1_outputs(1245)));
    layer2_outputs(1788) <= (layer1_outputs(2004)) and not (layer1_outputs(2039));
    layer2_outputs(1789) <= not(layer1_outputs(723)) or (layer1_outputs(1075));
    layer2_outputs(1790) <= not(layer1_outputs(1850));
    layer2_outputs(1791) <= (layer1_outputs(17)) or (layer1_outputs(2005));
    layer2_outputs(1792) <= layer1_outputs(1298);
    layer2_outputs(1793) <= (layer1_outputs(1715)) and (layer1_outputs(623));
    layer2_outputs(1794) <= not(layer1_outputs(1967)) or (layer1_outputs(2547));
    layer2_outputs(1795) <= layer1_outputs(2043);
    layer2_outputs(1796) <= (layer1_outputs(57)) or (layer1_outputs(37));
    layer2_outputs(1797) <= layer1_outputs(1779);
    layer2_outputs(1798) <= not((layer1_outputs(693)) xor (layer1_outputs(1368)));
    layer2_outputs(1799) <= not(layer1_outputs(345));
    layer2_outputs(1800) <= layer1_outputs(1654);
    layer2_outputs(1801) <= not(layer1_outputs(1505)) or (layer1_outputs(1731));
    layer2_outputs(1802) <= layer1_outputs(1002);
    layer2_outputs(1803) <= not(layer1_outputs(2081)) or (layer1_outputs(1721));
    layer2_outputs(1804) <= not(layer1_outputs(630));
    layer2_outputs(1805) <= layer1_outputs(1584);
    layer2_outputs(1806) <= not(layer1_outputs(1431));
    layer2_outputs(1807) <= not(layer1_outputs(921)) or (layer1_outputs(606));
    layer2_outputs(1808) <= not(layer1_outputs(1228));
    layer2_outputs(1809) <= not(layer1_outputs(1558));
    layer2_outputs(1810) <= layer1_outputs(1032);
    layer2_outputs(1811) <= (layer1_outputs(869)) xor (layer1_outputs(155));
    layer2_outputs(1812) <= layer1_outputs(305);
    layer2_outputs(1813) <= not((layer1_outputs(1229)) and (layer1_outputs(1212)));
    layer2_outputs(1814) <= (layer1_outputs(261)) and not (layer1_outputs(1998));
    layer2_outputs(1815) <= not(layer1_outputs(961)) or (layer1_outputs(1588));
    layer2_outputs(1816) <= (layer1_outputs(2092)) and not (layer1_outputs(1053));
    layer2_outputs(1817) <= not(layer1_outputs(2008));
    layer2_outputs(1818) <= layer1_outputs(146);
    layer2_outputs(1819) <= not(layer1_outputs(268)) or (layer1_outputs(362));
    layer2_outputs(1820) <= layer1_outputs(2134);
    layer2_outputs(1821) <= (layer1_outputs(745)) or (layer1_outputs(1255));
    layer2_outputs(1822) <= layer1_outputs(1166);
    layer2_outputs(1823) <= (layer1_outputs(344)) and not (layer1_outputs(1713));
    layer2_outputs(1824) <= layer1_outputs(1184);
    layer2_outputs(1825) <= layer1_outputs(2542);
    layer2_outputs(1826) <= not((layer1_outputs(2247)) xor (layer1_outputs(1747)));
    layer2_outputs(1827) <= not(layer1_outputs(713)) or (layer1_outputs(2355));
    layer2_outputs(1828) <= not(layer1_outputs(2219));
    layer2_outputs(1829) <= not(layer1_outputs(2019));
    layer2_outputs(1830) <= not(layer1_outputs(486)) or (layer1_outputs(624));
    layer2_outputs(1831) <= layer1_outputs(2326);
    layer2_outputs(1832) <= not((layer1_outputs(2166)) and (layer1_outputs(2366)));
    layer2_outputs(1833) <= (layer1_outputs(2531)) and not (layer1_outputs(2166));
    layer2_outputs(1834) <= (layer1_outputs(832)) and not (layer1_outputs(1665));
    layer2_outputs(1835) <= not(layer1_outputs(1363)) or (layer1_outputs(1199));
    layer2_outputs(1836) <= not((layer1_outputs(1600)) or (layer1_outputs(2064)));
    layer2_outputs(1837) <= not((layer1_outputs(1531)) xor (layer1_outputs(1334)));
    layer2_outputs(1838) <= not(layer1_outputs(1512)) or (layer1_outputs(1375));
    layer2_outputs(1839) <= not(layer1_outputs(1862)) or (layer1_outputs(2014));
    layer2_outputs(1840) <= not(layer1_outputs(2156)) or (layer1_outputs(348));
    layer2_outputs(1841) <= (layer1_outputs(904)) or (layer1_outputs(1090));
    layer2_outputs(1842) <= (layer1_outputs(1337)) and not (layer1_outputs(1696));
    layer2_outputs(1843) <= layer1_outputs(844);
    layer2_outputs(1844) <= '0';
    layer2_outputs(1845) <= not(layer1_outputs(1286)) or (layer1_outputs(1330));
    layer2_outputs(1846) <= layer1_outputs(769);
    layer2_outputs(1847) <= (layer1_outputs(1047)) and not (layer1_outputs(1160));
    layer2_outputs(1848) <= not((layer1_outputs(1911)) and (layer1_outputs(930)));
    layer2_outputs(1849) <= not(layer1_outputs(492)) or (layer1_outputs(1471));
    layer2_outputs(1850) <= not(layer1_outputs(30));
    layer2_outputs(1851) <= not(layer1_outputs(993)) or (layer1_outputs(150));
    layer2_outputs(1852) <= layer1_outputs(1461);
    layer2_outputs(1853) <= not(layer1_outputs(2464));
    layer2_outputs(1854) <= not(layer1_outputs(2188));
    layer2_outputs(1855) <= not(layer1_outputs(2383));
    layer2_outputs(1856) <= not(layer1_outputs(1574));
    layer2_outputs(1857) <= (layer1_outputs(2096)) and not (layer1_outputs(1948));
    layer2_outputs(1858) <= not(layer1_outputs(2205));
    layer2_outputs(1859) <= layer1_outputs(547);
    layer2_outputs(1860) <= (layer1_outputs(2378)) and not (layer1_outputs(953));
    layer2_outputs(1861) <= layer1_outputs(455);
    layer2_outputs(1862) <= '1';
    layer2_outputs(1863) <= not(layer1_outputs(1461)) or (layer1_outputs(2209));
    layer2_outputs(1864) <= layer1_outputs(1513);
    layer2_outputs(1865) <= layer1_outputs(732);
    layer2_outputs(1866) <= layer1_outputs(632);
    layer2_outputs(1867) <= layer1_outputs(2423);
    layer2_outputs(1868) <= not(layer1_outputs(41));
    layer2_outputs(1869) <= not((layer1_outputs(973)) or (layer1_outputs(561)));
    layer2_outputs(1870) <= not(layer1_outputs(1265)) or (layer1_outputs(1475));
    layer2_outputs(1871) <= not((layer1_outputs(1925)) xor (layer1_outputs(1244)));
    layer2_outputs(1872) <= not(layer1_outputs(1517));
    layer2_outputs(1873) <= (layer1_outputs(2459)) and not (layer1_outputs(1570));
    layer2_outputs(1874) <= (layer1_outputs(36)) and not (layer1_outputs(1753));
    layer2_outputs(1875) <= '0';
    layer2_outputs(1876) <= (layer1_outputs(2556)) and not (layer1_outputs(1607));
    layer2_outputs(1877) <= not(layer1_outputs(1547));
    layer2_outputs(1878) <= not(layer1_outputs(1665)) or (layer1_outputs(1693));
    layer2_outputs(1879) <= not((layer1_outputs(2114)) and (layer1_outputs(1246)));
    layer2_outputs(1880) <= (layer1_outputs(1136)) and not (layer1_outputs(1361));
    layer2_outputs(1881) <= not(layer1_outputs(570));
    layer2_outputs(1882) <= layer1_outputs(697);
    layer2_outputs(1883) <= not((layer1_outputs(1348)) and (layer1_outputs(162)));
    layer2_outputs(1884) <= (layer1_outputs(2221)) and not (layer1_outputs(549));
    layer2_outputs(1885) <= not(layer1_outputs(1097));
    layer2_outputs(1886) <= not(layer1_outputs(383));
    layer2_outputs(1887) <= layer1_outputs(990);
    layer2_outputs(1888) <= (layer1_outputs(1045)) or (layer1_outputs(447));
    layer2_outputs(1889) <= not(layer1_outputs(1739));
    layer2_outputs(1890) <= (layer1_outputs(1622)) and not (layer1_outputs(2224));
    layer2_outputs(1891) <= layer1_outputs(1367);
    layer2_outputs(1892) <= not(layer1_outputs(1087));
    layer2_outputs(1893) <= not(layer1_outputs(2043));
    layer2_outputs(1894) <= layer1_outputs(79);
    layer2_outputs(1895) <= not(layer1_outputs(1209));
    layer2_outputs(1896) <= not(layer1_outputs(2498));
    layer2_outputs(1897) <= '0';
    layer2_outputs(1898) <= (layer1_outputs(1778)) or (layer1_outputs(15));
    layer2_outputs(1899) <= not(layer1_outputs(1079));
    layer2_outputs(1900) <= not(layer1_outputs(722));
    layer2_outputs(1901) <= not((layer1_outputs(1290)) and (layer1_outputs(459)));
    layer2_outputs(1902) <= layer1_outputs(1951);
    layer2_outputs(1903) <= not(layer1_outputs(1608)) or (layer1_outputs(221));
    layer2_outputs(1904) <= layer1_outputs(1807);
    layer2_outputs(1905) <= not((layer1_outputs(1591)) or (layer1_outputs(1484)));
    layer2_outputs(1906) <= not(layer1_outputs(1696));
    layer2_outputs(1907) <= not((layer1_outputs(2237)) or (layer1_outputs(2113)));
    layer2_outputs(1908) <= not(layer1_outputs(2111));
    layer2_outputs(1909) <= not((layer1_outputs(1309)) or (layer1_outputs(1355)));
    layer2_outputs(1910) <= not(layer1_outputs(1183));
    layer2_outputs(1911) <= (layer1_outputs(1611)) or (layer1_outputs(2444));
    layer2_outputs(1912) <= (layer1_outputs(615)) and not (layer1_outputs(2361));
    layer2_outputs(1913) <= (layer1_outputs(410)) or (layer1_outputs(2533));
    layer2_outputs(1914) <= not(layer1_outputs(1443));
    layer2_outputs(1915) <= layer1_outputs(350);
    layer2_outputs(1916) <= not(layer1_outputs(421));
    layer2_outputs(1917) <= not((layer1_outputs(12)) or (layer1_outputs(682)));
    layer2_outputs(1918) <= not((layer1_outputs(747)) xor (layer1_outputs(2553)));
    layer2_outputs(1919) <= layer1_outputs(1620);
    layer2_outputs(1920) <= (layer1_outputs(2490)) and not (layer1_outputs(848));
    layer2_outputs(1921) <= not((layer1_outputs(1527)) xor (layer1_outputs(249)));
    layer2_outputs(1922) <= layer1_outputs(1480);
    layer2_outputs(1923) <= not(layer1_outputs(1250));
    layer2_outputs(1924) <= layer1_outputs(1791);
    layer2_outputs(1925) <= layer1_outputs(1985);
    layer2_outputs(1926) <= '1';
    layer2_outputs(1927) <= layer1_outputs(1327);
    layer2_outputs(1928) <= layer1_outputs(141);
    layer2_outputs(1929) <= (layer1_outputs(1984)) and not (layer1_outputs(1182));
    layer2_outputs(1930) <= (layer1_outputs(2252)) and (layer1_outputs(2488));
    layer2_outputs(1931) <= layer1_outputs(2517);
    layer2_outputs(1932) <= (layer1_outputs(2519)) and (layer1_outputs(2110));
    layer2_outputs(1933) <= layer1_outputs(2002);
    layer2_outputs(1934) <= not(layer1_outputs(1217));
    layer2_outputs(1935) <= not(layer1_outputs(1680));
    layer2_outputs(1936) <= (layer1_outputs(2072)) and not (layer1_outputs(2037));
    layer2_outputs(1937) <= layer1_outputs(2034);
    layer2_outputs(1938) <= (layer1_outputs(607)) and not (layer1_outputs(2325));
    layer2_outputs(1939) <= layer1_outputs(2323);
    layer2_outputs(1940) <= not((layer1_outputs(565)) or (layer1_outputs(1803)));
    layer2_outputs(1941) <= layer1_outputs(948);
    layer2_outputs(1942) <= not(layer1_outputs(319));
    layer2_outputs(1943) <= not(layer1_outputs(384)) or (layer1_outputs(2429));
    layer2_outputs(1944) <= layer1_outputs(1309);
    layer2_outputs(1945) <= not(layer1_outputs(463));
    layer2_outputs(1946) <= layer1_outputs(160);
    layer2_outputs(1947) <= (layer1_outputs(112)) and not (layer1_outputs(564));
    layer2_outputs(1948) <= not(layer1_outputs(218));
    layer2_outputs(1949) <= not(layer1_outputs(2520));
    layer2_outputs(1950) <= layer1_outputs(608);
    layer2_outputs(1951) <= (layer1_outputs(1395)) or (layer1_outputs(1564));
    layer2_outputs(1952) <= not(layer1_outputs(2354)) or (layer1_outputs(1380));
    layer2_outputs(1953) <= (layer1_outputs(934)) and not (layer1_outputs(400));
    layer2_outputs(1954) <= not(layer1_outputs(726));
    layer2_outputs(1955) <= not(layer1_outputs(2480));
    layer2_outputs(1956) <= not(layer1_outputs(1895)) or (layer1_outputs(665));
    layer2_outputs(1957) <= not(layer1_outputs(2449));
    layer2_outputs(1958) <= (layer1_outputs(1414)) or (layer1_outputs(563));
    layer2_outputs(1959) <= not(layer1_outputs(1003));
    layer2_outputs(1960) <= not(layer1_outputs(2049));
    layer2_outputs(1961) <= not(layer1_outputs(878));
    layer2_outputs(1962) <= not(layer1_outputs(1328));
    layer2_outputs(1963) <= (layer1_outputs(1198)) and (layer1_outputs(2027));
    layer2_outputs(1964) <= '0';
    layer2_outputs(1965) <= not((layer1_outputs(1869)) and (layer1_outputs(280)));
    layer2_outputs(1966) <= not(layer1_outputs(960));
    layer2_outputs(1967) <= not((layer1_outputs(135)) or (layer1_outputs(1689)));
    layer2_outputs(1968) <= not(layer1_outputs(1708));
    layer2_outputs(1969) <= not(layer1_outputs(1627));
    layer2_outputs(1970) <= layer1_outputs(110);
    layer2_outputs(1971) <= not(layer1_outputs(2187));
    layer2_outputs(1972) <= not((layer1_outputs(590)) and (layer1_outputs(1346)));
    layer2_outputs(1973) <= not(layer1_outputs(1623));
    layer2_outputs(1974) <= (layer1_outputs(896)) or (layer1_outputs(2046));
    layer2_outputs(1975) <= not(layer1_outputs(2182));
    layer2_outputs(1976) <= layer1_outputs(919);
    layer2_outputs(1977) <= (layer1_outputs(1303)) and not (layer1_outputs(753));
    layer2_outputs(1978) <= (layer1_outputs(1300)) and (layer1_outputs(103));
    layer2_outputs(1979) <= not(layer1_outputs(794));
    layer2_outputs(1980) <= layer1_outputs(481);
    layer2_outputs(1981) <= not((layer1_outputs(704)) or (layer1_outputs(1041)));
    layer2_outputs(1982) <= layer1_outputs(1890);
    layer2_outputs(1983) <= not(layer1_outputs(218)) or (layer1_outputs(2148));
    layer2_outputs(1984) <= (layer1_outputs(1589)) or (layer1_outputs(1700));
    layer2_outputs(1985) <= (layer1_outputs(1769)) and not (layer1_outputs(1401));
    layer2_outputs(1986) <= (layer1_outputs(869)) and (layer1_outputs(1638));
    layer2_outputs(1987) <= not(layer1_outputs(1480));
    layer2_outputs(1988) <= not(layer1_outputs(563));
    layer2_outputs(1989) <= not(layer1_outputs(2023));
    layer2_outputs(1990) <= not((layer1_outputs(974)) and (layer1_outputs(688)));
    layer2_outputs(1991) <= (layer1_outputs(2424)) and not (layer1_outputs(1705));
    layer2_outputs(1992) <= layer1_outputs(2408);
    layer2_outputs(1993) <= layer1_outputs(471);
    layer2_outputs(1994) <= layer1_outputs(2086);
    layer2_outputs(1995) <= (layer1_outputs(822)) and (layer1_outputs(1081));
    layer2_outputs(1996) <= not(layer1_outputs(1010));
    layer2_outputs(1997) <= (layer1_outputs(2423)) or (layer1_outputs(1104));
    layer2_outputs(1998) <= not(layer1_outputs(988)) or (layer1_outputs(898));
    layer2_outputs(1999) <= (layer1_outputs(1719)) and not (layer1_outputs(216));
    layer2_outputs(2000) <= not((layer1_outputs(1200)) or (layer1_outputs(2092)));
    layer2_outputs(2001) <= layer1_outputs(1707);
    layer2_outputs(2002) <= '0';
    layer2_outputs(2003) <= (layer1_outputs(431)) and not (layer1_outputs(2161));
    layer2_outputs(2004) <= not(layer1_outputs(1434));
    layer2_outputs(2005) <= not(layer1_outputs(351));
    layer2_outputs(2006) <= layer1_outputs(2016);
    layer2_outputs(2007) <= not(layer1_outputs(1634));
    layer2_outputs(2008) <= (layer1_outputs(1514)) xor (layer1_outputs(1546));
    layer2_outputs(2009) <= (layer1_outputs(2455)) or (layer1_outputs(530));
    layer2_outputs(2010) <= not(layer1_outputs(1619));
    layer2_outputs(2011) <= (layer1_outputs(729)) and not (layer1_outputs(1797));
    layer2_outputs(2012) <= not(layer1_outputs(1384));
    layer2_outputs(2013) <= not(layer1_outputs(125));
    layer2_outputs(2014) <= not(layer1_outputs(1318));
    layer2_outputs(2015) <= not(layer1_outputs(1089));
    layer2_outputs(2016) <= not(layer1_outputs(2306)) or (layer1_outputs(429));
    layer2_outputs(2017) <= (layer1_outputs(1991)) and (layer1_outputs(55));
    layer2_outputs(2018) <= (layer1_outputs(52)) and not (layer1_outputs(1672));
    layer2_outputs(2019) <= not(layer1_outputs(1804)) or (layer1_outputs(171));
    layer2_outputs(2020) <= not((layer1_outputs(480)) and (layer1_outputs(2186)));
    layer2_outputs(2021) <= not(layer1_outputs(2123));
    layer2_outputs(2022) <= not(layer1_outputs(1343));
    layer2_outputs(2023) <= (layer1_outputs(1834)) or (layer1_outputs(1961));
    layer2_outputs(2024) <= not(layer1_outputs(2352));
    layer2_outputs(2025) <= not(layer1_outputs(261));
    layer2_outputs(2026) <= not((layer1_outputs(1984)) or (layer1_outputs(131)));
    layer2_outputs(2027) <= layer1_outputs(341);
    layer2_outputs(2028) <= not(layer1_outputs(1299));
    layer2_outputs(2029) <= not(layer1_outputs(175)) or (layer1_outputs(540));
    layer2_outputs(2030) <= (layer1_outputs(878)) and not (layer1_outputs(391));
    layer2_outputs(2031) <= layer1_outputs(923);
    layer2_outputs(2032) <= (layer1_outputs(1928)) or (layer1_outputs(1725));
    layer2_outputs(2033) <= not(layer1_outputs(2225));
    layer2_outputs(2034) <= not(layer1_outputs(660));
    layer2_outputs(2035) <= layer1_outputs(2375);
    layer2_outputs(2036) <= not((layer1_outputs(154)) or (layer1_outputs(2253)));
    layer2_outputs(2037) <= not(layer1_outputs(1866));
    layer2_outputs(2038) <= layer1_outputs(1279);
    layer2_outputs(2039) <= layer1_outputs(1603);
    layer2_outputs(2040) <= layer1_outputs(342);
    layer2_outputs(2041) <= not(layer1_outputs(585));
    layer2_outputs(2042) <= not(layer1_outputs(1318));
    layer2_outputs(2043) <= not((layer1_outputs(2394)) or (layer1_outputs(1452)));
    layer2_outputs(2044) <= (layer1_outputs(1910)) and not (layer1_outputs(1063));
    layer2_outputs(2045) <= layer1_outputs(33);
    layer2_outputs(2046) <= not(layer1_outputs(1294)) or (layer1_outputs(1394));
    layer2_outputs(2047) <= (layer1_outputs(700)) xor (layer1_outputs(868));
    layer2_outputs(2048) <= (layer1_outputs(1516)) or (layer1_outputs(2074));
    layer2_outputs(2049) <= not(layer1_outputs(1953));
    layer2_outputs(2050) <= not(layer1_outputs(220));
    layer2_outputs(2051) <= layer1_outputs(2308);
    layer2_outputs(2052) <= (layer1_outputs(166)) and (layer1_outputs(856));
    layer2_outputs(2053) <= layer1_outputs(1351);
    layer2_outputs(2054) <= not(layer1_outputs(1411)) or (layer1_outputs(1223));
    layer2_outputs(2055) <= (layer1_outputs(1170)) and (layer1_outputs(2546));
    layer2_outputs(2056) <= (layer1_outputs(864)) and not (layer1_outputs(1723));
    layer2_outputs(2057) <= (layer1_outputs(1633)) and (layer1_outputs(2426));
    layer2_outputs(2058) <= (layer1_outputs(2217)) or (layer1_outputs(913));
    layer2_outputs(2059) <= layer1_outputs(283);
    layer2_outputs(2060) <= not((layer1_outputs(1456)) and (layer1_outputs(774)));
    layer2_outputs(2061) <= layer1_outputs(1359);
    layer2_outputs(2062) <= not((layer1_outputs(994)) or (layer1_outputs(569)));
    layer2_outputs(2063) <= not(layer1_outputs(2301));
    layer2_outputs(2064) <= layer1_outputs(2173);
    layer2_outputs(2065) <= layer1_outputs(1286);
    layer2_outputs(2066) <= (layer1_outputs(174)) and not (layer1_outputs(2314));
    layer2_outputs(2067) <= (layer1_outputs(683)) or (layer1_outputs(1055));
    layer2_outputs(2068) <= not(layer1_outputs(379)) or (layer1_outputs(1583));
    layer2_outputs(2069) <= layer1_outputs(1905);
    layer2_outputs(2070) <= (layer1_outputs(2496)) and not (layer1_outputs(1113));
    layer2_outputs(2071) <= layer1_outputs(320);
    layer2_outputs(2072) <= not(layer1_outputs(1950));
    layer2_outputs(2073) <= not(layer1_outputs(2266)) or (layer1_outputs(2244));
    layer2_outputs(2074) <= not(layer1_outputs(499));
    layer2_outputs(2075) <= layer1_outputs(2412);
    layer2_outputs(2076) <= not(layer1_outputs(1043));
    layer2_outputs(2077) <= not((layer1_outputs(946)) or (layer1_outputs(251)));
    layer2_outputs(2078) <= not((layer1_outputs(1186)) or (layer1_outputs(1865)));
    layer2_outputs(2079) <= not((layer1_outputs(686)) or (layer1_outputs(2417)));
    layer2_outputs(2080) <= not(layer1_outputs(537)) or (layer1_outputs(2338));
    layer2_outputs(2081) <= (layer1_outputs(295)) and not (layer1_outputs(2147));
    layer2_outputs(2082) <= (layer1_outputs(356)) or (layer1_outputs(22));
    layer2_outputs(2083) <= (layer1_outputs(263)) and not (layer1_outputs(1987));
    layer2_outputs(2084) <= not(layer1_outputs(209));
    layer2_outputs(2085) <= (layer1_outputs(559)) and (layer1_outputs(1987));
    layer2_outputs(2086) <= not((layer1_outputs(743)) and (layer1_outputs(524)));
    layer2_outputs(2087) <= not(layer1_outputs(1447));
    layer2_outputs(2088) <= not(layer1_outputs(1258));
    layer2_outputs(2089) <= not((layer1_outputs(1198)) and (layer1_outputs(2444)));
    layer2_outputs(2090) <= not(layer1_outputs(183));
    layer2_outputs(2091) <= not(layer1_outputs(35)) or (layer1_outputs(1443));
    layer2_outputs(2092) <= not(layer1_outputs(1132));
    layer2_outputs(2093) <= not(layer1_outputs(241)) or (layer1_outputs(8));
    layer2_outputs(2094) <= not(layer1_outputs(962));
    layer2_outputs(2095) <= layer1_outputs(445);
    layer2_outputs(2096) <= (layer1_outputs(1894)) and not (layer1_outputs(418));
    layer2_outputs(2097) <= not(layer1_outputs(1332)) or (layer1_outputs(244));
    layer2_outputs(2098) <= not((layer1_outputs(653)) and (layer1_outputs(1861)));
    layer2_outputs(2099) <= not((layer1_outputs(359)) xor (layer1_outputs(1861)));
    layer2_outputs(2100) <= not(layer1_outputs(690)) or (layer1_outputs(1211));
    layer2_outputs(2101) <= layer1_outputs(1209);
    layer2_outputs(2102) <= (layer1_outputs(271)) and (layer1_outputs(2365));
    layer2_outputs(2103) <= layer1_outputs(2335);
    layer2_outputs(2104) <= not(layer1_outputs(2035));
    layer2_outputs(2105) <= not(layer1_outputs(2122)) or (layer1_outputs(1542));
    layer2_outputs(2106) <= not(layer1_outputs(2)) or (layer1_outputs(1449));
    layer2_outputs(2107) <= not((layer1_outputs(688)) and (layer1_outputs(757)));
    layer2_outputs(2108) <= not(layer1_outputs(418));
    layer2_outputs(2109) <= layer1_outputs(1030);
    layer2_outputs(2110) <= (layer1_outputs(39)) and not (layer1_outputs(1666));
    layer2_outputs(2111) <= not(layer1_outputs(147));
    layer2_outputs(2112) <= layer1_outputs(635);
    layer2_outputs(2113) <= (layer1_outputs(2450)) and (layer1_outputs(1384));
    layer2_outputs(2114) <= not(layer1_outputs(2425));
    layer2_outputs(2115) <= not((layer1_outputs(1247)) and (layer1_outputs(1494)));
    layer2_outputs(2116) <= (layer1_outputs(824)) and (layer1_outputs(437));
    layer2_outputs(2117) <= not((layer1_outputs(142)) or (layer1_outputs(176)));
    layer2_outputs(2118) <= not((layer1_outputs(906)) or (layer1_outputs(531)));
    layer2_outputs(2119) <= not(layer1_outputs(2482));
    layer2_outputs(2120) <= (layer1_outputs(914)) and not (layer1_outputs(2313));
    layer2_outputs(2121) <= layer1_outputs(879);
    layer2_outputs(2122) <= (layer1_outputs(106)) or (layer1_outputs(1172));
    layer2_outputs(2123) <= not((layer1_outputs(1578)) or (layer1_outputs(1274)));
    layer2_outputs(2124) <= layer1_outputs(1629);
    layer2_outputs(2125) <= not(layer1_outputs(70)) or (layer1_outputs(2496));
    layer2_outputs(2126) <= (layer1_outputs(2539)) and (layer1_outputs(1778));
    layer2_outputs(2127) <= layer1_outputs(1481);
    layer2_outputs(2128) <= '0';
    layer2_outputs(2129) <= layer1_outputs(641);
    layer2_outputs(2130) <= not((layer1_outputs(1191)) xor (layer1_outputs(352)));
    layer2_outputs(2131) <= not((layer1_outputs(1034)) and (layer1_outputs(2491)));
    layer2_outputs(2132) <= layer1_outputs(2452);
    layer2_outputs(2133) <= (layer1_outputs(711)) and not (layer1_outputs(1779));
    layer2_outputs(2134) <= (layer1_outputs(2254)) and (layer1_outputs(91));
    layer2_outputs(2135) <= not((layer1_outputs(1007)) xor (layer1_outputs(38)));
    layer2_outputs(2136) <= not((layer1_outputs(1156)) xor (layer1_outputs(2189)));
    layer2_outputs(2137) <= not(layer1_outputs(2193));
    layer2_outputs(2138) <= not(layer1_outputs(1376)) or (layer1_outputs(2341));
    layer2_outputs(2139) <= not((layer1_outputs(856)) xor (layer1_outputs(567)));
    layer2_outputs(2140) <= layer1_outputs(50);
    layer2_outputs(2141) <= not((layer1_outputs(1405)) and (layer1_outputs(739)));
    layer2_outputs(2142) <= not(layer1_outputs(1021)) or (layer1_outputs(1566));
    layer2_outputs(2143) <= layer1_outputs(825);
    layer2_outputs(2144) <= (layer1_outputs(365)) or (layer1_outputs(2193));
    layer2_outputs(2145) <= not((layer1_outputs(1254)) and (layer1_outputs(1229)));
    layer2_outputs(2146) <= layer1_outputs(115);
    layer2_outputs(2147) <= not(layer1_outputs(1960));
    layer2_outputs(2148) <= (layer1_outputs(1635)) and not (layer1_outputs(1578));
    layer2_outputs(2149) <= not((layer1_outputs(1552)) or (layer1_outputs(1574)));
    layer2_outputs(2150) <= not((layer1_outputs(389)) or (layer1_outputs(242)));
    layer2_outputs(2151) <= not((layer1_outputs(2395)) or (layer1_outputs(654)));
    layer2_outputs(2152) <= (layer1_outputs(958)) or (layer1_outputs(2527));
    layer2_outputs(2153) <= not(layer1_outputs(2035));
    layer2_outputs(2154) <= (layer1_outputs(1411)) or (layer1_outputs(1475));
    layer2_outputs(2155) <= layer1_outputs(1940);
    layer2_outputs(2156) <= layer1_outputs(2293);
    layer2_outputs(2157) <= (layer1_outputs(2534)) and (layer1_outputs(1570));
    layer2_outputs(2158) <= not(layer1_outputs(2342));
    layer2_outputs(2159) <= (layer1_outputs(1906)) and (layer1_outputs(1403));
    layer2_outputs(2160) <= not(layer1_outputs(1211));
    layer2_outputs(2161) <= layer1_outputs(2551);
    layer2_outputs(2162) <= not(layer1_outputs(286));
    layer2_outputs(2163) <= not(layer1_outputs(1494)) or (layer1_outputs(1831));
    layer2_outputs(2164) <= layer1_outputs(1116);
    layer2_outputs(2165) <= not(layer1_outputs(1237));
    layer2_outputs(2166) <= not(layer1_outputs(1610)) or (layer1_outputs(2250));
    layer2_outputs(2167) <= '0';
    layer2_outputs(2168) <= not(layer1_outputs(2277)) or (layer1_outputs(604));
    layer2_outputs(2169) <= (layer1_outputs(1995)) and (layer1_outputs(1958));
    layer2_outputs(2170) <= not(layer1_outputs(719));
    layer2_outputs(2171) <= not((layer1_outputs(1470)) and (layer1_outputs(789)));
    layer2_outputs(2172) <= layer1_outputs(1993);
    layer2_outputs(2173) <= (layer1_outputs(1643)) or (layer1_outputs(1550));
    layer2_outputs(2174) <= not((layer1_outputs(2438)) and (layer1_outputs(468)));
    layer2_outputs(2175) <= (layer1_outputs(2300)) and not (layer1_outputs(2054));
    layer2_outputs(2176) <= not(layer1_outputs(833));
    layer2_outputs(2177) <= (layer1_outputs(146)) xor (layer1_outputs(1512));
    layer2_outputs(2178) <= (layer1_outputs(1732)) and not (layer1_outputs(1141));
    layer2_outputs(2179) <= not(layer1_outputs(334));
    layer2_outputs(2180) <= (layer1_outputs(2477)) and (layer1_outputs(177));
    layer2_outputs(2181) <= not(layer1_outputs(1888)) or (layer1_outputs(163));
    layer2_outputs(2182) <= not(layer1_outputs(816)) or (layer1_outputs(1971));
    layer2_outputs(2183) <= layer1_outputs(634);
    layer2_outputs(2184) <= not(layer1_outputs(472)) or (layer1_outputs(228));
    layer2_outputs(2185) <= not(layer1_outputs(1013)) or (layer1_outputs(2177));
    layer2_outputs(2186) <= (layer1_outputs(1125)) and not (layer1_outputs(784));
    layer2_outputs(2187) <= '0';
    layer2_outputs(2188) <= not(layer1_outputs(440));
    layer2_outputs(2189) <= layer1_outputs(1099);
    layer2_outputs(2190) <= layer1_outputs(2348);
    layer2_outputs(2191) <= (layer1_outputs(760)) and not (layer1_outputs(1699));
    layer2_outputs(2192) <= '1';
    layer2_outputs(2193) <= not(layer1_outputs(710));
    layer2_outputs(2194) <= (layer1_outputs(2465)) and not (layer1_outputs(2010));
    layer2_outputs(2195) <= (layer1_outputs(84)) xor (layer1_outputs(1611));
    layer2_outputs(2196) <= not(layer1_outputs(1662));
    layer2_outputs(2197) <= layer1_outputs(1285);
    layer2_outputs(2198) <= not(layer1_outputs(1969));
    layer2_outputs(2199) <= not(layer1_outputs(744)) or (layer1_outputs(1692));
    layer2_outputs(2200) <= '0';
    layer2_outputs(2201) <= not((layer1_outputs(1037)) xor (layer1_outputs(2177)));
    layer2_outputs(2202) <= not((layer1_outputs(974)) and (layer1_outputs(911)));
    layer2_outputs(2203) <= layer1_outputs(2135);
    layer2_outputs(2204) <= not(layer1_outputs(358));
    layer2_outputs(2205) <= (layer1_outputs(718)) and not (layer1_outputs(363));
    layer2_outputs(2206) <= not(layer1_outputs(266));
    layer2_outputs(2207) <= not(layer1_outputs(3));
    layer2_outputs(2208) <= layer1_outputs(14);
    layer2_outputs(2209) <= not((layer1_outputs(662)) or (layer1_outputs(614)));
    layer2_outputs(2210) <= not((layer1_outputs(2136)) and (layer1_outputs(2385)));
    layer2_outputs(2211) <= (layer1_outputs(1926)) and not (layer1_outputs(1972));
    layer2_outputs(2212) <= layer1_outputs(1603);
    layer2_outputs(2213) <= not(layer1_outputs(699));
    layer2_outputs(2214) <= layer1_outputs(939);
    layer2_outputs(2215) <= layer1_outputs(1540);
    layer2_outputs(2216) <= (layer1_outputs(2508)) and not (layer1_outputs(1118));
    layer2_outputs(2217) <= (layer1_outputs(1490)) and not (layer1_outputs(2083));
    layer2_outputs(2218) <= '0';
    layer2_outputs(2219) <= not(layer1_outputs(537)) or (layer1_outputs(2048));
    layer2_outputs(2220) <= not((layer1_outputs(2014)) or (layer1_outputs(1585)));
    layer2_outputs(2221) <= not((layer1_outputs(768)) and (layer1_outputs(1832)));
    layer2_outputs(2222) <= layer1_outputs(2251);
    layer2_outputs(2223) <= not((layer1_outputs(775)) and (layer1_outputs(1914)));
    layer2_outputs(2224) <= (layer1_outputs(2538)) or (layer1_outputs(1646));
    layer2_outputs(2225) <= layer1_outputs(2100);
    layer2_outputs(2226) <= layer1_outputs(1121);
    layer2_outputs(2227) <= not((layer1_outputs(1272)) and (layer1_outputs(955)));
    layer2_outputs(2228) <= layer1_outputs(961);
    layer2_outputs(2229) <= layer1_outputs(2487);
    layer2_outputs(2230) <= layer1_outputs(2085);
    layer2_outputs(2231) <= (layer1_outputs(2472)) or (layer1_outputs(333));
    layer2_outputs(2232) <= layer1_outputs(1347);
    layer2_outputs(2233) <= not(layer1_outputs(714));
    layer2_outputs(2234) <= (layer1_outputs(2197)) and not (layer1_outputs(157));
    layer2_outputs(2235) <= layer1_outputs(2332);
    layer2_outputs(2236) <= layer1_outputs(2249);
    layer2_outputs(2237) <= (layer1_outputs(1617)) and (layer1_outputs(1821));
    layer2_outputs(2238) <= not(layer1_outputs(1200));
    layer2_outputs(2239) <= layer1_outputs(9);
    layer2_outputs(2240) <= not(layer1_outputs(2133)) or (layer1_outputs(409));
    layer2_outputs(2241) <= not((layer1_outputs(1927)) or (layer1_outputs(1415)));
    layer2_outputs(2242) <= not(layer1_outputs(2104));
    layer2_outputs(2243) <= not(layer1_outputs(466));
    layer2_outputs(2244) <= layer1_outputs(1220);
    layer2_outputs(2245) <= not(layer1_outputs(696));
    layer2_outputs(2246) <= not(layer1_outputs(1701));
    layer2_outputs(2247) <= (layer1_outputs(932)) or (layer1_outputs(1189));
    layer2_outputs(2248) <= layer1_outputs(496);
    layer2_outputs(2249) <= '1';
    layer2_outputs(2250) <= layer1_outputs(318);
    layer2_outputs(2251) <= (layer1_outputs(782)) and (layer1_outputs(560));
    layer2_outputs(2252) <= not(layer1_outputs(118));
    layer2_outputs(2253) <= not((layer1_outputs(759)) and (layer1_outputs(1726)));
    layer2_outputs(2254) <= not((layer1_outputs(148)) and (layer1_outputs(2019)));
    layer2_outputs(2255) <= not(layer1_outputs(2213)) or (layer1_outputs(987));
    layer2_outputs(2256) <= not(layer1_outputs(1015));
    layer2_outputs(2257) <= layer1_outputs(203);
    layer2_outputs(2258) <= not(layer1_outputs(474));
    layer2_outputs(2259) <= not(layer1_outputs(2358));
    layer2_outputs(2260) <= not(layer1_outputs(76)) or (layer1_outputs(2454));
    layer2_outputs(2261) <= layer1_outputs(1553);
    layer2_outputs(2262) <= not(layer1_outputs(1077));
    layer2_outputs(2263) <= (layer1_outputs(894)) and not (layer1_outputs(428));
    layer2_outputs(2264) <= (layer1_outputs(454)) and (layer1_outputs(1350));
    layer2_outputs(2265) <= layer1_outputs(1124);
    layer2_outputs(2266) <= layer1_outputs(1847);
    layer2_outputs(2267) <= (layer1_outputs(551)) and not (layer1_outputs(1062));
    layer2_outputs(2268) <= not(layer1_outputs(136)) or (layer1_outputs(2374));
    layer2_outputs(2269) <= not(layer1_outputs(2404)) or (layer1_outputs(188));
    layer2_outputs(2270) <= (layer1_outputs(989)) and (layer1_outputs(2401));
    layer2_outputs(2271) <= (layer1_outputs(678)) or (layer1_outputs(2557));
    layer2_outputs(2272) <= not((layer1_outputs(2359)) and (layer1_outputs(1607)));
    layer2_outputs(2273) <= not((layer1_outputs(1425)) or (layer1_outputs(2226)));
    layer2_outputs(2274) <= not((layer1_outputs(2482)) or (layer1_outputs(1123)));
    layer2_outputs(2275) <= not(layer1_outputs(239)) or (layer1_outputs(1168));
    layer2_outputs(2276) <= not(layer1_outputs(1651));
    layer2_outputs(2277) <= (layer1_outputs(94)) and not (layer1_outputs(1305));
    layer2_outputs(2278) <= not(layer1_outputs(2238)) or (layer1_outputs(1833));
    layer2_outputs(2279) <= not(layer1_outputs(2376));
    layer2_outputs(2280) <= layer1_outputs(2024);
    layer2_outputs(2281) <= (layer1_outputs(293)) or (layer1_outputs(253));
    layer2_outputs(2282) <= layer1_outputs(2409);
    layer2_outputs(2283) <= not((layer1_outputs(684)) xor (layer1_outputs(1446)));
    layer2_outputs(2284) <= not(layer1_outputs(1652));
    layer2_outputs(2285) <= not(layer1_outputs(1448)) or (layer1_outputs(1080));
    layer2_outputs(2286) <= not(layer1_outputs(571));
    layer2_outputs(2287) <= (layer1_outputs(1911)) and not (layer1_outputs(1058));
    layer2_outputs(2288) <= not((layer1_outputs(957)) and (layer1_outputs(2468)));
    layer2_outputs(2289) <= not(layer1_outputs(1308));
    layer2_outputs(2290) <= not(layer1_outputs(269)) or (layer1_outputs(317));
    layer2_outputs(2291) <= '0';
    layer2_outputs(2292) <= (layer1_outputs(543)) and not (layer1_outputs(1519));
    layer2_outputs(2293) <= not(layer1_outputs(870));
    layer2_outputs(2294) <= layer1_outputs(2219);
    layer2_outputs(2295) <= not(layer1_outputs(345));
    layer2_outputs(2296) <= (layer1_outputs(1789)) and (layer1_outputs(1031));
    layer2_outputs(2297) <= not((layer1_outputs(644)) or (layer1_outputs(2033)));
    layer2_outputs(2298) <= (layer1_outputs(523)) or (layer1_outputs(808));
    layer2_outputs(2299) <= not(layer1_outputs(1205));
    layer2_outputs(2300) <= layer1_outputs(2171);
    layer2_outputs(2301) <= not(layer1_outputs(710)) or (layer1_outputs(200));
    layer2_outputs(2302) <= not((layer1_outputs(2222)) or (layer1_outputs(1851)));
    layer2_outputs(2303) <= (layer1_outputs(1400)) and not (layer1_outputs(441));
    layer2_outputs(2304) <= not(layer1_outputs(1647)) or (layer1_outputs(1129));
    layer2_outputs(2305) <= (layer1_outputs(691)) xor (layer1_outputs(642));
    layer2_outputs(2306) <= not(layer1_outputs(2456));
    layer2_outputs(2307) <= (layer1_outputs(2515)) and not (layer1_outputs(1182));
    layer2_outputs(2308) <= not(layer1_outputs(1219));
    layer2_outputs(2309) <= not(layer1_outputs(384)) or (layer1_outputs(970));
    layer2_outputs(2310) <= (layer1_outputs(2047)) and not (layer1_outputs(299));
    layer2_outputs(2311) <= not(layer1_outputs(1505));
    layer2_outputs(2312) <= (layer1_outputs(2181)) or (layer1_outputs(592));
    layer2_outputs(2313) <= (layer1_outputs(980)) and not (layer1_outputs(177));
    layer2_outputs(2314) <= not(layer1_outputs(266)) or (layer1_outputs(2422));
    layer2_outputs(2315) <= not((layer1_outputs(1431)) xor (layer1_outputs(877)));
    layer2_outputs(2316) <= (layer1_outputs(1085)) and not (layer1_outputs(836));
    layer2_outputs(2317) <= (layer1_outputs(2224)) and not (layer1_outputs(325));
    layer2_outputs(2318) <= layer1_outputs(978);
    layer2_outputs(2319) <= (layer1_outputs(1595)) and not (layer1_outputs(1032));
    layer2_outputs(2320) <= (layer1_outputs(143)) and (layer1_outputs(979));
    layer2_outputs(2321) <= '0';
    layer2_outputs(2322) <= not(layer1_outputs(655)) or (layer1_outputs(2282));
    layer2_outputs(2323) <= layer1_outputs(1240);
    layer2_outputs(2324) <= layer1_outputs(519);
    layer2_outputs(2325) <= layer1_outputs(1135);
    layer2_outputs(2326) <= layer1_outputs(25);
    layer2_outputs(2327) <= not(layer1_outputs(1975));
    layer2_outputs(2328) <= not(layer1_outputs(1985));
    layer2_outputs(2329) <= (layer1_outputs(944)) and not (layer1_outputs(1404));
    layer2_outputs(2330) <= layer1_outputs(27);
    layer2_outputs(2331) <= not(layer1_outputs(965));
    layer2_outputs(2332) <= not(layer1_outputs(2102));
    layer2_outputs(2333) <= not(layer1_outputs(1525));
    layer2_outputs(2334) <= not(layer1_outputs(1577)) or (layer1_outputs(988));
    layer2_outputs(2335) <= not(layer1_outputs(2155));
    layer2_outputs(2336) <= not(layer1_outputs(916)) or (layer1_outputs(2108));
    layer2_outputs(2337) <= layer1_outputs(735);
    layer2_outputs(2338) <= not((layer1_outputs(750)) or (layer1_outputs(983)));
    layer2_outputs(2339) <= layer1_outputs(273);
    layer2_outputs(2340) <= (layer1_outputs(1455)) and (layer1_outputs(1752));
    layer2_outputs(2341) <= not(layer1_outputs(2109)) or (layer1_outputs(457));
    layer2_outputs(2342) <= layer1_outputs(728);
    layer2_outputs(2343) <= not((layer1_outputs(1336)) or (layer1_outputs(490)));
    layer2_outputs(2344) <= not(layer1_outputs(197));
    layer2_outputs(2345) <= layer1_outputs(1433);
    layer2_outputs(2346) <= (layer1_outputs(153)) and not (layer1_outputs(897));
    layer2_outputs(2347) <= (layer1_outputs(835)) and (layer1_outputs(1052));
    layer2_outputs(2348) <= not(layer1_outputs(166));
    layer2_outputs(2349) <= layer1_outputs(1201);
    layer2_outputs(2350) <= not(layer1_outputs(2419)) or (layer1_outputs(69));
    layer2_outputs(2351) <= (layer1_outputs(2374)) and not (layer1_outputs(1266));
    layer2_outputs(2352) <= layer1_outputs(876);
    layer2_outputs(2353) <= (layer1_outputs(296)) or (layer1_outputs(1654));
    layer2_outputs(2354) <= not(layer1_outputs(544));
    layer2_outputs(2355) <= (layer1_outputs(1324)) and not (layer1_outputs(712));
    layer2_outputs(2356) <= layer1_outputs(1619);
    layer2_outputs(2357) <= not(layer1_outputs(1707));
    layer2_outputs(2358) <= (layer1_outputs(1788)) xor (layer1_outputs(1425));
    layer2_outputs(2359) <= not((layer1_outputs(2370)) or (layer1_outputs(1639)));
    layer2_outputs(2360) <= not((layer1_outputs(505)) or (layer1_outputs(543)));
    layer2_outputs(2361) <= layer1_outputs(2528);
    layer2_outputs(2362) <= (layer1_outputs(1822)) and (layer1_outputs(2228));
    layer2_outputs(2363) <= not(layer1_outputs(2538));
    layer2_outputs(2364) <= layer1_outputs(1887);
    layer2_outputs(2365) <= layer1_outputs(381);
    layer2_outputs(2366) <= (layer1_outputs(1682)) and not (layer1_outputs(473));
    layer2_outputs(2367) <= layer1_outputs(1872);
    layer2_outputs(2368) <= not(layer1_outputs(986)) or (layer1_outputs(1219));
    layer2_outputs(2369) <= not(layer1_outputs(621)) or (layer1_outputs(201));
    layer2_outputs(2370) <= (layer1_outputs(1915)) or (layer1_outputs(2269));
    layer2_outputs(2371) <= not(layer1_outputs(2272));
    layer2_outputs(2372) <= not(layer1_outputs(1014)) or (layer1_outputs(1084));
    layer2_outputs(2373) <= not(layer1_outputs(2441));
    layer2_outputs(2374) <= not((layer1_outputs(2194)) or (layer1_outputs(903)));
    layer2_outputs(2375) <= not((layer1_outputs(1324)) or (layer1_outputs(1381)));
    layer2_outputs(2376) <= layer1_outputs(402);
    layer2_outputs(2377) <= layer1_outputs(1040);
    layer2_outputs(2378) <= not(layer1_outputs(1003));
    layer2_outputs(2379) <= not((layer1_outputs(1390)) and (layer1_outputs(368)));
    layer2_outputs(2380) <= (layer1_outputs(129)) and (layer1_outputs(1830));
    layer2_outputs(2381) <= (layer1_outputs(2329)) and (layer1_outputs(388));
    layer2_outputs(2382) <= not(layer1_outputs(728));
    layer2_outputs(2383) <= layer1_outputs(1942);
    layer2_outputs(2384) <= not(layer1_outputs(225));
    layer2_outputs(2385) <= not((layer1_outputs(1120)) or (layer1_outputs(1075)));
    layer2_outputs(2386) <= layer1_outputs(888);
    layer2_outputs(2387) <= (layer1_outputs(1429)) and (layer1_outputs(310));
    layer2_outputs(2388) <= (layer1_outputs(227)) and (layer1_outputs(2126));
    layer2_outputs(2389) <= not(layer1_outputs(1931));
    layer2_outputs(2390) <= not((layer1_outputs(161)) and (layer1_outputs(954)));
    layer2_outputs(2391) <= not((layer1_outputs(1712)) and (layer1_outputs(385)));
    layer2_outputs(2392) <= (layer1_outputs(2447)) and not (layer1_outputs(2410));
    layer2_outputs(2393) <= not(layer1_outputs(197));
    layer2_outputs(2394) <= layer1_outputs(258);
    layer2_outputs(2395) <= '1';
    layer2_outputs(2396) <= not(layer1_outputs(2077)) or (layer1_outputs(2552));
    layer2_outputs(2397) <= not((layer1_outputs(727)) or (layer1_outputs(1835)));
    layer2_outputs(2398) <= (layer1_outputs(1697)) and not (layer1_outputs(419));
    layer2_outputs(2399) <= '1';
    layer2_outputs(2400) <= (layer1_outputs(1455)) and (layer1_outputs(175));
    layer2_outputs(2401) <= not(layer1_outputs(987));
    layer2_outputs(2402) <= not(layer1_outputs(820));
    layer2_outputs(2403) <= (layer1_outputs(2115)) and (layer1_outputs(354));
    layer2_outputs(2404) <= not(layer1_outputs(1215));
    layer2_outputs(2405) <= layer1_outputs(2263);
    layer2_outputs(2406) <= (layer1_outputs(246)) and not (layer1_outputs(1078));
    layer2_outputs(2407) <= layer1_outputs(2414);
    layer2_outputs(2408) <= layer1_outputs(1024);
    layer2_outputs(2409) <= (layer1_outputs(2345)) xor (layer1_outputs(2368));
    layer2_outputs(2410) <= layer1_outputs(62);
    layer2_outputs(2411) <= not(layer1_outputs(465));
    layer2_outputs(2412) <= not(layer1_outputs(582)) or (layer1_outputs(1794));
    layer2_outputs(2413) <= not(layer1_outputs(1205));
    layer2_outputs(2414) <= '1';
    layer2_outputs(2415) <= layer1_outputs(2151);
    layer2_outputs(2416) <= (layer1_outputs(1802)) and (layer1_outputs(2338));
    layer2_outputs(2417) <= not((layer1_outputs(471)) or (layer1_outputs(1257)));
    layer2_outputs(2418) <= (layer1_outputs(517)) and not (layer1_outputs(1735));
    layer2_outputs(2419) <= layer1_outputs(1105);
    layer2_outputs(2420) <= (layer1_outputs(1470)) and not (layer1_outputs(907));
    layer2_outputs(2421) <= not(layer1_outputs(599)) or (layer1_outputs(504));
    layer2_outputs(2422) <= (layer1_outputs(1357)) xor (layer1_outputs(2513));
    layer2_outputs(2423) <= not((layer1_outputs(91)) or (layer1_outputs(1878)));
    layer2_outputs(2424) <= not(layer1_outputs(1975)) or (layer1_outputs(393));
    layer2_outputs(2425) <= (layer1_outputs(98)) and not (layer1_outputs(386));
    layer2_outputs(2426) <= not((layer1_outputs(43)) and (layer1_outputs(272)));
    layer2_outputs(2427) <= layer1_outputs(872);
    layer2_outputs(2428) <= not(layer1_outputs(104));
    layer2_outputs(2429) <= not(layer1_outputs(42)) or (layer1_outputs(228));
    layer2_outputs(2430) <= '0';
    layer2_outputs(2431) <= (layer1_outputs(1340)) or (layer1_outputs(2218));
    layer2_outputs(2432) <= (layer1_outputs(991)) and not (layer1_outputs(1943));
    layer2_outputs(2433) <= (layer1_outputs(1386)) or (layer1_outputs(1353));
    layer2_outputs(2434) <= (layer1_outputs(2417)) or (layer1_outputs(1582));
    layer2_outputs(2435) <= not(layer1_outputs(168));
    layer2_outputs(2436) <= not(layer1_outputs(488));
    layer2_outputs(2437) <= (layer1_outputs(1559)) and not (layer1_outputs(1763));
    layer2_outputs(2438) <= not((layer1_outputs(2115)) and (layer1_outputs(752)));
    layer2_outputs(2439) <= (layer1_outputs(75)) or (layer1_outputs(1636));
    layer2_outputs(2440) <= not(layer1_outputs(2117)) or (layer1_outputs(2146));
    layer2_outputs(2441) <= not(layer1_outputs(929)) or (layer1_outputs(106));
    layer2_outputs(2442) <= not((layer1_outputs(376)) and (layer1_outputs(1497)));
    layer2_outputs(2443) <= not((layer1_outputs(108)) xor (layer1_outputs(1636)));
    layer2_outputs(2444) <= '1';
    layer2_outputs(2445) <= not(layer1_outputs(159));
    layer2_outputs(2446) <= not(layer1_outputs(542));
    layer2_outputs(2447) <= (layer1_outputs(265)) and not (layer1_outputs(1649));
    layer2_outputs(2448) <= layer1_outputs(2186);
    layer2_outputs(2449) <= layer1_outputs(880);
    layer2_outputs(2450) <= (layer1_outputs(2366)) and not (layer1_outputs(1006));
    layer2_outputs(2451) <= not((layer1_outputs(461)) and (layer1_outputs(1141)));
    layer2_outputs(2452) <= (layer1_outputs(1426)) and (layer1_outputs(1529));
    layer2_outputs(2453) <= not(layer1_outputs(554)) or (layer1_outputs(1345));
    layer2_outputs(2454) <= (layer1_outputs(458)) or (layer1_outputs(1533));
    layer2_outputs(2455) <= (layer1_outputs(204)) and (layer1_outputs(1909));
    layer2_outputs(2456) <= not(layer1_outputs(681));
    layer2_outputs(2457) <= not((layer1_outputs(462)) or (layer1_outputs(981)));
    layer2_outputs(2458) <= not(layer1_outputs(1966));
    layer2_outputs(2459) <= not((layer1_outputs(44)) or (layer1_outputs(600)));
    layer2_outputs(2460) <= (layer1_outputs(2145)) and (layer1_outputs(115));
    layer2_outputs(2461) <= (layer1_outputs(515)) xor (layer1_outputs(2448));
    layer2_outputs(2462) <= not(layer1_outputs(18));
    layer2_outputs(2463) <= (layer1_outputs(1990)) and (layer1_outputs(892));
    layer2_outputs(2464) <= not(layer1_outputs(1712)) or (layer1_outputs(1617));
    layer2_outputs(2465) <= layer1_outputs(643);
    layer2_outputs(2466) <= layer1_outputs(781);
    layer2_outputs(2467) <= not(layer1_outputs(1331)) or (layer1_outputs(285));
    layer2_outputs(2468) <= not(layer1_outputs(255)) or (layer1_outputs(2292));
    layer2_outputs(2469) <= layer1_outputs(778);
    layer2_outputs(2470) <= (layer1_outputs(1588)) xor (layer1_outputs(1241));
    layer2_outputs(2471) <= (layer1_outputs(2478)) and not (layer1_outputs(2298));
    layer2_outputs(2472) <= not((layer1_outputs(1604)) and (layer1_outputs(867)));
    layer2_outputs(2473) <= (layer1_outputs(2104)) and not (layer1_outputs(2051));
    layer2_outputs(2474) <= not(layer1_outputs(85)) or (layer1_outputs(767));
    layer2_outputs(2475) <= (layer1_outputs(664)) and not (layer1_outputs(2158));
    layer2_outputs(2476) <= '1';
    layer2_outputs(2477) <= not(layer1_outputs(2005));
    layer2_outputs(2478) <= layer1_outputs(33);
    layer2_outputs(2479) <= (layer1_outputs(1483)) and (layer1_outputs(1313));
    layer2_outputs(2480) <= '0';
    layer2_outputs(2481) <= not((layer1_outputs(1288)) or (layer1_outputs(415)));
    layer2_outputs(2482) <= layer1_outputs(2393);
    layer2_outputs(2483) <= (layer1_outputs(2529)) and not (layer1_outputs(1881));
    layer2_outputs(2484) <= (layer1_outputs(2143)) and not (layer1_outputs(1587));
    layer2_outputs(2485) <= (layer1_outputs(1530)) and not (layer1_outputs(2031));
    layer2_outputs(2486) <= not((layer1_outputs(1852)) or (layer1_outputs(1621)));
    layer2_outputs(2487) <= layer1_outputs(2206);
    layer2_outputs(2488) <= layer1_outputs(1618);
    layer2_outputs(2489) <= layer1_outputs(97);
    layer2_outputs(2490) <= layer1_outputs(1389);
    layer2_outputs(2491) <= (layer1_outputs(572)) and not (layer1_outputs(1819));
    layer2_outputs(2492) <= not((layer1_outputs(674)) or (layer1_outputs(1073)));
    layer2_outputs(2493) <= (layer1_outputs(1989)) and not (layer1_outputs(2507));
    layer2_outputs(2494) <= not(layer1_outputs(22));
    layer2_outputs(2495) <= layer1_outputs(355);
    layer2_outputs(2496) <= (layer1_outputs(2280)) and not (layer1_outputs(1519));
    layer2_outputs(2497) <= not((layer1_outputs(1755)) or (layer1_outputs(2489)));
    layer2_outputs(2498) <= not(layer1_outputs(846)) or (layer1_outputs(1839));
    layer2_outputs(2499) <= not(layer1_outputs(2507));
    layer2_outputs(2500) <= layer1_outputs(2418);
    layer2_outputs(2501) <= not(layer1_outputs(2331)) or (layer1_outputs(1148));
    layer2_outputs(2502) <= (layer1_outputs(1827)) and not (layer1_outputs(2020));
    layer2_outputs(2503) <= (layer1_outputs(2154)) and (layer1_outputs(1466));
    layer2_outputs(2504) <= not(layer1_outputs(1717)) or (layer1_outputs(2424));
    layer2_outputs(2505) <= not(layer1_outputs(1177));
    layer2_outputs(2506) <= layer1_outputs(1593);
    layer2_outputs(2507) <= (layer1_outputs(209)) xor (layer1_outputs(1447));
    layer2_outputs(2508) <= not(layer1_outputs(2327));
    layer2_outputs(2509) <= (layer1_outputs(1777)) and (layer1_outputs(1279));
    layer2_outputs(2510) <= layer1_outputs(449);
    layer2_outputs(2511) <= not((layer1_outputs(1168)) xor (layer1_outputs(1440)));
    layer2_outputs(2512) <= not(layer1_outputs(545)) or (layer1_outputs(446));
    layer2_outputs(2513) <= (layer1_outputs(588)) and not (layer1_outputs(1053));
    layer2_outputs(2514) <= not((layer1_outputs(335)) and (layer1_outputs(1983)));
    layer2_outputs(2515) <= (layer1_outputs(1158)) and (layer1_outputs(101));
    layer2_outputs(2516) <= (layer1_outputs(328)) and not (layer1_outputs(1412));
    layer2_outputs(2517) <= '0';
    layer2_outputs(2518) <= layer1_outputs(980);
    layer2_outputs(2519) <= layer1_outputs(278);
    layer2_outputs(2520) <= not(layer1_outputs(162));
    layer2_outputs(2521) <= not((layer1_outputs(1386)) or (layer1_outputs(1892)));
    layer2_outputs(2522) <= (layer1_outputs(918)) and not (layer1_outputs(1484));
    layer2_outputs(2523) <= not((layer1_outputs(1561)) and (layer1_outputs(1743)));
    layer2_outputs(2524) <= not(layer1_outputs(2004)) or (layer1_outputs(1354));
    layer2_outputs(2525) <= (layer1_outputs(2167)) and not (layer1_outputs(2211));
    layer2_outputs(2526) <= not((layer1_outputs(874)) or (layer1_outputs(2245)));
    layer2_outputs(2527) <= (layer1_outputs(1729)) and not (layer1_outputs(684));
    layer2_outputs(2528) <= layer1_outputs(346);
    layer2_outputs(2529) <= not(layer1_outputs(408)) or (layer1_outputs(831));
    layer2_outputs(2530) <= not((layer1_outputs(776)) and (layer1_outputs(625)));
    layer2_outputs(2531) <= (layer1_outputs(1293)) or (layer1_outputs(1563));
    layer2_outputs(2532) <= layer1_outputs(129);
    layer2_outputs(2533) <= (layer1_outputs(530)) or (layer1_outputs(1523));
    layer2_outputs(2534) <= not((layer1_outputs(370)) and (layer1_outputs(2330)));
    layer2_outputs(2535) <= (layer1_outputs(870)) and not (layer1_outputs(977));
    layer2_outputs(2536) <= not(layer1_outputs(102));
    layer2_outputs(2537) <= (layer1_outputs(1326)) or (layer1_outputs(831));
    layer2_outputs(2538) <= '0';
    layer2_outputs(2539) <= not(layer1_outputs(998));
    layer2_outputs(2540) <= not(layer1_outputs(609));
    layer2_outputs(2541) <= '1';
    layer2_outputs(2542) <= layer1_outputs(325);
    layer2_outputs(2543) <= not(layer1_outputs(262)) or (layer1_outputs(951));
    layer2_outputs(2544) <= (layer1_outputs(1329)) and (layer1_outputs(2416));
    layer2_outputs(2545) <= (layer1_outputs(764)) xor (layer1_outputs(369));
    layer2_outputs(2546) <= (layer1_outputs(979)) or (layer1_outputs(680));
    layer2_outputs(2547) <= (layer1_outputs(786)) and not (layer1_outputs(581));
    layer2_outputs(2548) <= not((layer1_outputs(2470)) and (layer1_outputs(807)));
    layer2_outputs(2549) <= (layer1_outputs(1537)) and not (layer1_outputs(801));
    layer2_outputs(2550) <= not((layer1_outputs(863)) xor (layer1_outputs(548)));
    layer2_outputs(2551) <= not((layer1_outputs(99)) xor (layer1_outputs(1738)));
    layer2_outputs(2552) <= not(layer1_outputs(1339));
    layer2_outputs(2553) <= not((layer1_outputs(1076)) xor (layer1_outputs(334)));
    layer2_outputs(2554) <= not((layer1_outputs(509)) and (layer1_outputs(2074)));
    layer2_outputs(2555) <= (layer1_outputs(1110)) xor (layer1_outputs(1520));
    layer2_outputs(2556) <= not(layer1_outputs(630));
    layer2_outputs(2557) <= layer1_outputs(1940);
    layer2_outputs(2558) <= (layer1_outputs(1023)) and (layer1_outputs(928));
    layer2_outputs(2559) <= not((layer1_outputs(818)) xor (layer1_outputs(259)));
    outputs(0) <= layer2_outputs(1257);
    outputs(1) <= (layer2_outputs(918)) and (layer2_outputs(1202));
    outputs(2) <= not(layer2_outputs(223)) or (layer2_outputs(729));
    outputs(3) <= layer2_outputs(1583);
    outputs(4) <= (layer2_outputs(1803)) and (layer2_outputs(730));
    outputs(5) <= layer2_outputs(643);
    outputs(6) <= not(layer2_outputs(91)) or (layer2_outputs(2215));
    outputs(7) <= not((layer2_outputs(307)) or (layer2_outputs(564)));
    outputs(8) <= layer2_outputs(556);
    outputs(9) <= not(layer2_outputs(2015));
    outputs(10) <= not(layer2_outputs(1815)) or (layer2_outputs(1905));
    outputs(11) <= (layer2_outputs(243)) xor (layer2_outputs(1420));
    outputs(12) <= layer2_outputs(2269);
    outputs(13) <= (layer2_outputs(75)) and not (layer2_outputs(1982));
    outputs(14) <= (layer2_outputs(1807)) xor (layer2_outputs(1052));
    outputs(15) <= not(layer2_outputs(1684));
    outputs(16) <= not(layer2_outputs(1291));
    outputs(17) <= (layer2_outputs(2173)) and (layer2_outputs(497));
    outputs(18) <= (layer2_outputs(746)) and (layer2_outputs(2138));
    outputs(19) <= (layer2_outputs(2256)) and not (layer2_outputs(2049));
    outputs(20) <= layer2_outputs(15);
    outputs(21) <= layer2_outputs(346);
    outputs(22) <= (layer2_outputs(450)) and not (layer2_outputs(1436));
    outputs(23) <= (layer2_outputs(1395)) and (layer2_outputs(355));
    outputs(24) <= not((layer2_outputs(1283)) or (layer2_outputs(1982)));
    outputs(25) <= layer2_outputs(1019);
    outputs(26) <= layer2_outputs(1845);
    outputs(27) <= not(layer2_outputs(2319));
    outputs(28) <= (layer2_outputs(327)) xor (layer2_outputs(793));
    outputs(29) <= (layer2_outputs(370)) and (layer2_outputs(2423));
    outputs(30) <= not(layer2_outputs(2515));
    outputs(31) <= not(layer2_outputs(885));
    outputs(32) <= not(layer2_outputs(1891));
    outputs(33) <= (layer2_outputs(1987)) or (layer2_outputs(2277));
    outputs(34) <= not((layer2_outputs(2365)) and (layer2_outputs(286)));
    outputs(35) <= not(layer2_outputs(1272));
    outputs(36) <= (layer2_outputs(2277)) or (layer2_outputs(1656));
    outputs(37) <= not(layer2_outputs(2163)) or (layer2_outputs(1690));
    outputs(38) <= not(layer2_outputs(844));
    outputs(39) <= not(layer2_outputs(2273));
    outputs(40) <= not(layer2_outputs(1545));
    outputs(41) <= layer2_outputs(926);
    outputs(42) <= layer2_outputs(354);
    outputs(43) <= not((layer2_outputs(2283)) and (layer2_outputs(2254)));
    outputs(44) <= layer2_outputs(74);
    outputs(45) <= not(layer2_outputs(517));
    outputs(46) <= not((layer2_outputs(511)) xor (layer2_outputs(853)));
    outputs(47) <= not(layer2_outputs(800)) or (layer2_outputs(785));
    outputs(48) <= (layer2_outputs(2197)) and (layer2_outputs(879));
    outputs(49) <= (layer2_outputs(55)) or (layer2_outputs(457));
    outputs(50) <= layer2_outputs(1192);
    outputs(51) <= layer2_outputs(1202);
    outputs(52) <= (layer2_outputs(2016)) and not (layer2_outputs(2288));
    outputs(53) <= not(layer2_outputs(309));
    outputs(54) <= not(layer2_outputs(212)) or (layer2_outputs(1838));
    outputs(55) <= not((layer2_outputs(1252)) and (layer2_outputs(1020)));
    outputs(56) <= (layer2_outputs(1413)) and not (layer2_outputs(204));
    outputs(57) <= layer2_outputs(2408);
    outputs(58) <= not(layer2_outputs(1302));
    outputs(59) <= not(layer2_outputs(108));
    outputs(60) <= not((layer2_outputs(296)) or (layer2_outputs(1529)));
    outputs(61) <= not((layer2_outputs(32)) and (layer2_outputs(2210)));
    outputs(62) <= (layer2_outputs(1244)) and (layer2_outputs(405));
    outputs(63) <= layer2_outputs(1385);
    outputs(64) <= layer2_outputs(1595);
    outputs(65) <= (layer2_outputs(1147)) and not (layer2_outputs(1973));
    outputs(66) <= layer2_outputs(111);
    outputs(67) <= layer2_outputs(128);
    outputs(68) <= not(layer2_outputs(1030));
    outputs(69) <= not(layer2_outputs(161));
    outputs(70) <= not((layer2_outputs(1664)) or (layer2_outputs(1914)));
    outputs(71) <= not(layer2_outputs(1419));
    outputs(72) <= layer2_outputs(2157);
    outputs(73) <= not(layer2_outputs(629));
    outputs(74) <= not(layer2_outputs(2427)) or (layer2_outputs(1894));
    outputs(75) <= not((layer2_outputs(1637)) xor (layer2_outputs(987)));
    outputs(76) <= not(layer2_outputs(1350)) or (layer2_outputs(2230));
    outputs(77) <= layer2_outputs(1147);
    outputs(78) <= not(layer2_outputs(667));
    outputs(79) <= layer2_outputs(1434);
    outputs(80) <= not(layer2_outputs(762));
    outputs(81) <= not(layer2_outputs(492));
    outputs(82) <= layer2_outputs(344);
    outputs(83) <= layer2_outputs(689);
    outputs(84) <= (layer2_outputs(1096)) and not (layer2_outputs(1195));
    outputs(85) <= (layer2_outputs(1002)) and not (layer2_outputs(612));
    outputs(86) <= (layer2_outputs(278)) and not (layer2_outputs(1804));
    outputs(87) <= layer2_outputs(551);
    outputs(88) <= not((layer2_outputs(1814)) or (layer2_outputs(1994)));
    outputs(89) <= not(layer2_outputs(2424));
    outputs(90) <= (layer2_outputs(251)) xor (layer2_outputs(1684));
    outputs(91) <= (layer2_outputs(1412)) and not (layer2_outputs(436));
    outputs(92) <= not(layer2_outputs(387));
    outputs(93) <= not((layer2_outputs(348)) or (layer2_outputs(778)));
    outputs(94) <= not(layer2_outputs(1937));
    outputs(95) <= layer2_outputs(2201);
    outputs(96) <= layer2_outputs(1230);
    outputs(97) <= layer2_outputs(1965);
    outputs(98) <= not(layer2_outputs(880));
    outputs(99) <= layer2_outputs(1415);
    outputs(100) <= layer2_outputs(1374);
    outputs(101) <= not((layer2_outputs(2232)) or (layer2_outputs(2535)));
    outputs(102) <= layer2_outputs(920);
    outputs(103) <= layer2_outputs(261);
    outputs(104) <= not(layer2_outputs(380));
    outputs(105) <= not(layer2_outputs(1274)) or (layer2_outputs(1817));
    outputs(106) <= layer2_outputs(386);
    outputs(107) <= not(layer2_outputs(1740));
    outputs(108) <= (layer2_outputs(1948)) and not (layer2_outputs(315));
    outputs(109) <= (layer2_outputs(1148)) xor (layer2_outputs(1725));
    outputs(110) <= not(layer2_outputs(1081));
    outputs(111) <= not(layer2_outputs(269));
    outputs(112) <= (layer2_outputs(45)) or (layer2_outputs(1239));
    outputs(113) <= (layer2_outputs(2006)) and (layer2_outputs(985));
    outputs(114) <= layer2_outputs(2215);
    outputs(115) <= not(layer2_outputs(1116));
    outputs(116) <= layer2_outputs(1547);
    outputs(117) <= not(layer2_outputs(1368));
    outputs(118) <= (layer2_outputs(825)) and (layer2_outputs(1125));
    outputs(119) <= layer2_outputs(121);
    outputs(120) <= (layer2_outputs(815)) and (layer2_outputs(934));
    outputs(121) <= layer2_outputs(1917);
    outputs(122) <= (layer2_outputs(561)) and not (layer2_outputs(1296));
    outputs(123) <= not((layer2_outputs(1342)) or (layer2_outputs(1683)));
    outputs(124) <= layer2_outputs(1547);
    outputs(125) <= not((layer2_outputs(2051)) xor (layer2_outputs(878)));
    outputs(126) <= (layer2_outputs(207)) and not (layer2_outputs(1429));
    outputs(127) <= not(layer2_outputs(602));
    outputs(128) <= not(layer2_outputs(461));
    outputs(129) <= layer2_outputs(258);
    outputs(130) <= layer2_outputs(1778);
    outputs(131) <= layer2_outputs(1580);
    outputs(132) <= not((layer2_outputs(1394)) xor (layer2_outputs(2538)));
    outputs(133) <= (layer2_outputs(449)) and (layer2_outputs(1607));
    outputs(134) <= not(layer2_outputs(1128)) or (layer2_outputs(2126));
    outputs(135) <= (layer2_outputs(658)) and not (layer2_outputs(1133));
    outputs(136) <= not(layer2_outputs(1836));
    outputs(137) <= not(layer2_outputs(900));
    outputs(138) <= layer2_outputs(1925);
    outputs(139) <= layer2_outputs(1733);
    outputs(140) <= not(layer2_outputs(891)) or (layer2_outputs(898));
    outputs(141) <= layer2_outputs(933);
    outputs(142) <= layer2_outputs(43);
    outputs(143) <= layer2_outputs(2463);
    outputs(144) <= (layer2_outputs(1951)) and not (layer2_outputs(1530));
    outputs(145) <= layer2_outputs(1402);
    outputs(146) <= (layer2_outputs(1791)) and (layer2_outputs(1687));
    outputs(147) <= not(layer2_outputs(1040));
    outputs(148) <= (layer2_outputs(982)) and not (layer2_outputs(394));
    outputs(149) <= (layer2_outputs(784)) and (layer2_outputs(854));
    outputs(150) <= not(layer2_outputs(2363));
    outputs(151) <= layer2_outputs(546);
    outputs(152) <= not(layer2_outputs(324));
    outputs(153) <= layer2_outputs(825);
    outputs(154) <= not(layer2_outputs(817));
    outputs(155) <= (layer2_outputs(1774)) and not (layer2_outputs(507));
    outputs(156) <= (layer2_outputs(1619)) and not (layer2_outputs(657));
    outputs(157) <= layer2_outputs(2213);
    outputs(158) <= not(layer2_outputs(741));
    outputs(159) <= not((layer2_outputs(1646)) or (layer2_outputs(2511)));
    outputs(160) <= (layer2_outputs(2012)) and not (layer2_outputs(1847));
    outputs(161) <= layer2_outputs(300);
    outputs(162) <= not(layer2_outputs(368));
    outputs(163) <= not((layer2_outputs(1401)) xor (layer2_outputs(2505)));
    outputs(164) <= not(layer2_outputs(151));
    outputs(165) <= not(layer2_outputs(1798));
    outputs(166) <= not(layer2_outputs(69)) or (layer2_outputs(1816));
    outputs(167) <= (layer2_outputs(946)) and not (layer2_outputs(394));
    outputs(168) <= not(layer2_outputs(662));
    outputs(169) <= layer2_outputs(1795);
    outputs(170) <= not(layer2_outputs(527));
    outputs(171) <= not((layer2_outputs(1539)) or (layer2_outputs(101)));
    outputs(172) <= not((layer2_outputs(1802)) xor (layer2_outputs(554)));
    outputs(173) <= not(layer2_outputs(564)) or (layer2_outputs(1764));
    outputs(174) <= (layer2_outputs(1623)) or (layer2_outputs(445));
    outputs(175) <= layer2_outputs(503);
    outputs(176) <= not(layer2_outputs(1223));
    outputs(177) <= not(layer2_outputs(2061));
    outputs(178) <= not(layer2_outputs(2474));
    outputs(179) <= not((layer2_outputs(2473)) or (layer2_outputs(1156)));
    outputs(180) <= (layer2_outputs(175)) and not (layer2_outputs(1787));
    outputs(181) <= not(layer2_outputs(964));
    outputs(182) <= (layer2_outputs(704)) or (layer2_outputs(546));
    outputs(183) <= (layer2_outputs(1022)) and (layer2_outputs(2156));
    outputs(184) <= (layer2_outputs(2453)) and not (layer2_outputs(2263));
    outputs(185) <= not((layer2_outputs(988)) or (layer2_outputs(2393)));
    outputs(186) <= layer2_outputs(897);
    outputs(187) <= not(layer2_outputs(229));
    outputs(188) <= not((layer2_outputs(1738)) and (layer2_outputs(599)));
    outputs(189) <= not(layer2_outputs(915));
    outputs(190) <= (layer2_outputs(1146)) and not (layer2_outputs(1648));
    outputs(191) <= layer2_outputs(1898);
    outputs(192) <= not(layer2_outputs(2067));
    outputs(193) <= not(layer2_outputs(454));
    outputs(194) <= layer2_outputs(1682);
    outputs(195) <= not(layer2_outputs(288));
    outputs(196) <= not(layer2_outputs(719)) or (layer2_outputs(190));
    outputs(197) <= (layer2_outputs(887)) and not (layer2_outputs(1259));
    outputs(198) <= layer2_outputs(1526);
    outputs(199) <= not(layer2_outputs(2554)) or (layer2_outputs(2389));
    outputs(200) <= not(layer2_outputs(2171));
    outputs(201) <= layer2_outputs(42);
    outputs(202) <= (layer2_outputs(2522)) or (layer2_outputs(503));
    outputs(203) <= not(layer2_outputs(1620)) or (layer2_outputs(645));
    outputs(204) <= not(layer2_outputs(651)) or (layer2_outputs(1168));
    outputs(205) <= not(layer2_outputs(1752)) or (layer2_outputs(1593));
    outputs(206) <= layer2_outputs(185);
    outputs(207) <= not(layer2_outputs(1106));
    outputs(208) <= not(layer2_outputs(141));
    outputs(209) <= (layer2_outputs(2440)) or (layer2_outputs(675));
    outputs(210) <= not((layer2_outputs(888)) or (layer2_outputs(642)));
    outputs(211) <= not(layer2_outputs(1309));
    outputs(212) <= layer2_outputs(1489);
    outputs(213) <= not(layer2_outputs(1114));
    outputs(214) <= layer2_outputs(217);
    outputs(215) <= (layer2_outputs(2048)) and not (layer2_outputs(1694));
    outputs(216) <= (layer2_outputs(563)) and not (layer2_outputs(1260));
    outputs(217) <= not((layer2_outputs(2481)) xor (layer2_outputs(2031)));
    outputs(218) <= not(layer2_outputs(1256));
    outputs(219) <= not(layer2_outputs(271));
    outputs(220) <= not((layer2_outputs(837)) xor (layer2_outputs(1812)));
    outputs(221) <= (layer2_outputs(116)) and not (layer2_outputs(1446));
    outputs(222) <= not(layer2_outputs(1178));
    outputs(223) <= not(layer2_outputs(861));
    outputs(224) <= not((layer2_outputs(1992)) xor (layer2_outputs(2116)));
    outputs(225) <= (layer2_outputs(2124)) or (layer2_outputs(1009));
    outputs(226) <= not(layer2_outputs(1928));
    outputs(227) <= not(layer2_outputs(1913));
    outputs(228) <= not(layer2_outputs(2340)) or (layer2_outputs(1978));
    outputs(229) <= (layer2_outputs(1402)) and not (layer2_outputs(1820));
    outputs(230) <= layer2_outputs(1067);
    outputs(231) <= not(layer2_outputs(2001));
    outputs(232) <= layer2_outputs(291);
    outputs(233) <= not(layer2_outputs(2328));
    outputs(234) <= not((layer2_outputs(1529)) and (layer2_outputs(255)));
    outputs(235) <= layer2_outputs(329);
    outputs(236) <= not(layer2_outputs(1937));
    outputs(237) <= layer2_outputs(103);
    outputs(238) <= (layer2_outputs(2534)) and not (layer2_outputs(218));
    outputs(239) <= not(layer2_outputs(1659)) or (layer2_outputs(645));
    outputs(240) <= not(layer2_outputs(425));
    outputs(241) <= not(layer2_outputs(1211)) or (layer2_outputs(1986));
    outputs(242) <= not(layer2_outputs(1426));
    outputs(243) <= not(layer2_outputs(1260));
    outputs(244) <= layer2_outputs(1251);
    outputs(245) <= (layer2_outputs(1057)) and not (layer2_outputs(157));
    outputs(246) <= (layer2_outputs(1329)) and (layer2_outputs(946));
    outputs(247) <= layer2_outputs(1089);
    outputs(248) <= (layer2_outputs(1593)) and (layer2_outputs(1775));
    outputs(249) <= not(layer2_outputs(2276));
    outputs(250) <= (layer2_outputs(580)) and not (layer2_outputs(1319));
    outputs(251) <= (layer2_outputs(1392)) and (layer2_outputs(1365));
    outputs(252) <= layer2_outputs(1662);
    outputs(253) <= not((layer2_outputs(2204)) or (layer2_outputs(2274)));
    outputs(254) <= (layer2_outputs(728)) and not (layer2_outputs(1100));
    outputs(255) <= layer2_outputs(1685);
    outputs(256) <= (layer2_outputs(914)) and not (layer2_outputs(1203));
    outputs(257) <= (layer2_outputs(521)) and not (layer2_outputs(326));
    outputs(258) <= layer2_outputs(2159);
    outputs(259) <= (layer2_outputs(702)) and not (layer2_outputs(1976));
    outputs(260) <= (layer2_outputs(2063)) and not (layer2_outputs(1380));
    outputs(261) <= not((layer2_outputs(1170)) or (layer2_outputs(424)));
    outputs(262) <= layer2_outputs(1842);
    outputs(263) <= not(layer2_outputs(491));
    outputs(264) <= (layer2_outputs(2320)) and not (layer2_outputs(2533));
    outputs(265) <= not(layer2_outputs(280));
    outputs(266) <= (layer2_outputs(1554)) and not (layer2_outputs(1806));
    outputs(267) <= not(layer2_outputs(1135));
    outputs(268) <= (layer2_outputs(1589)) and (layer2_outputs(469));
    outputs(269) <= layer2_outputs(1007);
    outputs(270) <= not((layer2_outputs(1784)) or (layer2_outputs(1591)));
    outputs(271) <= not((layer2_outputs(233)) or (layer2_outputs(398)));
    outputs(272) <= layer2_outputs(467);
    outputs(273) <= (layer2_outputs(1451)) and not (layer2_outputs(767));
    outputs(274) <= not((layer2_outputs(2181)) xor (layer2_outputs(2303)));
    outputs(275) <= not(layer2_outputs(1840));
    outputs(276) <= not((layer2_outputs(1510)) xor (layer2_outputs(293)));
    outputs(277) <= not((layer2_outputs(1218)) or (layer2_outputs(171)));
    outputs(278) <= (layer2_outputs(457)) and not (layer2_outputs(875));
    outputs(279) <= (layer2_outputs(2062)) or (layer2_outputs(243));
    outputs(280) <= (layer2_outputs(683)) and (layer2_outputs(2022));
    outputs(281) <= not(layer2_outputs(316));
    outputs(282) <= (layer2_outputs(896)) and not (layer2_outputs(2440));
    outputs(283) <= not((layer2_outputs(1313)) or (layer2_outputs(588)));
    outputs(284) <= (layer2_outputs(1815)) and (layer2_outputs(1079));
    outputs(285) <= layer2_outputs(734);
    outputs(286) <= (layer2_outputs(625)) and not (layer2_outputs(1983));
    outputs(287) <= not(layer2_outputs(1796));
    outputs(288) <= not((layer2_outputs(1838)) or (layer2_outputs(271)));
    outputs(289) <= not((layer2_outputs(1850)) or (layer2_outputs(2150)));
    outputs(290) <= (layer2_outputs(640)) and (layer2_outputs(1041));
    outputs(291) <= not((layer2_outputs(1092)) or (layer2_outputs(1119)));
    outputs(292) <= (layer2_outputs(1899)) and not (layer2_outputs(1828));
    outputs(293) <= (layer2_outputs(2331)) and not (layer2_outputs(371));
    outputs(294) <= (layer2_outputs(988)) and not (layer2_outputs(892));
    outputs(295) <= layer2_outputs(61);
    outputs(296) <= (layer2_outputs(1311)) and not (layer2_outputs(213));
    outputs(297) <= not(layer2_outputs(1334));
    outputs(298) <= not(layer2_outputs(1277));
    outputs(299) <= (layer2_outputs(912)) and not (layer2_outputs(1835));
    outputs(300) <= not(layer2_outputs(1618));
    outputs(301) <= (layer2_outputs(1085)) and (layer2_outputs(1327));
    outputs(302) <= layer2_outputs(957);
    outputs(303) <= not(layer2_outputs(1727));
    outputs(304) <= not(layer2_outputs(1951));
    outputs(305) <= (layer2_outputs(1005)) and not (layer2_outputs(145));
    outputs(306) <= (layer2_outputs(2113)) and (layer2_outputs(2170));
    outputs(307) <= (layer2_outputs(52)) and not (layer2_outputs(1990));
    outputs(308) <= not(layer2_outputs(67));
    outputs(309) <= (layer2_outputs(2482)) and not (layer2_outputs(828));
    outputs(310) <= not(layer2_outputs(326));
    outputs(311) <= not(layer2_outputs(1162));
    outputs(312) <= (layer2_outputs(547)) and not (layer2_outputs(490));
    outputs(313) <= (layer2_outputs(880)) and (layer2_outputs(2270));
    outputs(314) <= (layer2_outputs(1472)) and not (layer2_outputs(2241));
    outputs(315) <= not(layer2_outputs(2046));
    outputs(316) <= (layer2_outputs(1213)) and not (layer2_outputs(260));
    outputs(317) <= (layer2_outputs(1739)) and (layer2_outputs(1824));
    outputs(318) <= not((layer2_outputs(562)) and (layer2_outputs(2260)));
    outputs(319) <= (layer2_outputs(1558)) and not (layer2_outputs(1628));
    outputs(320) <= not(layer2_outputs(1777));
    outputs(321) <= not(layer2_outputs(1770));
    outputs(322) <= (layer2_outputs(1953)) and not (layer2_outputs(1939));
    outputs(323) <= layer2_outputs(2133);
    outputs(324) <= layer2_outputs(2465);
    outputs(325) <= not((layer2_outputs(2538)) or (layer2_outputs(1132)));
    outputs(326) <= (layer2_outputs(1869)) and not (layer2_outputs(754));
    outputs(327) <= (layer2_outputs(1229)) and not (layer2_outputs(777));
    outputs(328) <= (layer2_outputs(181)) and (layer2_outputs(981));
    outputs(329) <= (layer2_outputs(1950)) and (layer2_outputs(670));
    outputs(330) <= (layer2_outputs(1789)) and not (layer2_outputs(491));
    outputs(331) <= (layer2_outputs(1735)) and (layer2_outputs(760));
    outputs(332) <= not(layer2_outputs(1356));
    outputs(333) <= (layer2_outputs(440)) and not (layer2_outputs(708));
    outputs(334) <= (layer2_outputs(2151)) and (layer2_outputs(68));
    outputs(335) <= (layer2_outputs(198)) and not (layer2_outputs(2438));
    outputs(336) <= (layer2_outputs(494)) and (layer2_outputs(1722));
    outputs(337) <= (layer2_outputs(903)) and not (layer2_outputs(2039));
    outputs(338) <= layer2_outputs(755);
    outputs(339) <= (layer2_outputs(209)) and (layer2_outputs(1071));
    outputs(340) <= (layer2_outputs(2217)) and not (layer2_outputs(396));
    outputs(341) <= (layer2_outputs(2392)) and (layer2_outputs(2183));
    outputs(342) <= (layer2_outputs(1707)) and not (layer2_outputs(1817));
    outputs(343) <= not((layer2_outputs(1544)) xor (layer2_outputs(78)));
    outputs(344) <= (layer2_outputs(378)) and not (layer2_outputs(2143));
    outputs(345) <= not((layer2_outputs(2410)) xor (layer2_outputs(934)));
    outputs(346) <= layer2_outputs(2381);
    outputs(347) <= layer2_outputs(1427);
    outputs(348) <= (layer2_outputs(2070)) and (layer2_outputs(748));
    outputs(349) <= layer2_outputs(1991);
    outputs(350) <= (layer2_outputs(1883)) and (layer2_outputs(1879));
    outputs(351) <= (layer2_outputs(267)) and not (layer2_outputs(2226));
    outputs(352) <= (layer2_outputs(1140)) and not (layer2_outputs(13));
    outputs(353) <= layer2_outputs(476);
    outputs(354) <= layer2_outputs(1267);
    outputs(355) <= (layer2_outputs(1429)) and not (layer2_outputs(1328));
    outputs(356) <= not((layer2_outputs(2080)) xor (layer2_outputs(1314)));
    outputs(357) <= (layer2_outputs(32)) and not (layer2_outputs(2336));
    outputs(358) <= layer2_outputs(241);
    outputs(359) <= layer2_outputs(239);
    outputs(360) <= not(layer2_outputs(573));
    outputs(361) <= (layer2_outputs(558)) and not (layer2_outputs(144));
    outputs(362) <= (layer2_outputs(1632)) and not (layer2_outputs(390));
    outputs(363) <= (layer2_outputs(320)) and (layer2_outputs(2136));
    outputs(364) <= (layer2_outputs(2378)) and not (layer2_outputs(450));
    outputs(365) <= not(layer2_outputs(2223));
    outputs(366) <= not((layer2_outputs(1711)) or (layer2_outputs(2293)));
    outputs(367) <= (layer2_outputs(611)) and (layer2_outputs(1247));
    outputs(368) <= (layer2_outputs(2329)) and not (layer2_outputs(413));
    outputs(369) <= not((layer2_outputs(1096)) or (layer2_outputs(1159)));
    outputs(370) <= layer2_outputs(1134);
    outputs(371) <= not((layer2_outputs(2558)) xor (layer2_outputs(2076)));
    outputs(372) <= (layer2_outputs(1312)) and not (layer2_outputs(2018));
    outputs(373) <= (layer2_outputs(1416)) and not (layer2_outputs(30));
    outputs(374) <= not(layer2_outputs(1234));
    outputs(375) <= (layer2_outputs(2077)) and (layer2_outputs(2356));
    outputs(376) <= (layer2_outputs(1015)) and (layer2_outputs(2319));
    outputs(377) <= layer2_outputs(2556);
    outputs(378) <= not((layer2_outputs(942)) or (layer2_outputs(1370)));
    outputs(379) <= (layer2_outputs(964)) and not (layer2_outputs(1383));
    outputs(380) <= (layer2_outputs(1443)) and not (layer2_outputs(2285));
    outputs(381) <= not((layer2_outputs(1238)) or (layer2_outputs(1760)));
    outputs(382) <= (layer2_outputs(2526)) and not (layer2_outputs(585));
    outputs(383) <= layer2_outputs(682);
    outputs(384) <= (layer2_outputs(2366)) and (layer2_outputs(967));
    outputs(385) <= (layer2_outputs(653)) or (layer2_outputs(2071));
    outputs(386) <= layer2_outputs(1417);
    outputs(387) <= not(layer2_outputs(1851));
    outputs(388) <= layer2_outputs(194);
    outputs(389) <= not(layer2_outputs(1741));
    outputs(390) <= (layer2_outputs(2008)) and (layer2_outputs(1175));
    outputs(391) <= layer2_outputs(1005);
    outputs(392) <= (layer2_outputs(2377)) and not (layer2_outputs(2367));
    outputs(393) <= (layer2_outputs(709)) or (layer2_outputs(1186));
    outputs(394) <= (layer2_outputs(1634)) and not (layer2_outputs(106));
    outputs(395) <= (layer2_outputs(2033)) and not (layer2_outputs(1192));
    outputs(396) <= (layer2_outputs(1548)) xor (layer2_outputs(742));
    outputs(397) <= (layer2_outputs(2418)) and (layer2_outputs(2041));
    outputs(398) <= (layer2_outputs(1837)) and (layer2_outputs(899));
    outputs(399) <= (layer2_outputs(2435)) and not (layer2_outputs(1241));
    outputs(400) <= (layer2_outputs(2383)) and (layer2_outputs(761));
    outputs(401) <= (layer2_outputs(2479)) and (layer2_outputs(246));
    outputs(402) <= layer2_outputs(376);
    outputs(403) <= (layer2_outputs(804)) and (layer2_outputs(1444));
    outputs(404) <= (layer2_outputs(2003)) and not (layer2_outputs(1490));
    outputs(405) <= not((layer2_outputs(284)) or (layer2_outputs(1504)));
    outputs(406) <= (layer2_outputs(2113)) and not (layer2_outputs(2092));
    outputs(407) <= not((layer2_outputs(162)) or (layer2_outputs(733)));
    outputs(408) <= (layer2_outputs(2475)) xor (layer2_outputs(1037));
    outputs(409) <= not((layer2_outputs(273)) or (layer2_outputs(1540)));
    outputs(410) <= (layer2_outputs(1331)) and not (layer2_outputs(2213));
    outputs(411) <= not((layer2_outputs(1572)) or (layer2_outputs(1392)));
    outputs(412) <= layer2_outputs(1558);
    outputs(413) <= not(layer2_outputs(830));
    outputs(414) <= (layer2_outputs(240)) and (layer2_outputs(1258));
    outputs(415) <= not(layer2_outputs(2542));
    outputs(416) <= (layer2_outputs(269)) and (layer2_outputs(811));
    outputs(417) <= not(layer2_outputs(2314));
    outputs(418) <= (layer2_outputs(2118)) and not (layer2_outputs(1512));
    outputs(419) <= not((layer2_outputs(2548)) or (layer2_outputs(1203)));
    outputs(420) <= (layer2_outputs(301)) and (layer2_outputs(1620));
    outputs(421) <= (layer2_outputs(967)) and not (layer2_outputs(2154));
    outputs(422) <= (layer2_outputs(1232)) and (layer2_outputs(268));
    outputs(423) <= (layer2_outputs(2167)) or (layer2_outputs(1717));
    outputs(424) <= not(layer2_outputs(1870));
    outputs(425) <= not(layer2_outputs(364));
    outputs(426) <= (layer2_outputs(197)) and (layer2_outputs(647));
    outputs(427) <= (layer2_outputs(1642)) or (layer2_outputs(1248));
    outputs(428) <= (layer2_outputs(1622)) and not (layer2_outputs(487));
    outputs(429) <= layer2_outputs(2491);
    outputs(430) <= layer2_outputs(549);
    outputs(431) <= not((layer2_outputs(1609)) or (layer2_outputs(832)));
    outputs(432) <= layer2_outputs(216);
    outputs(433) <= not((layer2_outputs(1282)) or (layer2_outputs(1654)));
    outputs(434) <= not(layer2_outputs(79));
    outputs(435) <= not((layer2_outputs(1855)) or (layer2_outputs(538)));
    outputs(436) <= not((layer2_outputs(1131)) or (layer2_outputs(2)));
    outputs(437) <= not(layer2_outputs(1056));
    outputs(438) <= not((layer2_outputs(2348)) or (layer2_outputs(1391)));
    outputs(439) <= (layer2_outputs(593)) and not (layer2_outputs(1242));
    outputs(440) <= (layer2_outputs(1253)) and (layer2_outputs(1903));
    outputs(441) <= layer2_outputs(2097);
    outputs(442) <= (layer2_outputs(2335)) and not (layer2_outputs(1723));
    outputs(443) <= not(layer2_outputs(1679));
    outputs(444) <= (layer2_outputs(1615)) xor (layer2_outputs(356));
    outputs(445) <= (layer2_outputs(88)) and not (layer2_outputs(2334));
    outputs(446) <= (layer2_outputs(277)) xor (layer2_outputs(516));
    outputs(447) <= not((layer2_outputs(1015)) xor (layer2_outputs(1020)));
    outputs(448) <= (layer2_outputs(907)) and (layer2_outputs(1890));
    outputs(449) <= layer2_outputs(1305);
    outputs(450) <= layer2_outputs(717);
    outputs(451) <= layer2_outputs(1066);
    outputs(452) <= layer2_outputs(134);
    outputs(453) <= layer2_outputs(2216);
    outputs(454) <= not(layer2_outputs(1271));
    outputs(455) <= layer2_outputs(727);
    outputs(456) <= not(layer2_outputs(2512));
    outputs(457) <= not((layer2_outputs(1945)) or (layer2_outputs(264)));
    outputs(458) <= not((layer2_outputs(715)) or (layer2_outputs(2207)));
    outputs(459) <= not((layer2_outputs(944)) and (layer2_outputs(2536)));
    outputs(460) <= layer2_outputs(1290);
    outputs(461) <= (layer2_outputs(807)) and not (layer2_outputs(1217));
    outputs(462) <= not(layer2_outputs(1045));
    outputs(463) <= not((layer2_outputs(1794)) or (layer2_outputs(2483)));
    outputs(464) <= not(layer2_outputs(1734));
    outputs(465) <= not(layer2_outputs(480));
    outputs(466) <= not(layer2_outputs(2222));
    outputs(467) <= layer2_outputs(2247);
    outputs(468) <= layer2_outputs(2070);
    outputs(469) <= (layer2_outputs(1245)) and (layer2_outputs(736));
    outputs(470) <= layer2_outputs(134);
    outputs(471) <= not(layer2_outputs(2185));
    outputs(472) <= (layer2_outputs(819)) and not (layer2_outputs(90));
    outputs(473) <= layer2_outputs(1758);
    outputs(474) <= not(layer2_outputs(1200));
    outputs(475) <= not((layer2_outputs(550)) or (layer2_outputs(189)));
    outputs(476) <= not((layer2_outputs(2184)) or (layer2_outputs(1439)));
    outputs(477) <= (layer2_outputs(1021)) and not (layer2_outputs(188));
    outputs(478) <= not((layer2_outputs(256)) or (layer2_outputs(336)));
    outputs(479) <= (layer2_outputs(421)) and not (layer2_outputs(954));
    outputs(480) <= not(layer2_outputs(2059));
    outputs(481) <= not((layer2_outputs(788)) or (layer2_outputs(1251)));
    outputs(482) <= (layer2_outputs(1988)) and (layer2_outputs(62));
    outputs(483) <= not(layer2_outputs(688));
    outputs(484) <= not((layer2_outputs(1907)) or (layer2_outputs(992)));
    outputs(485) <= not((layer2_outputs(1337)) or (layer2_outputs(1391)));
    outputs(486) <= not(layer2_outputs(664));
    outputs(487) <= not((layer2_outputs(2487)) or (layer2_outputs(343)));
    outputs(488) <= not((layer2_outputs(1911)) or (layer2_outputs(729)));
    outputs(489) <= (layer2_outputs(700)) and not (layer2_outputs(393));
    outputs(490) <= not(layer2_outputs(949));
    outputs(491) <= not((layer2_outputs(2179)) xor (layer2_outputs(1534)));
    outputs(492) <= not(layer2_outputs(1144));
    outputs(493) <= (layer2_outputs(114)) and (layer2_outputs(690));
    outputs(494) <= (layer2_outputs(764)) and not (layer2_outputs(1334));
    outputs(495) <= (layer2_outputs(1151)) and not (layer2_outputs(1489));
    outputs(496) <= (layer2_outputs(1995)) and not (layer2_outputs(429));
    outputs(497) <= not(layer2_outputs(152));
    outputs(498) <= not(layer2_outputs(2082));
    outputs(499) <= not(layer2_outputs(1790)) or (layer2_outputs(1759));
    outputs(500) <= (layer2_outputs(2381)) and (layer2_outputs(456));
    outputs(501) <= (layer2_outputs(2510)) and not (layer2_outputs(283));
    outputs(502) <= (layer2_outputs(1396)) and not (layer2_outputs(2112));
    outputs(503) <= layer2_outputs(634);
    outputs(504) <= not((layer2_outputs(966)) xor (layer2_outputs(669)));
    outputs(505) <= layer2_outputs(1728);
    outputs(506) <= layer2_outputs(2258);
    outputs(507) <= not(layer2_outputs(2212));
    outputs(508) <= (layer2_outputs(2511)) and not (layer2_outputs(2066));
    outputs(509) <= (layer2_outputs(249)) xor (layer2_outputs(1115));
    outputs(510) <= not(layer2_outputs(170));
    outputs(511) <= layer2_outputs(1740);
    outputs(512) <= not(layer2_outputs(1116));
    outputs(513) <= not(layer2_outputs(735));
    outputs(514) <= not((layer2_outputs(46)) or (layer2_outputs(1210)));
    outputs(515) <= (layer2_outputs(1333)) xor (layer2_outputs(904));
    outputs(516) <= not(layer2_outputs(2161));
    outputs(517) <= not(layer2_outputs(514));
    outputs(518) <= not(layer2_outputs(1409));
    outputs(519) <= not(layer2_outputs(1997));
    outputs(520) <= layer2_outputs(1315);
    outputs(521) <= layer2_outputs(837);
    outputs(522) <= (layer2_outputs(2240)) and not (layer2_outputs(797));
    outputs(523) <= (layer2_outputs(1566)) xor (layer2_outputs(2401));
    outputs(524) <= (layer2_outputs(1067)) and not (layer2_outputs(1984));
    outputs(525) <= layer2_outputs(475);
    outputs(526) <= (layer2_outputs(1618)) and not (layer2_outputs(555));
    outputs(527) <= not(layer2_outputs(314));
    outputs(528) <= not(layer2_outputs(1029));
    outputs(529) <= (layer2_outputs(136)) or (layer2_outputs(1698));
    outputs(530) <= not(layer2_outputs(1344));
    outputs(531) <= (layer2_outputs(318)) and not (layer2_outputs(1109));
    outputs(532) <= layer2_outputs(523);
    outputs(533) <= (layer2_outputs(250)) and (layer2_outputs(2442));
    outputs(534) <= layer2_outputs(586);
    outputs(535) <= (layer2_outputs(876)) xor (layer2_outputs(759));
    outputs(536) <= not(layer2_outputs(1674));
    outputs(537) <= layer2_outputs(1692);
    outputs(538) <= layer2_outputs(674);
    outputs(539) <= (layer2_outputs(1966)) and (layer2_outputs(2203));
    outputs(540) <= not(layer2_outputs(504));
    outputs(541) <= (layer2_outputs(852)) xor (layer2_outputs(2355));
    outputs(542) <= (layer2_outputs(184)) xor (layer2_outputs(568));
    outputs(543) <= layer2_outputs(874);
    outputs(544) <= (layer2_outputs(2193)) and not (layer2_outputs(696));
    outputs(545) <= (layer2_outputs(2310)) and not (layer2_outputs(505));
    outputs(546) <= (layer2_outputs(2281)) and (layer2_outputs(866));
    outputs(547) <= not(layer2_outputs(1093));
    outputs(548) <= (layer2_outputs(1169)) and not (layer2_outputs(740));
    outputs(549) <= not((layer2_outputs(1400)) and (layer2_outputs(182)));
    outputs(550) <= not((layer2_outputs(1705)) xor (layer2_outputs(159)));
    outputs(551) <= (layer2_outputs(2153)) and not (layer2_outputs(706));
    outputs(552) <= (layer2_outputs(1376)) and not (layer2_outputs(2303));
    outputs(553) <= not(layer2_outputs(1839)) or (layer2_outputs(968));
    outputs(554) <= not((layer2_outputs(792)) xor (layer2_outputs(2386)));
    outputs(555) <= layer2_outputs(265);
    outputs(556) <= not(layer2_outputs(2123));
    outputs(557) <= not(layer2_outputs(389));
    outputs(558) <= not(layer2_outputs(86));
    outputs(559) <= not((layer2_outputs(123)) and (layer2_outputs(684)));
    outputs(560) <= (layer2_outputs(1819)) and not (layer2_outputs(1570));
    outputs(561) <= (layer2_outputs(1357)) and not (layer2_outputs(2052));
    outputs(562) <= not((layer2_outputs(2200)) xor (layer2_outputs(1917)));
    outputs(563) <= not(layer2_outputs(979));
    outputs(564) <= (layer2_outputs(1375)) and not (layer2_outputs(1134));
    outputs(565) <= not((layer2_outputs(252)) and (layer2_outputs(873)));
    outputs(566) <= not(layer2_outputs(1801));
    outputs(567) <= (layer2_outputs(1877)) and (layer2_outputs(1960));
    outputs(568) <= (layer2_outputs(1710)) or (layer2_outputs(2490));
    outputs(569) <= layer2_outputs(1233);
    outputs(570) <= not((layer2_outputs(373)) or (layer2_outputs(668)));
    outputs(571) <= layer2_outputs(747);
    outputs(572) <= not(layer2_outputs(2456));
    outputs(573) <= not((layer2_outputs(605)) xor (layer2_outputs(105)));
    outputs(574) <= layer2_outputs(1527);
    outputs(575) <= (layer2_outputs(1033)) or (layer2_outputs(2358));
    outputs(576) <= layer2_outputs(515);
    outputs(577) <= (layer2_outputs(231)) and not (layer2_outputs(161));
    outputs(578) <= (layer2_outputs(862)) and not (layer2_outputs(742));
    outputs(579) <= not(layer2_outputs(124));
    outputs(580) <= layer2_outputs(1396);
    outputs(581) <= not(layer2_outputs(1709)) or (layer2_outputs(2030));
    outputs(582) <= (layer2_outputs(2299)) or (layer2_outputs(2020));
    outputs(583) <= not(layer2_outputs(2390));
    outputs(584) <= not((layer2_outputs(1926)) xor (layer2_outputs(1778)));
    outputs(585) <= not((layer2_outputs(608)) or (layer2_outputs(2044)));
    outputs(586) <= not(layer2_outputs(689));
    outputs(587) <= (layer2_outputs(2360)) or (layer2_outputs(173));
    outputs(588) <= not((layer2_outputs(1766)) xor (layer2_outputs(906)));
    outputs(589) <= not((layer2_outputs(1871)) and (layer2_outputs(1189)));
    outputs(590) <= (layer2_outputs(1050)) or (layer2_outputs(998));
    outputs(591) <= not(layer2_outputs(1125)) or (layer2_outputs(803));
    outputs(592) <= layer2_outputs(1963);
    outputs(593) <= not(layer2_outputs(2270));
    outputs(594) <= not(layer2_outputs(1448));
    outputs(595) <= layer2_outputs(1438);
    outputs(596) <= layer2_outputs(749);
    outputs(597) <= not((layer2_outputs(298)) xor (layer2_outputs(2331)));
    outputs(598) <= (layer2_outputs(2548)) and (layer2_outputs(2164));
    outputs(599) <= not(layer2_outputs(2485));
    outputs(600) <= layer2_outputs(1009);
    outputs(601) <= (layer2_outputs(1193)) or (layer2_outputs(2420));
    outputs(602) <= not((layer2_outputs(26)) xor (layer2_outputs(1120)));
    outputs(603) <= not(layer2_outputs(89));
    outputs(604) <= not(layer2_outputs(1754));
    outputs(605) <= not(layer2_outputs(156));
    outputs(606) <= layer2_outputs(1910);
    outputs(607) <= layer2_outputs(499);
    outputs(608) <= not(layer2_outputs(812));
    outputs(609) <= not(layer2_outputs(1336)) or (layer2_outputs(656));
    outputs(610) <= layer2_outputs(1152);
    outputs(611) <= not(layer2_outputs(791));
    outputs(612) <= not((layer2_outputs(377)) or (layer2_outputs(2491)));
    outputs(613) <= not(layer2_outputs(92));
    outputs(614) <= (layer2_outputs(2239)) or (layer2_outputs(1193));
    outputs(615) <= layer2_outputs(204);
    outputs(616) <= layer2_outputs(874);
    outputs(617) <= (layer2_outputs(927)) xor (layer2_outputs(458));
    outputs(618) <= not(layer2_outputs(715));
    outputs(619) <= layer2_outputs(2398);
    outputs(620) <= not((layer2_outputs(610)) or (layer2_outputs(1813)));
    outputs(621) <= layer2_outputs(879);
    outputs(622) <= layer2_outputs(966);
    outputs(623) <= layer2_outputs(557);
    outputs(624) <= layer2_outputs(613);
    outputs(625) <= not((layer2_outputs(1674)) or (layer2_outputs(522)));
    outputs(626) <= layer2_outputs(77);
    outputs(627) <= (layer2_outputs(1856)) and not (layer2_outputs(38));
    outputs(628) <= not(layer2_outputs(2162));
    outputs(629) <= not((layer2_outputs(580)) and (layer2_outputs(1331)));
    outputs(630) <= not(layer2_outputs(1578));
    outputs(631) <= (layer2_outputs(1043)) and (layer2_outputs(114));
    outputs(632) <= not(layer2_outputs(2075));
    outputs(633) <= not(layer2_outputs(882));
    outputs(634) <= layer2_outputs(2552);
    outputs(635) <= (layer2_outputs(274)) and (layer2_outputs(231));
    outputs(636) <= not(layer2_outputs(1885)) or (layer2_outputs(1696));
    outputs(637) <= not((layer2_outputs(2391)) or (layer2_outputs(313)));
    outputs(638) <= not(layer2_outputs(455));
    outputs(639) <= layer2_outputs(1010);
    outputs(640) <= (layer2_outputs(1131)) or (layer2_outputs(849));
    outputs(641) <= not(layer2_outputs(270));
    outputs(642) <= (layer2_outputs(422)) and not (layer2_outputs(637));
    outputs(643) <= (layer2_outputs(819)) and not (layer2_outputs(1691));
    outputs(644) <= not(layer2_outputs(1874));
    outputs(645) <= (layer2_outputs(1107)) and (layer2_outputs(1989));
    outputs(646) <= not(layer2_outputs(731));
    outputs(647) <= (layer2_outputs(617)) and (layer2_outputs(318));
    outputs(648) <= (layer2_outputs(2312)) and (layer2_outputs(2160));
    outputs(649) <= layer2_outputs(1166);
    outputs(650) <= not(layer2_outputs(555));
    outputs(651) <= not(layer2_outputs(317));
    outputs(652) <= layer2_outputs(1303);
    outputs(653) <= layer2_outputs(976);
    outputs(654) <= (layer2_outputs(2149)) xor (layer2_outputs(2459));
    outputs(655) <= (layer2_outputs(2204)) and not (layer2_outputs(1737));
    outputs(656) <= not(layer2_outputs(1018)) or (layer2_outputs(1757));
    outputs(657) <= not(layer2_outputs(1854));
    outputs(658) <= layer2_outputs(2026);
    outputs(659) <= not((layer2_outputs(1330)) xor (layer2_outputs(1742)));
    outputs(660) <= not(layer2_outputs(1330));
    outputs(661) <= (layer2_outputs(1438)) and not (layer2_outputs(717));
    outputs(662) <= layer2_outputs(312);
    outputs(663) <= not(layer2_outputs(696));
    outputs(664) <= (layer2_outputs(707)) or (layer2_outputs(1256));
    outputs(665) <= layer2_outputs(962);
    outputs(666) <= layer2_outputs(1884);
    outputs(667) <= not((layer2_outputs(1846)) xor (layer2_outputs(563)));
    outputs(668) <= not(layer2_outputs(124)) or (layer2_outputs(1282));
    outputs(669) <= (layer2_outputs(2526)) and (layer2_outputs(302));
    outputs(670) <= (layer2_outputs(1525)) xor (layer2_outputs(388));
    outputs(671) <= (layer2_outputs(300)) or (layer2_outputs(2382));
    outputs(672) <= layer2_outputs(1830);
    outputs(673) <= not((layer2_outputs(463)) and (layer2_outputs(2384)));
    outputs(674) <= layer2_outputs(433);
    outputs(675) <= not(layer2_outputs(237));
    outputs(676) <= layer2_outputs(1597);
    outputs(677) <= not((layer2_outputs(459)) xor (layer2_outputs(2518)));
    outputs(678) <= not(layer2_outputs(812)) or (layer2_outputs(1773));
    outputs(679) <= not(layer2_outputs(2338));
    outputs(680) <= not(layer2_outputs(1550));
    outputs(681) <= not(layer2_outputs(834));
    outputs(682) <= (layer2_outputs(926)) and not (layer2_outputs(1389));
    outputs(683) <= not(layer2_outputs(107));
    outputs(684) <= (layer2_outputs(613)) and (layer2_outputs(569));
    outputs(685) <= (layer2_outputs(2441)) and not (layer2_outputs(991));
    outputs(686) <= not((layer2_outputs(1641)) xor (layer2_outputs(2383)));
    outputs(687) <= (layer2_outputs(2537)) and not (layer2_outputs(2531));
    outputs(688) <= not(layer2_outputs(1590));
    outputs(689) <= (layer2_outputs(2190)) and (layer2_outputs(2045));
    outputs(690) <= layer2_outputs(1745);
    outputs(691) <= not((layer2_outputs(1603)) and (layer2_outputs(1729)));
    outputs(692) <= (layer2_outputs(620)) and (layer2_outputs(552));
    outputs(693) <= layer2_outputs(1118);
    outputs(694) <= layer2_outputs(1666);
    outputs(695) <= not((layer2_outputs(583)) and (layer2_outputs(228)));
    outputs(696) <= not(layer2_outputs(1967));
    outputs(697) <= (layer2_outputs(870)) and not (layer2_outputs(1874));
    outputs(698) <= not(layer2_outputs(583));
    outputs(699) <= not((layer2_outputs(1075)) and (layer2_outputs(2372)));
    outputs(700) <= layer2_outputs(1568);
    outputs(701) <= not((layer2_outputs(2307)) and (layer2_outputs(2531)));
    outputs(702) <= not(layer2_outputs(44)) or (layer2_outputs(502));
    outputs(703) <= not(layer2_outputs(974));
    outputs(704) <= not(layer2_outputs(2294));
    outputs(705) <= not((layer2_outputs(2351)) or (layer2_outputs(973)));
    outputs(706) <= not(layer2_outputs(1543));
    outputs(707) <= not((layer2_outputs(2485)) or (layer2_outputs(30)));
    outputs(708) <= not(layer2_outputs(303));
    outputs(709) <= (layer2_outputs(1038)) and (layer2_outputs(2356));
    outputs(710) <= layer2_outputs(1394);
    outputs(711) <= layer2_outputs(1755);
    outputs(712) <= not(layer2_outputs(2379));
    outputs(713) <= (layer2_outputs(535)) and not (layer2_outputs(745));
    outputs(714) <= not(layer2_outputs(493));
    outputs(715) <= layer2_outputs(1756);
    outputs(716) <= (layer2_outputs(412)) and (layer2_outputs(802));
    outputs(717) <= layer2_outputs(532);
    outputs(718) <= not(layer2_outputs(581));
    outputs(719) <= not(layer2_outputs(1295));
    outputs(720) <= not(layer2_outputs(2025));
    outputs(721) <= not(layer2_outputs(1013));
    outputs(722) <= (layer2_outputs(798)) or (layer2_outputs(721));
    outputs(723) <= layer2_outputs(102);
    outputs(724) <= (layer2_outputs(1149)) xor (layer2_outputs(2371));
    outputs(725) <= not(layer2_outputs(2324));
    outputs(726) <= (layer2_outputs(2449)) and not (layer2_outputs(2513));
    outputs(727) <= layer2_outputs(1233);
    outputs(728) <= layer2_outputs(68);
    outputs(729) <= (layer2_outputs(1856)) or (layer2_outputs(2191));
    outputs(730) <= not((layer2_outputs(1056)) xor (layer2_outputs(814)));
    outputs(731) <= not(layer2_outputs(1288));
    outputs(732) <= (layer2_outputs(155)) xor (layer2_outputs(678));
    outputs(733) <= (layer2_outputs(1197)) xor (layer2_outputs(1730));
    outputs(734) <= layer2_outputs(1585);
    outputs(735) <= layer2_outputs(2191);
    outputs(736) <= not(layer2_outputs(1482));
    outputs(737) <= not((layer2_outputs(570)) and (layer2_outputs(1448)));
    outputs(738) <= not(layer2_outputs(2105));
    outputs(739) <= (layer2_outputs(760)) and (layer2_outputs(1966));
    outputs(740) <= not((layer2_outputs(2141)) and (layer2_outputs(1090)));
    outputs(741) <= layer2_outputs(1216);
    outputs(742) <= not(layer2_outputs(1831)) or (layer2_outputs(1204));
    outputs(743) <= not((layer2_outputs(1069)) or (layer2_outputs(1482)));
    outputs(744) <= not(layer2_outputs(2178)) or (layer2_outputs(1954));
    outputs(745) <= layer2_outputs(560);
    outputs(746) <= layer2_outputs(1145);
    outputs(747) <= layer2_outputs(1962);
    outputs(748) <= (layer2_outputs(28)) xor (layer2_outputs(1471));
    outputs(749) <= (layer2_outputs(743)) and not (layer2_outputs(1024));
    outputs(750) <= layer2_outputs(140);
    outputs(751) <= not(layer2_outputs(774));
    outputs(752) <= layer2_outputs(2496);
    outputs(753) <= not(layer2_outputs(1379));
    outputs(754) <= (layer2_outputs(498)) and not (layer2_outputs(2509));
    outputs(755) <= (layer2_outputs(21)) and not (layer2_outputs(2169));
    outputs(756) <= layer2_outputs(49);
    outputs(757) <= layer2_outputs(612);
    outputs(758) <= not((layer2_outputs(1907)) or (layer2_outputs(1501)));
    outputs(759) <= not(layer2_outputs(238));
    outputs(760) <= (layer2_outputs(1236)) and (layer2_outputs(1956));
    outputs(761) <= layer2_outputs(140);
    outputs(762) <= not(layer2_outputs(834));
    outputs(763) <= not(layer2_outputs(2543));
    outputs(764) <= layer2_outputs(763);
    outputs(765) <= layer2_outputs(1969);
    outputs(766) <= not(layer2_outputs(85)) or (layer2_outputs(582));
    outputs(767) <= layer2_outputs(325);
    outputs(768) <= not(layer2_outputs(1625));
    outputs(769) <= not(layer2_outputs(343));
    outputs(770) <= not(layer2_outputs(1146));
    outputs(771) <= not(layer2_outputs(214));
    outputs(772) <= not(layer2_outputs(2217));
    outputs(773) <= layer2_outputs(2472);
    outputs(774) <= not((layer2_outputs(628)) xor (layer2_outputs(1743)));
    outputs(775) <= layer2_outputs(193);
    outputs(776) <= (layer2_outputs(605)) and (layer2_outputs(1236));
    outputs(777) <= not((layer2_outputs(2370)) or (layer2_outputs(2428)));
    outputs(778) <= not((layer2_outputs(2037)) or (layer2_outputs(2261)));
    outputs(779) <= not((layer2_outputs(1243)) or (layer2_outputs(2005)));
    outputs(780) <= (layer2_outputs(660)) and not (layer2_outputs(2028));
    outputs(781) <= (layer2_outputs(122)) and not (layer2_outputs(202));
    outputs(782) <= not((layer2_outputs(1435)) or (layer2_outputs(2022)));
    outputs(783) <= (layer2_outputs(818)) and (layer2_outputs(2234));
    outputs(784) <= layer2_outputs(693);
    outputs(785) <= not((layer2_outputs(942)) or (layer2_outputs(384)));
    outputs(786) <= layer2_outputs(1180);
    outputs(787) <= not(layer2_outputs(909));
    outputs(788) <= (layer2_outputs(1476)) and (layer2_outputs(2053));
    outputs(789) <= (layer2_outputs(2196)) or (layer2_outputs(162));
    outputs(790) <= not((layer2_outputs(1369)) xor (layer2_outputs(476)));
    outputs(791) <= layer2_outputs(833);
    outputs(792) <= (layer2_outputs(328)) and not (layer2_outputs(1710));
    outputs(793) <= layer2_outputs(2018);
    outputs(794) <= layer2_outputs(1584);
    outputs(795) <= layer2_outputs(1970);
    outputs(796) <= not((layer2_outputs(1486)) or (layer2_outputs(2342)));
    outputs(797) <= (layer2_outputs(449)) and not (layer2_outputs(2153));
    outputs(798) <= layer2_outputs(1522);
    outputs(799) <= layer2_outputs(1697);
    outputs(800) <= (layer2_outputs(113)) and (layer2_outputs(1586));
    outputs(801) <= not(layer2_outputs(1843));
    outputs(802) <= (layer2_outputs(1194)) and not (layer2_outputs(2502));
    outputs(803) <= not(layer2_outputs(319));
    outputs(804) <= layer2_outputs(447);
    outputs(805) <= layer2_outputs(2532);
    outputs(806) <= not((layer2_outputs(998)) xor (layer2_outputs(519)));
    outputs(807) <= layer2_outputs(1941);
    outputs(808) <= layer2_outputs(1783);
    outputs(809) <= (layer2_outputs(1646)) and not (layer2_outputs(1168));
    outputs(810) <= layer2_outputs(922);
    outputs(811) <= layer2_outputs(2413);
    outputs(812) <= not(layer2_outputs(1467)) or (layer2_outputs(2187));
    outputs(813) <= layer2_outputs(435);
    outputs(814) <= not((layer2_outputs(494)) xor (layer2_outputs(1026)));
    outputs(815) <= (layer2_outputs(1537)) and not (layer2_outputs(1909));
    outputs(816) <= layer2_outputs(169);
    outputs(817) <= not(layer2_outputs(2168));
    outputs(818) <= not(layer2_outputs(170));
    outputs(819) <= layer2_outputs(2228);
    outputs(820) <= (layer2_outputs(596)) xor (layer2_outputs(1242));
    outputs(821) <= not(layer2_outputs(203));
    outputs(822) <= not((layer2_outputs(400)) or (layer2_outputs(958)));
    outputs(823) <= not(layer2_outputs(446));
    outputs(824) <= (layer2_outputs(720)) and not (layer2_outputs(2367));
    outputs(825) <= (layer2_outputs(1258)) xor (layer2_outputs(2393));
    outputs(826) <= not(layer2_outputs(773)) or (layer2_outputs(1460));
    outputs(827) <= not(layer2_outputs(261));
    outputs(828) <= layer2_outputs(1036);
    outputs(829) <= (layer2_outputs(1971)) and not (layer2_outputs(871));
    outputs(830) <= not(layer2_outputs(2332));
    outputs(831) <= layer2_outputs(1665);
    outputs(832) <= not(layer2_outputs(2448));
    outputs(833) <= not(layer2_outputs(764));
    outputs(834) <= layer2_outputs(910);
    outputs(835) <= not((layer2_outputs(69)) or (layer2_outputs(59)));
    outputs(836) <= layer2_outputs(2233);
    outputs(837) <= layer2_outputs(680);
    outputs(838) <= (layer2_outputs(195)) and (layer2_outputs(1044));
    outputs(839) <= (layer2_outputs(698)) and (layer2_outputs(2489));
    outputs(840) <= not((layer2_outputs(1320)) and (layer2_outputs(463)));
    outputs(841) <= (layer2_outputs(2016)) and not (layer2_outputs(0));
    outputs(842) <= (layer2_outputs(2225)) and not (layer2_outputs(2122));
    outputs(843) <= layer2_outputs(1829);
    outputs(844) <= not(layer2_outputs(1318));
    outputs(845) <= not((layer2_outputs(2289)) or (layer2_outputs(1717)));
    outputs(846) <= (layer2_outputs(1887)) and not (layer2_outputs(25));
    outputs(847) <= layer2_outputs(1882);
    outputs(848) <= not(layer2_outputs(143));
    outputs(849) <= layer2_outputs(2403);
    outputs(850) <= layer2_outputs(1783);
    outputs(851) <= (layer2_outputs(1979)) and (layer2_outputs(1368));
    outputs(852) <= (layer2_outputs(18)) and not (layer2_outputs(535));
    outputs(853) <= not(layer2_outputs(150));
    outputs(854) <= not((layer2_outputs(121)) or (layer2_outputs(737)));
    outputs(855) <= (layer2_outputs(2206)) xor (layer2_outputs(156));
    outputs(856) <= (layer2_outputs(531)) and not (layer2_outputs(150));
    outputs(857) <= not(layer2_outputs(2384));
    outputs(858) <= (layer2_outputs(694)) and (layer2_outputs(2155));
    outputs(859) <= (layer2_outputs(843)) and not (layer2_outputs(893));
    outputs(860) <= not(layer2_outputs(292));
    outputs(861) <= layer2_outputs(673);
    outputs(862) <= layer2_outputs(308);
    outputs(863) <= not(layer2_outputs(2009));
    outputs(864) <= (layer2_outputs(141)) and (layer2_outputs(131));
    outputs(865) <= not((layer2_outputs(788)) or (layer2_outputs(1541)));
    outputs(866) <= (layer2_outputs(2151)) and (layer2_outputs(1968));
    outputs(867) <= layer2_outputs(215);
    outputs(868) <= layer2_outputs(789);
    outputs(869) <= (layer2_outputs(1086)) and (layer2_outputs(1927));
    outputs(870) <= (layer2_outputs(859)) and not (layer2_outputs(453));
    outputs(871) <= (layer2_outputs(1769)) xor (layer2_outputs(458));
    outputs(872) <= (layer2_outputs(524)) and not (layer2_outputs(1902));
    outputs(873) <= not(layer2_outputs(1983)) or (layer2_outputs(939));
    outputs(874) <= not((layer2_outputs(661)) xor (layer2_outputs(1656)));
    outputs(875) <= not(layer2_outputs(1390));
    outputs(876) <= (layer2_outputs(2266)) and (layer2_outputs(944));
    outputs(877) <= (layer2_outputs(965)) and (layer2_outputs(1957));
    outputs(878) <= layer2_outputs(1609);
    outputs(879) <= not(layer2_outputs(2546));
    outputs(880) <= not((layer2_outputs(1748)) or (layer2_outputs(1810)));
    outputs(881) <= (layer2_outputs(1602)) and (layer2_outputs(1000));
    outputs(882) <= not((layer2_outputs(820)) or (layer2_outputs(403)));
    outputs(883) <= not((layer2_outputs(180)) or (layer2_outputs(71)));
    outputs(884) <= layer2_outputs(222);
    outputs(885) <= layer2_outputs(1858);
    outputs(886) <= (layer2_outputs(2515)) and not (layer2_outputs(1991));
    outputs(887) <= (layer2_outputs(1259)) and (layer2_outputs(2286));
    outputs(888) <= layer2_outputs(734);
    outputs(889) <= not(layer2_outputs(1478));
    outputs(890) <= not(layer2_outputs(2375));
    outputs(891) <= (layer2_outputs(1397)) and not (layer2_outputs(1133));
    outputs(892) <= (layer2_outputs(1807)) and not (layer2_outputs(1539));
    outputs(893) <= layer2_outputs(2230);
    outputs(894) <= layer2_outputs(2406);
    outputs(895) <= (layer2_outputs(2492)) and (layer2_outputs(712));
    outputs(896) <= (layer2_outputs(1889)) and not (layer2_outputs(2041));
    outputs(897) <= layer2_outputs(616);
    outputs(898) <= not((layer2_outputs(1492)) or (layer2_outputs(2288)));
    outputs(899) <= not(layer2_outputs(1061));
    outputs(900) <= (layer2_outputs(1239)) and (layer2_outputs(1931));
    outputs(901) <= not((layer2_outputs(2276)) or (layer2_outputs(1866)));
    outputs(902) <= layer2_outputs(890);
    outputs(903) <= layer2_outputs(2446);
    outputs(904) <= (layer2_outputs(1903)) and not (layer2_outputs(488));
    outputs(905) <= not(layer2_outputs(1896));
    outputs(906) <= not(layer2_outputs(2289));
    outputs(907) <= (layer2_outputs(2140)) and (layer2_outputs(1829));
    outputs(908) <= (layer2_outputs(868)) and not (layer2_outputs(250));
    outputs(909) <= (layer2_outputs(1151)) and (layer2_outputs(857));
    outputs(910) <= not((layer2_outputs(2502)) xor (layer2_outputs(1953)));
    outputs(911) <= layer2_outputs(2397);
    outputs(912) <= not(layer2_outputs(2353));
    outputs(913) <= layer2_outputs(2175);
    outputs(914) <= layer2_outputs(1183);
    outputs(915) <= not(layer2_outputs(138));
    outputs(916) <= not((layer2_outputs(2361)) or (layer2_outputs(489)));
    outputs(917) <= (layer2_outputs(750)) and not (layer2_outputs(736));
    outputs(918) <= (layer2_outputs(387)) or (layer2_outputs(1349));
    outputs(919) <= layer2_outputs(1530);
    outputs(920) <= (layer2_outputs(1882)) and not (layer2_outputs(1217));
    outputs(921) <= layer2_outputs(1458);
    outputs(922) <= not(layer2_outputs(348));
    outputs(923) <= not((layer2_outputs(1004)) xor (layer2_outputs(2523)));
    outputs(924) <= (layer2_outputs(1867)) and not (layer2_outputs(1564));
    outputs(925) <= not(layer2_outputs(1671)) or (layer2_outputs(1184));
    outputs(926) <= not(layer2_outputs(84));
    outputs(927) <= layer2_outputs(1388);
    outputs(928) <= layer2_outputs(1785);
    outputs(929) <= not(layer2_outputs(2279));
    outputs(930) <= (layer2_outputs(2351)) and not (layer2_outputs(135));
    outputs(931) <= not(layer2_outputs(920));
    outputs(932) <= layer2_outputs(151);
    outputs(933) <= not(layer2_outputs(1082));
    outputs(934) <= (layer2_outputs(118)) and not (layer2_outputs(319));
    outputs(935) <= not(layer2_outputs(60));
    outputs(936) <= not((layer2_outputs(1813)) or (layer2_outputs(842)));
    outputs(937) <= (layer2_outputs(205)) and not (layer2_outputs(4));
    outputs(938) <= layer2_outputs(1326);
    outputs(939) <= layer2_outputs(430);
    outputs(940) <= not(layer2_outputs(1604));
    outputs(941) <= not((layer2_outputs(332)) or (layer2_outputs(2104)));
    outputs(942) <= layer2_outputs(688);
    outputs(943) <= (layer2_outputs(1355)) and not (layer2_outputs(709));
    outputs(944) <= not(layer2_outputs(1419));
    outputs(945) <= not((layer2_outputs(401)) or (layer2_outputs(1073)));
    outputs(946) <= (layer2_outputs(791)) and not (layer2_outputs(919));
    outputs(947) <= not(layer2_outputs(1094));
    outputs(948) <= layer2_outputs(1977);
    outputs(949) <= not(layer2_outputs(2085));
    outputs(950) <= not(layer2_outputs(576));
    outputs(951) <= (layer2_outputs(17)) xor (layer2_outputs(2203));
    outputs(952) <= (layer2_outputs(779)) and (layer2_outputs(51));
    outputs(953) <= layer2_outputs(504);
    outputs(954) <= not(layer2_outputs(1390));
    outputs(955) <= not((layer2_outputs(198)) or (layer2_outputs(1793)));
    outputs(956) <= layer2_outputs(23);
    outputs(957) <= layer2_outputs(802);
    outputs(958) <= layer2_outputs(37);
    outputs(959) <= not(layer2_outputs(246));
    outputs(960) <= layer2_outputs(805);
    outputs(961) <= (layer2_outputs(1746)) and not (layer2_outputs(514));
    outputs(962) <= not(layer2_outputs(1857));
    outputs(963) <= layer2_outputs(2245);
    outputs(964) <= not(layer2_outputs(1462));
    outputs(965) <= (layer2_outputs(1184)) and not (layer2_outputs(357));
    outputs(966) <= not(layer2_outputs(2329));
    outputs(967) <= not((layer2_outputs(323)) or (layer2_outputs(2089)));
    outputs(968) <= not((layer2_outputs(2436)) or (layer2_outputs(705)));
    outputs(969) <= layer2_outputs(2115);
    outputs(970) <= not((layer2_outputs(1138)) xor (layer2_outputs(1346)));
    outputs(971) <= (layer2_outputs(2184)) or (layer2_outputs(2437));
    outputs(972) <= not(layer2_outputs(495));
    outputs(973) <= not(layer2_outputs(2373));
    outputs(974) <= not(layer2_outputs(1735)) or (layer2_outputs(664));
    outputs(975) <= (layer2_outputs(1670)) or (layer2_outputs(588));
    outputs(976) <= (layer2_outputs(1533)) xor (layer2_outputs(669));
    outputs(977) <= layer2_outputs(714);
    outputs(978) <= (layer2_outputs(1915)) and not (layer2_outputs(432));
    outputs(979) <= layer2_outputs(2225);
    outputs(980) <= (layer2_outputs(1519)) and (layer2_outputs(1939));
    outputs(981) <= (layer2_outputs(1463)) and (layer2_outputs(367));
    outputs(982) <= not(layer2_outputs(1701));
    outputs(983) <= layer2_outputs(863);
    outputs(984) <= (layer2_outputs(2482)) and not (layer2_outputs(1196));
    outputs(985) <= not((layer2_outputs(2192)) xor (layer2_outputs(1158)));
    outputs(986) <= not((layer2_outputs(2445)) or (layer2_outputs(813)));
    outputs(987) <= not(layer2_outputs(281));
    outputs(988) <= (layer2_outputs(2221)) xor (layer2_outputs(177));
    outputs(989) <= layer2_outputs(1823);
    outputs(990) <= (layer2_outputs(1594)) xor (layer2_outputs(1750));
    outputs(991) <= (layer2_outputs(2345)) xor (layer2_outputs(2080));
    outputs(992) <= layer2_outputs(2233);
    outputs(993) <= layer2_outputs(415);
    outputs(994) <= layer2_outputs(437);
    outputs(995) <= layer2_outputs(859);
    outputs(996) <= not((layer2_outputs(813)) and (layer2_outputs(1408)));
    outputs(997) <= (layer2_outputs(2411)) and not (layer2_outputs(1376));
    outputs(998) <= (layer2_outputs(2004)) and (layer2_outputs(1995));
    outputs(999) <= (layer2_outputs(1840)) and not (layer2_outputs(2457));
    outputs(1000) <= (layer2_outputs(2315)) and (layer2_outputs(1465));
    outputs(1001) <= layer2_outputs(2278);
    outputs(1002) <= layer2_outputs(757);
    outputs(1003) <= (layer2_outputs(1268)) and not (layer2_outputs(518));
    outputs(1004) <= layer2_outputs(687);
    outputs(1005) <= not(layer2_outputs(1792));
    outputs(1006) <= (layer2_outputs(571)) and not (layer2_outputs(1091));
    outputs(1007) <= not((layer2_outputs(276)) and (layer2_outputs(2311)));
    outputs(1008) <= layer2_outputs(1768);
    outputs(1009) <= not(layer2_outputs(1060));
    outputs(1010) <= (layer2_outputs(1051)) and not (layer2_outputs(1920));
    outputs(1011) <= layer2_outputs(424);
    outputs(1012) <= layer2_outputs(1582);
    outputs(1013) <= not(layer2_outputs(538));
    outputs(1014) <= (layer2_outputs(617)) and (layer2_outputs(863));
    outputs(1015) <= (layer2_outputs(757)) and not (layer2_outputs(2317));
    outputs(1016) <= not(layer2_outputs(855));
    outputs(1017) <= layer2_outputs(1888);
    outputs(1018) <= layer2_outputs(1083);
    outputs(1019) <= (layer2_outputs(997)) and (layer2_outputs(164));
    outputs(1020) <= layer2_outputs(2481);
    outputs(1021) <= layer2_outputs(398);
    outputs(1022) <= (layer2_outputs(2221)) and (layer2_outputs(594));
    outputs(1023) <= (layer2_outputs(1675)) and not (layer2_outputs(2195));
    outputs(1024) <= not((layer2_outputs(1395)) or (layer2_outputs(1703)));
    outputs(1025) <= not((layer2_outputs(1381)) or (layer2_outputs(1042)));
    outputs(1026) <= layer2_outputs(1012);
    outputs(1027) <= layer2_outputs(1496);
    outputs(1028) <= layer2_outputs(512);
    outputs(1029) <= not(layer2_outputs(27));
    outputs(1030) <= not(layer2_outputs(713));
    outputs(1031) <= (layer2_outputs(137)) and (layer2_outputs(2034));
    outputs(1032) <= layer2_outputs(1716);
    outputs(1033) <= not(layer2_outputs(937));
    outputs(1034) <= not(layer2_outputs(1972));
    outputs(1035) <= not((layer2_outputs(2235)) or (layer2_outputs(780)));
    outputs(1036) <= not(layer2_outputs(941));
    outputs(1037) <= not((layer2_outputs(1234)) or (layer2_outputs(1819)));
    outputs(1038) <= layer2_outputs(1377);
    outputs(1039) <= layer2_outputs(2533);
    outputs(1040) <= (layer2_outputs(1945)) and (layer2_outputs(700));
    outputs(1041) <= not((layer2_outputs(2088)) or (layer2_outputs(1214)));
    outputs(1042) <= not(layer2_outputs(416));
    outputs(1043) <= (layer2_outputs(2402)) and not (layer2_outputs(1912));
    outputs(1044) <= not((layer2_outputs(2403)) xor (layer2_outputs(805)));
    outputs(1045) <= (layer2_outputs(1386)) and not (layer2_outputs(131));
    outputs(1046) <= (layer2_outputs(2095)) and not (layer2_outputs(1485));
    outputs(1047) <= not(layer2_outputs(2558));
    outputs(1048) <= (layer2_outputs(845)) and (layer2_outputs(1262));
    outputs(1049) <= layer2_outputs(1047);
    outputs(1050) <= layer2_outputs(1967);
    outputs(1051) <= not(layer2_outputs(600));
    outputs(1052) <= not(layer2_outputs(330));
    outputs(1053) <= (layer2_outputs(1339)) or (layer2_outputs(488));
    outputs(1054) <= not(layer2_outputs(1031));
    outputs(1055) <= layer2_outputs(1195);
    outputs(1056) <= not(layer2_outputs(2427)) or (layer2_outputs(1892));
    outputs(1057) <= not(layer2_outputs(219));
    outputs(1058) <= not(layer2_outputs(2242));
    outputs(1059) <= (layer2_outputs(869)) and not (layer2_outputs(1457));
    outputs(1060) <= layer2_outputs(158);
    outputs(1061) <= (layer2_outputs(1836)) and not (layer2_outputs(109));
    outputs(1062) <= layer2_outputs(1449);
    outputs(1063) <= layer2_outputs(1163);
    outputs(1064) <= not((layer2_outputs(1655)) or (layer2_outputs(659)));
    outputs(1065) <= not((layer2_outputs(1153)) xor (layer2_outputs(1298)));
    outputs(1066) <= not((layer2_outputs(1273)) or (layer2_outputs(2120)));
    outputs(1067) <= layer2_outputs(139);
    outputs(1068) <= not(layer2_outputs(1077));
    outputs(1069) <= (layer2_outputs(1971)) and not (layer2_outputs(1044));
    outputs(1070) <= layer2_outputs(1001);
    outputs(1071) <= layer2_outputs(2493);
    outputs(1072) <= (layer2_outputs(211)) and (layer2_outputs(930));
    outputs(1073) <= not(layer2_outputs(1853));
    outputs(1074) <= (layer2_outputs(1167)) and not (layer2_outputs(1916));
    outputs(1075) <= layer2_outputs(2246);
    outputs(1076) <= not((layer2_outputs(656)) or (layer2_outputs(186)));
    outputs(1077) <= layer2_outputs(1407);
    outputs(1078) <= (layer2_outputs(1062)) and (layer2_outputs(1276));
    outputs(1079) <= not(layer2_outputs(730));
    outputs(1080) <= (layer2_outputs(599)) and (layer2_outputs(2096));
    outputs(1081) <= not(layer2_outputs(1308));
    outputs(1082) <= layer2_outputs(731);
    outputs(1083) <= not((layer2_outputs(562)) xor (layer2_outputs(1932)));
    outputs(1084) <= not(layer2_outputs(464)) or (layer2_outputs(841));
    outputs(1085) <= not(layer2_outputs(304));
    outputs(1086) <= not(layer2_outputs(2458)) or (layer2_outputs(1577));
    outputs(1087) <= layer2_outputs(2178);
    outputs(1088) <= not(layer2_outputs(2478));
    outputs(1089) <= layer2_outputs(1491);
    outputs(1090) <= layer2_outputs(2096);
    outputs(1091) <= layer2_outputs(53);
    outputs(1092) <= layer2_outputs(2332);
    outputs(1093) <= (layer2_outputs(770)) xor (layer2_outputs(208));
    outputs(1094) <= not(layer2_outputs(192)) or (layer2_outputs(466));
    outputs(1095) <= not((layer2_outputs(1696)) or (layer2_outputs(993)));
    outputs(1096) <= layer2_outputs(406);
    outputs(1097) <= not(layer2_outputs(1499));
    outputs(1098) <= not((layer2_outputs(1206)) or (layer2_outputs(355)));
    outputs(1099) <= not(layer2_outputs(330));
    outputs(1100) <= layer2_outputs(154);
    outputs(1101) <= not(layer2_outputs(551)) or (layer2_outputs(1012));
    outputs(1102) <= not((layer2_outputs(222)) and (layer2_outputs(938)));
    outputs(1103) <= layer2_outputs(111);
    outputs(1104) <= not(layer2_outputs(1338));
    outputs(1105) <= layer2_outputs(817);
    outputs(1106) <= (layer2_outputs(442)) or (layer2_outputs(906));
    outputs(1107) <= (layer2_outputs(985)) and not (layer2_outputs(193));
    outputs(1108) <= not(layer2_outputs(1022));
    outputs(1109) <= (layer2_outputs(1846)) or (layer2_outputs(1713));
    outputs(1110) <= not(layer2_outputs(1680));
    outputs(1111) <= not(layer2_outputs(1360));
    outputs(1112) <= layer2_outputs(2211);
    outputs(1113) <= layer2_outputs(133);
    outputs(1114) <= not((layer2_outputs(70)) or (layer2_outputs(2406)));
    outputs(1115) <= layer2_outputs(1764);
    outputs(1116) <= layer2_outputs(2325);
    outputs(1117) <= (layer2_outputs(1275)) and not (layer2_outputs(1507));
    outputs(1118) <= layer2_outputs(1159);
    outputs(1119) <= not(layer2_outputs(2038));
    outputs(1120) <= not(layer2_outputs(1649)) or (layer2_outputs(953));
    outputs(1121) <= layer2_outputs(1976);
    outputs(1122) <= not(layer2_outputs(1207));
    outputs(1123) <= not(layer2_outputs(359));
    outputs(1124) <= layer2_outputs(2445);
    outputs(1125) <= layer2_outputs(1987);
    outputs(1126) <= not(layer2_outputs(1858));
    outputs(1127) <= not(layer2_outputs(2490));
    outputs(1128) <= layer2_outputs(1876);
    outputs(1129) <= (layer2_outputs(2441)) and (layer2_outputs(548));
    outputs(1130) <= not(layer2_outputs(2534)) or (layer2_outputs(1821));
    outputs(1131) <= not(layer2_outputs(1399)) or (layer2_outputs(796));
    outputs(1132) <= layer2_outputs(225);
    outputs(1133) <= (layer2_outputs(1127)) and not (layer2_outputs(1745));
    outputs(1134) <= not(layer2_outputs(1040));
    outputs(1135) <= layer2_outputs(2094);
    outputs(1136) <= not((layer2_outputs(1469)) or (layer2_outputs(695)));
    outputs(1137) <= (layer2_outputs(1173)) and not (layer2_outputs(284));
    outputs(1138) <= (layer2_outputs(783)) xor (layer2_outputs(10));
    outputs(1139) <= not((layer2_outputs(470)) or (layer2_outputs(2415)));
    outputs(1140) <= layer2_outputs(2176);
    outputs(1141) <= layer2_outputs(1631);
    outputs(1142) <= layer2_outputs(133);
    outputs(1143) <= layer2_outputs(275);
    outputs(1144) <= layer2_outputs(129);
    outputs(1145) <= not(layer2_outputs(338));
    outputs(1146) <= not(layer2_outputs(606));
    outputs(1147) <= layer2_outputs(1552);
    outputs(1148) <= not((layer2_outputs(221)) xor (layer2_outputs(981)));
    outputs(1149) <= not(layer2_outputs(1719)) or (layer2_outputs(475));
    outputs(1150) <= not((layer2_outputs(220)) or (layer2_outputs(889)));
    outputs(1151) <= (layer2_outputs(2130)) and (layer2_outputs(1494));
    outputs(1152) <= not((layer2_outputs(691)) xor (layer2_outputs(2007)));
    outputs(1153) <= layer2_outputs(180);
    outputs(1154) <= not(layer2_outputs(218));
    outputs(1155) <= layer2_outputs(1406);
    outputs(1156) <= not((layer2_outputs(2420)) or (layer2_outputs(2298)));
    outputs(1157) <= layer2_outputs(1549);
    outputs(1158) <= (layer2_outputs(618)) and not (layer2_outputs(325));
    outputs(1159) <= layer2_outputs(2493);
    outputs(1160) <= not((layer2_outputs(1893)) xor (layer2_outputs(2414)));
    outputs(1161) <= not(layer2_outputs(2540));
    outputs(1162) <= not(layer2_outputs(549));
    outputs(1163) <= layer2_outputs(2510);
    outputs(1164) <= not(layer2_outputs(201));
    outputs(1165) <= not(layer2_outputs(1279));
    outputs(1166) <= not(layer2_outputs(1975));
    outputs(1167) <= layer2_outputs(2009);
    outputs(1168) <= (layer2_outputs(711)) and (layer2_outputs(2148));
    outputs(1169) <= not(layer2_outputs(1469));
    outputs(1170) <= layer2_outputs(2499);
    outputs(1171) <= not(layer2_outputs(1499));
    outputs(1172) <= not(layer2_outputs(1218));
    outputs(1173) <= not((layer2_outputs(2500)) or (layer2_outputs(1166)));
    outputs(1174) <= not(layer2_outputs(868));
    outputs(1175) <= not(layer2_outputs(305));
    outputs(1176) <= not(layer2_outputs(233));
    outputs(1177) <= not(layer2_outputs(1373));
    outputs(1178) <= not(layer2_outputs(2551));
    outputs(1179) <= not(layer2_outputs(383)) or (layer2_outputs(1010));
    outputs(1180) <= (layer2_outputs(2545)) and not (layer2_outputs(1452));
    outputs(1181) <= not((layer2_outputs(113)) or (layer2_outputs(1866)));
    outputs(1182) <= layer2_outputs(928);
    outputs(1183) <= layer2_outputs(886);
    outputs(1184) <= not(layer2_outputs(2197));
    outputs(1185) <= layer2_outputs(908);
    outputs(1186) <= layer2_outputs(1300);
    outputs(1187) <= layer2_outputs(444);
    outputs(1188) <= (layer2_outputs(2049)) and (layer2_outputs(1393));
    outputs(1189) <= not(layer2_outputs(207)) or (layer2_outputs(1339));
    outputs(1190) <= not(layer2_outputs(1992)) or (layer2_outputs(1579));
    outputs(1191) <= (layer2_outputs(917)) and not (layer2_outputs(607));
    outputs(1192) <= not((layer2_outputs(1000)) or (layer2_outputs(1565)));
    outputs(1193) <= (layer2_outputs(1531)) and not (layer2_outputs(2398));
    outputs(1194) <= not(layer2_outputs(49));
    outputs(1195) <= (layer2_outputs(1311)) and not (layer2_outputs(716));
    outputs(1196) <= (layer2_outputs(1027)) and (layer2_outputs(2031));
    outputs(1197) <= layer2_outputs(2387);
    outputs(1198) <= not(layer2_outputs(2416));
    outputs(1199) <= layer2_outputs(2236);
    outputs(1200) <= layer2_outputs(1111);
    outputs(1201) <= not(layer2_outputs(1536));
    outputs(1202) <= layer2_outputs(1113);
    outputs(1203) <= not((layer2_outputs(1695)) or (layer2_outputs(1207)));
    outputs(1204) <= not(layer2_outputs(1771));
    outputs(1205) <= not(layer2_outputs(876));
    outputs(1206) <= not((layer2_outputs(1142)) or (layer2_outputs(1944)));
    outputs(1207) <= not(layer2_outputs(692));
    outputs(1208) <= (layer2_outputs(80)) and not (layer2_outputs(614));
    outputs(1209) <= not((layer2_outputs(1248)) or (layer2_outputs(2295)));
    outputs(1210) <= not((layer2_outputs(827)) or (layer2_outputs(1500)));
    outputs(1211) <= not(layer2_outputs(460));
    outputs(1212) <= not(layer2_outputs(2117));
    outputs(1213) <= not(layer2_outputs(1604));
    outputs(1214) <= not(layer2_outputs(167));
    outputs(1215) <= not(layer2_outputs(2426));
    outputs(1216) <= not(layer2_outputs(1641));
    outputs(1217) <= not(layer2_outputs(41));
    outputs(1218) <= not((layer2_outputs(1532)) or (layer2_outputs(368)));
    outputs(1219) <= not(layer2_outputs(93));
    outputs(1220) <= not(layer2_outputs(39));
    outputs(1221) <= layer2_outputs(509);
    outputs(1222) <= layer2_outputs(663);
    outputs(1223) <= layer2_outputs(2182);
    outputs(1224) <= not(layer2_outputs(1362));
    outputs(1225) <= layer2_outputs(2507);
    outputs(1226) <= (layer2_outputs(1240)) and not (layer2_outputs(687));
    outputs(1227) <= not(layer2_outputs(793));
    outputs(1228) <= layer2_outputs(1552);
    outputs(1229) <= not(layer2_outputs(2262));
    outputs(1230) <= not(layer2_outputs(827));
    outputs(1231) <= (layer2_outputs(2535)) and not (layer2_outputs(1194));
    outputs(1232) <= not(layer2_outputs(130));
    outputs(1233) <= layer2_outputs(1135);
    outputs(1234) <= not(layer2_outputs(1143));
    outputs(1235) <= not(layer2_outputs(600));
    outputs(1236) <= not(layer2_outputs(922)) or (layer2_outputs(144));
    outputs(1237) <= layer2_outputs(60);
    outputs(1238) <= not(layer2_outputs(76));
    outputs(1239) <= not(layer2_outputs(2404)) or (layer2_outputs(311));
    outputs(1240) <= not(layer2_outputs(282));
    outputs(1241) <= (layer2_outputs(2333)) and not (layer2_outputs(1321));
    outputs(1242) <= not(layer2_outputs(992));
    outputs(1243) <= not((layer2_outputs(2152)) xor (layer2_outputs(2024)));
    outputs(1244) <= layer2_outputs(1834);
    outputs(1245) <= layer2_outputs(2318);
    outputs(1246) <= layer2_outputs(1854);
    outputs(1247) <= layer2_outputs(1769);
    outputs(1248) <= not(layer2_outputs(63));
    outputs(1249) <= (layer2_outputs(1411)) xor (layer2_outputs(2202));
    outputs(1250) <= layer2_outputs(1744);
    outputs(1251) <= not(layer2_outputs(844)) or (layer2_outputs(1388));
    outputs(1252) <= (layer2_outputs(1088)) and (layer2_outputs(1212));
    outputs(1253) <= (layer2_outputs(2391)) or (layer2_outputs(202));
    outputs(1254) <= not((layer2_outputs(1268)) and (layer2_outputs(1384)));
    outputs(1255) <= layer2_outputs(2439);
    outputs(1256) <= layer2_outputs(1049);
    outputs(1257) <= not(layer2_outputs(1852));
    outputs(1258) <= layer2_outputs(1372);
    outputs(1259) <= layer2_outputs(997);
    outputs(1260) <= not((layer2_outputs(1210)) xor (layer2_outputs(1660)));
    outputs(1261) <= (layer2_outputs(1101)) and not (layer2_outputs(274));
    outputs(1262) <= not(layer2_outputs(680));
    outputs(1263) <= not(layer2_outputs(596));
    outputs(1264) <= not((layer2_outputs(2119)) and (layer2_outputs(977)));
    outputs(1265) <= not(layer2_outputs(86));
    outputs(1266) <= (layer2_outputs(500)) xor (layer2_outputs(1875));
    outputs(1267) <= not(layer2_outputs(1546));
    outputs(1268) <= layer2_outputs(2552);
    outputs(1269) <= layer2_outputs(1647);
    outputs(1270) <= not((layer2_outputs(1581)) or (layer2_outputs(2017)));
    outputs(1271) <= layer2_outputs(633);
    outputs(1272) <= layer2_outputs(1291);
    outputs(1273) <= not(layer2_outputs(107));
    outputs(1274) <= not(layer2_outputs(1451));
    outputs(1275) <= not((layer2_outputs(1949)) or (layer2_outputs(1748)));
    outputs(1276) <= not(layer2_outputs(2508));
    outputs(1277) <= not((layer2_outputs(5)) or (layer2_outputs(2214)));
    outputs(1278) <= (layer2_outputs(1119)) and not (layer2_outputs(56));
    outputs(1279) <= layer2_outputs(1812);
    outputs(1280) <= layer2_outputs(347);
    outputs(1281) <= layer2_outputs(1667);
    outputs(1282) <= not(layer2_outputs(1068));
    outputs(1283) <= not((layer2_outputs(993)) or (layer2_outputs(1432)));
    outputs(1284) <= not((layer2_outputs(244)) or (layer2_outputs(71)));
    outputs(1285) <= not((layer2_outputs(36)) or (layer2_outputs(1582)));
    outputs(1286) <= not(layer2_outputs(1715));
    outputs(1287) <= not(layer2_outputs(1784));
    outputs(1288) <= not(layer2_outputs(1669));
    outputs(1289) <= not((layer2_outputs(1713)) or (layer2_outputs(1076)));
    outputs(1290) <= not(layer2_outputs(752));
    outputs(1291) <= (layer2_outputs(2431)) and not (layer2_outputs(302));
    outputs(1292) <= not(layer2_outputs(601)) or (layer2_outputs(2180));
    outputs(1293) <= not((layer2_outputs(1036)) xor (layer2_outputs(2518)));
    outputs(1294) <= (layer2_outputs(940)) and not (layer2_outputs(287));
    outputs(1295) <= (layer2_outputs(2148)) xor (layer2_outputs(1121));
    outputs(1296) <= not(layer2_outputs(894));
    outputs(1297) <= layer2_outputs(1799);
    outputs(1298) <= (layer2_outputs(1693)) and (layer2_outputs(2089));
    outputs(1299) <= layer2_outputs(75);
    outputs(1300) <= (layer2_outputs(522)) and (layer2_outputs(366));
    outputs(1301) <= (layer2_outputs(1473)) and (layer2_outputs(1857));
    outputs(1302) <= layer2_outputs(1270);
    outputs(1303) <= layer2_outputs(2253);
    outputs(1304) <= not((layer2_outputs(256)) or (layer2_outputs(875)));
    outputs(1305) <= layer2_outputs(314);
    outputs(1306) <= not(layer2_outputs(2461));
    outputs(1307) <= not(layer2_outputs(2411));
    outputs(1308) <= (layer2_outputs(783)) and (layer2_outputs(338));
    outputs(1309) <= layer2_outputs(2238);
    outputs(1310) <= (layer2_outputs(501)) xor (layer2_outputs(2513));
    outputs(1311) <= layer2_outputs(1181);
    outputs(1312) <= layer2_outputs(2000);
    outputs(1313) <= not(layer2_outputs(1601));
    outputs(1314) <= not((layer2_outputs(2050)) or (layer2_outputs(1346)));
    outputs(1315) <= (layer2_outputs(371)) and (layer2_outputs(1227));
    outputs(1316) <= (layer2_outputs(1070)) and not (layer2_outputs(1462));
    outputs(1317) <= not(layer2_outputs(412));
    outputs(1318) <= (layer2_outputs(120)) and not (layer2_outputs(2407));
    outputs(1319) <= not(layer2_outputs(810));
    outputs(1320) <= (layer2_outputs(3)) and not (layer2_outputs(12));
    outputs(1321) <= not(layer2_outputs(708));
    outputs(1322) <= (layer2_outputs(2244)) and not (layer2_outputs(2263));
    outputs(1323) <= not(layer2_outputs(593));
    outputs(1324) <= (layer2_outputs(973)) and (layer2_outputs(149));
    outputs(1325) <= (layer2_outputs(165)) and not (layer2_outputs(1152));
    outputs(1326) <= layer2_outputs(45);
    outputs(1327) <= (layer2_outputs(1635)) and (layer2_outputs(1423));
    outputs(1328) <= (layer2_outputs(1327)) and not (layer2_outputs(2478));
    outputs(1329) <= layer2_outputs(1414);
    outputs(1330) <= (layer2_outputs(1575)) and not (layer2_outputs(306));
    outputs(1331) <= (layer2_outputs(2480)) xor (layer2_outputs(2044));
    outputs(1332) <= layer2_outputs(253);
    outputs(1333) <= not(layer2_outputs(1744));
    outputs(1334) <= (layer2_outputs(1486)) and not (layer2_outputs(1614));
    outputs(1335) <= (layer2_outputs(409)) and not (layer2_outputs(1919));
    outputs(1336) <= (layer2_outputs(116)) and not (layer2_outputs(2337));
    outputs(1337) <= not(layer2_outputs(1288));
    outputs(1338) <= not((layer2_outputs(247)) or (layer2_outputs(539)));
    outputs(1339) <= not(layer2_outputs(1100));
    outputs(1340) <= not((layer2_outputs(968)) or (layer2_outputs(877)));
    outputs(1341) <= layer2_outputs(1414);
    outputs(1342) <= not(layer2_outputs(2449));
    outputs(1343) <= layer2_outputs(1136);
    outputs(1344) <= not(layer2_outputs(203)) or (layer2_outputs(1306));
    outputs(1345) <= (layer2_outputs(935)) and (layer2_outputs(904));
    outputs(1346) <= layer2_outputs(520);
    outputs(1347) <= (layer2_outputs(1736)) and not (layer2_outputs(1068));
    outputs(1348) <= not((layer2_outputs(1072)) xor (layer2_outputs(2100)));
    outputs(1349) <= not((layer2_outputs(565)) xor (layer2_outputs(2451)));
    outputs(1350) <= not(layer2_outputs(2250));
    outputs(1351) <= (layer2_outputs(129)) and not (layer2_outputs(1617));
    outputs(1352) <= not((layer2_outputs(2093)) or (layer2_outputs(758)));
    outputs(1353) <= (layer2_outputs(189)) xor (layer2_outputs(2436));
    outputs(1354) <= (layer2_outputs(823)) and (layer2_outputs(419));
    outputs(1355) <= layer2_outputs(1868);
    outputs(1356) <= not(layer2_outputs(1188));
    outputs(1357) <= not((layer2_outputs(1899)) xor (layer2_outputs(50)));
    outputs(1358) <= layer2_outputs(1972);
    outputs(1359) <= layer2_outputs(341);
    outputs(1360) <= not(layer2_outputs(1734));
    outputs(1361) <= not(layer2_outputs(2265));
    outputs(1362) <= layer2_outputs(901);
    outputs(1363) <= not(layer2_outputs(2109));
    outputs(1364) <= not(layer2_outputs(527)) or (layer2_outputs(1500));
    outputs(1365) <= not(layer2_outputs(2328));
    outputs(1366) <= layer2_outputs(1776);
    outputs(1367) <= (layer2_outputs(604)) and not (layer2_outputs(1378));
    outputs(1368) <= (layer2_outputs(1831)) and not (layer2_outputs(1509));
    outputs(1369) <= layer2_outputs(1809);
    outputs(1370) <= not(layer2_outputs(2334));
    outputs(1371) <= layer2_outputs(82);
    outputs(1372) <= (layer2_outputs(1687)) and not (layer2_outputs(534));
    outputs(1373) <= not((layer2_outputs(1820)) xor (layer2_outputs(2006)));
    outputs(1374) <= layer2_outputs(1845);
    outputs(1375) <= not((layer2_outputs(781)) or (layer2_outputs(1154)));
    outputs(1376) <= layer2_outputs(1024);
    outputs(1377) <= (layer2_outputs(1616)) and not (layer2_outputs(1204));
    outputs(1378) <= layer2_outputs(2422);
    outputs(1379) <= layer2_outputs(95);
    outputs(1380) <= (layer2_outputs(541)) and not (layer2_outputs(118));
    outputs(1381) <= layer2_outputs(2358);
    outputs(1382) <= layer2_outputs(435);
    outputs(1383) <= not(layer2_outputs(862)) or (layer2_outputs(1810));
    outputs(1384) <= layer2_outputs(85);
    outputs(1385) <= not(layer2_outputs(1104)) or (layer2_outputs(1075));
    outputs(1386) <= layer2_outputs(1006);
    outputs(1387) <= (layer2_outputs(1153)) and not (layer2_outputs(629));
    outputs(1388) <= layer2_outputs(377);
    outputs(1389) <= not(layer2_outputs(2421)) or (layer2_outputs(2271));
    outputs(1390) <= layer2_outputs(1458);
    outputs(1391) <= layer2_outputs(1057);
    outputs(1392) <= layer2_outputs(948);
    outputs(1393) <= not((layer2_outputs(953)) xor (layer2_outputs(1563)));
    outputs(1394) <= not(layer2_outputs(2412));
    outputs(1395) <= (layer2_outputs(382)) and not (layer2_outputs(1811));
    outputs(1396) <= not((layer2_outputs(544)) or (layer2_outputs(102)));
    outputs(1397) <= not(layer2_outputs(986));
    outputs(1398) <= not(layer2_outputs(828)) or (layer2_outputs(2273));
    outputs(1399) <= layer2_outputs(916);
    outputs(1400) <= layer2_outputs(66);
    outputs(1401) <= not(layer2_outputs(1287));
    outputs(1402) <= not(layer2_outputs(952));
    outputs(1403) <= layer2_outputs(936);
    outputs(1404) <= (layer2_outputs(88)) and not (layer2_outputs(238));
    outputs(1405) <= (layer2_outputs(191)) and not (layer2_outputs(425));
    outputs(1406) <= (layer2_outputs(1649)) and not (layer2_outputs(2245));
    outputs(1407) <= not(layer2_outputs(1527));
    outputs(1408) <= layer2_outputs(2422);
    outputs(1409) <= not((layer2_outputs(965)) xor (layer2_outputs(639)));
    outputs(1410) <= (layer2_outputs(990)) xor (layer2_outputs(1425));
    outputs(1411) <= not((layer2_outputs(1422)) xor (layer2_outputs(2509)));
    outputs(1412) <= not((layer2_outputs(2010)) or (layer2_outputs(1562)));
    outputs(1413) <= not(layer2_outputs(2171));
    outputs(1414) <= not((layer2_outputs(2394)) or (layer2_outputs(1905)));
    outputs(1415) <= not((layer2_outputs(1630)) xor (layer2_outputs(482)));
    outputs(1416) <= (layer2_outputs(683)) and not (layer2_outputs(1158));
    outputs(1417) <= layer2_outputs(1278);
    outputs(1418) <= not(layer2_outputs(1167));
    outputs(1419) <= (layer2_outputs(2175)) xor (layer2_outputs(2258));
    outputs(1420) <= not(layer2_outputs(1076));
    outputs(1421) <= not(layer2_outputs(1512));
    outputs(1422) <= not((layer2_outputs(1149)) xor (layer2_outputs(1969)));
    outputs(1423) <= not((layer2_outputs(340)) or (layer2_outputs(2084)));
    outputs(1424) <= not(layer2_outputs(239)) or (layer2_outputs(581));
    outputs(1425) <= not(layer2_outputs(2143));
    outputs(1426) <= not(layer2_outputs(1019));
    outputs(1427) <= not((layer2_outputs(1675)) and (layer2_outputs(2139)));
    outputs(1428) <= not(layer2_outputs(811)) or (layer2_outputs(90));
    outputs(1429) <= not(layer2_outputs(640));
    outputs(1430) <= layer2_outputs(1029);
    outputs(1431) <= (layer2_outputs(1824)) and (layer2_outputs(915));
    outputs(1432) <= not((layer2_outputs(1650)) xor (layer2_outputs(1749)));
    outputs(1433) <= not(layer2_outputs(2087));
    outputs(1434) <= not(layer2_outputs(947));
    outputs(1435) <= layer2_outputs(520);
    outputs(1436) <= not(layer2_outputs(1935));
    outputs(1437) <= not((layer2_outputs(83)) or (layer2_outputs(2274)));
    outputs(1438) <= (layer2_outputs(1053)) and (layer2_outputs(65));
    outputs(1439) <= layer2_outputs(1315);
    outputs(1440) <= not(layer2_outputs(1479));
    outputs(1441) <= (layer2_outputs(931)) or (layer2_outputs(567));
    outputs(1442) <= not((layer2_outputs(929)) or (layer2_outputs(721)));
    outputs(1443) <= (layer2_outputs(847)) and not (layer2_outputs(2469));
    outputs(1444) <= layer2_outputs(716);
    outputs(1445) <= (layer2_outputs(528)) and (layer2_outputs(1281));
    outputs(1446) <= not(layer2_outputs(1510));
    outputs(1447) <= (layer2_outputs(1459)) and not (layer2_outputs(1518));
    outputs(1448) <= not((layer2_outputs(718)) or (layer2_outputs(175)));
    outputs(1449) <= not((layer2_outputs(483)) or (layer2_outputs(1160)));
    outputs(1450) <= not(layer2_outputs(1061));
    outputs(1451) <= layer2_outputs(1626);
    outputs(1452) <= not(layer2_outputs(467)) or (layer2_outputs(1662));
    outputs(1453) <= (layer2_outputs(251)) xor (layer2_outputs(2019));
    outputs(1454) <= not(layer2_outputs(2248));
    outputs(1455) <= (layer2_outputs(1801)) and not (layer2_outputs(1415));
    outputs(1456) <= layer2_outputs(1427);
    outputs(1457) <= (layer2_outputs(471)) and not (layer2_outputs(913));
    outputs(1458) <= not((layer2_outputs(1535)) or (layer2_outputs(510)));
    outputs(1459) <= layer2_outputs(2106);
    outputs(1460) <= (layer2_outputs(1671)) and not (layer2_outputs(1890));
    outputs(1461) <= (layer2_outputs(1688)) and not (layer2_outputs(2501));
    outputs(1462) <= (layer2_outputs(1814)) xor (layer2_outputs(160));
    outputs(1463) <= not(layer2_outputs(2073));
    outputs(1464) <= (layer2_outputs(122)) xor (layer2_outputs(1599));
    outputs(1465) <= (layer2_outputs(2503)) and (layer2_outputs(378));
    outputs(1466) <= (layer2_outputs(2042)) and (layer2_outputs(7));
    outputs(1467) <= (layer2_outputs(2000)) and not (layer2_outputs(301));
    outputs(1468) <= not(layer2_outputs(2067));
    outputs(1469) <= not((layer2_outputs(1549)) and (layer2_outputs(1220)));
    outputs(1470) <= not((layer2_outputs(1034)) or (layer2_outputs(334)));
    outputs(1471) <= layer2_outputs(1946);
    outputs(1472) <= layer2_outputs(509);
    outputs(1473) <= (layer2_outputs(2172)) and not (layer2_outputs(2470));
    outputs(1474) <= layer2_outputs(1514);
    outputs(1475) <= (layer2_outputs(790)) and not (layer2_outputs(2348));
    outputs(1476) <= (layer2_outputs(1114)) and (layer2_outputs(1790));
    outputs(1477) <= not(layer2_outputs(2364));
    outputs(1478) <= (layer2_outputs(2052)) or (layer2_outputs(1616));
    outputs(1479) <= not(layer2_outputs(1463));
    outputs(1480) <= not(layer2_outputs(403));
    outputs(1481) <= layer2_outputs(1574);
    outputs(1482) <= not(layer2_outputs(1310)) or (layer2_outputs(1473));
    outputs(1483) <= not((layer2_outputs(2223)) xor (layer2_outputs(1215)));
    outputs(1484) <= (layer2_outputs(1551)) xor (layer2_outputs(1977));
    outputs(1485) <= (layer2_outputs(1070)) and not (layer2_outputs(2250));
    outputs(1486) <= not((layer2_outputs(1841)) xor (layer2_outputs(362)));
    outputs(1487) <= (layer2_outputs(1161)) and not (layer2_outputs(320));
    outputs(1488) <= not(layer2_outputs(1497)) or (layer2_outputs(508));
    outputs(1489) <= (layer2_outputs(1492)) xor (layer2_outputs(776));
    outputs(1490) <= not(layer2_outputs(1262));
    outputs(1491) <= not(layer2_outputs(2131));
    outputs(1492) <= (layer2_outputs(1275)) xor (layer2_outputs(1559));
    outputs(1493) <= (layer2_outputs(1122)) xor (layer2_outputs(1079));
    outputs(1494) <= layer2_outputs(2098);
    outputs(1495) <= (layer2_outputs(1320)) and (layer2_outputs(897));
    outputs(1496) <= (layer2_outputs(10)) and not (layer2_outputs(557));
    outputs(1497) <= (layer2_outputs(808)) xor (layer2_outputs(34));
    outputs(1498) <= not((layer2_outputs(275)) xor (layer2_outputs(1369)));
    outputs(1499) <= not(layer2_outputs(2050));
    outputs(1500) <= layer2_outputs(2477);
    outputs(1501) <= not(layer2_outputs(1142));
    outputs(1502) <= not(layer2_outputs(418));
    outputs(1503) <= not(layer2_outputs(1120));
    outputs(1504) <= (layer2_outputs(1826)) and not (layer2_outputs(2470));
    outputs(1505) <= not(layer2_outputs(1788));
    outputs(1506) <= not((layer2_outputs(333)) xor (layer2_outputs(925)));
    outputs(1507) <= not(layer2_outputs(1357));
    outputs(1508) <= not(layer2_outputs(2330));
    outputs(1509) <= not((layer2_outputs(1775)) or (layer2_outputs(290)));
    outputs(1510) <= (layer2_outputs(1681)) and not (layer2_outputs(2078));
    outputs(1511) <= (layer2_outputs(1069)) and (layer2_outputs(2255));
    outputs(1512) <= (layer2_outputs(901)) and (layer2_outputs(533));
    outputs(1513) <= (layer2_outputs(1956)) and not (layer2_outputs(603));
    outputs(1514) <= not(layer2_outputs(1676));
    outputs(1515) <= not(layer2_outputs(1782));
    outputs(1516) <= (layer2_outputs(2189)) and (layer2_outputs(1372));
    outputs(1517) <= (layer2_outputs(2298)) and (layer2_outputs(1352));
    outputs(1518) <= (layer2_outputs(1439)) or (layer2_outputs(2237));
    outputs(1519) <= not(layer2_outputs(352));
    outputs(1520) <= (layer2_outputs(1693)) and not (layer2_outputs(1043));
    outputs(1521) <= not((layer2_outputs(2023)) xor (layer2_outputs(262)));
    outputs(1522) <= (layer2_outputs(989)) or (layer2_outputs(342));
    outputs(1523) <= not(layer2_outputs(104)) or (layer2_outputs(1117));
    outputs(1524) <= (layer2_outputs(1796)) and not (layer2_outputs(2529));
    outputs(1525) <= not(layer2_outputs(1596));
    outputs(1526) <= layer2_outputs(1383);
    outputs(1527) <= (layer2_outputs(2116)) xor (layer2_outputs(1553));
    outputs(1528) <= not(layer2_outputs(1297));
    outputs(1529) <= not((layer2_outputs(1730)) xor (layer2_outputs(2313)));
    outputs(1530) <= not(layer2_outputs(1919));
    outputs(1531) <= (layer2_outputs(2547)) and not (layer2_outputs(803));
    outputs(1532) <= (layer2_outputs(547)) and not (layer2_outputs(1761));
    outputs(1533) <= (layer2_outputs(935)) and not (layer2_outputs(1445));
    outputs(1534) <= not(layer2_outputs(2292));
    outputs(1535) <= layer2_outputs(864);
    outputs(1536) <= layer2_outputs(658);
    outputs(1537) <= not(layer2_outputs(1336));
    outputs(1538) <= layer2_outputs(42);
    outputs(1539) <= layer2_outputs(1614);
    outputs(1540) <= layer2_outputs(1049);
    outputs(1541) <= not(layer2_outputs(2104));
    outputs(1542) <= layer2_outputs(1567);
    outputs(1543) <= (layer2_outputs(283)) and not (layer2_outputs(686));
    outputs(1544) <= not(layer2_outputs(840));
    outputs(1545) <= layer2_outputs(1063);
    outputs(1546) <= layer2_outputs(1543);
    outputs(1547) <= layer2_outputs(754);
    outputs(1548) <= not((layer2_outputs(2232)) or (layer2_outputs(328)));
    outputs(1549) <= (layer2_outputs(1122)) and not (layer2_outputs(826));
    outputs(1550) <= not(layer2_outputs(2108));
    outputs(1551) <= not((layer2_outputs(983)) or (layer2_outputs(777)));
    outputs(1552) <= not((layer2_outputs(1455)) or (layer2_outputs(751)));
    outputs(1553) <= not(layer2_outputs(2477));
    outputs(1554) <= layer2_outputs(57);
    outputs(1555) <= not((layer2_outputs(762)) and (layer2_outputs(2315)));
    outputs(1556) <= (layer2_outputs(598)) and (layer2_outputs(790));
    outputs(1557) <= (layer2_outputs(188)) and not (layer2_outputs(1688));
    outputs(1558) <= not(layer2_outputs(885));
    outputs(1559) <= (layer2_outputs(782)) and not (layer2_outputs(1447));
    outputs(1560) <= (layer2_outputs(1054)) and (layer2_outputs(2259));
    outputs(1561) <= layer2_outputs(2020);
    outputs(1562) <= not((layer2_outputs(2527)) xor (layer2_outputs(2494)));
    outputs(1563) <= layer2_outputs(389);
    outputs(1564) <= not(layer2_outputs(1644));
    outputs(1565) <= (layer2_outputs(1606)) and (layer2_outputs(2545));
    outputs(1566) <= layer2_outputs(2011);
    outputs(1567) <= not(layer2_outputs(1266));
    outputs(1568) <= layer2_outputs(2156);
    outputs(1569) <= not(layer2_outputs(1209));
    outputs(1570) <= (layer2_outputs(1884)) and not (layer2_outputs(1434));
    outputs(1571) <= layer2_outputs(1048);
    outputs(1572) <= not(layer2_outputs(6));
    outputs(1573) <= layer2_outputs(518);
    outputs(1574) <= layer2_outputs(1345);
    outputs(1575) <= (layer2_outputs(1613)) and not (layer2_outputs(2055));
    outputs(1576) <= layer2_outputs(2387);
    outputs(1577) <= not(layer2_outputs(2349));
    outputs(1578) <= (layer2_outputs(1780)) and (layer2_outputs(1643));
    outputs(1579) <= (layer2_outputs(2457)) and not (layer2_outputs(438));
    outputs(1580) <= not(layer2_outputs(117));
    outputs(1581) <= (layer2_outputs(29)) xor (layer2_outputs(2287));
    outputs(1582) <= not(layer2_outputs(1257));
    outputs(1583) <= (layer2_outputs(2488)) and (layer2_outputs(93));
    outputs(1584) <= layer2_outputs(2547);
    outputs(1585) <= (layer2_outputs(1449)) and (layer2_outputs(711));
    outputs(1586) <= not(layer2_outputs(1587));
    outputs(1587) <= (layer2_outputs(1474)) and not (layer2_outputs(1264));
    outputs(1588) <= (layer2_outputs(1400)) and not (layer2_outputs(1880));
    outputs(1589) <= not(layer2_outputs(402));
    outputs(1590) <= (layer2_outputs(1454)) xor (layer2_outputs(374));
    outputs(1591) <= layer2_outputs(1780);
    outputs(1592) <= not(layer2_outputs(1172));
    outputs(1593) <= layer2_outputs(1723);
    outputs(1594) <= (layer2_outputs(975)) and (layer2_outputs(2462));
    outputs(1595) <= not(layer2_outputs(146));
    outputs(1596) <= not(layer2_outputs(125));
    outputs(1597) <= (layer2_outputs(2359)) and not (layer2_outputs(537));
    outputs(1598) <= (layer2_outputs(1692)) and (layer2_outputs(2014));
    outputs(1599) <= layer2_outputs(822);
    outputs(1600) <= (layer2_outputs(1108)) and not (layer2_outputs(1809));
    outputs(1601) <= not((layer2_outputs(1860)) xor (layer2_outputs(1201)));
    outputs(1602) <= not((layer2_outputs(1113)) or (layer2_outputs(2516)));
    outputs(1603) <= not((layer2_outputs(1488)) and (layer2_outputs(2107)));
    outputs(1604) <= (layer2_outputs(2488)) and (layer2_outputs(2527));
    outputs(1605) <= not(layer2_outputs(223));
    outputs(1606) <= layer2_outputs(486);
    outputs(1607) <= not(layer2_outputs(956));
    outputs(1608) <= not(layer2_outputs(89)) or (layer2_outputs(995));
    outputs(1609) <= layer2_outputs(869);
    outputs(1610) <= (layer2_outputs(2357)) and not (layer2_outputs(2099));
    outputs(1611) <= (layer2_outputs(778)) xor (layer2_outputs(363));
    outputs(1612) <= (layer2_outputs(360)) and not (layer2_outputs(1501));
    outputs(1613) <= layer2_outputs(1437);
    outputs(1614) <= (layer2_outputs(335)) and (layer2_outputs(1428));
    outputs(1615) <= layer2_outputs(2032);
    outputs(1616) <= (layer2_outputs(307)) or (layer2_outputs(2030));
    outputs(1617) <= not(layer2_outputs(2216));
    outputs(1618) <= not((layer2_outputs(1822)) or (layer2_outputs(167)));
    outputs(1619) <= (layer2_outputs(1250)) xor (layer2_outputs(1350));
    outputs(1620) <= not((layer2_outputs(1286)) or (layer2_outputs(1720)));
    outputs(1621) <= not(layer2_outputs(796));
    outputs(1622) <= (layer2_outputs(1007)) and (layer2_outputs(1310));
    outputs(1623) <= layer2_outputs(1847);
    outputs(1624) <= not((layer2_outputs(2045)) and (layer2_outputs(1426)));
    outputs(1625) <= layer2_outputs(1886);
    outputs(1626) <= not(layer2_outputs(641));
    outputs(1627) <= (layer2_outputs(2224)) and not (layer2_outputs(1348));
    outputs(1628) <= layer2_outputs(448);
    outputs(1629) <= not(layer2_outputs(364)) or (layer2_outputs(1690));
    outputs(1630) <= not(layer2_outputs(1927)) or (layer2_outputs(2352));
    outputs(1631) <= not(layer2_outputs(291));
    outputs(1632) <= not(layer2_outputs(938));
    outputs(1633) <= (layer2_outputs(152)) and not (layer2_outputs(1834));
    outputs(1634) <= (layer2_outputs(543)) and not (layer2_outputs(313));
    outputs(1635) <= layer2_outputs(2081);
    outputs(1636) <= not(layer2_outputs(597)) or (layer2_outputs(1423));
    outputs(1637) <= layer2_outputs(50);
    outputs(1638) <= layer2_outputs(1216);
    outputs(1639) <= layer2_outputs(865);
    outputs(1640) <= not(layer2_outputs(545));
    outputs(1641) <= not(layer2_outputs(2442));
    outputs(1642) <= layer2_outputs(1046);
    outputs(1643) <= not(layer2_outputs(2486));
    outputs(1644) <= layer2_outputs(1002);
    outputs(1645) <= not(layer2_outputs(409));
    outputs(1646) <= layer2_outputs(569);
    outputs(1647) <= layer2_outputs(1886);
    outputs(1648) <= layer2_outputs(2188);
    outputs(1649) <= layer2_outputs(2247);
    outputs(1650) <= layer2_outputs(2158);
    outputs(1651) <= not(layer2_outputs(2004));
    outputs(1652) <= layer2_outputs(1101);
    outputs(1653) <= not((layer2_outputs(1912)) and (layer2_outputs(375)));
    outputs(1654) <= layer2_outputs(1341);
    outputs(1655) <= layer2_outputs(1477);
    outputs(1656) <= not((layer2_outputs(2437)) or (layer2_outputs(1191)));
    outputs(1657) <= not(layer2_outputs(462));
    outputs(1658) <= not(layer2_outputs(1130));
    outputs(1659) <= layer2_outputs(1493);
    outputs(1660) <= (layer2_outputs(628)) and not (layer2_outputs(2282));
    outputs(1661) <= not((layer2_outputs(110)) or (layer2_outputs(1078)));
    outputs(1662) <= not(layer2_outputs(794));
    outputs(1663) <= layer2_outputs(1942);
    outputs(1664) <= (layer2_outputs(774)) and not (layer2_outputs(537));
    outputs(1665) <= not((layer2_outputs(1092)) xor (layer2_outputs(665)));
    outputs(1666) <= layer2_outputs(308);
    outputs(1667) <= layer2_outputs(1141);
    outputs(1668) <= not(layer2_outputs(2115));
    outputs(1669) <= layer2_outputs(2345);
    outputs(1670) <= layer2_outputs(2496);
    outputs(1671) <= not(layer2_outputs(999)) or (layer2_outputs(67));
    outputs(1672) <= not(layer2_outputs(932));
    outputs(1673) <= not(layer2_outputs(1205));
    outputs(1674) <= layer2_outputs(47);
    outputs(1675) <= not(layer2_outputs(381));
    outputs(1676) <= not((layer2_outputs(1538)) or (layer2_outputs(1632)));
    outputs(1677) <= not(layer2_outputs(1244));
    outputs(1678) <= not((layer2_outputs(579)) or (layer2_outputs(257)));
    outputs(1679) <= not(layer2_outputs(1235));
    outputs(1680) <= layer2_outputs(1085);
    outputs(1681) <= layer2_outputs(921);
    outputs(1682) <= layer2_outputs(526);
    outputs(1683) <= layer2_outputs(631);
    outputs(1684) <= not(layer2_outputs(1097));
    outputs(1685) <= not((layer2_outputs(936)) and (layer2_outputs(676)));
    outputs(1686) <= not(layer2_outputs(1337));
    outputs(1687) <= not(layer2_outputs(2268));
    outputs(1688) <= not(layer2_outputs(2130));
    outputs(1689) <= not(layer2_outputs(971));
    outputs(1690) <= not((layer2_outputs(957)) or (layer2_outputs(178)));
    outputs(1691) <= layer2_outputs(1058);
    outputs(1692) <= layer2_outputs(143);
    outputs(1693) <= (layer2_outputs(1538)) xor (layer2_outputs(2421));
    outputs(1694) <= not((layer2_outputs(444)) or (layer2_outputs(187)));
    outputs(1695) <= (layer2_outputs(2432)) and not (layer2_outputs(1280));
    outputs(1696) <= layer2_outputs(1425);
    outputs(1697) <= (layer2_outputs(1409)) and not (layer2_outputs(1513));
    outputs(1698) <= not(layer2_outputs(719)) or (layer2_outputs(2492));
    outputs(1699) <= not(layer2_outputs(2464)) or (layer2_outputs(1673));
    outputs(1700) <= layer2_outputs(1863);
    outputs(1701) <= not(layer2_outputs(864));
    outputs(1702) <= not(layer2_outputs(524));
    outputs(1703) <= not(layer2_outputs(1212)) or (layer2_outputs(930));
    outputs(1704) <= (layer2_outputs(1573)) and not (layer2_outputs(2092));
    outputs(1705) <= not((layer2_outputs(2495)) or (layer2_outputs(36)));
    outputs(1706) <= (layer2_outputs(839)) and (layer2_outputs(530));
    outputs(1707) <= not(layer2_outputs(982));
    outputs(1708) <= layer2_outputs(2144);
    outputs(1709) <= (layer2_outputs(145)) or (layer2_outputs(12));
    outputs(1710) <= not((layer2_outputs(169)) or (layer2_outputs(1853)));
    outputs(1711) <= not(layer2_outputs(1485));
    outputs(1712) <= (layer2_outputs(2014)) and not (layer2_outputs(553));
    outputs(1713) <= not(layer2_outputs(1737));
    outputs(1714) <= not((layer2_outputs(247)) or (layer2_outputs(362)));
    outputs(1715) <= layer2_outputs(896);
    outputs(1716) <= (layer2_outputs(324)) and not (layer2_outputs(2385));
    outputs(1717) <= layer2_outputs(2134);
    outputs(1718) <= not(layer2_outputs(2486));
    outputs(1719) <= not(layer2_outputs(1851));
    outputs(1720) <= not(layer2_outputs(2068));
    outputs(1721) <= not(layer2_outputs(1358));
    outputs(1722) <= not(layer2_outputs(616));
    outputs(1723) <= (layer2_outputs(138)) and not (layer2_outputs(767));
    outputs(1724) <= layer2_outputs(455);
    outputs(1725) <= not(layer2_outputs(2137));
    outputs(1726) <= layer2_outputs(185);
    outputs(1727) <= not(layer2_outputs(770));
    outputs(1728) <= not(layer2_outputs(1241)) or (layer2_outputs(607));
    outputs(1729) <= not(layer2_outputs(1752));
    outputs(1730) <= (layer2_outputs(1733)) and not (layer2_outputs(2553));
    outputs(1731) <= (layer2_outputs(724)) and not (layer2_outputs(2447));
    outputs(1732) <= (layer2_outputs(1600)) and (layer2_outputs(453));
    outputs(1733) <= not(layer2_outputs(276)) or (layer2_outputs(289));
    outputs(1734) <= layer2_outputs(2346);
    outputs(1735) <= not(layer2_outputs(847));
    outputs(1736) <= layer2_outputs(1718);
    outputs(1737) <= (layer2_outputs(1)) xor (layer2_outputs(2084));
    outputs(1738) <= layer2_outputs(1859);
    outputs(1739) <= not(layer2_outputs(838));
    outputs(1740) <= not(layer2_outputs(94));
    outputs(1741) <= layer2_outputs(1506);
    outputs(1742) <= layer2_outputs(1182);
    outputs(1743) <= layer2_outputs(2048);
    outputs(1744) <= layer2_outputs(1940);
    outputs(1745) <= layer2_outputs(2083);
    outputs(1746) <= layer2_outputs(1185);
    outputs(1747) <= layer2_outputs(959);
    outputs(1748) <= (layer2_outputs(3)) xor (layer2_outputs(1955));
    outputs(1749) <= layer2_outputs(1249);
    outputs(1750) <= not(layer2_outputs(1343));
    outputs(1751) <= layer2_outputs(1793);
    outputs(1752) <= layer2_outputs(846);
    outputs(1753) <= not(layer2_outputs(2064));
    outputs(1754) <= not(layer2_outputs(39));
    outputs(1755) <= layer2_outputs(2346);
    outputs(1756) <= not((layer2_outputs(601)) or (layer2_outputs(647)));
    outputs(1757) <= not(layer2_outputs(1514));
    outputs(1758) <= layer2_outputs(2024);
    outputs(1759) <= not(layer2_outputs(1456));
    outputs(1760) <= layer2_outputs(1993);
    outputs(1761) <= not((layer2_outputs(1760)) or (layer2_outputs(567)));
    outputs(1762) <= not(layer2_outputs(1946));
    outputs(1763) <= layer2_outputs(1221);
    outputs(1764) <= not((layer2_outputs(1825)) or (layer2_outputs(1160)));
    outputs(1765) <= not((layer2_outputs(1873)) or (layer2_outputs(568)));
    outputs(1766) <= (layer2_outputs(163)) or (layer2_outputs(1636));
    outputs(1767) <= (layer2_outputs(747)) and not (layer2_outputs(539));
    outputs(1768) <= (layer2_outputs(2083)) and not (layer2_outputs(2471));
    outputs(1769) <= not(layer2_outputs(1441));
    outputs(1770) <= (layer2_outputs(642)) and not (layer2_outputs(466));
    outputs(1771) <= not(layer2_outputs(146)) or (layer2_outputs(978));
    outputs(1772) <= (layer2_outputs(877)) or (layer2_outputs(1700));
    outputs(1773) <= (layer2_outputs(1755)) and (layer2_outputs(2209));
    outputs(1774) <= (layer2_outputs(232)) and (layer2_outputs(1975));
    outputs(1775) <= (layer2_outputs(1832)) and not (layer2_outputs(1721));
    outputs(1776) <= layer2_outputs(1528);
    outputs(1777) <= (layer2_outputs(2472)) and (layer2_outputs(784));
    outputs(1778) <= layer2_outputs(1931);
    outputs(1779) <= (layer2_outputs(602)) xor (layer2_outputs(46));
    outputs(1780) <= not((layer2_outputs(1431)) or (layer2_outputs(1555)));
    outputs(1781) <= (layer2_outputs(995)) and (layer2_outputs(621));
    outputs(1782) <= layer2_outputs(59);
    outputs(1783) <= (layer2_outputs(2551)) and not (layer2_outputs(1731));
    outputs(1784) <= not((layer2_outputs(245)) or (layer2_outputs(1065)));
    outputs(1785) <= (layer2_outputs(331)) xor (layer2_outputs(950));
    outputs(1786) <= layer2_outputs(671);
    outputs(1787) <= (layer2_outputs(2069)) and not (layer2_outputs(2507));
    outputs(1788) <= (layer2_outputs(2316)) or (layer2_outputs(1739));
    outputs(1789) <= not(layer2_outputs(414));
    outputs(1790) <= not((layer2_outputs(1517)) or (layer2_outputs(2350)));
    outputs(1791) <= (layer2_outputs(506)) and not (layer2_outputs(2471));
    outputs(1792) <= (layer2_outputs(1017)) and (layer2_outputs(1178));
    outputs(1793) <= not(layer2_outputs(2446));
    outputs(1794) <= not((layer2_outputs(2251)) or (layer2_outputs(1356)));
    outputs(1795) <= (layer2_outputs(1220)) and not (layer2_outputs(1077));
    outputs(1796) <= not(layer2_outputs(2091));
    outputs(1797) <= not(layer2_outputs(1466));
    outputs(1798) <= not((layer2_outputs(2026)) or (layer2_outputs(2528)));
    outputs(1799) <= not(layer2_outputs(673));
    outputs(1800) <= layer2_outputs(2057);
    outputs(1801) <= (layer2_outputs(54)) and not (layer2_outputs(159));
    outputs(1802) <= (layer2_outputs(945)) and not (layer2_outputs(237));
    outputs(1803) <= (layer2_outputs(2412)) and not (layer2_outputs(787));
    outputs(1804) <= layer2_outputs(816);
    outputs(1805) <= not(layer2_outputs(360));
    outputs(1806) <= not(layer2_outputs(2264));
    outputs(1807) <= not(layer2_outputs(2537));
    outputs(1808) <= not(layer2_outputs(2373));
    outputs(1809) <= not(layer2_outputs(2379));
    outputs(1810) <= layer2_outputs(353);
    outputs(1811) <= layer2_outputs(1316);
    outputs(1812) <= not((layer2_outputs(2133)) or (layer2_outputs(1058)));
    outputs(1813) <= not(layer2_outputs(2114));
    outputs(1814) <= not((layer2_outputs(1227)) and (layer2_outputs(1586)));
    outputs(1815) <= (layer2_outputs(110)) or (layer2_outputs(2135));
    outputs(1816) <= (layer2_outputs(1924)) or (layer2_outputs(2443));
    outputs(1817) <= (layer2_outputs(1443)) and not (layer2_outputs(1470));
    outputs(1818) <= (layer2_outputs(1672)) and not (layer2_outputs(337));
    outputs(1819) <= (layer2_outputs(349)) and (layer2_outputs(1038));
    outputs(1820) <= not(layer2_outputs(1918));
    outputs(1821) <= (layer2_outputs(1906)) and not (layer2_outputs(1507));
    outputs(1822) <= layer2_outputs(513);
    outputs(1823) <= layer2_outputs(831);
    outputs(1824) <= not((layer2_outputs(635)) xor (layer2_outputs(1338)));
    outputs(1825) <= not(layer2_outputs(2032));
    outputs(1826) <= not(layer2_outputs(933));
    outputs(1827) <= layer2_outputs(976);
    outputs(1828) <= (layer2_outputs(1471)) and not (layer2_outputs(1706));
    outputs(1829) <= (layer2_outputs(1653)) xor (layer2_outputs(473));
    outputs(1830) <= not(layer2_outputs(2281));
    outputs(1831) <= not((layer2_outputs(1023)) or (layer2_outputs(1240)));
    outputs(1832) <= (layer2_outputs(2301)) and (layer2_outputs(2284));
    outputs(1833) <= (layer2_outputs(1254)) and not (layer2_outputs(2327));
    outputs(1834) <= not(layer2_outputs(2060));
    outputs(1835) <= layer2_outputs(1487);
    outputs(1836) <= (layer2_outputs(1444)) and not (layer2_outputs(2112));
    outputs(1837) <= layer2_outputs(1481);
    outputs(1838) <= (layer2_outputs(620)) and (layer2_outputs(24));
    outputs(1839) <= (layer2_outputs(426)) and (layer2_outputs(493));
    outputs(1840) <= layer2_outputs(727);
    outputs(1841) <= not((layer2_outputs(2253)) or (layer2_outputs(1786)));
    outputs(1842) <= (layer2_outputs(2362)) and not (layer2_outputs(585));
    outputs(1843) <= (layer2_outputs(221)) or (layer2_outputs(1922));
    outputs(1844) <= not((layer2_outputs(1333)) xor (layer2_outputs(277)));
    outputs(1845) <= not(layer2_outputs(1837));
    outputs(1846) <= layer2_outputs(230);
    outputs(1847) <= (layer2_outputs(1139)) and (layer2_outputs(2021));
    outputs(1848) <= layer2_outputs(87);
    outputs(1849) <= layer2_outputs(586);
    outputs(1850) <= (layer2_outputs(768)) and (layer2_outputs(72));
    outputs(1851) <= not((layer2_outputs(95)) or (layer2_outputs(2081)));
    outputs(1852) <= layer2_outputs(666);
    outputs(1853) <= (layer2_outputs(1537)) and (layer2_outputs(1441));
    outputs(1854) <= layer2_outputs(589);
    outputs(1855) <= not(layer2_outputs(16));
    outputs(1856) <= layer2_outputs(1629);
    outputs(1857) <= layer2_outputs(2043);
    outputs(1858) <= not(layer2_outputs(2300));
    outputs(1859) <= layer2_outputs(2349);
    outputs(1860) <= (layer2_outputs(1128)) and not (layer2_outputs(240));
    outputs(1861) <= layer2_outputs(2460);
    outputs(1862) <= layer2_outputs(61);
    outputs(1863) <= (layer2_outputs(2033)) and not (layer2_outputs(2140));
    outputs(1864) <= (layer2_outputs(571)) and (layer2_outputs(1544));
    outputs(1865) <= (layer2_outputs(1546)) and (layer2_outputs(1110));
    outputs(1866) <= not(layer2_outputs(1600)) or (layer2_outputs(1174));
    outputs(1867) <= layer2_outputs(1080);
    outputs(1868) <= (layer2_outputs(1359)) and not (layer2_outputs(1418));
    outputs(1869) <= not(layer2_outputs(2264));
    outputs(1870) <= (layer2_outputs(229)) and (layer2_outputs(2072));
    outputs(1871) <= (layer2_outputs(1753)) and (layer2_outputs(961));
    outputs(1872) <= (layer2_outputs(1803)) and (layer2_outputs(479));
    outputs(1873) <= layer2_outputs(2110);
    outputs(1874) <= not(layer2_outputs(1053));
    outputs(1875) <= not(layer2_outputs(19));
    outputs(1876) <= (layer2_outputs(2166)) and (layer2_outputs(18));
    outputs(1877) <= layer2_outputs(210);
    outputs(1878) <= (layer2_outputs(20)) xor (layer2_outputs(73));
    outputs(1879) <= not((layer2_outputs(699)) or (layer2_outputs(1031)));
    outputs(1880) <= layer2_outputs(2417);
    outputs(1881) <= (layer2_outputs(1935)) and not (layer2_outputs(1269));
    outputs(1882) <= not((layer2_outputs(1201)) or (layer2_outputs(213)));
    outputs(1883) <= not(layer2_outputs(2149));
    outputs(1884) <= layer2_outputs(1726);
    outputs(1885) <= not(layer2_outputs(2532));
    outputs(1886) <= layer2_outputs(230);
    outputs(1887) <= layer2_outputs(955);
    outputs(1888) <= (layer2_outputs(1603)) and (layer2_outputs(2525));
    outputs(1889) <= layer2_outputs(187);
    outputs(1890) <= (layer2_outputs(1871)) and not (layer2_outputs(47));
    outputs(1891) <= layer2_outputs(1998);
    outputs(1892) <= layer2_outputs(2519);
    outputs(1893) <= (layer2_outputs(306)) or (layer2_outputs(1124));
    outputs(1894) <= layer2_outputs(525);
    outputs(1895) <= layer2_outputs(1177);
    outputs(1896) <= not(layer2_outputs(2090));
    outputs(1897) <= not(layer2_outputs(419));
    outputs(1898) <= not(layer2_outputs(984));
    outputs(1899) <= layer2_outputs(923);
    outputs(1900) <= not(layer2_outputs(359));
    outputs(1901) <= (layer2_outputs(1084)) and (layer2_outputs(2341));
    outputs(1902) <= not(layer2_outputs(2498));
    outputs(1903) <= layer2_outputs(1947);
    outputs(1904) <= (layer2_outputs(1502)) and not (layer2_outputs(1345));
    outputs(1905) <= not(layer2_outputs(1137));
    outputs(1906) <= layer2_outputs(2357);
    outputs(1907) <= (layer2_outputs(1888)) xor (layer2_outputs(1498));
    outputs(1908) <= (layer2_outputs(2129)) and not (layer2_outputs(1478));
    outputs(1909) <= (layer2_outputs(531)) and not (layer2_outputs(1382));
    outputs(1910) <= not(layer2_outputs(916));
    outputs(1911) <= not(layer2_outputs(1353));
    outputs(1912) <= not(layer2_outputs(232));
    outputs(1913) <= not(layer2_outputs(1561));
    outputs(1914) <= (layer2_outputs(1442)) or (layer2_outputs(404));
    outputs(1915) <= (layer2_outputs(1095)) and (layer2_outputs(1648));
    outputs(1916) <= not((layer2_outputs(1617)) or (layer2_outputs(115)));
    outputs(1917) <= not((layer2_outputs(552)) and (layer2_outputs(78)));
    outputs(1918) <= not(layer2_outputs(311));
    outputs(1919) <= layer2_outputs(1001);
    outputs(1920) <= (layer2_outputs(2322)) and not (layer2_outputs(994));
    outputs(1921) <= layer2_outputs(1872);
    outputs(1922) <= (layer2_outputs(1354)) and not (layer2_outputs(1353));
    outputs(1923) <= (layer2_outputs(1298)) and (layer2_outputs(2186));
    outputs(1924) <= not((layer2_outputs(738)) xor (layer2_outputs(2487)));
    outputs(1925) <= (layer2_outputs(1613)) and not (layer2_outputs(1772));
    outputs(1926) <= layer2_outputs(542);
    outputs(1927) <= not(layer2_outputs(1689));
    outputs(1928) <= not(layer2_outputs(1962));
    outputs(1929) <= not(layer2_outputs(1232));
    outputs(1930) <= not(layer2_outputs(1827));
    outputs(1931) <= (layer2_outputs(1554)) and not (layer2_outputs(266));
    outputs(1932) <= layer2_outputs(532);
    outputs(1933) <= (layer2_outputs(1741)) and not (layer2_outputs(832));
    outputs(1934) <= not(layer2_outputs(1289));
    outputs(1935) <= (layer2_outputs(1864)) and not (layer2_outputs(1433));
    outputs(1936) <= not(layer2_outputs(618));
    outputs(1937) <= (layer2_outputs(1828)) xor (layer2_outputs(1615));
    outputs(1938) <= (layer2_outputs(1254)) and not (layer2_outputs(148));
    outputs(1939) <= layer2_outputs(1480);
    outputs(1940) <= not(layer2_outputs(2528));
    outputs(1941) <= (layer2_outputs(2344)) and not (layer2_outputs(842));
    outputs(1942) <= not((layer2_outputs(14)) or (layer2_outputs(1363)));
    outputs(1943) <= not(layer2_outputs(1832)) or (layer2_outputs(391));
    outputs(1944) <= (layer2_outputs(2065)) and not (layer2_outputs(1623));
    outputs(1945) <= (layer2_outputs(1105)) and (layer2_outputs(2267));
    outputs(1946) <= (layer2_outputs(272)) and not (layer2_outputs(153));
    outputs(1947) <= not(layer2_outputs(99));
    outputs(1948) <= (layer2_outputs(1768)) and not (layer2_outputs(1841));
    outputs(1949) <= (layer2_outputs(960)) or (layer2_outputs(610));
    outputs(1950) <= not((layer2_outputs(2522)) or (layer2_outputs(574)));
    outputs(1951) <= not(layer2_outputs(1560)) or (layer2_outputs(352));
    outputs(1952) <= layer2_outputs(160);
    outputs(1953) <= not((layer2_outputs(1269)) or (layer2_outputs(2122)));
    outputs(1954) <= (layer2_outputs(2037)) and not (layer2_outputs(1751));
    outputs(1955) <= not((layer2_outputs(1087)) or (layer2_outputs(1412)));
    outputs(1956) <= not(layer2_outputs(2504));
    outputs(1957) <= layer2_outputs(399);
    outputs(1958) <= (layer2_outputs(1686)) xor (layer2_outputs(1881));
    outputs(1959) <= (layer2_outputs(1235)) and not (layer2_outputs(1892));
    outputs(1960) <= layer2_outputs(806);
    outputs(1961) <= (layer2_outputs(429)) and not (layer2_outputs(147));
    outputs(1962) <= (layer2_outputs(1985)) and not (layer2_outputs(1347));
    outputs(1963) <= not(layer2_outputs(1198));
    outputs(1964) <= (layer2_outputs(33)) xor (layer2_outputs(649));
    outputs(1965) <= (layer2_outputs(690)) and not (layer2_outputs(609));
    outputs(1966) <= not((layer2_outputs(382)) and (layer2_outputs(905)));
    outputs(1967) <= not(layer2_outputs(109));
    outputs(1968) <= not(layer2_outputs(701));
    outputs(1969) <= layer2_outputs(2073);
    outputs(1970) <= layer2_outputs(665);
    outputs(1971) <= layer2_outputs(703);
    outputs(1972) <= not(layer2_outputs(578));
    outputs(1973) <= not((layer2_outputs(927)) or (layer2_outputs(1154)));
    outputs(1974) <= (layer2_outputs(258)) or (layer2_outputs(1580));
    outputs(1975) <= (layer2_outputs(1237)) and not (layer2_outputs(1835));
    outputs(1976) <= layer2_outputs(1954);
    outputs(1977) <= not(layer2_outputs(1450)) or (layer2_outputs(1556));
    outputs(1978) <= not(layer2_outputs(2198));
    outputs(1979) <= layer2_outputs(648);
    outputs(1980) <= not(layer2_outputs(918));
    outputs(1981) <= layer2_outputs(206);
    outputs(1982) <= not(layer2_outputs(2199));
    outputs(1983) <= layer2_outputs(194);
    outputs(1984) <= (layer2_outputs(2462)) xor (layer2_outputs(1440));
    outputs(1985) <= layer2_outputs(1596);
    outputs(1986) <= (layer2_outputs(196)) and not (layer2_outputs(2208));
    outputs(1987) <= (layer2_outputs(1566)) and not (layer2_outputs(148));
    outputs(1988) <= (layer2_outputs(2494)) and not (layer2_outputs(1323));
    outputs(1989) <= not((layer2_outputs(2306)) or (layer2_outputs(2290)));
    outputs(1990) <= not((layer2_outputs(1589)) or (layer2_outputs(2239)));
    outputs(1991) <= layer2_outputs(1431);
    outputs(1992) <= not(layer2_outputs(2451));
    outputs(1993) <= (layer2_outputs(2021)) and not (layer2_outputs(253));
    outputs(1994) <= (layer2_outputs(1635)) and not (layer2_outputs(1347));
    outputs(1995) <= (layer2_outputs(2542)) and (layer2_outputs(795));
    outputs(1996) <= (layer2_outputs(1761)) and not (layer2_outputs(801));
    outputs(1997) <= layer2_outputs(1753);
    outputs(1998) <= not((layer2_outputs(2514)) and (layer2_outputs(2468)));
    outputs(1999) <= not((layer2_outputs(780)) or (layer2_outputs(797)));
    outputs(2000) <= (layer2_outputs(1922)) and (layer2_outputs(983));
    outputs(2001) <= not(layer2_outputs(528));
    outputs(2002) <= (layer2_outputs(1542)) and not (layer2_outputs(2207));
    outputs(2003) <= (layer2_outputs(1852)) and not (layer2_outputs(1246));
    outputs(2004) <= not(layer2_outputs(2454));
    outputs(2005) <= not((layer2_outputs(829)) or (layer2_outputs(2244)));
    outputs(2006) <= not((layer2_outputs(615)) or (layer2_outputs(127)));
    outputs(2007) <= layer2_outputs(1084);
    outputs(2008) <= layer2_outputs(248);
    outputs(2009) <= layer2_outputs(1909);
    outputs(2010) <= layer2_outputs(870);
    outputs(2011) <= not((layer2_outputs(1689)) or (layer2_outputs(2042)));
    outputs(2012) <= not(layer2_outputs(1163));
    outputs(2013) <= (layer2_outputs(1398)) and not (layer2_outputs(701));
    outputs(2014) <= (layer2_outputs(1999)) and not (layer2_outputs(733));
    outputs(2015) <= (layer2_outputs(2402)) and not (layer2_outputs(994));
    outputs(2016) <= (layer2_outputs(1183)) and not (layer2_outputs(474));
    outputs(2017) <= (layer2_outputs(1127)) and not (layer2_outputs(1230));
    outputs(2018) <= (layer2_outputs(2405)) and not (layer2_outputs(1564));
    outputs(2019) <= not(layer2_outputs(1850));
    outputs(2020) <= not(layer2_outputs(1605));
    outputs(2021) <= (layer2_outputs(821)) and not (layer2_outputs(1072));
    outputs(2022) <= layer2_outputs(58);
    outputs(2023) <= not(layer2_outputs(2028));
    outputs(2024) <= layer2_outputs(350);
    outputs(2025) <= layer2_outputs(2085);
    outputs(2026) <= not((layer2_outputs(205)) xor (layer2_outputs(2484)));
    outputs(2027) <= layer2_outputs(1523);
    outputs(2028) <= (layer2_outputs(666)) and not (layer2_outputs(1944));
    outputs(2029) <= not((layer2_outputs(2541)) xor (layer2_outputs(1421)));
    outputs(2030) <= not((layer2_outputs(2461)) and (layer2_outputs(1108)));
    outputs(2031) <= not((layer2_outputs(911)) xor (layer2_outputs(766)));
    outputs(2032) <= not(layer2_outputs(2141));
    outputs(2033) <= (layer2_outputs(405)) and not (layer2_outputs(481));
    outputs(2034) <= not(layer2_outputs(2425));
    outputs(2035) <= layer2_outputs(41);
    outputs(2036) <= (layer2_outputs(943)) and (layer2_outputs(1238));
    outputs(2037) <= layer2_outputs(225);
    outputs(2038) <= (layer2_outputs(1008)) and not (layer2_outputs(914));
    outputs(2039) <= (layer2_outputs(72)) and not (layer2_outputs(924));
    outputs(2040) <= not(layer2_outputs(2354));
    outputs(2041) <= not(layer2_outputs(2027));
    outputs(2042) <= (layer2_outputs(902)) and not (layer2_outputs(1873));
    outputs(2043) <= not(layer2_outputs(1652));
    outputs(2044) <= not(layer2_outputs(775));
    outputs(2045) <= layer2_outputs(414);
    outputs(2046) <= not(layer2_outputs(5));
    outputs(2047) <= not((layer2_outputs(630)) or (layer2_outputs(1848)));
    outputs(2048) <= not((layer2_outputs(1199)) and (layer2_outputs(2139)));
    outputs(2049) <= (layer2_outputs(497)) and not (layer2_outputs(98));
    outputs(2050) <= layer2_outputs(2182);
    outputs(2051) <= (layer2_outputs(846)) xor (layer2_outputs(940));
    outputs(2052) <= (layer2_outputs(1643)) and (layer2_outputs(1942));
    outputs(2053) <= layer2_outputs(1099);
    outputs(2054) <= not(layer2_outputs(1676));
    outputs(2055) <= (layer2_outputs(1428)) and (layer2_outputs(1961));
    outputs(2056) <= layer2_outputs(2137);
    outputs(2057) <= not((layer2_outputs(384)) or (layer2_outputs(781)));
    outputs(2058) <= layer2_outputs(1281);
    outputs(2059) <= not((layer2_outputs(851)) or (layer2_outputs(763)));
    outputs(2060) <= layer2_outputs(2327);
    outputs(2061) <= not((layer2_outputs(530)) or (layer2_outputs(1190)));
    outputs(2062) <= not((layer2_outputs(1371)) xor (layer2_outputs(410)));
    outputs(2063) <= layer2_outputs(1171);
    outputs(2064) <= layer2_outputs(363);
    outputs(2065) <= not(layer2_outputs(671)) or (layer2_outputs(1960));
    outputs(2066) <= not(layer2_outputs(1354));
    outputs(2067) <= (layer2_outputs(1518)) xor (layer2_outputs(2377));
    outputs(2068) <= layer2_outputs(2423);
    outputs(2069) <= (layer2_outputs(1732)) and not (layer2_outputs(2251));
    outputs(2070) <= layer2_outputs(1765);
    outputs(2071) <= (layer2_outputs(900)) and (layer2_outputs(724));
    outputs(2072) <= not(layer2_outputs(1800));
    outputs(2073) <= not((layer2_outputs(2268)) and (layer2_outputs(1526)));
    outputs(2074) <= layer2_outputs(1502);
    outputs(2075) <= (layer2_outputs(130)) and not (layer2_outputs(1421));
    outputs(2076) <= layer2_outputs(1984);
    outputs(2077) <= not(layer2_outputs(411)) or (layer2_outputs(2292));
    outputs(2078) <= not((layer2_outputs(434)) or (layer2_outputs(208)));
    outputs(2079) <= (layer2_outputs(1849)) and (layer2_outputs(960));
    outputs(2080) <= not(layer2_outputs(1225));
    outputs(2081) <= not(layer2_outputs(686));
    outputs(2082) <= not(layer2_outputs(624));
    outputs(2083) <= not(layer2_outputs(506)) or (layer2_outputs(1064));
    outputs(2084) <= layer2_outputs(1701);
    outputs(2085) <= not(layer2_outputs(1363)) or (layer2_outputs(1804));
    outputs(2086) <= (layer2_outputs(638)) xor (layer2_outputs(2495));
    outputs(2087) <= not(layer2_outputs(1943));
    outputs(2088) <= not(layer2_outputs(2025));
    outputs(2089) <= (layer2_outputs(765)) xor (layer2_outputs(2497));
    outputs(2090) <= layer2_outputs(401);
    outputs(2091) <= not(layer2_outputs(1302));
    outputs(2092) <= not((layer2_outputs(421)) xor (layer2_outputs(554)));
    outputs(2093) <= layer2_outputs(1179);
    outputs(2094) <= not(layer2_outputs(739));
    outputs(2095) <= (layer2_outputs(1123)) and not (layer2_outputs(2553));
    outputs(2096) <= not((layer2_outputs(2185)) or (layer2_outputs(923)));
    outputs(2097) <= not(layer2_outputs(744)) or (layer2_outputs(1508));
    outputs(2098) <= not(layer2_outputs(1484));
    outputs(2099) <= (layer2_outputs(2147)) and not (layer2_outputs(2309));
    outputs(2100) <= not(layer2_outputs(1806));
    outputs(2101) <= not(layer2_outputs(1929));
    outputs(2102) <= layer2_outputs(1086);
    outputs(2103) <= layer2_outputs(1639);
    outputs(2104) <= (layer2_outputs(662)) and not (layer2_outputs(128));
    outputs(2105) <= layer2_outputs(794);
    outputs(2106) <= not(layer2_outputs(303));
    outputs(2107) <= not(layer2_outputs(2557));
    outputs(2108) <= layer2_outputs(1592);
    outputs(2109) <= not(layer2_outputs(174));
    outputs(2110) <= (layer2_outputs(469)) and not (layer2_outputs(1222));
    outputs(2111) <= layer2_outputs(1304);
    outputs(2112) <= (layer2_outputs(746)) and not (layer2_outputs(2157));
    outputs(2113) <= not((layer2_outputs(51)) or (layer2_outputs(1059)));
    outputs(2114) <= (layer2_outputs(1453)) or (layer2_outputs(397));
    outputs(2115) <= not(layer2_outputs(577)) or (layer2_outputs(1410));
    outputs(2116) <= layer2_outputs(1694);
    outputs(2117) <= layer2_outputs(1145);
    outputs(2118) <= layer2_outputs(775);
    outputs(2119) <= not(layer2_outputs(31));
    outputs(2120) <= not(layer2_outputs(1722));
    outputs(2121) <= not(layer2_outputs(759)) or (layer2_outputs(2135));
    outputs(2122) <= (layer2_outputs(954)) xor (layer2_outputs(1949));
    outputs(2123) <= not((layer2_outputs(2360)) xor (layer2_outputs(2312)));
    outputs(2124) <= (layer2_outputs(1296)) xor (layer2_outputs(1479));
    outputs(2125) <= not((layer2_outputs(1021)) or (layer2_outputs(477)));
    outputs(2126) <= layer2_outputs(2368);
    outputs(2127) <= (layer2_outputs(843)) and not (layer2_outputs(975));
    outputs(2128) <= not(layer2_outputs(1877));
    outputs(2129) <= layer2_outputs(2452);
    outputs(2130) <= not(layer2_outputs(758));
    outputs(2131) <= not(layer2_outputs(2145));
    outputs(2132) <= not(layer2_outputs(2146));
    outputs(2133) <= layer2_outputs(234);
    outputs(2134) <= layer2_outputs(64);
    outputs(2135) <= not(layer2_outputs(456));
    outputs(2136) <= (layer2_outputs(1920)) or (layer2_outputs(1446));
    outputs(2137) <= (layer2_outputs(168)) or (layer2_outputs(268));
    outputs(2138) <= not(layer2_outputs(1380));
    outputs(2139) <= (layer2_outputs(2539)) or (layer2_outputs(2103));
    outputs(2140) <= (layer2_outputs(1911)) and not (layer2_outputs(911));
    outputs(2141) <= (layer2_outputs(1104)) and not (layer2_outputs(2266));
    outputs(2142) <= (layer2_outputs(420)) or (layer2_outputs(1003));
    outputs(2143) <= (layer2_outputs(2354)) and (layer2_outputs(611));
    outputs(2144) <= not(layer2_outputs(399));
    outputs(2145) <= not(layer2_outputs(2165));
    outputs(2146) <= not(layer2_outputs(2183)) or (layer2_outputs(1226));
    outputs(2147) <= not(layer2_outputs(801)) or (layer2_outputs(2121));
    outputs(2148) <= (layer2_outputs(2034)) xor (layer2_outputs(1211));
    outputs(2149) <= layer2_outputs(2101);
    outputs(2150) <= layer2_outputs(536);
    outputs(2151) <= not(layer2_outputs(1915));
    outputs(2152) <= not(layer2_outputs(2326));
    outputs(2153) <= not(layer2_outputs(443));
    outputs(2154) <= layer2_outputs(606);
    outputs(2155) <= layer2_outputs(2452);
    outputs(2156) <= layer2_outputs(48);
    outputs(2157) <= not(layer2_outputs(103));
    outputs(2158) <= (layer2_outputs(1640)) and not (layer2_outputs(322));
    outputs(2159) <= not(layer2_outputs(1081)) or (layer2_outputs(1453));
    outputs(2160) <= not(layer2_outputs(1465));
    outputs(2161) <= not(layer2_outputs(210));
    outputs(2162) <= layer2_outputs(2368);
    outputs(2163) <= not((layer2_outputs(594)) and (layer2_outputs(426)));
    outputs(2164) <= not((layer2_outputs(1378)) xor (layer2_outputs(2027)));
    outputs(2165) <= not(layer2_outputs(2029));
    outputs(2166) <= (layer2_outputs(0)) xor (layer2_outputs(2291));
    outputs(2167) <= (layer2_outputs(472)) and not (layer2_outputs(739));
    outputs(2168) <= not((layer2_outputs(2279)) or (layer2_outputs(2077)));
    outputs(2169) <= (layer2_outputs(1791)) and (layer2_outputs(410));
    outputs(2170) <= (layer2_outputs(590)) or (layer2_outputs(1638));
    outputs(2171) <= (layer2_outputs(406)) and not (layer2_outputs(907));
    outputs(2172) <= layer2_outputs(267);
    outputs(2173) <= not(layer2_outputs(164));
    outputs(2174) <= (layer2_outputs(1373)) and not (layer2_outputs(646));
    outputs(2175) <= not((layer2_outputs(1403)) or (layer2_outputs(2236)));
    outputs(2176) <= not(layer2_outputs(106)) or (layer2_outputs(1808));
    outputs(2177) <= (layer2_outputs(1849)) and not (layer2_outputs(980));
    outputs(2178) <= layer2_outputs(591);
    outputs(2179) <= (layer2_outputs(2536)) and (layer2_outputs(765));
    outputs(2180) <= layer2_outputs(266);
    outputs(2181) <= not(layer2_outputs(1842));
    outputs(2182) <= (layer2_outputs(1996)) xor (layer2_outputs(2337));
    outputs(2183) <= layer2_outputs(2336);
    outputs(2184) <= not(layer2_outputs(1933));
    outputs(2185) <= layer2_outputs(1112);
    outputs(2186) <= (layer2_outputs(977)) or (layer2_outputs(2120));
    outputs(2187) <= not(layer2_outputs(2159));
    outputs(2188) <= not(layer2_outputs(756));
    outputs(2189) <= not(layer2_outputs(1324));
    outputs(2190) <= (layer2_outputs(2121)) or (layer2_outputs(969));
    outputs(2191) <= (layer2_outputs(2172)) and not (layer2_outputs(1933));
    outputs(2192) <= (layer2_outputs(1078)) and not (layer2_outputs(841));
    outputs(2193) <= not((layer2_outputs(1716)) or (layer2_outputs(1553)));
    outputs(2194) <= not(layer2_outputs(127));
    outputs(2195) <= not(layer2_outputs(1749));
    outputs(2196) <= (layer2_outputs(2069)) and (layer2_outputs(1013));
    outputs(2197) <= not((layer2_outputs(2550)) or (layer2_outputs(99)));
    outputs(2198) <= layer2_outputs(1521);
    outputs(2199) <= not(layer2_outputs(1878));
    outputs(2200) <= (layer2_outputs(891)) and not (layer2_outputs(710));
    outputs(2201) <= not((layer2_outputs(1139)) xor (layer2_outputs(1936)));
    outputs(2202) <= (layer2_outputs(1916)) and not (layer2_outputs(1993));
    outputs(2203) <= not(layer2_outputs(1285));
    outputs(2204) <= not(layer2_outputs(2029));
    outputs(2205) <= not(layer2_outputs(391));
    outputs(2206) <= not((layer2_outputs(428)) xor (layer2_outputs(304)));
    outputs(2207) <= not(layer2_outputs(468));
    outputs(2208) <= (layer2_outputs(979)) xor (layer2_outputs(2035));
    outputs(2209) <= not((layer2_outputs(751)) and (layer2_outputs(1011)));
    outputs(2210) <= (layer2_outputs(1264)) xor (layer2_outputs(1283));
    outputs(2211) <= not(layer2_outputs(2301)) or (layer2_outputs(1176));
    outputs(2212) <= (layer2_outputs(1685)) and (layer2_outputs(1343));
    outputs(2213) <= layer2_outputs(856);
    outputs(2214) <= layer2_outputs(971);
    outputs(2215) <= layer2_outputs(590);
    outputs(2216) <= (layer2_outputs(895)) and not (layer2_outputs(725));
    outputs(2217) <= not(layer2_outputs(1263));
    outputs(2218) <= not((layer2_outputs(1963)) or (layer2_outputs(2428)));
    outputs(2219) <= layer2_outputs(332);
    outputs(2220) <= not(layer2_outputs(632)) or (layer2_outputs(1306));
    outputs(2221) <= (layer2_outputs(63)) and not (layer2_outputs(2450));
    outputs(2222) <= not((layer2_outputs(1843)) xor (layer2_outputs(1352)));
    outputs(2223) <= (layer2_outputs(1025)) and not (layer2_outputs(1773));
    outputs(2224) <= not(layer2_outputs(744));
    outputs(2225) <= not(layer2_outputs(2308));
    outputs(2226) <= layer2_outputs(1082);
    outputs(2227) <= (layer2_outputs(2015)) and (layer2_outputs(1255));
    outputs(2228) <= not(layer2_outputs(534));
    outputs(2229) <= (layer2_outputs(961)) and not (layer2_outputs(1981));
    outputs(2230) <= (layer2_outputs(894)) or (layer2_outputs(1695));
    outputs(2231) <= not(layer2_outputs(171));
    outputs(2232) <= not(layer2_outputs(1860));
    outputs(2233) <= not((layer2_outputs(2359)) xor (layer2_outputs(1708)));
    outputs(2234) <= not((layer2_outputs(1219)) xor (layer2_outputs(1017)));
    outputs(2235) <= (layer2_outputs(2142)) and not (layer2_outputs(1321));
    outputs(2236) <= (layer2_outputs(1657)) or (layer2_outputs(1317));
    outputs(2237) <= not((layer2_outputs(1677)) or (layer2_outputs(2364)));
    outputs(2238) <= not(layer2_outputs(2086));
    outputs(2239) <= (layer2_outputs(1802)) and not (layer2_outputs(1351));
    outputs(2240) <= not(layer2_outputs(227)) or (layer2_outputs(2110));
    outputs(2241) <= not(layer2_outputs(1222));
    outputs(2242) <= not(layer2_outputs(2342));
    outputs(2243) <= (layer2_outputs(1610)) xor (layer2_outputs(298));
    outputs(2244) <= not(layer2_outputs(1669));
    outputs(2245) <= not(layer2_outputs(76)) or (layer2_outputs(219));
    outputs(2246) <= not((layer2_outputs(1329)) or (layer2_outputs(2108)));
    outputs(2247) <= not(layer2_outputs(1712));
    outputs(2248) <= not((layer2_outputs(2508)) and (layer2_outputs(570)));
    outputs(2249) <= not(layer2_outputs(1126));
    outputs(2250) <= not(layer2_outputs(2429));
    outputs(2251) <= not(layer2_outputs(1569));
    outputs(2252) <= layer2_outputs(1625);
    outputs(2253) <= (layer2_outputs(1137)) and not (layer2_outputs(1224));
    outputs(2254) <= not((layer2_outputs(2347)) or (layer2_outputs(769)));
    outputs(2255) <= layer2_outputs(1464);
    outputs(2256) <= not(layer2_outputs(1895));
    outputs(2257) <= not(layer2_outputs(2405));
    outputs(2258) <= layer2_outputs(465);
    outputs(2259) <= not((layer2_outputs(344)) xor (layer2_outputs(643)));
    outputs(2260) <= not(layer2_outputs(956));
    outputs(2261) <= layer2_outputs(1295);
    outputs(2262) <= layer2_outputs(1180);
    outputs(2263) <= not((layer2_outputs(1294)) and (layer2_outputs(1818)));
    outputs(2264) <= layer2_outputs(1602);
    outputs(2265) <= layer2_outputs(1918);
    outputs(2266) <= layer2_outputs(2219);
    outputs(2267) <= not(layer2_outputs(1779));
    outputs(2268) <= layer2_outputs(650);
    outputs(2269) <= (layer2_outputs(737)) or (layer2_outputs(2400));
    outputs(2270) <= layer2_outputs(101);
    outputs(2271) <= (layer2_outputs(1367)) and not (layer2_outputs(2102));
    outputs(2272) <= not((layer2_outputs(413)) xor (layer2_outputs(407)));
    outputs(2273) <= not(layer2_outputs(1626)) or (layer2_outputs(2174));
    outputs(2274) <= layer2_outputs(2544);
    outputs(2275) <= layer2_outputs(1176);
    outputs(2276) <= not(layer2_outputs(1712));
    outputs(2277) <= (layer2_outputs(2061)) and not (layer2_outputs(1575));
    outputs(2278) <= not((layer2_outputs(2347)) or (layer2_outputs(2455)));
    outputs(2279) <= not(layer2_outputs(423));
    outputs(2280) <= not((layer2_outputs(471)) xor (layer2_outputs(1599)));
    outputs(2281) <= layer2_outputs(2313);
    outputs(2282) <= layer2_outputs(969);
    outputs(2283) <= not(layer2_outputs(1867));
    outputs(2284) <= (layer2_outputs(66)) and (layer2_outputs(1658));
    outputs(2285) <= not(layer2_outputs(670));
    outputs(2286) <= (layer2_outputs(8)) and not (layer2_outputs(1284));
    outputs(2287) <= (layer2_outputs(2380)) xor (layer2_outputs(502));
    outputs(2288) <= layer2_outputs(1071);
    outputs(2289) <= not(layer2_outputs(2300));
    outputs(2290) <= (layer2_outputs(1117)) or (layer2_outputs(1273));
    outputs(2291) <= not(layer2_outputs(1697));
    outputs(2292) <= not(layer2_outputs(888));
    outputs(2293) <= (layer2_outputs(1576)) and (layer2_outputs(1470));
    outputs(2294) <= (layer2_outputs(853)) and not (layer2_outputs(2394));
    outputs(2295) <= (layer2_outputs(2059)) and not (layer2_outputs(1285));
    outputs(2296) <= not(layer2_outputs(485));
    outputs(2297) <= not((layer2_outputs(1110)) or (layer2_outputs(677)));
    outputs(2298) <= (layer2_outputs(442)) xor (layer2_outputs(871));
    outputs(2299) <= not((layer2_outputs(987)) or (layer2_outputs(1619)));
    outputs(2300) <= not(layer2_outputs(1187));
    outputs(2301) <= (layer2_outputs(1474)) and (layer2_outputs(2555));
    outputs(2302) <= (layer2_outputs(264)) and (layer2_outputs(1798));
    outputs(2303) <= not(layer2_outputs(244));
    outputs(2304) <= (layer2_outputs(566)) and not (layer2_outputs(459));
    outputs(2305) <= not((layer2_outputs(474)) or (layer2_outputs(1678)));
    outputs(2306) <= layer2_outputs(1865);
    outputs(2307) <= (layer2_outputs(339)) xor (layer2_outputs(1797));
    outputs(2308) <= layer2_outputs(1776);
    outputs(2309) <= (layer2_outputs(2056)) and not (layer2_outputs(1290));
    outputs(2310) <= layer2_outputs(226);
    outputs(2311) <= layer2_outputs(795);
    outputs(2312) <= not(layer2_outputs(1173)) or (layer2_outputs(2296));
    outputs(2313) <= not((layer2_outputs(1686)) or (layer2_outputs(2293)));
    outputs(2314) <= not((layer2_outputs(559)) and (layer2_outputs(235)));
    outputs(2315) <= not(layer2_outputs(2559));
    outputs(2316) <= not(layer2_outputs(82));
    outputs(2317) <= layer2_outputs(1442);
    outputs(2318) <= layer2_outputs(2362);
    outputs(2319) <= layer2_outputs(2516);
    outputs(2320) <= (layer2_outputs(1647)) and not (layer2_outputs(1455));
    outputs(2321) <= not((layer2_outputs(1665)) or (layer2_outputs(1190)));
    outputs(2322) <= not(layer2_outputs(1520));
    outputs(2323) <= (layer2_outputs(1999)) and (layer2_outputs(492));
    outputs(2324) <= not(layer2_outputs(27));
    outputs(2325) <= not(layer2_outputs(2433));
    outputs(2326) <= not(layer2_outputs(2097));
    outputs(2327) <= not((layer2_outputs(445)) or (layer2_outputs(2463)));
    outputs(2328) <= not(layer2_outputs(1450)) or (layer2_outputs(2150));
    outputs(2329) <= layer2_outputs(290);
    outputs(2330) <= not(layer2_outputs(2530));
    outputs(2331) <= (layer2_outputs(566)) and (layer2_outputs(779));
    outputs(2332) <= (layer2_outputs(1743)) and not (layer2_outputs(644));
    outputs(2333) <= not(layer2_outputs(2524)) or (layer2_outputs(1364));
    outputs(2334) <= not(layer2_outputs(1789));
    outputs(2335) <= (layer2_outputs(1659)) and not (layer2_outputs(743));
    outputs(2336) <= not(layer2_outputs(100));
    outputs(2337) <= (layer2_outputs(1729)) and (layer2_outputs(2350));
    outputs(2338) <= layer2_outputs(349);
    outputs(2339) <= not(layer2_outputs(1208));
    outputs(2340) <= layer2_outputs(1914);
    outputs(2341) <= layer2_outputs(2386);
    outputs(2342) <= (layer2_outputs(35)) xor (layer2_outputs(1742));
    outputs(2343) <= (layer2_outputs(1996)) and (layer2_outputs(65));
    outputs(2344) <= not((layer2_outputs(2152)) or (layer2_outputs(33)));
    outputs(2345) <= not((layer2_outputs(432)) or (layer2_outputs(285)));
    outputs(2346) <= (layer2_outputs(2036)) and not (layer2_outputs(2214));
    outputs(2347) <= (layer2_outputs(2222)) and not (layer2_outputs(561));
    outputs(2348) <= (layer2_outputs(2079)) and (layer2_outputs(821));
    outputs(2349) <= (layer2_outputs(2229)) and (layer2_outputs(2280));
    outputs(2350) <= not(layer2_outputs(984));
    outputs(2351) <= not((layer2_outputs(806)) xor (layer2_outputs(428)));
    outputs(2352) <= (layer2_outputs(2162)) and not (layer2_outputs(609));
    outputs(2353) <= not(layer2_outputs(478));
    outputs(2354) <= (layer2_outputs(224)) and not (layer2_outputs(1304));
    outputs(2355) <= not((layer2_outputs(511)) or (layer2_outputs(1422)));
    outputs(2356) <= not(layer2_outputs(2339));
    outputs(2357) <= layer2_outputs(1731);
    outputs(2358) <= (layer2_outputs(1955)) xor (layer2_outputs(452));
    outputs(2359) <= not(layer2_outputs(575));
    outputs(2360) <= (layer2_outputs(2467)) and (layer2_outputs(28));
    outputs(2361) <= not((layer2_outputs(1301)) or (layer2_outputs(807)));
    outputs(2362) <= not(layer2_outputs(200));
    outputs(2363) <= layer2_outputs(2521);
    outputs(2364) <= not(layer2_outputs(816));
    outputs(2365) <= not(layer2_outputs(1495));
    outputs(2366) <= not(layer2_outputs(726));
    outputs(2367) <= not(layer2_outputs(2138));
    outputs(2368) <= not(layer2_outputs(1588));
    outputs(2369) <= layer2_outputs(1115);
    outputs(2370) <= not((layer2_outputs(1198)) or (layer2_outputs(56)));
    outputs(2371) <= (layer2_outputs(769)) and not (layer2_outputs(1413));
    outputs(2372) <= (layer2_outputs(1095)) and not (layer2_outputs(1477));
    outputs(2373) <= (layer2_outputs(510)) and not (layer2_outputs(677));
    outputs(2374) <= layer2_outputs(2382);
    outputs(2375) <= (layer2_outputs(112)) and (layer2_outputs(835));
    outputs(2376) <= layer2_outputs(1503);
    outputs(2377) <= (layer2_outputs(1379)) and not (layer2_outputs(1208));
    outputs(2378) <= not((layer2_outputs(1932)) or (layer2_outputs(2058)));
    outputs(2379) <= (layer2_outputs(1089)) xor (layer2_outputs(2132));
    outputs(2380) <= not(layer2_outputs(2005));
    outputs(2381) <= layer2_outputs(693);
    outputs(2382) <= not(layer2_outputs(2378));
    outputs(2383) <= layer2_outputs(577);
    outputs(2384) <= not(layer2_outputs(878));
    outputs(2385) <= layer2_outputs(224);
    outputs(2386) <= not((layer2_outputs(745)) xor (layer2_outputs(7)));
    outputs(2387) <= not(layer2_outputs(2514));
    outputs(2388) <= not(layer2_outputs(540)) or (layer2_outputs(1509));
    outputs(2389) <= not((layer2_outputs(2109)) or (layer2_outputs(1185)));
    outputs(2390) <= (layer2_outputs(626)) and (layer2_outputs(1714));
    outputs(2391) <= not(layer2_outputs(631));
    outputs(2392) <= (layer2_outputs(1035)) and not (layer2_outputs(887));
    outputs(2393) <= not(layer2_outputs(1598));
    outputs(2394) <= (layer2_outputs(1008)) and not (layer2_outputs(1950));
    outputs(2395) <= not(layer2_outputs(431)) or (layer2_outputs(400));
    outputs(2396) <= not(layer2_outputs(1261));
    outputs(2397) <= not((layer2_outputs(2146)) or (layer2_outputs(2071)));
    outputs(2398) <= (layer2_outputs(1762)) and (layer2_outputs(1091));
    outputs(2399) <= layer2_outputs(1930);
    outputs(2400) <= not(layer2_outputs(1606)) or (layer2_outputs(1897));
    outputs(2401) <= not(layer2_outputs(2530));
    outputs(2402) <= (layer2_outputs(1028)) and (layer2_outputs(83));
    outputs(2403) <= (layer2_outputs(2154)) and not (layer2_outputs(1959));
    outputs(2404) <= not((layer2_outputs(1699)) or (layer2_outputs(1645)));
    outputs(2405) <= not(layer2_outputs(84));
    outputs(2406) <= layer2_outputs(299);
    outputs(2407) <= not((layer2_outputs(698)) and (layer2_outputs(2310)));
    outputs(2408) <= not((layer2_outputs(787)) or (layer2_outputs(407)));
    outputs(2409) <= not(layer2_outputs(1800));
    outputs(2410) <= not((layer2_outputs(1267)) or (layer2_outputs(87)));
    outputs(2411) <= layer2_outputs(1342);
    outputs(2412) <= not((layer2_outputs(1420)) or (layer2_outputs(1581)));
    outputs(2413) <= not(layer2_outputs(851));
    outputs(2414) <= layer2_outputs(655);
    outputs(2415) <= not(layer2_outputs(1569)) or (layer2_outputs(2489));
    outputs(2416) <= not(layer2_outputs(2434));
    outputs(2417) <= layer2_outputs(2111);
    outputs(2418) <= not((layer2_outputs(417)) or (layer2_outputs(1026)));
    outputs(2419) <= not(layer2_outputs(2265));
    outputs(2420) <= not((layer2_outputs(1403)) or (layer2_outputs(478)));
    outputs(2421) <= not(layer2_outputs(705));
    outputs(2422) <= (layer2_outputs(25)) and not (layer2_outputs(2455));
    outputs(2423) <= layer2_outputs(2226);
    outputs(2424) <= layer2_outputs(381);
    outputs(2425) <= not(layer2_outputs(1548));
    outputs(2426) <= not((layer2_outputs(824)) xor (layer2_outputs(1472)));
    outputs(2427) <= (layer2_outputs(2055)) xor (layer2_outputs(699));
    outputs(2428) <= (layer2_outputs(112)) and (layer2_outputs(214));
    outputs(2429) <= not((layer2_outputs(2290)) or (layer2_outputs(639)));
    outputs(2430) <= not(layer2_outputs(2271));
    outputs(2431) <= layer2_outputs(633);
    outputs(2432) <= layer2_outputs(682);
    outputs(2433) <= layer2_outputs(1974);
    outputs(2434) <= not(layer2_outputs(126));
    outputs(2435) <= (layer2_outputs(2466)) and not (layer2_outputs(2054));
    outputs(2436) <= layer2_outputs(1958);
    outputs(2437) <= layer2_outputs(2072);
    outputs(2438) <= not((layer2_outputs(1332)) or (layer2_outputs(2190)));
    outputs(2439) <= layer2_outputs(404);
    outputs(2440) <= not(layer2_outputs(2241));
    outputs(2441) <= layer2_outputs(1319);
    outputs(2442) <= (layer2_outputs(58)) and not (layer2_outputs(589));
    outputs(2443) <= not(layer2_outputs(1270));
    outputs(2444) <= layer2_outputs(119);
    outputs(2445) <= (layer2_outputs(636)) and (layer2_outputs(1229));
    outputs(2446) <= not(layer2_outputs(990));
    outputs(2447) <= (layer2_outputs(2129)) and not (layer2_outputs(285));
    outputs(2448) <= not(layer2_outputs(294));
    outputs(2449) <= (layer2_outputs(472)) and not (layer2_outputs(417));
    outputs(2450) <= not(layer2_outputs(183)) or (layer2_outputs(1611));
    outputs(2451) <= (layer2_outputs(2127)) and not (layer2_outputs(2234));
    outputs(2452) <= layer2_outputs(2036);
    outputs(2453) <= not(layer2_outputs(1293));
    outputs(2454) <= not(layer2_outputs(1557));
    outputs(2455) <= not(layer2_outputs(1430));
    outputs(2456) <= layer2_outputs(228);
    outputs(2457) <= (layer2_outputs(1601)) and not (layer2_outputs(1410));
    outputs(2458) <= not(layer2_outputs(1506));
    outputs(2459) <= layer2_outputs(1787);
    outputs(2460) <= not((layer2_outputs(499)) or (layer2_outputs(342)));
    outputs(2461) <= not(layer2_outputs(454));
    outputs(2462) <= layer2_outputs(1300);
    outputs(2463) <= not((layer2_outputs(482)) or (layer2_outputs(536)));
    outputs(2464) <= not(layer2_outputs(2433));
    outputs(2465) <= (layer2_outputs(1587)) and not (layer2_outputs(2011));
    outputs(2466) <= layer2_outputs(1579);
    outputs(2467) <= (layer2_outputs(1316)) and not (layer2_outputs(529));
    outputs(2468) <= not((layer2_outputs(356)) or (layer2_outputs(2447)));
    outputs(2469) <= not(layer2_outputs(2503));
    outputs(2470) <= layer2_outputs(902);
    outputs(2471) <= not(layer2_outputs(2396)) or (layer2_outputs(2068));
    outputs(2472) <= (layer2_outputs(1571)) and (layer2_outputs(2443));
    outputs(2473) <= (layer2_outputs(361)) and (layer2_outputs(1889));
    outputs(2474) <= layer2_outputs(1738);
    outputs(2475) <= not((layer2_outputs(1747)) and (layer2_outputs(1277)));
    outputs(2476) <= (layer2_outputs(1317)) and (layer2_outputs(367));
    outputs(2477) <= (layer2_outputs(917)) and not (layer2_outputs(1505));
    outputs(2478) <= not((layer2_outputs(1746)) and (layer2_outputs(1959)));
    outputs(2479) <= (layer2_outputs(1490)) and not (layer2_outputs(2380));
    outputs(2480) <= not(layer2_outputs(370));
    outputs(2481) <= (layer2_outputs(1668)) and not (layer2_outputs(543));
    outputs(2482) <= layer2_outputs(1679);
    outputs(2483) <= not(layer2_outputs(191));
    outputs(2484) <= not(layer2_outputs(830));
    outputs(2485) <= layer2_outputs(919);
    outputs(2486) <= (layer2_outputs(1896)) and not (layer2_outputs(2252));
    outputs(2487) <= not(layer2_outputs(345));
    outputs(2488) <= layer2_outputs(1556);
    outputs(2489) <= (layer2_outputs(2107)) and not (layer2_outputs(1908));
    outputs(2490) <= layer2_outputs(434);
    outputs(2491) <= not(layer2_outputs(1055));
    outputs(2492) <= layer2_outputs(766);
    outputs(2493) <= not(layer2_outputs(2091));
    outputs(2494) <= not((layer2_outputs(38)) or (layer2_outputs(1224)));
    outputs(2495) <= (layer2_outputs(1974)) or (layer2_outputs(1087));
    outputs(2496) <= not(layer2_outputs(2243));
    outputs(2497) <= not((layer2_outputs(1169)) or (layer2_outputs(281)));
    outputs(2498) <= not(layer2_outputs(2210));
    outputs(2499) <= not((layer2_outputs(1700)) or (layer2_outputs(2160)));
    outputs(2500) <= not(layer2_outputs(913));
    outputs(2501) <= layer2_outputs(1714);
    outputs(2502) <= (layer2_outputs(484)) and not (layer2_outputs(849));
    outputs(2503) <= not(layer2_outputs(1588));
    outputs(2504) <= not(layer2_outputs(1335));
    outputs(2505) <= layer2_outputs(572);
    outputs(2506) <= layer2_outputs(857);
    outputs(2507) <= not(layer2_outputs(365));
    outputs(2508) <= not((layer2_outputs(889)) or (layer2_outputs(659)));
    outputs(2509) <= layer2_outputs(321);
    outputs(2510) <= (layer2_outputs(259)) and (layer2_outputs(1165));
    outputs(2511) <= not(layer2_outputs(1952));
    outputs(2512) <= layer2_outputs(2376);
    outputs(2513) <= not(layer2_outputs(172)) or (layer2_outputs(1891));
    outputs(2514) <= layer2_outputs(1958);
    outputs(2515) <= layer2_outputs(16);
    outputs(2516) <= layer2_outputs(2306);
    outputs(2517) <= layer2_outputs(1265);
    outputs(2518) <= (layer2_outputs(2013)) and not (layer2_outputs(2040));
    outputs(2519) <= not((layer2_outputs(1782)) and (layer2_outputs(722)));
    outputs(2520) <= not(layer2_outputs(749)) or (layer2_outputs(1711));
    outputs(2521) <= layer2_outputs(2066);
    outputs(2522) <= not(layer2_outputs(1332));
    outputs(2523) <= layer2_outputs(1496);
    outputs(2524) <= not(layer2_outputs(646));
    outputs(2525) <= (layer2_outputs(1074)) and (layer2_outputs(1754));
    outputs(2526) <= not(layer2_outputs(1591));
    outputs(2527) <= (layer2_outputs(1228)) xor (layer2_outputs(809));
    outputs(2528) <= layer2_outputs(1362);
    outputs(2529) <= (layer2_outputs(92)) and (layer2_outputs(48));
    outputs(2530) <= not(layer2_outputs(1143)) or (layer2_outputs(1129));
    outputs(2531) <= not(layer2_outputs(822));
    outputs(2532) <= (layer2_outputs(490)) and not (layer2_outputs(1821));
    outputs(2533) <= not((layer2_outputs(713)) or (layer2_outputs(2483)));
    outputs(2534) <= layer2_outputs(1766);
    outputs(2535) <= (layer2_outputs(1461)) and not (layer2_outputs(595));
    outputs(2536) <= (layer2_outputs(2013)) and (layer2_outputs(1633));
    outputs(2537) <= not(layer2_outputs(2305));
    outputs(2538) <= not((layer2_outputs(1657)) or (layer2_outputs(786)));
    outputs(2539) <= not(layer2_outputs(1042));
    outputs(2540) <= not(layer2_outputs(55));
    outputs(2541) <= (layer2_outputs(2170)) and (layer2_outputs(1531));
    outputs(2542) <= not(layer2_outputs(297));
    outputs(2543) <= layer2_outputs(2087);
    outputs(2544) <= (layer2_outputs(1289)) and not (layer2_outputs(1532));
    outputs(2545) <= (layer2_outputs(626)) and not (layer2_outputs(1610));
    outputs(2546) <= (layer2_outputs(2254)) and not (layer2_outputs(592));
    outputs(2547) <= not(layer2_outputs(1859));
    outputs(2548) <= not(layer2_outputs(679));
    outputs(2549) <= not(layer2_outputs(1261));
    outputs(2550) <= layer2_outputs(2196);
    outputs(2551) <= (layer2_outputs(1570)) and (layer2_outputs(861));
    outputs(2552) <= layer2_outputs(831);
    outputs(2553) <= (layer2_outputs(2194)) and not (layer2_outputs(829));
    outputs(2554) <= layer2_outputs(986);
    outputs(2555) <= not(layer2_outputs(1404));
    outputs(2556) <= not((layer2_outputs(525)) xor (layer2_outputs(1111)));
    outputs(2557) <= not(layer2_outputs(1557));
    outputs(2558) <= (layer2_outputs(2361)) or (layer2_outputs(2409));
    outputs(2559) <= (layer2_outputs(2195)) and not (layer2_outputs(2017));

end Behavioral;
