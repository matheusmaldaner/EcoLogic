library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(12799 downto 0);
    signal layer1_outputs: std_logic_vector(12799 downto 0);
    signal layer2_outputs: std_logic_vector(12799 downto 0);

begin
    layer0_outputs(0) <= a or b;
    layer0_outputs(1) <= b and not a;
    layer0_outputs(2) <= a or b;
    layer0_outputs(3) <= not (a or b);
    layer0_outputs(4) <= not (a or b);
    layer0_outputs(5) <= b and not a;
    layer0_outputs(6) <= a or b;
    layer0_outputs(7) <= a xor b;
    layer0_outputs(8) <= a or b;
    layer0_outputs(9) <= b and not a;
    layer0_outputs(10) <= a and not b;
    layer0_outputs(11) <= a xor b;
    layer0_outputs(12) <= not a;
    layer0_outputs(13) <= not (a or b);
    layer0_outputs(14) <= not (a or b);
    layer0_outputs(15) <= a and b;
    layer0_outputs(16) <= not b or a;
    layer0_outputs(17) <= b and not a;
    layer0_outputs(18) <= not (a and b);
    layer0_outputs(19) <= b and not a;
    layer0_outputs(20) <= not b or a;
    layer0_outputs(21) <= not (a or b);
    layer0_outputs(22) <= a or b;
    layer0_outputs(23) <= not a or b;
    layer0_outputs(24) <= not a or b;
    layer0_outputs(25) <= not a or b;
    layer0_outputs(26) <= a and not b;
    layer0_outputs(27) <= not b;
    layer0_outputs(28) <= not b;
    layer0_outputs(29) <= not b;
    layer0_outputs(30) <= b and not a;
    layer0_outputs(31) <= b and not a;
    layer0_outputs(32) <= not (a xor b);
    layer0_outputs(33) <= a or b;
    layer0_outputs(34) <= b and not a;
    layer0_outputs(35) <= not (a xor b);
    layer0_outputs(36) <= b;
    layer0_outputs(37) <= a and b;
    layer0_outputs(38) <= a and not b;
    layer0_outputs(39) <= b;
    layer0_outputs(40) <= not b;
    layer0_outputs(41) <= not (a and b);
    layer0_outputs(42) <= not (a xor b);
    layer0_outputs(43) <= a;
    layer0_outputs(44) <= not (a xor b);
    layer0_outputs(45) <= not (a xor b);
    layer0_outputs(46) <= not (a xor b);
    layer0_outputs(47) <= b and not a;
    layer0_outputs(48) <= a and b;
    layer0_outputs(49) <= a;
    layer0_outputs(50) <= not b;
    layer0_outputs(51) <= a and not b;
    layer0_outputs(52) <= not (a or b);
    layer0_outputs(53) <= not (a xor b);
    layer0_outputs(54) <= a xor b;
    layer0_outputs(55) <= not b or a;
    layer0_outputs(56) <= b;
    layer0_outputs(57) <= not (a or b);
    layer0_outputs(58) <= a and b;
    layer0_outputs(59) <= b and not a;
    layer0_outputs(60) <= a or b;
    layer0_outputs(61) <= not a or b;
    layer0_outputs(62) <= a and b;
    layer0_outputs(63) <= 1'b0;
    layer0_outputs(64) <= a;
    layer0_outputs(65) <= not b or a;
    layer0_outputs(66) <= not (a or b);
    layer0_outputs(67) <= not a;
    layer0_outputs(68) <= a or b;
    layer0_outputs(69) <= a;
    layer0_outputs(70) <= a or b;
    layer0_outputs(71) <= not b or a;
    layer0_outputs(72) <= not (a xor b);
    layer0_outputs(73) <= a or b;
    layer0_outputs(74) <= a or b;
    layer0_outputs(75) <= not (a or b);
    layer0_outputs(76) <= b;
    layer0_outputs(77) <= not a or b;
    layer0_outputs(78) <= a or b;
    layer0_outputs(79) <= a xor b;
    layer0_outputs(80) <= not (a or b);
    layer0_outputs(81) <= a xor b;
    layer0_outputs(82) <= b;
    layer0_outputs(83) <= not a or b;
    layer0_outputs(84) <= not a;
    layer0_outputs(85) <= not b;
    layer0_outputs(86) <= not (a or b);
    layer0_outputs(87) <= not b or a;
    layer0_outputs(88) <= b;
    layer0_outputs(89) <= not b;
    layer0_outputs(90) <= a xor b;
    layer0_outputs(91) <= not a or b;
    layer0_outputs(92) <= not (a xor b);
    layer0_outputs(93) <= not b or a;
    layer0_outputs(94) <= b;
    layer0_outputs(95) <= not (a xor b);
    layer0_outputs(96) <= not (a xor b);
    layer0_outputs(97) <= not (a xor b);
    layer0_outputs(98) <= not a or b;
    layer0_outputs(99) <= not (a xor b);
    layer0_outputs(100) <= a;
    layer0_outputs(101) <= a and b;
    layer0_outputs(102) <= a or b;
    layer0_outputs(103) <= a;
    layer0_outputs(104) <= not (a xor b);
    layer0_outputs(105) <= a;
    layer0_outputs(106) <= a and b;
    layer0_outputs(107) <= a and not b;
    layer0_outputs(108) <= not a or b;
    layer0_outputs(109) <= a or b;
    layer0_outputs(110) <= a xor b;
    layer0_outputs(111) <= a and not b;
    layer0_outputs(112) <= not a or b;
    layer0_outputs(113) <= a xor b;
    layer0_outputs(114) <= a or b;
    layer0_outputs(115) <= b;
    layer0_outputs(116) <= a or b;
    layer0_outputs(117) <= a and b;
    layer0_outputs(118) <= 1'b1;
    layer0_outputs(119) <= not (a xor b);
    layer0_outputs(120) <= not b;
    layer0_outputs(121) <= b and not a;
    layer0_outputs(122) <= not a or b;
    layer0_outputs(123) <= a;
    layer0_outputs(124) <= a or b;
    layer0_outputs(125) <= not (a or b);
    layer0_outputs(126) <= a;
    layer0_outputs(127) <= a or b;
    layer0_outputs(128) <= not a;
    layer0_outputs(129) <= a;
    layer0_outputs(130) <= not b or a;
    layer0_outputs(131) <= not (a xor b);
    layer0_outputs(132) <= a;
    layer0_outputs(133) <= not (a xor b);
    layer0_outputs(134) <= not a;
    layer0_outputs(135) <= a;
    layer0_outputs(136) <= a;
    layer0_outputs(137) <= b;
    layer0_outputs(138) <= not (a or b);
    layer0_outputs(139) <= not (a or b);
    layer0_outputs(140) <= b and not a;
    layer0_outputs(141) <= not (a or b);
    layer0_outputs(142) <= a xor b;
    layer0_outputs(143) <= 1'b1;
    layer0_outputs(144) <= not b or a;
    layer0_outputs(145) <= a and not b;
    layer0_outputs(146) <= not (a or b);
    layer0_outputs(147) <= not a or b;
    layer0_outputs(148) <= a and b;
    layer0_outputs(149) <= not a;
    layer0_outputs(150) <= not (a or b);
    layer0_outputs(151) <= a or b;
    layer0_outputs(152) <= not b or a;
    layer0_outputs(153) <= a and not b;
    layer0_outputs(154) <= not (a xor b);
    layer0_outputs(155) <= 1'b0;
    layer0_outputs(156) <= b and not a;
    layer0_outputs(157) <= not (a or b);
    layer0_outputs(158) <= not (a or b);
    layer0_outputs(159) <= not (a xor b);
    layer0_outputs(160) <= not b;
    layer0_outputs(161) <= a or b;
    layer0_outputs(162) <= a or b;
    layer0_outputs(163) <= a and not b;
    layer0_outputs(164) <= not b or a;
    layer0_outputs(165) <= b;
    layer0_outputs(166) <= a or b;
    layer0_outputs(167) <= a;
    layer0_outputs(168) <= b;
    layer0_outputs(169) <= not b;
    layer0_outputs(170) <= a and b;
    layer0_outputs(171) <= not (a or b);
    layer0_outputs(172) <= not a;
    layer0_outputs(173) <= not a;
    layer0_outputs(174) <= a or b;
    layer0_outputs(175) <= not (a xor b);
    layer0_outputs(176) <= not (a and b);
    layer0_outputs(177) <= a;
    layer0_outputs(178) <= b and not a;
    layer0_outputs(179) <= not (a and b);
    layer0_outputs(180) <= a;
    layer0_outputs(181) <= a or b;
    layer0_outputs(182) <= a or b;
    layer0_outputs(183) <= a or b;
    layer0_outputs(184) <= a or b;
    layer0_outputs(185) <= a xor b;
    layer0_outputs(186) <= not (a or b);
    layer0_outputs(187) <= a xor b;
    layer0_outputs(188) <= not b or a;
    layer0_outputs(189) <= a;
    layer0_outputs(190) <= not (a or b);
    layer0_outputs(191) <= not b or a;
    layer0_outputs(192) <= not a or b;
    layer0_outputs(193) <= 1'b0;
    layer0_outputs(194) <= b and not a;
    layer0_outputs(195) <= not a;
    layer0_outputs(196) <= not a or b;
    layer0_outputs(197) <= not a;
    layer0_outputs(198) <= a and not b;
    layer0_outputs(199) <= 1'b0;
    layer0_outputs(200) <= a xor b;
    layer0_outputs(201) <= not b;
    layer0_outputs(202) <= not (a or b);
    layer0_outputs(203) <= not (a and b);
    layer0_outputs(204) <= not (a or b);
    layer0_outputs(205) <= a or b;
    layer0_outputs(206) <= a;
    layer0_outputs(207) <= not a or b;
    layer0_outputs(208) <= not b;
    layer0_outputs(209) <= not (a or b);
    layer0_outputs(210) <= not a;
    layer0_outputs(211) <= not b;
    layer0_outputs(212) <= not b or a;
    layer0_outputs(213) <= b;
    layer0_outputs(214) <= b and not a;
    layer0_outputs(215) <= b and not a;
    layer0_outputs(216) <= a and not b;
    layer0_outputs(217) <= a or b;
    layer0_outputs(218) <= not (a or b);
    layer0_outputs(219) <= not (a or b);
    layer0_outputs(220) <= not b;
    layer0_outputs(221) <= 1'b0;
    layer0_outputs(222) <= not (a xor b);
    layer0_outputs(223) <= not b or a;
    layer0_outputs(224) <= 1'b0;
    layer0_outputs(225) <= not (a xor b);
    layer0_outputs(226) <= not (a or b);
    layer0_outputs(227) <= a or b;
    layer0_outputs(228) <= not a;
    layer0_outputs(229) <= not (a or b);
    layer0_outputs(230) <= not b;
    layer0_outputs(231) <= not (a or b);
    layer0_outputs(232) <= b and not a;
    layer0_outputs(233) <= b;
    layer0_outputs(234) <= a and b;
    layer0_outputs(235) <= a and not b;
    layer0_outputs(236) <= a and b;
    layer0_outputs(237) <= b and not a;
    layer0_outputs(238) <= 1'b0;
    layer0_outputs(239) <= not (a or b);
    layer0_outputs(240) <= 1'b0;
    layer0_outputs(241) <= not a;
    layer0_outputs(242) <= b and not a;
    layer0_outputs(243) <= a;
    layer0_outputs(244) <= b and not a;
    layer0_outputs(245) <= not b or a;
    layer0_outputs(246) <= a and not b;
    layer0_outputs(247) <= b and not a;
    layer0_outputs(248) <= a;
    layer0_outputs(249) <= not a;
    layer0_outputs(250) <= not b;
    layer0_outputs(251) <= a;
    layer0_outputs(252) <= not a;
    layer0_outputs(253) <= a;
    layer0_outputs(254) <= a or b;
    layer0_outputs(255) <= not (a and b);
    layer0_outputs(256) <= a xor b;
    layer0_outputs(257) <= not b;
    layer0_outputs(258) <= not (a or b);
    layer0_outputs(259) <= not b or a;
    layer0_outputs(260) <= not a or b;
    layer0_outputs(261) <= not (a or b);
    layer0_outputs(262) <= a and not b;
    layer0_outputs(263) <= not a;
    layer0_outputs(264) <= a or b;
    layer0_outputs(265) <= not (a xor b);
    layer0_outputs(266) <= not (a or b);
    layer0_outputs(267) <= b;
    layer0_outputs(268) <= not a;
    layer0_outputs(269) <= 1'b1;
    layer0_outputs(270) <= a;
    layer0_outputs(271) <= not (a and b);
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= not (a or b);
    layer0_outputs(274) <= not b or a;
    layer0_outputs(275) <= a or b;
    layer0_outputs(276) <= b and not a;
    layer0_outputs(277) <= 1'b1;
    layer0_outputs(278) <= b;
    layer0_outputs(279) <= not b or a;
    layer0_outputs(280) <= not (a or b);
    layer0_outputs(281) <= b;
    layer0_outputs(282) <= not a or b;
    layer0_outputs(283) <= not b or a;
    layer0_outputs(284) <= a;
    layer0_outputs(285) <= not (a and b);
    layer0_outputs(286) <= not a;
    layer0_outputs(287) <= a or b;
    layer0_outputs(288) <= b;
    layer0_outputs(289) <= a or b;
    layer0_outputs(290) <= a xor b;
    layer0_outputs(291) <= not a;
    layer0_outputs(292) <= a;
    layer0_outputs(293) <= a xor b;
    layer0_outputs(294) <= a xor b;
    layer0_outputs(295) <= not b;
    layer0_outputs(296) <= not a or b;
    layer0_outputs(297) <= not (a or b);
    layer0_outputs(298) <= not b;
    layer0_outputs(299) <= a or b;
    layer0_outputs(300) <= a or b;
    layer0_outputs(301) <= a and b;
    layer0_outputs(302) <= not a;
    layer0_outputs(303) <= not a;
    layer0_outputs(304) <= not b or a;
    layer0_outputs(305) <= a xor b;
    layer0_outputs(306) <= not (a xor b);
    layer0_outputs(307) <= not b or a;
    layer0_outputs(308) <= a and not b;
    layer0_outputs(309) <= not a;
    layer0_outputs(310) <= b;
    layer0_outputs(311) <= not b;
    layer0_outputs(312) <= b and not a;
    layer0_outputs(313) <= a or b;
    layer0_outputs(314) <= not (a and b);
    layer0_outputs(315) <= 1'b0;
    layer0_outputs(316) <= a or b;
    layer0_outputs(317) <= not b or a;
    layer0_outputs(318) <= not b;
    layer0_outputs(319) <= not a;
    layer0_outputs(320) <= not b;
    layer0_outputs(321) <= not a;
    layer0_outputs(322) <= not a or b;
    layer0_outputs(323) <= b;
    layer0_outputs(324) <= not a or b;
    layer0_outputs(325) <= a and not b;
    layer0_outputs(326) <= not a or b;
    layer0_outputs(327) <= not a;
    layer0_outputs(328) <= not b or a;
    layer0_outputs(329) <= not a or b;
    layer0_outputs(330) <= b and not a;
    layer0_outputs(331) <= b;
    layer0_outputs(332) <= a or b;
    layer0_outputs(333) <= a or b;
    layer0_outputs(334) <= not a;
    layer0_outputs(335) <= not a;
    layer0_outputs(336) <= 1'b0;
    layer0_outputs(337) <= a or b;
    layer0_outputs(338) <= not a;
    layer0_outputs(339) <= not (a or b);
    layer0_outputs(340) <= not b or a;
    layer0_outputs(341) <= not b or a;
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= a and not b;
    layer0_outputs(344) <= a xor b;
    layer0_outputs(345) <= a and not b;
    layer0_outputs(346) <= not a or b;
    layer0_outputs(347) <= not (a xor b);
    layer0_outputs(348) <= not (a or b);
    layer0_outputs(349) <= b;
    layer0_outputs(350) <= a;
    layer0_outputs(351) <= not b;
    layer0_outputs(352) <= a xor b;
    layer0_outputs(353) <= a or b;
    layer0_outputs(354) <= not a or b;
    layer0_outputs(355) <= not (a or b);
    layer0_outputs(356) <= not b or a;
    layer0_outputs(357) <= not (a or b);
    layer0_outputs(358) <= a or b;
    layer0_outputs(359) <= b and not a;
    layer0_outputs(360) <= not (a xor b);
    layer0_outputs(361) <= not (a xor b);
    layer0_outputs(362) <= a and b;
    layer0_outputs(363) <= b and not a;
    layer0_outputs(364) <= a;
    layer0_outputs(365) <= 1'b0;
    layer0_outputs(366) <= b;
    layer0_outputs(367) <= not a;
    layer0_outputs(368) <= a or b;
    layer0_outputs(369) <= a xor b;
    layer0_outputs(370) <= a and not b;
    layer0_outputs(371) <= a or b;
    layer0_outputs(372) <= not (a and b);
    layer0_outputs(373) <= not (a and b);
    layer0_outputs(374) <= not (a or b);
    layer0_outputs(375) <= b;
    layer0_outputs(376) <= a xor b;
    layer0_outputs(377) <= not a;
    layer0_outputs(378) <= not (a or b);
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= not a;
    layer0_outputs(381) <= b;
    layer0_outputs(382) <= not a;
    layer0_outputs(383) <= not b or a;
    layer0_outputs(384) <= not (a xor b);
    layer0_outputs(385) <= a;
    layer0_outputs(386) <= not a;
    layer0_outputs(387) <= not b or a;
    layer0_outputs(388) <= a xor b;
    layer0_outputs(389) <= not b or a;
    layer0_outputs(390) <= not a;
    layer0_outputs(391) <= a xor b;
    layer0_outputs(392) <= not b or a;
    layer0_outputs(393) <= not (a or b);
    layer0_outputs(394) <= b;
    layer0_outputs(395) <= a;
    layer0_outputs(396) <= not b or a;
    layer0_outputs(397) <= not (a or b);
    layer0_outputs(398) <= not (a or b);
    layer0_outputs(399) <= a and not b;
    layer0_outputs(400) <= a or b;
    layer0_outputs(401) <= a or b;
    layer0_outputs(402) <= a or b;
    layer0_outputs(403) <= b and not a;
    layer0_outputs(404) <= b;
    layer0_outputs(405) <= not b;
    layer0_outputs(406) <= b and not a;
    layer0_outputs(407) <= not b or a;
    layer0_outputs(408) <= a xor b;
    layer0_outputs(409) <= b and not a;
    layer0_outputs(410) <= a or b;
    layer0_outputs(411) <= not (a or b);
    layer0_outputs(412) <= b and not a;
    layer0_outputs(413) <= a;
    layer0_outputs(414) <= not (a and b);
    layer0_outputs(415) <= 1'b0;
    layer0_outputs(416) <= not b or a;
    layer0_outputs(417) <= not (a or b);
    layer0_outputs(418) <= a or b;
    layer0_outputs(419) <= a and not b;
    layer0_outputs(420) <= a xor b;
    layer0_outputs(421) <= not b;
    layer0_outputs(422) <= b;
    layer0_outputs(423) <= a xor b;
    layer0_outputs(424) <= a or b;
    layer0_outputs(425) <= a xor b;
    layer0_outputs(426) <= b and not a;
    layer0_outputs(427) <= 1'b1;
    layer0_outputs(428) <= b and not a;
    layer0_outputs(429) <= not b or a;
    layer0_outputs(430) <= b;
    layer0_outputs(431) <= a xor b;
    layer0_outputs(432) <= not (a xor b);
    layer0_outputs(433) <= a or b;
    layer0_outputs(434) <= not (a or b);
    layer0_outputs(435) <= not a;
    layer0_outputs(436) <= not (a and b);
    layer0_outputs(437) <= not b;
    layer0_outputs(438) <= not (a and b);
    layer0_outputs(439) <= a;
    layer0_outputs(440) <= a or b;
    layer0_outputs(441) <= b;
    layer0_outputs(442) <= a and not b;
    layer0_outputs(443) <= not a;
    layer0_outputs(444) <= not (a or b);
    layer0_outputs(445) <= a or b;
    layer0_outputs(446) <= b;
    layer0_outputs(447) <= a or b;
    layer0_outputs(448) <= a;
    layer0_outputs(449) <= not b;
    layer0_outputs(450) <= a and not b;
    layer0_outputs(451) <= not a;
    layer0_outputs(452) <= b and not a;
    layer0_outputs(453) <= not (a and b);
    layer0_outputs(454) <= a and b;
    layer0_outputs(455) <= a or b;
    layer0_outputs(456) <= not (a or b);
    layer0_outputs(457) <= 1'b1;
    layer0_outputs(458) <= a or b;
    layer0_outputs(459) <= a;
    layer0_outputs(460) <= b and not a;
    layer0_outputs(461) <= a or b;
    layer0_outputs(462) <= 1'b1;
    layer0_outputs(463) <= not a;
    layer0_outputs(464) <= 1'b1;
    layer0_outputs(465) <= not b or a;
    layer0_outputs(466) <= not a or b;
    layer0_outputs(467) <= b and not a;
    layer0_outputs(468) <= a;
    layer0_outputs(469) <= not (a and b);
    layer0_outputs(470) <= not b or a;
    layer0_outputs(471) <= a;
    layer0_outputs(472) <= a or b;
    layer0_outputs(473) <= not b;
    layer0_outputs(474) <= a and not b;
    layer0_outputs(475) <= a xor b;
    layer0_outputs(476) <= a or b;
    layer0_outputs(477) <= not b or a;
    layer0_outputs(478) <= not (a xor b);
    layer0_outputs(479) <= b;
    layer0_outputs(480) <= not b or a;
    layer0_outputs(481) <= not (a xor b);
    layer0_outputs(482) <= a xor b;
    layer0_outputs(483) <= b;
    layer0_outputs(484) <= not a;
    layer0_outputs(485) <= a or b;
    layer0_outputs(486) <= a xor b;
    layer0_outputs(487) <= a and not b;
    layer0_outputs(488) <= not a;
    layer0_outputs(489) <= not a;
    layer0_outputs(490) <= a xor b;
    layer0_outputs(491) <= not a;
    layer0_outputs(492) <= not a;
    layer0_outputs(493) <= a xor b;
    layer0_outputs(494) <= not b or a;
    layer0_outputs(495) <= b;
    layer0_outputs(496) <= b;
    layer0_outputs(497) <= a and b;
    layer0_outputs(498) <= a and not b;
    layer0_outputs(499) <= a xor b;
    layer0_outputs(500) <= not (a or b);
    layer0_outputs(501) <= a;
    layer0_outputs(502) <= 1'b1;
    layer0_outputs(503) <= b;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= not a;
    layer0_outputs(506) <= not b or a;
    layer0_outputs(507) <= a or b;
    layer0_outputs(508) <= not (a or b);
    layer0_outputs(509) <= not a or b;
    layer0_outputs(510) <= not b;
    layer0_outputs(511) <= 1'b1;
    layer0_outputs(512) <= a and b;
    layer0_outputs(513) <= not b;
    layer0_outputs(514) <= a and b;
    layer0_outputs(515) <= not (a xor b);
    layer0_outputs(516) <= a or b;
    layer0_outputs(517) <= a xor b;
    layer0_outputs(518) <= not a or b;
    layer0_outputs(519) <= not b or a;
    layer0_outputs(520) <= not (a or b);
    layer0_outputs(521) <= not b;
    layer0_outputs(522) <= not a;
    layer0_outputs(523) <= a xor b;
    layer0_outputs(524) <= a;
    layer0_outputs(525) <= a or b;
    layer0_outputs(526) <= not a;
    layer0_outputs(527) <= a;
    layer0_outputs(528) <= a or b;
    layer0_outputs(529) <= not a or b;
    layer0_outputs(530) <= not (a or b);
    layer0_outputs(531) <= not b;
    layer0_outputs(532) <= a;
    layer0_outputs(533) <= not b or a;
    layer0_outputs(534) <= b and not a;
    layer0_outputs(535) <= a or b;
    layer0_outputs(536) <= not b or a;
    layer0_outputs(537) <= not (a or b);
    layer0_outputs(538) <= a xor b;
    layer0_outputs(539) <= not (a or b);
    layer0_outputs(540) <= b and not a;
    layer0_outputs(541) <= not (a or b);
    layer0_outputs(542) <= not a;
    layer0_outputs(543) <= a and not b;
    layer0_outputs(544) <= not b;
    layer0_outputs(545) <= not b;
    layer0_outputs(546) <= a xor b;
    layer0_outputs(547) <= not (a or b);
    layer0_outputs(548) <= a and b;
    layer0_outputs(549) <= a or b;
    layer0_outputs(550) <= not a or b;
    layer0_outputs(551) <= not a or b;
    layer0_outputs(552) <= not (a or b);
    layer0_outputs(553) <= b;
    layer0_outputs(554) <= a or b;
    layer0_outputs(555) <= a xor b;
    layer0_outputs(556) <= a xor b;
    layer0_outputs(557) <= a or b;
    layer0_outputs(558) <= not (a xor b);
    layer0_outputs(559) <= a xor b;
    layer0_outputs(560) <= not (a xor b);
    layer0_outputs(561) <= not (a or b);
    layer0_outputs(562) <= a or b;
    layer0_outputs(563) <= a xor b;
    layer0_outputs(564) <= b and not a;
    layer0_outputs(565) <= b and not a;
    layer0_outputs(566) <= not b or a;
    layer0_outputs(567) <= not a or b;
    layer0_outputs(568) <= not a or b;
    layer0_outputs(569) <= a xor b;
    layer0_outputs(570) <= a xor b;
    layer0_outputs(571) <= a or b;
    layer0_outputs(572) <= b and not a;
    layer0_outputs(573) <= a or b;
    layer0_outputs(574) <= not a;
    layer0_outputs(575) <= not a;
    layer0_outputs(576) <= not (a xor b);
    layer0_outputs(577) <= b;
    layer0_outputs(578) <= 1'b1;
    layer0_outputs(579) <= a;
    layer0_outputs(580) <= not a;
    layer0_outputs(581) <= a or b;
    layer0_outputs(582) <= 1'b1;
    layer0_outputs(583) <= not a;
    layer0_outputs(584) <= not b;
    layer0_outputs(585) <= not (a xor b);
    layer0_outputs(586) <= 1'b1;
    layer0_outputs(587) <= a and b;
    layer0_outputs(588) <= a and not b;
    layer0_outputs(589) <= a;
    layer0_outputs(590) <= 1'b0;
    layer0_outputs(591) <= a;
    layer0_outputs(592) <= not (a xor b);
    layer0_outputs(593) <= 1'b1;
    layer0_outputs(594) <= a and not b;
    layer0_outputs(595) <= not b;
    layer0_outputs(596) <= a xor b;
    layer0_outputs(597) <= not a;
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= a;
    layer0_outputs(600) <= not a;
    layer0_outputs(601) <= a or b;
    layer0_outputs(602) <= a;
    layer0_outputs(603) <= 1'b0;
    layer0_outputs(604) <= b;
    layer0_outputs(605) <= b;
    layer0_outputs(606) <= a and b;
    layer0_outputs(607) <= a xor b;
    layer0_outputs(608) <= a xor b;
    layer0_outputs(609) <= a;
    layer0_outputs(610) <= a and not b;
    layer0_outputs(611) <= a and b;
    layer0_outputs(612) <= a;
    layer0_outputs(613) <= not b;
    layer0_outputs(614) <= a and not b;
    layer0_outputs(615) <= b;
    layer0_outputs(616) <= a and b;
    layer0_outputs(617) <= not b or a;
    layer0_outputs(618) <= a and not b;
    layer0_outputs(619) <= not (a xor b);
    layer0_outputs(620) <= not (a or b);
    layer0_outputs(621) <= a;
    layer0_outputs(622) <= a and b;
    layer0_outputs(623) <= a or b;
    layer0_outputs(624) <= a or b;
    layer0_outputs(625) <= a;
    layer0_outputs(626) <= not (a xor b);
    layer0_outputs(627) <= a xor b;
    layer0_outputs(628) <= a xor b;
    layer0_outputs(629) <= a and not b;
    layer0_outputs(630) <= not a;
    layer0_outputs(631) <= a and not b;
    layer0_outputs(632) <= b;
    layer0_outputs(633) <= not (a xor b);
    layer0_outputs(634) <= not (a xor b);
    layer0_outputs(635) <= not (a or b);
    layer0_outputs(636) <= 1'b0;
    layer0_outputs(637) <= a or b;
    layer0_outputs(638) <= a xor b;
    layer0_outputs(639) <= a;
    layer0_outputs(640) <= not (a xor b);
    layer0_outputs(641) <= b and not a;
    layer0_outputs(642) <= not b or a;
    layer0_outputs(643) <= a;
    layer0_outputs(644) <= not b;
    layer0_outputs(645) <= a and b;
    layer0_outputs(646) <= b;
    layer0_outputs(647) <= 1'b1;
    layer0_outputs(648) <= a and b;
    layer0_outputs(649) <= a and b;
    layer0_outputs(650) <= a xor b;
    layer0_outputs(651) <= not b;
    layer0_outputs(652) <= not a or b;
    layer0_outputs(653) <= not b;
    layer0_outputs(654) <= b;
    layer0_outputs(655) <= a xor b;
    layer0_outputs(656) <= b;
    layer0_outputs(657) <= a or b;
    layer0_outputs(658) <= not b or a;
    layer0_outputs(659) <= b and not a;
    layer0_outputs(660) <= b;
    layer0_outputs(661) <= a;
    layer0_outputs(662) <= not (a or b);
    layer0_outputs(663) <= a xor b;
    layer0_outputs(664) <= not a or b;
    layer0_outputs(665) <= a or b;
    layer0_outputs(666) <= a and not b;
    layer0_outputs(667) <= a and not b;
    layer0_outputs(668) <= not a;
    layer0_outputs(669) <= a and not b;
    layer0_outputs(670) <= a;
    layer0_outputs(671) <= not a;
    layer0_outputs(672) <= a or b;
    layer0_outputs(673) <= not (a xor b);
    layer0_outputs(674) <= not (a or b);
    layer0_outputs(675) <= b;
    layer0_outputs(676) <= a;
    layer0_outputs(677) <= a or b;
    layer0_outputs(678) <= not b;
    layer0_outputs(679) <= not b;
    layer0_outputs(680) <= not (a or b);
    layer0_outputs(681) <= a or b;
    layer0_outputs(682) <= not b;
    layer0_outputs(683) <= not (a xor b);
    layer0_outputs(684) <= not b or a;
    layer0_outputs(685) <= not (a or b);
    layer0_outputs(686) <= not (a xor b);
    layer0_outputs(687) <= 1'b1;
    layer0_outputs(688) <= not (a or b);
    layer0_outputs(689) <= a and not b;
    layer0_outputs(690) <= not a;
    layer0_outputs(691) <= b and not a;
    layer0_outputs(692) <= b;
    layer0_outputs(693) <= 1'b0;
    layer0_outputs(694) <= b and not a;
    layer0_outputs(695) <= a and not b;
    layer0_outputs(696) <= not a or b;
    layer0_outputs(697) <= b;
    layer0_outputs(698) <= a xor b;
    layer0_outputs(699) <= a or b;
    layer0_outputs(700) <= not b or a;
    layer0_outputs(701) <= not (a or b);
    layer0_outputs(702) <= b and not a;
    layer0_outputs(703) <= b and not a;
    layer0_outputs(704) <= a;
    layer0_outputs(705) <= a xor b;
    layer0_outputs(706) <= not b;
    layer0_outputs(707) <= not (a or b);
    layer0_outputs(708) <= 1'b1;
    layer0_outputs(709) <= b;
    layer0_outputs(710) <= a and not b;
    layer0_outputs(711) <= not a;
    layer0_outputs(712) <= not b;
    layer0_outputs(713) <= not (a or b);
    layer0_outputs(714) <= not (a or b);
    layer0_outputs(715) <= not a;
    layer0_outputs(716) <= a and not b;
    layer0_outputs(717) <= not a or b;
    layer0_outputs(718) <= not (a or b);
    layer0_outputs(719) <= a and not b;
    layer0_outputs(720) <= b and not a;
    layer0_outputs(721) <= a xor b;
    layer0_outputs(722) <= not (a or b);
    layer0_outputs(723) <= a and not b;
    layer0_outputs(724) <= not (a xor b);
    layer0_outputs(725) <= b;
    layer0_outputs(726) <= a or b;
    layer0_outputs(727) <= a;
    layer0_outputs(728) <= a;
    layer0_outputs(729) <= not a;
    layer0_outputs(730) <= not (a xor b);
    layer0_outputs(731) <= b;
    layer0_outputs(732) <= a or b;
    layer0_outputs(733) <= not (a or b);
    layer0_outputs(734) <= a;
    layer0_outputs(735) <= not a or b;
    layer0_outputs(736) <= a;
    layer0_outputs(737) <= a xor b;
    layer0_outputs(738) <= a xor b;
    layer0_outputs(739) <= a and not b;
    layer0_outputs(740) <= not a;
    layer0_outputs(741) <= a;
    layer0_outputs(742) <= a and not b;
    layer0_outputs(743) <= not (a or b);
    layer0_outputs(744) <= not (a xor b);
    layer0_outputs(745) <= a xor b;
    layer0_outputs(746) <= a and b;
    layer0_outputs(747) <= a xor b;
    layer0_outputs(748) <= a and b;
    layer0_outputs(749) <= not b;
    layer0_outputs(750) <= a;
    layer0_outputs(751) <= not (a and b);
    layer0_outputs(752) <= 1'b1;
    layer0_outputs(753) <= b;
    layer0_outputs(754) <= b;
    layer0_outputs(755) <= not a;
    layer0_outputs(756) <= b;
    layer0_outputs(757) <= not (a and b);
    layer0_outputs(758) <= b and not a;
    layer0_outputs(759) <= not (a or b);
    layer0_outputs(760) <= not a or b;
    layer0_outputs(761) <= not (a xor b);
    layer0_outputs(762) <= a or b;
    layer0_outputs(763) <= not b;
    layer0_outputs(764) <= a and b;
    layer0_outputs(765) <= not a or b;
    layer0_outputs(766) <= not (a xor b);
    layer0_outputs(767) <= not a;
    layer0_outputs(768) <= not b or a;
    layer0_outputs(769) <= a and b;
    layer0_outputs(770) <= not (a and b);
    layer0_outputs(771) <= a or b;
    layer0_outputs(772) <= not a;
    layer0_outputs(773) <= b;
    layer0_outputs(774) <= b;
    layer0_outputs(775) <= not a or b;
    layer0_outputs(776) <= not b or a;
    layer0_outputs(777) <= not (a xor b);
    layer0_outputs(778) <= a and not b;
    layer0_outputs(779) <= not (a xor b);
    layer0_outputs(780) <= b;
    layer0_outputs(781) <= a;
    layer0_outputs(782) <= not b or a;
    layer0_outputs(783) <= b and not a;
    layer0_outputs(784) <= a xor b;
    layer0_outputs(785) <= not (a xor b);
    layer0_outputs(786) <= a or b;
    layer0_outputs(787) <= a xor b;
    layer0_outputs(788) <= a or b;
    layer0_outputs(789) <= not b;
    layer0_outputs(790) <= a;
    layer0_outputs(791) <= a xor b;
    layer0_outputs(792) <= not (a xor b);
    layer0_outputs(793) <= b;
    layer0_outputs(794) <= not (a or b);
    layer0_outputs(795) <= a and not b;
    layer0_outputs(796) <= a;
    layer0_outputs(797) <= not b or a;
    layer0_outputs(798) <= not a;
    layer0_outputs(799) <= not b;
    layer0_outputs(800) <= a;
    layer0_outputs(801) <= not (a or b);
    layer0_outputs(802) <= a or b;
    layer0_outputs(803) <= b and not a;
    layer0_outputs(804) <= not (a xor b);
    layer0_outputs(805) <= not b;
    layer0_outputs(806) <= a or b;
    layer0_outputs(807) <= not b;
    layer0_outputs(808) <= not (a or b);
    layer0_outputs(809) <= not a;
    layer0_outputs(810) <= not a or b;
    layer0_outputs(811) <= a or b;
    layer0_outputs(812) <= b and not a;
    layer0_outputs(813) <= not (a xor b);
    layer0_outputs(814) <= not (a or b);
    layer0_outputs(815) <= not b;
    layer0_outputs(816) <= not (a xor b);
    layer0_outputs(817) <= not a or b;
    layer0_outputs(818) <= a and b;
    layer0_outputs(819) <= not b;
    layer0_outputs(820) <= not a;
    layer0_outputs(821) <= not (a xor b);
    layer0_outputs(822) <= not a;
    layer0_outputs(823) <= a or b;
    layer0_outputs(824) <= a or b;
    layer0_outputs(825) <= not (a xor b);
    layer0_outputs(826) <= not a;
    layer0_outputs(827) <= b and not a;
    layer0_outputs(828) <= b and not a;
    layer0_outputs(829) <= not (a xor b);
    layer0_outputs(830) <= a and b;
    layer0_outputs(831) <= not (a or b);
    layer0_outputs(832) <= not b or a;
    layer0_outputs(833) <= not b or a;
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= not (a or b);
    layer0_outputs(836) <= not (a or b);
    layer0_outputs(837) <= a;
    layer0_outputs(838) <= a xor b;
    layer0_outputs(839) <= a;
    layer0_outputs(840) <= not (a xor b);
    layer0_outputs(841) <= a xor b;
    layer0_outputs(842) <= a or b;
    layer0_outputs(843) <= not b or a;
    layer0_outputs(844) <= b;
    layer0_outputs(845) <= 1'b0;
    layer0_outputs(846) <= not (a or b);
    layer0_outputs(847) <= a;
    layer0_outputs(848) <= not (a xor b);
    layer0_outputs(849) <= b;
    layer0_outputs(850) <= a or b;
    layer0_outputs(851) <= a;
    layer0_outputs(852) <= b;
    layer0_outputs(853) <= not (a or b);
    layer0_outputs(854) <= 1'b0;
    layer0_outputs(855) <= not a or b;
    layer0_outputs(856) <= not a or b;
    layer0_outputs(857) <= not a;
    layer0_outputs(858) <= a xor b;
    layer0_outputs(859) <= not a;
    layer0_outputs(860) <= not (a and b);
    layer0_outputs(861) <= a;
    layer0_outputs(862) <= not a;
    layer0_outputs(863) <= a or b;
    layer0_outputs(864) <= a and not b;
    layer0_outputs(865) <= not a;
    layer0_outputs(866) <= not a;
    layer0_outputs(867) <= b;
    layer0_outputs(868) <= a xor b;
    layer0_outputs(869) <= not b or a;
    layer0_outputs(870) <= not (a and b);
    layer0_outputs(871) <= a or b;
    layer0_outputs(872) <= not (a xor b);
    layer0_outputs(873) <= a and not b;
    layer0_outputs(874) <= a;
    layer0_outputs(875) <= not a;
    layer0_outputs(876) <= a xor b;
    layer0_outputs(877) <= a or b;
    layer0_outputs(878) <= not a;
    layer0_outputs(879) <= b;
    layer0_outputs(880) <= b and not a;
    layer0_outputs(881) <= not b or a;
    layer0_outputs(882) <= a or b;
    layer0_outputs(883) <= not a or b;
    layer0_outputs(884) <= not (a xor b);
    layer0_outputs(885) <= not (a or b);
    layer0_outputs(886) <= a or b;
    layer0_outputs(887) <= not (a or b);
    layer0_outputs(888) <= not b or a;
    layer0_outputs(889) <= not a;
    layer0_outputs(890) <= not (a and b);
    layer0_outputs(891) <= not a;
    layer0_outputs(892) <= not b;
    layer0_outputs(893) <= not a;
    layer0_outputs(894) <= b;
    layer0_outputs(895) <= not b or a;
    layer0_outputs(896) <= not b;
    layer0_outputs(897) <= a xor b;
    layer0_outputs(898) <= a or b;
    layer0_outputs(899) <= b and not a;
    layer0_outputs(900) <= not (a xor b);
    layer0_outputs(901) <= b;
    layer0_outputs(902) <= not b;
    layer0_outputs(903) <= a;
    layer0_outputs(904) <= 1'b0;
    layer0_outputs(905) <= a and not b;
    layer0_outputs(906) <= not (a or b);
    layer0_outputs(907) <= not (a or b);
    layer0_outputs(908) <= a or b;
    layer0_outputs(909) <= a xor b;
    layer0_outputs(910) <= b;
    layer0_outputs(911) <= not a;
    layer0_outputs(912) <= not a;
    layer0_outputs(913) <= a and b;
    layer0_outputs(914) <= not b or a;
    layer0_outputs(915) <= not a;
    layer0_outputs(916) <= a;
    layer0_outputs(917) <= a and not b;
    layer0_outputs(918) <= not b or a;
    layer0_outputs(919) <= not a;
    layer0_outputs(920) <= not (a or b);
    layer0_outputs(921) <= b;
    layer0_outputs(922) <= b;
    layer0_outputs(923) <= 1'b1;
    layer0_outputs(924) <= not (a xor b);
    layer0_outputs(925) <= not b or a;
    layer0_outputs(926) <= not a or b;
    layer0_outputs(927) <= a or b;
    layer0_outputs(928) <= not b or a;
    layer0_outputs(929) <= a and b;
    layer0_outputs(930) <= not (a or b);
    layer0_outputs(931) <= not b or a;
    layer0_outputs(932) <= not (a xor b);
    layer0_outputs(933) <= not (a or b);
    layer0_outputs(934) <= a;
    layer0_outputs(935) <= not a or b;
    layer0_outputs(936) <= a or b;
    layer0_outputs(937) <= not b or a;
    layer0_outputs(938) <= not a;
    layer0_outputs(939) <= a or b;
    layer0_outputs(940) <= not (a xor b);
    layer0_outputs(941) <= not (a xor b);
    layer0_outputs(942) <= not b;
    layer0_outputs(943) <= a or b;
    layer0_outputs(944) <= not b or a;
    layer0_outputs(945) <= not (a or b);
    layer0_outputs(946) <= a or b;
    layer0_outputs(947) <= b;
    layer0_outputs(948) <= not (a xor b);
    layer0_outputs(949) <= b and not a;
    layer0_outputs(950) <= not (a xor b);
    layer0_outputs(951) <= b;
    layer0_outputs(952) <= not (a or b);
    layer0_outputs(953) <= a or b;
    layer0_outputs(954) <= not b or a;
    layer0_outputs(955) <= not (a xor b);
    layer0_outputs(956) <= a and not b;
    layer0_outputs(957) <= a xor b;
    layer0_outputs(958) <= not (a or b);
    layer0_outputs(959) <= b;
    layer0_outputs(960) <= a or b;
    layer0_outputs(961) <= b;
    layer0_outputs(962) <= not (a xor b);
    layer0_outputs(963) <= not (a or b);
    layer0_outputs(964) <= a and not b;
    layer0_outputs(965) <= b;
    layer0_outputs(966) <= not (a and b);
    layer0_outputs(967) <= b;
    layer0_outputs(968) <= a;
    layer0_outputs(969) <= not a;
    layer0_outputs(970) <= a;
    layer0_outputs(971) <= 1'b1;
    layer0_outputs(972) <= a and not b;
    layer0_outputs(973) <= a or b;
    layer0_outputs(974) <= not (a and b);
    layer0_outputs(975) <= not b or a;
    layer0_outputs(976) <= a and not b;
    layer0_outputs(977) <= not (a xor b);
    layer0_outputs(978) <= a xor b;
    layer0_outputs(979) <= not a;
    layer0_outputs(980) <= a;
    layer0_outputs(981) <= b;
    layer0_outputs(982) <= a or b;
    layer0_outputs(983) <= a;
    layer0_outputs(984) <= not (a xor b);
    layer0_outputs(985) <= not b or a;
    layer0_outputs(986) <= not b or a;
    layer0_outputs(987) <= a and not b;
    layer0_outputs(988) <= not (a xor b);
    layer0_outputs(989) <= not a;
    layer0_outputs(990) <= a or b;
    layer0_outputs(991) <= not a;
    layer0_outputs(992) <= a or b;
    layer0_outputs(993) <= a xor b;
    layer0_outputs(994) <= not a;
    layer0_outputs(995) <= not (a xor b);
    layer0_outputs(996) <= a xor b;
    layer0_outputs(997) <= not (a xor b);
    layer0_outputs(998) <= not a;
    layer0_outputs(999) <= a or b;
    layer0_outputs(1000) <= not b;
    layer0_outputs(1001) <= not a or b;
    layer0_outputs(1002) <= b;
    layer0_outputs(1003) <= a and not b;
    layer0_outputs(1004) <= a xor b;
    layer0_outputs(1005) <= a or b;
    layer0_outputs(1006) <= not b or a;
    layer0_outputs(1007) <= a and b;
    layer0_outputs(1008) <= a xor b;
    layer0_outputs(1009) <= not b;
    layer0_outputs(1010) <= a or b;
    layer0_outputs(1011) <= a and not b;
    layer0_outputs(1012) <= a xor b;
    layer0_outputs(1013) <= not (a or b);
    layer0_outputs(1014) <= 1'b0;
    layer0_outputs(1015) <= a;
    layer0_outputs(1016) <= a or b;
    layer0_outputs(1017) <= a;
    layer0_outputs(1018) <= a;
    layer0_outputs(1019) <= 1'b0;
    layer0_outputs(1020) <= not (a and b);
    layer0_outputs(1021) <= not b or a;
    layer0_outputs(1022) <= b;
    layer0_outputs(1023) <= 1'b0;
    layer0_outputs(1024) <= a or b;
    layer0_outputs(1025) <= not b or a;
    layer0_outputs(1026) <= not (a xor b);
    layer0_outputs(1027) <= a or b;
    layer0_outputs(1028) <= not a or b;
    layer0_outputs(1029) <= not b;
    layer0_outputs(1030) <= a or b;
    layer0_outputs(1031) <= b;
    layer0_outputs(1032) <= not a or b;
    layer0_outputs(1033) <= not b;
    layer0_outputs(1034) <= a xor b;
    layer0_outputs(1035) <= b and not a;
    layer0_outputs(1036) <= a and not b;
    layer0_outputs(1037) <= not (a or b);
    layer0_outputs(1038) <= not (a xor b);
    layer0_outputs(1039) <= not (a xor b);
    layer0_outputs(1040) <= not b;
    layer0_outputs(1041) <= not (a xor b);
    layer0_outputs(1042) <= a xor b;
    layer0_outputs(1043) <= a and b;
    layer0_outputs(1044) <= not a or b;
    layer0_outputs(1045) <= not b or a;
    layer0_outputs(1046) <= not a;
    layer0_outputs(1047) <= b;
    layer0_outputs(1048) <= a;
    layer0_outputs(1049) <= not b;
    layer0_outputs(1050) <= a or b;
    layer0_outputs(1051) <= not (a and b);
    layer0_outputs(1052) <= not b or a;
    layer0_outputs(1053) <= not a or b;
    layer0_outputs(1054) <= not (a and b);
    layer0_outputs(1055) <= not (a xor b);
    layer0_outputs(1056) <= 1'b0;
    layer0_outputs(1057) <= not a;
    layer0_outputs(1058) <= not a or b;
    layer0_outputs(1059) <= not (a or b);
    layer0_outputs(1060) <= not a or b;
    layer0_outputs(1061) <= a;
    layer0_outputs(1062) <= a and not b;
    layer0_outputs(1063) <= a or b;
    layer0_outputs(1064) <= not (a and b);
    layer0_outputs(1065) <= a or b;
    layer0_outputs(1066) <= a xor b;
    layer0_outputs(1067) <= a and not b;
    layer0_outputs(1068) <= not a or b;
    layer0_outputs(1069) <= a and b;
    layer0_outputs(1070) <= a or b;
    layer0_outputs(1071) <= a or b;
    layer0_outputs(1072) <= not a or b;
    layer0_outputs(1073) <= not (a xor b);
    layer0_outputs(1074) <= b and not a;
    layer0_outputs(1075) <= a xor b;
    layer0_outputs(1076) <= not b;
    layer0_outputs(1077) <= b and not a;
    layer0_outputs(1078) <= not (a or b);
    layer0_outputs(1079) <= not (a or b);
    layer0_outputs(1080) <= not (a or b);
    layer0_outputs(1081) <= not (a or b);
    layer0_outputs(1082) <= not (a xor b);
    layer0_outputs(1083) <= not a;
    layer0_outputs(1084) <= not (a or b);
    layer0_outputs(1085) <= a or b;
    layer0_outputs(1086) <= a xor b;
    layer0_outputs(1087) <= a xor b;
    layer0_outputs(1088) <= not b or a;
    layer0_outputs(1089) <= not a;
    layer0_outputs(1090) <= a and b;
    layer0_outputs(1091) <= a;
    layer0_outputs(1092) <= a or b;
    layer0_outputs(1093) <= not a;
    layer0_outputs(1094) <= not (a or b);
    layer0_outputs(1095) <= not (a or b);
    layer0_outputs(1096) <= a xor b;
    layer0_outputs(1097) <= not a;
    layer0_outputs(1098) <= not (a xor b);
    layer0_outputs(1099) <= b;
    layer0_outputs(1100) <= a and not b;
    layer0_outputs(1101) <= a;
    layer0_outputs(1102) <= not a;
    layer0_outputs(1103) <= not (a or b);
    layer0_outputs(1104) <= b and not a;
    layer0_outputs(1105) <= not (a or b);
    layer0_outputs(1106) <= b;
    layer0_outputs(1107) <= 1'b1;
    layer0_outputs(1108) <= b and not a;
    layer0_outputs(1109) <= a and not b;
    layer0_outputs(1110) <= not (a xor b);
    layer0_outputs(1111) <= not b or a;
    layer0_outputs(1112) <= b and not a;
    layer0_outputs(1113) <= b;
    layer0_outputs(1114) <= not (a or b);
    layer0_outputs(1115) <= b;
    layer0_outputs(1116) <= b and not a;
    layer0_outputs(1117) <= 1'b0;
    layer0_outputs(1118) <= not b;
    layer0_outputs(1119) <= not b;
    layer0_outputs(1120) <= a xor b;
    layer0_outputs(1121) <= a or b;
    layer0_outputs(1122) <= not b;
    layer0_outputs(1123) <= a or b;
    layer0_outputs(1124) <= not a;
    layer0_outputs(1125) <= a or b;
    layer0_outputs(1126) <= not b;
    layer0_outputs(1127) <= a;
    layer0_outputs(1128) <= a or b;
    layer0_outputs(1129) <= not (a or b);
    layer0_outputs(1130) <= not (a xor b);
    layer0_outputs(1131) <= a xor b;
    layer0_outputs(1132) <= a or b;
    layer0_outputs(1133) <= not b or a;
    layer0_outputs(1134) <= not b or a;
    layer0_outputs(1135) <= not a;
    layer0_outputs(1136) <= not a or b;
    layer0_outputs(1137) <= a or b;
    layer0_outputs(1138) <= not b;
    layer0_outputs(1139) <= not (a or b);
    layer0_outputs(1140) <= b;
    layer0_outputs(1141) <= not (a xor b);
    layer0_outputs(1142) <= not (a or b);
    layer0_outputs(1143) <= a xor b;
    layer0_outputs(1144) <= not b;
    layer0_outputs(1145) <= not a or b;
    layer0_outputs(1146) <= not b;
    layer0_outputs(1147) <= a xor b;
    layer0_outputs(1148) <= a xor b;
    layer0_outputs(1149) <= a or b;
    layer0_outputs(1150) <= not (a or b);
    layer0_outputs(1151) <= not a;
    layer0_outputs(1152) <= b;
    layer0_outputs(1153) <= not (a or b);
    layer0_outputs(1154) <= not a;
    layer0_outputs(1155) <= a;
    layer0_outputs(1156) <= b;
    layer0_outputs(1157) <= not b or a;
    layer0_outputs(1158) <= a;
    layer0_outputs(1159) <= not a or b;
    layer0_outputs(1160) <= not b;
    layer0_outputs(1161) <= a;
    layer0_outputs(1162) <= not (a xor b);
    layer0_outputs(1163) <= not (a and b);
    layer0_outputs(1164) <= a or b;
    layer0_outputs(1165) <= not b;
    layer0_outputs(1166) <= a;
    layer0_outputs(1167) <= a and not b;
    layer0_outputs(1168) <= not (a xor b);
    layer0_outputs(1169) <= b;
    layer0_outputs(1170) <= b;
    layer0_outputs(1171) <= not (a or b);
    layer0_outputs(1172) <= not b or a;
    layer0_outputs(1173) <= a;
    layer0_outputs(1174) <= a xor b;
    layer0_outputs(1175) <= b;
    layer0_outputs(1176) <= a;
    layer0_outputs(1177) <= b;
    layer0_outputs(1178) <= a or b;
    layer0_outputs(1179) <= a;
    layer0_outputs(1180) <= b;
    layer0_outputs(1181) <= not (a or b);
    layer0_outputs(1182) <= 1'b1;
    layer0_outputs(1183) <= a or b;
    layer0_outputs(1184) <= b;
    layer0_outputs(1185) <= a xor b;
    layer0_outputs(1186) <= not b;
    layer0_outputs(1187) <= b and not a;
    layer0_outputs(1188) <= not (a xor b);
    layer0_outputs(1189) <= not (a or b);
    layer0_outputs(1190) <= not a or b;
    layer0_outputs(1191) <= a and not b;
    layer0_outputs(1192) <= not b or a;
    layer0_outputs(1193) <= not (a or b);
    layer0_outputs(1194) <= not (a xor b);
    layer0_outputs(1195) <= not a or b;
    layer0_outputs(1196) <= a xor b;
    layer0_outputs(1197) <= a or b;
    layer0_outputs(1198) <= not (a or b);
    layer0_outputs(1199) <= not (a xor b);
    layer0_outputs(1200) <= not a or b;
    layer0_outputs(1201) <= not a;
    layer0_outputs(1202) <= a and not b;
    layer0_outputs(1203) <= not b;
    layer0_outputs(1204) <= not a;
    layer0_outputs(1205) <= a xor b;
    layer0_outputs(1206) <= b;
    layer0_outputs(1207) <= a xor b;
    layer0_outputs(1208) <= b;
    layer0_outputs(1209) <= b;
    layer0_outputs(1210) <= b;
    layer0_outputs(1211) <= not (a or b);
    layer0_outputs(1212) <= b and not a;
    layer0_outputs(1213) <= not a or b;
    layer0_outputs(1214) <= not (a or b);
    layer0_outputs(1215) <= not b;
    layer0_outputs(1216) <= not a;
    layer0_outputs(1217) <= 1'b1;
    layer0_outputs(1218) <= not (a xor b);
    layer0_outputs(1219) <= b and not a;
    layer0_outputs(1220) <= 1'b1;
    layer0_outputs(1221) <= b and not a;
    layer0_outputs(1222) <= not a;
    layer0_outputs(1223) <= not (a and b);
    layer0_outputs(1224) <= not (a xor b);
    layer0_outputs(1225) <= a and not b;
    layer0_outputs(1226) <= not b;
    layer0_outputs(1227) <= not (a or b);
    layer0_outputs(1228) <= a or b;
    layer0_outputs(1229) <= b and not a;
    layer0_outputs(1230) <= not a;
    layer0_outputs(1231) <= a or b;
    layer0_outputs(1232) <= not (a xor b);
    layer0_outputs(1233) <= not a or b;
    layer0_outputs(1234) <= not b or a;
    layer0_outputs(1235) <= not (a or b);
    layer0_outputs(1236) <= not b or a;
    layer0_outputs(1237) <= a xor b;
    layer0_outputs(1238) <= not b or a;
    layer0_outputs(1239) <= not (a or b);
    layer0_outputs(1240) <= not b or a;
    layer0_outputs(1241) <= a xor b;
    layer0_outputs(1242) <= not a or b;
    layer0_outputs(1243) <= a or b;
    layer0_outputs(1244) <= not a;
    layer0_outputs(1245) <= not (a xor b);
    layer0_outputs(1246) <= not (a or b);
    layer0_outputs(1247) <= a and not b;
    layer0_outputs(1248) <= not a or b;
    layer0_outputs(1249) <= b;
    layer0_outputs(1250) <= not b;
    layer0_outputs(1251) <= not (a or b);
    layer0_outputs(1252) <= b;
    layer0_outputs(1253) <= not (a or b);
    layer0_outputs(1254) <= not (a xor b);
    layer0_outputs(1255) <= b;
    layer0_outputs(1256) <= not (a and b);
    layer0_outputs(1257) <= a;
    layer0_outputs(1258) <= a or b;
    layer0_outputs(1259) <= not b or a;
    layer0_outputs(1260) <= a;
    layer0_outputs(1261) <= not a or b;
    layer0_outputs(1262) <= not a;
    layer0_outputs(1263) <= b;
    layer0_outputs(1264) <= not (a or b);
    layer0_outputs(1265) <= b and not a;
    layer0_outputs(1266) <= not a or b;
    layer0_outputs(1267) <= a and b;
    layer0_outputs(1268) <= not (a xor b);
    layer0_outputs(1269) <= not (a or b);
    layer0_outputs(1270) <= a and b;
    layer0_outputs(1271) <= b;
    layer0_outputs(1272) <= not a or b;
    layer0_outputs(1273) <= not (a xor b);
    layer0_outputs(1274) <= 1'b1;
    layer0_outputs(1275) <= not (a and b);
    layer0_outputs(1276) <= a or b;
    layer0_outputs(1277) <= not (a xor b);
    layer0_outputs(1278) <= not a;
    layer0_outputs(1279) <= a;
    layer0_outputs(1280) <= not b;
    layer0_outputs(1281) <= not (a or b);
    layer0_outputs(1282) <= not a;
    layer0_outputs(1283) <= a and not b;
    layer0_outputs(1284) <= a and not b;
    layer0_outputs(1285) <= a and not b;
    layer0_outputs(1286) <= a or b;
    layer0_outputs(1287) <= not b;
    layer0_outputs(1288) <= a;
    layer0_outputs(1289) <= not (a xor b);
    layer0_outputs(1290) <= not a or b;
    layer0_outputs(1291) <= a xor b;
    layer0_outputs(1292) <= 1'b0;
    layer0_outputs(1293) <= b;
    layer0_outputs(1294) <= a and not b;
    layer0_outputs(1295) <= not b;
    layer0_outputs(1296) <= a or b;
    layer0_outputs(1297) <= a or b;
    layer0_outputs(1298) <= not a or b;
    layer0_outputs(1299) <= not b;
    layer0_outputs(1300) <= not (a xor b);
    layer0_outputs(1301) <= not (a xor b);
    layer0_outputs(1302) <= not (a xor b);
    layer0_outputs(1303) <= not a or b;
    layer0_outputs(1304) <= a or b;
    layer0_outputs(1305) <= a;
    layer0_outputs(1306) <= not a or b;
    layer0_outputs(1307) <= not a or b;
    layer0_outputs(1308) <= not a;
    layer0_outputs(1309) <= b and not a;
    layer0_outputs(1310) <= not (a or b);
    layer0_outputs(1311) <= b;
    layer0_outputs(1312) <= b and not a;
    layer0_outputs(1313) <= not (a or b);
    layer0_outputs(1314) <= a xor b;
    layer0_outputs(1315) <= a and b;
    layer0_outputs(1316) <= not (a xor b);
    layer0_outputs(1317) <= a or b;
    layer0_outputs(1318) <= not a;
    layer0_outputs(1319) <= a or b;
    layer0_outputs(1320) <= not b;
    layer0_outputs(1321) <= a xor b;
    layer0_outputs(1322) <= b and not a;
    layer0_outputs(1323) <= a xor b;
    layer0_outputs(1324) <= a or b;
    layer0_outputs(1325) <= not (a xor b);
    layer0_outputs(1326) <= a xor b;
    layer0_outputs(1327) <= 1'b0;
    layer0_outputs(1328) <= a and not b;
    layer0_outputs(1329) <= not a;
    layer0_outputs(1330) <= b and not a;
    layer0_outputs(1331) <= a xor b;
    layer0_outputs(1332) <= b;
    layer0_outputs(1333) <= b and not a;
    layer0_outputs(1334) <= not (a or b);
    layer0_outputs(1335) <= a xor b;
    layer0_outputs(1336) <= a or b;
    layer0_outputs(1337) <= a;
    layer0_outputs(1338) <= 1'b1;
    layer0_outputs(1339) <= b and not a;
    layer0_outputs(1340) <= not a;
    layer0_outputs(1341) <= b;
    layer0_outputs(1342) <= not b or a;
    layer0_outputs(1343) <= b;
    layer0_outputs(1344) <= a or b;
    layer0_outputs(1345) <= not (a or b);
    layer0_outputs(1346) <= not (a xor b);
    layer0_outputs(1347) <= a or b;
    layer0_outputs(1348) <= a xor b;
    layer0_outputs(1349) <= a or b;
    layer0_outputs(1350) <= a or b;
    layer0_outputs(1351) <= not a;
    layer0_outputs(1352) <= not a;
    layer0_outputs(1353) <= a and b;
    layer0_outputs(1354) <= b and not a;
    layer0_outputs(1355) <= a or b;
    layer0_outputs(1356) <= not b;
    layer0_outputs(1357) <= not (a xor b);
    layer0_outputs(1358) <= b;
    layer0_outputs(1359) <= a and b;
    layer0_outputs(1360) <= a xor b;
    layer0_outputs(1361) <= a or b;
    layer0_outputs(1362) <= 1'b1;
    layer0_outputs(1363) <= not a or b;
    layer0_outputs(1364) <= not a;
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= not b;
    layer0_outputs(1367) <= a or b;
    layer0_outputs(1368) <= not (a and b);
    layer0_outputs(1369) <= not a or b;
    layer0_outputs(1370) <= not (a xor b);
    layer0_outputs(1371) <= b;
    layer0_outputs(1372) <= not (a xor b);
    layer0_outputs(1373) <= not (a or b);
    layer0_outputs(1374) <= b;
    layer0_outputs(1375) <= a;
    layer0_outputs(1376) <= a xor b;
    layer0_outputs(1377) <= not (a xor b);
    layer0_outputs(1378) <= a;
    layer0_outputs(1379) <= not (a xor b);
    layer0_outputs(1380) <= a or b;
    layer0_outputs(1381) <= a or b;
    layer0_outputs(1382) <= not b or a;
    layer0_outputs(1383) <= not a;
    layer0_outputs(1384) <= a;
    layer0_outputs(1385) <= a and not b;
    layer0_outputs(1386) <= not b or a;
    layer0_outputs(1387) <= not (a xor b);
    layer0_outputs(1388) <= b and not a;
    layer0_outputs(1389) <= not b or a;
    layer0_outputs(1390) <= not (a and b);
    layer0_outputs(1391) <= a or b;
    layer0_outputs(1392) <= a and not b;
    layer0_outputs(1393) <= not b;
    layer0_outputs(1394) <= not b;
    layer0_outputs(1395) <= not b;
    layer0_outputs(1396) <= not b or a;
    layer0_outputs(1397) <= not (a and b);
    layer0_outputs(1398) <= not a or b;
    layer0_outputs(1399) <= a xor b;
    layer0_outputs(1400) <= not (a or b);
    layer0_outputs(1401) <= b;
    layer0_outputs(1402) <= a;
    layer0_outputs(1403) <= a and not b;
    layer0_outputs(1404) <= a;
    layer0_outputs(1405) <= not b or a;
    layer0_outputs(1406) <= a and not b;
    layer0_outputs(1407) <= not b;
    layer0_outputs(1408) <= not a;
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= a and b;
    layer0_outputs(1411) <= not a;
    layer0_outputs(1412) <= not a;
    layer0_outputs(1413) <= not (a xor b);
    layer0_outputs(1414) <= a or b;
    layer0_outputs(1415) <= 1'b0;
    layer0_outputs(1416) <= a and not b;
    layer0_outputs(1417) <= not b;
    layer0_outputs(1418) <= not a;
    layer0_outputs(1419) <= not a;
    layer0_outputs(1420) <= not a;
    layer0_outputs(1421) <= a or b;
    layer0_outputs(1422) <= a or b;
    layer0_outputs(1423) <= not b;
    layer0_outputs(1424) <= 1'b1;
    layer0_outputs(1425) <= not (a and b);
    layer0_outputs(1426) <= not (a or b);
    layer0_outputs(1427) <= a xor b;
    layer0_outputs(1428) <= not (a or b);
    layer0_outputs(1429) <= 1'b0;
    layer0_outputs(1430) <= a and not b;
    layer0_outputs(1431) <= b;
    layer0_outputs(1432) <= not a or b;
    layer0_outputs(1433) <= a;
    layer0_outputs(1434) <= b;
    layer0_outputs(1435) <= b;
    layer0_outputs(1436) <= not a;
    layer0_outputs(1437) <= not (a xor b);
    layer0_outputs(1438) <= a and not b;
    layer0_outputs(1439) <= not a or b;
    layer0_outputs(1440) <= not b;
    layer0_outputs(1441) <= b;
    layer0_outputs(1442) <= 1'b1;
    layer0_outputs(1443) <= not a or b;
    layer0_outputs(1444) <= 1'b0;
    layer0_outputs(1445) <= not b or a;
    layer0_outputs(1446) <= not a or b;
    layer0_outputs(1447) <= a or b;
    layer0_outputs(1448) <= b;
    layer0_outputs(1449) <= not a;
    layer0_outputs(1450) <= a or b;
    layer0_outputs(1451) <= not b;
    layer0_outputs(1452) <= a xor b;
    layer0_outputs(1453) <= a or b;
    layer0_outputs(1454) <= not (a or b);
    layer0_outputs(1455) <= not (a or b);
    layer0_outputs(1456) <= a and not b;
    layer0_outputs(1457) <= b and not a;
    layer0_outputs(1458) <= a or b;
    layer0_outputs(1459) <= a or b;
    layer0_outputs(1460) <= a xor b;
    layer0_outputs(1461) <= not (a or b);
    layer0_outputs(1462) <= b and not a;
    layer0_outputs(1463) <= a xor b;
    layer0_outputs(1464) <= not a;
    layer0_outputs(1465) <= a;
    layer0_outputs(1466) <= not (a xor b);
    layer0_outputs(1467) <= not a or b;
    layer0_outputs(1468) <= not (a xor b);
    layer0_outputs(1469) <= not a or b;
    layer0_outputs(1470) <= a and b;
    layer0_outputs(1471) <= not b or a;
    layer0_outputs(1472) <= not (a or b);
    layer0_outputs(1473) <= not (a xor b);
    layer0_outputs(1474) <= not b;
    layer0_outputs(1475) <= a xor b;
    layer0_outputs(1476) <= not b or a;
    layer0_outputs(1477) <= 1'b1;
    layer0_outputs(1478) <= a and not b;
    layer0_outputs(1479) <= b;
    layer0_outputs(1480) <= not a or b;
    layer0_outputs(1481) <= not (a xor b);
    layer0_outputs(1482) <= a or b;
    layer0_outputs(1483) <= 1'b1;
    layer0_outputs(1484) <= not a;
    layer0_outputs(1485) <= 1'b1;
    layer0_outputs(1486) <= a and not b;
    layer0_outputs(1487) <= not b;
    layer0_outputs(1488) <= b and not a;
    layer0_outputs(1489) <= a and b;
    layer0_outputs(1490) <= not a or b;
    layer0_outputs(1491) <= a or b;
    layer0_outputs(1492) <= not (a or b);
    layer0_outputs(1493) <= a xor b;
    layer0_outputs(1494) <= a or b;
    layer0_outputs(1495) <= not b or a;
    layer0_outputs(1496) <= b;
    layer0_outputs(1497) <= a;
    layer0_outputs(1498) <= a xor b;
    layer0_outputs(1499) <= a;
    layer0_outputs(1500) <= a xor b;
    layer0_outputs(1501) <= not (a xor b);
    layer0_outputs(1502) <= not b;
    layer0_outputs(1503) <= b;
    layer0_outputs(1504) <= not b;
    layer0_outputs(1505) <= not (a or b);
    layer0_outputs(1506) <= not a or b;
    layer0_outputs(1507) <= b;
    layer0_outputs(1508) <= a and not b;
    layer0_outputs(1509) <= not b or a;
    layer0_outputs(1510) <= not b;
    layer0_outputs(1511) <= not a;
    layer0_outputs(1512) <= not (a xor b);
    layer0_outputs(1513) <= a and not b;
    layer0_outputs(1514) <= not (a xor b);
    layer0_outputs(1515) <= 1'b0;
    layer0_outputs(1516) <= a xor b;
    layer0_outputs(1517) <= b;
    layer0_outputs(1518) <= a and not b;
    layer0_outputs(1519) <= not (a or b);
    layer0_outputs(1520) <= a xor b;
    layer0_outputs(1521) <= not (a and b);
    layer0_outputs(1522) <= not (a or b);
    layer0_outputs(1523) <= not b;
    layer0_outputs(1524) <= a or b;
    layer0_outputs(1525) <= a;
    layer0_outputs(1526) <= not a or b;
    layer0_outputs(1527) <= not (a xor b);
    layer0_outputs(1528) <= not b or a;
    layer0_outputs(1529) <= 1'b0;
    layer0_outputs(1530) <= b and not a;
    layer0_outputs(1531) <= not b;
    layer0_outputs(1532) <= not a;
    layer0_outputs(1533) <= a or b;
    layer0_outputs(1534) <= not (a or b);
    layer0_outputs(1535) <= not b or a;
    layer0_outputs(1536) <= not (a xor b);
    layer0_outputs(1537) <= a or b;
    layer0_outputs(1538) <= not b or a;
    layer0_outputs(1539) <= a and not b;
    layer0_outputs(1540) <= not b;
    layer0_outputs(1541) <= not (a xor b);
    layer0_outputs(1542) <= b and not a;
    layer0_outputs(1543) <= 1'b1;
    layer0_outputs(1544) <= not a;
    layer0_outputs(1545) <= not (a and b);
    layer0_outputs(1546) <= a xor b;
    layer0_outputs(1547) <= a and b;
    layer0_outputs(1548) <= not a;
    layer0_outputs(1549) <= a and not b;
    layer0_outputs(1550) <= not b or a;
    layer0_outputs(1551) <= 1'b0;
    layer0_outputs(1552) <= not (a or b);
    layer0_outputs(1553) <= not a;
    layer0_outputs(1554) <= not (a xor b);
    layer0_outputs(1555) <= b and not a;
    layer0_outputs(1556) <= b;
    layer0_outputs(1557) <= b;
    layer0_outputs(1558) <= a xor b;
    layer0_outputs(1559) <= 1'b1;
    layer0_outputs(1560) <= not a;
    layer0_outputs(1561) <= b;
    layer0_outputs(1562) <= not b or a;
    layer0_outputs(1563) <= a xor b;
    layer0_outputs(1564) <= not b or a;
    layer0_outputs(1565) <= not a or b;
    layer0_outputs(1566) <= b;
    layer0_outputs(1567) <= a and not b;
    layer0_outputs(1568) <= not b;
    layer0_outputs(1569) <= not b or a;
    layer0_outputs(1570) <= not b;
    layer0_outputs(1571) <= not (a or b);
    layer0_outputs(1572) <= not b;
    layer0_outputs(1573) <= not b;
    layer0_outputs(1574) <= not a or b;
    layer0_outputs(1575) <= b;
    layer0_outputs(1576) <= not b;
    layer0_outputs(1577) <= not (a xor b);
    layer0_outputs(1578) <= 1'b0;
    layer0_outputs(1579) <= a and not b;
    layer0_outputs(1580) <= not (a or b);
    layer0_outputs(1581) <= a xor b;
    layer0_outputs(1582) <= a xor b;
    layer0_outputs(1583) <= b;
    layer0_outputs(1584) <= not b;
    layer0_outputs(1585) <= 1'b1;
    layer0_outputs(1586) <= b and not a;
    layer0_outputs(1587) <= a and b;
    layer0_outputs(1588) <= 1'b0;
    layer0_outputs(1589) <= not (a xor b);
    layer0_outputs(1590) <= b;
    layer0_outputs(1591) <= b;
    layer0_outputs(1592) <= a xor b;
    layer0_outputs(1593) <= not a or b;
    layer0_outputs(1594) <= not b or a;
    layer0_outputs(1595) <= not a;
    layer0_outputs(1596) <= not b;
    layer0_outputs(1597) <= not b or a;
    layer0_outputs(1598) <= a or b;
    layer0_outputs(1599) <= a or b;
    layer0_outputs(1600) <= not a or b;
    layer0_outputs(1601) <= 1'b1;
    layer0_outputs(1602) <= a;
    layer0_outputs(1603) <= b;
    layer0_outputs(1604) <= not (a xor b);
    layer0_outputs(1605) <= not b or a;
    layer0_outputs(1606) <= a xor b;
    layer0_outputs(1607) <= not (a or b);
    layer0_outputs(1608) <= not b;
    layer0_outputs(1609) <= a and not b;
    layer0_outputs(1610) <= not (a or b);
    layer0_outputs(1611) <= b;
    layer0_outputs(1612) <= not (a and b);
    layer0_outputs(1613) <= a or b;
    layer0_outputs(1614) <= 1'b1;
    layer0_outputs(1615) <= not a;
    layer0_outputs(1616) <= not (a xor b);
    layer0_outputs(1617) <= b;
    layer0_outputs(1618) <= a or b;
    layer0_outputs(1619) <= b and not a;
    layer0_outputs(1620) <= a;
    layer0_outputs(1621) <= a or b;
    layer0_outputs(1622) <= b and not a;
    layer0_outputs(1623) <= not b or a;
    layer0_outputs(1624) <= a and not b;
    layer0_outputs(1625) <= not (a or b);
    layer0_outputs(1626) <= a;
    layer0_outputs(1627) <= a xor b;
    layer0_outputs(1628) <= not a;
    layer0_outputs(1629) <= a;
    layer0_outputs(1630) <= not b;
    layer0_outputs(1631) <= not (a or b);
    layer0_outputs(1632) <= not (a and b);
    layer0_outputs(1633) <= not (a or b);
    layer0_outputs(1634) <= a xor b;
    layer0_outputs(1635) <= not a or b;
    layer0_outputs(1636) <= not b or a;
    layer0_outputs(1637) <= not b;
    layer0_outputs(1638) <= not a;
    layer0_outputs(1639) <= a xor b;
    layer0_outputs(1640) <= a or b;
    layer0_outputs(1641) <= a and not b;
    layer0_outputs(1642) <= a or b;
    layer0_outputs(1643) <= a and not b;
    layer0_outputs(1644) <= not a or b;
    layer0_outputs(1645) <= not (a and b);
    layer0_outputs(1646) <= b;
    layer0_outputs(1647) <= a xor b;
    layer0_outputs(1648) <= a xor b;
    layer0_outputs(1649) <= a xor b;
    layer0_outputs(1650) <= b;
    layer0_outputs(1651) <= b;
    layer0_outputs(1652) <= 1'b0;
    layer0_outputs(1653) <= a and not b;
    layer0_outputs(1654) <= a or b;
    layer0_outputs(1655) <= a xor b;
    layer0_outputs(1656) <= not (a xor b);
    layer0_outputs(1657) <= not (a xor b);
    layer0_outputs(1658) <= b and not a;
    layer0_outputs(1659) <= not a or b;
    layer0_outputs(1660) <= a;
    layer0_outputs(1661) <= a and b;
    layer0_outputs(1662) <= not a or b;
    layer0_outputs(1663) <= a xor b;
    layer0_outputs(1664) <= not a;
    layer0_outputs(1665) <= not (a or b);
    layer0_outputs(1666) <= not b or a;
    layer0_outputs(1667) <= b;
    layer0_outputs(1668) <= b;
    layer0_outputs(1669) <= not b or a;
    layer0_outputs(1670) <= a and b;
    layer0_outputs(1671) <= not b or a;
    layer0_outputs(1672) <= not b or a;
    layer0_outputs(1673) <= b;
    layer0_outputs(1674) <= not b;
    layer0_outputs(1675) <= not (a xor b);
    layer0_outputs(1676) <= not (a or b);
    layer0_outputs(1677) <= not (a or b);
    layer0_outputs(1678) <= a;
    layer0_outputs(1679) <= not b or a;
    layer0_outputs(1680) <= 1'b0;
    layer0_outputs(1681) <= a or b;
    layer0_outputs(1682) <= not a or b;
    layer0_outputs(1683) <= a and not b;
    layer0_outputs(1684) <= not b;
    layer0_outputs(1685) <= not b or a;
    layer0_outputs(1686) <= not b;
    layer0_outputs(1687) <= a xor b;
    layer0_outputs(1688) <= not b;
    layer0_outputs(1689) <= not (a xor b);
    layer0_outputs(1690) <= a;
    layer0_outputs(1691) <= a xor b;
    layer0_outputs(1692) <= a;
    layer0_outputs(1693) <= b;
    layer0_outputs(1694) <= not b or a;
    layer0_outputs(1695) <= a and b;
    layer0_outputs(1696) <= not (a or b);
    layer0_outputs(1697) <= not (a or b);
    layer0_outputs(1698) <= not a or b;
    layer0_outputs(1699) <= a;
    layer0_outputs(1700) <= a and not b;
    layer0_outputs(1701) <= not a or b;
    layer0_outputs(1702) <= b;
    layer0_outputs(1703) <= not (a and b);
    layer0_outputs(1704) <= not (a xor b);
    layer0_outputs(1705) <= a and not b;
    layer0_outputs(1706) <= b and not a;
    layer0_outputs(1707) <= a and not b;
    layer0_outputs(1708) <= a or b;
    layer0_outputs(1709) <= a and not b;
    layer0_outputs(1710) <= a and not b;
    layer0_outputs(1711) <= not a;
    layer0_outputs(1712) <= b and not a;
    layer0_outputs(1713) <= not b;
    layer0_outputs(1714) <= a;
    layer0_outputs(1715) <= a;
    layer0_outputs(1716) <= b;
    layer0_outputs(1717) <= b;
    layer0_outputs(1718) <= b;
    layer0_outputs(1719) <= not b;
    layer0_outputs(1720) <= a or b;
    layer0_outputs(1721) <= a;
    layer0_outputs(1722) <= a or b;
    layer0_outputs(1723) <= b;
    layer0_outputs(1724) <= not a or b;
    layer0_outputs(1725) <= a xor b;
    layer0_outputs(1726) <= a or b;
    layer0_outputs(1727) <= not a;
    layer0_outputs(1728) <= not (a or b);
    layer0_outputs(1729) <= a and not b;
    layer0_outputs(1730) <= a or b;
    layer0_outputs(1731) <= not (a or b);
    layer0_outputs(1732) <= not (a or b);
    layer0_outputs(1733) <= a or b;
    layer0_outputs(1734) <= b;
    layer0_outputs(1735) <= a xor b;
    layer0_outputs(1736) <= a and not b;
    layer0_outputs(1737) <= not b or a;
    layer0_outputs(1738) <= not a;
    layer0_outputs(1739) <= not (a xor b);
    layer0_outputs(1740) <= a;
    layer0_outputs(1741) <= not (a or b);
    layer0_outputs(1742) <= a or b;
    layer0_outputs(1743) <= a and not b;
    layer0_outputs(1744) <= not b or a;
    layer0_outputs(1745) <= not (a or b);
    layer0_outputs(1746) <= not b or a;
    layer0_outputs(1747) <= not (a or b);
    layer0_outputs(1748) <= b and not a;
    layer0_outputs(1749) <= a or b;
    layer0_outputs(1750) <= b and not a;
    layer0_outputs(1751) <= not (a or b);
    layer0_outputs(1752) <= not (a or b);
    layer0_outputs(1753) <= b;
    layer0_outputs(1754) <= not (a xor b);
    layer0_outputs(1755) <= not (a or b);
    layer0_outputs(1756) <= not b;
    layer0_outputs(1757) <= a xor b;
    layer0_outputs(1758) <= not b;
    layer0_outputs(1759) <= not a or b;
    layer0_outputs(1760) <= a and not b;
    layer0_outputs(1761) <= a xor b;
    layer0_outputs(1762) <= a xor b;
    layer0_outputs(1763) <= a;
    layer0_outputs(1764) <= a or b;
    layer0_outputs(1765) <= not b;
    layer0_outputs(1766) <= not (a or b);
    layer0_outputs(1767) <= not a;
    layer0_outputs(1768) <= a and not b;
    layer0_outputs(1769) <= not b or a;
    layer0_outputs(1770) <= a and not b;
    layer0_outputs(1771) <= not b or a;
    layer0_outputs(1772) <= a;
    layer0_outputs(1773) <= not a;
    layer0_outputs(1774) <= not (a xor b);
    layer0_outputs(1775) <= a or b;
    layer0_outputs(1776) <= not b;
    layer0_outputs(1777) <= not a;
    layer0_outputs(1778) <= a or b;
    layer0_outputs(1779) <= a and not b;
    layer0_outputs(1780) <= a;
    layer0_outputs(1781) <= a or b;
    layer0_outputs(1782) <= not (a and b);
    layer0_outputs(1783) <= not b;
    layer0_outputs(1784) <= not (a or b);
    layer0_outputs(1785) <= a and not b;
    layer0_outputs(1786) <= b;
    layer0_outputs(1787) <= not b;
    layer0_outputs(1788) <= a xor b;
    layer0_outputs(1789) <= a xor b;
    layer0_outputs(1790) <= a or b;
    layer0_outputs(1791) <= not (a and b);
    layer0_outputs(1792) <= 1'b0;
    layer0_outputs(1793) <= a or b;
    layer0_outputs(1794) <= a and b;
    layer0_outputs(1795) <= not (a xor b);
    layer0_outputs(1796) <= a xor b;
    layer0_outputs(1797) <= not (a or b);
    layer0_outputs(1798) <= a or b;
    layer0_outputs(1799) <= not a;
    layer0_outputs(1800) <= not (a or b);
    layer0_outputs(1801) <= a and not b;
    layer0_outputs(1802) <= a and not b;
    layer0_outputs(1803) <= not (a or b);
    layer0_outputs(1804) <= not (a or b);
    layer0_outputs(1805) <= not a;
    layer0_outputs(1806) <= not b;
    layer0_outputs(1807) <= not a or b;
    layer0_outputs(1808) <= a and not b;
    layer0_outputs(1809) <= a or b;
    layer0_outputs(1810) <= a or b;
    layer0_outputs(1811) <= 1'b0;
    layer0_outputs(1812) <= not a or b;
    layer0_outputs(1813) <= a and b;
    layer0_outputs(1814) <= b and not a;
    layer0_outputs(1815) <= a and not b;
    layer0_outputs(1816) <= b;
    layer0_outputs(1817) <= b;
    layer0_outputs(1818) <= a;
    layer0_outputs(1819) <= not a or b;
    layer0_outputs(1820) <= a;
    layer0_outputs(1821) <= a xor b;
    layer0_outputs(1822) <= a xor b;
    layer0_outputs(1823) <= not b;
    layer0_outputs(1824) <= not (a xor b);
    layer0_outputs(1825) <= 1'b1;
    layer0_outputs(1826) <= not (a xor b);
    layer0_outputs(1827) <= not (a or b);
    layer0_outputs(1828) <= b;
    layer0_outputs(1829) <= b and not a;
    layer0_outputs(1830) <= b and not a;
    layer0_outputs(1831) <= not b;
    layer0_outputs(1832) <= not a;
    layer0_outputs(1833) <= a and b;
    layer0_outputs(1834) <= not b or a;
    layer0_outputs(1835) <= a xor b;
    layer0_outputs(1836) <= not (a and b);
    layer0_outputs(1837) <= not a or b;
    layer0_outputs(1838) <= not b or a;
    layer0_outputs(1839) <= not a;
    layer0_outputs(1840) <= a or b;
    layer0_outputs(1841) <= not b;
    layer0_outputs(1842) <= 1'b1;
    layer0_outputs(1843) <= b and not a;
    layer0_outputs(1844) <= not a or b;
    layer0_outputs(1845) <= not (a or b);
    layer0_outputs(1846) <= not a or b;
    layer0_outputs(1847) <= a;
    layer0_outputs(1848) <= not a;
    layer0_outputs(1849) <= a or b;
    layer0_outputs(1850) <= not (a or b);
    layer0_outputs(1851) <= a;
    layer0_outputs(1852) <= a or b;
    layer0_outputs(1853) <= b;
    layer0_outputs(1854) <= b and not a;
    layer0_outputs(1855) <= b;
    layer0_outputs(1856) <= 1'b0;
    layer0_outputs(1857) <= b;
    layer0_outputs(1858) <= b;
    layer0_outputs(1859) <= not (a xor b);
    layer0_outputs(1860) <= not (a or b);
    layer0_outputs(1861) <= not (a or b);
    layer0_outputs(1862) <= not (a or b);
    layer0_outputs(1863) <= 1'b1;
    layer0_outputs(1864) <= b;
    layer0_outputs(1865) <= not b;
    layer0_outputs(1866) <= not b;
    layer0_outputs(1867) <= a and not b;
    layer0_outputs(1868) <= a;
    layer0_outputs(1869) <= a xor b;
    layer0_outputs(1870) <= b and not a;
    layer0_outputs(1871) <= not (a xor b);
    layer0_outputs(1872) <= a and not b;
    layer0_outputs(1873) <= not (a or b);
    layer0_outputs(1874) <= not b;
    layer0_outputs(1875) <= b and not a;
    layer0_outputs(1876) <= a or b;
    layer0_outputs(1877) <= not (a xor b);
    layer0_outputs(1878) <= a and not b;
    layer0_outputs(1879) <= not a or b;
    layer0_outputs(1880) <= not a or b;
    layer0_outputs(1881) <= not (a xor b);
    layer0_outputs(1882) <= 1'b1;
    layer0_outputs(1883) <= not b or a;
    layer0_outputs(1884) <= not (a and b);
    layer0_outputs(1885) <= not (a or b);
    layer0_outputs(1886) <= a xor b;
    layer0_outputs(1887) <= a;
    layer0_outputs(1888) <= a or b;
    layer0_outputs(1889) <= not a or b;
    layer0_outputs(1890) <= not (a or b);
    layer0_outputs(1891) <= not a or b;
    layer0_outputs(1892) <= a or b;
    layer0_outputs(1893) <= not a;
    layer0_outputs(1894) <= a and b;
    layer0_outputs(1895) <= not (a or b);
    layer0_outputs(1896) <= 1'b0;
    layer0_outputs(1897) <= not (a and b);
    layer0_outputs(1898) <= a and b;
    layer0_outputs(1899) <= not (a xor b);
    layer0_outputs(1900) <= not (a xor b);
    layer0_outputs(1901) <= a;
    layer0_outputs(1902) <= 1'b0;
    layer0_outputs(1903) <= 1'b0;
    layer0_outputs(1904) <= not (a or b);
    layer0_outputs(1905) <= a and not b;
    layer0_outputs(1906) <= not (a or b);
    layer0_outputs(1907) <= b;
    layer0_outputs(1908) <= not (a or b);
    layer0_outputs(1909) <= not b;
    layer0_outputs(1910) <= not b;
    layer0_outputs(1911) <= not b;
    layer0_outputs(1912) <= not a;
    layer0_outputs(1913) <= a xor b;
    layer0_outputs(1914) <= b and not a;
    layer0_outputs(1915) <= a or b;
    layer0_outputs(1916) <= b;
    layer0_outputs(1917) <= not b or a;
    layer0_outputs(1918) <= not b;
    layer0_outputs(1919) <= a and not b;
    layer0_outputs(1920) <= not b;
    layer0_outputs(1921) <= a or b;
    layer0_outputs(1922) <= not b or a;
    layer0_outputs(1923) <= 1'b0;
    layer0_outputs(1924) <= b;
    layer0_outputs(1925) <= not (a xor b);
    layer0_outputs(1926) <= not a or b;
    layer0_outputs(1927) <= not b or a;
    layer0_outputs(1928) <= a and b;
    layer0_outputs(1929) <= b;
    layer0_outputs(1930) <= b;
    layer0_outputs(1931) <= not b or a;
    layer0_outputs(1932) <= a and not b;
    layer0_outputs(1933) <= not b or a;
    layer0_outputs(1934) <= not (a xor b);
    layer0_outputs(1935) <= not (a xor b);
    layer0_outputs(1936) <= not a or b;
    layer0_outputs(1937) <= b;
    layer0_outputs(1938) <= not a or b;
    layer0_outputs(1939) <= not b or a;
    layer0_outputs(1940) <= 1'b1;
    layer0_outputs(1941) <= a;
    layer0_outputs(1942) <= a xor b;
    layer0_outputs(1943) <= b and not a;
    layer0_outputs(1944) <= a and b;
    layer0_outputs(1945) <= not b;
    layer0_outputs(1946) <= a or b;
    layer0_outputs(1947) <= 1'b0;
    layer0_outputs(1948) <= a xor b;
    layer0_outputs(1949) <= not (a or b);
    layer0_outputs(1950) <= not b;
    layer0_outputs(1951) <= not (a xor b);
    layer0_outputs(1952) <= a and not b;
    layer0_outputs(1953) <= b;
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= a xor b;
    layer0_outputs(1956) <= a;
    layer0_outputs(1957) <= not b or a;
    layer0_outputs(1958) <= not (a or b);
    layer0_outputs(1959) <= a or b;
    layer0_outputs(1960) <= a or b;
    layer0_outputs(1961) <= b and not a;
    layer0_outputs(1962) <= not a or b;
    layer0_outputs(1963) <= a xor b;
    layer0_outputs(1964) <= not b or a;
    layer0_outputs(1965) <= not b;
    layer0_outputs(1966) <= not a or b;
    layer0_outputs(1967) <= a and b;
    layer0_outputs(1968) <= 1'b0;
    layer0_outputs(1969) <= not b or a;
    layer0_outputs(1970) <= not a;
    layer0_outputs(1971) <= b;
    layer0_outputs(1972) <= b and not a;
    layer0_outputs(1973) <= a xor b;
    layer0_outputs(1974) <= not b;
    layer0_outputs(1975) <= a or b;
    layer0_outputs(1976) <= a or b;
    layer0_outputs(1977) <= a and b;
    layer0_outputs(1978) <= not (a or b);
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a or b;
    layer0_outputs(1981) <= not (a and b);
    layer0_outputs(1982) <= b and not a;
    layer0_outputs(1983) <= a xor b;
    layer0_outputs(1984) <= not (a xor b);
    layer0_outputs(1985) <= not b or a;
    layer0_outputs(1986) <= a or b;
    layer0_outputs(1987) <= not (a or b);
    layer0_outputs(1988) <= not a;
    layer0_outputs(1989) <= a and b;
    layer0_outputs(1990) <= a xor b;
    layer0_outputs(1991) <= not b;
    layer0_outputs(1992) <= 1'b1;
    layer0_outputs(1993) <= 1'b0;
    layer0_outputs(1994) <= not a or b;
    layer0_outputs(1995) <= not (a xor b);
    layer0_outputs(1996) <= a and not b;
    layer0_outputs(1997) <= not (a xor b);
    layer0_outputs(1998) <= a and not b;
    layer0_outputs(1999) <= a xor b;
    layer0_outputs(2000) <= a xor b;
    layer0_outputs(2001) <= a and not b;
    layer0_outputs(2002) <= not (a or b);
    layer0_outputs(2003) <= not a or b;
    layer0_outputs(2004) <= not (a or b);
    layer0_outputs(2005) <= a or b;
    layer0_outputs(2006) <= 1'b1;
    layer0_outputs(2007) <= b and not a;
    layer0_outputs(2008) <= a or b;
    layer0_outputs(2009) <= not a or b;
    layer0_outputs(2010) <= b and not a;
    layer0_outputs(2011) <= a;
    layer0_outputs(2012) <= a xor b;
    layer0_outputs(2013) <= 1'b0;
    layer0_outputs(2014) <= a xor b;
    layer0_outputs(2015) <= 1'b1;
    layer0_outputs(2016) <= not a or b;
    layer0_outputs(2017) <= not a;
    layer0_outputs(2018) <= a and not b;
    layer0_outputs(2019) <= not (a or b);
    layer0_outputs(2020) <= 1'b0;
    layer0_outputs(2021) <= a or b;
    layer0_outputs(2022) <= not a or b;
    layer0_outputs(2023) <= a and not b;
    layer0_outputs(2024) <= a and not b;
    layer0_outputs(2025) <= not (a xor b);
    layer0_outputs(2026) <= b and not a;
    layer0_outputs(2027) <= not b or a;
    layer0_outputs(2028) <= not (a xor b);
    layer0_outputs(2029) <= a or b;
    layer0_outputs(2030) <= a or b;
    layer0_outputs(2031) <= not b or a;
    layer0_outputs(2032) <= not (a or b);
    layer0_outputs(2033) <= 1'b0;
    layer0_outputs(2034) <= not a or b;
    layer0_outputs(2035) <= a;
    layer0_outputs(2036) <= 1'b1;
    layer0_outputs(2037) <= 1'b0;
    layer0_outputs(2038) <= not (a or b);
    layer0_outputs(2039) <= not (a and b);
    layer0_outputs(2040) <= not a;
    layer0_outputs(2041) <= a xor b;
    layer0_outputs(2042) <= not (a xor b);
    layer0_outputs(2043) <= a and b;
    layer0_outputs(2044) <= a or b;
    layer0_outputs(2045) <= a;
    layer0_outputs(2046) <= b and not a;
    layer0_outputs(2047) <= not (a or b);
    layer0_outputs(2048) <= not (a or b);
    layer0_outputs(2049) <= a and not b;
    layer0_outputs(2050) <= not a;
    layer0_outputs(2051) <= a or b;
    layer0_outputs(2052) <= b;
    layer0_outputs(2053) <= a xor b;
    layer0_outputs(2054) <= b;
    layer0_outputs(2055) <= a;
    layer0_outputs(2056) <= not b or a;
    layer0_outputs(2057) <= a or b;
    layer0_outputs(2058) <= b;
    layer0_outputs(2059) <= b;
    layer0_outputs(2060) <= a and not b;
    layer0_outputs(2061) <= 1'b1;
    layer0_outputs(2062) <= a or b;
    layer0_outputs(2063) <= a;
    layer0_outputs(2064) <= not b or a;
    layer0_outputs(2065) <= b;
    layer0_outputs(2066) <= a or b;
    layer0_outputs(2067) <= a or b;
    layer0_outputs(2068) <= not (a xor b);
    layer0_outputs(2069) <= not a or b;
    layer0_outputs(2070) <= not a or b;
    layer0_outputs(2071) <= 1'b1;
    layer0_outputs(2072) <= not (a xor b);
    layer0_outputs(2073) <= b;
    layer0_outputs(2074) <= a or b;
    layer0_outputs(2075) <= b and not a;
    layer0_outputs(2076) <= a or b;
    layer0_outputs(2077) <= a xor b;
    layer0_outputs(2078) <= not (a xor b);
    layer0_outputs(2079) <= a or b;
    layer0_outputs(2080) <= not b or a;
    layer0_outputs(2081) <= not (a xor b);
    layer0_outputs(2082) <= b and not a;
    layer0_outputs(2083) <= not b or a;
    layer0_outputs(2084) <= not (a xor b);
    layer0_outputs(2085) <= not b or a;
    layer0_outputs(2086) <= 1'b1;
    layer0_outputs(2087) <= 1'b1;
    layer0_outputs(2088) <= 1'b1;
    layer0_outputs(2089) <= a and not b;
    layer0_outputs(2090) <= a or b;
    layer0_outputs(2091) <= b;
    layer0_outputs(2092) <= a or b;
    layer0_outputs(2093) <= 1'b1;
    layer0_outputs(2094) <= a xor b;
    layer0_outputs(2095) <= not (a xor b);
    layer0_outputs(2096) <= b;
    layer0_outputs(2097) <= a or b;
    layer0_outputs(2098) <= not a or b;
    layer0_outputs(2099) <= not b or a;
    layer0_outputs(2100) <= a;
    layer0_outputs(2101) <= not b;
    layer0_outputs(2102) <= a xor b;
    layer0_outputs(2103) <= not (a or b);
    layer0_outputs(2104) <= not a;
    layer0_outputs(2105) <= not (a xor b);
    layer0_outputs(2106) <= not (a xor b);
    layer0_outputs(2107) <= a and b;
    layer0_outputs(2108) <= b;
    layer0_outputs(2109) <= not b;
    layer0_outputs(2110) <= a;
    layer0_outputs(2111) <= a xor b;
    layer0_outputs(2112) <= not (a or b);
    layer0_outputs(2113) <= a and not b;
    layer0_outputs(2114) <= not (a or b);
    layer0_outputs(2115) <= not a;
    layer0_outputs(2116) <= b and not a;
    layer0_outputs(2117) <= not a or b;
    layer0_outputs(2118) <= not b or a;
    layer0_outputs(2119) <= not (a or b);
    layer0_outputs(2120) <= not (a xor b);
    layer0_outputs(2121) <= b;
    layer0_outputs(2122) <= not a or b;
    layer0_outputs(2123) <= a;
    layer0_outputs(2124) <= a;
    layer0_outputs(2125) <= not b;
    layer0_outputs(2126) <= not b or a;
    layer0_outputs(2127) <= not a;
    layer0_outputs(2128) <= not (a xor b);
    layer0_outputs(2129) <= b;
    layer0_outputs(2130) <= a or b;
    layer0_outputs(2131) <= not (a or b);
    layer0_outputs(2132) <= a and b;
    layer0_outputs(2133) <= not b;
    layer0_outputs(2134) <= b;
    layer0_outputs(2135) <= a and not b;
    layer0_outputs(2136) <= not (a or b);
    layer0_outputs(2137) <= a or b;
    layer0_outputs(2138) <= not (a xor b);
    layer0_outputs(2139) <= a xor b;
    layer0_outputs(2140) <= a or b;
    layer0_outputs(2141) <= not a;
    layer0_outputs(2142) <= not (a or b);
    layer0_outputs(2143) <= a or b;
    layer0_outputs(2144) <= a or b;
    layer0_outputs(2145) <= a and not b;
    layer0_outputs(2146) <= a or b;
    layer0_outputs(2147) <= a and b;
    layer0_outputs(2148) <= b and not a;
    layer0_outputs(2149) <= not b or a;
    layer0_outputs(2150) <= a or b;
    layer0_outputs(2151) <= not (a or b);
    layer0_outputs(2152) <= a and not b;
    layer0_outputs(2153) <= not (a or b);
    layer0_outputs(2154) <= a xor b;
    layer0_outputs(2155) <= a;
    layer0_outputs(2156) <= not (a xor b);
    layer0_outputs(2157) <= not b or a;
    layer0_outputs(2158) <= b and not a;
    layer0_outputs(2159) <= not (a xor b);
    layer0_outputs(2160) <= a and not b;
    layer0_outputs(2161) <= not (a or b);
    layer0_outputs(2162) <= a or b;
    layer0_outputs(2163) <= a;
    layer0_outputs(2164) <= not b or a;
    layer0_outputs(2165) <= not b or a;
    layer0_outputs(2166) <= not b or a;
    layer0_outputs(2167) <= a and not b;
    layer0_outputs(2168) <= a or b;
    layer0_outputs(2169) <= not a or b;
    layer0_outputs(2170) <= not b;
    layer0_outputs(2171) <= a;
    layer0_outputs(2172) <= a or b;
    layer0_outputs(2173) <= not b;
    layer0_outputs(2174) <= a;
    layer0_outputs(2175) <= not (a or b);
    layer0_outputs(2176) <= b;
    layer0_outputs(2177) <= not (a or b);
    layer0_outputs(2178) <= a or b;
    layer0_outputs(2179) <= a xor b;
    layer0_outputs(2180) <= a and not b;
    layer0_outputs(2181) <= not a;
    layer0_outputs(2182) <= 1'b1;
    layer0_outputs(2183) <= not a or b;
    layer0_outputs(2184) <= not b;
    layer0_outputs(2185) <= b and not a;
    layer0_outputs(2186) <= a and b;
    layer0_outputs(2187) <= not a;
    layer0_outputs(2188) <= a or b;
    layer0_outputs(2189) <= b and not a;
    layer0_outputs(2190) <= not a;
    layer0_outputs(2191) <= not b or a;
    layer0_outputs(2192) <= b;
    layer0_outputs(2193) <= a and not b;
    layer0_outputs(2194) <= a or b;
    layer0_outputs(2195) <= a xor b;
    layer0_outputs(2196) <= b and not a;
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= not (a or b);
    layer0_outputs(2199) <= b;
    layer0_outputs(2200) <= a xor b;
    layer0_outputs(2201) <= a xor b;
    layer0_outputs(2202) <= not (a or b);
    layer0_outputs(2203) <= not b;
    layer0_outputs(2204) <= not b;
    layer0_outputs(2205) <= a or b;
    layer0_outputs(2206) <= a or b;
    layer0_outputs(2207) <= not a or b;
    layer0_outputs(2208) <= a xor b;
    layer0_outputs(2209) <= not b;
    layer0_outputs(2210) <= not b or a;
    layer0_outputs(2211) <= a xor b;
    layer0_outputs(2212) <= a and not b;
    layer0_outputs(2213) <= 1'b0;
    layer0_outputs(2214) <= not a or b;
    layer0_outputs(2215) <= a and b;
    layer0_outputs(2216) <= not a;
    layer0_outputs(2217) <= not (a or b);
    layer0_outputs(2218) <= not (a or b);
    layer0_outputs(2219) <= not a or b;
    layer0_outputs(2220) <= a or b;
    layer0_outputs(2221) <= not b;
    layer0_outputs(2222) <= a or b;
    layer0_outputs(2223) <= not b or a;
    layer0_outputs(2224) <= 1'b1;
    layer0_outputs(2225) <= not (a xor b);
    layer0_outputs(2226) <= not (a xor b);
    layer0_outputs(2227) <= b;
    layer0_outputs(2228) <= not b or a;
    layer0_outputs(2229) <= a;
    layer0_outputs(2230) <= a xor b;
    layer0_outputs(2231) <= not (a and b);
    layer0_outputs(2232) <= not (a or b);
    layer0_outputs(2233) <= b;
    layer0_outputs(2234) <= a xor b;
    layer0_outputs(2235) <= 1'b0;
    layer0_outputs(2236) <= a and not b;
    layer0_outputs(2237) <= not a or b;
    layer0_outputs(2238) <= not b;
    layer0_outputs(2239) <= b;
    layer0_outputs(2240) <= a and not b;
    layer0_outputs(2241) <= b and not a;
    layer0_outputs(2242) <= not b or a;
    layer0_outputs(2243) <= not a or b;
    layer0_outputs(2244) <= not a;
    layer0_outputs(2245) <= not a or b;
    layer0_outputs(2246) <= a and not b;
    layer0_outputs(2247) <= a and not b;
    layer0_outputs(2248) <= not (a xor b);
    layer0_outputs(2249) <= a or b;
    layer0_outputs(2250) <= b;
    layer0_outputs(2251) <= not b;
    layer0_outputs(2252) <= not b;
    layer0_outputs(2253) <= b and not a;
    layer0_outputs(2254) <= 1'b1;
    layer0_outputs(2255) <= b and not a;
    layer0_outputs(2256) <= a;
    layer0_outputs(2257) <= a and not b;
    layer0_outputs(2258) <= a;
    layer0_outputs(2259) <= a;
    layer0_outputs(2260) <= not a or b;
    layer0_outputs(2261) <= a;
    layer0_outputs(2262) <= b;
    layer0_outputs(2263) <= not b or a;
    layer0_outputs(2264) <= not (a xor b);
    layer0_outputs(2265) <= not a;
    layer0_outputs(2266) <= b;
    layer0_outputs(2267) <= 1'b1;
    layer0_outputs(2268) <= not (a or b);
    layer0_outputs(2269) <= not (a xor b);
    layer0_outputs(2270) <= not a;
    layer0_outputs(2271) <= not (a or b);
    layer0_outputs(2272) <= a xor b;
    layer0_outputs(2273) <= not a;
    layer0_outputs(2274) <= not (a xor b);
    layer0_outputs(2275) <= 1'b1;
    layer0_outputs(2276) <= a;
    layer0_outputs(2277) <= not (a xor b);
    layer0_outputs(2278) <= not b;
    layer0_outputs(2279) <= not (a or b);
    layer0_outputs(2280) <= not a or b;
    layer0_outputs(2281) <= a or b;
    layer0_outputs(2282) <= not (a xor b);
    layer0_outputs(2283) <= not (a xor b);
    layer0_outputs(2284) <= a xor b;
    layer0_outputs(2285) <= a;
    layer0_outputs(2286) <= not (a xor b);
    layer0_outputs(2287) <= not b or a;
    layer0_outputs(2288) <= a and not b;
    layer0_outputs(2289) <= not a;
    layer0_outputs(2290) <= b and not a;
    layer0_outputs(2291) <= 1'b0;
    layer0_outputs(2292) <= not (a xor b);
    layer0_outputs(2293) <= a;
    layer0_outputs(2294) <= not (a or b);
    layer0_outputs(2295) <= not b or a;
    layer0_outputs(2296) <= 1'b1;
    layer0_outputs(2297) <= b;
    layer0_outputs(2298) <= 1'b1;
    layer0_outputs(2299) <= a;
    layer0_outputs(2300) <= b and not a;
    layer0_outputs(2301) <= a and not b;
    layer0_outputs(2302) <= a and not b;
    layer0_outputs(2303) <= a xor b;
    layer0_outputs(2304) <= a xor b;
    layer0_outputs(2305) <= not a;
    layer0_outputs(2306) <= b;
    layer0_outputs(2307) <= a xor b;
    layer0_outputs(2308) <= not b or a;
    layer0_outputs(2309) <= 1'b0;
    layer0_outputs(2310) <= a or b;
    layer0_outputs(2311) <= b;
    layer0_outputs(2312) <= not a;
    layer0_outputs(2313) <= not (a or b);
    layer0_outputs(2314) <= a;
    layer0_outputs(2315) <= a xor b;
    layer0_outputs(2316) <= not (a or b);
    layer0_outputs(2317) <= not (a or b);
    layer0_outputs(2318) <= not a;
    layer0_outputs(2319) <= b;
    layer0_outputs(2320) <= b;
    layer0_outputs(2321) <= b;
    layer0_outputs(2322) <= a;
    layer0_outputs(2323) <= a and not b;
    layer0_outputs(2324) <= not b;
    layer0_outputs(2325) <= 1'b1;
    layer0_outputs(2326) <= not a;
    layer0_outputs(2327) <= not a or b;
    layer0_outputs(2328) <= a xor b;
    layer0_outputs(2329) <= a or b;
    layer0_outputs(2330) <= b and not a;
    layer0_outputs(2331) <= a and not b;
    layer0_outputs(2332) <= b;
    layer0_outputs(2333) <= not a;
    layer0_outputs(2334) <= a xor b;
    layer0_outputs(2335) <= not (a xor b);
    layer0_outputs(2336) <= a;
    layer0_outputs(2337) <= not (a or b);
    layer0_outputs(2338) <= a or b;
    layer0_outputs(2339) <= not b or a;
    layer0_outputs(2340) <= not a;
    layer0_outputs(2341) <= b and not a;
    layer0_outputs(2342) <= a xor b;
    layer0_outputs(2343) <= 1'b1;
    layer0_outputs(2344) <= not a or b;
    layer0_outputs(2345) <= a;
    layer0_outputs(2346) <= b;
    layer0_outputs(2347) <= a or b;
    layer0_outputs(2348) <= a or b;
    layer0_outputs(2349) <= 1'b0;
    layer0_outputs(2350) <= not (a or b);
    layer0_outputs(2351) <= b;
    layer0_outputs(2352) <= a and not b;
    layer0_outputs(2353) <= not b;
    layer0_outputs(2354) <= a xor b;
    layer0_outputs(2355) <= not (a and b);
    layer0_outputs(2356) <= not a or b;
    layer0_outputs(2357) <= not b;
    layer0_outputs(2358) <= b;
    layer0_outputs(2359) <= b and not a;
    layer0_outputs(2360) <= not b or a;
    layer0_outputs(2361) <= not (a and b);
    layer0_outputs(2362) <= not (a xor b);
    layer0_outputs(2363) <= not b;
    layer0_outputs(2364) <= not b or a;
    layer0_outputs(2365) <= b and not a;
    layer0_outputs(2366) <= a or b;
    layer0_outputs(2367) <= not a or b;
    layer0_outputs(2368) <= not a;
    layer0_outputs(2369) <= b and not a;
    layer0_outputs(2370) <= not (a xor b);
    layer0_outputs(2371) <= not b or a;
    layer0_outputs(2372) <= a or b;
    layer0_outputs(2373) <= not (a or b);
    layer0_outputs(2374) <= b;
    layer0_outputs(2375) <= a or b;
    layer0_outputs(2376) <= not b or a;
    layer0_outputs(2377) <= not b;
    layer0_outputs(2378) <= b and not a;
    layer0_outputs(2379) <= not b;
    layer0_outputs(2380) <= a or b;
    layer0_outputs(2381) <= a xor b;
    layer0_outputs(2382) <= b;
    layer0_outputs(2383) <= a xor b;
    layer0_outputs(2384) <= a and not b;
    layer0_outputs(2385) <= a xor b;
    layer0_outputs(2386) <= 1'b0;
    layer0_outputs(2387) <= not a or b;
    layer0_outputs(2388) <= a or b;
    layer0_outputs(2389) <= not b or a;
    layer0_outputs(2390) <= 1'b1;
    layer0_outputs(2391) <= a xor b;
    layer0_outputs(2392) <= a;
    layer0_outputs(2393) <= not a;
    layer0_outputs(2394) <= a xor b;
    layer0_outputs(2395) <= a or b;
    layer0_outputs(2396) <= b;
    layer0_outputs(2397) <= a and b;
    layer0_outputs(2398) <= not b or a;
    layer0_outputs(2399) <= not (a and b);
    layer0_outputs(2400) <= a;
    layer0_outputs(2401) <= not b or a;
    layer0_outputs(2402) <= not (a xor b);
    layer0_outputs(2403) <= not (a or b);
    layer0_outputs(2404) <= not a;
    layer0_outputs(2405) <= a;
    layer0_outputs(2406) <= not (a xor b);
    layer0_outputs(2407) <= not a or b;
    layer0_outputs(2408) <= a and not b;
    layer0_outputs(2409) <= not (a and b);
    layer0_outputs(2410) <= not b;
    layer0_outputs(2411) <= a;
    layer0_outputs(2412) <= not (a and b);
    layer0_outputs(2413) <= not (a xor b);
    layer0_outputs(2414) <= not (a or b);
    layer0_outputs(2415) <= not a;
    layer0_outputs(2416) <= a xor b;
    layer0_outputs(2417) <= not b;
    layer0_outputs(2418) <= 1'b1;
    layer0_outputs(2419) <= not b;
    layer0_outputs(2420) <= 1'b0;
    layer0_outputs(2421) <= not (a and b);
    layer0_outputs(2422) <= a and not b;
    layer0_outputs(2423) <= not a;
    layer0_outputs(2424) <= b and not a;
    layer0_outputs(2425) <= a;
    layer0_outputs(2426) <= not b or a;
    layer0_outputs(2427) <= b and not a;
    layer0_outputs(2428) <= not (a xor b);
    layer0_outputs(2429) <= 1'b0;
    layer0_outputs(2430) <= a and not b;
    layer0_outputs(2431) <= a and b;
    layer0_outputs(2432) <= not a;
    layer0_outputs(2433) <= 1'b1;
    layer0_outputs(2434) <= not (a xor b);
    layer0_outputs(2435) <= not b or a;
    layer0_outputs(2436) <= a xor b;
    layer0_outputs(2437) <= not (a or b);
    layer0_outputs(2438) <= not b;
    layer0_outputs(2439) <= b and not a;
    layer0_outputs(2440) <= a or b;
    layer0_outputs(2441) <= not b or a;
    layer0_outputs(2442) <= a and b;
    layer0_outputs(2443) <= a;
    layer0_outputs(2444) <= b and not a;
    layer0_outputs(2445) <= not (a xor b);
    layer0_outputs(2446) <= not (a xor b);
    layer0_outputs(2447) <= not b or a;
    layer0_outputs(2448) <= a and not b;
    layer0_outputs(2449) <= b;
    layer0_outputs(2450) <= not b;
    layer0_outputs(2451) <= a and b;
    layer0_outputs(2452) <= not (a or b);
    layer0_outputs(2453) <= not (a xor b);
    layer0_outputs(2454) <= not a or b;
    layer0_outputs(2455) <= not (a xor b);
    layer0_outputs(2456) <= a xor b;
    layer0_outputs(2457) <= not (a xor b);
    layer0_outputs(2458) <= not (a or b);
    layer0_outputs(2459) <= a and not b;
    layer0_outputs(2460) <= not a or b;
    layer0_outputs(2461) <= not (a or b);
    layer0_outputs(2462) <= a;
    layer0_outputs(2463) <= a or b;
    layer0_outputs(2464) <= not b;
    layer0_outputs(2465) <= not (a or b);
    layer0_outputs(2466) <= not a or b;
    layer0_outputs(2467) <= not b;
    layer0_outputs(2468) <= a or b;
    layer0_outputs(2469) <= not a;
    layer0_outputs(2470) <= a;
    layer0_outputs(2471) <= not b;
    layer0_outputs(2472) <= a or b;
    layer0_outputs(2473) <= a and b;
    layer0_outputs(2474) <= not (a or b);
    layer0_outputs(2475) <= 1'b1;
    layer0_outputs(2476) <= not (a or b);
    layer0_outputs(2477) <= not (a xor b);
    layer0_outputs(2478) <= b and not a;
    layer0_outputs(2479) <= not b;
    layer0_outputs(2480) <= a;
    layer0_outputs(2481) <= a or b;
    layer0_outputs(2482) <= not (a xor b);
    layer0_outputs(2483) <= a;
    layer0_outputs(2484) <= not a or b;
    layer0_outputs(2485) <= not a or b;
    layer0_outputs(2486) <= a xor b;
    layer0_outputs(2487) <= not b or a;
    layer0_outputs(2488) <= a or b;
    layer0_outputs(2489) <= a and not b;
    layer0_outputs(2490) <= not a;
    layer0_outputs(2491) <= b;
    layer0_outputs(2492) <= a or b;
    layer0_outputs(2493) <= b;
    layer0_outputs(2494) <= not (a and b);
    layer0_outputs(2495) <= not a;
    layer0_outputs(2496) <= not b or a;
    layer0_outputs(2497) <= not a or b;
    layer0_outputs(2498) <= not a;
    layer0_outputs(2499) <= b;
    layer0_outputs(2500) <= b;
    layer0_outputs(2501) <= not a or b;
    layer0_outputs(2502) <= not b or a;
    layer0_outputs(2503) <= not a;
    layer0_outputs(2504) <= a;
    layer0_outputs(2505) <= not b or a;
    layer0_outputs(2506) <= not (a xor b);
    layer0_outputs(2507) <= a;
    layer0_outputs(2508) <= b;
    layer0_outputs(2509) <= not a or b;
    layer0_outputs(2510) <= a xor b;
    layer0_outputs(2511) <= a and b;
    layer0_outputs(2512) <= a or b;
    layer0_outputs(2513) <= not (a xor b);
    layer0_outputs(2514) <= a and not b;
    layer0_outputs(2515) <= not a or b;
    layer0_outputs(2516) <= a xor b;
    layer0_outputs(2517) <= not b;
    layer0_outputs(2518) <= not (a or b);
    layer0_outputs(2519) <= a or b;
    layer0_outputs(2520) <= a or b;
    layer0_outputs(2521) <= b and not a;
    layer0_outputs(2522) <= a or b;
    layer0_outputs(2523) <= a and b;
    layer0_outputs(2524) <= not b;
    layer0_outputs(2525) <= a or b;
    layer0_outputs(2526) <= not b or a;
    layer0_outputs(2527) <= a and not b;
    layer0_outputs(2528) <= not (a or b);
    layer0_outputs(2529) <= not (a xor b);
    layer0_outputs(2530) <= not a;
    layer0_outputs(2531) <= not a;
    layer0_outputs(2532) <= b and not a;
    layer0_outputs(2533) <= a xor b;
    layer0_outputs(2534) <= a or b;
    layer0_outputs(2535) <= not a or b;
    layer0_outputs(2536) <= b;
    layer0_outputs(2537) <= not (a and b);
    layer0_outputs(2538) <= not a;
    layer0_outputs(2539) <= b;
    layer0_outputs(2540) <= not b;
    layer0_outputs(2541) <= not b or a;
    layer0_outputs(2542) <= b and not a;
    layer0_outputs(2543) <= not (a and b);
    layer0_outputs(2544) <= not (a and b);
    layer0_outputs(2545) <= b and not a;
    layer0_outputs(2546) <= a or b;
    layer0_outputs(2547) <= not a or b;
    layer0_outputs(2548) <= b;
    layer0_outputs(2549) <= not (a or b);
    layer0_outputs(2550) <= b;
    layer0_outputs(2551) <= a;
    layer0_outputs(2552) <= not (a or b);
    layer0_outputs(2553) <= b;
    layer0_outputs(2554) <= not (a xor b);
    layer0_outputs(2555) <= 1'b0;
    layer0_outputs(2556) <= not b or a;
    layer0_outputs(2557) <= not (a and b);
    layer0_outputs(2558) <= not a;
    layer0_outputs(2559) <= not b;
    layer0_outputs(2560) <= not b or a;
    layer0_outputs(2561) <= not (a xor b);
    layer0_outputs(2562) <= not (a or b);
    layer0_outputs(2563) <= b;
    layer0_outputs(2564) <= not a;
    layer0_outputs(2565) <= not (a xor b);
    layer0_outputs(2566) <= not b;
    layer0_outputs(2567) <= a or b;
    layer0_outputs(2568) <= b;
    layer0_outputs(2569) <= a;
    layer0_outputs(2570) <= not a or b;
    layer0_outputs(2571) <= a;
    layer0_outputs(2572) <= not b;
    layer0_outputs(2573) <= a or b;
    layer0_outputs(2574) <= a or b;
    layer0_outputs(2575) <= not a;
    layer0_outputs(2576) <= not (a xor b);
    layer0_outputs(2577) <= not a;
    layer0_outputs(2578) <= a;
    layer0_outputs(2579) <= not (a or b);
    layer0_outputs(2580) <= not a;
    layer0_outputs(2581) <= not (a xor b);
    layer0_outputs(2582) <= not (a or b);
    layer0_outputs(2583) <= not b;
    layer0_outputs(2584) <= b and not a;
    layer0_outputs(2585) <= not a or b;
    layer0_outputs(2586) <= a;
    layer0_outputs(2587) <= not (a xor b);
    layer0_outputs(2588) <= a or b;
    layer0_outputs(2589) <= not (a xor b);
    layer0_outputs(2590) <= a or b;
    layer0_outputs(2591) <= a and not b;
    layer0_outputs(2592) <= b;
    layer0_outputs(2593) <= a and not b;
    layer0_outputs(2594) <= not a or b;
    layer0_outputs(2595) <= not (a or b);
    layer0_outputs(2596) <= b and not a;
    layer0_outputs(2597) <= a xor b;
    layer0_outputs(2598) <= not b or a;
    layer0_outputs(2599) <= not (a xor b);
    layer0_outputs(2600) <= a xor b;
    layer0_outputs(2601) <= a and not b;
    layer0_outputs(2602) <= not a;
    layer0_outputs(2603) <= not (a or b);
    layer0_outputs(2604) <= not (a xor b);
    layer0_outputs(2605) <= not (a xor b);
    layer0_outputs(2606) <= not (a xor b);
    layer0_outputs(2607) <= not b;
    layer0_outputs(2608) <= a and b;
    layer0_outputs(2609) <= a;
    layer0_outputs(2610) <= not b or a;
    layer0_outputs(2611) <= not b;
    layer0_outputs(2612) <= 1'b1;
    layer0_outputs(2613) <= not a;
    layer0_outputs(2614) <= a or b;
    layer0_outputs(2615) <= a and not b;
    layer0_outputs(2616) <= a and not b;
    layer0_outputs(2617) <= a or b;
    layer0_outputs(2618) <= not a;
    layer0_outputs(2619) <= a and b;
    layer0_outputs(2620) <= not b;
    layer0_outputs(2621) <= not b or a;
    layer0_outputs(2622) <= a or b;
    layer0_outputs(2623) <= not b;
    layer0_outputs(2624) <= not (a or b);
    layer0_outputs(2625) <= a or b;
    layer0_outputs(2626) <= not b;
    layer0_outputs(2627) <= not (a xor b);
    layer0_outputs(2628) <= a;
    layer0_outputs(2629) <= a;
    layer0_outputs(2630) <= not a or b;
    layer0_outputs(2631) <= not a or b;
    layer0_outputs(2632) <= a xor b;
    layer0_outputs(2633) <= a xor b;
    layer0_outputs(2634) <= a or b;
    layer0_outputs(2635) <= b and not a;
    layer0_outputs(2636) <= not (a xor b);
    layer0_outputs(2637) <= not b or a;
    layer0_outputs(2638) <= a xor b;
    layer0_outputs(2639) <= not (a and b);
    layer0_outputs(2640) <= not (a or b);
    layer0_outputs(2641) <= not b;
    layer0_outputs(2642) <= not b;
    layer0_outputs(2643) <= not (a or b);
    layer0_outputs(2644) <= a and b;
    layer0_outputs(2645) <= not (a or b);
    layer0_outputs(2646) <= a or b;
    layer0_outputs(2647) <= not (a and b);
    layer0_outputs(2648) <= a or b;
    layer0_outputs(2649) <= b;
    layer0_outputs(2650) <= not (a or b);
    layer0_outputs(2651) <= not b;
    layer0_outputs(2652) <= a;
    layer0_outputs(2653) <= not (a xor b);
    layer0_outputs(2654) <= not a or b;
    layer0_outputs(2655) <= a;
    layer0_outputs(2656) <= a;
    layer0_outputs(2657) <= not (a or b);
    layer0_outputs(2658) <= a xor b;
    layer0_outputs(2659) <= a;
    layer0_outputs(2660) <= 1'b1;
    layer0_outputs(2661) <= not a;
    layer0_outputs(2662) <= b and not a;
    layer0_outputs(2663) <= b;
    layer0_outputs(2664) <= a and b;
    layer0_outputs(2665) <= a;
    layer0_outputs(2666) <= not (a or b);
    layer0_outputs(2667) <= not b;
    layer0_outputs(2668) <= a or b;
    layer0_outputs(2669) <= a or b;
    layer0_outputs(2670) <= not b;
    layer0_outputs(2671) <= not a or b;
    layer0_outputs(2672) <= not a;
    layer0_outputs(2673) <= not b;
    layer0_outputs(2674) <= not (a or b);
    layer0_outputs(2675) <= a xor b;
    layer0_outputs(2676) <= not a or b;
    layer0_outputs(2677) <= not (a xor b);
    layer0_outputs(2678) <= not b;
    layer0_outputs(2679) <= a or b;
    layer0_outputs(2680) <= not (a xor b);
    layer0_outputs(2681) <= a or b;
    layer0_outputs(2682) <= a xor b;
    layer0_outputs(2683) <= b;
    layer0_outputs(2684) <= not (a and b);
    layer0_outputs(2685) <= not (a and b);
    layer0_outputs(2686) <= a or b;
    layer0_outputs(2687) <= not (a or b);
    layer0_outputs(2688) <= b;
    layer0_outputs(2689) <= not b;
    layer0_outputs(2690) <= not (a or b);
    layer0_outputs(2691) <= not a;
    layer0_outputs(2692) <= not a;
    layer0_outputs(2693) <= not a;
    layer0_outputs(2694) <= a and not b;
    layer0_outputs(2695) <= a xor b;
    layer0_outputs(2696) <= not (a and b);
    layer0_outputs(2697) <= not (a and b);
    layer0_outputs(2698) <= not a;
    layer0_outputs(2699) <= not a or b;
    layer0_outputs(2700) <= not (a or b);
    layer0_outputs(2701) <= a;
    layer0_outputs(2702) <= not (a xor b);
    layer0_outputs(2703) <= not (a xor b);
    layer0_outputs(2704) <= b and not a;
    layer0_outputs(2705) <= not a or b;
    layer0_outputs(2706) <= a xor b;
    layer0_outputs(2707) <= 1'b0;
    layer0_outputs(2708) <= not a;
    layer0_outputs(2709) <= a and b;
    layer0_outputs(2710) <= a and b;
    layer0_outputs(2711) <= not b;
    layer0_outputs(2712) <= b;
    layer0_outputs(2713) <= a;
    layer0_outputs(2714) <= a and not b;
    layer0_outputs(2715) <= not (a or b);
    layer0_outputs(2716) <= a or b;
    layer0_outputs(2717) <= 1'b1;
    layer0_outputs(2718) <= a xor b;
    layer0_outputs(2719) <= not b or a;
    layer0_outputs(2720) <= 1'b0;
    layer0_outputs(2721) <= not b;
    layer0_outputs(2722) <= a or b;
    layer0_outputs(2723) <= not (a or b);
    layer0_outputs(2724) <= not (a xor b);
    layer0_outputs(2725) <= a;
    layer0_outputs(2726) <= not b;
    layer0_outputs(2727) <= a xor b;
    layer0_outputs(2728) <= not (a or b);
    layer0_outputs(2729) <= b and not a;
    layer0_outputs(2730) <= a xor b;
    layer0_outputs(2731) <= b and not a;
    layer0_outputs(2732) <= b and not a;
    layer0_outputs(2733) <= a or b;
    layer0_outputs(2734) <= not (a or b);
    layer0_outputs(2735) <= a or b;
    layer0_outputs(2736) <= not (a or b);
    layer0_outputs(2737) <= a xor b;
    layer0_outputs(2738) <= a xor b;
    layer0_outputs(2739) <= not (a or b);
    layer0_outputs(2740) <= a xor b;
    layer0_outputs(2741) <= not (a or b);
    layer0_outputs(2742) <= not (a and b);
    layer0_outputs(2743) <= not (a or b);
    layer0_outputs(2744) <= not b or a;
    layer0_outputs(2745) <= not (a or b);
    layer0_outputs(2746) <= a xor b;
    layer0_outputs(2747) <= b;
    layer0_outputs(2748) <= not a;
    layer0_outputs(2749) <= not (a and b);
    layer0_outputs(2750) <= a or b;
    layer0_outputs(2751) <= b and not a;
    layer0_outputs(2752) <= a;
    layer0_outputs(2753) <= not a;
    layer0_outputs(2754) <= b and not a;
    layer0_outputs(2755) <= a xor b;
    layer0_outputs(2756) <= b;
    layer0_outputs(2757) <= a;
    layer0_outputs(2758) <= a;
    layer0_outputs(2759) <= a xor b;
    layer0_outputs(2760) <= a or b;
    layer0_outputs(2761) <= 1'b0;
    layer0_outputs(2762) <= a or b;
    layer0_outputs(2763) <= not (a xor b);
    layer0_outputs(2764) <= a or b;
    layer0_outputs(2765) <= a or b;
    layer0_outputs(2766) <= not (a or b);
    layer0_outputs(2767) <= not b;
    layer0_outputs(2768) <= not a;
    layer0_outputs(2769) <= not a;
    layer0_outputs(2770) <= not b or a;
    layer0_outputs(2771) <= a;
    layer0_outputs(2772) <= a;
    layer0_outputs(2773) <= not b or a;
    layer0_outputs(2774) <= a;
    layer0_outputs(2775) <= 1'b1;
    layer0_outputs(2776) <= not b or a;
    layer0_outputs(2777) <= a and b;
    layer0_outputs(2778) <= b;
    layer0_outputs(2779) <= a or b;
    layer0_outputs(2780) <= not (a xor b);
    layer0_outputs(2781) <= not (a and b);
    layer0_outputs(2782) <= 1'b1;
    layer0_outputs(2783) <= a and b;
    layer0_outputs(2784) <= not (a or b);
    layer0_outputs(2785) <= not a;
    layer0_outputs(2786) <= not b;
    layer0_outputs(2787) <= not a or b;
    layer0_outputs(2788) <= not (a or b);
    layer0_outputs(2789) <= a or b;
    layer0_outputs(2790) <= not a or b;
    layer0_outputs(2791) <= b;
    layer0_outputs(2792) <= a;
    layer0_outputs(2793) <= b and not a;
    layer0_outputs(2794) <= not a;
    layer0_outputs(2795) <= a;
    layer0_outputs(2796) <= not (a and b);
    layer0_outputs(2797) <= b;
    layer0_outputs(2798) <= not (a xor b);
    layer0_outputs(2799) <= not a;
    layer0_outputs(2800) <= a and not b;
    layer0_outputs(2801) <= b and not a;
    layer0_outputs(2802) <= not a or b;
    layer0_outputs(2803) <= not (a xor b);
    layer0_outputs(2804) <= not (a or b);
    layer0_outputs(2805) <= not a or b;
    layer0_outputs(2806) <= not b or a;
    layer0_outputs(2807) <= not a or b;
    layer0_outputs(2808) <= b and not a;
    layer0_outputs(2809) <= not (a or b);
    layer0_outputs(2810) <= not (a xor b);
    layer0_outputs(2811) <= not b or a;
    layer0_outputs(2812) <= b and not a;
    layer0_outputs(2813) <= not a;
    layer0_outputs(2814) <= not (a or b);
    layer0_outputs(2815) <= a and not b;
    layer0_outputs(2816) <= not (a xor b);
    layer0_outputs(2817) <= not (a xor b);
    layer0_outputs(2818) <= a xor b;
    layer0_outputs(2819) <= not b;
    layer0_outputs(2820) <= a;
    layer0_outputs(2821) <= not b or a;
    layer0_outputs(2822) <= not b;
    layer0_outputs(2823) <= not (a and b);
    layer0_outputs(2824) <= a or b;
    layer0_outputs(2825) <= b and not a;
    layer0_outputs(2826) <= not a;
    layer0_outputs(2827) <= not b or a;
    layer0_outputs(2828) <= b;
    layer0_outputs(2829) <= a and not b;
    layer0_outputs(2830) <= a;
    layer0_outputs(2831) <= a and not b;
    layer0_outputs(2832) <= not b;
    layer0_outputs(2833) <= b and not a;
    layer0_outputs(2834) <= b;
    layer0_outputs(2835) <= b;
    layer0_outputs(2836) <= a;
    layer0_outputs(2837) <= a or b;
    layer0_outputs(2838) <= not a or b;
    layer0_outputs(2839) <= not b;
    layer0_outputs(2840) <= not (a xor b);
    layer0_outputs(2841) <= not (a xor b);
    layer0_outputs(2842) <= 1'b0;
    layer0_outputs(2843) <= not a;
    layer0_outputs(2844) <= not (a xor b);
    layer0_outputs(2845) <= not (a or b);
    layer0_outputs(2846) <= not (a or b);
    layer0_outputs(2847) <= not (a and b);
    layer0_outputs(2848) <= not b;
    layer0_outputs(2849) <= not a;
    layer0_outputs(2850) <= 1'b0;
    layer0_outputs(2851) <= not b;
    layer0_outputs(2852) <= a;
    layer0_outputs(2853) <= not (a xor b);
    layer0_outputs(2854) <= 1'b0;
    layer0_outputs(2855) <= not (a and b);
    layer0_outputs(2856) <= a xor b;
    layer0_outputs(2857) <= a or b;
    layer0_outputs(2858) <= not (a or b);
    layer0_outputs(2859) <= b;
    layer0_outputs(2860) <= not b;
    layer0_outputs(2861) <= b;
    layer0_outputs(2862) <= a xor b;
    layer0_outputs(2863) <= a;
    layer0_outputs(2864) <= a xor b;
    layer0_outputs(2865) <= b and not a;
    layer0_outputs(2866) <= not b;
    layer0_outputs(2867) <= not a;
    layer0_outputs(2868) <= b and not a;
    layer0_outputs(2869) <= not b;
    layer0_outputs(2870) <= b;
    layer0_outputs(2871) <= a xor b;
    layer0_outputs(2872) <= not b or a;
    layer0_outputs(2873) <= not (a xor b);
    layer0_outputs(2874) <= a or b;
    layer0_outputs(2875) <= not (a xor b);
    layer0_outputs(2876) <= not b;
    layer0_outputs(2877) <= not b;
    layer0_outputs(2878) <= b and not a;
    layer0_outputs(2879) <= b and not a;
    layer0_outputs(2880) <= a xor b;
    layer0_outputs(2881) <= not b or a;
    layer0_outputs(2882) <= not a;
    layer0_outputs(2883) <= not (a or b);
    layer0_outputs(2884) <= not (a or b);
    layer0_outputs(2885) <= not (a xor b);
    layer0_outputs(2886) <= a and b;
    layer0_outputs(2887) <= not (a or b);
    layer0_outputs(2888) <= not (a or b);
    layer0_outputs(2889) <= not (a or b);
    layer0_outputs(2890) <= a or b;
    layer0_outputs(2891) <= not a or b;
    layer0_outputs(2892) <= a;
    layer0_outputs(2893) <= not a or b;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= b and not a;
    layer0_outputs(2896) <= a and not b;
    layer0_outputs(2897) <= not b or a;
    layer0_outputs(2898) <= a or b;
    layer0_outputs(2899) <= not (a and b);
    layer0_outputs(2900) <= not (a or b);
    layer0_outputs(2901) <= a and not b;
    layer0_outputs(2902) <= a or b;
    layer0_outputs(2903) <= a xor b;
    layer0_outputs(2904) <= not (a and b);
    layer0_outputs(2905) <= a xor b;
    layer0_outputs(2906) <= not (a or b);
    layer0_outputs(2907) <= not (a xor b);
    layer0_outputs(2908) <= not (a xor b);
    layer0_outputs(2909) <= b;
    layer0_outputs(2910) <= a;
    layer0_outputs(2911) <= not b or a;
    layer0_outputs(2912) <= not (a xor b);
    layer0_outputs(2913) <= b and not a;
    layer0_outputs(2914) <= b and not a;
    layer0_outputs(2915) <= not (a xor b);
    layer0_outputs(2916) <= a;
    layer0_outputs(2917) <= not b or a;
    layer0_outputs(2918) <= not (a or b);
    layer0_outputs(2919) <= not b or a;
    layer0_outputs(2920) <= a xor b;
    layer0_outputs(2921) <= a or b;
    layer0_outputs(2922) <= 1'b0;
    layer0_outputs(2923) <= not a;
    layer0_outputs(2924) <= a and not b;
    layer0_outputs(2925) <= a xor b;
    layer0_outputs(2926) <= not (a and b);
    layer0_outputs(2927) <= a or b;
    layer0_outputs(2928) <= not a;
    layer0_outputs(2929) <= b and not a;
    layer0_outputs(2930) <= a;
    layer0_outputs(2931) <= b and not a;
    layer0_outputs(2932) <= a or b;
    layer0_outputs(2933) <= b;
    layer0_outputs(2934) <= not b or a;
    layer0_outputs(2935) <= a and not b;
    layer0_outputs(2936) <= b;
    layer0_outputs(2937) <= not b or a;
    layer0_outputs(2938) <= b and not a;
    layer0_outputs(2939) <= not b;
    layer0_outputs(2940) <= not a or b;
    layer0_outputs(2941) <= 1'b0;
    layer0_outputs(2942) <= a;
    layer0_outputs(2943) <= not a or b;
    layer0_outputs(2944) <= a;
    layer0_outputs(2945) <= a or b;
    layer0_outputs(2946) <= b;
    layer0_outputs(2947) <= not (a or b);
    layer0_outputs(2948) <= a and not b;
    layer0_outputs(2949) <= a xor b;
    layer0_outputs(2950) <= a xor b;
    layer0_outputs(2951) <= not (a or b);
    layer0_outputs(2952) <= a;
    layer0_outputs(2953) <= not a;
    layer0_outputs(2954) <= a and not b;
    layer0_outputs(2955) <= not a;
    layer0_outputs(2956) <= a and not b;
    layer0_outputs(2957) <= not a;
    layer0_outputs(2958) <= b and not a;
    layer0_outputs(2959) <= not a or b;
    layer0_outputs(2960) <= a and b;
    layer0_outputs(2961) <= 1'b0;
    layer0_outputs(2962) <= b;
    layer0_outputs(2963) <= a and not b;
    layer0_outputs(2964) <= not a;
    layer0_outputs(2965) <= not a or b;
    layer0_outputs(2966) <= a or b;
    layer0_outputs(2967) <= a;
    layer0_outputs(2968) <= not b;
    layer0_outputs(2969) <= a;
    layer0_outputs(2970) <= a xor b;
    layer0_outputs(2971) <= not (a or b);
    layer0_outputs(2972) <= not (a xor b);
    layer0_outputs(2973) <= not a;
    layer0_outputs(2974) <= a xor b;
    layer0_outputs(2975) <= not b;
    layer0_outputs(2976) <= a and b;
    layer0_outputs(2977) <= a and not b;
    layer0_outputs(2978) <= a or b;
    layer0_outputs(2979) <= a xor b;
    layer0_outputs(2980) <= not (a or b);
    layer0_outputs(2981) <= not a;
    layer0_outputs(2982) <= not a;
    layer0_outputs(2983) <= b and not a;
    layer0_outputs(2984) <= not (a or b);
    layer0_outputs(2985) <= a or b;
    layer0_outputs(2986) <= a or b;
    layer0_outputs(2987) <= not b;
    layer0_outputs(2988) <= a or b;
    layer0_outputs(2989) <= a;
    layer0_outputs(2990) <= not a or b;
    layer0_outputs(2991) <= a;
    layer0_outputs(2992) <= a or b;
    layer0_outputs(2993) <= a xor b;
    layer0_outputs(2994) <= not (a or b);
    layer0_outputs(2995) <= b;
    layer0_outputs(2996) <= not a;
    layer0_outputs(2997) <= not b;
    layer0_outputs(2998) <= a or b;
    layer0_outputs(2999) <= not (a or b);
    layer0_outputs(3000) <= b;
    layer0_outputs(3001) <= b and not a;
    layer0_outputs(3002) <= a or b;
    layer0_outputs(3003) <= not a or b;
    layer0_outputs(3004) <= not (a xor b);
    layer0_outputs(3005) <= a or b;
    layer0_outputs(3006) <= a xor b;
    layer0_outputs(3007) <= not (a or b);
    layer0_outputs(3008) <= not b;
    layer0_outputs(3009) <= not b or a;
    layer0_outputs(3010) <= a and not b;
    layer0_outputs(3011) <= not b;
    layer0_outputs(3012) <= a or b;
    layer0_outputs(3013) <= not b or a;
    layer0_outputs(3014) <= a and b;
    layer0_outputs(3015) <= not (a xor b);
    layer0_outputs(3016) <= a xor b;
    layer0_outputs(3017) <= a or b;
    layer0_outputs(3018) <= not (a or b);
    layer0_outputs(3019) <= not (a and b);
    layer0_outputs(3020) <= not (a xor b);
    layer0_outputs(3021) <= not (a xor b);
    layer0_outputs(3022) <= 1'b0;
    layer0_outputs(3023) <= not a or b;
    layer0_outputs(3024) <= b;
    layer0_outputs(3025) <= b and not a;
    layer0_outputs(3026) <= a or b;
    layer0_outputs(3027) <= not a;
    layer0_outputs(3028) <= 1'b1;
    layer0_outputs(3029) <= a or b;
    layer0_outputs(3030) <= not a or b;
    layer0_outputs(3031) <= b;
    layer0_outputs(3032) <= a and b;
    layer0_outputs(3033) <= not b;
    layer0_outputs(3034) <= a or b;
    layer0_outputs(3035) <= a or b;
    layer0_outputs(3036) <= b and not a;
    layer0_outputs(3037) <= a and b;
    layer0_outputs(3038) <= not (a xor b);
    layer0_outputs(3039) <= a xor b;
    layer0_outputs(3040) <= 1'b0;
    layer0_outputs(3041) <= not a;
    layer0_outputs(3042) <= a xor b;
    layer0_outputs(3043) <= not (a xor b);
    layer0_outputs(3044) <= not b or a;
    layer0_outputs(3045) <= not (a xor b);
    layer0_outputs(3046) <= b and not a;
    layer0_outputs(3047) <= not a;
    layer0_outputs(3048) <= 1'b0;
    layer0_outputs(3049) <= not b or a;
    layer0_outputs(3050) <= a xor b;
    layer0_outputs(3051) <= not a or b;
    layer0_outputs(3052) <= a;
    layer0_outputs(3053) <= not b;
    layer0_outputs(3054) <= not b or a;
    layer0_outputs(3055) <= not (a xor b);
    layer0_outputs(3056) <= b;
    layer0_outputs(3057) <= not (a or b);
    layer0_outputs(3058) <= not b;
    layer0_outputs(3059) <= not b or a;
    layer0_outputs(3060) <= a;
    layer0_outputs(3061) <= a;
    layer0_outputs(3062) <= b and not a;
    layer0_outputs(3063) <= not a;
    layer0_outputs(3064) <= a;
    layer0_outputs(3065) <= a xor b;
    layer0_outputs(3066) <= not a or b;
    layer0_outputs(3067) <= a or b;
    layer0_outputs(3068) <= 1'b0;
    layer0_outputs(3069) <= a xor b;
    layer0_outputs(3070) <= not a;
    layer0_outputs(3071) <= 1'b1;
    layer0_outputs(3072) <= a and b;
    layer0_outputs(3073) <= a xor b;
    layer0_outputs(3074) <= b and not a;
    layer0_outputs(3075) <= a and not b;
    layer0_outputs(3076) <= a xor b;
    layer0_outputs(3077) <= a and not b;
    layer0_outputs(3078) <= a and b;
    layer0_outputs(3079) <= a;
    layer0_outputs(3080) <= not a;
    layer0_outputs(3081) <= not (a or b);
    layer0_outputs(3082) <= not b or a;
    layer0_outputs(3083) <= 1'b0;
    layer0_outputs(3084) <= not a;
    layer0_outputs(3085) <= not b or a;
    layer0_outputs(3086) <= a xor b;
    layer0_outputs(3087) <= a xor b;
    layer0_outputs(3088) <= b and not a;
    layer0_outputs(3089) <= not (a and b);
    layer0_outputs(3090) <= not b;
    layer0_outputs(3091) <= not (a or b);
    layer0_outputs(3092) <= a;
    layer0_outputs(3093) <= a xor b;
    layer0_outputs(3094) <= not a;
    layer0_outputs(3095) <= b and not a;
    layer0_outputs(3096) <= not (a xor b);
    layer0_outputs(3097) <= 1'b1;
    layer0_outputs(3098) <= a;
    layer0_outputs(3099) <= a xor b;
    layer0_outputs(3100) <= not (a and b);
    layer0_outputs(3101) <= a or b;
    layer0_outputs(3102) <= not b;
    layer0_outputs(3103) <= not b;
    layer0_outputs(3104) <= not (a and b);
    layer0_outputs(3105) <= b;
    layer0_outputs(3106) <= a xor b;
    layer0_outputs(3107) <= not (a xor b);
    layer0_outputs(3108) <= b and not a;
    layer0_outputs(3109) <= not (a or b);
    layer0_outputs(3110) <= a xor b;
    layer0_outputs(3111) <= b and not a;
    layer0_outputs(3112) <= not a or b;
    layer0_outputs(3113) <= not a;
    layer0_outputs(3114) <= b;
    layer0_outputs(3115) <= b;
    layer0_outputs(3116) <= a or b;
    layer0_outputs(3117) <= not a or b;
    layer0_outputs(3118) <= a xor b;
    layer0_outputs(3119) <= not a or b;
    layer0_outputs(3120) <= a or b;
    layer0_outputs(3121) <= b;
    layer0_outputs(3122) <= not (a or b);
    layer0_outputs(3123) <= b and not a;
    layer0_outputs(3124) <= not (a or b);
    layer0_outputs(3125) <= a or b;
    layer0_outputs(3126) <= not a or b;
    layer0_outputs(3127) <= b and not a;
    layer0_outputs(3128) <= not a;
    layer0_outputs(3129) <= a and b;
    layer0_outputs(3130) <= a xor b;
    layer0_outputs(3131) <= not b;
    layer0_outputs(3132) <= not a;
    layer0_outputs(3133) <= a;
    layer0_outputs(3134) <= not b or a;
    layer0_outputs(3135) <= not a;
    layer0_outputs(3136) <= not b or a;
    layer0_outputs(3137) <= not a or b;
    layer0_outputs(3138) <= a xor b;
    layer0_outputs(3139) <= not a or b;
    layer0_outputs(3140) <= not a;
    layer0_outputs(3141) <= b and not a;
    layer0_outputs(3142) <= not a;
    layer0_outputs(3143) <= not b;
    layer0_outputs(3144) <= not (a or b);
    layer0_outputs(3145) <= not (a or b);
    layer0_outputs(3146) <= a xor b;
    layer0_outputs(3147) <= a and b;
    layer0_outputs(3148) <= not a;
    layer0_outputs(3149) <= not a or b;
    layer0_outputs(3150) <= b;
    layer0_outputs(3151) <= a;
    layer0_outputs(3152) <= a and not b;
    layer0_outputs(3153) <= not b;
    layer0_outputs(3154) <= b and not a;
    layer0_outputs(3155) <= b;
    layer0_outputs(3156) <= not (a or b);
    layer0_outputs(3157) <= not (a xor b);
    layer0_outputs(3158) <= not a or b;
    layer0_outputs(3159) <= a xor b;
    layer0_outputs(3160) <= a and not b;
    layer0_outputs(3161) <= b;
    layer0_outputs(3162) <= not (a and b);
    layer0_outputs(3163) <= b;
    layer0_outputs(3164) <= not (a or b);
    layer0_outputs(3165) <= not b;
    layer0_outputs(3166) <= not (a xor b);
    layer0_outputs(3167) <= b and not a;
    layer0_outputs(3168) <= a xor b;
    layer0_outputs(3169) <= not (a or b);
    layer0_outputs(3170) <= not (a or b);
    layer0_outputs(3171) <= not b or a;
    layer0_outputs(3172) <= b;
    layer0_outputs(3173) <= not a;
    layer0_outputs(3174) <= a;
    layer0_outputs(3175) <= not (a or b);
    layer0_outputs(3176) <= not (a xor b);
    layer0_outputs(3177) <= a and b;
    layer0_outputs(3178) <= a or b;
    layer0_outputs(3179) <= not (a or b);
    layer0_outputs(3180) <= not (a xor b);
    layer0_outputs(3181) <= b and not a;
    layer0_outputs(3182) <= a xor b;
    layer0_outputs(3183) <= b and not a;
    layer0_outputs(3184) <= not (a xor b);
    layer0_outputs(3185) <= not b;
    layer0_outputs(3186) <= not b;
    layer0_outputs(3187) <= a;
    layer0_outputs(3188) <= not b;
    layer0_outputs(3189) <= b;
    layer0_outputs(3190) <= not (a or b);
    layer0_outputs(3191) <= not (a or b);
    layer0_outputs(3192) <= not (a xor b);
    layer0_outputs(3193) <= not (a or b);
    layer0_outputs(3194) <= a and not b;
    layer0_outputs(3195) <= b;
    layer0_outputs(3196) <= a xor b;
    layer0_outputs(3197) <= not (a xor b);
    layer0_outputs(3198) <= b and not a;
    layer0_outputs(3199) <= not a or b;
    layer0_outputs(3200) <= b and not a;
    layer0_outputs(3201) <= not (a or b);
    layer0_outputs(3202) <= not a or b;
    layer0_outputs(3203) <= b;
    layer0_outputs(3204) <= b;
    layer0_outputs(3205) <= a;
    layer0_outputs(3206) <= a or b;
    layer0_outputs(3207) <= not b or a;
    layer0_outputs(3208) <= a and not b;
    layer0_outputs(3209) <= 1'b0;
    layer0_outputs(3210) <= not (a xor b);
    layer0_outputs(3211) <= a or b;
    layer0_outputs(3212) <= b;
    layer0_outputs(3213) <= not (a and b);
    layer0_outputs(3214) <= a xor b;
    layer0_outputs(3215) <= a or b;
    layer0_outputs(3216) <= not a;
    layer0_outputs(3217) <= a or b;
    layer0_outputs(3218) <= not (a or b);
    layer0_outputs(3219) <= a or b;
    layer0_outputs(3220) <= b;
    layer0_outputs(3221) <= not b;
    layer0_outputs(3222) <= not b;
    layer0_outputs(3223) <= a and b;
    layer0_outputs(3224) <= a or b;
    layer0_outputs(3225) <= not (a or b);
    layer0_outputs(3226) <= 1'b0;
    layer0_outputs(3227) <= a or b;
    layer0_outputs(3228) <= b and not a;
    layer0_outputs(3229) <= not (a xor b);
    layer0_outputs(3230) <= not (a xor b);
    layer0_outputs(3231) <= not (a xor b);
    layer0_outputs(3232) <= not b;
    layer0_outputs(3233) <= not b or a;
    layer0_outputs(3234) <= a xor b;
    layer0_outputs(3235) <= a and not b;
    layer0_outputs(3236) <= not a or b;
    layer0_outputs(3237) <= 1'b1;
    layer0_outputs(3238) <= b;
    layer0_outputs(3239) <= a xor b;
    layer0_outputs(3240) <= not (a or b);
    layer0_outputs(3241) <= a or b;
    layer0_outputs(3242) <= not a;
    layer0_outputs(3243) <= a or b;
    layer0_outputs(3244) <= not (a xor b);
    layer0_outputs(3245) <= 1'b1;
    layer0_outputs(3246) <= not (a and b);
    layer0_outputs(3247) <= a or b;
    layer0_outputs(3248) <= a and not b;
    layer0_outputs(3249) <= a or b;
    layer0_outputs(3250) <= not a;
    layer0_outputs(3251) <= not a;
    layer0_outputs(3252) <= not (a xor b);
    layer0_outputs(3253) <= b;
    layer0_outputs(3254) <= a or b;
    layer0_outputs(3255) <= not (a or b);
    layer0_outputs(3256) <= not a or b;
    layer0_outputs(3257) <= not a or b;
    layer0_outputs(3258) <= a and not b;
    layer0_outputs(3259) <= not (a or b);
    layer0_outputs(3260) <= a and not b;
    layer0_outputs(3261) <= not (a or b);
    layer0_outputs(3262) <= a xor b;
    layer0_outputs(3263) <= not a or b;
    layer0_outputs(3264) <= a and not b;
    layer0_outputs(3265) <= b;
    layer0_outputs(3266) <= a and not b;
    layer0_outputs(3267) <= a and not b;
    layer0_outputs(3268) <= not b or a;
    layer0_outputs(3269) <= a and b;
    layer0_outputs(3270) <= a and b;
    layer0_outputs(3271) <= not b or a;
    layer0_outputs(3272) <= a and b;
    layer0_outputs(3273) <= b;
    layer0_outputs(3274) <= a or b;
    layer0_outputs(3275) <= not b;
    layer0_outputs(3276) <= not b or a;
    layer0_outputs(3277) <= a;
    layer0_outputs(3278) <= not (a or b);
    layer0_outputs(3279) <= not (a or b);
    layer0_outputs(3280) <= not b or a;
    layer0_outputs(3281) <= a or b;
    layer0_outputs(3282) <= b;
    layer0_outputs(3283) <= not a or b;
    layer0_outputs(3284) <= a and not b;
    layer0_outputs(3285) <= not (a or b);
    layer0_outputs(3286) <= not a or b;
    layer0_outputs(3287) <= not (a or b);
    layer0_outputs(3288) <= a;
    layer0_outputs(3289) <= not (a or b);
    layer0_outputs(3290) <= not a;
    layer0_outputs(3291) <= a or b;
    layer0_outputs(3292) <= not b;
    layer0_outputs(3293) <= not (a or b);
    layer0_outputs(3294) <= a or b;
    layer0_outputs(3295) <= not (a or b);
    layer0_outputs(3296) <= a and b;
    layer0_outputs(3297) <= b and not a;
    layer0_outputs(3298) <= b;
    layer0_outputs(3299) <= b;
    layer0_outputs(3300) <= not (a xor b);
    layer0_outputs(3301) <= not a or b;
    layer0_outputs(3302) <= not a or b;
    layer0_outputs(3303) <= a and not b;
    layer0_outputs(3304) <= not b or a;
    layer0_outputs(3305) <= a or b;
    layer0_outputs(3306) <= not (a or b);
    layer0_outputs(3307) <= a xor b;
    layer0_outputs(3308) <= a or b;
    layer0_outputs(3309) <= not b or a;
    layer0_outputs(3310) <= 1'b1;
    layer0_outputs(3311) <= b;
    layer0_outputs(3312) <= not b or a;
    layer0_outputs(3313) <= b and not a;
    layer0_outputs(3314) <= not (a or b);
    layer0_outputs(3315) <= b;
    layer0_outputs(3316) <= a xor b;
    layer0_outputs(3317) <= a or b;
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= not a or b;
    layer0_outputs(3320) <= a and not b;
    layer0_outputs(3321) <= b and not a;
    layer0_outputs(3322) <= not a or b;
    layer0_outputs(3323) <= a or b;
    layer0_outputs(3324) <= a;
    layer0_outputs(3325) <= not a;
    layer0_outputs(3326) <= not a or b;
    layer0_outputs(3327) <= b;
    layer0_outputs(3328) <= a xor b;
    layer0_outputs(3329) <= not b or a;
    layer0_outputs(3330) <= not b;
    layer0_outputs(3331) <= not b;
    layer0_outputs(3332) <= 1'b0;
    layer0_outputs(3333) <= not (a or b);
    layer0_outputs(3334) <= b;
    layer0_outputs(3335) <= a;
    layer0_outputs(3336) <= a or b;
    layer0_outputs(3337) <= b and not a;
    layer0_outputs(3338) <= not (a or b);
    layer0_outputs(3339) <= a and not b;
    layer0_outputs(3340) <= b;
    layer0_outputs(3341) <= a and not b;
    layer0_outputs(3342) <= b;
    layer0_outputs(3343) <= not (a or b);
    layer0_outputs(3344) <= not (a xor b);
    layer0_outputs(3345) <= not b;
    layer0_outputs(3346) <= not a or b;
    layer0_outputs(3347) <= not a;
    layer0_outputs(3348) <= not (a or b);
    layer0_outputs(3349) <= not (a or b);
    layer0_outputs(3350) <= a;
    layer0_outputs(3351) <= a and not b;
    layer0_outputs(3352) <= b;
    layer0_outputs(3353) <= not (a or b);
    layer0_outputs(3354) <= not a or b;
    layer0_outputs(3355) <= b and not a;
    layer0_outputs(3356) <= not (a or b);
    layer0_outputs(3357) <= a and not b;
    layer0_outputs(3358) <= b;
    layer0_outputs(3359) <= not (a xor b);
    layer0_outputs(3360) <= a and not b;
    layer0_outputs(3361) <= not (a xor b);
    layer0_outputs(3362) <= a or b;
    layer0_outputs(3363) <= not b;
    layer0_outputs(3364) <= a and not b;
    layer0_outputs(3365) <= b;
    layer0_outputs(3366) <= b and not a;
    layer0_outputs(3367) <= not b or a;
    layer0_outputs(3368) <= a or b;
    layer0_outputs(3369) <= b and not a;
    layer0_outputs(3370) <= not b;
    layer0_outputs(3371) <= not b;
    layer0_outputs(3372) <= not (a xor b);
    layer0_outputs(3373) <= b and not a;
    layer0_outputs(3374) <= not (a or b);
    layer0_outputs(3375) <= not (a and b);
    layer0_outputs(3376) <= a or b;
    layer0_outputs(3377) <= a or b;
    layer0_outputs(3378) <= a or b;
    layer0_outputs(3379) <= not a or b;
    layer0_outputs(3380) <= not a;
    layer0_outputs(3381) <= not (a or b);
    layer0_outputs(3382) <= a;
    layer0_outputs(3383) <= 1'b1;
    layer0_outputs(3384) <= not (a and b);
    layer0_outputs(3385) <= b;
    layer0_outputs(3386) <= a or b;
    layer0_outputs(3387) <= a or b;
    layer0_outputs(3388) <= a xor b;
    layer0_outputs(3389) <= a xor b;
    layer0_outputs(3390) <= 1'b0;
    layer0_outputs(3391) <= not a;
    layer0_outputs(3392) <= a or b;
    layer0_outputs(3393) <= a xor b;
    layer0_outputs(3394) <= not a or b;
    layer0_outputs(3395) <= not (a xor b);
    layer0_outputs(3396) <= not a;
    layer0_outputs(3397) <= a and not b;
    layer0_outputs(3398) <= not (a or b);
    layer0_outputs(3399) <= a;
    layer0_outputs(3400) <= not a or b;
    layer0_outputs(3401) <= b;
    layer0_outputs(3402) <= not (a xor b);
    layer0_outputs(3403) <= not b or a;
    layer0_outputs(3404) <= not a;
    layer0_outputs(3405) <= not (a and b);
    layer0_outputs(3406) <= not a;
    layer0_outputs(3407) <= b;
    layer0_outputs(3408) <= not b;
    layer0_outputs(3409) <= not b;
    layer0_outputs(3410) <= b and not a;
    layer0_outputs(3411) <= not (a xor b);
    layer0_outputs(3412) <= a or b;
    layer0_outputs(3413) <= a or b;
    layer0_outputs(3414) <= a and b;
    layer0_outputs(3415) <= not (a xor b);
    layer0_outputs(3416) <= a xor b;
    layer0_outputs(3417) <= not a;
    layer0_outputs(3418) <= b and not a;
    layer0_outputs(3419) <= 1'b0;
    layer0_outputs(3420) <= a;
    layer0_outputs(3421) <= b and not a;
    layer0_outputs(3422) <= b and not a;
    layer0_outputs(3423) <= not (a or b);
    layer0_outputs(3424) <= a or b;
    layer0_outputs(3425) <= a and not b;
    layer0_outputs(3426) <= a xor b;
    layer0_outputs(3427) <= not (a xor b);
    layer0_outputs(3428) <= not (a and b);
    layer0_outputs(3429) <= not (a xor b);
    layer0_outputs(3430) <= not (a or b);
    layer0_outputs(3431) <= a and b;
    layer0_outputs(3432) <= a or b;
    layer0_outputs(3433) <= not (a xor b);
    layer0_outputs(3434) <= not (a and b);
    layer0_outputs(3435) <= a and not b;
    layer0_outputs(3436) <= a xor b;
    layer0_outputs(3437) <= a xor b;
    layer0_outputs(3438) <= not a;
    layer0_outputs(3439) <= 1'b1;
    layer0_outputs(3440) <= not a or b;
    layer0_outputs(3441) <= b;
    layer0_outputs(3442) <= b;
    layer0_outputs(3443) <= not (a xor b);
    layer0_outputs(3444) <= 1'b1;
    layer0_outputs(3445) <= a and not b;
    layer0_outputs(3446) <= a and not b;
    layer0_outputs(3447) <= not b;
    layer0_outputs(3448) <= 1'b1;
    layer0_outputs(3449) <= not a;
    layer0_outputs(3450) <= a and not b;
    layer0_outputs(3451) <= not a;
    layer0_outputs(3452) <= a xor b;
    layer0_outputs(3453) <= b;
    layer0_outputs(3454) <= a or b;
    layer0_outputs(3455) <= not a;
    layer0_outputs(3456) <= a or b;
    layer0_outputs(3457) <= not b or a;
    layer0_outputs(3458) <= b and not a;
    layer0_outputs(3459) <= b and not a;
    layer0_outputs(3460) <= b and not a;
    layer0_outputs(3461) <= not b or a;
    layer0_outputs(3462) <= not b or a;
    layer0_outputs(3463) <= a xor b;
    layer0_outputs(3464) <= not a;
    layer0_outputs(3465) <= a or b;
    layer0_outputs(3466) <= not a or b;
    layer0_outputs(3467) <= a or b;
    layer0_outputs(3468) <= a or b;
    layer0_outputs(3469) <= a xor b;
    layer0_outputs(3470) <= 1'b0;
    layer0_outputs(3471) <= a;
    layer0_outputs(3472) <= a and not b;
    layer0_outputs(3473) <= not b or a;
    layer0_outputs(3474) <= not a or b;
    layer0_outputs(3475) <= not (a xor b);
    layer0_outputs(3476) <= a and not b;
    layer0_outputs(3477) <= 1'b1;
    layer0_outputs(3478) <= a xor b;
    layer0_outputs(3479) <= not (a xor b);
    layer0_outputs(3480) <= a and b;
    layer0_outputs(3481) <= not (a xor b);
    layer0_outputs(3482) <= not b;
    layer0_outputs(3483) <= a xor b;
    layer0_outputs(3484) <= not (a xor b);
    layer0_outputs(3485) <= not a or b;
    layer0_outputs(3486) <= a;
    layer0_outputs(3487) <= not (a or b);
    layer0_outputs(3488) <= a or b;
    layer0_outputs(3489) <= a xor b;
    layer0_outputs(3490) <= a xor b;
    layer0_outputs(3491) <= not (a or b);
    layer0_outputs(3492) <= not b;
    layer0_outputs(3493) <= not (a or b);
    layer0_outputs(3494) <= a and not b;
    layer0_outputs(3495) <= not b or a;
    layer0_outputs(3496) <= a and not b;
    layer0_outputs(3497) <= a;
    layer0_outputs(3498) <= not b;
    layer0_outputs(3499) <= not b or a;
    layer0_outputs(3500) <= b;
    layer0_outputs(3501) <= not a;
    layer0_outputs(3502) <= a;
    layer0_outputs(3503) <= b and not a;
    layer0_outputs(3504) <= a or b;
    layer0_outputs(3505) <= not (a or b);
    layer0_outputs(3506) <= 1'b1;
    layer0_outputs(3507) <= b;
    layer0_outputs(3508) <= b;
    layer0_outputs(3509) <= 1'b1;
    layer0_outputs(3510) <= not (a or b);
    layer0_outputs(3511) <= b;
    layer0_outputs(3512) <= not (a xor b);
    layer0_outputs(3513) <= a and b;
    layer0_outputs(3514) <= not a;
    layer0_outputs(3515) <= a or b;
    layer0_outputs(3516) <= b and not a;
    layer0_outputs(3517) <= not (a or b);
    layer0_outputs(3518) <= not (a xor b);
    layer0_outputs(3519) <= not (a or b);
    layer0_outputs(3520) <= a xor b;
    layer0_outputs(3521) <= not b;
    layer0_outputs(3522) <= not a or b;
    layer0_outputs(3523) <= not (a or b);
    layer0_outputs(3524) <= not (a xor b);
    layer0_outputs(3525) <= 1'b0;
    layer0_outputs(3526) <= not a or b;
    layer0_outputs(3527) <= not a;
    layer0_outputs(3528) <= a xor b;
    layer0_outputs(3529) <= b;
    layer0_outputs(3530) <= not (a and b);
    layer0_outputs(3531) <= not (a xor b);
    layer0_outputs(3532) <= b;
    layer0_outputs(3533) <= not (a or b);
    layer0_outputs(3534) <= not (a xor b);
    layer0_outputs(3535) <= a or b;
    layer0_outputs(3536) <= a;
    layer0_outputs(3537) <= not (a xor b);
    layer0_outputs(3538) <= not a;
    layer0_outputs(3539) <= not (a xor b);
    layer0_outputs(3540) <= not (a or b);
    layer0_outputs(3541) <= not a or b;
    layer0_outputs(3542) <= not b or a;
    layer0_outputs(3543) <= a and not b;
    layer0_outputs(3544) <= 1'b0;
    layer0_outputs(3545) <= not a or b;
    layer0_outputs(3546) <= a or b;
    layer0_outputs(3547) <= b and not a;
    layer0_outputs(3548) <= not (a xor b);
    layer0_outputs(3549) <= not (a or b);
    layer0_outputs(3550) <= not b or a;
    layer0_outputs(3551) <= a and not b;
    layer0_outputs(3552) <= not b or a;
    layer0_outputs(3553) <= a xor b;
    layer0_outputs(3554) <= a;
    layer0_outputs(3555) <= 1'b1;
    layer0_outputs(3556) <= not (a or b);
    layer0_outputs(3557) <= not b;
    layer0_outputs(3558) <= not b;
    layer0_outputs(3559) <= b and not a;
    layer0_outputs(3560) <= not (a xor b);
    layer0_outputs(3561) <= not (a xor b);
    layer0_outputs(3562) <= not (a or b);
    layer0_outputs(3563) <= a;
    layer0_outputs(3564) <= 1'b1;
    layer0_outputs(3565) <= 1'b1;
    layer0_outputs(3566) <= not a or b;
    layer0_outputs(3567) <= not (a or b);
    layer0_outputs(3568) <= not (a or b);
    layer0_outputs(3569) <= not a;
    layer0_outputs(3570) <= a and not b;
    layer0_outputs(3571) <= not (a or b);
    layer0_outputs(3572) <= not b;
    layer0_outputs(3573) <= a or b;
    layer0_outputs(3574) <= 1'b0;
    layer0_outputs(3575) <= not (a and b);
    layer0_outputs(3576) <= not (a or b);
    layer0_outputs(3577) <= b;
    layer0_outputs(3578) <= not b;
    layer0_outputs(3579) <= not (a xor b);
    layer0_outputs(3580) <= a and not b;
    layer0_outputs(3581) <= not (a or b);
    layer0_outputs(3582) <= not (a xor b);
    layer0_outputs(3583) <= not (a or b);
    layer0_outputs(3584) <= b and not a;
    layer0_outputs(3585) <= not b;
    layer0_outputs(3586) <= a;
    layer0_outputs(3587) <= b;
    layer0_outputs(3588) <= b and not a;
    layer0_outputs(3589) <= a or b;
    layer0_outputs(3590) <= not a or b;
    layer0_outputs(3591) <= a;
    layer0_outputs(3592) <= a xor b;
    layer0_outputs(3593) <= not b or a;
    layer0_outputs(3594) <= not a or b;
    layer0_outputs(3595) <= a and not b;
    layer0_outputs(3596) <= b;
    layer0_outputs(3597) <= not (a or b);
    layer0_outputs(3598) <= not (a or b);
    layer0_outputs(3599) <= not b or a;
    layer0_outputs(3600) <= a and b;
    layer0_outputs(3601) <= a;
    layer0_outputs(3602) <= a or b;
    layer0_outputs(3603) <= not a or b;
    layer0_outputs(3604) <= a or b;
    layer0_outputs(3605) <= not (a xor b);
    layer0_outputs(3606) <= a or b;
    layer0_outputs(3607) <= not b;
    layer0_outputs(3608) <= not b or a;
    layer0_outputs(3609) <= 1'b0;
    layer0_outputs(3610) <= a xor b;
    layer0_outputs(3611) <= a xor b;
    layer0_outputs(3612) <= b and not a;
    layer0_outputs(3613) <= not b or a;
    layer0_outputs(3614) <= a;
    layer0_outputs(3615) <= a xor b;
    layer0_outputs(3616) <= not (a xor b);
    layer0_outputs(3617) <= b;
    layer0_outputs(3618) <= a;
    layer0_outputs(3619) <= a or b;
    layer0_outputs(3620) <= b;
    layer0_outputs(3621) <= a or b;
    layer0_outputs(3622) <= not (a xor b);
    layer0_outputs(3623) <= not (a or b);
    layer0_outputs(3624) <= a or b;
    layer0_outputs(3625) <= b;
    layer0_outputs(3626) <= 1'b0;
    layer0_outputs(3627) <= b and not a;
    layer0_outputs(3628) <= not (a or b);
    layer0_outputs(3629) <= a or b;
    layer0_outputs(3630) <= 1'b0;
    layer0_outputs(3631) <= not b or a;
    layer0_outputs(3632) <= not (a xor b);
    layer0_outputs(3633) <= a or b;
    layer0_outputs(3634) <= a;
    layer0_outputs(3635) <= not b or a;
    layer0_outputs(3636) <= not (a xor b);
    layer0_outputs(3637) <= not b or a;
    layer0_outputs(3638) <= a;
    layer0_outputs(3639) <= a and b;
    layer0_outputs(3640) <= not a or b;
    layer0_outputs(3641) <= not (a or b);
    layer0_outputs(3642) <= a xor b;
    layer0_outputs(3643) <= a or b;
    layer0_outputs(3644) <= a or b;
    layer0_outputs(3645) <= not (a xor b);
    layer0_outputs(3646) <= a or b;
    layer0_outputs(3647) <= not b or a;
    layer0_outputs(3648) <= not a or b;
    layer0_outputs(3649) <= not (a or b);
    layer0_outputs(3650) <= a and not b;
    layer0_outputs(3651) <= not b;
    layer0_outputs(3652) <= not (a or b);
    layer0_outputs(3653) <= not (a xor b);
    layer0_outputs(3654) <= not a;
    layer0_outputs(3655) <= not (a or b);
    layer0_outputs(3656) <= not a;
    layer0_outputs(3657) <= a or b;
    layer0_outputs(3658) <= not a or b;
    layer0_outputs(3659) <= a xor b;
    layer0_outputs(3660) <= not a or b;
    layer0_outputs(3661) <= not (a xor b);
    layer0_outputs(3662) <= a or b;
    layer0_outputs(3663) <= a;
    layer0_outputs(3664) <= b and not a;
    layer0_outputs(3665) <= a or b;
    layer0_outputs(3666) <= not (a or b);
    layer0_outputs(3667) <= a;
    layer0_outputs(3668) <= 1'b0;
    layer0_outputs(3669) <= a or b;
    layer0_outputs(3670) <= a and b;
    layer0_outputs(3671) <= not a or b;
    layer0_outputs(3672) <= not (a xor b);
    layer0_outputs(3673) <= b and not a;
    layer0_outputs(3674) <= not a;
    layer0_outputs(3675) <= a xor b;
    layer0_outputs(3676) <= a or b;
    layer0_outputs(3677) <= not a or b;
    layer0_outputs(3678) <= not a;
    layer0_outputs(3679) <= not b or a;
    layer0_outputs(3680) <= b and not a;
    layer0_outputs(3681) <= not a;
    layer0_outputs(3682) <= a xor b;
    layer0_outputs(3683) <= a or b;
    layer0_outputs(3684) <= not (a xor b);
    layer0_outputs(3685) <= not (a or b);
    layer0_outputs(3686) <= a and not b;
    layer0_outputs(3687) <= not (a or b);
    layer0_outputs(3688) <= not (a or b);
    layer0_outputs(3689) <= not (a or b);
    layer0_outputs(3690) <= not b or a;
    layer0_outputs(3691) <= b;
    layer0_outputs(3692) <= a xor b;
    layer0_outputs(3693) <= not (a or b);
    layer0_outputs(3694) <= not b or a;
    layer0_outputs(3695) <= not (a or b);
    layer0_outputs(3696) <= not (a or b);
    layer0_outputs(3697) <= a;
    layer0_outputs(3698) <= not b;
    layer0_outputs(3699) <= b and not a;
    layer0_outputs(3700) <= a and b;
    layer0_outputs(3701) <= b;
    layer0_outputs(3702) <= a xor b;
    layer0_outputs(3703) <= b;
    layer0_outputs(3704) <= not b or a;
    layer0_outputs(3705) <= not (a and b);
    layer0_outputs(3706) <= a xor b;
    layer0_outputs(3707) <= a or b;
    layer0_outputs(3708) <= a or b;
    layer0_outputs(3709) <= not b or a;
    layer0_outputs(3710) <= a or b;
    layer0_outputs(3711) <= b;
    layer0_outputs(3712) <= b and not a;
    layer0_outputs(3713) <= a;
    layer0_outputs(3714) <= b;
    layer0_outputs(3715) <= not a or b;
    layer0_outputs(3716) <= a and b;
    layer0_outputs(3717) <= not a or b;
    layer0_outputs(3718) <= not a;
    layer0_outputs(3719) <= a xor b;
    layer0_outputs(3720) <= not (a xor b);
    layer0_outputs(3721) <= not (a xor b);
    layer0_outputs(3722) <= not a;
    layer0_outputs(3723) <= not a;
    layer0_outputs(3724) <= a and not b;
    layer0_outputs(3725) <= a;
    layer0_outputs(3726) <= b;
    layer0_outputs(3727) <= not b or a;
    layer0_outputs(3728) <= not (a and b);
    layer0_outputs(3729) <= a or b;
    layer0_outputs(3730) <= 1'b1;
    layer0_outputs(3731) <= b and not a;
    layer0_outputs(3732) <= 1'b1;
    layer0_outputs(3733) <= not (a or b);
    layer0_outputs(3734) <= a;
    layer0_outputs(3735) <= a xor b;
    layer0_outputs(3736) <= b;
    layer0_outputs(3737) <= not a or b;
    layer0_outputs(3738) <= a;
    layer0_outputs(3739) <= a or b;
    layer0_outputs(3740) <= not a or b;
    layer0_outputs(3741) <= a;
    layer0_outputs(3742) <= a and not b;
    layer0_outputs(3743) <= a and not b;
    layer0_outputs(3744) <= not (a xor b);
    layer0_outputs(3745) <= not a or b;
    layer0_outputs(3746) <= b and not a;
    layer0_outputs(3747) <= not (a or b);
    layer0_outputs(3748) <= 1'b1;
    layer0_outputs(3749) <= not b;
    layer0_outputs(3750) <= b and not a;
    layer0_outputs(3751) <= b;
    layer0_outputs(3752) <= not b or a;
    layer0_outputs(3753) <= b;
    layer0_outputs(3754) <= 1'b1;
    layer0_outputs(3755) <= not a;
    layer0_outputs(3756) <= a and b;
    layer0_outputs(3757) <= not b;
    layer0_outputs(3758) <= a or b;
    layer0_outputs(3759) <= not (a xor b);
    layer0_outputs(3760) <= a or b;
    layer0_outputs(3761) <= a xor b;
    layer0_outputs(3762) <= a or b;
    layer0_outputs(3763) <= not (a xor b);
    layer0_outputs(3764) <= b;
    layer0_outputs(3765) <= b and not a;
    layer0_outputs(3766) <= not b or a;
    layer0_outputs(3767) <= a xor b;
    layer0_outputs(3768) <= b;
    layer0_outputs(3769) <= a;
    layer0_outputs(3770) <= not (a or b);
    layer0_outputs(3771) <= 1'b1;
    layer0_outputs(3772) <= 1'b1;
    layer0_outputs(3773) <= not a;
    layer0_outputs(3774) <= a and not b;
    layer0_outputs(3775) <= a;
    layer0_outputs(3776) <= b;
    layer0_outputs(3777) <= a or b;
    layer0_outputs(3778) <= a xor b;
    layer0_outputs(3779) <= a or b;
    layer0_outputs(3780) <= a and not b;
    layer0_outputs(3781) <= not b;
    layer0_outputs(3782) <= b;
    layer0_outputs(3783) <= a;
    layer0_outputs(3784) <= a or b;
    layer0_outputs(3785) <= not (a xor b);
    layer0_outputs(3786) <= a or b;
    layer0_outputs(3787) <= not a;
    layer0_outputs(3788) <= not a;
    layer0_outputs(3789) <= a;
    layer0_outputs(3790) <= a and b;
    layer0_outputs(3791) <= not (a or b);
    layer0_outputs(3792) <= not a or b;
    layer0_outputs(3793) <= 1'b1;
    layer0_outputs(3794) <= not (a xor b);
    layer0_outputs(3795) <= not (a or b);
    layer0_outputs(3796) <= not (a or b);
    layer0_outputs(3797) <= b;
    layer0_outputs(3798) <= not (a xor b);
    layer0_outputs(3799) <= a and not b;
    layer0_outputs(3800) <= b and not a;
    layer0_outputs(3801) <= a;
    layer0_outputs(3802) <= not b;
    layer0_outputs(3803) <= a xor b;
    layer0_outputs(3804) <= b;
    layer0_outputs(3805) <= a or b;
    layer0_outputs(3806) <= a and b;
    layer0_outputs(3807) <= not (a and b);
    layer0_outputs(3808) <= a xor b;
    layer0_outputs(3809) <= not a;
    layer0_outputs(3810) <= not (a xor b);
    layer0_outputs(3811) <= a and not b;
    layer0_outputs(3812) <= a or b;
    layer0_outputs(3813) <= not b;
    layer0_outputs(3814) <= a or b;
    layer0_outputs(3815) <= a xor b;
    layer0_outputs(3816) <= a or b;
    layer0_outputs(3817) <= a xor b;
    layer0_outputs(3818) <= b and not a;
    layer0_outputs(3819) <= not (a or b);
    layer0_outputs(3820) <= a xor b;
    layer0_outputs(3821) <= not a;
    layer0_outputs(3822) <= a;
    layer0_outputs(3823) <= not (a xor b);
    layer0_outputs(3824) <= b and not a;
    layer0_outputs(3825) <= not a;
    layer0_outputs(3826) <= not a or b;
    layer0_outputs(3827) <= a xor b;
    layer0_outputs(3828) <= not a or b;
    layer0_outputs(3829) <= a xor b;
    layer0_outputs(3830) <= a xor b;
    layer0_outputs(3831) <= not a or b;
    layer0_outputs(3832) <= a or b;
    layer0_outputs(3833) <= a and not b;
    layer0_outputs(3834) <= a;
    layer0_outputs(3835) <= not (a xor b);
    layer0_outputs(3836) <= not (a or b);
    layer0_outputs(3837) <= not (a xor b);
    layer0_outputs(3838) <= not b;
    layer0_outputs(3839) <= not a or b;
    layer0_outputs(3840) <= a xor b;
    layer0_outputs(3841) <= not (a and b);
    layer0_outputs(3842) <= not b;
    layer0_outputs(3843) <= not b or a;
    layer0_outputs(3844) <= a or b;
    layer0_outputs(3845) <= a xor b;
    layer0_outputs(3846) <= not (a xor b);
    layer0_outputs(3847) <= a or b;
    layer0_outputs(3848) <= not (a or b);
    layer0_outputs(3849) <= a or b;
    layer0_outputs(3850) <= a and b;
    layer0_outputs(3851) <= b and not a;
    layer0_outputs(3852) <= a and not b;
    layer0_outputs(3853) <= a or b;
    layer0_outputs(3854) <= not (a xor b);
    layer0_outputs(3855) <= not (a or b);
    layer0_outputs(3856) <= not (a or b);
    layer0_outputs(3857) <= a and b;
    layer0_outputs(3858) <= 1'b1;
    layer0_outputs(3859) <= not (a or b);
    layer0_outputs(3860) <= not a;
    layer0_outputs(3861) <= a or b;
    layer0_outputs(3862) <= a or b;
    layer0_outputs(3863) <= b;
    layer0_outputs(3864) <= b and not a;
    layer0_outputs(3865) <= not a;
    layer0_outputs(3866) <= not a or b;
    layer0_outputs(3867) <= not (a xor b);
    layer0_outputs(3868) <= not (a or b);
    layer0_outputs(3869) <= a xor b;
    layer0_outputs(3870) <= a or b;
    layer0_outputs(3871) <= not b or a;
    layer0_outputs(3872) <= not a;
    layer0_outputs(3873) <= not b;
    layer0_outputs(3874) <= a and not b;
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= not b;
    layer0_outputs(3877) <= b and not a;
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= a and not b;
    layer0_outputs(3880) <= a;
    layer0_outputs(3881) <= not b;
    layer0_outputs(3882) <= a and not b;
    layer0_outputs(3883) <= not (a xor b);
    layer0_outputs(3884) <= a or b;
    layer0_outputs(3885) <= a xor b;
    layer0_outputs(3886) <= a or b;
    layer0_outputs(3887) <= a xor b;
    layer0_outputs(3888) <= not (a or b);
    layer0_outputs(3889) <= not (a or b);
    layer0_outputs(3890) <= a xor b;
    layer0_outputs(3891) <= not a or b;
    layer0_outputs(3892) <= b;
    layer0_outputs(3893) <= not b or a;
    layer0_outputs(3894) <= not (a or b);
    layer0_outputs(3895) <= a;
    layer0_outputs(3896) <= a and not b;
    layer0_outputs(3897) <= not (a xor b);
    layer0_outputs(3898) <= a and not b;
    layer0_outputs(3899) <= not (a or b);
    layer0_outputs(3900) <= a or b;
    layer0_outputs(3901) <= not (a or b);
    layer0_outputs(3902) <= not b;
    layer0_outputs(3903) <= a xor b;
    layer0_outputs(3904) <= not b;
    layer0_outputs(3905) <= not a;
    layer0_outputs(3906) <= not b;
    layer0_outputs(3907) <= not (a xor b);
    layer0_outputs(3908) <= a or b;
    layer0_outputs(3909) <= not (a xor b);
    layer0_outputs(3910) <= not b;
    layer0_outputs(3911) <= b;
    layer0_outputs(3912) <= not a;
    layer0_outputs(3913) <= not (a and b);
    layer0_outputs(3914) <= b;
    layer0_outputs(3915) <= not (a xor b);
    layer0_outputs(3916) <= a and b;
    layer0_outputs(3917) <= a xor b;
    layer0_outputs(3918) <= not a;
    layer0_outputs(3919) <= a or b;
    layer0_outputs(3920) <= not a;
    layer0_outputs(3921) <= not (a xor b);
    layer0_outputs(3922) <= not (a xor b);
    layer0_outputs(3923) <= not (a and b);
    layer0_outputs(3924) <= b;
    layer0_outputs(3925) <= not b or a;
    layer0_outputs(3926) <= not (a or b);
    layer0_outputs(3927) <= a or b;
    layer0_outputs(3928) <= not a or b;
    layer0_outputs(3929) <= a;
    layer0_outputs(3930) <= a or b;
    layer0_outputs(3931) <= not (a or b);
    layer0_outputs(3932) <= a;
    layer0_outputs(3933) <= not b;
    layer0_outputs(3934) <= not a;
    layer0_outputs(3935) <= a and not b;
    layer0_outputs(3936) <= b and not a;
    layer0_outputs(3937) <= not b or a;
    layer0_outputs(3938) <= a and not b;
    layer0_outputs(3939) <= a xor b;
    layer0_outputs(3940) <= a and b;
    layer0_outputs(3941) <= not (a or b);
    layer0_outputs(3942) <= a and b;
    layer0_outputs(3943) <= 1'b0;
    layer0_outputs(3944) <= a and not b;
    layer0_outputs(3945) <= not a or b;
    layer0_outputs(3946) <= b;
    layer0_outputs(3947) <= a or b;
    layer0_outputs(3948) <= b and not a;
    layer0_outputs(3949) <= not b or a;
    layer0_outputs(3950) <= a and b;
    layer0_outputs(3951) <= not b or a;
    layer0_outputs(3952) <= b and not a;
    layer0_outputs(3953) <= a or b;
    layer0_outputs(3954) <= b;
    layer0_outputs(3955) <= not a;
    layer0_outputs(3956) <= not b;
    layer0_outputs(3957) <= 1'b0;
    layer0_outputs(3958) <= not (a and b);
    layer0_outputs(3959) <= a or b;
    layer0_outputs(3960) <= not a;
    layer0_outputs(3961) <= not b or a;
    layer0_outputs(3962) <= not a;
    layer0_outputs(3963) <= 1'b0;
    layer0_outputs(3964) <= b;
    layer0_outputs(3965) <= a and b;
    layer0_outputs(3966) <= not b or a;
    layer0_outputs(3967) <= not b or a;
    layer0_outputs(3968) <= a;
    layer0_outputs(3969) <= b and not a;
    layer0_outputs(3970) <= not b or a;
    layer0_outputs(3971) <= not a or b;
    layer0_outputs(3972) <= not b or a;
    layer0_outputs(3973) <= 1'b0;
    layer0_outputs(3974) <= not b or a;
    layer0_outputs(3975) <= a and b;
    layer0_outputs(3976) <= not (a xor b);
    layer0_outputs(3977) <= not a;
    layer0_outputs(3978) <= b;
    layer0_outputs(3979) <= a xor b;
    layer0_outputs(3980) <= 1'b0;
    layer0_outputs(3981) <= b and not a;
    layer0_outputs(3982) <= a or b;
    layer0_outputs(3983) <= a or b;
    layer0_outputs(3984) <= not b or a;
    layer0_outputs(3985) <= not b or a;
    layer0_outputs(3986) <= not b;
    layer0_outputs(3987) <= not b or a;
    layer0_outputs(3988) <= a;
    layer0_outputs(3989) <= b;
    layer0_outputs(3990) <= b;
    layer0_outputs(3991) <= a or b;
    layer0_outputs(3992) <= not (a or b);
    layer0_outputs(3993) <= a xor b;
    layer0_outputs(3994) <= 1'b0;
    layer0_outputs(3995) <= not a or b;
    layer0_outputs(3996) <= a or b;
    layer0_outputs(3997) <= not a;
    layer0_outputs(3998) <= not (a xor b);
    layer0_outputs(3999) <= a xor b;
    layer0_outputs(4000) <= a or b;
    layer0_outputs(4001) <= not (a or b);
    layer0_outputs(4002) <= not b;
    layer0_outputs(4003) <= b and not a;
    layer0_outputs(4004) <= a xor b;
    layer0_outputs(4005) <= not b or a;
    layer0_outputs(4006) <= not b;
    layer0_outputs(4007) <= not a;
    layer0_outputs(4008) <= a and not b;
    layer0_outputs(4009) <= a and not b;
    layer0_outputs(4010) <= b;
    layer0_outputs(4011) <= not (a and b);
    layer0_outputs(4012) <= not a;
    layer0_outputs(4013) <= not b;
    layer0_outputs(4014) <= not a;
    layer0_outputs(4015) <= not (a or b);
    layer0_outputs(4016) <= b and not a;
    layer0_outputs(4017) <= a and not b;
    layer0_outputs(4018) <= not a or b;
    layer0_outputs(4019) <= a;
    layer0_outputs(4020) <= not b or a;
    layer0_outputs(4021) <= a and not b;
    layer0_outputs(4022) <= a or b;
    layer0_outputs(4023) <= not b or a;
    layer0_outputs(4024) <= not (a xor b);
    layer0_outputs(4025) <= not b or a;
    layer0_outputs(4026) <= not b or a;
    layer0_outputs(4027) <= not (a xor b);
    layer0_outputs(4028) <= not b or a;
    layer0_outputs(4029) <= 1'b1;
    layer0_outputs(4030) <= a and not b;
    layer0_outputs(4031) <= not (a or b);
    layer0_outputs(4032) <= b and not a;
    layer0_outputs(4033) <= not a;
    layer0_outputs(4034) <= not a;
    layer0_outputs(4035) <= b and not a;
    layer0_outputs(4036) <= a xor b;
    layer0_outputs(4037) <= not a or b;
    layer0_outputs(4038) <= a or b;
    layer0_outputs(4039) <= 1'b0;
    layer0_outputs(4040) <= a xor b;
    layer0_outputs(4041) <= 1'b1;
    layer0_outputs(4042) <= not (a or b);
    layer0_outputs(4043) <= a or b;
    layer0_outputs(4044) <= a and b;
    layer0_outputs(4045) <= not a or b;
    layer0_outputs(4046) <= a or b;
    layer0_outputs(4047) <= not b or a;
    layer0_outputs(4048) <= not b or a;
    layer0_outputs(4049) <= b;
    layer0_outputs(4050) <= a or b;
    layer0_outputs(4051) <= not b or a;
    layer0_outputs(4052) <= not (a xor b);
    layer0_outputs(4053) <= not (a or b);
    layer0_outputs(4054) <= a or b;
    layer0_outputs(4055) <= not (a or b);
    layer0_outputs(4056) <= 1'b1;
    layer0_outputs(4057) <= not (a xor b);
    layer0_outputs(4058) <= not b;
    layer0_outputs(4059) <= a or b;
    layer0_outputs(4060) <= a and not b;
    layer0_outputs(4061) <= not b or a;
    layer0_outputs(4062) <= a or b;
    layer0_outputs(4063) <= a xor b;
    layer0_outputs(4064) <= a or b;
    layer0_outputs(4065) <= not (a and b);
    layer0_outputs(4066) <= not b or a;
    layer0_outputs(4067) <= not b or a;
    layer0_outputs(4068) <= not (a or b);
    layer0_outputs(4069) <= a;
    layer0_outputs(4070) <= b and not a;
    layer0_outputs(4071) <= b;
    layer0_outputs(4072) <= not b or a;
    layer0_outputs(4073) <= a xor b;
    layer0_outputs(4074) <= a and b;
    layer0_outputs(4075) <= not b or a;
    layer0_outputs(4076) <= a and not b;
    layer0_outputs(4077) <= 1'b1;
    layer0_outputs(4078) <= a xor b;
    layer0_outputs(4079) <= a xor b;
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= not a or b;
    layer0_outputs(4082) <= not (a xor b);
    layer0_outputs(4083) <= a and b;
    layer0_outputs(4084) <= b;
    layer0_outputs(4085) <= not a;
    layer0_outputs(4086) <= not (a or b);
    layer0_outputs(4087) <= not a or b;
    layer0_outputs(4088) <= not b;
    layer0_outputs(4089) <= not b or a;
    layer0_outputs(4090) <= not (a xor b);
    layer0_outputs(4091) <= a or b;
    layer0_outputs(4092) <= b and not a;
    layer0_outputs(4093) <= not b;
    layer0_outputs(4094) <= not (a xor b);
    layer0_outputs(4095) <= not a;
    layer0_outputs(4096) <= b;
    layer0_outputs(4097) <= not a;
    layer0_outputs(4098) <= not a;
    layer0_outputs(4099) <= 1'b1;
    layer0_outputs(4100) <= a xor b;
    layer0_outputs(4101) <= not b;
    layer0_outputs(4102) <= not (a xor b);
    layer0_outputs(4103) <= not (a or b);
    layer0_outputs(4104) <= not (a or b);
    layer0_outputs(4105) <= b and not a;
    layer0_outputs(4106) <= not (a xor b);
    layer0_outputs(4107) <= not (a xor b);
    layer0_outputs(4108) <= b;
    layer0_outputs(4109) <= a and not b;
    layer0_outputs(4110) <= not (a or b);
    layer0_outputs(4111) <= b and not a;
    layer0_outputs(4112) <= a xor b;
    layer0_outputs(4113) <= a;
    layer0_outputs(4114) <= not a or b;
    layer0_outputs(4115) <= not (a or b);
    layer0_outputs(4116) <= not (a or b);
    layer0_outputs(4117) <= a and b;
    layer0_outputs(4118) <= not a;
    layer0_outputs(4119) <= a or b;
    layer0_outputs(4120) <= not a;
    layer0_outputs(4121) <= a;
    layer0_outputs(4122) <= b and not a;
    layer0_outputs(4123) <= not (a and b);
    layer0_outputs(4124) <= a xor b;
    layer0_outputs(4125) <= b and not a;
    layer0_outputs(4126) <= not (a or b);
    layer0_outputs(4127) <= 1'b1;
    layer0_outputs(4128) <= not (a or b);
    layer0_outputs(4129) <= a;
    layer0_outputs(4130) <= not (a and b);
    layer0_outputs(4131) <= not b;
    layer0_outputs(4132) <= a and not b;
    layer0_outputs(4133) <= a or b;
    layer0_outputs(4134) <= b and not a;
    layer0_outputs(4135) <= not (a xor b);
    layer0_outputs(4136) <= a xor b;
    layer0_outputs(4137) <= not a or b;
    layer0_outputs(4138) <= b and not a;
    layer0_outputs(4139) <= not a or b;
    layer0_outputs(4140) <= 1'b0;
    layer0_outputs(4141) <= b and not a;
    layer0_outputs(4142) <= 1'b1;
    layer0_outputs(4143) <= not (a or b);
    layer0_outputs(4144) <= not a or b;
    layer0_outputs(4145) <= a;
    layer0_outputs(4146) <= not b or a;
    layer0_outputs(4147) <= not b;
    layer0_outputs(4148) <= a and not b;
    layer0_outputs(4149) <= a;
    layer0_outputs(4150) <= b;
    layer0_outputs(4151) <= not a or b;
    layer0_outputs(4152) <= a xor b;
    layer0_outputs(4153) <= not (a xor b);
    layer0_outputs(4154) <= not a;
    layer0_outputs(4155) <= a and b;
    layer0_outputs(4156) <= a and not b;
    layer0_outputs(4157) <= a xor b;
    layer0_outputs(4158) <= b and not a;
    layer0_outputs(4159) <= not (a or b);
    layer0_outputs(4160) <= a or b;
    layer0_outputs(4161) <= not (a or b);
    layer0_outputs(4162) <= not (a xor b);
    layer0_outputs(4163) <= b and not a;
    layer0_outputs(4164) <= b;
    layer0_outputs(4165) <= not (a xor b);
    layer0_outputs(4166) <= b;
    layer0_outputs(4167) <= a or b;
    layer0_outputs(4168) <= a and b;
    layer0_outputs(4169) <= a;
    layer0_outputs(4170) <= not (a or b);
    layer0_outputs(4171) <= not (a or b);
    layer0_outputs(4172) <= not b or a;
    layer0_outputs(4173) <= not (a or b);
    layer0_outputs(4174) <= not (a or b);
    layer0_outputs(4175) <= b;
    layer0_outputs(4176) <= a xor b;
    layer0_outputs(4177) <= a and not b;
    layer0_outputs(4178) <= b and not a;
    layer0_outputs(4179) <= a;
    layer0_outputs(4180) <= not (a or b);
    layer0_outputs(4181) <= a and not b;
    layer0_outputs(4182) <= not (a or b);
    layer0_outputs(4183) <= b and not a;
    layer0_outputs(4184) <= not (a xor b);
    layer0_outputs(4185) <= not (a or b);
    layer0_outputs(4186) <= not (a or b);
    layer0_outputs(4187) <= b;
    layer0_outputs(4188) <= not (a xor b);
    layer0_outputs(4189) <= b and not a;
    layer0_outputs(4190) <= not (a or b);
    layer0_outputs(4191) <= not b or a;
    layer0_outputs(4192) <= not (a xor b);
    layer0_outputs(4193) <= not (a and b);
    layer0_outputs(4194) <= not (a and b);
    layer0_outputs(4195) <= 1'b0;
    layer0_outputs(4196) <= a or b;
    layer0_outputs(4197) <= b;
    layer0_outputs(4198) <= a xor b;
    layer0_outputs(4199) <= a xor b;
    layer0_outputs(4200) <= not (a or b);
    layer0_outputs(4201) <= not (a and b);
    layer0_outputs(4202) <= not (a and b);
    layer0_outputs(4203) <= not b or a;
    layer0_outputs(4204) <= 1'b1;
    layer0_outputs(4205) <= a and not b;
    layer0_outputs(4206) <= b;
    layer0_outputs(4207) <= 1'b0;
    layer0_outputs(4208) <= a and not b;
    layer0_outputs(4209) <= not (a and b);
    layer0_outputs(4210) <= not (a xor b);
    layer0_outputs(4211) <= not (a or b);
    layer0_outputs(4212) <= not b or a;
    layer0_outputs(4213) <= a or b;
    layer0_outputs(4214) <= not (a or b);
    layer0_outputs(4215) <= not b or a;
    layer0_outputs(4216) <= a and not b;
    layer0_outputs(4217) <= a xor b;
    layer0_outputs(4218) <= a or b;
    layer0_outputs(4219) <= not (a and b);
    layer0_outputs(4220) <= not a;
    layer0_outputs(4221) <= b;
    layer0_outputs(4222) <= a and not b;
    layer0_outputs(4223) <= not (a xor b);
    layer0_outputs(4224) <= not b or a;
    layer0_outputs(4225) <= a or b;
    layer0_outputs(4226) <= a or b;
    layer0_outputs(4227) <= not (a or b);
    layer0_outputs(4228) <= a and not b;
    layer0_outputs(4229) <= not (a or b);
    layer0_outputs(4230) <= not (a or b);
    layer0_outputs(4231) <= b;
    layer0_outputs(4232) <= not a;
    layer0_outputs(4233) <= not a;
    layer0_outputs(4234) <= not a;
    layer0_outputs(4235) <= a and b;
    layer0_outputs(4236) <= a or b;
    layer0_outputs(4237) <= a or b;
    layer0_outputs(4238) <= a xor b;
    layer0_outputs(4239) <= not (a or b);
    layer0_outputs(4240) <= 1'b1;
    layer0_outputs(4241) <= a and not b;
    layer0_outputs(4242) <= b and not a;
    layer0_outputs(4243) <= not (a and b);
    layer0_outputs(4244) <= not (a or b);
    layer0_outputs(4245) <= not (a or b);
    layer0_outputs(4246) <= a or b;
    layer0_outputs(4247) <= a or b;
    layer0_outputs(4248) <= not (a xor b);
    layer0_outputs(4249) <= not (a or b);
    layer0_outputs(4250) <= not b;
    layer0_outputs(4251) <= a xor b;
    layer0_outputs(4252) <= b and not a;
    layer0_outputs(4253) <= 1'b1;
    layer0_outputs(4254) <= b and not a;
    layer0_outputs(4255) <= a;
    layer0_outputs(4256) <= a xor b;
    layer0_outputs(4257) <= not b or a;
    layer0_outputs(4258) <= not a;
    layer0_outputs(4259) <= not (a xor b);
    layer0_outputs(4260) <= not a or b;
    layer0_outputs(4261) <= b;
    layer0_outputs(4262) <= not b;
    layer0_outputs(4263) <= not a;
    layer0_outputs(4264) <= not b or a;
    layer0_outputs(4265) <= not a;
    layer0_outputs(4266) <= a and not b;
    layer0_outputs(4267) <= not (a xor b);
    layer0_outputs(4268) <= not a or b;
    layer0_outputs(4269) <= not (a xor b);
    layer0_outputs(4270) <= not (a xor b);
    layer0_outputs(4271) <= b and not a;
    layer0_outputs(4272) <= a;
    layer0_outputs(4273) <= a or b;
    layer0_outputs(4274) <= not (a xor b);
    layer0_outputs(4275) <= not (a xor b);
    layer0_outputs(4276) <= not a;
    layer0_outputs(4277) <= not (a or b);
    layer0_outputs(4278) <= 1'b0;
    layer0_outputs(4279) <= not a;
    layer0_outputs(4280) <= a and b;
    layer0_outputs(4281) <= b;
    layer0_outputs(4282) <= b and not a;
    layer0_outputs(4283) <= not b or a;
    layer0_outputs(4284) <= b;
    layer0_outputs(4285) <= a and not b;
    layer0_outputs(4286) <= not a or b;
    layer0_outputs(4287) <= not (a xor b);
    layer0_outputs(4288) <= b;
    layer0_outputs(4289) <= not a or b;
    layer0_outputs(4290) <= not (a or b);
    layer0_outputs(4291) <= b;
    layer0_outputs(4292) <= not (a or b);
    layer0_outputs(4293) <= not a or b;
    layer0_outputs(4294) <= not b or a;
    layer0_outputs(4295) <= not b or a;
    layer0_outputs(4296) <= a;
    layer0_outputs(4297) <= b;
    layer0_outputs(4298) <= not a or b;
    layer0_outputs(4299) <= a or b;
    layer0_outputs(4300) <= not b or a;
    layer0_outputs(4301) <= not b;
    layer0_outputs(4302) <= a and b;
    layer0_outputs(4303) <= a;
    layer0_outputs(4304) <= a;
    layer0_outputs(4305) <= not (a or b);
    layer0_outputs(4306) <= not (a or b);
    layer0_outputs(4307) <= 1'b1;
    layer0_outputs(4308) <= not b or a;
    layer0_outputs(4309) <= not (a or b);
    layer0_outputs(4310) <= not a or b;
    layer0_outputs(4311) <= a xor b;
    layer0_outputs(4312) <= not b;
    layer0_outputs(4313) <= b;
    layer0_outputs(4314) <= b and not a;
    layer0_outputs(4315) <= a xor b;
    layer0_outputs(4316) <= a;
    layer0_outputs(4317) <= not b;
    layer0_outputs(4318) <= not (a xor b);
    layer0_outputs(4319) <= a xor b;
    layer0_outputs(4320) <= not (a xor b);
    layer0_outputs(4321) <= not b or a;
    layer0_outputs(4322) <= not (a xor b);
    layer0_outputs(4323) <= b;
    layer0_outputs(4324) <= not a;
    layer0_outputs(4325) <= b and not a;
    layer0_outputs(4326) <= b and not a;
    layer0_outputs(4327) <= not (a or b);
    layer0_outputs(4328) <= a or b;
    layer0_outputs(4329) <= a xor b;
    layer0_outputs(4330) <= not (a or b);
    layer0_outputs(4331) <= not (a xor b);
    layer0_outputs(4332) <= b;
    layer0_outputs(4333) <= not b or a;
    layer0_outputs(4334) <= a or b;
    layer0_outputs(4335) <= not (a or b);
    layer0_outputs(4336) <= not b;
    layer0_outputs(4337) <= not a;
    layer0_outputs(4338) <= a xor b;
    layer0_outputs(4339) <= not (a xor b);
    layer0_outputs(4340) <= a xor b;
    layer0_outputs(4341) <= a and not b;
    layer0_outputs(4342) <= not (a and b);
    layer0_outputs(4343) <= not (a or b);
    layer0_outputs(4344) <= not (a xor b);
    layer0_outputs(4345) <= b and not a;
    layer0_outputs(4346) <= b and not a;
    layer0_outputs(4347) <= not a;
    layer0_outputs(4348) <= not b;
    layer0_outputs(4349) <= b and not a;
    layer0_outputs(4350) <= not b or a;
    layer0_outputs(4351) <= a xor b;
    layer0_outputs(4352) <= not (a and b);
    layer0_outputs(4353) <= a and not b;
    layer0_outputs(4354) <= a xor b;
    layer0_outputs(4355) <= not (a or b);
    layer0_outputs(4356) <= not a or b;
    layer0_outputs(4357) <= not (a or b);
    layer0_outputs(4358) <= not (a and b);
    layer0_outputs(4359) <= not (a or b);
    layer0_outputs(4360) <= a and not b;
    layer0_outputs(4361) <= a;
    layer0_outputs(4362) <= a and not b;
    layer0_outputs(4363) <= a and not b;
    layer0_outputs(4364) <= not (a xor b);
    layer0_outputs(4365) <= a xor b;
    layer0_outputs(4366) <= a xor b;
    layer0_outputs(4367) <= not (a xor b);
    layer0_outputs(4368) <= b and not a;
    layer0_outputs(4369) <= not b;
    layer0_outputs(4370) <= a and not b;
    layer0_outputs(4371) <= not b;
    layer0_outputs(4372) <= a;
    layer0_outputs(4373) <= not (a xor b);
    layer0_outputs(4374) <= a or b;
    layer0_outputs(4375) <= not a;
    layer0_outputs(4376) <= b;
    layer0_outputs(4377) <= not (a xor b);
    layer0_outputs(4378) <= not b or a;
    layer0_outputs(4379) <= 1'b1;
    layer0_outputs(4380) <= not a;
    layer0_outputs(4381) <= b;
    layer0_outputs(4382) <= a xor b;
    layer0_outputs(4383) <= 1'b0;
    layer0_outputs(4384) <= a or b;
    layer0_outputs(4385) <= not (a xor b);
    layer0_outputs(4386) <= not (a and b);
    layer0_outputs(4387) <= a and not b;
    layer0_outputs(4388) <= a xor b;
    layer0_outputs(4389) <= a and not b;
    layer0_outputs(4390) <= a and not b;
    layer0_outputs(4391) <= b;
    layer0_outputs(4392) <= a or b;
    layer0_outputs(4393) <= a;
    layer0_outputs(4394) <= b and not a;
    layer0_outputs(4395) <= not (a or b);
    layer0_outputs(4396) <= a and b;
    layer0_outputs(4397) <= a or b;
    layer0_outputs(4398) <= not a or b;
    layer0_outputs(4399) <= a and not b;
    layer0_outputs(4400) <= a;
    layer0_outputs(4401) <= b;
    layer0_outputs(4402) <= not (a or b);
    layer0_outputs(4403) <= b;
    layer0_outputs(4404) <= not (a or b);
    layer0_outputs(4405) <= not (a or b);
    layer0_outputs(4406) <= 1'b1;
    layer0_outputs(4407) <= a;
    layer0_outputs(4408) <= b;
    layer0_outputs(4409) <= not a or b;
    layer0_outputs(4410) <= b and not a;
    layer0_outputs(4411) <= not (a xor b);
    layer0_outputs(4412) <= not b;
    layer0_outputs(4413) <= a and b;
    layer0_outputs(4414) <= b and not a;
    layer0_outputs(4415) <= not (a or b);
    layer0_outputs(4416) <= not (a xor b);
    layer0_outputs(4417) <= a;
    layer0_outputs(4418) <= b;
    layer0_outputs(4419) <= not a;
    layer0_outputs(4420) <= a or b;
    layer0_outputs(4421) <= not (a xor b);
    layer0_outputs(4422) <= not a;
    layer0_outputs(4423) <= not (a or b);
    layer0_outputs(4424) <= 1'b1;
    layer0_outputs(4425) <= not (a xor b);
    layer0_outputs(4426) <= not a;
    layer0_outputs(4427) <= b and not a;
    layer0_outputs(4428) <= a or b;
    layer0_outputs(4429) <= not b;
    layer0_outputs(4430) <= not a;
    layer0_outputs(4431) <= a or b;
    layer0_outputs(4432) <= not (a or b);
    layer0_outputs(4433) <= 1'b1;
    layer0_outputs(4434) <= a or b;
    layer0_outputs(4435) <= not (a or b);
    layer0_outputs(4436) <= not a;
    layer0_outputs(4437) <= a and not b;
    layer0_outputs(4438) <= a or b;
    layer0_outputs(4439) <= not (a and b);
    layer0_outputs(4440) <= a;
    layer0_outputs(4441) <= not b;
    layer0_outputs(4442) <= a and b;
    layer0_outputs(4443) <= a or b;
    layer0_outputs(4444) <= a;
    layer0_outputs(4445) <= not (a xor b);
    layer0_outputs(4446) <= a;
    layer0_outputs(4447) <= not b or a;
    layer0_outputs(4448) <= a xor b;
    layer0_outputs(4449) <= a and not b;
    layer0_outputs(4450) <= a and b;
    layer0_outputs(4451) <= a and b;
    layer0_outputs(4452) <= a and not b;
    layer0_outputs(4453) <= a;
    layer0_outputs(4454) <= not b;
    layer0_outputs(4455) <= not b or a;
    layer0_outputs(4456) <= not (a xor b);
    layer0_outputs(4457) <= not (a or b);
    layer0_outputs(4458) <= not b;
    layer0_outputs(4459) <= a xor b;
    layer0_outputs(4460) <= a or b;
    layer0_outputs(4461) <= 1'b0;
    layer0_outputs(4462) <= not a;
    layer0_outputs(4463) <= not (a or b);
    layer0_outputs(4464) <= a xor b;
    layer0_outputs(4465) <= a;
    layer0_outputs(4466) <= a xor b;
    layer0_outputs(4467) <= b and not a;
    layer0_outputs(4468) <= 1'b0;
    layer0_outputs(4469) <= not b or a;
    layer0_outputs(4470) <= b and not a;
    layer0_outputs(4471) <= a or b;
    layer0_outputs(4472) <= not a or b;
    layer0_outputs(4473) <= not b or a;
    layer0_outputs(4474) <= a;
    layer0_outputs(4475) <= b;
    layer0_outputs(4476) <= a;
    layer0_outputs(4477) <= not b or a;
    layer0_outputs(4478) <= b;
    layer0_outputs(4479) <= a;
    layer0_outputs(4480) <= not (a xor b);
    layer0_outputs(4481) <= a or b;
    layer0_outputs(4482) <= not (a or b);
    layer0_outputs(4483) <= not a or b;
    layer0_outputs(4484) <= not b or a;
    layer0_outputs(4485) <= not a;
    layer0_outputs(4486) <= a xor b;
    layer0_outputs(4487) <= a xor b;
    layer0_outputs(4488) <= not (a or b);
    layer0_outputs(4489) <= not b or a;
    layer0_outputs(4490) <= 1'b1;
    layer0_outputs(4491) <= not b;
    layer0_outputs(4492) <= not b or a;
    layer0_outputs(4493) <= b and not a;
    layer0_outputs(4494) <= not (a xor b);
    layer0_outputs(4495) <= not b;
    layer0_outputs(4496) <= 1'b0;
    layer0_outputs(4497) <= a or b;
    layer0_outputs(4498) <= b;
    layer0_outputs(4499) <= not b;
    layer0_outputs(4500) <= a or b;
    layer0_outputs(4501) <= b;
    layer0_outputs(4502) <= not (a xor b);
    layer0_outputs(4503) <= 1'b1;
    layer0_outputs(4504) <= 1'b0;
    layer0_outputs(4505) <= a or b;
    layer0_outputs(4506) <= not (a xor b);
    layer0_outputs(4507) <= a;
    layer0_outputs(4508) <= not (a xor b);
    layer0_outputs(4509) <= not a or b;
    layer0_outputs(4510) <= a;
    layer0_outputs(4511) <= b;
    layer0_outputs(4512) <= a and not b;
    layer0_outputs(4513) <= a or b;
    layer0_outputs(4514) <= 1'b1;
    layer0_outputs(4515) <= a xor b;
    layer0_outputs(4516) <= a and not b;
    layer0_outputs(4517) <= b;
    layer0_outputs(4518) <= a and not b;
    layer0_outputs(4519) <= not (a or b);
    layer0_outputs(4520) <= b;
    layer0_outputs(4521) <= a;
    layer0_outputs(4522) <= not (a xor b);
    layer0_outputs(4523) <= a or b;
    layer0_outputs(4524) <= a;
    layer0_outputs(4525) <= a or b;
    layer0_outputs(4526) <= 1'b1;
    layer0_outputs(4527) <= not a;
    layer0_outputs(4528) <= not (a xor b);
    layer0_outputs(4529) <= 1'b0;
    layer0_outputs(4530) <= a xor b;
    layer0_outputs(4531) <= a;
    layer0_outputs(4532) <= a;
    layer0_outputs(4533) <= not a;
    layer0_outputs(4534) <= a and not b;
    layer0_outputs(4535) <= b;
    layer0_outputs(4536) <= not (a or b);
    layer0_outputs(4537) <= not b;
    layer0_outputs(4538) <= not (a xor b);
    layer0_outputs(4539) <= b;
    layer0_outputs(4540) <= a or b;
    layer0_outputs(4541) <= not (a and b);
    layer0_outputs(4542) <= not (a or b);
    layer0_outputs(4543) <= not (a or b);
    layer0_outputs(4544) <= not a;
    layer0_outputs(4545) <= a and b;
    layer0_outputs(4546) <= not b or a;
    layer0_outputs(4547) <= a or b;
    layer0_outputs(4548) <= not (a xor b);
    layer0_outputs(4549) <= b;
    layer0_outputs(4550) <= a;
    layer0_outputs(4551) <= b and not a;
    layer0_outputs(4552) <= a and not b;
    layer0_outputs(4553) <= not b or a;
    layer0_outputs(4554) <= a or b;
    layer0_outputs(4555) <= a xor b;
    layer0_outputs(4556) <= b and not a;
    layer0_outputs(4557) <= not (a and b);
    layer0_outputs(4558) <= not b;
    layer0_outputs(4559) <= not (a or b);
    layer0_outputs(4560) <= a xor b;
    layer0_outputs(4561) <= not (a or b);
    layer0_outputs(4562) <= not a;
    layer0_outputs(4563) <= a xor b;
    layer0_outputs(4564) <= b and not a;
    layer0_outputs(4565) <= not b or a;
    layer0_outputs(4566) <= b and not a;
    layer0_outputs(4567) <= not b or a;
    layer0_outputs(4568) <= a xor b;
    layer0_outputs(4569) <= not a or b;
    layer0_outputs(4570) <= not (a xor b);
    layer0_outputs(4571) <= b;
    layer0_outputs(4572) <= not (a or b);
    layer0_outputs(4573) <= a xor b;
    layer0_outputs(4574) <= not a or b;
    layer0_outputs(4575) <= not a or b;
    layer0_outputs(4576) <= not a or b;
    layer0_outputs(4577) <= a xor b;
    layer0_outputs(4578) <= a or b;
    layer0_outputs(4579) <= not b;
    layer0_outputs(4580) <= not b;
    layer0_outputs(4581) <= not (a xor b);
    layer0_outputs(4582) <= not (a or b);
    layer0_outputs(4583) <= not b;
    layer0_outputs(4584) <= a xor b;
    layer0_outputs(4585) <= a xor b;
    layer0_outputs(4586) <= not a;
    layer0_outputs(4587) <= not b or a;
    layer0_outputs(4588) <= not b or a;
    layer0_outputs(4589) <= a xor b;
    layer0_outputs(4590) <= not a;
    layer0_outputs(4591) <= a and not b;
    layer0_outputs(4592) <= a xor b;
    layer0_outputs(4593) <= a xor b;
    layer0_outputs(4594) <= b and not a;
    layer0_outputs(4595) <= a and b;
    layer0_outputs(4596) <= a xor b;
    layer0_outputs(4597) <= not (a xor b);
    layer0_outputs(4598) <= not (a or b);
    layer0_outputs(4599) <= not b;
    layer0_outputs(4600) <= a or b;
    layer0_outputs(4601) <= b;
    layer0_outputs(4602) <= not (a or b);
    layer0_outputs(4603) <= a and b;
    layer0_outputs(4604) <= a and b;
    layer0_outputs(4605) <= b;
    layer0_outputs(4606) <= a or b;
    layer0_outputs(4607) <= a or b;
    layer0_outputs(4608) <= a and not b;
    layer0_outputs(4609) <= not a or b;
    layer0_outputs(4610) <= a;
    layer0_outputs(4611) <= a or b;
    layer0_outputs(4612) <= a xor b;
    layer0_outputs(4613) <= a or b;
    layer0_outputs(4614) <= not (a or b);
    layer0_outputs(4615) <= not (a xor b);
    layer0_outputs(4616) <= not b or a;
    layer0_outputs(4617) <= a and b;
    layer0_outputs(4618) <= a and not b;
    layer0_outputs(4619) <= a;
    layer0_outputs(4620) <= not b or a;
    layer0_outputs(4621) <= b;
    layer0_outputs(4622) <= not a;
    layer0_outputs(4623) <= a;
    layer0_outputs(4624) <= not (a xor b);
    layer0_outputs(4625) <= b and not a;
    layer0_outputs(4626) <= not (a xor b);
    layer0_outputs(4627) <= not (a or b);
    layer0_outputs(4628) <= not b or a;
    layer0_outputs(4629) <= not b or a;
    layer0_outputs(4630) <= not (a xor b);
    layer0_outputs(4631) <= a xor b;
    layer0_outputs(4632) <= b and not a;
    layer0_outputs(4633) <= not (a or b);
    layer0_outputs(4634) <= not (a and b);
    layer0_outputs(4635) <= not a;
    layer0_outputs(4636) <= not (a xor b);
    layer0_outputs(4637) <= not (a xor b);
    layer0_outputs(4638) <= not a;
    layer0_outputs(4639) <= 1'b0;
    layer0_outputs(4640) <= not (a or b);
    layer0_outputs(4641) <= not (a and b);
    layer0_outputs(4642) <= not (a xor b);
    layer0_outputs(4643) <= not b or a;
    layer0_outputs(4644) <= a and b;
    layer0_outputs(4645) <= not (a or b);
    layer0_outputs(4646) <= not a;
    layer0_outputs(4647) <= not (a or b);
    layer0_outputs(4648) <= a xor b;
    layer0_outputs(4649) <= b;
    layer0_outputs(4650) <= not (a xor b);
    layer0_outputs(4651) <= not (a or b);
    layer0_outputs(4652) <= b;
    layer0_outputs(4653) <= b and not a;
    layer0_outputs(4654) <= a or b;
    layer0_outputs(4655) <= a or b;
    layer0_outputs(4656) <= not (a xor b);
    layer0_outputs(4657) <= b;
    layer0_outputs(4658) <= not a or b;
    layer0_outputs(4659) <= 1'b1;
    layer0_outputs(4660) <= not (a or b);
    layer0_outputs(4661) <= not b or a;
    layer0_outputs(4662) <= not (a or b);
    layer0_outputs(4663) <= not (a or b);
    layer0_outputs(4664) <= not b;
    layer0_outputs(4665) <= not b or a;
    layer0_outputs(4666) <= not b;
    layer0_outputs(4667) <= a or b;
    layer0_outputs(4668) <= not b;
    layer0_outputs(4669) <= 1'b1;
    layer0_outputs(4670) <= a and b;
    layer0_outputs(4671) <= 1'b0;
    layer0_outputs(4672) <= not (a or b);
    layer0_outputs(4673) <= a or b;
    layer0_outputs(4674) <= not b;
    layer0_outputs(4675) <= not (a or b);
    layer0_outputs(4676) <= a;
    layer0_outputs(4677) <= a or b;
    layer0_outputs(4678) <= not b;
    layer0_outputs(4679) <= b;
    layer0_outputs(4680) <= not (a xor b);
    layer0_outputs(4681) <= not (a or b);
    layer0_outputs(4682) <= not a;
    layer0_outputs(4683) <= not b;
    layer0_outputs(4684) <= a xor b;
    layer0_outputs(4685) <= a and not b;
    layer0_outputs(4686) <= not b;
    layer0_outputs(4687) <= a and not b;
    layer0_outputs(4688) <= not (a or b);
    layer0_outputs(4689) <= not a or b;
    layer0_outputs(4690) <= not a;
    layer0_outputs(4691) <= a;
    layer0_outputs(4692) <= not b or a;
    layer0_outputs(4693) <= not a;
    layer0_outputs(4694) <= 1'b1;
    layer0_outputs(4695) <= not b;
    layer0_outputs(4696) <= not b;
    layer0_outputs(4697) <= not b;
    layer0_outputs(4698) <= not (a or b);
    layer0_outputs(4699) <= a xor b;
    layer0_outputs(4700) <= not a or b;
    layer0_outputs(4701) <= not (a xor b);
    layer0_outputs(4702) <= not a or b;
    layer0_outputs(4703) <= a or b;
    layer0_outputs(4704) <= a and b;
    layer0_outputs(4705) <= not (a xor b);
    layer0_outputs(4706) <= not a or b;
    layer0_outputs(4707) <= a;
    layer0_outputs(4708) <= a and b;
    layer0_outputs(4709) <= a;
    layer0_outputs(4710) <= not (a and b);
    layer0_outputs(4711) <= b and not a;
    layer0_outputs(4712) <= a xor b;
    layer0_outputs(4713) <= not (a xor b);
    layer0_outputs(4714) <= not a;
    layer0_outputs(4715) <= a xor b;
    layer0_outputs(4716) <= not b or a;
    layer0_outputs(4717) <= a and not b;
    layer0_outputs(4718) <= a xor b;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= not a or b;
    layer0_outputs(4721) <= not (a or b);
    layer0_outputs(4722) <= not (a or b);
    layer0_outputs(4723) <= b and not a;
    layer0_outputs(4724) <= b and not a;
    layer0_outputs(4725) <= a or b;
    layer0_outputs(4726) <= not (a or b);
    layer0_outputs(4727) <= not a;
    layer0_outputs(4728) <= not a or b;
    layer0_outputs(4729) <= a or b;
    layer0_outputs(4730) <= not a or b;
    layer0_outputs(4731) <= not (a or b);
    layer0_outputs(4732) <= not a or b;
    layer0_outputs(4733) <= a and b;
    layer0_outputs(4734) <= b and not a;
    layer0_outputs(4735) <= a and b;
    layer0_outputs(4736) <= not b or a;
    layer0_outputs(4737) <= a;
    layer0_outputs(4738) <= a;
    layer0_outputs(4739) <= 1'b0;
    layer0_outputs(4740) <= a or b;
    layer0_outputs(4741) <= not b or a;
    layer0_outputs(4742) <= not a;
    layer0_outputs(4743) <= a and not b;
    layer0_outputs(4744) <= not a;
    layer0_outputs(4745) <= not b or a;
    layer0_outputs(4746) <= not b;
    layer0_outputs(4747) <= not (a xor b);
    layer0_outputs(4748) <= 1'b0;
    layer0_outputs(4749) <= not a;
    layer0_outputs(4750) <= a;
    layer0_outputs(4751) <= b;
    layer0_outputs(4752) <= b and not a;
    layer0_outputs(4753) <= a xor b;
    layer0_outputs(4754) <= not b;
    layer0_outputs(4755) <= not b or a;
    layer0_outputs(4756) <= not b;
    layer0_outputs(4757) <= a xor b;
    layer0_outputs(4758) <= not b;
    layer0_outputs(4759) <= a or b;
    layer0_outputs(4760) <= not a;
    layer0_outputs(4761) <= not (a or b);
    layer0_outputs(4762) <= b;
    layer0_outputs(4763) <= b and not a;
    layer0_outputs(4764) <= a or b;
    layer0_outputs(4765) <= not (a xor b);
    layer0_outputs(4766) <= b;
    layer0_outputs(4767) <= not b;
    layer0_outputs(4768) <= a and not b;
    layer0_outputs(4769) <= a or b;
    layer0_outputs(4770) <= not (a or b);
    layer0_outputs(4771) <= not b or a;
    layer0_outputs(4772) <= not (a and b);
    layer0_outputs(4773) <= a;
    layer0_outputs(4774) <= b;
    layer0_outputs(4775) <= not b or a;
    layer0_outputs(4776) <= not a;
    layer0_outputs(4777) <= a and not b;
    layer0_outputs(4778) <= b;
    layer0_outputs(4779) <= not (a xor b);
    layer0_outputs(4780) <= a or b;
    layer0_outputs(4781) <= not b or a;
    layer0_outputs(4782) <= b;
    layer0_outputs(4783) <= not (a xor b);
    layer0_outputs(4784) <= a or b;
    layer0_outputs(4785) <= not a or b;
    layer0_outputs(4786) <= not (a or b);
    layer0_outputs(4787) <= not a;
    layer0_outputs(4788) <= not b or a;
    layer0_outputs(4789) <= not b;
    layer0_outputs(4790) <= not (a or b);
    layer0_outputs(4791) <= not (a and b);
    layer0_outputs(4792) <= not (a xor b);
    layer0_outputs(4793) <= a or b;
    layer0_outputs(4794) <= b;
    layer0_outputs(4795) <= not (a or b);
    layer0_outputs(4796) <= a and b;
    layer0_outputs(4797) <= b;
    layer0_outputs(4798) <= not b or a;
    layer0_outputs(4799) <= a;
    layer0_outputs(4800) <= not b;
    layer0_outputs(4801) <= not b;
    layer0_outputs(4802) <= not (a xor b);
    layer0_outputs(4803) <= not (a xor b);
    layer0_outputs(4804) <= a;
    layer0_outputs(4805) <= a or b;
    layer0_outputs(4806) <= a or b;
    layer0_outputs(4807) <= not (a xor b);
    layer0_outputs(4808) <= not a or b;
    layer0_outputs(4809) <= not (a or b);
    layer0_outputs(4810) <= 1'b0;
    layer0_outputs(4811) <= a or b;
    layer0_outputs(4812) <= not (a xor b);
    layer0_outputs(4813) <= a or b;
    layer0_outputs(4814) <= 1'b0;
    layer0_outputs(4815) <= a and not b;
    layer0_outputs(4816) <= a xor b;
    layer0_outputs(4817) <= not a;
    layer0_outputs(4818) <= a xor b;
    layer0_outputs(4819) <= a or b;
    layer0_outputs(4820) <= a or b;
    layer0_outputs(4821) <= a and not b;
    layer0_outputs(4822) <= a xor b;
    layer0_outputs(4823) <= not a;
    layer0_outputs(4824) <= not a or b;
    layer0_outputs(4825) <= not a;
    layer0_outputs(4826) <= not a or b;
    layer0_outputs(4827) <= not (a or b);
    layer0_outputs(4828) <= not (a xor b);
    layer0_outputs(4829) <= a and not b;
    layer0_outputs(4830) <= a and not b;
    layer0_outputs(4831) <= not a;
    layer0_outputs(4832) <= a and not b;
    layer0_outputs(4833) <= 1'b1;
    layer0_outputs(4834) <= a xor b;
    layer0_outputs(4835) <= a and not b;
    layer0_outputs(4836) <= a or b;
    layer0_outputs(4837) <= not (a xor b);
    layer0_outputs(4838) <= a or b;
    layer0_outputs(4839) <= a;
    layer0_outputs(4840) <= not b;
    layer0_outputs(4841) <= not (a xor b);
    layer0_outputs(4842) <= b;
    layer0_outputs(4843) <= not (a or b);
    layer0_outputs(4844) <= a xor b;
    layer0_outputs(4845) <= not (a xor b);
    layer0_outputs(4846) <= not (a xor b);
    layer0_outputs(4847) <= b;
    layer0_outputs(4848) <= not b or a;
    layer0_outputs(4849) <= not b or a;
    layer0_outputs(4850) <= not (a or b);
    layer0_outputs(4851) <= b and not a;
    layer0_outputs(4852) <= not (a xor b);
    layer0_outputs(4853) <= a;
    layer0_outputs(4854) <= a and not b;
    layer0_outputs(4855) <= not (a xor b);
    layer0_outputs(4856) <= not b;
    layer0_outputs(4857) <= not (a or b);
    layer0_outputs(4858) <= a xor b;
    layer0_outputs(4859) <= a;
    layer0_outputs(4860) <= not a or b;
    layer0_outputs(4861) <= a and not b;
    layer0_outputs(4862) <= b and not a;
    layer0_outputs(4863) <= a or b;
    layer0_outputs(4864) <= a;
    layer0_outputs(4865) <= a or b;
    layer0_outputs(4866) <= a xor b;
    layer0_outputs(4867) <= a xor b;
    layer0_outputs(4868) <= not b or a;
    layer0_outputs(4869) <= not (a or b);
    layer0_outputs(4870) <= not (a xor b);
    layer0_outputs(4871) <= b and not a;
    layer0_outputs(4872) <= not b or a;
    layer0_outputs(4873) <= not (a or b);
    layer0_outputs(4874) <= not a;
    layer0_outputs(4875) <= a or b;
    layer0_outputs(4876) <= not (a or b);
    layer0_outputs(4877) <= not b or a;
    layer0_outputs(4878) <= not a;
    layer0_outputs(4879) <= b;
    layer0_outputs(4880) <= not (a or b);
    layer0_outputs(4881) <= a;
    layer0_outputs(4882) <= b;
    layer0_outputs(4883) <= b and not a;
    layer0_outputs(4884) <= not b;
    layer0_outputs(4885) <= not (a xor b);
    layer0_outputs(4886) <= b;
    layer0_outputs(4887) <= not b;
    layer0_outputs(4888) <= a or b;
    layer0_outputs(4889) <= b and not a;
    layer0_outputs(4890) <= a or b;
    layer0_outputs(4891) <= not b or a;
    layer0_outputs(4892) <= not a or b;
    layer0_outputs(4893) <= a and b;
    layer0_outputs(4894) <= not (a and b);
    layer0_outputs(4895) <= b;
    layer0_outputs(4896) <= a xor b;
    layer0_outputs(4897) <= a;
    layer0_outputs(4898) <= not b;
    layer0_outputs(4899) <= not b;
    layer0_outputs(4900) <= a or b;
    layer0_outputs(4901) <= b and not a;
    layer0_outputs(4902) <= not a;
    layer0_outputs(4903) <= a and b;
    layer0_outputs(4904) <= not b;
    layer0_outputs(4905) <= a xor b;
    layer0_outputs(4906) <= b;
    layer0_outputs(4907) <= not (a or b);
    layer0_outputs(4908) <= b and not a;
    layer0_outputs(4909) <= a or b;
    layer0_outputs(4910) <= not (a or b);
    layer0_outputs(4911) <= a or b;
    layer0_outputs(4912) <= not a;
    layer0_outputs(4913) <= not b;
    layer0_outputs(4914) <= not b;
    layer0_outputs(4915) <= a;
    layer0_outputs(4916) <= not (a xor b);
    layer0_outputs(4917) <= a or b;
    layer0_outputs(4918) <= not a or b;
    layer0_outputs(4919) <= a or b;
    layer0_outputs(4920) <= not a or b;
    layer0_outputs(4921) <= not a;
    layer0_outputs(4922) <= a or b;
    layer0_outputs(4923) <= not (a or b);
    layer0_outputs(4924) <= not b or a;
    layer0_outputs(4925) <= not b or a;
    layer0_outputs(4926) <= a;
    layer0_outputs(4927) <= 1'b1;
    layer0_outputs(4928) <= a or b;
    layer0_outputs(4929) <= a or b;
    layer0_outputs(4930) <= not (a or b);
    layer0_outputs(4931) <= not a;
    layer0_outputs(4932) <= b and not a;
    layer0_outputs(4933) <= not (a or b);
    layer0_outputs(4934) <= not a;
    layer0_outputs(4935) <= not a;
    layer0_outputs(4936) <= not (a xor b);
    layer0_outputs(4937) <= a;
    layer0_outputs(4938) <= not (a xor b);
    layer0_outputs(4939) <= b and not a;
    layer0_outputs(4940) <= b and not a;
    layer0_outputs(4941) <= a or b;
    layer0_outputs(4942) <= a or b;
    layer0_outputs(4943) <= a xor b;
    layer0_outputs(4944) <= a or b;
    layer0_outputs(4945) <= not (a xor b);
    layer0_outputs(4946) <= not (a or b);
    layer0_outputs(4947) <= a or b;
    layer0_outputs(4948) <= b;
    layer0_outputs(4949) <= not (a or b);
    layer0_outputs(4950) <= a or b;
    layer0_outputs(4951) <= a and not b;
    layer0_outputs(4952) <= not (a or b);
    layer0_outputs(4953) <= a xor b;
    layer0_outputs(4954) <= not a or b;
    layer0_outputs(4955) <= b and not a;
    layer0_outputs(4956) <= not a or b;
    layer0_outputs(4957) <= not a or b;
    layer0_outputs(4958) <= not a;
    layer0_outputs(4959) <= 1'b1;
    layer0_outputs(4960) <= a and not b;
    layer0_outputs(4961) <= a;
    layer0_outputs(4962) <= a xor b;
    layer0_outputs(4963) <= 1'b0;
    layer0_outputs(4964) <= b;
    layer0_outputs(4965) <= a xor b;
    layer0_outputs(4966) <= not b or a;
    layer0_outputs(4967) <= not a or b;
    layer0_outputs(4968) <= not (a xor b);
    layer0_outputs(4969) <= not b;
    layer0_outputs(4970) <= a;
    layer0_outputs(4971) <= a or b;
    layer0_outputs(4972) <= not b;
    layer0_outputs(4973) <= b;
    layer0_outputs(4974) <= b;
    layer0_outputs(4975) <= a;
    layer0_outputs(4976) <= a;
    layer0_outputs(4977) <= b and not a;
    layer0_outputs(4978) <= not (a xor b);
    layer0_outputs(4979) <= a;
    layer0_outputs(4980) <= not b or a;
    layer0_outputs(4981) <= b and not a;
    layer0_outputs(4982) <= not (a or b);
    layer0_outputs(4983) <= a xor b;
    layer0_outputs(4984) <= not a or b;
    layer0_outputs(4985) <= not (a or b);
    layer0_outputs(4986) <= a or b;
    layer0_outputs(4987) <= a;
    layer0_outputs(4988) <= a and b;
    layer0_outputs(4989) <= b and not a;
    layer0_outputs(4990) <= a;
    layer0_outputs(4991) <= not b or a;
    layer0_outputs(4992) <= b;
    layer0_outputs(4993) <= 1'b1;
    layer0_outputs(4994) <= not b or a;
    layer0_outputs(4995) <= a xor b;
    layer0_outputs(4996) <= b;
    layer0_outputs(4997) <= a and not b;
    layer0_outputs(4998) <= b and not a;
    layer0_outputs(4999) <= not b or a;
    layer0_outputs(5000) <= not (a or b);
    layer0_outputs(5001) <= not b;
    layer0_outputs(5002) <= not (a xor b);
    layer0_outputs(5003) <= a or b;
    layer0_outputs(5004) <= a xor b;
    layer0_outputs(5005) <= b and not a;
    layer0_outputs(5006) <= not b;
    layer0_outputs(5007) <= a and b;
    layer0_outputs(5008) <= not (a or b);
    layer0_outputs(5009) <= b;
    layer0_outputs(5010) <= not (a or b);
    layer0_outputs(5011) <= b;
    layer0_outputs(5012) <= a xor b;
    layer0_outputs(5013) <= a or b;
    layer0_outputs(5014) <= not (a or b);
    layer0_outputs(5015) <= a and not b;
    layer0_outputs(5016) <= not a or b;
    layer0_outputs(5017) <= a xor b;
    layer0_outputs(5018) <= a and b;
    layer0_outputs(5019) <= a and b;
    layer0_outputs(5020) <= a xor b;
    layer0_outputs(5021) <= not a;
    layer0_outputs(5022) <= not (a or b);
    layer0_outputs(5023) <= b;
    layer0_outputs(5024) <= not (a xor b);
    layer0_outputs(5025) <= b;
    layer0_outputs(5026) <= not (a xor b);
    layer0_outputs(5027) <= a;
    layer0_outputs(5028) <= a or b;
    layer0_outputs(5029) <= b and not a;
    layer0_outputs(5030) <= not b;
    layer0_outputs(5031) <= not (a xor b);
    layer0_outputs(5032) <= not a or b;
    layer0_outputs(5033) <= not a;
    layer0_outputs(5034) <= not a or b;
    layer0_outputs(5035) <= b;
    layer0_outputs(5036) <= not a;
    layer0_outputs(5037) <= a or b;
    layer0_outputs(5038) <= a and not b;
    layer0_outputs(5039) <= not (a xor b);
    layer0_outputs(5040) <= not b or a;
    layer0_outputs(5041) <= a xor b;
    layer0_outputs(5042) <= b;
    layer0_outputs(5043) <= not a or b;
    layer0_outputs(5044) <= not b;
    layer0_outputs(5045) <= a xor b;
    layer0_outputs(5046) <= not (a xor b);
    layer0_outputs(5047) <= not (a xor b);
    layer0_outputs(5048) <= not a or b;
    layer0_outputs(5049) <= not (a xor b);
    layer0_outputs(5050) <= b;
    layer0_outputs(5051) <= a and not b;
    layer0_outputs(5052) <= not b;
    layer0_outputs(5053) <= not (a xor b);
    layer0_outputs(5054) <= not (a or b);
    layer0_outputs(5055) <= not a or b;
    layer0_outputs(5056) <= not a;
    layer0_outputs(5057) <= not a;
    layer0_outputs(5058) <= 1'b1;
    layer0_outputs(5059) <= 1'b0;
    layer0_outputs(5060) <= not (a xor b);
    layer0_outputs(5061) <= 1'b1;
    layer0_outputs(5062) <= a xor b;
    layer0_outputs(5063) <= not (a xor b);
    layer0_outputs(5064) <= not a;
    layer0_outputs(5065) <= a or b;
    layer0_outputs(5066) <= b and not a;
    layer0_outputs(5067) <= b and not a;
    layer0_outputs(5068) <= 1'b1;
    layer0_outputs(5069) <= not (a and b);
    layer0_outputs(5070) <= not a or b;
    layer0_outputs(5071) <= b;
    layer0_outputs(5072) <= not a or b;
    layer0_outputs(5073) <= a;
    layer0_outputs(5074) <= not (a or b);
    layer0_outputs(5075) <= a or b;
    layer0_outputs(5076) <= a xor b;
    layer0_outputs(5077) <= not (a or b);
    layer0_outputs(5078) <= b and not a;
    layer0_outputs(5079) <= not a;
    layer0_outputs(5080) <= not b;
    layer0_outputs(5081) <= not (a or b);
    layer0_outputs(5082) <= b and not a;
    layer0_outputs(5083) <= a and not b;
    layer0_outputs(5084) <= a or b;
    layer0_outputs(5085) <= not a;
    layer0_outputs(5086) <= b and not a;
    layer0_outputs(5087) <= not a or b;
    layer0_outputs(5088) <= not (a or b);
    layer0_outputs(5089) <= not (a xor b);
    layer0_outputs(5090) <= a or b;
    layer0_outputs(5091) <= not a;
    layer0_outputs(5092) <= a;
    layer0_outputs(5093) <= b;
    layer0_outputs(5094) <= a and not b;
    layer0_outputs(5095) <= not a or b;
    layer0_outputs(5096) <= not b;
    layer0_outputs(5097) <= not b or a;
    layer0_outputs(5098) <= not b;
    layer0_outputs(5099) <= not (a xor b);
    layer0_outputs(5100) <= not (a and b);
    layer0_outputs(5101) <= a xor b;
    layer0_outputs(5102) <= not a or b;
    layer0_outputs(5103) <= not (a xor b);
    layer0_outputs(5104) <= not b;
    layer0_outputs(5105) <= not (a or b);
    layer0_outputs(5106) <= b and not a;
    layer0_outputs(5107) <= b and not a;
    layer0_outputs(5108) <= a;
    layer0_outputs(5109) <= not b;
    layer0_outputs(5110) <= a xor b;
    layer0_outputs(5111) <= not (a and b);
    layer0_outputs(5112) <= a xor b;
    layer0_outputs(5113) <= b and not a;
    layer0_outputs(5114) <= not a;
    layer0_outputs(5115) <= 1'b1;
    layer0_outputs(5116) <= b and not a;
    layer0_outputs(5117) <= not a;
    layer0_outputs(5118) <= not (a or b);
    layer0_outputs(5119) <= a or b;
    layer0_outputs(5120) <= not (a or b);
    layer0_outputs(5121) <= not b;
    layer0_outputs(5122) <= a and b;
    layer0_outputs(5123) <= b;
    layer0_outputs(5124) <= a xor b;
    layer0_outputs(5125) <= a or b;
    layer0_outputs(5126) <= not (a or b);
    layer0_outputs(5127) <= a;
    layer0_outputs(5128) <= not a or b;
    layer0_outputs(5129) <= not a or b;
    layer0_outputs(5130) <= not b;
    layer0_outputs(5131) <= b and not a;
    layer0_outputs(5132) <= a;
    layer0_outputs(5133) <= not b;
    layer0_outputs(5134) <= not b;
    layer0_outputs(5135) <= a xor b;
    layer0_outputs(5136) <= not (a xor b);
    layer0_outputs(5137) <= not (a and b);
    layer0_outputs(5138) <= b;
    layer0_outputs(5139) <= a and not b;
    layer0_outputs(5140) <= not (a or b);
    layer0_outputs(5141) <= b;
    layer0_outputs(5142) <= a xor b;
    layer0_outputs(5143) <= b;
    layer0_outputs(5144) <= not (a xor b);
    layer0_outputs(5145) <= not a or b;
    layer0_outputs(5146) <= a or b;
    layer0_outputs(5147) <= not b or a;
    layer0_outputs(5148) <= not a;
    layer0_outputs(5149) <= not (a xor b);
    layer0_outputs(5150) <= a and not b;
    layer0_outputs(5151) <= not (a and b);
    layer0_outputs(5152) <= a or b;
    layer0_outputs(5153) <= not b or a;
    layer0_outputs(5154) <= a or b;
    layer0_outputs(5155) <= a or b;
    layer0_outputs(5156) <= not b;
    layer0_outputs(5157) <= a or b;
    layer0_outputs(5158) <= a or b;
    layer0_outputs(5159) <= a and b;
    layer0_outputs(5160) <= not (a xor b);
    layer0_outputs(5161) <= not a or b;
    layer0_outputs(5162) <= not (a or b);
    layer0_outputs(5163) <= not (a xor b);
    layer0_outputs(5164) <= not b;
    layer0_outputs(5165) <= a or b;
    layer0_outputs(5166) <= a or b;
    layer0_outputs(5167) <= not b;
    layer0_outputs(5168) <= not b;
    layer0_outputs(5169) <= a xor b;
    layer0_outputs(5170) <= not b;
    layer0_outputs(5171) <= not (a or b);
    layer0_outputs(5172) <= a and not b;
    layer0_outputs(5173) <= not b or a;
    layer0_outputs(5174) <= a or b;
    layer0_outputs(5175) <= not b;
    layer0_outputs(5176) <= a xor b;
    layer0_outputs(5177) <= not (a xor b);
    layer0_outputs(5178) <= a;
    layer0_outputs(5179) <= b;
    layer0_outputs(5180) <= b;
    layer0_outputs(5181) <= not (a xor b);
    layer0_outputs(5182) <= not b or a;
    layer0_outputs(5183) <= not a;
    layer0_outputs(5184) <= a and not b;
    layer0_outputs(5185) <= a and not b;
    layer0_outputs(5186) <= a and not b;
    layer0_outputs(5187) <= not a;
    layer0_outputs(5188) <= b;
    layer0_outputs(5189) <= a and b;
    layer0_outputs(5190) <= not (a or b);
    layer0_outputs(5191) <= not b or a;
    layer0_outputs(5192) <= not (a xor b);
    layer0_outputs(5193) <= not (a or b);
    layer0_outputs(5194) <= a or b;
    layer0_outputs(5195) <= b and not a;
    layer0_outputs(5196) <= not b or a;
    layer0_outputs(5197) <= a or b;
    layer0_outputs(5198) <= a or b;
    layer0_outputs(5199) <= not (a xor b);
    layer0_outputs(5200) <= not a or b;
    layer0_outputs(5201) <= not a or b;
    layer0_outputs(5202) <= not a;
    layer0_outputs(5203) <= b;
    layer0_outputs(5204) <= a;
    layer0_outputs(5205) <= a and not b;
    layer0_outputs(5206) <= a or b;
    layer0_outputs(5207) <= not (a and b);
    layer0_outputs(5208) <= b;
    layer0_outputs(5209) <= not b or a;
    layer0_outputs(5210) <= a;
    layer0_outputs(5211) <= not a or b;
    layer0_outputs(5212) <= not (a xor b);
    layer0_outputs(5213) <= not b or a;
    layer0_outputs(5214) <= not (a or b);
    layer0_outputs(5215) <= not b or a;
    layer0_outputs(5216) <= not (a or b);
    layer0_outputs(5217) <= not a or b;
    layer0_outputs(5218) <= not (a xor b);
    layer0_outputs(5219) <= b and not a;
    layer0_outputs(5220) <= not (a or b);
    layer0_outputs(5221) <= not a or b;
    layer0_outputs(5222) <= b;
    layer0_outputs(5223) <= 1'b0;
    layer0_outputs(5224) <= a xor b;
    layer0_outputs(5225) <= not a or b;
    layer0_outputs(5226) <= a and b;
    layer0_outputs(5227) <= a and b;
    layer0_outputs(5228) <= not (a xor b);
    layer0_outputs(5229) <= not (a or b);
    layer0_outputs(5230) <= not b or a;
    layer0_outputs(5231) <= a;
    layer0_outputs(5232) <= a;
    layer0_outputs(5233) <= not (a xor b);
    layer0_outputs(5234) <= not b or a;
    layer0_outputs(5235) <= a or b;
    layer0_outputs(5236) <= b and not a;
    layer0_outputs(5237) <= a;
    layer0_outputs(5238) <= not a;
    layer0_outputs(5239) <= a xor b;
    layer0_outputs(5240) <= a and not b;
    layer0_outputs(5241) <= not a;
    layer0_outputs(5242) <= not a;
    layer0_outputs(5243) <= not b or a;
    layer0_outputs(5244) <= not (a xor b);
    layer0_outputs(5245) <= not (a or b);
    layer0_outputs(5246) <= not a or b;
    layer0_outputs(5247) <= not (a and b);
    layer0_outputs(5248) <= not a;
    layer0_outputs(5249) <= b and not a;
    layer0_outputs(5250) <= not (a xor b);
    layer0_outputs(5251) <= a xor b;
    layer0_outputs(5252) <= not (a xor b);
    layer0_outputs(5253) <= a or b;
    layer0_outputs(5254) <= not b or a;
    layer0_outputs(5255) <= a and not b;
    layer0_outputs(5256) <= b and not a;
    layer0_outputs(5257) <= b and not a;
    layer0_outputs(5258) <= b and not a;
    layer0_outputs(5259) <= not a or b;
    layer0_outputs(5260) <= a and not b;
    layer0_outputs(5261) <= not a or b;
    layer0_outputs(5262) <= not (a xor b);
    layer0_outputs(5263) <= not (a xor b);
    layer0_outputs(5264) <= a;
    layer0_outputs(5265) <= not b;
    layer0_outputs(5266) <= a and not b;
    layer0_outputs(5267) <= a xor b;
    layer0_outputs(5268) <= not a or b;
    layer0_outputs(5269) <= not a or b;
    layer0_outputs(5270) <= a or b;
    layer0_outputs(5271) <= a and not b;
    layer0_outputs(5272) <= a or b;
    layer0_outputs(5273) <= a and not b;
    layer0_outputs(5274) <= not a or b;
    layer0_outputs(5275) <= not (a or b);
    layer0_outputs(5276) <= not (a xor b);
    layer0_outputs(5277) <= b;
    layer0_outputs(5278) <= a or b;
    layer0_outputs(5279) <= b;
    layer0_outputs(5280) <= a and b;
    layer0_outputs(5281) <= b and not a;
    layer0_outputs(5282) <= not a;
    layer0_outputs(5283) <= a xor b;
    layer0_outputs(5284) <= b;
    layer0_outputs(5285) <= a or b;
    layer0_outputs(5286) <= not (a or b);
    layer0_outputs(5287) <= a xor b;
    layer0_outputs(5288) <= a and b;
    layer0_outputs(5289) <= not b;
    layer0_outputs(5290) <= not a;
    layer0_outputs(5291) <= a;
    layer0_outputs(5292) <= not a;
    layer0_outputs(5293) <= a;
    layer0_outputs(5294) <= 1'b1;
    layer0_outputs(5295) <= a and b;
    layer0_outputs(5296) <= not (a or b);
    layer0_outputs(5297) <= a and not b;
    layer0_outputs(5298) <= b and not a;
    layer0_outputs(5299) <= b;
    layer0_outputs(5300) <= not (a or b);
    layer0_outputs(5301) <= b;
    layer0_outputs(5302) <= a;
    layer0_outputs(5303) <= a or b;
    layer0_outputs(5304) <= not b or a;
    layer0_outputs(5305) <= a and not b;
    layer0_outputs(5306) <= a xor b;
    layer0_outputs(5307) <= not b or a;
    layer0_outputs(5308) <= a and not b;
    layer0_outputs(5309) <= not (a xor b);
    layer0_outputs(5310) <= not b or a;
    layer0_outputs(5311) <= not (a or b);
    layer0_outputs(5312) <= b;
    layer0_outputs(5313) <= a or b;
    layer0_outputs(5314) <= b and not a;
    layer0_outputs(5315) <= b;
    layer0_outputs(5316) <= not a or b;
    layer0_outputs(5317) <= not a or b;
    layer0_outputs(5318) <= not b;
    layer0_outputs(5319) <= a and b;
    layer0_outputs(5320) <= a;
    layer0_outputs(5321) <= not (a xor b);
    layer0_outputs(5322) <= 1'b1;
    layer0_outputs(5323) <= a or b;
    layer0_outputs(5324) <= a or b;
    layer0_outputs(5325) <= not a or b;
    layer0_outputs(5326) <= not b;
    layer0_outputs(5327) <= not (a or b);
    layer0_outputs(5328) <= not a;
    layer0_outputs(5329) <= not a or b;
    layer0_outputs(5330) <= a or b;
    layer0_outputs(5331) <= a and not b;
    layer0_outputs(5332) <= not (a or b);
    layer0_outputs(5333) <= not (a or b);
    layer0_outputs(5334) <= not b or a;
    layer0_outputs(5335) <= not a or b;
    layer0_outputs(5336) <= a and b;
    layer0_outputs(5337) <= 1'b0;
    layer0_outputs(5338) <= a;
    layer0_outputs(5339) <= a or b;
    layer0_outputs(5340) <= a;
    layer0_outputs(5341) <= b;
    layer0_outputs(5342) <= a xor b;
    layer0_outputs(5343) <= a;
    layer0_outputs(5344) <= a and b;
    layer0_outputs(5345) <= a;
    layer0_outputs(5346) <= a;
    layer0_outputs(5347) <= a or b;
    layer0_outputs(5348) <= not (a xor b);
    layer0_outputs(5349) <= a;
    layer0_outputs(5350) <= b and not a;
    layer0_outputs(5351) <= not (a xor b);
    layer0_outputs(5352) <= 1'b0;
    layer0_outputs(5353) <= a or b;
    layer0_outputs(5354) <= not (a or b);
    layer0_outputs(5355) <= not b or a;
    layer0_outputs(5356) <= a or b;
    layer0_outputs(5357) <= a or b;
    layer0_outputs(5358) <= a and b;
    layer0_outputs(5359) <= 1'b0;
    layer0_outputs(5360) <= not a;
    layer0_outputs(5361) <= not b or a;
    layer0_outputs(5362) <= b;
    layer0_outputs(5363) <= b and not a;
    layer0_outputs(5364) <= a;
    layer0_outputs(5365) <= 1'b1;
    layer0_outputs(5366) <= a;
    layer0_outputs(5367) <= not (a and b);
    layer0_outputs(5368) <= not (a xor b);
    layer0_outputs(5369) <= not (a xor b);
    layer0_outputs(5370) <= a;
    layer0_outputs(5371) <= b and not a;
    layer0_outputs(5372) <= not b;
    layer0_outputs(5373) <= a and not b;
    layer0_outputs(5374) <= not a;
    layer0_outputs(5375) <= not b or a;
    layer0_outputs(5376) <= not a or b;
    layer0_outputs(5377) <= not a;
    layer0_outputs(5378) <= a xor b;
    layer0_outputs(5379) <= not (a or b);
    layer0_outputs(5380) <= not b or a;
    layer0_outputs(5381) <= not a;
    layer0_outputs(5382) <= not a or b;
    layer0_outputs(5383) <= a or b;
    layer0_outputs(5384) <= b;
    layer0_outputs(5385) <= a;
    layer0_outputs(5386) <= a and not b;
    layer0_outputs(5387) <= a xor b;
    layer0_outputs(5388) <= not b or a;
    layer0_outputs(5389) <= not (a or b);
    layer0_outputs(5390) <= not (a xor b);
    layer0_outputs(5391) <= 1'b0;
    layer0_outputs(5392) <= a and b;
    layer0_outputs(5393) <= a or b;
    layer0_outputs(5394) <= not (a xor b);
    layer0_outputs(5395) <= a and not b;
    layer0_outputs(5396) <= not (a xor b);
    layer0_outputs(5397) <= a xor b;
    layer0_outputs(5398) <= b and not a;
    layer0_outputs(5399) <= not (a or b);
    layer0_outputs(5400) <= a xor b;
    layer0_outputs(5401) <= 1'b1;
    layer0_outputs(5402) <= not (a or b);
    layer0_outputs(5403) <= a xor b;
    layer0_outputs(5404) <= b;
    layer0_outputs(5405) <= not a;
    layer0_outputs(5406) <= a xor b;
    layer0_outputs(5407) <= not b;
    layer0_outputs(5408) <= a and b;
    layer0_outputs(5409) <= not (a or b);
    layer0_outputs(5410) <= not (a xor b);
    layer0_outputs(5411) <= a xor b;
    layer0_outputs(5412) <= a;
    layer0_outputs(5413) <= not b or a;
    layer0_outputs(5414) <= b and not a;
    layer0_outputs(5415) <= not b;
    layer0_outputs(5416) <= not b or a;
    layer0_outputs(5417) <= a xor b;
    layer0_outputs(5418) <= 1'b0;
    layer0_outputs(5419) <= not a;
    layer0_outputs(5420) <= 1'b1;
    layer0_outputs(5421) <= a xor b;
    layer0_outputs(5422) <= b and not a;
    layer0_outputs(5423) <= b and not a;
    layer0_outputs(5424) <= not (a xor b);
    layer0_outputs(5425) <= not b;
    layer0_outputs(5426) <= not b;
    layer0_outputs(5427) <= a and not b;
    layer0_outputs(5428) <= a xor b;
    layer0_outputs(5429) <= 1'b0;
    layer0_outputs(5430) <= not b or a;
    layer0_outputs(5431) <= not b or a;
    layer0_outputs(5432) <= not (a xor b);
    layer0_outputs(5433) <= 1'b0;
    layer0_outputs(5434) <= not (a or b);
    layer0_outputs(5435) <= a or b;
    layer0_outputs(5436) <= b and not a;
    layer0_outputs(5437) <= not a;
    layer0_outputs(5438) <= not (a xor b);
    layer0_outputs(5439) <= not b or a;
    layer0_outputs(5440) <= not a;
    layer0_outputs(5441) <= a xor b;
    layer0_outputs(5442) <= not a or b;
    layer0_outputs(5443) <= not b;
    layer0_outputs(5444) <= not b or a;
    layer0_outputs(5445) <= a or b;
    layer0_outputs(5446) <= not b or a;
    layer0_outputs(5447) <= not a or b;
    layer0_outputs(5448) <= a or b;
    layer0_outputs(5449) <= 1'b0;
    layer0_outputs(5450) <= not (a and b);
    layer0_outputs(5451) <= not (a or b);
    layer0_outputs(5452) <= a;
    layer0_outputs(5453) <= a xor b;
    layer0_outputs(5454) <= a and b;
    layer0_outputs(5455) <= b;
    layer0_outputs(5456) <= a or b;
    layer0_outputs(5457) <= 1'b1;
    layer0_outputs(5458) <= a and not b;
    layer0_outputs(5459) <= not (a or b);
    layer0_outputs(5460) <= b and not a;
    layer0_outputs(5461) <= not a or b;
    layer0_outputs(5462) <= not (a xor b);
    layer0_outputs(5463) <= a or b;
    layer0_outputs(5464) <= not (a or b);
    layer0_outputs(5465) <= a;
    layer0_outputs(5466) <= not a;
    layer0_outputs(5467) <= not a;
    layer0_outputs(5468) <= b;
    layer0_outputs(5469) <= a or b;
    layer0_outputs(5470) <= not b or a;
    layer0_outputs(5471) <= not a;
    layer0_outputs(5472) <= a;
    layer0_outputs(5473) <= not b;
    layer0_outputs(5474) <= a or b;
    layer0_outputs(5475) <= not (a and b);
    layer0_outputs(5476) <= not a;
    layer0_outputs(5477) <= not (a or b);
    layer0_outputs(5478) <= not b;
    layer0_outputs(5479) <= a or b;
    layer0_outputs(5480) <= a;
    layer0_outputs(5481) <= 1'b1;
    layer0_outputs(5482) <= b;
    layer0_outputs(5483) <= 1'b1;
    layer0_outputs(5484) <= 1'b1;
    layer0_outputs(5485) <= not a or b;
    layer0_outputs(5486) <= not a;
    layer0_outputs(5487) <= not (a xor b);
    layer0_outputs(5488) <= a and not b;
    layer0_outputs(5489) <= not (a or b);
    layer0_outputs(5490) <= not a or b;
    layer0_outputs(5491) <= b and not a;
    layer0_outputs(5492) <= a;
    layer0_outputs(5493) <= not a;
    layer0_outputs(5494) <= not (a or b);
    layer0_outputs(5495) <= not b;
    layer0_outputs(5496) <= not (a xor b);
    layer0_outputs(5497) <= a or b;
    layer0_outputs(5498) <= not (a xor b);
    layer0_outputs(5499) <= not (a xor b);
    layer0_outputs(5500) <= a xor b;
    layer0_outputs(5501) <= a and b;
    layer0_outputs(5502) <= not a or b;
    layer0_outputs(5503) <= 1'b1;
    layer0_outputs(5504) <= not a;
    layer0_outputs(5505) <= not (a xor b);
    layer0_outputs(5506) <= a or b;
    layer0_outputs(5507) <= b;
    layer0_outputs(5508) <= not b or a;
    layer0_outputs(5509) <= b and not a;
    layer0_outputs(5510) <= a and not b;
    layer0_outputs(5511) <= b and not a;
    layer0_outputs(5512) <= b;
    layer0_outputs(5513) <= a;
    layer0_outputs(5514) <= not a or b;
    layer0_outputs(5515) <= b;
    layer0_outputs(5516) <= a xor b;
    layer0_outputs(5517) <= not (a or b);
    layer0_outputs(5518) <= a xor b;
    layer0_outputs(5519) <= not a;
    layer0_outputs(5520) <= a or b;
    layer0_outputs(5521) <= b;
    layer0_outputs(5522) <= not b;
    layer0_outputs(5523) <= a or b;
    layer0_outputs(5524) <= a xor b;
    layer0_outputs(5525) <= not b or a;
    layer0_outputs(5526) <= a;
    layer0_outputs(5527) <= not b or a;
    layer0_outputs(5528) <= a or b;
    layer0_outputs(5529) <= a xor b;
    layer0_outputs(5530) <= b;
    layer0_outputs(5531) <= a and b;
    layer0_outputs(5532) <= not b;
    layer0_outputs(5533) <= b and not a;
    layer0_outputs(5534) <= not (a or b);
    layer0_outputs(5535) <= b and not a;
    layer0_outputs(5536) <= not b or a;
    layer0_outputs(5537) <= not a;
    layer0_outputs(5538) <= not a or b;
    layer0_outputs(5539) <= not b;
    layer0_outputs(5540) <= 1'b0;
    layer0_outputs(5541) <= not b;
    layer0_outputs(5542) <= not a or b;
    layer0_outputs(5543) <= not (a xor b);
    layer0_outputs(5544) <= a;
    layer0_outputs(5545) <= a;
    layer0_outputs(5546) <= not b;
    layer0_outputs(5547) <= not (a or b);
    layer0_outputs(5548) <= not (a or b);
    layer0_outputs(5549) <= a and b;
    layer0_outputs(5550) <= b;
    layer0_outputs(5551) <= a or b;
    layer0_outputs(5552) <= a;
    layer0_outputs(5553) <= not a or b;
    layer0_outputs(5554) <= not a or b;
    layer0_outputs(5555) <= 1'b1;
    layer0_outputs(5556) <= not a or b;
    layer0_outputs(5557) <= a;
    layer0_outputs(5558) <= not (a xor b);
    layer0_outputs(5559) <= not (a or b);
    layer0_outputs(5560) <= a or b;
    layer0_outputs(5561) <= a xor b;
    layer0_outputs(5562) <= a or b;
    layer0_outputs(5563) <= not a or b;
    layer0_outputs(5564) <= a;
    layer0_outputs(5565) <= a and not b;
    layer0_outputs(5566) <= a and b;
    layer0_outputs(5567) <= b and not a;
    layer0_outputs(5568) <= not (a or b);
    layer0_outputs(5569) <= a or b;
    layer0_outputs(5570) <= a;
    layer0_outputs(5571) <= a;
    layer0_outputs(5572) <= a and not b;
    layer0_outputs(5573) <= not a;
    layer0_outputs(5574) <= not (a xor b);
    layer0_outputs(5575) <= not a;
    layer0_outputs(5576) <= not a;
    layer0_outputs(5577) <= not a;
    layer0_outputs(5578) <= not (a xor b);
    layer0_outputs(5579) <= not (a xor b);
    layer0_outputs(5580) <= not (a or b);
    layer0_outputs(5581) <= a xor b;
    layer0_outputs(5582) <= not b or a;
    layer0_outputs(5583) <= a xor b;
    layer0_outputs(5584) <= not a;
    layer0_outputs(5585) <= a or b;
    layer0_outputs(5586) <= not b or a;
    layer0_outputs(5587) <= not a;
    layer0_outputs(5588) <= b and not a;
    layer0_outputs(5589) <= not (a xor b);
    layer0_outputs(5590) <= b;
    layer0_outputs(5591) <= not a or b;
    layer0_outputs(5592) <= not (a or b);
    layer0_outputs(5593) <= not (a xor b);
    layer0_outputs(5594) <= a or b;
    layer0_outputs(5595) <= a;
    layer0_outputs(5596) <= b and not a;
    layer0_outputs(5597) <= a xor b;
    layer0_outputs(5598) <= a;
    layer0_outputs(5599) <= not b or a;
    layer0_outputs(5600) <= not (a xor b);
    layer0_outputs(5601) <= a or b;
    layer0_outputs(5602) <= a xor b;
    layer0_outputs(5603) <= not (a xor b);
    layer0_outputs(5604) <= not a or b;
    layer0_outputs(5605) <= a;
    layer0_outputs(5606) <= a and not b;
    layer0_outputs(5607) <= a xor b;
    layer0_outputs(5608) <= not a;
    layer0_outputs(5609) <= a;
    layer0_outputs(5610) <= 1'b1;
    layer0_outputs(5611) <= a;
    layer0_outputs(5612) <= b and not a;
    layer0_outputs(5613) <= not (a or b);
    layer0_outputs(5614) <= not (a xor b);
    layer0_outputs(5615) <= not (a and b);
    layer0_outputs(5616) <= a and not b;
    layer0_outputs(5617) <= a or b;
    layer0_outputs(5618) <= a xor b;
    layer0_outputs(5619) <= a and b;
    layer0_outputs(5620) <= b;
    layer0_outputs(5621) <= a and b;
    layer0_outputs(5622) <= a;
    layer0_outputs(5623) <= not (a or b);
    layer0_outputs(5624) <= 1'b1;
    layer0_outputs(5625) <= b and not a;
    layer0_outputs(5626) <= a or b;
    layer0_outputs(5627) <= not b;
    layer0_outputs(5628) <= a xor b;
    layer0_outputs(5629) <= a or b;
    layer0_outputs(5630) <= not (a or b);
    layer0_outputs(5631) <= a;
    layer0_outputs(5632) <= a or b;
    layer0_outputs(5633) <= a;
    layer0_outputs(5634) <= not a or b;
    layer0_outputs(5635) <= a and b;
    layer0_outputs(5636) <= a and not b;
    layer0_outputs(5637) <= 1'b0;
    layer0_outputs(5638) <= not (a xor b);
    layer0_outputs(5639) <= not (a or b);
    layer0_outputs(5640) <= not b;
    layer0_outputs(5641) <= a;
    layer0_outputs(5642) <= 1'b1;
    layer0_outputs(5643) <= not a or b;
    layer0_outputs(5644) <= a and not b;
    layer0_outputs(5645) <= a or b;
    layer0_outputs(5646) <= 1'b0;
    layer0_outputs(5647) <= not b;
    layer0_outputs(5648) <= a or b;
    layer0_outputs(5649) <= not a or b;
    layer0_outputs(5650) <= b;
    layer0_outputs(5651) <= not b;
    layer0_outputs(5652) <= not a or b;
    layer0_outputs(5653) <= not (a xor b);
    layer0_outputs(5654) <= a xor b;
    layer0_outputs(5655) <= b and not a;
    layer0_outputs(5656) <= b;
    layer0_outputs(5657) <= a xor b;
    layer0_outputs(5658) <= not a or b;
    layer0_outputs(5659) <= a;
    layer0_outputs(5660) <= a and b;
    layer0_outputs(5661) <= a xor b;
    layer0_outputs(5662) <= not (a and b);
    layer0_outputs(5663) <= not (a or b);
    layer0_outputs(5664) <= not a or b;
    layer0_outputs(5665) <= not a;
    layer0_outputs(5666) <= a or b;
    layer0_outputs(5667) <= not (a or b);
    layer0_outputs(5668) <= a;
    layer0_outputs(5669) <= not (a or b);
    layer0_outputs(5670) <= a;
    layer0_outputs(5671) <= not a;
    layer0_outputs(5672) <= not (a or b);
    layer0_outputs(5673) <= a xor b;
    layer0_outputs(5674) <= a or b;
    layer0_outputs(5675) <= b and not a;
    layer0_outputs(5676) <= not a or b;
    layer0_outputs(5677) <= not (a xor b);
    layer0_outputs(5678) <= b and not a;
    layer0_outputs(5679) <= a and not b;
    layer0_outputs(5680) <= a;
    layer0_outputs(5681) <= b and not a;
    layer0_outputs(5682) <= a xor b;
    layer0_outputs(5683) <= not a or b;
    layer0_outputs(5684) <= 1'b1;
    layer0_outputs(5685) <= not (a or b);
    layer0_outputs(5686) <= b;
    layer0_outputs(5687) <= not (a or b);
    layer0_outputs(5688) <= not (a or b);
    layer0_outputs(5689) <= not a;
    layer0_outputs(5690) <= b;
    layer0_outputs(5691) <= b;
    layer0_outputs(5692) <= not a or b;
    layer0_outputs(5693) <= not a or b;
    layer0_outputs(5694) <= not (a xor b);
    layer0_outputs(5695) <= 1'b0;
    layer0_outputs(5696) <= not b or a;
    layer0_outputs(5697) <= 1'b0;
    layer0_outputs(5698) <= not a or b;
    layer0_outputs(5699) <= a or b;
    layer0_outputs(5700) <= a or b;
    layer0_outputs(5701) <= not b or a;
    layer0_outputs(5702) <= a;
    layer0_outputs(5703) <= b;
    layer0_outputs(5704) <= a;
    layer0_outputs(5705) <= a and b;
    layer0_outputs(5706) <= not (a and b);
    layer0_outputs(5707) <= b and not a;
    layer0_outputs(5708) <= b;
    layer0_outputs(5709) <= not b;
    layer0_outputs(5710) <= not (a or b);
    layer0_outputs(5711) <= a or b;
    layer0_outputs(5712) <= b;
    layer0_outputs(5713) <= 1'b0;
    layer0_outputs(5714) <= a;
    layer0_outputs(5715) <= not (a xor b);
    layer0_outputs(5716) <= a;
    layer0_outputs(5717) <= not (a xor b);
    layer0_outputs(5718) <= not b;
    layer0_outputs(5719) <= a xor b;
    layer0_outputs(5720) <= not b or a;
    layer0_outputs(5721) <= a xor b;
    layer0_outputs(5722) <= not a or b;
    layer0_outputs(5723) <= b;
    layer0_outputs(5724) <= a or b;
    layer0_outputs(5725) <= not b;
    layer0_outputs(5726) <= not (a xor b);
    layer0_outputs(5727) <= 1'b1;
    layer0_outputs(5728) <= not (a or b);
    layer0_outputs(5729) <= a or b;
    layer0_outputs(5730) <= not a;
    layer0_outputs(5731) <= not a or b;
    layer0_outputs(5732) <= not (a or b);
    layer0_outputs(5733) <= not (a and b);
    layer0_outputs(5734) <= a xor b;
    layer0_outputs(5735) <= a;
    layer0_outputs(5736) <= b and not a;
    layer0_outputs(5737) <= not a or b;
    layer0_outputs(5738) <= b and not a;
    layer0_outputs(5739) <= not b;
    layer0_outputs(5740) <= not (a xor b);
    layer0_outputs(5741) <= not (a xor b);
    layer0_outputs(5742) <= a xor b;
    layer0_outputs(5743) <= not (a xor b);
    layer0_outputs(5744) <= not (a or b);
    layer0_outputs(5745) <= not a;
    layer0_outputs(5746) <= not a;
    layer0_outputs(5747) <= b;
    layer0_outputs(5748) <= 1'b0;
    layer0_outputs(5749) <= 1'b0;
    layer0_outputs(5750) <= a;
    layer0_outputs(5751) <= not b;
    layer0_outputs(5752) <= not (a xor b);
    layer0_outputs(5753) <= not a or b;
    layer0_outputs(5754) <= not a;
    layer0_outputs(5755) <= 1'b0;
    layer0_outputs(5756) <= a xor b;
    layer0_outputs(5757) <= not b;
    layer0_outputs(5758) <= 1'b1;
    layer0_outputs(5759) <= a;
    layer0_outputs(5760) <= a;
    layer0_outputs(5761) <= not (a xor b);
    layer0_outputs(5762) <= 1'b1;
    layer0_outputs(5763) <= not (a or b);
    layer0_outputs(5764) <= not (a or b);
    layer0_outputs(5765) <= a and not b;
    layer0_outputs(5766) <= not a;
    layer0_outputs(5767) <= b and not a;
    layer0_outputs(5768) <= not a;
    layer0_outputs(5769) <= not b;
    layer0_outputs(5770) <= b and not a;
    layer0_outputs(5771) <= b;
    layer0_outputs(5772) <= 1'b1;
    layer0_outputs(5773) <= a or b;
    layer0_outputs(5774) <= not (a or b);
    layer0_outputs(5775) <= not (a xor b);
    layer0_outputs(5776) <= b;
    layer0_outputs(5777) <= b;
    layer0_outputs(5778) <= not b or a;
    layer0_outputs(5779) <= not (a xor b);
    layer0_outputs(5780) <= not (a xor b);
    layer0_outputs(5781) <= not (a xor b);
    layer0_outputs(5782) <= b and not a;
    layer0_outputs(5783) <= a or b;
    layer0_outputs(5784) <= a;
    layer0_outputs(5785) <= a;
    layer0_outputs(5786) <= 1'b0;
    layer0_outputs(5787) <= not b;
    layer0_outputs(5788) <= b;
    layer0_outputs(5789) <= a xor b;
    layer0_outputs(5790) <= a and b;
    layer0_outputs(5791) <= a and not b;
    layer0_outputs(5792) <= a or b;
    layer0_outputs(5793) <= not (a or b);
    layer0_outputs(5794) <= not a;
    layer0_outputs(5795) <= a or b;
    layer0_outputs(5796) <= not (a and b);
    layer0_outputs(5797) <= not a or b;
    layer0_outputs(5798) <= not (a and b);
    layer0_outputs(5799) <= b;
    layer0_outputs(5800) <= b and not a;
    layer0_outputs(5801) <= not a;
    layer0_outputs(5802) <= a xor b;
    layer0_outputs(5803) <= not (a xor b);
    layer0_outputs(5804) <= not a or b;
    layer0_outputs(5805) <= b and not a;
    layer0_outputs(5806) <= not a or b;
    layer0_outputs(5807) <= not b;
    layer0_outputs(5808) <= a;
    layer0_outputs(5809) <= a xor b;
    layer0_outputs(5810) <= b and not a;
    layer0_outputs(5811) <= 1'b1;
    layer0_outputs(5812) <= b and not a;
    layer0_outputs(5813) <= a and not b;
    layer0_outputs(5814) <= not b;
    layer0_outputs(5815) <= not b;
    layer0_outputs(5816) <= not (a xor b);
    layer0_outputs(5817) <= a or b;
    layer0_outputs(5818) <= not (a xor b);
    layer0_outputs(5819) <= a or b;
    layer0_outputs(5820) <= b and not a;
    layer0_outputs(5821) <= not b;
    layer0_outputs(5822) <= b and not a;
    layer0_outputs(5823) <= b;
    layer0_outputs(5824) <= not b;
    layer0_outputs(5825) <= not b;
    layer0_outputs(5826) <= not (a or b);
    layer0_outputs(5827) <= a;
    layer0_outputs(5828) <= 1'b1;
    layer0_outputs(5829) <= not (a xor b);
    layer0_outputs(5830) <= a and b;
    layer0_outputs(5831) <= not b or a;
    layer0_outputs(5832) <= a xor b;
    layer0_outputs(5833) <= a and b;
    layer0_outputs(5834) <= not b or a;
    layer0_outputs(5835) <= a or b;
    layer0_outputs(5836) <= 1'b0;
    layer0_outputs(5837) <= a or b;
    layer0_outputs(5838) <= a or b;
    layer0_outputs(5839) <= a;
    layer0_outputs(5840) <= not (a or b);
    layer0_outputs(5841) <= b;
    layer0_outputs(5842) <= a;
    layer0_outputs(5843) <= not a or b;
    layer0_outputs(5844) <= a and b;
    layer0_outputs(5845) <= b and not a;
    layer0_outputs(5846) <= not b;
    layer0_outputs(5847) <= b and not a;
    layer0_outputs(5848) <= a or b;
    layer0_outputs(5849) <= a and not b;
    layer0_outputs(5850) <= a and not b;
    layer0_outputs(5851) <= not b;
    layer0_outputs(5852) <= not a;
    layer0_outputs(5853) <= not b or a;
    layer0_outputs(5854) <= not (a or b);
    layer0_outputs(5855) <= b;
    layer0_outputs(5856) <= not b or a;
    layer0_outputs(5857) <= a or b;
    layer0_outputs(5858) <= a and not b;
    layer0_outputs(5859) <= not (a xor b);
    layer0_outputs(5860) <= not (a or b);
    layer0_outputs(5861) <= not b;
    layer0_outputs(5862) <= not b;
    layer0_outputs(5863) <= b;
    layer0_outputs(5864) <= a and not b;
    layer0_outputs(5865) <= not (a or b);
    layer0_outputs(5866) <= not (a or b);
    layer0_outputs(5867) <= b and not a;
    layer0_outputs(5868) <= a xor b;
    layer0_outputs(5869) <= a or b;
    layer0_outputs(5870) <= a xor b;
    layer0_outputs(5871) <= not (a and b);
    layer0_outputs(5872) <= a and not b;
    layer0_outputs(5873) <= a and not b;
    layer0_outputs(5874) <= not b;
    layer0_outputs(5875) <= not b or a;
    layer0_outputs(5876) <= not b or a;
    layer0_outputs(5877) <= b and not a;
    layer0_outputs(5878) <= not a;
    layer0_outputs(5879) <= not a;
    layer0_outputs(5880) <= not (a or b);
    layer0_outputs(5881) <= not (a xor b);
    layer0_outputs(5882) <= a;
    layer0_outputs(5883) <= a xor b;
    layer0_outputs(5884) <= b;
    layer0_outputs(5885) <= 1'b0;
    layer0_outputs(5886) <= b;
    layer0_outputs(5887) <= b;
    layer0_outputs(5888) <= not a;
    layer0_outputs(5889) <= not (a or b);
    layer0_outputs(5890) <= a and not b;
    layer0_outputs(5891) <= not b;
    layer0_outputs(5892) <= 1'b1;
    layer0_outputs(5893) <= not (a or b);
    layer0_outputs(5894) <= a and not b;
    layer0_outputs(5895) <= a or b;
    layer0_outputs(5896) <= a xor b;
    layer0_outputs(5897) <= a;
    layer0_outputs(5898) <= a;
    layer0_outputs(5899) <= not a;
    layer0_outputs(5900) <= b and not a;
    layer0_outputs(5901) <= a xor b;
    layer0_outputs(5902) <= not b or a;
    layer0_outputs(5903) <= not (a xor b);
    layer0_outputs(5904) <= 1'b1;
    layer0_outputs(5905) <= not (a or b);
    layer0_outputs(5906) <= 1'b0;
    layer0_outputs(5907) <= a;
    layer0_outputs(5908) <= not (a xor b);
    layer0_outputs(5909) <= not a;
    layer0_outputs(5910) <= b and not a;
    layer0_outputs(5911) <= not a or b;
    layer0_outputs(5912) <= b;
    layer0_outputs(5913) <= 1'b1;
    layer0_outputs(5914) <= not a;
    layer0_outputs(5915) <= b and not a;
    layer0_outputs(5916) <= not a;
    layer0_outputs(5917) <= a xor b;
    layer0_outputs(5918) <= not (a xor b);
    layer0_outputs(5919) <= not b or a;
    layer0_outputs(5920) <= b and not a;
    layer0_outputs(5921) <= a or b;
    layer0_outputs(5922) <= not (a or b);
    layer0_outputs(5923) <= a or b;
    layer0_outputs(5924) <= not (a and b);
    layer0_outputs(5925) <= not a or b;
    layer0_outputs(5926) <= not b or a;
    layer0_outputs(5927) <= not (a or b);
    layer0_outputs(5928) <= not (a or b);
    layer0_outputs(5929) <= not (a xor b);
    layer0_outputs(5930) <= 1'b0;
    layer0_outputs(5931) <= not a or b;
    layer0_outputs(5932) <= not (a or b);
    layer0_outputs(5933) <= a xor b;
    layer0_outputs(5934) <= not b or a;
    layer0_outputs(5935) <= a xor b;
    layer0_outputs(5936) <= not b;
    layer0_outputs(5937) <= a or b;
    layer0_outputs(5938) <= not a or b;
    layer0_outputs(5939) <= not b or a;
    layer0_outputs(5940) <= a and not b;
    layer0_outputs(5941) <= not (a or b);
    layer0_outputs(5942) <= not a or b;
    layer0_outputs(5943) <= a;
    layer0_outputs(5944) <= a or b;
    layer0_outputs(5945) <= not (a and b);
    layer0_outputs(5946) <= a;
    layer0_outputs(5947) <= not a or b;
    layer0_outputs(5948) <= a or b;
    layer0_outputs(5949) <= a xor b;
    layer0_outputs(5950) <= not a;
    layer0_outputs(5951) <= not b;
    layer0_outputs(5952) <= not (a xor b);
    layer0_outputs(5953) <= not a or b;
    layer0_outputs(5954) <= not (a or b);
    layer0_outputs(5955) <= 1'b0;
    layer0_outputs(5956) <= b and not a;
    layer0_outputs(5957) <= a and b;
    layer0_outputs(5958) <= not b;
    layer0_outputs(5959) <= not (a and b);
    layer0_outputs(5960) <= not a;
    layer0_outputs(5961) <= b and not a;
    layer0_outputs(5962) <= b;
    layer0_outputs(5963) <= a and not b;
    layer0_outputs(5964) <= b;
    layer0_outputs(5965) <= not (a xor b);
    layer0_outputs(5966) <= not a or b;
    layer0_outputs(5967) <= not b;
    layer0_outputs(5968) <= not b or a;
    layer0_outputs(5969) <= b;
    layer0_outputs(5970) <= not (a xor b);
    layer0_outputs(5971) <= 1'b1;
    layer0_outputs(5972) <= not (a xor b);
    layer0_outputs(5973) <= b;
    layer0_outputs(5974) <= a and not b;
    layer0_outputs(5975) <= not (a or b);
    layer0_outputs(5976) <= not (a xor b);
    layer0_outputs(5977) <= b and not a;
    layer0_outputs(5978) <= a and not b;
    layer0_outputs(5979) <= 1'b1;
    layer0_outputs(5980) <= a or b;
    layer0_outputs(5981) <= b and not a;
    layer0_outputs(5982) <= not (a xor b);
    layer0_outputs(5983) <= b;
    layer0_outputs(5984) <= a or b;
    layer0_outputs(5985) <= a xor b;
    layer0_outputs(5986) <= b and not a;
    layer0_outputs(5987) <= b;
    layer0_outputs(5988) <= not b or a;
    layer0_outputs(5989) <= a xor b;
    layer0_outputs(5990) <= 1'b0;
    layer0_outputs(5991) <= not (a and b);
    layer0_outputs(5992) <= 1'b0;
    layer0_outputs(5993) <= a and not b;
    layer0_outputs(5994) <= not a;
    layer0_outputs(5995) <= not (a and b);
    layer0_outputs(5996) <= not b;
    layer0_outputs(5997) <= not b or a;
    layer0_outputs(5998) <= not b or a;
    layer0_outputs(5999) <= not a;
    layer0_outputs(6000) <= a and not b;
    layer0_outputs(6001) <= not a or b;
    layer0_outputs(6002) <= a or b;
    layer0_outputs(6003) <= a and not b;
    layer0_outputs(6004) <= a xor b;
    layer0_outputs(6005) <= not (a xor b);
    layer0_outputs(6006) <= a or b;
    layer0_outputs(6007) <= not b;
    layer0_outputs(6008) <= not (a or b);
    layer0_outputs(6009) <= 1'b0;
    layer0_outputs(6010) <= not a;
    layer0_outputs(6011) <= a xor b;
    layer0_outputs(6012) <= a and not b;
    layer0_outputs(6013) <= not b or a;
    layer0_outputs(6014) <= not a;
    layer0_outputs(6015) <= not b;
    layer0_outputs(6016) <= not (a or b);
    layer0_outputs(6017) <= a;
    layer0_outputs(6018) <= not (a xor b);
    layer0_outputs(6019) <= b and not a;
    layer0_outputs(6020) <= not (a or b);
    layer0_outputs(6021) <= a;
    layer0_outputs(6022) <= a and b;
    layer0_outputs(6023) <= a;
    layer0_outputs(6024) <= not a or b;
    layer0_outputs(6025) <= 1'b0;
    layer0_outputs(6026) <= a and not b;
    layer0_outputs(6027) <= not a;
    layer0_outputs(6028) <= b and not a;
    layer0_outputs(6029) <= a and b;
    layer0_outputs(6030) <= a or b;
    layer0_outputs(6031) <= 1'b1;
    layer0_outputs(6032) <= a or b;
    layer0_outputs(6033) <= a or b;
    layer0_outputs(6034) <= not a;
    layer0_outputs(6035) <= b and not a;
    layer0_outputs(6036) <= a or b;
    layer0_outputs(6037) <= 1'b0;
    layer0_outputs(6038) <= a;
    layer0_outputs(6039) <= 1'b0;
    layer0_outputs(6040) <= not (a or b);
    layer0_outputs(6041) <= b and not a;
    layer0_outputs(6042) <= a and not b;
    layer0_outputs(6043) <= b;
    layer0_outputs(6044) <= a and not b;
    layer0_outputs(6045) <= a or b;
    layer0_outputs(6046) <= b and not a;
    layer0_outputs(6047) <= a or b;
    layer0_outputs(6048) <= not (a xor b);
    layer0_outputs(6049) <= not b;
    layer0_outputs(6050) <= not (a xor b);
    layer0_outputs(6051) <= not a or b;
    layer0_outputs(6052) <= b and not a;
    layer0_outputs(6053) <= 1'b1;
    layer0_outputs(6054) <= a and b;
    layer0_outputs(6055) <= b;
    layer0_outputs(6056) <= not a or b;
    layer0_outputs(6057) <= a xor b;
    layer0_outputs(6058) <= a xor b;
    layer0_outputs(6059) <= a and not b;
    layer0_outputs(6060) <= not a;
    layer0_outputs(6061) <= 1'b1;
    layer0_outputs(6062) <= a or b;
    layer0_outputs(6063) <= a;
    layer0_outputs(6064) <= 1'b1;
    layer0_outputs(6065) <= a;
    layer0_outputs(6066) <= 1'b0;
    layer0_outputs(6067) <= a or b;
    layer0_outputs(6068) <= a and not b;
    layer0_outputs(6069) <= b;
    layer0_outputs(6070) <= 1'b0;
    layer0_outputs(6071) <= not a;
    layer0_outputs(6072) <= not (a and b);
    layer0_outputs(6073) <= a xor b;
    layer0_outputs(6074) <= not b;
    layer0_outputs(6075) <= a or b;
    layer0_outputs(6076) <= b;
    layer0_outputs(6077) <= not (a xor b);
    layer0_outputs(6078) <= b;
    layer0_outputs(6079) <= b and not a;
    layer0_outputs(6080) <= a xor b;
    layer0_outputs(6081) <= not b;
    layer0_outputs(6082) <= a;
    layer0_outputs(6083) <= a and not b;
    layer0_outputs(6084) <= a and b;
    layer0_outputs(6085) <= not (a or b);
    layer0_outputs(6086) <= a;
    layer0_outputs(6087) <= not (a or b);
    layer0_outputs(6088) <= a or b;
    layer0_outputs(6089) <= b;
    layer0_outputs(6090) <= not a;
    layer0_outputs(6091) <= not (a or b);
    layer0_outputs(6092) <= 1'b0;
    layer0_outputs(6093) <= a xor b;
    layer0_outputs(6094) <= b;
    layer0_outputs(6095) <= 1'b1;
    layer0_outputs(6096) <= not (a or b);
    layer0_outputs(6097) <= b and not a;
    layer0_outputs(6098) <= not b;
    layer0_outputs(6099) <= not (a or b);
    layer0_outputs(6100) <= b and not a;
    layer0_outputs(6101) <= not a or b;
    layer0_outputs(6102) <= 1'b0;
    layer0_outputs(6103) <= b;
    layer0_outputs(6104) <= b;
    layer0_outputs(6105) <= a;
    layer0_outputs(6106) <= not a;
    layer0_outputs(6107) <= a or b;
    layer0_outputs(6108) <= not (a xor b);
    layer0_outputs(6109) <= not (a xor b);
    layer0_outputs(6110) <= a and not b;
    layer0_outputs(6111) <= not a;
    layer0_outputs(6112) <= b;
    layer0_outputs(6113) <= a and not b;
    layer0_outputs(6114) <= a and b;
    layer0_outputs(6115) <= not a;
    layer0_outputs(6116) <= a and not b;
    layer0_outputs(6117) <= a and not b;
    layer0_outputs(6118) <= not (a and b);
    layer0_outputs(6119) <= a xor b;
    layer0_outputs(6120) <= not (a or b);
    layer0_outputs(6121) <= not b or a;
    layer0_outputs(6122) <= a or b;
    layer0_outputs(6123) <= a xor b;
    layer0_outputs(6124) <= not a;
    layer0_outputs(6125) <= a and not b;
    layer0_outputs(6126) <= a and not b;
    layer0_outputs(6127) <= a or b;
    layer0_outputs(6128) <= not (a xor b);
    layer0_outputs(6129) <= b;
    layer0_outputs(6130) <= a and b;
    layer0_outputs(6131) <= not (a or b);
    layer0_outputs(6132) <= 1'b0;
    layer0_outputs(6133) <= not b;
    layer0_outputs(6134) <= not (a xor b);
    layer0_outputs(6135) <= not (a xor b);
    layer0_outputs(6136) <= not b or a;
    layer0_outputs(6137) <= a and not b;
    layer0_outputs(6138) <= not b;
    layer0_outputs(6139) <= not (a xor b);
    layer0_outputs(6140) <= b;
    layer0_outputs(6141) <= 1'b0;
    layer0_outputs(6142) <= a;
    layer0_outputs(6143) <= a and not b;
    layer0_outputs(6144) <= not a;
    layer0_outputs(6145) <= not (a and b);
    layer0_outputs(6146) <= a or b;
    layer0_outputs(6147) <= not (a xor b);
    layer0_outputs(6148) <= a and not b;
    layer0_outputs(6149) <= not a or b;
    layer0_outputs(6150) <= a or b;
    layer0_outputs(6151) <= not (a and b);
    layer0_outputs(6152) <= b;
    layer0_outputs(6153) <= a and not b;
    layer0_outputs(6154) <= a or b;
    layer0_outputs(6155) <= not a or b;
    layer0_outputs(6156) <= not (a or b);
    layer0_outputs(6157) <= not (a or b);
    layer0_outputs(6158) <= not a or b;
    layer0_outputs(6159) <= not a;
    layer0_outputs(6160) <= a or b;
    layer0_outputs(6161) <= a xor b;
    layer0_outputs(6162) <= a or b;
    layer0_outputs(6163) <= 1'b1;
    layer0_outputs(6164) <= not (a xor b);
    layer0_outputs(6165) <= a xor b;
    layer0_outputs(6166) <= b;
    layer0_outputs(6167) <= a and b;
    layer0_outputs(6168) <= not (a or b);
    layer0_outputs(6169) <= not (a xor b);
    layer0_outputs(6170) <= a xor b;
    layer0_outputs(6171) <= b;
    layer0_outputs(6172) <= not a;
    layer0_outputs(6173) <= a and b;
    layer0_outputs(6174) <= b;
    layer0_outputs(6175) <= b;
    layer0_outputs(6176) <= b;
    layer0_outputs(6177) <= not (a xor b);
    layer0_outputs(6178) <= a or b;
    layer0_outputs(6179) <= b and not a;
    layer0_outputs(6180) <= a xor b;
    layer0_outputs(6181) <= a or b;
    layer0_outputs(6182) <= a;
    layer0_outputs(6183) <= a or b;
    layer0_outputs(6184) <= not (a or b);
    layer0_outputs(6185) <= not (a xor b);
    layer0_outputs(6186) <= a xor b;
    layer0_outputs(6187) <= not (a and b);
    layer0_outputs(6188) <= not (a or b);
    layer0_outputs(6189) <= not a;
    layer0_outputs(6190) <= b;
    layer0_outputs(6191) <= a xor b;
    layer0_outputs(6192) <= not b;
    layer0_outputs(6193) <= a xor b;
    layer0_outputs(6194) <= b;
    layer0_outputs(6195) <= not a;
    layer0_outputs(6196) <= a;
    layer0_outputs(6197) <= a and b;
    layer0_outputs(6198) <= not (a or b);
    layer0_outputs(6199) <= a or b;
    layer0_outputs(6200) <= a and not b;
    layer0_outputs(6201) <= a xor b;
    layer0_outputs(6202) <= b;
    layer0_outputs(6203) <= b;
    layer0_outputs(6204) <= a;
    layer0_outputs(6205) <= a xor b;
    layer0_outputs(6206) <= not b or a;
    layer0_outputs(6207) <= not (a xor b);
    layer0_outputs(6208) <= a;
    layer0_outputs(6209) <= a;
    layer0_outputs(6210) <= not b;
    layer0_outputs(6211) <= not (a xor b);
    layer0_outputs(6212) <= a or b;
    layer0_outputs(6213) <= not a;
    layer0_outputs(6214) <= a;
    layer0_outputs(6215) <= not (a or b);
    layer0_outputs(6216) <= not (a xor b);
    layer0_outputs(6217) <= not (a xor b);
    layer0_outputs(6218) <= not b;
    layer0_outputs(6219) <= a;
    layer0_outputs(6220) <= a xor b;
    layer0_outputs(6221) <= not (a or b);
    layer0_outputs(6222) <= a or b;
    layer0_outputs(6223) <= not a or b;
    layer0_outputs(6224) <= not (a xor b);
    layer0_outputs(6225) <= not a or b;
    layer0_outputs(6226) <= 1'b0;
    layer0_outputs(6227) <= a xor b;
    layer0_outputs(6228) <= not a;
    layer0_outputs(6229) <= not b or a;
    layer0_outputs(6230) <= not (a xor b);
    layer0_outputs(6231) <= a and not b;
    layer0_outputs(6232) <= a;
    layer0_outputs(6233) <= not a;
    layer0_outputs(6234) <= a and not b;
    layer0_outputs(6235) <= a or b;
    layer0_outputs(6236) <= a xor b;
    layer0_outputs(6237) <= b;
    layer0_outputs(6238) <= b and not a;
    layer0_outputs(6239) <= a or b;
    layer0_outputs(6240) <= b and not a;
    layer0_outputs(6241) <= a or b;
    layer0_outputs(6242) <= not a or b;
    layer0_outputs(6243) <= a xor b;
    layer0_outputs(6244) <= a and not b;
    layer0_outputs(6245) <= not (a and b);
    layer0_outputs(6246) <= not (a xor b);
    layer0_outputs(6247) <= a xor b;
    layer0_outputs(6248) <= a or b;
    layer0_outputs(6249) <= a and not b;
    layer0_outputs(6250) <= a or b;
    layer0_outputs(6251) <= b and not a;
    layer0_outputs(6252) <= a;
    layer0_outputs(6253) <= not b or a;
    layer0_outputs(6254) <= a;
    layer0_outputs(6255) <= not (a xor b);
    layer0_outputs(6256) <= a;
    layer0_outputs(6257) <= not (a xor b);
    layer0_outputs(6258) <= not a;
    layer0_outputs(6259) <= not a or b;
    layer0_outputs(6260) <= not a;
    layer0_outputs(6261) <= a xor b;
    layer0_outputs(6262) <= not b or a;
    layer0_outputs(6263) <= not (a xor b);
    layer0_outputs(6264) <= a or b;
    layer0_outputs(6265) <= 1'b1;
    layer0_outputs(6266) <= a or b;
    layer0_outputs(6267) <= a xor b;
    layer0_outputs(6268) <= a;
    layer0_outputs(6269) <= not (a or b);
    layer0_outputs(6270) <= not (a xor b);
    layer0_outputs(6271) <= not (a xor b);
    layer0_outputs(6272) <= not a;
    layer0_outputs(6273) <= b and not a;
    layer0_outputs(6274) <= not (a or b);
    layer0_outputs(6275) <= not (a or b);
    layer0_outputs(6276) <= not (a or b);
    layer0_outputs(6277) <= a xor b;
    layer0_outputs(6278) <= not b or a;
    layer0_outputs(6279) <= a or b;
    layer0_outputs(6280) <= a or b;
    layer0_outputs(6281) <= a xor b;
    layer0_outputs(6282) <= b;
    layer0_outputs(6283) <= a and not b;
    layer0_outputs(6284) <= not a;
    layer0_outputs(6285) <= a and not b;
    layer0_outputs(6286) <= not (a or b);
    layer0_outputs(6287) <= not a;
    layer0_outputs(6288) <= not (a xor b);
    layer0_outputs(6289) <= not (a or b);
    layer0_outputs(6290) <= a;
    layer0_outputs(6291) <= not b;
    layer0_outputs(6292) <= a;
    layer0_outputs(6293) <= b;
    layer0_outputs(6294) <= a;
    layer0_outputs(6295) <= not (a xor b);
    layer0_outputs(6296) <= 1'b0;
    layer0_outputs(6297) <= not (a xor b);
    layer0_outputs(6298) <= not (a xor b);
    layer0_outputs(6299) <= not b or a;
    layer0_outputs(6300) <= 1'b1;
    layer0_outputs(6301) <= a xor b;
    layer0_outputs(6302) <= a or b;
    layer0_outputs(6303) <= a xor b;
    layer0_outputs(6304) <= not a;
    layer0_outputs(6305) <= not (a or b);
    layer0_outputs(6306) <= a;
    layer0_outputs(6307) <= not (a xor b);
    layer0_outputs(6308) <= a xor b;
    layer0_outputs(6309) <= a xor b;
    layer0_outputs(6310) <= a or b;
    layer0_outputs(6311) <= a xor b;
    layer0_outputs(6312) <= not b;
    layer0_outputs(6313) <= not (a xor b);
    layer0_outputs(6314) <= a or b;
    layer0_outputs(6315) <= not b or a;
    layer0_outputs(6316) <= not (a or b);
    layer0_outputs(6317) <= a and not b;
    layer0_outputs(6318) <= not b;
    layer0_outputs(6319) <= not (a and b);
    layer0_outputs(6320) <= 1'b1;
    layer0_outputs(6321) <= a xor b;
    layer0_outputs(6322) <= a or b;
    layer0_outputs(6323) <= b and not a;
    layer0_outputs(6324) <= a or b;
    layer0_outputs(6325) <= not a or b;
    layer0_outputs(6326) <= a or b;
    layer0_outputs(6327) <= a and not b;
    layer0_outputs(6328) <= not (a or b);
    layer0_outputs(6329) <= a;
    layer0_outputs(6330) <= not a;
    layer0_outputs(6331) <= not (a or b);
    layer0_outputs(6332) <= not a or b;
    layer0_outputs(6333) <= not a;
    layer0_outputs(6334) <= a;
    layer0_outputs(6335) <= not a;
    layer0_outputs(6336) <= a;
    layer0_outputs(6337) <= a;
    layer0_outputs(6338) <= not a or b;
    layer0_outputs(6339) <= a and b;
    layer0_outputs(6340) <= not (a xor b);
    layer0_outputs(6341) <= a or b;
    layer0_outputs(6342) <= not (a xor b);
    layer0_outputs(6343) <= not (a xor b);
    layer0_outputs(6344) <= a or b;
    layer0_outputs(6345) <= a xor b;
    layer0_outputs(6346) <= not b or a;
    layer0_outputs(6347) <= not a;
    layer0_outputs(6348) <= a xor b;
    layer0_outputs(6349) <= not a or b;
    layer0_outputs(6350) <= a;
    layer0_outputs(6351) <= not a;
    layer0_outputs(6352) <= a and b;
    layer0_outputs(6353) <= not (a and b);
    layer0_outputs(6354) <= a or b;
    layer0_outputs(6355) <= not (a xor b);
    layer0_outputs(6356) <= 1'b1;
    layer0_outputs(6357) <= not b or a;
    layer0_outputs(6358) <= 1'b1;
    layer0_outputs(6359) <= b and not a;
    layer0_outputs(6360) <= not b or a;
    layer0_outputs(6361) <= a or b;
    layer0_outputs(6362) <= not b;
    layer0_outputs(6363) <= not (a or b);
    layer0_outputs(6364) <= 1'b1;
    layer0_outputs(6365) <= not (a xor b);
    layer0_outputs(6366) <= not a or b;
    layer0_outputs(6367) <= not a or b;
    layer0_outputs(6368) <= a;
    layer0_outputs(6369) <= 1'b0;
    layer0_outputs(6370) <= a xor b;
    layer0_outputs(6371) <= b and not a;
    layer0_outputs(6372) <= a and not b;
    layer0_outputs(6373) <= not (a xor b);
    layer0_outputs(6374) <= a and not b;
    layer0_outputs(6375) <= not (a or b);
    layer0_outputs(6376) <= not (a xor b);
    layer0_outputs(6377) <= not b;
    layer0_outputs(6378) <= not a;
    layer0_outputs(6379) <= not (a xor b);
    layer0_outputs(6380) <= a xor b;
    layer0_outputs(6381) <= not (a or b);
    layer0_outputs(6382) <= a xor b;
    layer0_outputs(6383) <= not a or b;
    layer0_outputs(6384) <= 1'b0;
    layer0_outputs(6385) <= not a or b;
    layer0_outputs(6386) <= a or b;
    layer0_outputs(6387) <= not b;
    layer0_outputs(6388) <= not a or b;
    layer0_outputs(6389) <= a and b;
    layer0_outputs(6390) <= a and not b;
    layer0_outputs(6391) <= not (a xor b);
    layer0_outputs(6392) <= not (a or b);
    layer0_outputs(6393) <= not b;
    layer0_outputs(6394) <= 1'b1;
    layer0_outputs(6395) <= b;
    layer0_outputs(6396) <= not (a xor b);
    layer0_outputs(6397) <= a or b;
    layer0_outputs(6398) <= 1'b1;
    layer0_outputs(6399) <= not (a and b);
    layer0_outputs(6400) <= b and not a;
    layer0_outputs(6401) <= a;
    layer0_outputs(6402) <= not (a or b);
    layer0_outputs(6403) <= b and not a;
    layer0_outputs(6404) <= not (a xor b);
    layer0_outputs(6405) <= not a;
    layer0_outputs(6406) <= a or b;
    layer0_outputs(6407) <= not a;
    layer0_outputs(6408) <= a;
    layer0_outputs(6409) <= not (a or b);
    layer0_outputs(6410) <= a xor b;
    layer0_outputs(6411) <= not (a xor b);
    layer0_outputs(6412) <= not (a or b);
    layer0_outputs(6413) <= a and not b;
    layer0_outputs(6414) <= not (a xor b);
    layer0_outputs(6415) <= a xor b;
    layer0_outputs(6416) <= b;
    layer0_outputs(6417) <= a xor b;
    layer0_outputs(6418) <= not b;
    layer0_outputs(6419) <= 1'b0;
    layer0_outputs(6420) <= a xor b;
    layer0_outputs(6421) <= b;
    layer0_outputs(6422) <= not (a xor b);
    layer0_outputs(6423) <= b and not a;
    layer0_outputs(6424) <= a;
    layer0_outputs(6425) <= a xor b;
    layer0_outputs(6426) <= a or b;
    layer0_outputs(6427) <= a or b;
    layer0_outputs(6428) <= not b;
    layer0_outputs(6429) <= not b or a;
    layer0_outputs(6430) <= a or b;
    layer0_outputs(6431) <= a or b;
    layer0_outputs(6432) <= not (a and b);
    layer0_outputs(6433) <= not (a xor b);
    layer0_outputs(6434) <= not (a or b);
    layer0_outputs(6435) <= not a;
    layer0_outputs(6436) <= not a;
    layer0_outputs(6437) <= a or b;
    layer0_outputs(6438) <= not (a or b);
    layer0_outputs(6439) <= not (a or b);
    layer0_outputs(6440) <= a or b;
    layer0_outputs(6441) <= a or b;
    layer0_outputs(6442) <= not b or a;
    layer0_outputs(6443) <= b and not a;
    layer0_outputs(6444) <= a and not b;
    layer0_outputs(6445) <= a xor b;
    layer0_outputs(6446) <= b;
    layer0_outputs(6447) <= a or b;
    layer0_outputs(6448) <= not b;
    layer0_outputs(6449) <= a;
    layer0_outputs(6450) <= not a;
    layer0_outputs(6451) <= not (a xor b);
    layer0_outputs(6452) <= a or b;
    layer0_outputs(6453) <= a and b;
    layer0_outputs(6454) <= not a or b;
    layer0_outputs(6455) <= not (a or b);
    layer0_outputs(6456) <= a and b;
    layer0_outputs(6457) <= b;
    layer0_outputs(6458) <= not b or a;
    layer0_outputs(6459) <= a xor b;
    layer0_outputs(6460) <= not b or a;
    layer0_outputs(6461) <= a and not b;
    layer0_outputs(6462) <= a xor b;
    layer0_outputs(6463) <= a;
    layer0_outputs(6464) <= not (a or b);
    layer0_outputs(6465) <= a or b;
    layer0_outputs(6466) <= not a;
    layer0_outputs(6467) <= not (a or b);
    layer0_outputs(6468) <= not (a xor b);
    layer0_outputs(6469) <= not a or b;
    layer0_outputs(6470) <= a;
    layer0_outputs(6471) <= not (a or b);
    layer0_outputs(6472) <= not (a and b);
    layer0_outputs(6473) <= a xor b;
    layer0_outputs(6474) <= not (a xor b);
    layer0_outputs(6475) <= 1'b1;
    layer0_outputs(6476) <= not (a xor b);
    layer0_outputs(6477) <= not (a xor b);
    layer0_outputs(6478) <= a or b;
    layer0_outputs(6479) <= b and not a;
    layer0_outputs(6480) <= not b;
    layer0_outputs(6481) <= b;
    layer0_outputs(6482) <= a and not b;
    layer0_outputs(6483) <= b and not a;
    layer0_outputs(6484) <= 1'b1;
    layer0_outputs(6485) <= not a or b;
    layer0_outputs(6486) <= not (a and b);
    layer0_outputs(6487) <= not a or b;
    layer0_outputs(6488) <= not b or a;
    layer0_outputs(6489) <= a xor b;
    layer0_outputs(6490) <= not a;
    layer0_outputs(6491) <= a;
    layer0_outputs(6492) <= b and not a;
    layer0_outputs(6493) <= not (a or b);
    layer0_outputs(6494) <= not a;
    layer0_outputs(6495) <= not (a and b);
    layer0_outputs(6496) <= 1'b1;
    layer0_outputs(6497) <= a and not b;
    layer0_outputs(6498) <= a xor b;
    layer0_outputs(6499) <= a or b;
    layer0_outputs(6500) <= not (a and b);
    layer0_outputs(6501) <= not b;
    layer0_outputs(6502) <= not b or a;
    layer0_outputs(6503) <= not (a xor b);
    layer0_outputs(6504) <= not a;
    layer0_outputs(6505) <= not (a or b);
    layer0_outputs(6506) <= a or b;
    layer0_outputs(6507) <= not b;
    layer0_outputs(6508) <= not (a xor b);
    layer0_outputs(6509) <= not (a xor b);
    layer0_outputs(6510) <= b;
    layer0_outputs(6511) <= not (a xor b);
    layer0_outputs(6512) <= not b or a;
    layer0_outputs(6513) <= b and not a;
    layer0_outputs(6514) <= not b;
    layer0_outputs(6515) <= a;
    layer0_outputs(6516) <= not a or b;
    layer0_outputs(6517) <= not a or b;
    layer0_outputs(6518) <= b;
    layer0_outputs(6519) <= a or b;
    layer0_outputs(6520) <= not b or a;
    layer0_outputs(6521) <= a and not b;
    layer0_outputs(6522) <= a and not b;
    layer0_outputs(6523) <= not a;
    layer0_outputs(6524) <= a or b;
    layer0_outputs(6525) <= not (a or b);
    layer0_outputs(6526) <= a xor b;
    layer0_outputs(6527) <= a xor b;
    layer0_outputs(6528) <= a xor b;
    layer0_outputs(6529) <= a xor b;
    layer0_outputs(6530) <= not (a or b);
    layer0_outputs(6531) <= not a;
    layer0_outputs(6532) <= a or b;
    layer0_outputs(6533) <= a;
    layer0_outputs(6534) <= b;
    layer0_outputs(6535) <= a and not b;
    layer0_outputs(6536) <= not b or a;
    layer0_outputs(6537) <= not b or a;
    layer0_outputs(6538) <= a xor b;
    layer0_outputs(6539) <= not (a xor b);
    layer0_outputs(6540) <= a;
    layer0_outputs(6541) <= not a or b;
    layer0_outputs(6542) <= not b;
    layer0_outputs(6543) <= a xor b;
    layer0_outputs(6544) <= not a or b;
    layer0_outputs(6545) <= not (a xor b);
    layer0_outputs(6546) <= a xor b;
    layer0_outputs(6547) <= b and not a;
    layer0_outputs(6548) <= not (a or b);
    layer0_outputs(6549) <= a;
    layer0_outputs(6550) <= 1'b1;
    layer0_outputs(6551) <= not a or b;
    layer0_outputs(6552) <= not b;
    layer0_outputs(6553) <= not a;
    layer0_outputs(6554) <= a xor b;
    layer0_outputs(6555) <= a;
    layer0_outputs(6556) <= a or b;
    layer0_outputs(6557) <= not (a and b);
    layer0_outputs(6558) <= a or b;
    layer0_outputs(6559) <= a or b;
    layer0_outputs(6560) <= not a or b;
    layer0_outputs(6561) <= b;
    layer0_outputs(6562) <= not b or a;
    layer0_outputs(6563) <= not b;
    layer0_outputs(6564) <= a and not b;
    layer0_outputs(6565) <= a and not b;
    layer0_outputs(6566) <= not (a xor b);
    layer0_outputs(6567) <= a or b;
    layer0_outputs(6568) <= not (a xor b);
    layer0_outputs(6569) <= b and not a;
    layer0_outputs(6570) <= a and not b;
    layer0_outputs(6571) <= a xor b;
    layer0_outputs(6572) <= not (a or b);
    layer0_outputs(6573) <= b and not a;
    layer0_outputs(6574) <= a and b;
    layer0_outputs(6575) <= a and not b;
    layer0_outputs(6576) <= not (a xor b);
    layer0_outputs(6577) <= b and not a;
    layer0_outputs(6578) <= not (a xor b);
    layer0_outputs(6579) <= 1'b0;
    layer0_outputs(6580) <= b;
    layer0_outputs(6581) <= not a;
    layer0_outputs(6582) <= 1'b0;
    layer0_outputs(6583) <= b;
    layer0_outputs(6584) <= a and not b;
    layer0_outputs(6585) <= not (a or b);
    layer0_outputs(6586) <= a;
    layer0_outputs(6587) <= not a or b;
    layer0_outputs(6588) <= not b;
    layer0_outputs(6589) <= a or b;
    layer0_outputs(6590) <= not a;
    layer0_outputs(6591) <= not b;
    layer0_outputs(6592) <= a;
    layer0_outputs(6593) <= b;
    layer0_outputs(6594) <= not a or b;
    layer0_outputs(6595) <= not a;
    layer0_outputs(6596) <= b;
    layer0_outputs(6597) <= b;
    layer0_outputs(6598) <= b;
    layer0_outputs(6599) <= not (a or b);
    layer0_outputs(6600) <= not (a xor b);
    layer0_outputs(6601) <= b and not a;
    layer0_outputs(6602) <= not b;
    layer0_outputs(6603) <= a or b;
    layer0_outputs(6604) <= not (a xor b);
    layer0_outputs(6605) <= not a or b;
    layer0_outputs(6606) <= not (a or b);
    layer0_outputs(6607) <= 1'b0;
    layer0_outputs(6608) <= a and not b;
    layer0_outputs(6609) <= not a;
    layer0_outputs(6610) <= a and b;
    layer0_outputs(6611) <= not (a or b);
    layer0_outputs(6612) <= not (a and b);
    layer0_outputs(6613) <= not b or a;
    layer0_outputs(6614) <= 1'b0;
    layer0_outputs(6615) <= a xor b;
    layer0_outputs(6616) <= a and not b;
    layer0_outputs(6617) <= a xor b;
    layer0_outputs(6618) <= not (a or b);
    layer0_outputs(6619) <= a;
    layer0_outputs(6620) <= not a;
    layer0_outputs(6621) <= a or b;
    layer0_outputs(6622) <= not (a xor b);
    layer0_outputs(6623) <= a;
    layer0_outputs(6624) <= a;
    layer0_outputs(6625) <= b;
    layer0_outputs(6626) <= not (a xor b);
    layer0_outputs(6627) <= a;
    layer0_outputs(6628) <= not (a and b);
    layer0_outputs(6629) <= a and not b;
    layer0_outputs(6630) <= a or b;
    layer0_outputs(6631) <= a or b;
    layer0_outputs(6632) <= not (a xor b);
    layer0_outputs(6633) <= not b;
    layer0_outputs(6634) <= a or b;
    layer0_outputs(6635) <= not (a xor b);
    layer0_outputs(6636) <= not (a xor b);
    layer0_outputs(6637) <= not b;
    layer0_outputs(6638) <= not b or a;
    layer0_outputs(6639) <= not (a or b);
    layer0_outputs(6640) <= not (a and b);
    layer0_outputs(6641) <= not a or b;
    layer0_outputs(6642) <= a and b;
    layer0_outputs(6643) <= 1'b0;
    layer0_outputs(6644) <= a xor b;
    layer0_outputs(6645) <= a or b;
    layer0_outputs(6646) <= not (a xor b);
    layer0_outputs(6647) <= a or b;
    layer0_outputs(6648) <= not (a or b);
    layer0_outputs(6649) <= not a or b;
    layer0_outputs(6650) <= not (a or b);
    layer0_outputs(6651) <= not b or a;
    layer0_outputs(6652) <= a and b;
    layer0_outputs(6653) <= b;
    layer0_outputs(6654) <= not b;
    layer0_outputs(6655) <= a or b;
    layer0_outputs(6656) <= b and not a;
    layer0_outputs(6657) <= a;
    layer0_outputs(6658) <= not a or b;
    layer0_outputs(6659) <= not (a or b);
    layer0_outputs(6660) <= not (a xor b);
    layer0_outputs(6661) <= not a;
    layer0_outputs(6662) <= not (a and b);
    layer0_outputs(6663) <= not (a or b);
    layer0_outputs(6664) <= not a;
    layer0_outputs(6665) <= not a;
    layer0_outputs(6666) <= b and not a;
    layer0_outputs(6667) <= 1'b1;
    layer0_outputs(6668) <= not (a or b);
    layer0_outputs(6669) <= a and b;
    layer0_outputs(6670) <= not a;
    layer0_outputs(6671) <= not b or a;
    layer0_outputs(6672) <= a and not b;
    layer0_outputs(6673) <= not (a or b);
    layer0_outputs(6674) <= not (a or b);
    layer0_outputs(6675) <= not (a and b);
    layer0_outputs(6676) <= b;
    layer0_outputs(6677) <= a and not b;
    layer0_outputs(6678) <= b;
    layer0_outputs(6679) <= 1'b1;
    layer0_outputs(6680) <= b;
    layer0_outputs(6681) <= not (a or b);
    layer0_outputs(6682) <= a or b;
    layer0_outputs(6683) <= a or b;
    layer0_outputs(6684) <= not (a or b);
    layer0_outputs(6685) <= not b or a;
    layer0_outputs(6686) <= not (a xor b);
    layer0_outputs(6687) <= a xor b;
    layer0_outputs(6688) <= not b or a;
    layer0_outputs(6689) <= a or b;
    layer0_outputs(6690) <= a or b;
    layer0_outputs(6691) <= not (a xor b);
    layer0_outputs(6692) <= not a or b;
    layer0_outputs(6693) <= a;
    layer0_outputs(6694) <= not a;
    layer0_outputs(6695) <= not (a or b);
    layer0_outputs(6696) <= a and not b;
    layer0_outputs(6697) <= not (a xor b);
    layer0_outputs(6698) <= not a or b;
    layer0_outputs(6699) <= a or b;
    layer0_outputs(6700) <= a and not b;
    layer0_outputs(6701) <= b;
    layer0_outputs(6702) <= not (a or b);
    layer0_outputs(6703) <= a or b;
    layer0_outputs(6704) <= a;
    layer0_outputs(6705) <= a xor b;
    layer0_outputs(6706) <= a xor b;
    layer0_outputs(6707) <= a xor b;
    layer0_outputs(6708) <= a xor b;
    layer0_outputs(6709) <= not (a xor b);
    layer0_outputs(6710) <= a and not b;
    layer0_outputs(6711) <= a or b;
    layer0_outputs(6712) <= b and not a;
    layer0_outputs(6713) <= b and not a;
    layer0_outputs(6714) <= not b or a;
    layer0_outputs(6715) <= a;
    layer0_outputs(6716) <= not b;
    layer0_outputs(6717) <= not a;
    layer0_outputs(6718) <= not (a or b);
    layer0_outputs(6719) <= 1'b1;
    layer0_outputs(6720) <= not a or b;
    layer0_outputs(6721) <= not (a or b);
    layer0_outputs(6722) <= not a or b;
    layer0_outputs(6723) <= a and not b;
    layer0_outputs(6724) <= a or b;
    layer0_outputs(6725) <= not (a xor b);
    layer0_outputs(6726) <= a;
    layer0_outputs(6727) <= b and not a;
    layer0_outputs(6728) <= a or b;
    layer0_outputs(6729) <= a;
    layer0_outputs(6730) <= a or b;
    layer0_outputs(6731) <= not b or a;
    layer0_outputs(6732) <= not b;
    layer0_outputs(6733) <= not a or b;
    layer0_outputs(6734) <= not a or b;
    layer0_outputs(6735) <= a and b;
    layer0_outputs(6736) <= not a or b;
    layer0_outputs(6737) <= not b;
    layer0_outputs(6738) <= not (a or b);
    layer0_outputs(6739) <= not a or b;
    layer0_outputs(6740) <= b;
    layer0_outputs(6741) <= b;
    layer0_outputs(6742) <= a or b;
    layer0_outputs(6743) <= not (a xor b);
    layer0_outputs(6744) <= a xor b;
    layer0_outputs(6745) <= 1'b1;
    layer0_outputs(6746) <= not b;
    layer0_outputs(6747) <= a;
    layer0_outputs(6748) <= not a;
    layer0_outputs(6749) <= a and not b;
    layer0_outputs(6750) <= not b;
    layer0_outputs(6751) <= not (a xor b);
    layer0_outputs(6752) <= a or b;
    layer0_outputs(6753) <= not a or b;
    layer0_outputs(6754) <= a and not b;
    layer0_outputs(6755) <= a;
    layer0_outputs(6756) <= b and not a;
    layer0_outputs(6757) <= a or b;
    layer0_outputs(6758) <= not a;
    layer0_outputs(6759) <= not a or b;
    layer0_outputs(6760) <= b and not a;
    layer0_outputs(6761) <= not b or a;
    layer0_outputs(6762) <= not a;
    layer0_outputs(6763) <= a and not b;
    layer0_outputs(6764) <= b and not a;
    layer0_outputs(6765) <= not (a xor b);
    layer0_outputs(6766) <= not (a xor b);
    layer0_outputs(6767) <= a and not b;
    layer0_outputs(6768) <= a or b;
    layer0_outputs(6769) <= a xor b;
    layer0_outputs(6770) <= not (a and b);
    layer0_outputs(6771) <= a or b;
    layer0_outputs(6772) <= not a;
    layer0_outputs(6773) <= a or b;
    layer0_outputs(6774) <= not (a or b);
    layer0_outputs(6775) <= a and not b;
    layer0_outputs(6776) <= not (a and b);
    layer0_outputs(6777) <= not (a or b);
    layer0_outputs(6778) <= a xor b;
    layer0_outputs(6779) <= b;
    layer0_outputs(6780) <= a xor b;
    layer0_outputs(6781) <= a or b;
    layer0_outputs(6782) <= a and not b;
    layer0_outputs(6783) <= b;
    layer0_outputs(6784) <= not a;
    layer0_outputs(6785) <= not b;
    layer0_outputs(6786) <= a xor b;
    layer0_outputs(6787) <= not (a or b);
    layer0_outputs(6788) <= a xor b;
    layer0_outputs(6789) <= not b or a;
    layer0_outputs(6790) <= a xor b;
    layer0_outputs(6791) <= 1'b1;
    layer0_outputs(6792) <= a xor b;
    layer0_outputs(6793) <= a and b;
    layer0_outputs(6794) <= not b;
    layer0_outputs(6795) <= not (a and b);
    layer0_outputs(6796) <= not (a or b);
    layer0_outputs(6797) <= 1'b0;
    layer0_outputs(6798) <= a;
    layer0_outputs(6799) <= a or b;
    layer0_outputs(6800) <= a xor b;
    layer0_outputs(6801) <= not (a xor b);
    layer0_outputs(6802) <= not a or b;
    layer0_outputs(6803) <= a xor b;
    layer0_outputs(6804) <= not b or a;
    layer0_outputs(6805) <= not b or a;
    layer0_outputs(6806) <= b and not a;
    layer0_outputs(6807) <= b and not a;
    layer0_outputs(6808) <= a or b;
    layer0_outputs(6809) <= b and not a;
    layer0_outputs(6810) <= not b;
    layer0_outputs(6811) <= a;
    layer0_outputs(6812) <= not a or b;
    layer0_outputs(6813) <= a xor b;
    layer0_outputs(6814) <= a xor b;
    layer0_outputs(6815) <= a or b;
    layer0_outputs(6816) <= b;
    layer0_outputs(6817) <= b and not a;
    layer0_outputs(6818) <= a;
    layer0_outputs(6819) <= a and not b;
    layer0_outputs(6820) <= a xor b;
    layer0_outputs(6821) <= not b;
    layer0_outputs(6822) <= a or b;
    layer0_outputs(6823) <= b;
    layer0_outputs(6824) <= a xor b;
    layer0_outputs(6825) <= a;
    layer0_outputs(6826) <= not (a or b);
    layer0_outputs(6827) <= not (a xor b);
    layer0_outputs(6828) <= not (a xor b);
    layer0_outputs(6829) <= a xor b;
    layer0_outputs(6830) <= not a or b;
    layer0_outputs(6831) <= not a or b;
    layer0_outputs(6832) <= a or b;
    layer0_outputs(6833) <= not (a or b);
    layer0_outputs(6834) <= a and not b;
    layer0_outputs(6835) <= 1'b1;
    layer0_outputs(6836) <= not b or a;
    layer0_outputs(6837) <= not b;
    layer0_outputs(6838) <= not (a or b);
    layer0_outputs(6839) <= not (a or b);
    layer0_outputs(6840) <= not b or a;
    layer0_outputs(6841) <= not a;
    layer0_outputs(6842) <= not b or a;
    layer0_outputs(6843) <= not (a or b);
    layer0_outputs(6844) <= not (a or b);
    layer0_outputs(6845) <= a xor b;
    layer0_outputs(6846) <= a or b;
    layer0_outputs(6847) <= not (a xor b);
    layer0_outputs(6848) <= b;
    layer0_outputs(6849) <= b;
    layer0_outputs(6850) <= a;
    layer0_outputs(6851) <= a or b;
    layer0_outputs(6852) <= not (a or b);
    layer0_outputs(6853) <= a;
    layer0_outputs(6854) <= not a;
    layer0_outputs(6855) <= b and not a;
    layer0_outputs(6856) <= 1'b1;
    layer0_outputs(6857) <= a or b;
    layer0_outputs(6858) <= not (a xor b);
    layer0_outputs(6859) <= a xor b;
    layer0_outputs(6860) <= not (a xor b);
    layer0_outputs(6861) <= 1'b1;
    layer0_outputs(6862) <= a and not b;
    layer0_outputs(6863) <= not a or b;
    layer0_outputs(6864) <= a and b;
    layer0_outputs(6865) <= a and b;
    layer0_outputs(6866) <= not b;
    layer0_outputs(6867) <= not b or a;
    layer0_outputs(6868) <= a or b;
    layer0_outputs(6869) <= not a or b;
    layer0_outputs(6870) <= 1'b1;
    layer0_outputs(6871) <= not b or a;
    layer0_outputs(6872) <= a and not b;
    layer0_outputs(6873) <= not a;
    layer0_outputs(6874) <= not (a or b);
    layer0_outputs(6875) <= not a;
    layer0_outputs(6876) <= a xor b;
    layer0_outputs(6877) <= not b or a;
    layer0_outputs(6878) <= not (a and b);
    layer0_outputs(6879) <= a or b;
    layer0_outputs(6880) <= not b;
    layer0_outputs(6881) <= not (a xor b);
    layer0_outputs(6882) <= not (a xor b);
    layer0_outputs(6883) <= not (a or b);
    layer0_outputs(6884) <= b and not a;
    layer0_outputs(6885) <= a xor b;
    layer0_outputs(6886) <= not (a or b);
    layer0_outputs(6887) <= a xor b;
    layer0_outputs(6888) <= a and not b;
    layer0_outputs(6889) <= a or b;
    layer0_outputs(6890) <= not (a xor b);
    layer0_outputs(6891) <= b;
    layer0_outputs(6892) <= a;
    layer0_outputs(6893) <= 1'b1;
    layer0_outputs(6894) <= a and not b;
    layer0_outputs(6895) <= a and not b;
    layer0_outputs(6896) <= not a or b;
    layer0_outputs(6897) <= not b;
    layer0_outputs(6898) <= not b or a;
    layer0_outputs(6899) <= not (a xor b);
    layer0_outputs(6900) <= b;
    layer0_outputs(6901) <= not (a or b);
    layer0_outputs(6902) <= a and not b;
    layer0_outputs(6903) <= not (a xor b);
    layer0_outputs(6904) <= not (a and b);
    layer0_outputs(6905) <= not a;
    layer0_outputs(6906) <= not (a or b);
    layer0_outputs(6907) <= a xor b;
    layer0_outputs(6908) <= not a;
    layer0_outputs(6909) <= not b or a;
    layer0_outputs(6910) <= a xor b;
    layer0_outputs(6911) <= a or b;
    layer0_outputs(6912) <= not (a or b);
    layer0_outputs(6913) <= a xor b;
    layer0_outputs(6914) <= not b or a;
    layer0_outputs(6915) <= a or b;
    layer0_outputs(6916) <= not (a xor b);
    layer0_outputs(6917) <= a;
    layer0_outputs(6918) <= not (a xor b);
    layer0_outputs(6919) <= not a or b;
    layer0_outputs(6920) <= a xor b;
    layer0_outputs(6921) <= b;
    layer0_outputs(6922) <= a;
    layer0_outputs(6923) <= not b or a;
    layer0_outputs(6924) <= not (a or b);
    layer0_outputs(6925) <= a or b;
    layer0_outputs(6926) <= not b;
    layer0_outputs(6927) <= not b or a;
    layer0_outputs(6928) <= not b;
    layer0_outputs(6929) <= not (a xor b);
    layer0_outputs(6930) <= 1'b0;
    layer0_outputs(6931) <= not (a xor b);
    layer0_outputs(6932) <= a and not b;
    layer0_outputs(6933) <= a xor b;
    layer0_outputs(6934) <= not (a and b);
    layer0_outputs(6935) <= a or b;
    layer0_outputs(6936) <= b and not a;
    layer0_outputs(6937) <= a or b;
    layer0_outputs(6938) <= not b or a;
    layer0_outputs(6939) <= 1'b0;
    layer0_outputs(6940) <= not b;
    layer0_outputs(6941) <= not (a xor b);
    layer0_outputs(6942) <= not (a xor b);
    layer0_outputs(6943) <= not (a xor b);
    layer0_outputs(6944) <= a xor b;
    layer0_outputs(6945) <= a or b;
    layer0_outputs(6946) <= not (a or b);
    layer0_outputs(6947) <= a xor b;
    layer0_outputs(6948) <= 1'b1;
    layer0_outputs(6949) <= not (a xor b);
    layer0_outputs(6950) <= not (a xor b);
    layer0_outputs(6951) <= 1'b1;
    layer0_outputs(6952) <= not (a or b);
    layer0_outputs(6953) <= a;
    layer0_outputs(6954) <= not (a or b);
    layer0_outputs(6955) <= a or b;
    layer0_outputs(6956) <= not (a or b);
    layer0_outputs(6957) <= not a or b;
    layer0_outputs(6958) <= a xor b;
    layer0_outputs(6959) <= not a or b;
    layer0_outputs(6960) <= a xor b;
    layer0_outputs(6961) <= not (a xor b);
    layer0_outputs(6962) <= b;
    layer0_outputs(6963) <= b;
    layer0_outputs(6964) <= not (a or b);
    layer0_outputs(6965) <= not b or a;
    layer0_outputs(6966) <= a xor b;
    layer0_outputs(6967) <= a xor b;
    layer0_outputs(6968) <= not (a and b);
    layer0_outputs(6969) <= not (a or b);
    layer0_outputs(6970) <= a or b;
    layer0_outputs(6971) <= a xor b;
    layer0_outputs(6972) <= a xor b;
    layer0_outputs(6973) <= a and b;
    layer0_outputs(6974) <= not (a xor b);
    layer0_outputs(6975) <= a xor b;
    layer0_outputs(6976) <= a or b;
    layer0_outputs(6977) <= a or b;
    layer0_outputs(6978) <= not b;
    layer0_outputs(6979) <= not a or b;
    layer0_outputs(6980) <= not b;
    layer0_outputs(6981) <= not (a xor b);
    layer0_outputs(6982) <= not (a xor b);
    layer0_outputs(6983) <= not a;
    layer0_outputs(6984) <= not (a or b);
    layer0_outputs(6985) <= a or b;
    layer0_outputs(6986) <= a or b;
    layer0_outputs(6987) <= b;
    layer0_outputs(6988) <= not (a or b);
    layer0_outputs(6989) <= not (a or b);
    layer0_outputs(6990) <= not a or b;
    layer0_outputs(6991) <= b;
    layer0_outputs(6992) <= not b;
    layer0_outputs(6993) <= a xor b;
    layer0_outputs(6994) <= a and not b;
    layer0_outputs(6995) <= not b or a;
    layer0_outputs(6996) <= not a or b;
    layer0_outputs(6997) <= not b or a;
    layer0_outputs(6998) <= a or b;
    layer0_outputs(6999) <= not a or b;
    layer0_outputs(7000) <= 1'b0;
    layer0_outputs(7001) <= b;
    layer0_outputs(7002) <= not a;
    layer0_outputs(7003) <= a xor b;
    layer0_outputs(7004) <= not (a or b);
    layer0_outputs(7005) <= a or b;
    layer0_outputs(7006) <= b and not a;
    layer0_outputs(7007) <= b;
    layer0_outputs(7008) <= not a;
    layer0_outputs(7009) <= b;
    layer0_outputs(7010) <= a or b;
    layer0_outputs(7011) <= a xor b;
    layer0_outputs(7012) <= b and not a;
    layer0_outputs(7013) <= a xor b;
    layer0_outputs(7014) <= not b or a;
    layer0_outputs(7015) <= a;
    layer0_outputs(7016) <= not (a or b);
    layer0_outputs(7017) <= a xor b;
    layer0_outputs(7018) <= not b or a;
    layer0_outputs(7019) <= a;
    layer0_outputs(7020) <= not a;
    layer0_outputs(7021) <= 1'b0;
    layer0_outputs(7022) <= a and not b;
    layer0_outputs(7023) <= not a or b;
    layer0_outputs(7024) <= not (a or b);
    layer0_outputs(7025) <= a or b;
    layer0_outputs(7026) <= a or b;
    layer0_outputs(7027) <= a xor b;
    layer0_outputs(7028) <= not a or b;
    layer0_outputs(7029) <= not b or a;
    layer0_outputs(7030) <= not (a xor b);
    layer0_outputs(7031) <= not b or a;
    layer0_outputs(7032) <= not a or b;
    layer0_outputs(7033) <= 1'b1;
    layer0_outputs(7034) <= not a;
    layer0_outputs(7035) <= a and not b;
    layer0_outputs(7036) <= not b;
    layer0_outputs(7037) <= b and not a;
    layer0_outputs(7038) <= a xor b;
    layer0_outputs(7039) <= a or b;
    layer0_outputs(7040) <= not (a xor b);
    layer0_outputs(7041) <= b and not a;
    layer0_outputs(7042) <= not a;
    layer0_outputs(7043) <= a xor b;
    layer0_outputs(7044) <= not b or a;
    layer0_outputs(7045) <= a xor b;
    layer0_outputs(7046) <= not b;
    layer0_outputs(7047) <= not (a xor b);
    layer0_outputs(7048) <= not (a or b);
    layer0_outputs(7049) <= not a;
    layer0_outputs(7050) <= 1'b0;
    layer0_outputs(7051) <= b;
    layer0_outputs(7052) <= a or b;
    layer0_outputs(7053) <= 1'b1;
    layer0_outputs(7054) <= not (a or b);
    layer0_outputs(7055) <= a and b;
    layer0_outputs(7056) <= not (a xor b);
    layer0_outputs(7057) <= a or b;
    layer0_outputs(7058) <= not (a or b);
    layer0_outputs(7059) <= b;
    layer0_outputs(7060) <= a;
    layer0_outputs(7061) <= a xor b;
    layer0_outputs(7062) <= not (a and b);
    layer0_outputs(7063) <= not (a or b);
    layer0_outputs(7064) <= a;
    layer0_outputs(7065) <= a or b;
    layer0_outputs(7066) <= not (a xor b);
    layer0_outputs(7067) <= not a or b;
    layer0_outputs(7068) <= a xor b;
    layer0_outputs(7069) <= not (a and b);
    layer0_outputs(7070) <= b and not a;
    layer0_outputs(7071) <= a or b;
    layer0_outputs(7072) <= not (a xor b);
    layer0_outputs(7073) <= a xor b;
    layer0_outputs(7074) <= 1'b0;
    layer0_outputs(7075) <= not (a or b);
    layer0_outputs(7076) <= b;
    layer0_outputs(7077) <= a or b;
    layer0_outputs(7078) <= b;
    layer0_outputs(7079) <= a and not b;
    layer0_outputs(7080) <= a xor b;
    layer0_outputs(7081) <= not (a xor b);
    layer0_outputs(7082) <= a xor b;
    layer0_outputs(7083) <= not a;
    layer0_outputs(7084) <= a;
    layer0_outputs(7085) <= b;
    layer0_outputs(7086) <= a and b;
    layer0_outputs(7087) <= not b or a;
    layer0_outputs(7088) <= a;
    layer0_outputs(7089) <= not (a xor b);
    layer0_outputs(7090) <= a and not b;
    layer0_outputs(7091) <= not (a or b);
    layer0_outputs(7092) <= a or b;
    layer0_outputs(7093) <= not (a xor b);
    layer0_outputs(7094) <= not a or b;
    layer0_outputs(7095) <= 1'b1;
    layer0_outputs(7096) <= b;
    layer0_outputs(7097) <= a and not b;
    layer0_outputs(7098) <= not a or b;
    layer0_outputs(7099) <= not (a xor b);
    layer0_outputs(7100) <= a or b;
    layer0_outputs(7101) <= not b or a;
    layer0_outputs(7102) <= not a or b;
    layer0_outputs(7103) <= not a or b;
    layer0_outputs(7104) <= not a or b;
    layer0_outputs(7105) <= not (a or b);
    layer0_outputs(7106) <= 1'b0;
    layer0_outputs(7107) <= not b;
    layer0_outputs(7108) <= b and not a;
    layer0_outputs(7109) <= 1'b1;
    layer0_outputs(7110) <= not b;
    layer0_outputs(7111) <= b;
    layer0_outputs(7112) <= not b or a;
    layer0_outputs(7113) <= 1'b0;
    layer0_outputs(7114) <= b;
    layer0_outputs(7115) <= not b;
    layer0_outputs(7116) <= a or b;
    layer0_outputs(7117) <= a and b;
    layer0_outputs(7118) <= not (a or b);
    layer0_outputs(7119) <= not (a xor b);
    layer0_outputs(7120) <= not b;
    layer0_outputs(7121) <= not a or b;
    layer0_outputs(7122) <= not a;
    layer0_outputs(7123) <= not (a xor b);
    layer0_outputs(7124) <= 1'b0;
    layer0_outputs(7125) <= a xor b;
    layer0_outputs(7126) <= not b;
    layer0_outputs(7127) <= not (a or b);
    layer0_outputs(7128) <= not (a or b);
    layer0_outputs(7129) <= b;
    layer0_outputs(7130) <= b;
    layer0_outputs(7131) <= a;
    layer0_outputs(7132) <= not b;
    layer0_outputs(7133) <= not b;
    layer0_outputs(7134) <= not b;
    layer0_outputs(7135) <= a or b;
    layer0_outputs(7136) <= a xor b;
    layer0_outputs(7137) <= a;
    layer0_outputs(7138) <= a;
    layer0_outputs(7139) <= not a;
    layer0_outputs(7140) <= not b;
    layer0_outputs(7141) <= not (a xor b);
    layer0_outputs(7142) <= a or b;
    layer0_outputs(7143) <= not (a and b);
    layer0_outputs(7144) <= a xor b;
    layer0_outputs(7145) <= a and b;
    layer0_outputs(7146) <= not a or b;
    layer0_outputs(7147) <= not a or b;
    layer0_outputs(7148) <= not (a and b);
    layer0_outputs(7149) <= a or b;
    layer0_outputs(7150) <= a xor b;
    layer0_outputs(7151) <= not a or b;
    layer0_outputs(7152) <= a or b;
    layer0_outputs(7153) <= b and not a;
    layer0_outputs(7154) <= not (a and b);
    layer0_outputs(7155) <= a xor b;
    layer0_outputs(7156) <= a or b;
    layer0_outputs(7157) <= a or b;
    layer0_outputs(7158) <= 1'b0;
    layer0_outputs(7159) <= not b or a;
    layer0_outputs(7160) <= not b or a;
    layer0_outputs(7161) <= b and not a;
    layer0_outputs(7162) <= not (a xor b);
    layer0_outputs(7163) <= not b or a;
    layer0_outputs(7164) <= a or b;
    layer0_outputs(7165) <= not b or a;
    layer0_outputs(7166) <= a or b;
    layer0_outputs(7167) <= 1'b0;
    layer0_outputs(7168) <= not (a or b);
    layer0_outputs(7169) <= not (a xor b);
    layer0_outputs(7170) <= not (a xor b);
    layer0_outputs(7171) <= a;
    layer0_outputs(7172) <= b and not a;
    layer0_outputs(7173) <= a and not b;
    layer0_outputs(7174) <= not b or a;
    layer0_outputs(7175) <= not a;
    layer0_outputs(7176) <= b and not a;
    layer0_outputs(7177) <= not b or a;
    layer0_outputs(7178) <= not (a or b);
    layer0_outputs(7179) <= a xor b;
    layer0_outputs(7180) <= 1'b1;
    layer0_outputs(7181) <= not (a or b);
    layer0_outputs(7182) <= a or b;
    layer0_outputs(7183) <= not (a and b);
    layer0_outputs(7184) <= 1'b1;
    layer0_outputs(7185) <= not b;
    layer0_outputs(7186) <= a xor b;
    layer0_outputs(7187) <= not a or b;
    layer0_outputs(7188) <= not b;
    layer0_outputs(7189) <= not b;
    layer0_outputs(7190) <= not (a xor b);
    layer0_outputs(7191) <= not (a xor b);
    layer0_outputs(7192) <= b;
    layer0_outputs(7193) <= not (a or b);
    layer0_outputs(7194) <= not (a or b);
    layer0_outputs(7195) <= a or b;
    layer0_outputs(7196) <= not (a xor b);
    layer0_outputs(7197) <= a and not b;
    layer0_outputs(7198) <= a and b;
    layer0_outputs(7199) <= not a or b;
    layer0_outputs(7200) <= a;
    layer0_outputs(7201) <= a or b;
    layer0_outputs(7202) <= 1'b1;
    layer0_outputs(7203) <= a;
    layer0_outputs(7204) <= b and not a;
    layer0_outputs(7205) <= a xor b;
    layer0_outputs(7206) <= b and not a;
    layer0_outputs(7207) <= b and not a;
    layer0_outputs(7208) <= a;
    layer0_outputs(7209) <= not b;
    layer0_outputs(7210) <= b;
    layer0_outputs(7211) <= a xor b;
    layer0_outputs(7212) <= a or b;
    layer0_outputs(7213) <= not b;
    layer0_outputs(7214) <= b and not a;
    layer0_outputs(7215) <= 1'b1;
    layer0_outputs(7216) <= a xor b;
    layer0_outputs(7217) <= b and not a;
    layer0_outputs(7218) <= a or b;
    layer0_outputs(7219) <= a xor b;
    layer0_outputs(7220) <= not (a or b);
    layer0_outputs(7221) <= a and not b;
    layer0_outputs(7222) <= not a or b;
    layer0_outputs(7223) <= not (a or b);
    layer0_outputs(7224) <= not b;
    layer0_outputs(7225) <= a xor b;
    layer0_outputs(7226) <= a xor b;
    layer0_outputs(7227) <= not (a xor b);
    layer0_outputs(7228) <= not (a and b);
    layer0_outputs(7229) <= a xor b;
    layer0_outputs(7230) <= not (a xor b);
    layer0_outputs(7231) <= a;
    layer0_outputs(7232) <= not a;
    layer0_outputs(7233) <= b and not a;
    layer0_outputs(7234) <= not (a or b);
    layer0_outputs(7235) <= a and not b;
    layer0_outputs(7236) <= a and not b;
    layer0_outputs(7237) <= a xor b;
    layer0_outputs(7238) <= not (a xor b);
    layer0_outputs(7239) <= not b;
    layer0_outputs(7240) <= not b;
    layer0_outputs(7241) <= not b;
    layer0_outputs(7242) <= a or b;
    layer0_outputs(7243) <= not b or a;
    layer0_outputs(7244) <= not b;
    layer0_outputs(7245) <= not (a or b);
    layer0_outputs(7246) <= not b or a;
    layer0_outputs(7247) <= not (a or b);
    layer0_outputs(7248) <= 1'b1;
    layer0_outputs(7249) <= b;
    layer0_outputs(7250) <= not (a xor b);
    layer0_outputs(7251) <= a or b;
    layer0_outputs(7252) <= a and not b;
    layer0_outputs(7253) <= not (a xor b);
    layer0_outputs(7254) <= not b or a;
    layer0_outputs(7255) <= not (a xor b);
    layer0_outputs(7256) <= b and not a;
    layer0_outputs(7257) <= not a or b;
    layer0_outputs(7258) <= a and not b;
    layer0_outputs(7259) <= b and not a;
    layer0_outputs(7260) <= not a or b;
    layer0_outputs(7261) <= not (a or b);
    layer0_outputs(7262) <= not b;
    layer0_outputs(7263) <= not a;
    layer0_outputs(7264) <= not (a or b);
    layer0_outputs(7265) <= not (a or b);
    layer0_outputs(7266) <= not a or b;
    layer0_outputs(7267) <= not (a or b);
    layer0_outputs(7268) <= not (a or b);
    layer0_outputs(7269) <= a or b;
    layer0_outputs(7270) <= a or b;
    layer0_outputs(7271) <= b and not a;
    layer0_outputs(7272) <= a or b;
    layer0_outputs(7273) <= b and not a;
    layer0_outputs(7274) <= b;
    layer0_outputs(7275) <= b;
    layer0_outputs(7276) <= not b or a;
    layer0_outputs(7277) <= b and not a;
    layer0_outputs(7278) <= not a;
    layer0_outputs(7279) <= a;
    layer0_outputs(7280) <= not a;
    layer0_outputs(7281) <= not (a or b);
    layer0_outputs(7282) <= a;
    layer0_outputs(7283) <= not (a or b);
    layer0_outputs(7284) <= a xor b;
    layer0_outputs(7285) <= not b;
    layer0_outputs(7286) <= not a or b;
    layer0_outputs(7287) <= not (a and b);
    layer0_outputs(7288) <= not b or a;
    layer0_outputs(7289) <= a or b;
    layer0_outputs(7290) <= not a or b;
    layer0_outputs(7291) <= a or b;
    layer0_outputs(7292) <= not a or b;
    layer0_outputs(7293) <= not (a and b);
    layer0_outputs(7294) <= not a;
    layer0_outputs(7295) <= not (a xor b);
    layer0_outputs(7296) <= b and not a;
    layer0_outputs(7297) <= a or b;
    layer0_outputs(7298) <= a xor b;
    layer0_outputs(7299) <= not a;
    layer0_outputs(7300) <= not b;
    layer0_outputs(7301) <= a;
    layer0_outputs(7302) <= a or b;
    layer0_outputs(7303) <= not (a or b);
    layer0_outputs(7304) <= not (a xor b);
    layer0_outputs(7305) <= not b or a;
    layer0_outputs(7306) <= not b or a;
    layer0_outputs(7307) <= not b or a;
    layer0_outputs(7308) <= a xor b;
    layer0_outputs(7309) <= a xor b;
    layer0_outputs(7310) <= b;
    layer0_outputs(7311) <= a xor b;
    layer0_outputs(7312) <= a;
    layer0_outputs(7313) <= not a;
    layer0_outputs(7314) <= not (a or b);
    layer0_outputs(7315) <= not (a xor b);
    layer0_outputs(7316) <= not (a xor b);
    layer0_outputs(7317) <= b and not a;
    layer0_outputs(7318) <= not (a xor b);
    layer0_outputs(7319) <= not (a xor b);
    layer0_outputs(7320) <= 1'b1;
    layer0_outputs(7321) <= not b or a;
    layer0_outputs(7322) <= b and not a;
    layer0_outputs(7323) <= not b or a;
    layer0_outputs(7324) <= 1'b0;
    layer0_outputs(7325) <= not b;
    layer0_outputs(7326) <= b and not a;
    layer0_outputs(7327) <= b and not a;
    layer0_outputs(7328) <= not a or b;
    layer0_outputs(7329) <= not b;
    layer0_outputs(7330) <= not (a or b);
    layer0_outputs(7331) <= b;
    layer0_outputs(7332) <= not b;
    layer0_outputs(7333) <= b and not a;
    layer0_outputs(7334) <= b and not a;
    layer0_outputs(7335) <= b;
    layer0_outputs(7336) <= b;
    layer0_outputs(7337) <= a and not b;
    layer0_outputs(7338) <= a xor b;
    layer0_outputs(7339) <= not (a or b);
    layer0_outputs(7340) <= a or b;
    layer0_outputs(7341) <= not (a or b);
    layer0_outputs(7342) <= b and not a;
    layer0_outputs(7343) <= a and not b;
    layer0_outputs(7344) <= not b or a;
    layer0_outputs(7345) <= not b;
    layer0_outputs(7346) <= a or b;
    layer0_outputs(7347) <= not (a or b);
    layer0_outputs(7348) <= a and not b;
    layer0_outputs(7349) <= not (a or b);
    layer0_outputs(7350) <= not a;
    layer0_outputs(7351) <= not (a or b);
    layer0_outputs(7352) <= not b;
    layer0_outputs(7353) <= b and not a;
    layer0_outputs(7354) <= not b;
    layer0_outputs(7355) <= a;
    layer0_outputs(7356) <= 1'b0;
    layer0_outputs(7357) <= not (a or b);
    layer0_outputs(7358) <= b;
    layer0_outputs(7359) <= a;
    layer0_outputs(7360) <= not a or b;
    layer0_outputs(7361) <= a xor b;
    layer0_outputs(7362) <= not (a or b);
    layer0_outputs(7363) <= a or b;
    layer0_outputs(7364) <= not (a xor b);
    layer0_outputs(7365) <= a or b;
    layer0_outputs(7366) <= not a or b;
    layer0_outputs(7367) <= b;
    layer0_outputs(7368) <= a;
    layer0_outputs(7369) <= not b or a;
    layer0_outputs(7370) <= a or b;
    layer0_outputs(7371) <= not b or a;
    layer0_outputs(7372) <= not (a or b);
    layer0_outputs(7373) <= 1'b0;
    layer0_outputs(7374) <= not b or a;
    layer0_outputs(7375) <= not (a or b);
    layer0_outputs(7376) <= not b or a;
    layer0_outputs(7377) <= not (a or b);
    layer0_outputs(7378) <= b;
    layer0_outputs(7379) <= a and b;
    layer0_outputs(7380) <= not b;
    layer0_outputs(7381) <= a;
    layer0_outputs(7382) <= a or b;
    layer0_outputs(7383) <= a or b;
    layer0_outputs(7384) <= not (a xor b);
    layer0_outputs(7385) <= 1'b1;
    layer0_outputs(7386) <= not (a xor b);
    layer0_outputs(7387) <= not b or a;
    layer0_outputs(7388) <= a or b;
    layer0_outputs(7389) <= b;
    layer0_outputs(7390) <= a or b;
    layer0_outputs(7391) <= not a;
    layer0_outputs(7392) <= not (a or b);
    layer0_outputs(7393) <= b;
    layer0_outputs(7394) <= not (a or b);
    layer0_outputs(7395) <= a;
    layer0_outputs(7396) <= not b or a;
    layer0_outputs(7397) <= a and b;
    layer0_outputs(7398) <= not (a or b);
    layer0_outputs(7399) <= not a;
    layer0_outputs(7400) <= b and not a;
    layer0_outputs(7401) <= not b or a;
    layer0_outputs(7402) <= a;
    layer0_outputs(7403) <= 1'b1;
    layer0_outputs(7404) <= not a or b;
    layer0_outputs(7405) <= not (a and b);
    layer0_outputs(7406) <= not a or b;
    layer0_outputs(7407) <= a xor b;
    layer0_outputs(7408) <= a xor b;
    layer0_outputs(7409) <= not (a xor b);
    layer0_outputs(7410) <= a or b;
    layer0_outputs(7411) <= not b;
    layer0_outputs(7412) <= a or b;
    layer0_outputs(7413) <= not b;
    layer0_outputs(7414) <= a;
    layer0_outputs(7415) <= a and not b;
    layer0_outputs(7416) <= not b or a;
    layer0_outputs(7417) <= not (a or b);
    layer0_outputs(7418) <= not a or b;
    layer0_outputs(7419) <= not b;
    layer0_outputs(7420) <= a;
    layer0_outputs(7421) <= not a;
    layer0_outputs(7422) <= not b or a;
    layer0_outputs(7423) <= a xor b;
    layer0_outputs(7424) <= not b or a;
    layer0_outputs(7425) <= not (a xor b);
    layer0_outputs(7426) <= b;
    layer0_outputs(7427) <= b and not a;
    layer0_outputs(7428) <= a or b;
    layer0_outputs(7429) <= 1'b1;
    layer0_outputs(7430) <= 1'b0;
    layer0_outputs(7431) <= a xor b;
    layer0_outputs(7432) <= not (a or b);
    layer0_outputs(7433) <= not (a or b);
    layer0_outputs(7434) <= not a or b;
    layer0_outputs(7435) <= not a;
    layer0_outputs(7436) <= a or b;
    layer0_outputs(7437) <= not a or b;
    layer0_outputs(7438) <= not (a xor b);
    layer0_outputs(7439) <= not b or a;
    layer0_outputs(7440) <= 1'b1;
    layer0_outputs(7441) <= b and not a;
    layer0_outputs(7442) <= a or b;
    layer0_outputs(7443) <= not (a or b);
    layer0_outputs(7444) <= not (a and b);
    layer0_outputs(7445) <= a or b;
    layer0_outputs(7446) <= a or b;
    layer0_outputs(7447) <= a xor b;
    layer0_outputs(7448) <= a and not b;
    layer0_outputs(7449) <= b and not a;
    layer0_outputs(7450) <= not (a xor b);
    layer0_outputs(7451) <= b and not a;
    layer0_outputs(7452) <= not b;
    layer0_outputs(7453) <= a xor b;
    layer0_outputs(7454) <= a or b;
    layer0_outputs(7455) <= not b;
    layer0_outputs(7456) <= 1'b0;
    layer0_outputs(7457) <= not (a xor b);
    layer0_outputs(7458) <= not a or b;
    layer0_outputs(7459) <= not (a and b);
    layer0_outputs(7460) <= not (a and b);
    layer0_outputs(7461) <= not (a or b);
    layer0_outputs(7462) <= not a;
    layer0_outputs(7463) <= a and b;
    layer0_outputs(7464) <= b and not a;
    layer0_outputs(7465) <= a xor b;
    layer0_outputs(7466) <= a or b;
    layer0_outputs(7467) <= a xor b;
    layer0_outputs(7468) <= not a or b;
    layer0_outputs(7469) <= not (a or b);
    layer0_outputs(7470) <= not b;
    layer0_outputs(7471) <= not (a or b);
    layer0_outputs(7472) <= not a or b;
    layer0_outputs(7473) <= not a or b;
    layer0_outputs(7474) <= not b;
    layer0_outputs(7475) <= not a or b;
    layer0_outputs(7476) <= not b or a;
    layer0_outputs(7477) <= b;
    layer0_outputs(7478) <= a;
    layer0_outputs(7479) <= 1'b0;
    layer0_outputs(7480) <= not (a or b);
    layer0_outputs(7481) <= a or b;
    layer0_outputs(7482) <= b;
    layer0_outputs(7483) <= not b or a;
    layer0_outputs(7484) <= a and b;
    layer0_outputs(7485) <= not a or b;
    layer0_outputs(7486) <= not (a or b);
    layer0_outputs(7487) <= a;
    layer0_outputs(7488) <= a xor b;
    layer0_outputs(7489) <= not (a or b);
    layer0_outputs(7490) <= a;
    layer0_outputs(7491) <= not (a or b);
    layer0_outputs(7492) <= a xor b;
    layer0_outputs(7493) <= not (a and b);
    layer0_outputs(7494) <= a and b;
    layer0_outputs(7495) <= a;
    layer0_outputs(7496) <= b and not a;
    layer0_outputs(7497) <= b;
    layer0_outputs(7498) <= not b;
    layer0_outputs(7499) <= b;
    layer0_outputs(7500) <= a or b;
    layer0_outputs(7501) <= not (a or b);
    layer0_outputs(7502) <= not a or b;
    layer0_outputs(7503) <= a xor b;
    layer0_outputs(7504) <= not (a xor b);
    layer0_outputs(7505) <= not (a xor b);
    layer0_outputs(7506) <= b and not a;
    layer0_outputs(7507) <= a and b;
    layer0_outputs(7508) <= b and not a;
    layer0_outputs(7509) <= a or b;
    layer0_outputs(7510) <= not b or a;
    layer0_outputs(7511) <= b and not a;
    layer0_outputs(7512) <= b;
    layer0_outputs(7513) <= not a;
    layer0_outputs(7514) <= not b;
    layer0_outputs(7515) <= not b;
    layer0_outputs(7516) <= a or b;
    layer0_outputs(7517) <= a xor b;
    layer0_outputs(7518) <= not b;
    layer0_outputs(7519) <= b;
    layer0_outputs(7520) <= a xor b;
    layer0_outputs(7521) <= a;
    layer0_outputs(7522) <= b;
    layer0_outputs(7523) <= 1'b0;
    layer0_outputs(7524) <= a;
    layer0_outputs(7525) <= a or b;
    layer0_outputs(7526) <= not (a or b);
    layer0_outputs(7527) <= a xor b;
    layer0_outputs(7528) <= not (a or b);
    layer0_outputs(7529) <= a xor b;
    layer0_outputs(7530) <= 1'b0;
    layer0_outputs(7531) <= b and not a;
    layer0_outputs(7532) <= b;
    layer0_outputs(7533) <= not b;
    layer0_outputs(7534) <= not a;
    layer0_outputs(7535) <= a or b;
    layer0_outputs(7536) <= not (a xor b);
    layer0_outputs(7537) <= not a;
    layer0_outputs(7538) <= not (a xor b);
    layer0_outputs(7539) <= not (a or b);
    layer0_outputs(7540) <= b and not a;
    layer0_outputs(7541) <= a and not b;
    layer0_outputs(7542) <= not (a xor b);
    layer0_outputs(7543) <= not b;
    layer0_outputs(7544) <= b;
    layer0_outputs(7545) <= a or b;
    layer0_outputs(7546) <= a and not b;
    layer0_outputs(7547) <= 1'b0;
    layer0_outputs(7548) <= not b or a;
    layer0_outputs(7549) <= a or b;
    layer0_outputs(7550) <= a;
    layer0_outputs(7551) <= a or b;
    layer0_outputs(7552) <= not b or a;
    layer0_outputs(7553) <= a xor b;
    layer0_outputs(7554) <= a and not b;
    layer0_outputs(7555) <= b;
    layer0_outputs(7556) <= b;
    layer0_outputs(7557) <= a or b;
    layer0_outputs(7558) <= not a or b;
    layer0_outputs(7559) <= b;
    layer0_outputs(7560) <= not (a or b);
    layer0_outputs(7561) <= a xor b;
    layer0_outputs(7562) <= 1'b0;
    layer0_outputs(7563) <= not a;
    layer0_outputs(7564) <= not b or a;
    layer0_outputs(7565) <= not a;
    layer0_outputs(7566) <= a xor b;
    layer0_outputs(7567) <= a xor b;
    layer0_outputs(7568) <= not (a and b);
    layer0_outputs(7569) <= not b;
    layer0_outputs(7570) <= not b;
    layer0_outputs(7571) <= not (a or b);
    layer0_outputs(7572) <= not (a or b);
    layer0_outputs(7573) <= a and not b;
    layer0_outputs(7574) <= not b or a;
    layer0_outputs(7575) <= a xor b;
    layer0_outputs(7576) <= 1'b1;
    layer0_outputs(7577) <= a or b;
    layer0_outputs(7578) <= a and not b;
    layer0_outputs(7579) <= 1'b0;
    layer0_outputs(7580) <= not (a or b);
    layer0_outputs(7581) <= not (a or b);
    layer0_outputs(7582) <= a xor b;
    layer0_outputs(7583) <= a and not b;
    layer0_outputs(7584) <= a or b;
    layer0_outputs(7585) <= not b or a;
    layer0_outputs(7586) <= not a;
    layer0_outputs(7587) <= a and not b;
    layer0_outputs(7588) <= not (a or b);
    layer0_outputs(7589) <= not a;
    layer0_outputs(7590) <= not (a xor b);
    layer0_outputs(7591) <= 1'b1;
    layer0_outputs(7592) <= b;
    layer0_outputs(7593) <= a and not b;
    layer0_outputs(7594) <= not b;
    layer0_outputs(7595) <= not b or a;
    layer0_outputs(7596) <= not (a and b);
    layer0_outputs(7597) <= not (a and b);
    layer0_outputs(7598) <= a and b;
    layer0_outputs(7599) <= not (a xor b);
    layer0_outputs(7600) <= a and not b;
    layer0_outputs(7601) <= a or b;
    layer0_outputs(7602) <= a or b;
    layer0_outputs(7603) <= not a;
    layer0_outputs(7604) <= not (a or b);
    layer0_outputs(7605) <= not a;
    layer0_outputs(7606) <= not b;
    layer0_outputs(7607) <= not (a xor b);
    layer0_outputs(7608) <= a or b;
    layer0_outputs(7609) <= not (a or b);
    layer0_outputs(7610) <= b and not a;
    layer0_outputs(7611) <= not (a or b);
    layer0_outputs(7612) <= not b or a;
    layer0_outputs(7613) <= not (a or b);
    layer0_outputs(7614) <= not a or b;
    layer0_outputs(7615) <= 1'b0;
    layer0_outputs(7616) <= not (a or b);
    layer0_outputs(7617) <= a and not b;
    layer0_outputs(7618) <= not (a or b);
    layer0_outputs(7619) <= a xor b;
    layer0_outputs(7620) <= not b;
    layer0_outputs(7621) <= not b or a;
    layer0_outputs(7622) <= a and b;
    layer0_outputs(7623) <= a and not b;
    layer0_outputs(7624) <= b and not a;
    layer0_outputs(7625) <= not a;
    layer0_outputs(7626) <= not a or b;
    layer0_outputs(7627) <= a;
    layer0_outputs(7628) <= not (a or b);
    layer0_outputs(7629) <= not (a or b);
    layer0_outputs(7630) <= a;
    layer0_outputs(7631) <= a xor b;
    layer0_outputs(7632) <= a xor b;
    layer0_outputs(7633) <= 1'b1;
    layer0_outputs(7634) <= not (a xor b);
    layer0_outputs(7635) <= not b or a;
    layer0_outputs(7636) <= a;
    layer0_outputs(7637) <= not (a or b);
    layer0_outputs(7638) <= a or b;
    layer0_outputs(7639) <= 1'b0;
    layer0_outputs(7640) <= a and not b;
    layer0_outputs(7641) <= not b or a;
    layer0_outputs(7642) <= a or b;
    layer0_outputs(7643) <= not b;
    layer0_outputs(7644) <= a or b;
    layer0_outputs(7645) <= a or b;
    layer0_outputs(7646) <= a or b;
    layer0_outputs(7647) <= not (a or b);
    layer0_outputs(7648) <= a;
    layer0_outputs(7649) <= not (a or b);
    layer0_outputs(7650) <= a or b;
    layer0_outputs(7651) <= not (a or b);
    layer0_outputs(7652) <= a;
    layer0_outputs(7653) <= not (a xor b);
    layer0_outputs(7654) <= a;
    layer0_outputs(7655) <= not (a or b);
    layer0_outputs(7656) <= not a;
    layer0_outputs(7657) <= a or b;
    layer0_outputs(7658) <= not (a xor b);
    layer0_outputs(7659) <= b and not a;
    layer0_outputs(7660) <= 1'b0;
    layer0_outputs(7661) <= a;
    layer0_outputs(7662) <= a or b;
    layer0_outputs(7663) <= not a or b;
    layer0_outputs(7664) <= a xor b;
    layer0_outputs(7665) <= not a;
    layer0_outputs(7666) <= not (a or b);
    layer0_outputs(7667) <= a or b;
    layer0_outputs(7668) <= not a or b;
    layer0_outputs(7669) <= b;
    layer0_outputs(7670) <= not (a or b);
    layer0_outputs(7671) <= not (a xor b);
    layer0_outputs(7672) <= b and not a;
    layer0_outputs(7673) <= a and not b;
    layer0_outputs(7674) <= a;
    layer0_outputs(7675) <= not a;
    layer0_outputs(7676) <= not (a or b);
    layer0_outputs(7677) <= not (a xor b);
    layer0_outputs(7678) <= not (a xor b);
    layer0_outputs(7679) <= not b or a;
    layer0_outputs(7680) <= b and not a;
    layer0_outputs(7681) <= b;
    layer0_outputs(7682) <= not a;
    layer0_outputs(7683) <= not (a xor b);
    layer0_outputs(7684) <= not a;
    layer0_outputs(7685) <= a;
    layer0_outputs(7686) <= a xor b;
    layer0_outputs(7687) <= not b or a;
    layer0_outputs(7688) <= not a;
    layer0_outputs(7689) <= not (a xor b);
    layer0_outputs(7690) <= a or b;
    layer0_outputs(7691) <= b;
    layer0_outputs(7692) <= a or b;
    layer0_outputs(7693) <= a;
    layer0_outputs(7694) <= not (a and b);
    layer0_outputs(7695) <= b and not a;
    layer0_outputs(7696) <= not (a xor b);
    layer0_outputs(7697) <= 1'b0;
    layer0_outputs(7698) <= not (a xor b);
    layer0_outputs(7699) <= 1'b0;
    layer0_outputs(7700) <= a and b;
    layer0_outputs(7701) <= not a or b;
    layer0_outputs(7702) <= not (a xor b);
    layer0_outputs(7703) <= b;
    layer0_outputs(7704) <= a or b;
    layer0_outputs(7705) <= not b or a;
    layer0_outputs(7706) <= not a;
    layer0_outputs(7707) <= not a;
    layer0_outputs(7708) <= 1'b1;
    layer0_outputs(7709) <= a or b;
    layer0_outputs(7710) <= not (a or b);
    layer0_outputs(7711) <= not (a or b);
    layer0_outputs(7712) <= not a or b;
    layer0_outputs(7713) <= a;
    layer0_outputs(7714) <= not b;
    layer0_outputs(7715) <= not (a or b);
    layer0_outputs(7716) <= not b;
    layer0_outputs(7717) <= a xor b;
    layer0_outputs(7718) <= b;
    layer0_outputs(7719) <= 1'b0;
    layer0_outputs(7720) <= a and not b;
    layer0_outputs(7721) <= not a;
    layer0_outputs(7722) <= a and not b;
    layer0_outputs(7723) <= not a or b;
    layer0_outputs(7724) <= not a or b;
    layer0_outputs(7725) <= a or b;
    layer0_outputs(7726) <= b;
    layer0_outputs(7727) <= a or b;
    layer0_outputs(7728) <= not (a xor b);
    layer0_outputs(7729) <= a xor b;
    layer0_outputs(7730) <= a xor b;
    layer0_outputs(7731) <= not a or b;
    layer0_outputs(7732) <= a xor b;
    layer0_outputs(7733) <= a;
    layer0_outputs(7734) <= not (a or b);
    layer0_outputs(7735) <= not (a or b);
    layer0_outputs(7736) <= a xor b;
    layer0_outputs(7737) <= not (a or b);
    layer0_outputs(7738) <= not (a xor b);
    layer0_outputs(7739) <= not (a xor b);
    layer0_outputs(7740) <= a and b;
    layer0_outputs(7741) <= a xor b;
    layer0_outputs(7742) <= not b or a;
    layer0_outputs(7743) <= a xor b;
    layer0_outputs(7744) <= a and not b;
    layer0_outputs(7745) <= 1'b1;
    layer0_outputs(7746) <= a or b;
    layer0_outputs(7747) <= not a or b;
    layer0_outputs(7748) <= b;
    layer0_outputs(7749) <= a or b;
    layer0_outputs(7750) <= not b;
    layer0_outputs(7751) <= a xor b;
    layer0_outputs(7752) <= a xor b;
    layer0_outputs(7753) <= not (a or b);
    layer0_outputs(7754) <= not a;
    layer0_outputs(7755) <= not (a or b);
    layer0_outputs(7756) <= not b or a;
    layer0_outputs(7757) <= a or b;
    layer0_outputs(7758) <= b;
    layer0_outputs(7759) <= not (a and b);
    layer0_outputs(7760) <= not (a or b);
    layer0_outputs(7761) <= not b or a;
    layer0_outputs(7762) <= not (a and b);
    layer0_outputs(7763) <= b;
    layer0_outputs(7764) <= not a or b;
    layer0_outputs(7765) <= a and b;
    layer0_outputs(7766) <= not a or b;
    layer0_outputs(7767) <= not a;
    layer0_outputs(7768) <= not (a or b);
    layer0_outputs(7769) <= a or b;
    layer0_outputs(7770) <= b;
    layer0_outputs(7771) <= 1'b1;
    layer0_outputs(7772) <= not b or a;
    layer0_outputs(7773) <= not (a or b);
    layer0_outputs(7774) <= a or b;
    layer0_outputs(7775) <= not a;
    layer0_outputs(7776) <= b and not a;
    layer0_outputs(7777) <= b and not a;
    layer0_outputs(7778) <= b and not a;
    layer0_outputs(7779) <= b and not a;
    layer0_outputs(7780) <= 1'b1;
    layer0_outputs(7781) <= not (a or b);
    layer0_outputs(7782) <= b and not a;
    layer0_outputs(7783) <= not (a xor b);
    layer0_outputs(7784) <= 1'b1;
    layer0_outputs(7785) <= not (a and b);
    layer0_outputs(7786) <= a;
    layer0_outputs(7787) <= a xor b;
    layer0_outputs(7788) <= a;
    layer0_outputs(7789) <= not b or a;
    layer0_outputs(7790) <= a and b;
    layer0_outputs(7791) <= b;
    layer0_outputs(7792) <= a;
    layer0_outputs(7793) <= not b;
    layer0_outputs(7794) <= b and not a;
    layer0_outputs(7795) <= not (a and b);
    layer0_outputs(7796) <= a and not b;
    layer0_outputs(7797) <= a or b;
    layer0_outputs(7798) <= a;
    layer0_outputs(7799) <= a;
    layer0_outputs(7800) <= 1'b0;
    layer0_outputs(7801) <= not (a or b);
    layer0_outputs(7802) <= not a;
    layer0_outputs(7803) <= not a or b;
    layer0_outputs(7804) <= not (a or b);
    layer0_outputs(7805) <= a and not b;
    layer0_outputs(7806) <= not b or a;
    layer0_outputs(7807) <= not a or b;
    layer0_outputs(7808) <= b;
    layer0_outputs(7809) <= a and b;
    layer0_outputs(7810) <= a;
    layer0_outputs(7811) <= not b or a;
    layer0_outputs(7812) <= b;
    layer0_outputs(7813) <= not (a or b);
    layer0_outputs(7814) <= not b or a;
    layer0_outputs(7815) <= a or b;
    layer0_outputs(7816) <= b;
    layer0_outputs(7817) <= a or b;
    layer0_outputs(7818) <= not b;
    layer0_outputs(7819) <= not a;
    layer0_outputs(7820) <= not a;
    layer0_outputs(7821) <= a;
    layer0_outputs(7822) <= b;
    layer0_outputs(7823) <= a or b;
    layer0_outputs(7824) <= a or b;
    layer0_outputs(7825) <= not (a xor b);
    layer0_outputs(7826) <= a xor b;
    layer0_outputs(7827) <= not a or b;
    layer0_outputs(7828) <= not (a or b);
    layer0_outputs(7829) <= not b;
    layer0_outputs(7830) <= not (a or b);
    layer0_outputs(7831) <= a xor b;
    layer0_outputs(7832) <= b;
    layer0_outputs(7833) <= a xor b;
    layer0_outputs(7834) <= not (a or b);
    layer0_outputs(7835) <= not (a and b);
    layer0_outputs(7836) <= a xor b;
    layer0_outputs(7837) <= a or b;
    layer0_outputs(7838) <= b;
    layer0_outputs(7839) <= a or b;
    layer0_outputs(7840) <= not b;
    layer0_outputs(7841) <= b;
    layer0_outputs(7842) <= a or b;
    layer0_outputs(7843) <= 1'b1;
    layer0_outputs(7844) <= not (a and b);
    layer0_outputs(7845) <= a or b;
    layer0_outputs(7846) <= a xor b;
    layer0_outputs(7847) <= b;
    layer0_outputs(7848) <= not (a and b);
    layer0_outputs(7849) <= not (a xor b);
    layer0_outputs(7850) <= a or b;
    layer0_outputs(7851) <= a or b;
    layer0_outputs(7852) <= 1'b1;
    layer0_outputs(7853) <= b and not a;
    layer0_outputs(7854) <= a;
    layer0_outputs(7855) <= a;
    layer0_outputs(7856) <= a;
    layer0_outputs(7857) <= a and not b;
    layer0_outputs(7858) <= a;
    layer0_outputs(7859) <= a or b;
    layer0_outputs(7860) <= a or b;
    layer0_outputs(7861) <= a xor b;
    layer0_outputs(7862) <= a and b;
    layer0_outputs(7863) <= not (a or b);
    layer0_outputs(7864) <= not a;
    layer0_outputs(7865) <= a xor b;
    layer0_outputs(7866) <= a xor b;
    layer0_outputs(7867) <= not (a or b);
    layer0_outputs(7868) <= not (a or b);
    layer0_outputs(7869) <= not (a xor b);
    layer0_outputs(7870) <= b and not a;
    layer0_outputs(7871) <= a or b;
    layer0_outputs(7872) <= a and b;
    layer0_outputs(7873) <= a and not b;
    layer0_outputs(7874) <= a and not b;
    layer0_outputs(7875) <= not (a and b);
    layer0_outputs(7876) <= a;
    layer0_outputs(7877) <= b and not a;
    layer0_outputs(7878) <= not b or a;
    layer0_outputs(7879) <= b;
    layer0_outputs(7880) <= not (a or b);
    layer0_outputs(7881) <= b;
    layer0_outputs(7882) <= a or b;
    layer0_outputs(7883) <= b;
    layer0_outputs(7884) <= 1'b1;
    layer0_outputs(7885) <= not (a or b);
    layer0_outputs(7886) <= 1'b1;
    layer0_outputs(7887) <= not (a xor b);
    layer0_outputs(7888) <= not b or a;
    layer0_outputs(7889) <= a;
    layer0_outputs(7890) <= not a or b;
    layer0_outputs(7891) <= not b or a;
    layer0_outputs(7892) <= a and b;
    layer0_outputs(7893) <= a and not b;
    layer0_outputs(7894) <= b;
    layer0_outputs(7895) <= not (a xor b);
    layer0_outputs(7896) <= a and b;
    layer0_outputs(7897) <= a;
    layer0_outputs(7898) <= b;
    layer0_outputs(7899) <= not (a or b);
    layer0_outputs(7900) <= b and not a;
    layer0_outputs(7901) <= not a;
    layer0_outputs(7902) <= a and not b;
    layer0_outputs(7903) <= b and not a;
    layer0_outputs(7904) <= a xor b;
    layer0_outputs(7905) <= a;
    layer0_outputs(7906) <= a xor b;
    layer0_outputs(7907) <= b and not a;
    layer0_outputs(7908) <= a xor b;
    layer0_outputs(7909) <= a or b;
    layer0_outputs(7910) <= a and not b;
    layer0_outputs(7911) <= a and b;
    layer0_outputs(7912) <= not (a and b);
    layer0_outputs(7913) <= not (a or b);
    layer0_outputs(7914) <= not b;
    layer0_outputs(7915) <= a and not b;
    layer0_outputs(7916) <= not (a or b);
    layer0_outputs(7917) <= not b;
    layer0_outputs(7918) <= a or b;
    layer0_outputs(7919) <= not b or a;
    layer0_outputs(7920) <= not (a or b);
    layer0_outputs(7921) <= not a or b;
    layer0_outputs(7922) <= a and not b;
    layer0_outputs(7923) <= a xor b;
    layer0_outputs(7924) <= a and not b;
    layer0_outputs(7925) <= not (a or b);
    layer0_outputs(7926) <= not a;
    layer0_outputs(7927) <= a or b;
    layer0_outputs(7928) <= not b or a;
    layer0_outputs(7929) <= a or b;
    layer0_outputs(7930) <= 1'b1;
    layer0_outputs(7931) <= not (a and b);
    layer0_outputs(7932) <= 1'b0;
    layer0_outputs(7933) <= a xor b;
    layer0_outputs(7934) <= not b;
    layer0_outputs(7935) <= not (a or b);
    layer0_outputs(7936) <= a;
    layer0_outputs(7937) <= not (a or b);
    layer0_outputs(7938) <= a or b;
    layer0_outputs(7939) <= b and not a;
    layer0_outputs(7940) <= not b or a;
    layer0_outputs(7941) <= b and not a;
    layer0_outputs(7942) <= b and not a;
    layer0_outputs(7943) <= b;
    layer0_outputs(7944) <= 1'b1;
    layer0_outputs(7945) <= b;
    layer0_outputs(7946) <= b;
    layer0_outputs(7947) <= not b or a;
    layer0_outputs(7948) <= not (a xor b);
    layer0_outputs(7949) <= a or b;
    layer0_outputs(7950) <= not b;
    layer0_outputs(7951) <= b and not a;
    layer0_outputs(7952) <= not (a or b);
    layer0_outputs(7953) <= 1'b1;
    layer0_outputs(7954) <= not a;
    layer0_outputs(7955) <= a and not b;
    layer0_outputs(7956) <= not b;
    layer0_outputs(7957) <= not (a or b);
    layer0_outputs(7958) <= not b or a;
    layer0_outputs(7959) <= a xor b;
    layer0_outputs(7960) <= a xor b;
    layer0_outputs(7961) <= b;
    layer0_outputs(7962) <= a and b;
    layer0_outputs(7963) <= not a;
    layer0_outputs(7964) <= not (a and b);
    layer0_outputs(7965) <= not a or b;
    layer0_outputs(7966) <= not (a xor b);
    layer0_outputs(7967) <= not (a or b);
    layer0_outputs(7968) <= not b;
    layer0_outputs(7969) <= a;
    layer0_outputs(7970) <= not (a or b);
    layer0_outputs(7971) <= a or b;
    layer0_outputs(7972) <= not b or a;
    layer0_outputs(7973) <= a;
    layer0_outputs(7974) <= not b or a;
    layer0_outputs(7975) <= a or b;
    layer0_outputs(7976) <= b;
    layer0_outputs(7977) <= not (a xor b);
    layer0_outputs(7978) <= not a;
    layer0_outputs(7979) <= not (a xor b);
    layer0_outputs(7980) <= not b;
    layer0_outputs(7981) <= not (a or b);
    layer0_outputs(7982) <= not (a or b);
    layer0_outputs(7983) <= not (a and b);
    layer0_outputs(7984) <= not (a xor b);
    layer0_outputs(7985) <= a or b;
    layer0_outputs(7986) <= a or b;
    layer0_outputs(7987) <= b and not a;
    layer0_outputs(7988) <= 1'b0;
    layer0_outputs(7989) <= not b or a;
    layer0_outputs(7990) <= a or b;
    layer0_outputs(7991) <= not b or a;
    layer0_outputs(7992) <= not (a or b);
    layer0_outputs(7993) <= 1'b0;
    layer0_outputs(7994) <= not (a xor b);
    layer0_outputs(7995) <= a and not b;
    layer0_outputs(7996) <= a and not b;
    layer0_outputs(7997) <= not a;
    layer0_outputs(7998) <= b;
    layer0_outputs(7999) <= not (a and b);
    layer0_outputs(8000) <= not (a or b);
    layer0_outputs(8001) <= not (a or b);
    layer0_outputs(8002) <= not b or a;
    layer0_outputs(8003) <= a xor b;
    layer0_outputs(8004) <= not (a xor b);
    layer0_outputs(8005) <= not b or a;
    layer0_outputs(8006) <= a;
    layer0_outputs(8007) <= a;
    layer0_outputs(8008) <= not (a xor b);
    layer0_outputs(8009) <= a or b;
    layer0_outputs(8010) <= a xor b;
    layer0_outputs(8011) <= not (a or b);
    layer0_outputs(8012) <= not (a or b);
    layer0_outputs(8013) <= not b or a;
    layer0_outputs(8014) <= not b or a;
    layer0_outputs(8015) <= a xor b;
    layer0_outputs(8016) <= not (a or b);
    layer0_outputs(8017) <= not (a or b);
    layer0_outputs(8018) <= a;
    layer0_outputs(8019) <= not b;
    layer0_outputs(8020) <= not (a and b);
    layer0_outputs(8021) <= not b;
    layer0_outputs(8022) <= a and b;
    layer0_outputs(8023) <= not a or b;
    layer0_outputs(8024) <= b;
    layer0_outputs(8025) <= 1'b0;
    layer0_outputs(8026) <= b and not a;
    layer0_outputs(8027) <= not b;
    layer0_outputs(8028) <= b and not a;
    layer0_outputs(8029) <= a xor b;
    layer0_outputs(8030) <= a;
    layer0_outputs(8031) <= a or b;
    layer0_outputs(8032) <= not b or a;
    layer0_outputs(8033) <= a xor b;
    layer0_outputs(8034) <= a or b;
    layer0_outputs(8035) <= a and not b;
    layer0_outputs(8036) <= a or b;
    layer0_outputs(8037) <= not (a or b);
    layer0_outputs(8038) <= 1'b0;
    layer0_outputs(8039) <= a xor b;
    layer0_outputs(8040) <= b and not a;
    layer0_outputs(8041) <= b;
    layer0_outputs(8042) <= not (a and b);
    layer0_outputs(8043) <= a xor b;
    layer0_outputs(8044) <= not a or b;
    layer0_outputs(8045) <= b;
    layer0_outputs(8046) <= a;
    layer0_outputs(8047) <= not (a or b);
    layer0_outputs(8048) <= not (a xor b);
    layer0_outputs(8049) <= not (a or b);
    layer0_outputs(8050) <= not (a xor b);
    layer0_outputs(8051) <= not a;
    layer0_outputs(8052) <= a xor b;
    layer0_outputs(8053) <= not a or b;
    layer0_outputs(8054) <= not (a or b);
    layer0_outputs(8055) <= not (a or b);
    layer0_outputs(8056) <= not b or a;
    layer0_outputs(8057) <= a;
    layer0_outputs(8058) <= a xor b;
    layer0_outputs(8059) <= not a;
    layer0_outputs(8060) <= a xor b;
    layer0_outputs(8061) <= a xor b;
    layer0_outputs(8062) <= not b;
    layer0_outputs(8063) <= not (a or b);
    layer0_outputs(8064) <= not (a xor b);
    layer0_outputs(8065) <= b and not a;
    layer0_outputs(8066) <= not (a xor b);
    layer0_outputs(8067) <= a;
    layer0_outputs(8068) <= not a or b;
    layer0_outputs(8069) <= not (a or b);
    layer0_outputs(8070) <= not b;
    layer0_outputs(8071) <= not (a or b);
    layer0_outputs(8072) <= not a;
    layer0_outputs(8073) <= not a;
    layer0_outputs(8074) <= not b or a;
    layer0_outputs(8075) <= not (a xor b);
    layer0_outputs(8076) <= 1'b1;
    layer0_outputs(8077) <= not (a or b);
    layer0_outputs(8078) <= not a or b;
    layer0_outputs(8079) <= b and not a;
    layer0_outputs(8080) <= a xor b;
    layer0_outputs(8081) <= a;
    layer0_outputs(8082) <= a;
    layer0_outputs(8083) <= a xor b;
    layer0_outputs(8084) <= not (a and b);
    layer0_outputs(8085) <= not a;
    layer0_outputs(8086) <= not (a xor b);
    layer0_outputs(8087) <= not b;
    layer0_outputs(8088) <= not a;
    layer0_outputs(8089) <= not a or b;
    layer0_outputs(8090) <= a and not b;
    layer0_outputs(8091) <= a;
    layer0_outputs(8092) <= b;
    layer0_outputs(8093) <= not b or a;
    layer0_outputs(8094) <= a xor b;
    layer0_outputs(8095) <= a or b;
    layer0_outputs(8096) <= a and b;
    layer0_outputs(8097) <= not (a or b);
    layer0_outputs(8098) <= not (a or b);
    layer0_outputs(8099) <= not (a or b);
    layer0_outputs(8100) <= a and b;
    layer0_outputs(8101) <= a xor b;
    layer0_outputs(8102) <= not (a or b);
    layer0_outputs(8103) <= a and not b;
    layer0_outputs(8104) <= not (a or b);
    layer0_outputs(8105) <= not (a or b);
    layer0_outputs(8106) <= not b;
    layer0_outputs(8107) <= not a or b;
    layer0_outputs(8108) <= a and b;
    layer0_outputs(8109) <= b and not a;
    layer0_outputs(8110) <= b;
    layer0_outputs(8111) <= not a or b;
    layer0_outputs(8112) <= not a or b;
    layer0_outputs(8113) <= a;
    layer0_outputs(8114) <= a and not b;
    layer0_outputs(8115) <= not a or b;
    layer0_outputs(8116) <= a and b;
    layer0_outputs(8117) <= a;
    layer0_outputs(8118) <= a;
    layer0_outputs(8119) <= not b;
    layer0_outputs(8120) <= a;
    layer0_outputs(8121) <= a and not b;
    layer0_outputs(8122) <= a xor b;
    layer0_outputs(8123) <= a;
    layer0_outputs(8124) <= a and not b;
    layer0_outputs(8125) <= not b or a;
    layer0_outputs(8126) <= a or b;
    layer0_outputs(8127) <= 1'b0;
    layer0_outputs(8128) <= not a or b;
    layer0_outputs(8129) <= 1'b1;
    layer0_outputs(8130) <= not b or a;
    layer0_outputs(8131) <= not (a xor b);
    layer0_outputs(8132) <= a or b;
    layer0_outputs(8133) <= a or b;
    layer0_outputs(8134) <= b and not a;
    layer0_outputs(8135) <= not a or b;
    layer0_outputs(8136) <= not b or a;
    layer0_outputs(8137) <= not a or b;
    layer0_outputs(8138) <= a xor b;
    layer0_outputs(8139) <= not b or a;
    layer0_outputs(8140) <= not (a and b);
    layer0_outputs(8141) <= not (a xor b);
    layer0_outputs(8142) <= not a or b;
    layer0_outputs(8143) <= a and b;
    layer0_outputs(8144) <= b;
    layer0_outputs(8145) <= not (a xor b);
    layer0_outputs(8146) <= b and not a;
    layer0_outputs(8147) <= not a or b;
    layer0_outputs(8148) <= not b or a;
    layer0_outputs(8149) <= not (a or b);
    layer0_outputs(8150) <= not (a or b);
    layer0_outputs(8151) <= a or b;
    layer0_outputs(8152) <= a;
    layer0_outputs(8153) <= 1'b1;
    layer0_outputs(8154) <= not (a or b);
    layer0_outputs(8155) <= not a;
    layer0_outputs(8156) <= a and not b;
    layer0_outputs(8157) <= a or b;
    layer0_outputs(8158) <= b and not a;
    layer0_outputs(8159) <= a or b;
    layer0_outputs(8160) <= a or b;
    layer0_outputs(8161) <= not (a or b);
    layer0_outputs(8162) <= a and not b;
    layer0_outputs(8163) <= not (a xor b);
    layer0_outputs(8164) <= a xor b;
    layer0_outputs(8165) <= not a;
    layer0_outputs(8166) <= b;
    layer0_outputs(8167) <= a;
    layer0_outputs(8168) <= not a;
    layer0_outputs(8169) <= b;
    layer0_outputs(8170) <= a and not b;
    layer0_outputs(8171) <= b;
    layer0_outputs(8172) <= b;
    layer0_outputs(8173) <= b and not a;
    layer0_outputs(8174) <= a xor b;
    layer0_outputs(8175) <= not (a or b);
    layer0_outputs(8176) <= not (a or b);
    layer0_outputs(8177) <= not (a or b);
    layer0_outputs(8178) <= a and not b;
    layer0_outputs(8179) <= not b;
    layer0_outputs(8180) <= a xor b;
    layer0_outputs(8181) <= b;
    layer0_outputs(8182) <= not (a and b);
    layer0_outputs(8183) <= a xor b;
    layer0_outputs(8184) <= not a;
    layer0_outputs(8185) <= not b;
    layer0_outputs(8186) <= not a;
    layer0_outputs(8187) <= not (a xor b);
    layer0_outputs(8188) <= a;
    layer0_outputs(8189) <= not a or b;
    layer0_outputs(8190) <= b;
    layer0_outputs(8191) <= not (a or b);
    layer0_outputs(8192) <= not a;
    layer0_outputs(8193) <= a or b;
    layer0_outputs(8194) <= not (a xor b);
    layer0_outputs(8195) <= a and not b;
    layer0_outputs(8196) <= b and not a;
    layer0_outputs(8197) <= not (a and b);
    layer0_outputs(8198) <= a xor b;
    layer0_outputs(8199) <= b;
    layer0_outputs(8200) <= a or b;
    layer0_outputs(8201) <= not b;
    layer0_outputs(8202) <= 1'b1;
    layer0_outputs(8203) <= a;
    layer0_outputs(8204) <= not (a xor b);
    layer0_outputs(8205) <= not b or a;
    layer0_outputs(8206) <= not (a xor b);
    layer0_outputs(8207) <= not (a xor b);
    layer0_outputs(8208) <= not (a xor b);
    layer0_outputs(8209) <= a xor b;
    layer0_outputs(8210) <= a and b;
    layer0_outputs(8211) <= 1'b1;
    layer0_outputs(8212) <= a and not b;
    layer0_outputs(8213) <= b;
    layer0_outputs(8214) <= b;
    layer0_outputs(8215) <= not b or a;
    layer0_outputs(8216) <= a;
    layer0_outputs(8217) <= a;
    layer0_outputs(8218) <= a and not b;
    layer0_outputs(8219) <= not a;
    layer0_outputs(8220) <= not (a or b);
    layer0_outputs(8221) <= 1'b1;
    layer0_outputs(8222) <= 1'b0;
    layer0_outputs(8223) <= b and not a;
    layer0_outputs(8224) <= not b;
    layer0_outputs(8225) <= 1'b1;
    layer0_outputs(8226) <= not a;
    layer0_outputs(8227) <= b and not a;
    layer0_outputs(8228) <= not (a xor b);
    layer0_outputs(8229) <= a xor b;
    layer0_outputs(8230) <= not a;
    layer0_outputs(8231) <= a;
    layer0_outputs(8232) <= a xor b;
    layer0_outputs(8233) <= a xor b;
    layer0_outputs(8234) <= a and not b;
    layer0_outputs(8235) <= b;
    layer0_outputs(8236) <= a and not b;
    layer0_outputs(8237) <= a or b;
    layer0_outputs(8238) <= not (a or b);
    layer0_outputs(8239) <= not a or b;
    layer0_outputs(8240) <= a;
    layer0_outputs(8241) <= not b;
    layer0_outputs(8242) <= a and not b;
    layer0_outputs(8243) <= not (a or b);
    layer0_outputs(8244) <= a and not b;
    layer0_outputs(8245) <= b and not a;
    layer0_outputs(8246) <= not a or b;
    layer0_outputs(8247) <= not (a or b);
    layer0_outputs(8248) <= not (a or b);
    layer0_outputs(8249) <= not (a or b);
    layer0_outputs(8250) <= b and not a;
    layer0_outputs(8251) <= a xor b;
    layer0_outputs(8252) <= a and not b;
    layer0_outputs(8253) <= not b or a;
    layer0_outputs(8254) <= not (a or b);
    layer0_outputs(8255) <= not b;
    layer0_outputs(8256) <= 1'b1;
    layer0_outputs(8257) <= b;
    layer0_outputs(8258) <= 1'b1;
    layer0_outputs(8259) <= not a;
    layer0_outputs(8260) <= a xor b;
    layer0_outputs(8261) <= not (a or b);
    layer0_outputs(8262) <= not (a and b);
    layer0_outputs(8263) <= not (a xor b);
    layer0_outputs(8264) <= a or b;
    layer0_outputs(8265) <= a;
    layer0_outputs(8266) <= not a;
    layer0_outputs(8267) <= a or b;
    layer0_outputs(8268) <= not (a or b);
    layer0_outputs(8269) <= a or b;
    layer0_outputs(8270) <= not a or b;
    layer0_outputs(8271) <= a or b;
    layer0_outputs(8272) <= a and b;
    layer0_outputs(8273) <= b;
    layer0_outputs(8274) <= not b;
    layer0_outputs(8275) <= not (a or b);
    layer0_outputs(8276) <= 1'b1;
    layer0_outputs(8277) <= not a;
    layer0_outputs(8278) <= a;
    layer0_outputs(8279) <= not (a or b);
    layer0_outputs(8280) <= a xor b;
    layer0_outputs(8281) <= not a;
    layer0_outputs(8282) <= not a;
    layer0_outputs(8283) <= b and not a;
    layer0_outputs(8284) <= a or b;
    layer0_outputs(8285) <= 1'b0;
    layer0_outputs(8286) <= not a;
    layer0_outputs(8287) <= 1'b0;
    layer0_outputs(8288) <= a;
    layer0_outputs(8289) <= not a;
    layer0_outputs(8290) <= not (a xor b);
    layer0_outputs(8291) <= not b or a;
    layer0_outputs(8292) <= b and not a;
    layer0_outputs(8293) <= a and b;
    layer0_outputs(8294) <= not b;
    layer0_outputs(8295) <= b and not a;
    layer0_outputs(8296) <= 1'b1;
    layer0_outputs(8297) <= not b or a;
    layer0_outputs(8298) <= not (a or b);
    layer0_outputs(8299) <= 1'b1;
    layer0_outputs(8300) <= a or b;
    layer0_outputs(8301) <= a xor b;
    layer0_outputs(8302) <= not a;
    layer0_outputs(8303) <= a or b;
    layer0_outputs(8304) <= not b or a;
    layer0_outputs(8305) <= not b;
    layer0_outputs(8306) <= a or b;
    layer0_outputs(8307) <= not a or b;
    layer0_outputs(8308) <= 1'b1;
    layer0_outputs(8309) <= a or b;
    layer0_outputs(8310) <= a and not b;
    layer0_outputs(8311) <= a and b;
    layer0_outputs(8312) <= a or b;
    layer0_outputs(8313) <= not a;
    layer0_outputs(8314) <= not (a or b);
    layer0_outputs(8315) <= 1'b1;
    layer0_outputs(8316) <= not b;
    layer0_outputs(8317) <= a xor b;
    layer0_outputs(8318) <= not b;
    layer0_outputs(8319) <= not (a xor b);
    layer0_outputs(8320) <= not (a xor b);
    layer0_outputs(8321) <= not b;
    layer0_outputs(8322) <= not (a or b);
    layer0_outputs(8323) <= 1'b1;
    layer0_outputs(8324) <= not (a xor b);
    layer0_outputs(8325) <= b;
    layer0_outputs(8326) <= not (a or b);
    layer0_outputs(8327) <= not (a xor b);
    layer0_outputs(8328) <= b and not a;
    layer0_outputs(8329) <= not a;
    layer0_outputs(8330) <= a or b;
    layer0_outputs(8331) <= not (a xor b);
    layer0_outputs(8332) <= not (a or b);
    layer0_outputs(8333) <= not a;
    layer0_outputs(8334) <= b and not a;
    layer0_outputs(8335) <= b;
    layer0_outputs(8336) <= not (a or b);
    layer0_outputs(8337) <= a;
    layer0_outputs(8338) <= a xor b;
    layer0_outputs(8339) <= a and not b;
    layer0_outputs(8340) <= a xor b;
    layer0_outputs(8341) <= b;
    layer0_outputs(8342) <= not a or b;
    layer0_outputs(8343) <= not b;
    layer0_outputs(8344) <= not (a or b);
    layer0_outputs(8345) <= not (a and b);
    layer0_outputs(8346) <= b and not a;
    layer0_outputs(8347) <= not (a and b);
    layer0_outputs(8348) <= a xor b;
    layer0_outputs(8349) <= a and not b;
    layer0_outputs(8350) <= a or b;
    layer0_outputs(8351) <= b and not a;
    layer0_outputs(8352) <= b;
    layer0_outputs(8353) <= b and not a;
    layer0_outputs(8354) <= not (a or b);
    layer0_outputs(8355) <= a or b;
    layer0_outputs(8356) <= not b;
    layer0_outputs(8357) <= b;
    layer0_outputs(8358) <= a;
    layer0_outputs(8359) <= a and not b;
    layer0_outputs(8360) <= a and b;
    layer0_outputs(8361) <= b and not a;
    layer0_outputs(8362) <= a or b;
    layer0_outputs(8363) <= 1'b0;
    layer0_outputs(8364) <= a or b;
    layer0_outputs(8365) <= not (a and b);
    layer0_outputs(8366) <= b and not a;
    layer0_outputs(8367) <= a;
    layer0_outputs(8368) <= not b or a;
    layer0_outputs(8369) <= not (a or b);
    layer0_outputs(8370) <= a;
    layer0_outputs(8371) <= not b or a;
    layer0_outputs(8372) <= not b;
    layer0_outputs(8373) <= a;
    layer0_outputs(8374) <= a and not b;
    layer0_outputs(8375) <= a xor b;
    layer0_outputs(8376) <= not b;
    layer0_outputs(8377) <= not (a or b);
    layer0_outputs(8378) <= not (a or b);
    layer0_outputs(8379) <= a or b;
    layer0_outputs(8380) <= not a or b;
    layer0_outputs(8381) <= not b;
    layer0_outputs(8382) <= not (a or b);
    layer0_outputs(8383) <= a xor b;
    layer0_outputs(8384) <= not (a and b);
    layer0_outputs(8385) <= not (a xor b);
    layer0_outputs(8386) <= not b;
    layer0_outputs(8387) <= not (a xor b);
    layer0_outputs(8388) <= not (a or b);
    layer0_outputs(8389) <= not a;
    layer0_outputs(8390) <= a xor b;
    layer0_outputs(8391) <= not (a and b);
    layer0_outputs(8392) <= b;
    layer0_outputs(8393) <= not (a or b);
    layer0_outputs(8394) <= not a or b;
    layer0_outputs(8395) <= not (a or b);
    layer0_outputs(8396) <= not (a or b);
    layer0_outputs(8397) <= not a or b;
    layer0_outputs(8398) <= 1'b1;
    layer0_outputs(8399) <= 1'b0;
    layer0_outputs(8400) <= not b or a;
    layer0_outputs(8401) <= a;
    layer0_outputs(8402) <= a and b;
    layer0_outputs(8403) <= a and not b;
    layer0_outputs(8404) <= a or b;
    layer0_outputs(8405) <= not (a xor b);
    layer0_outputs(8406) <= b and not a;
    layer0_outputs(8407) <= a and not b;
    layer0_outputs(8408) <= not (a xor b);
    layer0_outputs(8409) <= not (a xor b);
    layer0_outputs(8410) <= a and not b;
    layer0_outputs(8411) <= not b;
    layer0_outputs(8412) <= not (a and b);
    layer0_outputs(8413) <= a xor b;
    layer0_outputs(8414) <= 1'b1;
    layer0_outputs(8415) <= not a;
    layer0_outputs(8416) <= a or b;
    layer0_outputs(8417) <= not (a or b);
    layer0_outputs(8418) <= not (a xor b);
    layer0_outputs(8419) <= not (a or b);
    layer0_outputs(8420) <= not a or b;
    layer0_outputs(8421) <= a xor b;
    layer0_outputs(8422) <= 1'b0;
    layer0_outputs(8423) <= not (a xor b);
    layer0_outputs(8424) <= not b or a;
    layer0_outputs(8425) <= a;
    layer0_outputs(8426) <= not a or b;
    layer0_outputs(8427) <= not b;
    layer0_outputs(8428) <= not (a xor b);
    layer0_outputs(8429) <= not a;
    layer0_outputs(8430) <= a and not b;
    layer0_outputs(8431) <= a and b;
    layer0_outputs(8432) <= a and not b;
    layer0_outputs(8433) <= not (a and b);
    layer0_outputs(8434) <= not b or a;
    layer0_outputs(8435) <= a xor b;
    layer0_outputs(8436) <= not b;
    layer0_outputs(8437) <= b and not a;
    layer0_outputs(8438) <= not b or a;
    layer0_outputs(8439) <= not a or b;
    layer0_outputs(8440) <= not (a or b);
    layer0_outputs(8441) <= not a;
    layer0_outputs(8442) <= not a;
    layer0_outputs(8443) <= not a;
    layer0_outputs(8444) <= b and not a;
    layer0_outputs(8445) <= not (a xor b);
    layer0_outputs(8446) <= a xor b;
    layer0_outputs(8447) <= a and not b;
    layer0_outputs(8448) <= not b;
    layer0_outputs(8449) <= not a;
    layer0_outputs(8450) <= a xor b;
    layer0_outputs(8451) <= not (a or b);
    layer0_outputs(8452) <= a;
    layer0_outputs(8453) <= a or b;
    layer0_outputs(8454) <= not (a or b);
    layer0_outputs(8455) <= not a or b;
    layer0_outputs(8456) <= a or b;
    layer0_outputs(8457) <= a or b;
    layer0_outputs(8458) <= a or b;
    layer0_outputs(8459) <= b and not a;
    layer0_outputs(8460) <= not (a xor b);
    layer0_outputs(8461) <= not (a or b);
    layer0_outputs(8462) <= a or b;
    layer0_outputs(8463) <= a;
    layer0_outputs(8464) <= 1'b0;
    layer0_outputs(8465) <= not (a and b);
    layer0_outputs(8466) <= not (a or b);
    layer0_outputs(8467) <= a xor b;
    layer0_outputs(8468) <= a xor b;
    layer0_outputs(8469) <= 1'b1;
    layer0_outputs(8470) <= not (a xor b);
    layer0_outputs(8471) <= not a or b;
    layer0_outputs(8472) <= b;
    layer0_outputs(8473) <= not (a or b);
    layer0_outputs(8474) <= not b or a;
    layer0_outputs(8475) <= not b;
    layer0_outputs(8476) <= 1'b1;
    layer0_outputs(8477) <= a or b;
    layer0_outputs(8478) <= a or b;
    layer0_outputs(8479) <= not b;
    layer0_outputs(8480) <= a or b;
    layer0_outputs(8481) <= not (a xor b);
    layer0_outputs(8482) <= 1'b1;
    layer0_outputs(8483) <= not b;
    layer0_outputs(8484) <= not b;
    layer0_outputs(8485) <= not a;
    layer0_outputs(8486) <= 1'b0;
    layer0_outputs(8487) <= not b or a;
    layer0_outputs(8488) <= b;
    layer0_outputs(8489) <= not a;
    layer0_outputs(8490) <= not (a or b);
    layer0_outputs(8491) <= not (a or b);
    layer0_outputs(8492) <= not b or a;
    layer0_outputs(8493) <= b;
    layer0_outputs(8494) <= not b;
    layer0_outputs(8495) <= not a or b;
    layer0_outputs(8496) <= a or b;
    layer0_outputs(8497) <= not b or a;
    layer0_outputs(8498) <= a;
    layer0_outputs(8499) <= a and b;
    layer0_outputs(8500) <= not a;
    layer0_outputs(8501) <= not a or b;
    layer0_outputs(8502) <= a and not b;
    layer0_outputs(8503) <= a xor b;
    layer0_outputs(8504) <= b and not a;
    layer0_outputs(8505) <= not a or b;
    layer0_outputs(8506) <= not a or b;
    layer0_outputs(8507) <= not b;
    layer0_outputs(8508) <= not (a xor b);
    layer0_outputs(8509) <= a;
    layer0_outputs(8510) <= not a;
    layer0_outputs(8511) <= not b or a;
    layer0_outputs(8512) <= a or b;
    layer0_outputs(8513) <= a or b;
    layer0_outputs(8514) <= a and not b;
    layer0_outputs(8515) <= not (a xor b);
    layer0_outputs(8516) <= not b or a;
    layer0_outputs(8517) <= not (a xor b);
    layer0_outputs(8518) <= a or b;
    layer0_outputs(8519) <= b;
    layer0_outputs(8520) <= not a or b;
    layer0_outputs(8521) <= a xor b;
    layer0_outputs(8522) <= a xor b;
    layer0_outputs(8523) <= not a or b;
    layer0_outputs(8524) <= not (a or b);
    layer0_outputs(8525) <= a and not b;
    layer0_outputs(8526) <= a;
    layer0_outputs(8527) <= b;
    layer0_outputs(8528) <= a or b;
    layer0_outputs(8529) <= a or b;
    layer0_outputs(8530) <= not b;
    layer0_outputs(8531) <= not a or b;
    layer0_outputs(8532) <= a and not b;
    layer0_outputs(8533) <= not (a xor b);
    layer0_outputs(8534) <= b and not a;
    layer0_outputs(8535) <= not b;
    layer0_outputs(8536) <= a and not b;
    layer0_outputs(8537) <= b;
    layer0_outputs(8538) <= not a;
    layer0_outputs(8539) <= not a or b;
    layer0_outputs(8540) <= not (a or b);
    layer0_outputs(8541) <= not (a and b);
    layer0_outputs(8542) <= a xor b;
    layer0_outputs(8543) <= b;
    layer0_outputs(8544) <= not (a xor b);
    layer0_outputs(8545) <= a or b;
    layer0_outputs(8546) <= not (a or b);
    layer0_outputs(8547) <= b and not a;
    layer0_outputs(8548) <= not (a or b);
    layer0_outputs(8549) <= a and not b;
    layer0_outputs(8550) <= not (a xor b);
    layer0_outputs(8551) <= not a;
    layer0_outputs(8552) <= not (a or b);
    layer0_outputs(8553) <= not b or a;
    layer0_outputs(8554) <= 1'b1;
    layer0_outputs(8555) <= b;
    layer0_outputs(8556) <= b;
    layer0_outputs(8557) <= not b;
    layer0_outputs(8558) <= a;
    layer0_outputs(8559) <= a and not b;
    layer0_outputs(8560) <= not (a or b);
    layer0_outputs(8561) <= a xor b;
    layer0_outputs(8562) <= a and not b;
    layer0_outputs(8563) <= b and not a;
    layer0_outputs(8564) <= a and not b;
    layer0_outputs(8565) <= a and not b;
    layer0_outputs(8566) <= not (a xor b);
    layer0_outputs(8567) <= a and b;
    layer0_outputs(8568) <= b and not a;
    layer0_outputs(8569) <= a xor b;
    layer0_outputs(8570) <= a and not b;
    layer0_outputs(8571) <= a and not b;
    layer0_outputs(8572) <= not a or b;
    layer0_outputs(8573) <= a or b;
    layer0_outputs(8574) <= not a;
    layer0_outputs(8575) <= not (a or b);
    layer0_outputs(8576) <= a or b;
    layer0_outputs(8577) <= a and b;
    layer0_outputs(8578) <= not b or a;
    layer0_outputs(8579) <= not (a or b);
    layer0_outputs(8580) <= not a;
    layer0_outputs(8581) <= a or b;
    layer0_outputs(8582) <= a and not b;
    layer0_outputs(8583) <= 1'b0;
    layer0_outputs(8584) <= a and b;
    layer0_outputs(8585) <= not b or a;
    layer0_outputs(8586) <= not b;
    layer0_outputs(8587) <= a or b;
    layer0_outputs(8588) <= a;
    layer0_outputs(8589) <= not (a and b);
    layer0_outputs(8590) <= 1'b0;
    layer0_outputs(8591) <= a xor b;
    layer0_outputs(8592) <= not b;
    layer0_outputs(8593) <= b;
    layer0_outputs(8594) <= a xor b;
    layer0_outputs(8595) <= not a;
    layer0_outputs(8596) <= a xor b;
    layer0_outputs(8597) <= not a;
    layer0_outputs(8598) <= a or b;
    layer0_outputs(8599) <= b and not a;
    layer0_outputs(8600) <= b;
    layer0_outputs(8601) <= a xor b;
    layer0_outputs(8602) <= not a or b;
    layer0_outputs(8603) <= a xor b;
    layer0_outputs(8604) <= b;
    layer0_outputs(8605) <= not (a xor b);
    layer0_outputs(8606) <= not (a and b);
    layer0_outputs(8607) <= b;
    layer0_outputs(8608) <= not (a or b);
    layer0_outputs(8609) <= a or b;
    layer0_outputs(8610) <= a and b;
    layer0_outputs(8611) <= not (a and b);
    layer0_outputs(8612) <= not (a or b);
    layer0_outputs(8613) <= a and not b;
    layer0_outputs(8614) <= not a or b;
    layer0_outputs(8615) <= not (a or b);
    layer0_outputs(8616) <= a or b;
    layer0_outputs(8617) <= a or b;
    layer0_outputs(8618) <= not b;
    layer0_outputs(8619) <= not (a or b);
    layer0_outputs(8620) <= a or b;
    layer0_outputs(8621) <= a or b;
    layer0_outputs(8622) <= b and not a;
    layer0_outputs(8623) <= a or b;
    layer0_outputs(8624) <= a;
    layer0_outputs(8625) <= not (a xor b);
    layer0_outputs(8626) <= b;
    layer0_outputs(8627) <= not a or b;
    layer0_outputs(8628) <= a and not b;
    layer0_outputs(8629) <= not b or a;
    layer0_outputs(8630) <= not (a xor b);
    layer0_outputs(8631) <= not (a or b);
    layer0_outputs(8632) <= a xor b;
    layer0_outputs(8633) <= a and not b;
    layer0_outputs(8634) <= not b;
    layer0_outputs(8635) <= not (a or b);
    layer0_outputs(8636) <= not (a xor b);
    layer0_outputs(8637) <= not b or a;
    layer0_outputs(8638) <= not (a or b);
    layer0_outputs(8639) <= not b;
    layer0_outputs(8640) <= a;
    layer0_outputs(8641) <= b;
    layer0_outputs(8642) <= not b;
    layer0_outputs(8643) <= a;
    layer0_outputs(8644) <= not (a or b);
    layer0_outputs(8645) <= not a or b;
    layer0_outputs(8646) <= not b;
    layer0_outputs(8647) <= not a;
    layer0_outputs(8648) <= not (a or b);
    layer0_outputs(8649) <= a and b;
    layer0_outputs(8650) <= a or b;
    layer0_outputs(8651) <= a and b;
    layer0_outputs(8652) <= b and not a;
    layer0_outputs(8653) <= not (a or b);
    layer0_outputs(8654) <= a xor b;
    layer0_outputs(8655) <= not b or a;
    layer0_outputs(8656) <= not b;
    layer0_outputs(8657) <= a xor b;
    layer0_outputs(8658) <= a or b;
    layer0_outputs(8659) <= not b;
    layer0_outputs(8660) <= not a or b;
    layer0_outputs(8661) <= a and b;
    layer0_outputs(8662) <= 1'b1;
    layer0_outputs(8663) <= not (a or b);
    layer0_outputs(8664) <= not a;
    layer0_outputs(8665) <= a xor b;
    layer0_outputs(8666) <= not (a and b);
    layer0_outputs(8667) <= not a;
    layer0_outputs(8668) <= not (a or b);
    layer0_outputs(8669) <= 1'b1;
    layer0_outputs(8670) <= not b or a;
    layer0_outputs(8671) <= a xor b;
    layer0_outputs(8672) <= a and not b;
    layer0_outputs(8673) <= not (a or b);
    layer0_outputs(8674) <= not b or a;
    layer0_outputs(8675) <= not b or a;
    layer0_outputs(8676) <= b;
    layer0_outputs(8677) <= a or b;
    layer0_outputs(8678) <= not b;
    layer0_outputs(8679) <= a xor b;
    layer0_outputs(8680) <= not (a or b);
    layer0_outputs(8681) <= a and not b;
    layer0_outputs(8682) <= a and not b;
    layer0_outputs(8683) <= a and not b;
    layer0_outputs(8684) <= a or b;
    layer0_outputs(8685) <= not (a xor b);
    layer0_outputs(8686) <= b and not a;
    layer0_outputs(8687) <= not (a or b);
    layer0_outputs(8688) <= a xor b;
    layer0_outputs(8689) <= a and not b;
    layer0_outputs(8690) <= not a;
    layer0_outputs(8691) <= a or b;
    layer0_outputs(8692) <= a and not b;
    layer0_outputs(8693) <= a or b;
    layer0_outputs(8694) <= not a or b;
    layer0_outputs(8695) <= not (a or b);
    layer0_outputs(8696) <= not (a or b);
    layer0_outputs(8697) <= a or b;
    layer0_outputs(8698) <= not a;
    layer0_outputs(8699) <= b;
    layer0_outputs(8700) <= a or b;
    layer0_outputs(8701) <= not (a and b);
    layer0_outputs(8702) <= a xor b;
    layer0_outputs(8703) <= not b;
    layer0_outputs(8704) <= not a;
    layer0_outputs(8705) <= 1'b1;
    layer0_outputs(8706) <= not b or a;
    layer0_outputs(8707) <= b;
    layer0_outputs(8708) <= a and not b;
    layer0_outputs(8709) <= not b;
    layer0_outputs(8710) <= a xor b;
    layer0_outputs(8711) <= b;
    layer0_outputs(8712) <= a or b;
    layer0_outputs(8713) <= b;
    layer0_outputs(8714) <= not a;
    layer0_outputs(8715) <= b and not a;
    layer0_outputs(8716) <= a or b;
    layer0_outputs(8717) <= not (a xor b);
    layer0_outputs(8718) <= b and not a;
    layer0_outputs(8719) <= not (a xor b);
    layer0_outputs(8720) <= a;
    layer0_outputs(8721) <= not b;
    layer0_outputs(8722) <= not (a or b);
    layer0_outputs(8723) <= not b;
    layer0_outputs(8724) <= a or b;
    layer0_outputs(8725) <= not (a xor b);
    layer0_outputs(8726) <= a;
    layer0_outputs(8727) <= b;
    layer0_outputs(8728) <= b and not a;
    layer0_outputs(8729) <= not (a xor b);
    layer0_outputs(8730) <= not a or b;
    layer0_outputs(8731) <= a and not b;
    layer0_outputs(8732) <= a xor b;
    layer0_outputs(8733) <= not b;
    layer0_outputs(8734) <= a or b;
    layer0_outputs(8735) <= b and not a;
    layer0_outputs(8736) <= not b or a;
    layer0_outputs(8737) <= b and not a;
    layer0_outputs(8738) <= a xor b;
    layer0_outputs(8739) <= a xor b;
    layer0_outputs(8740) <= a or b;
    layer0_outputs(8741) <= a;
    layer0_outputs(8742) <= a;
    layer0_outputs(8743) <= not (a or b);
    layer0_outputs(8744) <= not a;
    layer0_outputs(8745) <= a and b;
    layer0_outputs(8746) <= not b or a;
    layer0_outputs(8747) <= a or b;
    layer0_outputs(8748) <= b and not a;
    layer0_outputs(8749) <= not b;
    layer0_outputs(8750) <= not a or b;
    layer0_outputs(8751) <= a and not b;
    layer0_outputs(8752) <= not (a or b);
    layer0_outputs(8753) <= a and not b;
    layer0_outputs(8754) <= a and not b;
    layer0_outputs(8755) <= not (a and b);
    layer0_outputs(8756) <= a xor b;
    layer0_outputs(8757) <= not a or b;
    layer0_outputs(8758) <= not a or b;
    layer0_outputs(8759) <= a;
    layer0_outputs(8760) <= not a;
    layer0_outputs(8761) <= b;
    layer0_outputs(8762) <= a xor b;
    layer0_outputs(8763) <= not a or b;
    layer0_outputs(8764) <= a or b;
    layer0_outputs(8765) <= not b;
    layer0_outputs(8766) <= b;
    layer0_outputs(8767) <= a or b;
    layer0_outputs(8768) <= a and b;
    layer0_outputs(8769) <= 1'b0;
    layer0_outputs(8770) <= not (a xor b);
    layer0_outputs(8771) <= a or b;
    layer0_outputs(8772) <= a or b;
    layer0_outputs(8773) <= b and not a;
    layer0_outputs(8774) <= a and b;
    layer0_outputs(8775) <= b;
    layer0_outputs(8776) <= b and not a;
    layer0_outputs(8777) <= not a;
    layer0_outputs(8778) <= not b or a;
    layer0_outputs(8779) <= not b;
    layer0_outputs(8780) <= a and b;
    layer0_outputs(8781) <= 1'b0;
    layer0_outputs(8782) <= b and not a;
    layer0_outputs(8783) <= not a or b;
    layer0_outputs(8784) <= a or b;
    layer0_outputs(8785) <= not (a xor b);
    layer0_outputs(8786) <= a xor b;
    layer0_outputs(8787) <= a;
    layer0_outputs(8788) <= a or b;
    layer0_outputs(8789) <= a and not b;
    layer0_outputs(8790) <= b and not a;
    layer0_outputs(8791) <= not (a xor b);
    layer0_outputs(8792) <= not (a xor b);
    layer0_outputs(8793) <= not b or a;
    layer0_outputs(8794) <= a xor b;
    layer0_outputs(8795) <= not b;
    layer0_outputs(8796) <= not b or a;
    layer0_outputs(8797) <= not (a or b);
    layer0_outputs(8798) <= 1'b1;
    layer0_outputs(8799) <= a and not b;
    layer0_outputs(8800) <= a xor b;
    layer0_outputs(8801) <= b;
    layer0_outputs(8802) <= not (a xor b);
    layer0_outputs(8803) <= a and not b;
    layer0_outputs(8804) <= not (a or b);
    layer0_outputs(8805) <= not (a or b);
    layer0_outputs(8806) <= not a;
    layer0_outputs(8807) <= not a or b;
    layer0_outputs(8808) <= not (a and b);
    layer0_outputs(8809) <= b;
    layer0_outputs(8810) <= a and not b;
    layer0_outputs(8811) <= not (a or b);
    layer0_outputs(8812) <= not a;
    layer0_outputs(8813) <= a and b;
    layer0_outputs(8814) <= a or b;
    layer0_outputs(8815) <= 1'b1;
    layer0_outputs(8816) <= not a;
    layer0_outputs(8817) <= a or b;
    layer0_outputs(8818) <= a xor b;
    layer0_outputs(8819) <= a and not b;
    layer0_outputs(8820) <= a or b;
    layer0_outputs(8821) <= b;
    layer0_outputs(8822) <= not b;
    layer0_outputs(8823) <= not (a or b);
    layer0_outputs(8824) <= not b;
    layer0_outputs(8825) <= not a;
    layer0_outputs(8826) <= b and not a;
    layer0_outputs(8827) <= not a;
    layer0_outputs(8828) <= not a;
    layer0_outputs(8829) <= not a;
    layer0_outputs(8830) <= a;
    layer0_outputs(8831) <= a xor b;
    layer0_outputs(8832) <= not (a or b);
    layer0_outputs(8833) <= a and not b;
    layer0_outputs(8834) <= a or b;
    layer0_outputs(8835) <= b;
    layer0_outputs(8836) <= a and not b;
    layer0_outputs(8837) <= a xor b;
    layer0_outputs(8838) <= b;
    layer0_outputs(8839) <= a and not b;
    layer0_outputs(8840) <= a or b;
    layer0_outputs(8841) <= b;
    layer0_outputs(8842) <= not b;
    layer0_outputs(8843) <= a or b;
    layer0_outputs(8844) <= not a;
    layer0_outputs(8845) <= not b;
    layer0_outputs(8846) <= a or b;
    layer0_outputs(8847) <= a or b;
    layer0_outputs(8848) <= not (a xor b);
    layer0_outputs(8849) <= not (a and b);
    layer0_outputs(8850) <= not (a or b);
    layer0_outputs(8851) <= a;
    layer0_outputs(8852) <= b and not a;
    layer0_outputs(8853) <= a or b;
    layer0_outputs(8854) <= not a or b;
    layer0_outputs(8855) <= b;
    layer0_outputs(8856) <= a and b;
    layer0_outputs(8857) <= not (a xor b);
    layer0_outputs(8858) <= a or b;
    layer0_outputs(8859) <= b and not a;
    layer0_outputs(8860) <= b;
    layer0_outputs(8861) <= not (a or b);
    layer0_outputs(8862) <= not b;
    layer0_outputs(8863) <= b;
    layer0_outputs(8864) <= not a or b;
    layer0_outputs(8865) <= not b;
    layer0_outputs(8866) <= b and not a;
    layer0_outputs(8867) <= a xor b;
    layer0_outputs(8868) <= a;
    layer0_outputs(8869) <= not a;
    layer0_outputs(8870) <= a;
    layer0_outputs(8871) <= not (a or b);
    layer0_outputs(8872) <= not (a or b);
    layer0_outputs(8873) <= 1'b1;
    layer0_outputs(8874) <= not b;
    layer0_outputs(8875) <= not b;
    layer0_outputs(8876) <= not a or b;
    layer0_outputs(8877) <= not a;
    layer0_outputs(8878) <= a xor b;
    layer0_outputs(8879) <= a and b;
    layer0_outputs(8880) <= not (a xor b);
    layer0_outputs(8881) <= not b or a;
    layer0_outputs(8882) <= not (a xor b);
    layer0_outputs(8883) <= not b;
    layer0_outputs(8884) <= not a;
    layer0_outputs(8885) <= b and not a;
    layer0_outputs(8886) <= b and not a;
    layer0_outputs(8887) <= not a;
    layer0_outputs(8888) <= not b or a;
    layer0_outputs(8889) <= b and not a;
    layer0_outputs(8890) <= b;
    layer0_outputs(8891) <= a or b;
    layer0_outputs(8892) <= not b or a;
    layer0_outputs(8893) <= a and not b;
    layer0_outputs(8894) <= not (a or b);
    layer0_outputs(8895) <= not (a xor b);
    layer0_outputs(8896) <= b;
    layer0_outputs(8897) <= not b or a;
    layer0_outputs(8898) <= b;
    layer0_outputs(8899) <= a or b;
    layer0_outputs(8900) <= a and not b;
    layer0_outputs(8901) <= a xor b;
    layer0_outputs(8902) <= b and not a;
    layer0_outputs(8903) <= not (a or b);
    layer0_outputs(8904) <= not a;
    layer0_outputs(8905) <= not (a or b);
    layer0_outputs(8906) <= not (a or b);
    layer0_outputs(8907) <= not (a or b);
    layer0_outputs(8908) <= not (a xor b);
    layer0_outputs(8909) <= a xor b;
    layer0_outputs(8910) <= not a;
    layer0_outputs(8911) <= not (a and b);
    layer0_outputs(8912) <= not (a xor b);
    layer0_outputs(8913) <= 1'b1;
    layer0_outputs(8914) <= not b;
    layer0_outputs(8915) <= a and not b;
    layer0_outputs(8916) <= a and not b;
    layer0_outputs(8917) <= a;
    layer0_outputs(8918) <= not a;
    layer0_outputs(8919) <= a;
    layer0_outputs(8920) <= not a;
    layer0_outputs(8921) <= not b;
    layer0_outputs(8922) <= not a;
    layer0_outputs(8923) <= not b;
    layer0_outputs(8924) <= not a;
    layer0_outputs(8925) <= not b or a;
    layer0_outputs(8926) <= b and not a;
    layer0_outputs(8927) <= b and not a;
    layer0_outputs(8928) <= b and not a;
    layer0_outputs(8929) <= not a or b;
    layer0_outputs(8930) <= b;
    layer0_outputs(8931) <= a or b;
    layer0_outputs(8932) <= a and not b;
    layer0_outputs(8933) <= a or b;
    layer0_outputs(8934) <= not b or a;
    layer0_outputs(8935) <= not (a or b);
    layer0_outputs(8936) <= 1'b0;
    layer0_outputs(8937) <= a;
    layer0_outputs(8938) <= a xor b;
    layer0_outputs(8939) <= not a or b;
    layer0_outputs(8940) <= a or b;
    layer0_outputs(8941) <= a xor b;
    layer0_outputs(8942) <= a or b;
    layer0_outputs(8943) <= a and b;
    layer0_outputs(8944) <= not (a and b);
    layer0_outputs(8945) <= a and b;
    layer0_outputs(8946) <= not a;
    layer0_outputs(8947) <= a;
    layer0_outputs(8948) <= not (a and b);
    layer0_outputs(8949) <= b;
    layer0_outputs(8950) <= a;
    layer0_outputs(8951) <= a or b;
    layer0_outputs(8952) <= not a;
    layer0_outputs(8953) <= a or b;
    layer0_outputs(8954) <= a;
    layer0_outputs(8955) <= not a;
    layer0_outputs(8956) <= a and b;
    layer0_outputs(8957) <= not (a or b);
    layer0_outputs(8958) <= not (a or b);
    layer0_outputs(8959) <= a and not b;
    layer0_outputs(8960) <= not b or a;
    layer0_outputs(8961) <= a and not b;
    layer0_outputs(8962) <= a;
    layer0_outputs(8963) <= 1'b1;
    layer0_outputs(8964) <= not (a or b);
    layer0_outputs(8965) <= not b or a;
    layer0_outputs(8966) <= a or b;
    layer0_outputs(8967) <= not a;
    layer0_outputs(8968) <= not b or a;
    layer0_outputs(8969) <= not b;
    layer0_outputs(8970) <= not b;
    layer0_outputs(8971) <= not b;
    layer0_outputs(8972) <= a xor b;
    layer0_outputs(8973) <= not a;
    layer0_outputs(8974) <= not (a or b);
    layer0_outputs(8975) <= not (a or b);
    layer0_outputs(8976) <= not (a xor b);
    layer0_outputs(8977) <= not (a xor b);
    layer0_outputs(8978) <= not (a and b);
    layer0_outputs(8979) <= a;
    layer0_outputs(8980) <= b;
    layer0_outputs(8981) <= a or b;
    layer0_outputs(8982) <= a or b;
    layer0_outputs(8983) <= not (a xor b);
    layer0_outputs(8984) <= b;
    layer0_outputs(8985) <= not (a or b);
    layer0_outputs(8986) <= a;
    layer0_outputs(8987) <= a or b;
    layer0_outputs(8988) <= a;
    layer0_outputs(8989) <= b and not a;
    layer0_outputs(8990) <= a and not b;
    layer0_outputs(8991) <= not (a or b);
    layer0_outputs(8992) <= not (a or b);
    layer0_outputs(8993) <= a;
    layer0_outputs(8994) <= not b;
    layer0_outputs(8995) <= a;
    layer0_outputs(8996) <= not b or a;
    layer0_outputs(8997) <= not (a xor b);
    layer0_outputs(8998) <= a or b;
    layer0_outputs(8999) <= a xor b;
    layer0_outputs(9000) <= 1'b0;
    layer0_outputs(9001) <= not a or b;
    layer0_outputs(9002) <= not (a or b);
    layer0_outputs(9003) <= not (a xor b);
    layer0_outputs(9004) <= not (a xor b);
    layer0_outputs(9005) <= a and not b;
    layer0_outputs(9006) <= not a;
    layer0_outputs(9007) <= 1'b1;
    layer0_outputs(9008) <= a;
    layer0_outputs(9009) <= a;
    layer0_outputs(9010) <= a;
    layer0_outputs(9011) <= b;
    layer0_outputs(9012) <= not (a or b);
    layer0_outputs(9013) <= not a;
    layer0_outputs(9014) <= not a or b;
    layer0_outputs(9015) <= 1'b0;
    layer0_outputs(9016) <= b;
    layer0_outputs(9017) <= not (a xor b);
    layer0_outputs(9018) <= a or b;
    layer0_outputs(9019) <= not b;
    layer0_outputs(9020) <= a xor b;
    layer0_outputs(9021) <= not (a or b);
    layer0_outputs(9022) <= b;
    layer0_outputs(9023) <= a xor b;
    layer0_outputs(9024) <= a;
    layer0_outputs(9025) <= b;
    layer0_outputs(9026) <= a or b;
    layer0_outputs(9027) <= 1'b0;
    layer0_outputs(9028) <= not b;
    layer0_outputs(9029) <= a or b;
    layer0_outputs(9030) <= b;
    layer0_outputs(9031) <= not (a or b);
    layer0_outputs(9032) <= a and b;
    layer0_outputs(9033) <= not (a or b);
    layer0_outputs(9034) <= not a or b;
    layer0_outputs(9035) <= not (a or b);
    layer0_outputs(9036) <= a or b;
    layer0_outputs(9037) <= not (a xor b);
    layer0_outputs(9038) <= not (a or b);
    layer0_outputs(9039) <= not b or a;
    layer0_outputs(9040) <= not b;
    layer0_outputs(9041) <= not (a xor b);
    layer0_outputs(9042) <= a and b;
    layer0_outputs(9043) <= a and not b;
    layer0_outputs(9044) <= a and not b;
    layer0_outputs(9045) <= not (a or b);
    layer0_outputs(9046) <= not b;
    layer0_outputs(9047) <= not (a or b);
    layer0_outputs(9048) <= a;
    layer0_outputs(9049) <= not (a or b);
    layer0_outputs(9050) <= a;
    layer0_outputs(9051) <= not (a xor b);
    layer0_outputs(9052) <= b and not a;
    layer0_outputs(9053) <= a or b;
    layer0_outputs(9054) <= b;
    layer0_outputs(9055) <= not a;
    layer0_outputs(9056) <= not b or a;
    layer0_outputs(9057) <= a or b;
    layer0_outputs(9058) <= not (a xor b);
    layer0_outputs(9059) <= b and not a;
    layer0_outputs(9060) <= a xor b;
    layer0_outputs(9061) <= not b;
    layer0_outputs(9062) <= not (a xor b);
    layer0_outputs(9063) <= a or b;
    layer0_outputs(9064) <= not b;
    layer0_outputs(9065) <= a xor b;
    layer0_outputs(9066) <= a and not b;
    layer0_outputs(9067) <= a;
    layer0_outputs(9068) <= a;
    layer0_outputs(9069) <= a and b;
    layer0_outputs(9070) <= a and b;
    layer0_outputs(9071) <= not (a xor b);
    layer0_outputs(9072) <= not a or b;
    layer0_outputs(9073) <= not a;
    layer0_outputs(9074) <= not (a xor b);
    layer0_outputs(9075) <= not a;
    layer0_outputs(9076) <= 1'b1;
    layer0_outputs(9077) <= b;
    layer0_outputs(9078) <= not (a and b);
    layer0_outputs(9079) <= a or b;
    layer0_outputs(9080) <= a or b;
    layer0_outputs(9081) <= not a;
    layer0_outputs(9082) <= not (a xor b);
    layer0_outputs(9083) <= a or b;
    layer0_outputs(9084) <= a xor b;
    layer0_outputs(9085) <= b;
    layer0_outputs(9086) <= a or b;
    layer0_outputs(9087) <= b;
    layer0_outputs(9088) <= not a or b;
    layer0_outputs(9089) <= b and not a;
    layer0_outputs(9090) <= not a;
    layer0_outputs(9091) <= b;
    layer0_outputs(9092) <= a;
    layer0_outputs(9093) <= not (a or b);
    layer0_outputs(9094) <= a and not b;
    layer0_outputs(9095) <= not (a xor b);
    layer0_outputs(9096) <= not a or b;
    layer0_outputs(9097) <= a xor b;
    layer0_outputs(9098) <= a xor b;
    layer0_outputs(9099) <= a;
    layer0_outputs(9100) <= not b;
    layer0_outputs(9101) <= not (a xor b);
    layer0_outputs(9102) <= not (a xor b);
    layer0_outputs(9103) <= not (a or b);
    layer0_outputs(9104) <= not (a or b);
    layer0_outputs(9105) <= not a or b;
    layer0_outputs(9106) <= b and not a;
    layer0_outputs(9107) <= not a;
    layer0_outputs(9108) <= 1'b1;
    layer0_outputs(9109) <= 1'b0;
    layer0_outputs(9110) <= not a;
    layer0_outputs(9111) <= b and not a;
    layer0_outputs(9112) <= a xor b;
    layer0_outputs(9113) <= a xor b;
    layer0_outputs(9114) <= not b;
    layer0_outputs(9115) <= a xor b;
    layer0_outputs(9116) <= not b;
    layer0_outputs(9117) <= a or b;
    layer0_outputs(9118) <= a or b;
    layer0_outputs(9119) <= b;
    layer0_outputs(9120) <= not (a or b);
    layer0_outputs(9121) <= not (a xor b);
    layer0_outputs(9122) <= a or b;
    layer0_outputs(9123) <= b;
    layer0_outputs(9124) <= a xor b;
    layer0_outputs(9125) <= a or b;
    layer0_outputs(9126) <= a xor b;
    layer0_outputs(9127) <= a or b;
    layer0_outputs(9128) <= b and not a;
    layer0_outputs(9129) <= b;
    layer0_outputs(9130) <= b and not a;
    layer0_outputs(9131) <= not (a or b);
    layer0_outputs(9132) <= not a;
    layer0_outputs(9133) <= not b;
    layer0_outputs(9134) <= not b;
    layer0_outputs(9135) <= not (a and b);
    layer0_outputs(9136) <= b;
    layer0_outputs(9137) <= a or b;
    layer0_outputs(9138) <= not b or a;
    layer0_outputs(9139) <= a xor b;
    layer0_outputs(9140) <= a and not b;
    layer0_outputs(9141) <= not (a or b);
    layer0_outputs(9142) <= a or b;
    layer0_outputs(9143) <= not (a or b);
    layer0_outputs(9144) <= not a;
    layer0_outputs(9145) <= not (a and b);
    layer0_outputs(9146) <= a or b;
    layer0_outputs(9147) <= b;
    layer0_outputs(9148) <= not (a or b);
    layer0_outputs(9149) <= not (a or b);
    layer0_outputs(9150) <= 1'b1;
    layer0_outputs(9151) <= not a or b;
    layer0_outputs(9152) <= b and not a;
    layer0_outputs(9153) <= a or b;
    layer0_outputs(9154) <= 1'b1;
    layer0_outputs(9155) <= a or b;
    layer0_outputs(9156) <= a or b;
    layer0_outputs(9157) <= not b;
    layer0_outputs(9158) <= not b or a;
    layer0_outputs(9159) <= a or b;
    layer0_outputs(9160) <= not a;
    layer0_outputs(9161) <= a and not b;
    layer0_outputs(9162) <= a and b;
    layer0_outputs(9163) <= not a;
    layer0_outputs(9164) <= a xor b;
    layer0_outputs(9165) <= not (a xor b);
    layer0_outputs(9166) <= a or b;
    layer0_outputs(9167) <= not (a xor b);
    layer0_outputs(9168) <= b;
    layer0_outputs(9169) <= a or b;
    layer0_outputs(9170) <= a xor b;
    layer0_outputs(9171) <= a and not b;
    layer0_outputs(9172) <= a;
    layer0_outputs(9173) <= a;
    layer0_outputs(9174) <= not (a or b);
    layer0_outputs(9175) <= not a;
    layer0_outputs(9176) <= not b or a;
    layer0_outputs(9177) <= 1'b1;
    layer0_outputs(9178) <= b;
    layer0_outputs(9179) <= a and not b;
    layer0_outputs(9180) <= a and not b;
    layer0_outputs(9181) <= not (a or b);
    layer0_outputs(9182) <= a xor b;
    layer0_outputs(9183) <= a;
    layer0_outputs(9184) <= a or b;
    layer0_outputs(9185) <= not a;
    layer0_outputs(9186) <= a xor b;
    layer0_outputs(9187) <= not b;
    layer0_outputs(9188) <= a xor b;
    layer0_outputs(9189) <= not (a xor b);
    layer0_outputs(9190) <= a or b;
    layer0_outputs(9191) <= 1'b1;
    layer0_outputs(9192) <= not a or b;
    layer0_outputs(9193) <= not b;
    layer0_outputs(9194) <= not a or b;
    layer0_outputs(9195) <= not a or b;
    layer0_outputs(9196) <= not (a or b);
    layer0_outputs(9197) <= not (a or b);
    layer0_outputs(9198) <= not (a or b);
    layer0_outputs(9199) <= 1'b0;
    layer0_outputs(9200) <= not (a xor b);
    layer0_outputs(9201) <= b and not a;
    layer0_outputs(9202) <= b and not a;
    layer0_outputs(9203) <= a and not b;
    layer0_outputs(9204) <= a xor b;
    layer0_outputs(9205) <= a or b;
    layer0_outputs(9206) <= not (a or b);
    layer0_outputs(9207) <= not (a and b);
    layer0_outputs(9208) <= not (a or b);
    layer0_outputs(9209) <= not (a or b);
    layer0_outputs(9210) <= not (a or b);
    layer0_outputs(9211) <= not (a or b);
    layer0_outputs(9212) <= not (a or b);
    layer0_outputs(9213) <= 1'b0;
    layer0_outputs(9214) <= not a or b;
    layer0_outputs(9215) <= a;
    layer0_outputs(9216) <= a xor b;
    layer0_outputs(9217) <= not (a xor b);
    layer0_outputs(9218) <= not a;
    layer0_outputs(9219) <= not (a or b);
    layer0_outputs(9220) <= not b or a;
    layer0_outputs(9221) <= a;
    layer0_outputs(9222) <= not (a xor b);
    layer0_outputs(9223) <= a or b;
    layer0_outputs(9224) <= a or b;
    layer0_outputs(9225) <= not a;
    layer0_outputs(9226) <= not (a and b);
    layer0_outputs(9227) <= b;
    layer0_outputs(9228) <= a;
    layer0_outputs(9229) <= not (a xor b);
    layer0_outputs(9230) <= a;
    layer0_outputs(9231) <= a;
    layer0_outputs(9232) <= not a;
    layer0_outputs(9233) <= not (a or b);
    layer0_outputs(9234) <= a;
    layer0_outputs(9235) <= a and not b;
    layer0_outputs(9236) <= not (a xor b);
    layer0_outputs(9237) <= not b or a;
    layer0_outputs(9238) <= not (a xor b);
    layer0_outputs(9239) <= not b or a;
    layer0_outputs(9240) <= a;
    layer0_outputs(9241) <= a xor b;
    layer0_outputs(9242) <= a and not b;
    layer0_outputs(9243) <= a or b;
    layer0_outputs(9244) <= a;
    layer0_outputs(9245) <= a and b;
    layer0_outputs(9246) <= not (a xor b);
    layer0_outputs(9247) <= b and not a;
    layer0_outputs(9248) <= a xor b;
    layer0_outputs(9249) <= 1'b0;
    layer0_outputs(9250) <= not (a or b);
    layer0_outputs(9251) <= not b or a;
    layer0_outputs(9252) <= not a;
    layer0_outputs(9253) <= not a;
    layer0_outputs(9254) <= not a or b;
    layer0_outputs(9255) <= a xor b;
    layer0_outputs(9256) <= a xor b;
    layer0_outputs(9257) <= not (a and b);
    layer0_outputs(9258) <= not a;
    layer0_outputs(9259) <= a or b;
    layer0_outputs(9260) <= a and not b;
    layer0_outputs(9261) <= not b or a;
    layer0_outputs(9262) <= b and not a;
    layer0_outputs(9263) <= a xor b;
    layer0_outputs(9264) <= not a or b;
    layer0_outputs(9265) <= b and not a;
    layer0_outputs(9266) <= not a;
    layer0_outputs(9267) <= not b or a;
    layer0_outputs(9268) <= b;
    layer0_outputs(9269) <= a xor b;
    layer0_outputs(9270) <= a or b;
    layer0_outputs(9271) <= not a or b;
    layer0_outputs(9272) <= not a or b;
    layer0_outputs(9273) <= 1'b0;
    layer0_outputs(9274) <= b;
    layer0_outputs(9275) <= a or b;
    layer0_outputs(9276) <= not b;
    layer0_outputs(9277) <= not (a xor b);
    layer0_outputs(9278) <= not a or b;
    layer0_outputs(9279) <= not (a and b);
    layer0_outputs(9280) <= a;
    layer0_outputs(9281) <= b and not a;
    layer0_outputs(9282) <= b;
    layer0_outputs(9283) <= a and not b;
    layer0_outputs(9284) <= not (a xor b);
    layer0_outputs(9285) <= a;
    layer0_outputs(9286) <= a;
    layer0_outputs(9287) <= a xor b;
    layer0_outputs(9288) <= not (a or b);
    layer0_outputs(9289) <= a and b;
    layer0_outputs(9290) <= a;
    layer0_outputs(9291) <= not b;
    layer0_outputs(9292) <= a;
    layer0_outputs(9293) <= a and not b;
    layer0_outputs(9294) <= b and not a;
    layer0_outputs(9295) <= a or b;
    layer0_outputs(9296) <= not a or b;
    layer0_outputs(9297) <= not (a and b);
    layer0_outputs(9298) <= not (a or b);
    layer0_outputs(9299) <= a;
    layer0_outputs(9300) <= not a or b;
    layer0_outputs(9301) <= b;
    layer0_outputs(9302) <= not (a xor b);
    layer0_outputs(9303) <= not (a xor b);
    layer0_outputs(9304) <= not (a or b);
    layer0_outputs(9305) <= a xor b;
    layer0_outputs(9306) <= b and not a;
    layer0_outputs(9307) <= a or b;
    layer0_outputs(9308) <= not b or a;
    layer0_outputs(9309) <= not (a and b);
    layer0_outputs(9310) <= a or b;
    layer0_outputs(9311) <= b;
    layer0_outputs(9312) <= a and b;
    layer0_outputs(9313) <= b;
    layer0_outputs(9314) <= a;
    layer0_outputs(9315) <= 1'b1;
    layer0_outputs(9316) <= a or b;
    layer0_outputs(9317) <= not b;
    layer0_outputs(9318) <= a xor b;
    layer0_outputs(9319) <= a and not b;
    layer0_outputs(9320) <= a;
    layer0_outputs(9321) <= not a or b;
    layer0_outputs(9322) <= b;
    layer0_outputs(9323) <= not (a xor b);
    layer0_outputs(9324) <= not b;
    layer0_outputs(9325) <= not (a or b);
    layer0_outputs(9326) <= 1'b0;
    layer0_outputs(9327) <= b;
    layer0_outputs(9328) <= not a or b;
    layer0_outputs(9329) <= not b;
    layer0_outputs(9330) <= a xor b;
    layer0_outputs(9331) <= a;
    layer0_outputs(9332) <= not (a or b);
    layer0_outputs(9333) <= a and not b;
    layer0_outputs(9334) <= 1'b1;
    layer0_outputs(9335) <= a xor b;
    layer0_outputs(9336) <= b and not a;
    layer0_outputs(9337) <= a and b;
    layer0_outputs(9338) <= a xor b;
    layer0_outputs(9339) <= not a or b;
    layer0_outputs(9340) <= a and not b;
    layer0_outputs(9341) <= a xor b;
    layer0_outputs(9342) <= a xor b;
    layer0_outputs(9343) <= not a;
    layer0_outputs(9344) <= a;
    layer0_outputs(9345) <= a xor b;
    layer0_outputs(9346) <= not b;
    layer0_outputs(9347) <= not (a or b);
    layer0_outputs(9348) <= a;
    layer0_outputs(9349) <= not (a or b);
    layer0_outputs(9350) <= not a;
    layer0_outputs(9351) <= b and not a;
    layer0_outputs(9352) <= a or b;
    layer0_outputs(9353) <= b;
    layer0_outputs(9354) <= a and not b;
    layer0_outputs(9355) <= a;
    layer0_outputs(9356) <= not (a xor b);
    layer0_outputs(9357) <= not a or b;
    layer0_outputs(9358) <= not (a xor b);
    layer0_outputs(9359) <= a and b;
    layer0_outputs(9360) <= a or b;
    layer0_outputs(9361) <= b and not a;
    layer0_outputs(9362) <= b and not a;
    layer0_outputs(9363) <= a or b;
    layer0_outputs(9364) <= a and b;
    layer0_outputs(9365) <= not (a or b);
    layer0_outputs(9366) <= not a or b;
    layer0_outputs(9367) <= a and not b;
    layer0_outputs(9368) <= a or b;
    layer0_outputs(9369) <= b and not a;
    layer0_outputs(9370) <= not b;
    layer0_outputs(9371) <= a xor b;
    layer0_outputs(9372) <= not b;
    layer0_outputs(9373) <= a and b;
    layer0_outputs(9374) <= a and not b;
    layer0_outputs(9375) <= b and not a;
    layer0_outputs(9376) <= not (a xor b);
    layer0_outputs(9377) <= not (a or b);
    layer0_outputs(9378) <= not (a or b);
    layer0_outputs(9379) <= b;
    layer0_outputs(9380) <= a xor b;
    layer0_outputs(9381) <= not a or b;
    layer0_outputs(9382) <= a;
    layer0_outputs(9383) <= not b;
    layer0_outputs(9384) <= not (a xor b);
    layer0_outputs(9385) <= a and not b;
    layer0_outputs(9386) <= a and b;
    layer0_outputs(9387) <= not (a or b);
    layer0_outputs(9388) <= a or b;
    layer0_outputs(9389) <= not b or a;
    layer0_outputs(9390) <= a or b;
    layer0_outputs(9391) <= not a;
    layer0_outputs(9392) <= not b;
    layer0_outputs(9393) <= not a;
    layer0_outputs(9394) <= not (a or b);
    layer0_outputs(9395) <= a and b;
    layer0_outputs(9396) <= not b or a;
    layer0_outputs(9397) <= a or b;
    layer0_outputs(9398) <= not (a xor b);
    layer0_outputs(9399) <= not a;
    layer0_outputs(9400) <= a or b;
    layer0_outputs(9401) <= a;
    layer0_outputs(9402) <= not b;
    layer0_outputs(9403) <= not (a or b);
    layer0_outputs(9404) <= a xor b;
    layer0_outputs(9405) <= not (a and b);
    layer0_outputs(9406) <= not b or a;
    layer0_outputs(9407) <= b and not a;
    layer0_outputs(9408) <= not a or b;
    layer0_outputs(9409) <= not (a xor b);
    layer0_outputs(9410) <= a and b;
    layer0_outputs(9411) <= not a;
    layer0_outputs(9412) <= a or b;
    layer0_outputs(9413) <= not b;
    layer0_outputs(9414) <= not b or a;
    layer0_outputs(9415) <= not b or a;
    layer0_outputs(9416) <= 1'b0;
    layer0_outputs(9417) <= a and b;
    layer0_outputs(9418) <= not (a xor b);
    layer0_outputs(9419) <= a xor b;
    layer0_outputs(9420) <= a or b;
    layer0_outputs(9421) <= not (a xor b);
    layer0_outputs(9422) <= a and not b;
    layer0_outputs(9423) <= a and b;
    layer0_outputs(9424) <= not a or b;
    layer0_outputs(9425) <= a or b;
    layer0_outputs(9426) <= not (a xor b);
    layer0_outputs(9427) <= a and b;
    layer0_outputs(9428) <= 1'b1;
    layer0_outputs(9429) <= not (a xor b);
    layer0_outputs(9430) <= b;
    layer0_outputs(9431) <= not (a and b);
    layer0_outputs(9432) <= a xor b;
    layer0_outputs(9433) <= 1'b0;
    layer0_outputs(9434) <= a or b;
    layer0_outputs(9435) <= not a;
    layer0_outputs(9436) <= a or b;
    layer0_outputs(9437) <= b;
    layer0_outputs(9438) <= a or b;
    layer0_outputs(9439) <= a or b;
    layer0_outputs(9440) <= a and b;
    layer0_outputs(9441) <= not (a xor b);
    layer0_outputs(9442) <= not b;
    layer0_outputs(9443) <= not (a xor b);
    layer0_outputs(9444) <= a xor b;
    layer0_outputs(9445) <= b;
    layer0_outputs(9446) <= not b or a;
    layer0_outputs(9447) <= not a;
    layer0_outputs(9448) <= not (a and b);
    layer0_outputs(9449) <= not a;
    layer0_outputs(9450) <= not a;
    layer0_outputs(9451) <= a xor b;
    layer0_outputs(9452) <= b and not a;
    layer0_outputs(9453) <= not a;
    layer0_outputs(9454) <= a or b;
    layer0_outputs(9455) <= a xor b;
    layer0_outputs(9456) <= not (a xor b);
    layer0_outputs(9457) <= not a;
    layer0_outputs(9458) <= a and not b;
    layer0_outputs(9459) <= b and not a;
    layer0_outputs(9460) <= a or b;
    layer0_outputs(9461) <= a;
    layer0_outputs(9462) <= not (a xor b);
    layer0_outputs(9463) <= a or b;
    layer0_outputs(9464) <= a;
    layer0_outputs(9465) <= a xor b;
    layer0_outputs(9466) <= 1'b0;
    layer0_outputs(9467) <= a or b;
    layer0_outputs(9468) <= not a or b;
    layer0_outputs(9469) <= not (a xor b);
    layer0_outputs(9470) <= not a;
    layer0_outputs(9471) <= not b or a;
    layer0_outputs(9472) <= not (a or b);
    layer0_outputs(9473) <= not (a xor b);
    layer0_outputs(9474) <= not (a and b);
    layer0_outputs(9475) <= a and not b;
    layer0_outputs(9476) <= not b;
    layer0_outputs(9477) <= b;
    layer0_outputs(9478) <= a or b;
    layer0_outputs(9479) <= not (a or b);
    layer0_outputs(9480) <= not a;
    layer0_outputs(9481) <= b and not a;
    layer0_outputs(9482) <= a and b;
    layer0_outputs(9483) <= not a or b;
    layer0_outputs(9484) <= a;
    layer0_outputs(9485) <= not a or b;
    layer0_outputs(9486) <= b and not a;
    layer0_outputs(9487) <= not (a or b);
    layer0_outputs(9488) <= not (a and b);
    layer0_outputs(9489) <= not (a and b);
    layer0_outputs(9490) <= b;
    layer0_outputs(9491) <= a and not b;
    layer0_outputs(9492) <= not b or a;
    layer0_outputs(9493) <= not (a xor b);
    layer0_outputs(9494) <= not a;
    layer0_outputs(9495) <= a;
    layer0_outputs(9496) <= a xor b;
    layer0_outputs(9497) <= not a;
    layer0_outputs(9498) <= a and b;
    layer0_outputs(9499) <= b;
    layer0_outputs(9500) <= b;
    layer0_outputs(9501) <= a xor b;
    layer0_outputs(9502) <= not a;
    layer0_outputs(9503) <= a xor b;
    layer0_outputs(9504) <= b and not a;
    layer0_outputs(9505) <= not b or a;
    layer0_outputs(9506) <= b and not a;
    layer0_outputs(9507) <= a or b;
    layer0_outputs(9508) <= not (a or b);
    layer0_outputs(9509) <= not (a or b);
    layer0_outputs(9510) <= b;
    layer0_outputs(9511) <= not b;
    layer0_outputs(9512) <= not (a or b);
    layer0_outputs(9513) <= a xor b;
    layer0_outputs(9514) <= a and b;
    layer0_outputs(9515) <= not a;
    layer0_outputs(9516) <= b and not a;
    layer0_outputs(9517) <= not a;
    layer0_outputs(9518) <= b;
    layer0_outputs(9519) <= 1'b1;
    layer0_outputs(9520) <= b;
    layer0_outputs(9521) <= not (a and b);
    layer0_outputs(9522) <= not a;
    layer0_outputs(9523) <= b and not a;
    layer0_outputs(9524) <= not (a and b);
    layer0_outputs(9525) <= a;
    layer0_outputs(9526) <= b;
    layer0_outputs(9527) <= not a or b;
    layer0_outputs(9528) <= not b;
    layer0_outputs(9529) <= a or b;
    layer0_outputs(9530) <= not (a xor b);
    layer0_outputs(9531) <= b and not a;
    layer0_outputs(9532) <= not (a xor b);
    layer0_outputs(9533) <= a xor b;
    layer0_outputs(9534) <= not b;
    layer0_outputs(9535) <= b;
    layer0_outputs(9536) <= a or b;
    layer0_outputs(9537) <= not b or a;
    layer0_outputs(9538) <= b;
    layer0_outputs(9539) <= not (a xor b);
    layer0_outputs(9540) <= a xor b;
    layer0_outputs(9541) <= b;
    layer0_outputs(9542) <= b and not a;
    layer0_outputs(9543) <= a xor b;
    layer0_outputs(9544) <= a;
    layer0_outputs(9545) <= a xor b;
    layer0_outputs(9546) <= a or b;
    layer0_outputs(9547) <= 1'b1;
    layer0_outputs(9548) <= a;
    layer0_outputs(9549) <= not a or b;
    layer0_outputs(9550) <= not (a or b);
    layer0_outputs(9551) <= a and b;
    layer0_outputs(9552) <= not b;
    layer0_outputs(9553) <= not b or a;
    layer0_outputs(9554) <= not a or b;
    layer0_outputs(9555) <= not a;
    layer0_outputs(9556) <= a or b;
    layer0_outputs(9557) <= a or b;
    layer0_outputs(9558) <= b and not a;
    layer0_outputs(9559) <= a xor b;
    layer0_outputs(9560) <= not b or a;
    layer0_outputs(9561) <= b;
    layer0_outputs(9562) <= not a or b;
    layer0_outputs(9563) <= not a;
    layer0_outputs(9564) <= not b;
    layer0_outputs(9565) <= not (a xor b);
    layer0_outputs(9566) <= not a;
    layer0_outputs(9567) <= b and not a;
    layer0_outputs(9568) <= a and b;
    layer0_outputs(9569) <= a or b;
    layer0_outputs(9570) <= not (a and b);
    layer0_outputs(9571) <= a or b;
    layer0_outputs(9572) <= b and not a;
    layer0_outputs(9573) <= not (a xor b);
    layer0_outputs(9574) <= not b or a;
    layer0_outputs(9575) <= not a or b;
    layer0_outputs(9576) <= b and not a;
    layer0_outputs(9577) <= not (a xor b);
    layer0_outputs(9578) <= a and b;
    layer0_outputs(9579) <= a xor b;
    layer0_outputs(9580) <= not (a and b);
    layer0_outputs(9581) <= a xor b;
    layer0_outputs(9582) <= not (a xor b);
    layer0_outputs(9583) <= not a or b;
    layer0_outputs(9584) <= b and not a;
    layer0_outputs(9585) <= a xor b;
    layer0_outputs(9586) <= not (a xor b);
    layer0_outputs(9587) <= 1'b0;
    layer0_outputs(9588) <= b and not a;
    layer0_outputs(9589) <= 1'b1;
    layer0_outputs(9590) <= a;
    layer0_outputs(9591) <= not b or a;
    layer0_outputs(9592) <= a xor b;
    layer0_outputs(9593) <= not (a xor b);
    layer0_outputs(9594) <= not (a or b);
    layer0_outputs(9595) <= 1'b0;
    layer0_outputs(9596) <= not a;
    layer0_outputs(9597) <= a;
    layer0_outputs(9598) <= a xor b;
    layer0_outputs(9599) <= a and not b;
    layer0_outputs(9600) <= a xor b;
    layer0_outputs(9601) <= a or b;
    layer0_outputs(9602) <= not (a xor b);
    layer0_outputs(9603) <= a xor b;
    layer0_outputs(9604) <= a;
    layer0_outputs(9605) <= a xor b;
    layer0_outputs(9606) <= not (a and b);
    layer0_outputs(9607) <= not a;
    layer0_outputs(9608) <= not (a or b);
    layer0_outputs(9609) <= not a;
    layer0_outputs(9610) <= not (a and b);
    layer0_outputs(9611) <= b;
    layer0_outputs(9612) <= a;
    layer0_outputs(9613) <= a and b;
    layer0_outputs(9614) <= not (a xor b);
    layer0_outputs(9615) <= not b or a;
    layer0_outputs(9616) <= a xor b;
    layer0_outputs(9617) <= a xor b;
    layer0_outputs(9618) <= a and not b;
    layer0_outputs(9619) <= a xor b;
    layer0_outputs(9620) <= not (a or b);
    layer0_outputs(9621) <= not b;
    layer0_outputs(9622) <= not a;
    layer0_outputs(9623) <= b;
    layer0_outputs(9624) <= not b;
    layer0_outputs(9625) <= a or b;
    layer0_outputs(9626) <= a or b;
    layer0_outputs(9627) <= a xor b;
    layer0_outputs(9628) <= a or b;
    layer0_outputs(9629) <= b;
    layer0_outputs(9630) <= not (a or b);
    layer0_outputs(9631) <= a;
    layer0_outputs(9632) <= not a;
    layer0_outputs(9633) <= not (a or b);
    layer0_outputs(9634) <= not (a or b);
    layer0_outputs(9635) <= 1'b1;
    layer0_outputs(9636) <= b;
    layer0_outputs(9637) <= not (a or b);
    layer0_outputs(9638) <= not a or b;
    layer0_outputs(9639) <= not (a xor b);
    layer0_outputs(9640) <= not (a or b);
    layer0_outputs(9641) <= a xor b;
    layer0_outputs(9642) <= not (a xor b);
    layer0_outputs(9643) <= not (a or b);
    layer0_outputs(9644) <= a or b;
    layer0_outputs(9645) <= a xor b;
    layer0_outputs(9646) <= a;
    layer0_outputs(9647) <= not a or b;
    layer0_outputs(9648) <= not (a xor b);
    layer0_outputs(9649) <= not a;
    layer0_outputs(9650) <= b and not a;
    layer0_outputs(9651) <= not (a or b);
    layer0_outputs(9652) <= not b or a;
    layer0_outputs(9653) <= b and not a;
    layer0_outputs(9654) <= a or b;
    layer0_outputs(9655) <= not b or a;
    layer0_outputs(9656) <= not b;
    layer0_outputs(9657) <= not b or a;
    layer0_outputs(9658) <= a or b;
    layer0_outputs(9659) <= not b;
    layer0_outputs(9660) <= not b;
    layer0_outputs(9661) <= not (a or b);
    layer0_outputs(9662) <= not (a or b);
    layer0_outputs(9663) <= b;
    layer0_outputs(9664) <= not a;
    layer0_outputs(9665) <= not (a xor b);
    layer0_outputs(9666) <= not (a xor b);
    layer0_outputs(9667) <= a xor b;
    layer0_outputs(9668) <= not (a or b);
    layer0_outputs(9669) <= not (a or b);
    layer0_outputs(9670) <= a or b;
    layer0_outputs(9671) <= not (a or b);
    layer0_outputs(9672) <= 1'b0;
    layer0_outputs(9673) <= not b or a;
    layer0_outputs(9674) <= a xor b;
    layer0_outputs(9675) <= not b;
    layer0_outputs(9676) <= b;
    layer0_outputs(9677) <= not a or b;
    layer0_outputs(9678) <= not a or b;
    layer0_outputs(9679) <= not a;
    layer0_outputs(9680) <= a xor b;
    layer0_outputs(9681) <= not a or b;
    layer0_outputs(9682) <= a and not b;
    layer0_outputs(9683) <= not a or b;
    layer0_outputs(9684) <= a;
    layer0_outputs(9685) <= not b or a;
    layer0_outputs(9686) <= a and not b;
    layer0_outputs(9687) <= not b;
    layer0_outputs(9688) <= b and not a;
    layer0_outputs(9689) <= b and not a;
    layer0_outputs(9690) <= 1'b1;
    layer0_outputs(9691) <= a xor b;
    layer0_outputs(9692) <= not a;
    layer0_outputs(9693) <= a xor b;
    layer0_outputs(9694) <= a xor b;
    layer0_outputs(9695) <= 1'b0;
    layer0_outputs(9696) <= b;
    layer0_outputs(9697) <= not (a or b);
    layer0_outputs(9698) <= a;
    layer0_outputs(9699) <= not (a or b);
    layer0_outputs(9700) <= not (a or b);
    layer0_outputs(9701) <= a or b;
    layer0_outputs(9702) <= a xor b;
    layer0_outputs(9703) <= not a or b;
    layer0_outputs(9704) <= a;
    layer0_outputs(9705) <= a xor b;
    layer0_outputs(9706) <= not b or a;
    layer0_outputs(9707) <= not (a or b);
    layer0_outputs(9708) <= not a or b;
    layer0_outputs(9709) <= a xor b;
    layer0_outputs(9710) <= b and not a;
    layer0_outputs(9711) <= a xor b;
    layer0_outputs(9712) <= not a;
    layer0_outputs(9713) <= not (a or b);
    layer0_outputs(9714) <= a and not b;
    layer0_outputs(9715) <= not (a or b);
    layer0_outputs(9716) <= b and not a;
    layer0_outputs(9717) <= a and not b;
    layer0_outputs(9718) <= b;
    layer0_outputs(9719) <= a xor b;
    layer0_outputs(9720) <= not (a or b);
    layer0_outputs(9721) <= not a;
    layer0_outputs(9722) <= a or b;
    layer0_outputs(9723) <= a or b;
    layer0_outputs(9724) <= not (a xor b);
    layer0_outputs(9725) <= not a;
    layer0_outputs(9726) <= a or b;
    layer0_outputs(9727) <= not (a or b);
    layer0_outputs(9728) <= a and not b;
    layer0_outputs(9729) <= not (a or b);
    layer0_outputs(9730) <= not (a xor b);
    layer0_outputs(9731) <= not (a or b);
    layer0_outputs(9732) <= not a or b;
    layer0_outputs(9733) <= a or b;
    layer0_outputs(9734) <= not (a xor b);
    layer0_outputs(9735) <= a and b;
    layer0_outputs(9736) <= not (a and b);
    layer0_outputs(9737) <= not (a or b);
    layer0_outputs(9738) <= not a;
    layer0_outputs(9739) <= not a;
    layer0_outputs(9740) <= 1'b0;
    layer0_outputs(9741) <= not a;
    layer0_outputs(9742) <= a and not b;
    layer0_outputs(9743) <= not a or b;
    layer0_outputs(9744) <= b;
    layer0_outputs(9745) <= not (a xor b);
    layer0_outputs(9746) <= a and not b;
    layer0_outputs(9747) <= not b or a;
    layer0_outputs(9748) <= not b;
    layer0_outputs(9749) <= a or b;
    layer0_outputs(9750) <= b and not a;
    layer0_outputs(9751) <= b and not a;
    layer0_outputs(9752) <= a or b;
    layer0_outputs(9753) <= not b;
    layer0_outputs(9754) <= a;
    layer0_outputs(9755) <= not a;
    layer0_outputs(9756) <= 1'b0;
    layer0_outputs(9757) <= not (a or b);
    layer0_outputs(9758) <= a and not b;
    layer0_outputs(9759) <= a or b;
    layer0_outputs(9760) <= 1'b0;
    layer0_outputs(9761) <= a xor b;
    layer0_outputs(9762) <= a or b;
    layer0_outputs(9763) <= not a;
    layer0_outputs(9764) <= 1'b1;
    layer0_outputs(9765) <= a and b;
    layer0_outputs(9766) <= not (a xor b);
    layer0_outputs(9767) <= a or b;
    layer0_outputs(9768) <= a and not b;
    layer0_outputs(9769) <= a or b;
    layer0_outputs(9770) <= not (a or b);
    layer0_outputs(9771) <= a or b;
    layer0_outputs(9772) <= b;
    layer0_outputs(9773) <= a;
    layer0_outputs(9774) <= a and b;
    layer0_outputs(9775) <= not (a or b);
    layer0_outputs(9776) <= b;
    layer0_outputs(9777) <= a and not b;
    layer0_outputs(9778) <= not a;
    layer0_outputs(9779) <= b and not a;
    layer0_outputs(9780) <= not b;
    layer0_outputs(9781) <= not (a xor b);
    layer0_outputs(9782) <= not a;
    layer0_outputs(9783) <= a;
    layer0_outputs(9784) <= not b or a;
    layer0_outputs(9785) <= not b;
    layer0_outputs(9786) <= b and not a;
    layer0_outputs(9787) <= not (a or b);
    layer0_outputs(9788) <= b and not a;
    layer0_outputs(9789) <= not (a xor b);
    layer0_outputs(9790) <= not (a or b);
    layer0_outputs(9791) <= a and not b;
    layer0_outputs(9792) <= not b or a;
    layer0_outputs(9793) <= not b;
    layer0_outputs(9794) <= not a or b;
    layer0_outputs(9795) <= not (a or b);
    layer0_outputs(9796) <= not a;
    layer0_outputs(9797) <= a or b;
    layer0_outputs(9798) <= not a;
    layer0_outputs(9799) <= not a;
    layer0_outputs(9800) <= not a or b;
    layer0_outputs(9801) <= not b;
    layer0_outputs(9802) <= not b;
    layer0_outputs(9803) <= not (a xor b);
    layer0_outputs(9804) <= not (a xor b);
    layer0_outputs(9805) <= a and not b;
    layer0_outputs(9806) <= not a or b;
    layer0_outputs(9807) <= b;
    layer0_outputs(9808) <= b and not a;
    layer0_outputs(9809) <= a or b;
    layer0_outputs(9810) <= a;
    layer0_outputs(9811) <= b and not a;
    layer0_outputs(9812) <= not a or b;
    layer0_outputs(9813) <= a xor b;
    layer0_outputs(9814) <= a;
    layer0_outputs(9815) <= not (a and b);
    layer0_outputs(9816) <= not a;
    layer0_outputs(9817) <= not (a xor b);
    layer0_outputs(9818) <= not b;
    layer0_outputs(9819) <= a and not b;
    layer0_outputs(9820) <= not (a or b);
    layer0_outputs(9821) <= b;
    layer0_outputs(9822) <= not (a xor b);
    layer0_outputs(9823) <= not (a xor b);
    layer0_outputs(9824) <= a and not b;
    layer0_outputs(9825) <= not b;
    layer0_outputs(9826) <= b;
    layer0_outputs(9827) <= a;
    layer0_outputs(9828) <= b;
    layer0_outputs(9829) <= a xor b;
    layer0_outputs(9830) <= not (a or b);
    layer0_outputs(9831) <= a and not b;
    layer0_outputs(9832) <= not a;
    layer0_outputs(9833) <= a or b;
    layer0_outputs(9834) <= b;
    layer0_outputs(9835) <= a and not b;
    layer0_outputs(9836) <= a xor b;
    layer0_outputs(9837) <= a xor b;
    layer0_outputs(9838) <= a or b;
    layer0_outputs(9839) <= not a;
    layer0_outputs(9840) <= not b;
    layer0_outputs(9841) <= b;
    layer0_outputs(9842) <= not (a xor b);
    layer0_outputs(9843) <= a or b;
    layer0_outputs(9844) <= not (a or b);
    layer0_outputs(9845) <= not (a xor b);
    layer0_outputs(9846) <= not (a or b);
    layer0_outputs(9847) <= b and not a;
    layer0_outputs(9848) <= b and not a;
    layer0_outputs(9849) <= not b or a;
    layer0_outputs(9850) <= not (a xor b);
    layer0_outputs(9851) <= not (a xor b);
    layer0_outputs(9852) <= a or b;
    layer0_outputs(9853) <= not a;
    layer0_outputs(9854) <= a;
    layer0_outputs(9855) <= not (a or b);
    layer0_outputs(9856) <= not b;
    layer0_outputs(9857) <= 1'b1;
    layer0_outputs(9858) <= b and not a;
    layer0_outputs(9859) <= b and not a;
    layer0_outputs(9860) <= not b;
    layer0_outputs(9861) <= a xor b;
    layer0_outputs(9862) <= not (a or b);
    layer0_outputs(9863) <= not b;
    layer0_outputs(9864) <= not b;
    layer0_outputs(9865) <= a xor b;
    layer0_outputs(9866) <= 1'b1;
    layer0_outputs(9867) <= a;
    layer0_outputs(9868) <= a xor b;
    layer0_outputs(9869) <= not (a or b);
    layer0_outputs(9870) <= not a;
    layer0_outputs(9871) <= not b;
    layer0_outputs(9872) <= a and not b;
    layer0_outputs(9873) <= a;
    layer0_outputs(9874) <= 1'b1;
    layer0_outputs(9875) <= b and not a;
    layer0_outputs(9876) <= not (a and b);
    layer0_outputs(9877) <= not (a or b);
    layer0_outputs(9878) <= not a;
    layer0_outputs(9879) <= not (a or b);
    layer0_outputs(9880) <= a and not b;
    layer0_outputs(9881) <= a or b;
    layer0_outputs(9882) <= not a or b;
    layer0_outputs(9883) <= a xor b;
    layer0_outputs(9884) <= a or b;
    layer0_outputs(9885) <= not (a or b);
    layer0_outputs(9886) <= b and not a;
    layer0_outputs(9887) <= not a;
    layer0_outputs(9888) <= not b or a;
    layer0_outputs(9889) <= b;
    layer0_outputs(9890) <= not (a or b);
    layer0_outputs(9891) <= a xor b;
    layer0_outputs(9892) <= a or b;
    layer0_outputs(9893) <= not (a xor b);
    layer0_outputs(9894) <= a or b;
    layer0_outputs(9895) <= a xor b;
    layer0_outputs(9896) <= b and not a;
    layer0_outputs(9897) <= b;
    layer0_outputs(9898) <= not (a xor b);
    layer0_outputs(9899) <= a or b;
    layer0_outputs(9900) <= a and not b;
    layer0_outputs(9901) <= b;
    layer0_outputs(9902) <= not (a or b);
    layer0_outputs(9903) <= not b or a;
    layer0_outputs(9904) <= a and not b;
    layer0_outputs(9905) <= not (a or b);
    layer0_outputs(9906) <= not a or b;
    layer0_outputs(9907) <= a and b;
    layer0_outputs(9908) <= not (a or b);
    layer0_outputs(9909) <= a and not b;
    layer0_outputs(9910) <= a xor b;
    layer0_outputs(9911) <= a xor b;
    layer0_outputs(9912) <= 1'b0;
    layer0_outputs(9913) <= a xor b;
    layer0_outputs(9914) <= not a;
    layer0_outputs(9915) <= 1'b1;
    layer0_outputs(9916) <= not (a or b);
    layer0_outputs(9917) <= a or b;
    layer0_outputs(9918) <= not b;
    layer0_outputs(9919) <= not (a or b);
    layer0_outputs(9920) <= not (a xor b);
    layer0_outputs(9921) <= b and not a;
    layer0_outputs(9922) <= not b;
    layer0_outputs(9923) <= not (a or b);
    layer0_outputs(9924) <= not b;
    layer0_outputs(9925) <= not b or a;
    layer0_outputs(9926) <= not b or a;
    layer0_outputs(9927) <= a;
    layer0_outputs(9928) <= b and not a;
    layer0_outputs(9929) <= not (a or b);
    layer0_outputs(9930) <= not a or b;
    layer0_outputs(9931) <= not (a xor b);
    layer0_outputs(9932) <= a and not b;
    layer0_outputs(9933) <= not b or a;
    layer0_outputs(9934) <= a and b;
    layer0_outputs(9935) <= a;
    layer0_outputs(9936) <= not (a xor b);
    layer0_outputs(9937) <= a;
    layer0_outputs(9938) <= not a or b;
    layer0_outputs(9939) <= not b or a;
    layer0_outputs(9940) <= a xor b;
    layer0_outputs(9941) <= not a;
    layer0_outputs(9942) <= not a;
    layer0_outputs(9943) <= 1'b0;
    layer0_outputs(9944) <= not b or a;
    layer0_outputs(9945) <= not b;
    layer0_outputs(9946) <= not a or b;
    layer0_outputs(9947) <= b;
    layer0_outputs(9948) <= not b;
    layer0_outputs(9949) <= not (a or b);
    layer0_outputs(9950) <= not a or b;
    layer0_outputs(9951) <= not (a xor b);
    layer0_outputs(9952) <= not (a or b);
    layer0_outputs(9953) <= a and not b;
    layer0_outputs(9954) <= not b;
    layer0_outputs(9955) <= not (a xor b);
    layer0_outputs(9956) <= not (a or b);
    layer0_outputs(9957) <= a or b;
    layer0_outputs(9958) <= not (a or b);
    layer0_outputs(9959) <= b and not a;
    layer0_outputs(9960) <= a;
    layer0_outputs(9961) <= a xor b;
    layer0_outputs(9962) <= not (a xor b);
    layer0_outputs(9963) <= b;
    layer0_outputs(9964) <= not a or b;
    layer0_outputs(9965) <= b and not a;
    layer0_outputs(9966) <= not (a and b);
    layer0_outputs(9967) <= a or b;
    layer0_outputs(9968) <= not a or b;
    layer0_outputs(9969) <= a or b;
    layer0_outputs(9970) <= b and not a;
    layer0_outputs(9971) <= not (a xor b);
    layer0_outputs(9972) <= not b or a;
    layer0_outputs(9973) <= not b;
    layer0_outputs(9974) <= not (a xor b);
    layer0_outputs(9975) <= a or b;
    layer0_outputs(9976) <= not (a or b);
    layer0_outputs(9977) <= not (a and b);
    layer0_outputs(9978) <= not (a and b);
    layer0_outputs(9979) <= not b;
    layer0_outputs(9980) <= not (a or b);
    layer0_outputs(9981) <= a;
    layer0_outputs(9982) <= b;
    layer0_outputs(9983) <= not a;
    layer0_outputs(9984) <= 1'b0;
    layer0_outputs(9985) <= not b or a;
    layer0_outputs(9986) <= not (a or b);
    layer0_outputs(9987) <= b;
    layer0_outputs(9988) <= not a or b;
    layer0_outputs(9989) <= a xor b;
    layer0_outputs(9990) <= not b;
    layer0_outputs(9991) <= a and b;
    layer0_outputs(9992) <= a or b;
    layer0_outputs(9993) <= b and not a;
    layer0_outputs(9994) <= not a;
    layer0_outputs(9995) <= a and b;
    layer0_outputs(9996) <= a xor b;
    layer0_outputs(9997) <= not (a xor b);
    layer0_outputs(9998) <= not a or b;
    layer0_outputs(9999) <= not a;
    layer0_outputs(10000) <= a;
    layer0_outputs(10001) <= not (a or b);
    layer0_outputs(10002) <= b and not a;
    layer0_outputs(10003) <= a or b;
    layer0_outputs(10004) <= not (a or b);
    layer0_outputs(10005) <= not b;
    layer0_outputs(10006) <= not (a or b);
    layer0_outputs(10007) <= not a;
    layer0_outputs(10008) <= a xor b;
    layer0_outputs(10009) <= a or b;
    layer0_outputs(10010) <= not (a or b);
    layer0_outputs(10011) <= not a;
    layer0_outputs(10012) <= not (a and b);
    layer0_outputs(10013) <= a or b;
    layer0_outputs(10014) <= b;
    layer0_outputs(10015) <= a xor b;
    layer0_outputs(10016) <= 1'b1;
    layer0_outputs(10017) <= 1'b0;
    layer0_outputs(10018) <= not (a xor b);
    layer0_outputs(10019) <= a and b;
    layer0_outputs(10020) <= not b or a;
    layer0_outputs(10021) <= a;
    layer0_outputs(10022) <= not (a xor b);
    layer0_outputs(10023) <= a and b;
    layer0_outputs(10024) <= a;
    layer0_outputs(10025) <= a and not b;
    layer0_outputs(10026) <= a or b;
    layer0_outputs(10027) <= a;
    layer0_outputs(10028) <= a or b;
    layer0_outputs(10029) <= not b;
    layer0_outputs(10030) <= not b;
    layer0_outputs(10031) <= 1'b0;
    layer0_outputs(10032) <= a and not b;
    layer0_outputs(10033) <= a xor b;
    layer0_outputs(10034) <= not b or a;
    layer0_outputs(10035) <= b;
    layer0_outputs(10036) <= a and not b;
    layer0_outputs(10037) <= b and not a;
    layer0_outputs(10038) <= not a;
    layer0_outputs(10039) <= not b;
    layer0_outputs(10040) <= a xor b;
    layer0_outputs(10041) <= not (a xor b);
    layer0_outputs(10042) <= b and not a;
    layer0_outputs(10043) <= b;
    layer0_outputs(10044) <= a or b;
    layer0_outputs(10045) <= b;
    layer0_outputs(10046) <= not b or a;
    layer0_outputs(10047) <= a or b;
    layer0_outputs(10048) <= a or b;
    layer0_outputs(10049) <= b and not a;
    layer0_outputs(10050) <= a;
    layer0_outputs(10051) <= not (a xor b);
    layer0_outputs(10052) <= not a or b;
    layer0_outputs(10053) <= not (a xor b);
    layer0_outputs(10054) <= not (a xor b);
    layer0_outputs(10055) <= not (a or b);
    layer0_outputs(10056) <= b and not a;
    layer0_outputs(10057) <= not (a xor b);
    layer0_outputs(10058) <= not (a or b);
    layer0_outputs(10059) <= b;
    layer0_outputs(10060) <= a and b;
    layer0_outputs(10061) <= not a;
    layer0_outputs(10062) <= 1'b1;
    layer0_outputs(10063) <= not a or b;
    layer0_outputs(10064) <= not (a xor b);
    layer0_outputs(10065) <= a and b;
    layer0_outputs(10066) <= a and b;
    layer0_outputs(10067) <= a xor b;
    layer0_outputs(10068) <= not (a or b);
    layer0_outputs(10069) <= not a or b;
    layer0_outputs(10070) <= not a or b;
    layer0_outputs(10071) <= not (a or b);
    layer0_outputs(10072) <= a and not b;
    layer0_outputs(10073) <= a and b;
    layer0_outputs(10074) <= not a;
    layer0_outputs(10075) <= a or b;
    layer0_outputs(10076) <= not (a or b);
    layer0_outputs(10077) <= not (a xor b);
    layer0_outputs(10078) <= a and b;
    layer0_outputs(10079) <= not (a and b);
    layer0_outputs(10080) <= b;
    layer0_outputs(10081) <= not b or a;
    layer0_outputs(10082) <= b;
    layer0_outputs(10083) <= not b;
    layer0_outputs(10084) <= a;
    layer0_outputs(10085) <= not a;
    layer0_outputs(10086) <= not b;
    layer0_outputs(10087) <= a or b;
    layer0_outputs(10088) <= 1'b1;
    layer0_outputs(10089) <= a or b;
    layer0_outputs(10090) <= not a;
    layer0_outputs(10091) <= not b;
    layer0_outputs(10092) <= a xor b;
    layer0_outputs(10093) <= not (a or b);
    layer0_outputs(10094) <= b and not a;
    layer0_outputs(10095) <= 1'b1;
    layer0_outputs(10096) <= b and not a;
    layer0_outputs(10097) <= not (a xor b);
    layer0_outputs(10098) <= a or b;
    layer0_outputs(10099) <= not b;
    layer0_outputs(10100) <= a xor b;
    layer0_outputs(10101) <= not b or a;
    layer0_outputs(10102) <= a;
    layer0_outputs(10103) <= a and not b;
    layer0_outputs(10104) <= 1'b1;
    layer0_outputs(10105) <= b and not a;
    layer0_outputs(10106) <= a;
    layer0_outputs(10107) <= a and b;
    layer0_outputs(10108) <= not (a xor b);
    layer0_outputs(10109) <= a or b;
    layer0_outputs(10110) <= b and not a;
    layer0_outputs(10111) <= a or b;
    layer0_outputs(10112) <= not a or b;
    layer0_outputs(10113) <= b;
    layer0_outputs(10114) <= a or b;
    layer0_outputs(10115) <= b and not a;
    layer0_outputs(10116) <= 1'b1;
    layer0_outputs(10117) <= a or b;
    layer0_outputs(10118) <= b;
    layer0_outputs(10119) <= a and not b;
    layer0_outputs(10120) <= not (a or b);
    layer0_outputs(10121) <= not (a xor b);
    layer0_outputs(10122) <= not (a or b);
    layer0_outputs(10123) <= not (a xor b);
    layer0_outputs(10124) <= a and not b;
    layer0_outputs(10125) <= b;
    layer0_outputs(10126) <= a;
    layer0_outputs(10127) <= not b or a;
    layer0_outputs(10128) <= not a or b;
    layer0_outputs(10129) <= not (a or b);
    layer0_outputs(10130) <= a;
    layer0_outputs(10131) <= a xor b;
    layer0_outputs(10132) <= a and not b;
    layer0_outputs(10133) <= a or b;
    layer0_outputs(10134) <= not a;
    layer0_outputs(10135) <= b and not a;
    layer0_outputs(10136) <= b and not a;
    layer0_outputs(10137) <= not (a xor b);
    layer0_outputs(10138) <= not b or a;
    layer0_outputs(10139) <= b;
    layer0_outputs(10140) <= not (a or b);
    layer0_outputs(10141) <= not (a xor b);
    layer0_outputs(10142) <= a xor b;
    layer0_outputs(10143) <= b and not a;
    layer0_outputs(10144) <= not (a or b);
    layer0_outputs(10145) <= not b or a;
    layer0_outputs(10146) <= not (a xor b);
    layer0_outputs(10147) <= b;
    layer0_outputs(10148) <= a and not b;
    layer0_outputs(10149) <= not a;
    layer0_outputs(10150) <= not (a xor b);
    layer0_outputs(10151) <= a;
    layer0_outputs(10152) <= not (a xor b);
    layer0_outputs(10153) <= a xor b;
    layer0_outputs(10154) <= a or b;
    layer0_outputs(10155) <= a xor b;
    layer0_outputs(10156) <= not (a xor b);
    layer0_outputs(10157) <= not (a or b);
    layer0_outputs(10158) <= not b or a;
    layer0_outputs(10159) <= a or b;
    layer0_outputs(10160) <= not (a or b);
    layer0_outputs(10161) <= not (a or b);
    layer0_outputs(10162) <= a or b;
    layer0_outputs(10163) <= not (a or b);
    layer0_outputs(10164) <= a;
    layer0_outputs(10165) <= a or b;
    layer0_outputs(10166) <= a or b;
    layer0_outputs(10167) <= a and not b;
    layer0_outputs(10168) <= a xor b;
    layer0_outputs(10169) <= not (a or b);
    layer0_outputs(10170) <= 1'b0;
    layer0_outputs(10171) <= a and b;
    layer0_outputs(10172) <= a xor b;
    layer0_outputs(10173) <= not b or a;
    layer0_outputs(10174) <= a xor b;
    layer0_outputs(10175) <= not (a or b);
    layer0_outputs(10176) <= not a or b;
    layer0_outputs(10177) <= a and not b;
    layer0_outputs(10178) <= a xor b;
    layer0_outputs(10179) <= b and not a;
    layer0_outputs(10180) <= a or b;
    layer0_outputs(10181) <= not (a or b);
    layer0_outputs(10182) <= a or b;
    layer0_outputs(10183) <= a xor b;
    layer0_outputs(10184) <= not a or b;
    layer0_outputs(10185) <= a and b;
    layer0_outputs(10186) <= not a;
    layer0_outputs(10187) <= a xor b;
    layer0_outputs(10188) <= b and not a;
    layer0_outputs(10189) <= 1'b1;
    layer0_outputs(10190) <= a or b;
    layer0_outputs(10191) <= a or b;
    layer0_outputs(10192) <= a or b;
    layer0_outputs(10193) <= a;
    layer0_outputs(10194) <= a;
    layer0_outputs(10195) <= a or b;
    layer0_outputs(10196) <= not (a xor b);
    layer0_outputs(10197) <= a xor b;
    layer0_outputs(10198) <= a and not b;
    layer0_outputs(10199) <= a;
    layer0_outputs(10200) <= not b;
    layer0_outputs(10201) <= not a;
    layer0_outputs(10202) <= not (a or b);
    layer0_outputs(10203) <= not (a or b);
    layer0_outputs(10204) <= b and not a;
    layer0_outputs(10205) <= 1'b0;
    layer0_outputs(10206) <= 1'b0;
    layer0_outputs(10207) <= 1'b1;
    layer0_outputs(10208) <= not (a and b);
    layer0_outputs(10209) <= not b;
    layer0_outputs(10210) <= not (a or b);
    layer0_outputs(10211) <= not a or b;
    layer0_outputs(10212) <= 1'b0;
    layer0_outputs(10213) <= not b or a;
    layer0_outputs(10214) <= not (a xor b);
    layer0_outputs(10215) <= not a or b;
    layer0_outputs(10216) <= not (a or b);
    layer0_outputs(10217) <= 1'b1;
    layer0_outputs(10218) <= not b;
    layer0_outputs(10219) <= not (a or b);
    layer0_outputs(10220) <= a and not b;
    layer0_outputs(10221) <= a and not b;
    layer0_outputs(10222) <= not b or a;
    layer0_outputs(10223) <= not a;
    layer0_outputs(10224) <= a or b;
    layer0_outputs(10225) <= a;
    layer0_outputs(10226) <= not (a or b);
    layer0_outputs(10227) <= not (a xor b);
    layer0_outputs(10228) <= a and not b;
    layer0_outputs(10229) <= a;
    layer0_outputs(10230) <= a and not b;
    layer0_outputs(10231) <= not (a and b);
    layer0_outputs(10232) <= not b;
    layer0_outputs(10233) <= a xor b;
    layer0_outputs(10234) <= not (a xor b);
    layer0_outputs(10235) <= not b or a;
    layer0_outputs(10236) <= not (a and b);
    layer0_outputs(10237) <= 1'b1;
    layer0_outputs(10238) <= b and not a;
    layer0_outputs(10239) <= b and not a;
    layer0_outputs(10240) <= not b;
    layer0_outputs(10241) <= not a;
    layer0_outputs(10242) <= a xor b;
    layer0_outputs(10243) <= b and not a;
    layer0_outputs(10244) <= b;
    layer0_outputs(10245) <= a xor b;
    layer0_outputs(10246) <= a or b;
    layer0_outputs(10247) <= not b or a;
    layer0_outputs(10248) <= not a or b;
    layer0_outputs(10249) <= a xor b;
    layer0_outputs(10250) <= a and not b;
    layer0_outputs(10251) <= a and b;
    layer0_outputs(10252) <= a;
    layer0_outputs(10253) <= not b;
    layer0_outputs(10254) <= b and not a;
    layer0_outputs(10255) <= a or b;
    layer0_outputs(10256) <= a xor b;
    layer0_outputs(10257) <= b;
    layer0_outputs(10258) <= a or b;
    layer0_outputs(10259) <= not (a xor b);
    layer0_outputs(10260) <= b;
    layer0_outputs(10261) <= a and not b;
    layer0_outputs(10262) <= not a or b;
    layer0_outputs(10263) <= a;
    layer0_outputs(10264) <= b and not a;
    layer0_outputs(10265) <= not a;
    layer0_outputs(10266) <= not (a and b);
    layer0_outputs(10267) <= not a;
    layer0_outputs(10268) <= not a;
    layer0_outputs(10269) <= not (a xor b);
    layer0_outputs(10270) <= not (a xor b);
    layer0_outputs(10271) <= b and not a;
    layer0_outputs(10272) <= not (a xor b);
    layer0_outputs(10273) <= not (a or b);
    layer0_outputs(10274) <= a or b;
    layer0_outputs(10275) <= not (a xor b);
    layer0_outputs(10276) <= a xor b;
    layer0_outputs(10277) <= 1'b1;
    layer0_outputs(10278) <= b and not a;
    layer0_outputs(10279) <= a or b;
    layer0_outputs(10280) <= not a;
    layer0_outputs(10281) <= not a or b;
    layer0_outputs(10282) <= a and b;
    layer0_outputs(10283) <= not (a xor b);
    layer0_outputs(10284) <= not (a xor b);
    layer0_outputs(10285) <= not b or a;
    layer0_outputs(10286) <= b and not a;
    layer0_outputs(10287) <= not (a and b);
    layer0_outputs(10288) <= a xor b;
    layer0_outputs(10289) <= 1'b1;
    layer0_outputs(10290) <= b;
    layer0_outputs(10291) <= not (a and b);
    layer0_outputs(10292) <= not a;
    layer0_outputs(10293) <= b and not a;
    layer0_outputs(10294) <= a and b;
    layer0_outputs(10295) <= a;
    layer0_outputs(10296) <= not (a or b);
    layer0_outputs(10297) <= not b;
    layer0_outputs(10298) <= not (a xor b);
    layer0_outputs(10299) <= not (a or b);
    layer0_outputs(10300) <= a or b;
    layer0_outputs(10301) <= a or b;
    layer0_outputs(10302) <= a or b;
    layer0_outputs(10303) <= 1'b1;
    layer0_outputs(10304) <= not (a xor b);
    layer0_outputs(10305) <= a or b;
    layer0_outputs(10306) <= not (a or b);
    layer0_outputs(10307) <= not (a or b);
    layer0_outputs(10308) <= not b or a;
    layer0_outputs(10309) <= b and not a;
    layer0_outputs(10310) <= not a or b;
    layer0_outputs(10311) <= not (a xor b);
    layer0_outputs(10312) <= a or b;
    layer0_outputs(10313) <= not (a or b);
    layer0_outputs(10314) <= not a;
    layer0_outputs(10315) <= not a or b;
    layer0_outputs(10316) <= not (a or b);
    layer0_outputs(10317) <= a xor b;
    layer0_outputs(10318) <= not (a xor b);
    layer0_outputs(10319) <= not (a or b);
    layer0_outputs(10320) <= not a;
    layer0_outputs(10321) <= not a or b;
    layer0_outputs(10322) <= a or b;
    layer0_outputs(10323) <= not b;
    layer0_outputs(10324) <= b and not a;
    layer0_outputs(10325) <= not (a and b);
    layer0_outputs(10326) <= b and not a;
    layer0_outputs(10327) <= b;
    layer0_outputs(10328) <= not (a or b);
    layer0_outputs(10329) <= b;
    layer0_outputs(10330) <= a xor b;
    layer0_outputs(10331) <= not (a and b);
    layer0_outputs(10332) <= a or b;
    layer0_outputs(10333) <= not (a xor b);
    layer0_outputs(10334) <= b;
    layer0_outputs(10335) <= 1'b1;
    layer0_outputs(10336) <= b and not a;
    layer0_outputs(10337) <= a xor b;
    layer0_outputs(10338) <= a and not b;
    layer0_outputs(10339) <= b and not a;
    layer0_outputs(10340) <= not b or a;
    layer0_outputs(10341) <= not a or b;
    layer0_outputs(10342) <= not (a or b);
    layer0_outputs(10343) <= a xor b;
    layer0_outputs(10344) <= a;
    layer0_outputs(10345) <= not a;
    layer0_outputs(10346) <= not (a xor b);
    layer0_outputs(10347) <= 1'b0;
    layer0_outputs(10348) <= not (a or b);
    layer0_outputs(10349) <= not b;
    layer0_outputs(10350) <= a xor b;
    layer0_outputs(10351) <= a and b;
    layer0_outputs(10352) <= b;
    layer0_outputs(10353) <= a and b;
    layer0_outputs(10354) <= a and not b;
    layer0_outputs(10355) <= not b or a;
    layer0_outputs(10356) <= 1'b1;
    layer0_outputs(10357) <= not b or a;
    layer0_outputs(10358) <= not b;
    layer0_outputs(10359) <= a;
    layer0_outputs(10360) <= a or b;
    layer0_outputs(10361) <= not (a xor b);
    layer0_outputs(10362) <= not b or a;
    layer0_outputs(10363) <= b;
    layer0_outputs(10364) <= not (a and b);
    layer0_outputs(10365) <= not a or b;
    layer0_outputs(10366) <= a xor b;
    layer0_outputs(10367) <= not b;
    layer0_outputs(10368) <= a or b;
    layer0_outputs(10369) <= 1'b1;
    layer0_outputs(10370) <= b and not a;
    layer0_outputs(10371) <= not b or a;
    layer0_outputs(10372) <= not a or b;
    layer0_outputs(10373) <= a;
    layer0_outputs(10374) <= 1'b0;
    layer0_outputs(10375) <= b and not a;
    layer0_outputs(10376) <= a xor b;
    layer0_outputs(10377) <= a or b;
    layer0_outputs(10378) <= not (a or b);
    layer0_outputs(10379) <= a or b;
    layer0_outputs(10380) <= not a;
    layer0_outputs(10381) <= not (a or b);
    layer0_outputs(10382) <= b;
    layer0_outputs(10383) <= not (a xor b);
    layer0_outputs(10384) <= not a;
    layer0_outputs(10385) <= a or b;
    layer0_outputs(10386) <= b and not a;
    layer0_outputs(10387) <= not a or b;
    layer0_outputs(10388) <= not b;
    layer0_outputs(10389) <= a xor b;
    layer0_outputs(10390) <= a xor b;
    layer0_outputs(10391) <= not b;
    layer0_outputs(10392) <= not b or a;
    layer0_outputs(10393) <= b;
    layer0_outputs(10394) <= a;
    layer0_outputs(10395) <= b;
    layer0_outputs(10396) <= not (a or b);
    layer0_outputs(10397) <= a or b;
    layer0_outputs(10398) <= a xor b;
    layer0_outputs(10399) <= 1'b0;
    layer0_outputs(10400) <= b and not a;
    layer0_outputs(10401) <= not b or a;
    layer0_outputs(10402) <= not a or b;
    layer0_outputs(10403) <= not a or b;
    layer0_outputs(10404) <= not a;
    layer0_outputs(10405) <= not a or b;
    layer0_outputs(10406) <= a or b;
    layer0_outputs(10407) <= a and not b;
    layer0_outputs(10408) <= not b or a;
    layer0_outputs(10409) <= a and not b;
    layer0_outputs(10410) <= a or b;
    layer0_outputs(10411) <= a;
    layer0_outputs(10412) <= a and not b;
    layer0_outputs(10413) <= a and b;
    layer0_outputs(10414) <= not (a or b);
    layer0_outputs(10415) <= not a or b;
    layer0_outputs(10416) <= a and not b;
    layer0_outputs(10417) <= a or b;
    layer0_outputs(10418) <= a and b;
    layer0_outputs(10419) <= not a or b;
    layer0_outputs(10420) <= a and b;
    layer0_outputs(10421) <= not b;
    layer0_outputs(10422) <= a or b;
    layer0_outputs(10423) <= a xor b;
    layer0_outputs(10424) <= not (a xor b);
    layer0_outputs(10425) <= a and not b;
    layer0_outputs(10426) <= not b;
    layer0_outputs(10427) <= a xor b;
    layer0_outputs(10428) <= not (a xor b);
    layer0_outputs(10429) <= not (a and b);
    layer0_outputs(10430) <= not b;
    layer0_outputs(10431) <= b;
    layer0_outputs(10432) <= not (a and b);
    layer0_outputs(10433) <= b;
    layer0_outputs(10434) <= a or b;
    layer0_outputs(10435) <= not b;
    layer0_outputs(10436) <= b;
    layer0_outputs(10437) <= not b or a;
    layer0_outputs(10438) <= 1'b1;
    layer0_outputs(10439) <= a xor b;
    layer0_outputs(10440) <= not (a xor b);
    layer0_outputs(10441) <= a;
    layer0_outputs(10442) <= not (a and b);
    layer0_outputs(10443) <= a xor b;
    layer0_outputs(10444) <= a and not b;
    layer0_outputs(10445) <= not a or b;
    layer0_outputs(10446) <= not (a and b);
    layer0_outputs(10447) <= not a or b;
    layer0_outputs(10448) <= not (a or b);
    layer0_outputs(10449) <= not (a or b);
    layer0_outputs(10450) <= a or b;
    layer0_outputs(10451) <= not (a or b);
    layer0_outputs(10452) <= b;
    layer0_outputs(10453) <= not (a or b);
    layer0_outputs(10454) <= a and not b;
    layer0_outputs(10455) <= not b;
    layer0_outputs(10456) <= b and not a;
    layer0_outputs(10457) <= a or b;
    layer0_outputs(10458) <= not (a xor b);
    layer0_outputs(10459) <= a;
    layer0_outputs(10460) <= a and not b;
    layer0_outputs(10461) <= a and not b;
    layer0_outputs(10462) <= a;
    layer0_outputs(10463) <= not (a xor b);
    layer0_outputs(10464) <= not b;
    layer0_outputs(10465) <= not (a or b);
    layer0_outputs(10466) <= a xor b;
    layer0_outputs(10467) <= not b or a;
    layer0_outputs(10468) <= 1'b0;
    layer0_outputs(10469) <= 1'b0;
    layer0_outputs(10470) <= b and not a;
    layer0_outputs(10471) <= not (a xor b);
    layer0_outputs(10472) <= not (a or b);
    layer0_outputs(10473) <= not b;
    layer0_outputs(10474) <= not (a xor b);
    layer0_outputs(10475) <= 1'b1;
    layer0_outputs(10476) <= b;
    layer0_outputs(10477) <= not (a xor b);
    layer0_outputs(10478) <= not a or b;
    layer0_outputs(10479) <= not (a xor b);
    layer0_outputs(10480) <= b and not a;
    layer0_outputs(10481) <= b and not a;
    layer0_outputs(10482) <= not (a xor b);
    layer0_outputs(10483) <= not (a or b);
    layer0_outputs(10484) <= a xor b;
    layer0_outputs(10485) <= not (a or b);
    layer0_outputs(10486) <= not (a or b);
    layer0_outputs(10487) <= not a;
    layer0_outputs(10488) <= not (a or b);
    layer0_outputs(10489) <= not (a xor b);
    layer0_outputs(10490) <= a;
    layer0_outputs(10491) <= a xor b;
    layer0_outputs(10492) <= not a or b;
    layer0_outputs(10493) <= a or b;
    layer0_outputs(10494) <= not (a or b);
    layer0_outputs(10495) <= not a or b;
    layer0_outputs(10496) <= not (a xor b);
    layer0_outputs(10497) <= not a;
    layer0_outputs(10498) <= not (a xor b);
    layer0_outputs(10499) <= a and not b;
    layer0_outputs(10500) <= b and not a;
    layer0_outputs(10501) <= a xor b;
    layer0_outputs(10502) <= a or b;
    layer0_outputs(10503) <= not b;
    layer0_outputs(10504) <= b and not a;
    layer0_outputs(10505) <= not a or b;
    layer0_outputs(10506) <= not b or a;
    layer0_outputs(10507) <= not a or b;
    layer0_outputs(10508) <= a xor b;
    layer0_outputs(10509) <= a xor b;
    layer0_outputs(10510) <= a xor b;
    layer0_outputs(10511) <= b and not a;
    layer0_outputs(10512) <= a and not b;
    layer0_outputs(10513) <= not (a or b);
    layer0_outputs(10514) <= a xor b;
    layer0_outputs(10515) <= not (a or b);
    layer0_outputs(10516) <= a and b;
    layer0_outputs(10517) <= not (a xor b);
    layer0_outputs(10518) <= a or b;
    layer0_outputs(10519) <= not a;
    layer0_outputs(10520) <= not (a xor b);
    layer0_outputs(10521) <= a and b;
    layer0_outputs(10522) <= not (a or b);
    layer0_outputs(10523) <= b;
    layer0_outputs(10524) <= a;
    layer0_outputs(10525) <= not (a xor b);
    layer0_outputs(10526) <= not a or b;
    layer0_outputs(10527) <= b;
    layer0_outputs(10528) <= not (a xor b);
    layer0_outputs(10529) <= not a;
    layer0_outputs(10530) <= not (a xor b);
    layer0_outputs(10531) <= not a;
    layer0_outputs(10532) <= a;
    layer0_outputs(10533) <= 1'b1;
    layer0_outputs(10534) <= not a or b;
    layer0_outputs(10535) <= not (a or b);
    layer0_outputs(10536) <= b;
    layer0_outputs(10537) <= not (a or b);
    layer0_outputs(10538) <= a xor b;
    layer0_outputs(10539) <= a;
    layer0_outputs(10540) <= a;
    layer0_outputs(10541) <= a and b;
    layer0_outputs(10542) <= a and b;
    layer0_outputs(10543) <= 1'b0;
    layer0_outputs(10544) <= b;
    layer0_outputs(10545) <= a xor b;
    layer0_outputs(10546) <= not a or b;
    layer0_outputs(10547) <= a or b;
    layer0_outputs(10548) <= a or b;
    layer0_outputs(10549) <= a or b;
    layer0_outputs(10550) <= a xor b;
    layer0_outputs(10551) <= not b;
    layer0_outputs(10552) <= b;
    layer0_outputs(10553) <= a and b;
    layer0_outputs(10554) <= not (a xor b);
    layer0_outputs(10555) <= a;
    layer0_outputs(10556) <= not b or a;
    layer0_outputs(10557) <= b and not a;
    layer0_outputs(10558) <= 1'b1;
    layer0_outputs(10559) <= not (a or b);
    layer0_outputs(10560) <= a xor b;
    layer0_outputs(10561) <= not (a xor b);
    layer0_outputs(10562) <= a and not b;
    layer0_outputs(10563) <= not (a and b);
    layer0_outputs(10564) <= not b;
    layer0_outputs(10565) <= a or b;
    layer0_outputs(10566) <= not b or a;
    layer0_outputs(10567) <= not a or b;
    layer0_outputs(10568) <= a xor b;
    layer0_outputs(10569) <= a or b;
    layer0_outputs(10570) <= b;
    layer0_outputs(10571) <= not b or a;
    layer0_outputs(10572) <= not (a xor b);
    layer0_outputs(10573) <= b;
    layer0_outputs(10574) <= a and not b;
    layer0_outputs(10575) <= not (a or b);
    layer0_outputs(10576) <= a or b;
    layer0_outputs(10577) <= a or b;
    layer0_outputs(10578) <= not a;
    layer0_outputs(10579) <= not b or a;
    layer0_outputs(10580) <= not b;
    layer0_outputs(10581) <= not (a xor b);
    layer0_outputs(10582) <= not (a xor b);
    layer0_outputs(10583) <= not b or a;
    layer0_outputs(10584) <= not b or a;
    layer0_outputs(10585) <= b;
    layer0_outputs(10586) <= 1'b0;
    layer0_outputs(10587) <= a xor b;
    layer0_outputs(10588) <= not a or b;
    layer0_outputs(10589) <= a;
    layer0_outputs(10590) <= not (a and b);
    layer0_outputs(10591) <= not (a xor b);
    layer0_outputs(10592) <= a;
    layer0_outputs(10593) <= a xor b;
    layer0_outputs(10594) <= not a;
    layer0_outputs(10595) <= not (a or b);
    layer0_outputs(10596) <= a;
    layer0_outputs(10597) <= a or b;
    layer0_outputs(10598) <= not a;
    layer0_outputs(10599) <= not (a and b);
    layer0_outputs(10600) <= not (a xor b);
    layer0_outputs(10601) <= a or b;
    layer0_outputs(10602) <= not (a xor b);
    layer0_outputs(10603) <= not b or a;
    layer0_outputs(10604) <= a and not b;
    layer0_outputs(10605) <= 1'b0;
    layer0_outputs(10606) <= b and not a;
    layer0_outputs(10607) <= not (a xor b);
    layer0_outputs(10608) <= a;
    layer0_outputs(10609) <= b and not a;
    layer0_outputs(10610) <= a;
    layer0_outputs(10611) <= a xor b;
    layer0_outputs(10612) <= b and not a;
    layer0_outputs(10613) <= a;
    layer0_outputs(10614) <= a;
    layer0_outputs(10615) <= b;
    layer0_outputs(10616) <= not (a xor b);
    layer0_outputs(10617) <= a and not b;
    layer0_outputs(10618) <= not (a and b);
    layer0_outputs(10619) <= a xor b;
    layer0_outputs(10620) <= a and not b;
    layer0_outputs(10621) <= b;
    layer0_outputs(10622) <= b;
    layer0_outputs(10623) <= not (a xor b);
    layer0_outputs(10624) <= not (a xor b);
    layer0_outputs(10625) <= not a;
    layer0_outputs(10626) <= a or b;
    layer0_outputs(10627) <= a or b;
    layer0_outputs(10628) <= a xor b;
    layer0_outputs(10629) <= not (a xor b);
    layer0_outputs(10630) <= b and not a;
    layer0_outputs(10631) <= b and not a;
    layer0_outputs(10632) <= a xor b;
    layer0_outputs(10633) <= a or b;
    layer0_outputs(10634) <= a or b;
    layer0_outputs(10635) <= not b;
    layer0_outputs(10636) <= not a or b;
    layer0_outputs(10637) <= not (a or b);
    layer0_outputs(10638) <= a and not b;
    layer0_outputs(10639) <= not (a and b);
    layer0_outputs(10640) <= not a;
    layer0_outputs(10641) <= not (a or b);
    layer0_outputs(10642) <= not b or a;
    layer0_outputs(10643) <= a and b;
    layer0_outputs(10644) <= not a or b;
    layer0_outputs(10645) <= a and not b;
    layer0_outputs(10646) <= a xor b;
    layer0_outputs(10647) <= a;
    layer0_outputs(10648) <= b;
    layer0_outputs(10649) <= not b;
    layer0_outputs(10650) <= a and not b;
    layer0_outputs(10651) <= b;
    layer0_outputs(10652) <= b;
    layer0_outputs(10653) <= b;
    layer0_outputs(10654) <= not a or b;
    layer0_outputs(10655) <= not a;
    layer0_outputs(10656) <= not (a or b);
    layer0_outputs(10657) <= not (a xor b);
    layer0_outputs(10658) <= not (a and b);
    layer0_outputs(10659) <= not (a or b);
    layer0_outputs(10660) <= not (a or b);
    layer0_outputs(10661) <= not a or b;
    layer0_outputs(10662) <= a and not b;
    layer0_outputs(10663) <= a xor b;
    layer0_outputs(10664) <= a and b;
    layer0_outputs(10665) <= not (a or b);
    layer0_outputs(10666) <= b and not a;
    layer0_outputs(10667) <= not (a xor b);
    layer0_outputs(10668) <= a xor b;
    layer0_outputs(10669) <= not b;
    layer0_outputs(10670) <= not b;
    layer0_outputs(10671) <= 1'b1;
    layer0_outputs(10672) <= a;
    layer0_outputs(10673) <= not a;
    layer0_outputs(10674) <= not (a or b);
    layer0_outputs(10675) <= not (a xor b);
    layer0_outputs(10676) <= not a;
    layer0_outputs(10677) <= not a;
    layer0_outputs(10678) <= b;
    layer0_outputs(10679) <= not b;
    layer0_outputs(10680) <= a or b;
    layer0_outputs(10681) <= a xor b;
    layer0_outputs(10682) <= a;
    layer0_outputs(10683) <= b;
    layer0_outputs(10684) <= not (a or b);
    layer0_outputs(10685) <= a xor b;
    layer0_outputs(10686) <= not (a or b);
    layer0_outputs(10687) <= a;
    layer0_outputs(10688) <= b and not a;
    layer0_outputs(10689) <= not (a xor b);
    layer0_outputs(10690) <= not (a or b);
    layer0_outputs(10691) <= not a or b;
    layer0_outputs(10692) <= b;
    layer0_outputs(10693) <= a;
    layer0_outputs(10694) <= b;
    layer0_outputs(10695) <= b and not a;
    layer0_outputs(10696) <= not (a and b);
    layer0_outputs(10697) <= not b;
    layer0_outputs(10698) <= 1'b1;
    layer0_outputs(10699) <= a and b;
    layer0_outputs(10700) <= not a;
    layer0_outputs(10701) <= not b or a;
    layer0_outputs(10702) <= a or b;
    layer0_outputs(10703) <= a or b;
    layer0_outputs(10704) <= a or b;
    layer0_outputs(10705) <= not b;
    layer0_outputs(10706) <= not b;
    layer0_outputs(10707) <= not b;
    layer0_outputs(10708) <= not b;
    layer0_outputs(10709) <= a or b;
    layer0_outputs(10710) <= 1'b0;
    layer0_outputs(10711) <= a or b;
    layer0_outputs(10712) <= not (a or b);
    layer0_outputs(10713) <= not (a or b);
    layer0_outputs(10714) <= a;
    layer0_outputs(10715) <= not (a xor b);
    layer0_outputs(10716) <= not a;
    layer0_outputs(10717) <= not a or b;
    layer0_outputs(10718) <= a xor b;
    layer0_outputs(10719) <= a xor b;
    layer0_outputs(10720) <= a or b;
    layer0_outputs(10721) <= not b;
    layer0_outputs(10722) <= not (a or b);
    layer0_outputs(10723) <= not (a or b);
    layer0_outputs(10724) <= not (a xor b);
    layer0_outputs(10725) <= a;
    layer0_outputs(10726) <= a or b;
    layer0_outputs(10727) <= a or b;
    layer0_outputs(10728) <= b and not a;
    layer0_outputs(10729) <= not (a or b);
    layer0_outputs(10730) <= a and b;
    layer0_outputs(10731) <= not (a or b);
    layer0_outputs(10732) <= not (a xor b);
    layer0_outputs(10733) <= not a or b;
    layer0_outputs(10734) <= not a;
    layer0_outputs(10735) <= not b or a;
    layer0_outputs(10736) <= b and not a;
    layer0_outputs(10737) <= a or b;
    layer0_outputs(10738) <= b and not a;
    layer0_outputs(10739) <= not (a or b);
    layer0_outputs(10740) <= not a or b;
    layer0_outputs(10741) <= not b or a;
    layer0_outputs(10742) <= not a or b;
    layer0_outputs(10743) <= a xor b;
    layer0_outputs(10744) <= not b;
    layer0_outputs(10745) <= 1'b1;
    layer0_outputs(10746) <= not b or a;
    layer0_outputs(10747) <= a xor b;
    layer0_outputs(10748) <= not a;
    layer0_outputs(10749) <= not (a and b);
    layer0_outputs(10750) <= b and not a;
    layer0_outputs(10751) <= not a;
    layer0_outputs(10752) <= a or b;
    layer0_outputs(10753) <= not a;
    layer0_outputs(10754) <= b and not a;
    layer0_outputs(10755) <= a and not b;
    layer0_outputs(10756) <= not (a and b);
    layer0_outputs(10757) <= 1'b0;
    layer0_outputs(10758) <= a or b;
    layer0_outputs(10759) <= a or b;
    layer0_outputs(10760) <= not b;
    layer0_outputs(10761) <= not (a xor b);
    layer0_outputs(10762) <= not a;
    layer0_outputs(10763) <= a and not b;
    layer0_outputs(10764) <= not (a xor b);
    layer0_outputs(10765) <= b;
    layer0_outputs(10766) <= a;
    layer0_outputs(10767) <= a or b;
    layer0_outputs(10768) <= a and not b;
    layer0_outputs(10769) <= 1'b1;
    layer0_outputs(10770) <= a;
    layer0_outputs(10771) <= not a or b;
    layer0_outputs(10772) <= not b;
    layer0_outputs(10773) <= not b;
    layer0_outputs(10774) <= not a or b;
    layer0_outputs(10775) <= not a;
    layer0_outputs(10776) <= a xor b;
    layer0_outputs(10777) <= not a;
    layer0_outputs(10778) <= not (a xor b);
    layer0_outputs(10779) <= not b;
    layer0_outputs(10780) <= a and not b;
    layer0_outputs(10781) <= a xor b;
    layer0_outputs(10782) <= not a;
    layer0_outputs(10783) <= not (a or b);
    layer0_outputs(10784) <= a xor b;
    layer0_outputs(10785) <= not (a or b);
    layer0_outputs(10786) <= not (a xor b);
    layer0_outputs(10787) <= b;
    layer0_outputs(10788) <= a xor b;
    layer0_outputs(10789) <= 1'b0;
    layer0_outputs(10790) <= a and b;
    layer0_outputs(10791) <= b and not a;
    layer0_outputs(10792) <= a or b;
    layer0_outputs(10793) <= a;
    layer0_outputs(10794) <= a;
    layer0_outputs(10795) <= a or b;
    layer0_outputs(10796) <= b and not a;
    layer0_outputs(10797) <= not b;
    layer0_outputs(10798) <= not a or b;
    layer0_outputs(10799) <= b;
    layer0_outputs(10800) <= not b or a;
    layer0_outputs(10801) <= a or b;
    layer0_outputs(10802) <= not (a xor b);
    layer0_outputs(10803) <= a or b;
    layer0_outputs(10804) <= a;
    layer0_outputs(10805) <= b;
    layer0_outputs(10806) <= b and not a;
    layer0_outputs(10807) <= not (a xor b);
    layer0_outputs(10808) <= a and not b;
    layer0_outputs(10809) <= a and not b;
    layer0_outputs(10810) <= a xor b;
    layer0_outputs(10811) <= a or b;
    layer0_outputs(10812) <= not (a xor b);
    layer0_outputs(10813) <= not b;
    layer0_outputs(10814) <= not b;
    layer0_outputs(10815) <= b and not a;
    layer0_outputs(10816) <= not a or b;
    layer0_outputs(10817) <= not b;
    layer0_outputs(10818) <= b and not a;
    layer0_outputs(10819) <= not b or a;
    layer0_outputs(10820) <= not (a xor b);
    layer0_outputs(10821) <= b and not a;
    layer0_outputs(10822) <= a xor b;
    layer0_outputs(10823) <= a xor b;
    layer0_outputs(10824) <= not b;
    layer0_outputs(10825) <= not b;
    layer0_outputs(10826) <= not (a or b);
    layer0_outputs(10827) <= not (a xor b);
    layer0_outputs(10828) <= not a;
    layer0_outputs(10829) <= not a;
    layer0_outputs(10830) <= a;
    layer0_outputs(10831) <= not a or b;
    layer0_outputs(10832) <= a or b;
    layer0_outputs(10833) <= not (a and b);
    layer0_outputs(10834) <= not a or b;
    layer0_outputs(10835) <= b and not a;
    layer0_outputs(10836) <= b;
    layer0_outputs(10837) <= not a;
    layer0_outputs(10838) <= 1'b1;
    layer0_outputs(10839) <= a or b;
    layer0_outputs(10840) <= not b;
    layer0_outputs(10841) <= not b or a;
    layer0_outputs(10842) <= a xor b;
    layer0_outputs(10843) <= b;
    layer0_outputs(10844) <= b and not a;
    layer0_outputs(10845) <= not (a or b);
    layer0_outputs(10846) <= not b or a;
    layer0_outputs(10847) <= b and not a;
    layer0_outputs(10848) <= not a or b;
    layer0_outputs(10849) <= not a;
    layer0_outputs(10850) <= a;
    layer0_outputs(10851) <= not a;
    layer0_outputs(10852) <= a or b;
    layer0_outputs(10853) <= not a or b;
    layer0_outputs(10854) <= not (a or b);
    layer0_outputs(10855) <= not (a or b);
    layer0_outputs(10856) <= not (a and b);
    layer0_outputs(10857) <= b;
    layer0_outputs(10858) <= not (a or b);
    layer0_outputs(10859) <= not a or b;
    layer0_outputs(10860) <= not (a or b);
    layer0_outputs(10861) <= not b or a;
    layer0_outputs(10862) <= b and not a;
    layer0_outputs(10863) <= not b or a;
    layer0_outputs(10864) <= 1'b0;
    layer0_outputs(10865) <= a and b;
    layer0_outputs(10866) <= a xor b;
    layer0_outputs(10867) <= not (a and b);
    layer0_outputs(10868) <= b;
    layer0_outputs(10869) <= b and not a;
    layer0_outputs(10870) <= not (a or b);
    layer0_outputs(10871) <= not b or a;
    layer0_outputs(10872) <= a and b;
    layer0_outputs(10873) <= b;
    layer0_outputs(10874) <= a or b;
    layer0_outputs(10875) <= not b or a;
    layer0_outputs(10876) <= not (a or b);
    layer0_outputs(10877) <= b;
    layer0_outputs(10878) <= a xor b;
    layer0_outputs(10879) <= a and not b;
    layer0_outputs(10880) <= not a;
    layer0_outputs(10881) <= not b;
    layer0_outputs(10882) <= a;
    layer0_outputs(10883) <= a or b;
    layer0_outputs(10884) <= b;
    layer0_outputs(10885) <= b and not a;
    layer0_outputs(10886) <= a;
    layer0_outputs(10887) <= b and not a;
    layer0_outputs(10888) <= a;
    layer0_outputs(10889) <= a xor b;
    layer0_outputs(10890) <= not a or b;
    layer0_outputs(10891) <= not (a or b);
    layer0_outputs(10892) <= not (a or b);
    layer0_outputs(10893) <= not a;
    layer0_outputs(10894) <= b;
    layer0_outputs(10895) <= not (a or b);
    layer0_outputs(10896) <= a and not b;
    layer0_outputs(10897) <= not (a xor b);
    layer0_outputs(10898) <= not b or a;
    layer0_outputs(10899) <= not (a xor b);
    layer0_outputs(10900) <= a xor b;
    layer0_outputs(10901) <= 1'b1;
    layer0_outputs(10902) <= not b;
    layer0_outputs(10903) <= not a;
    layer0_outputs(10904) <= a or b;
    layer0_outputs(10905) <= a xor b;
    layer0_outputs(10906) <= not b or a;
    layer0_outputs(10907) <= not (a or b);
    layer0_outputs(10908) <= not (a or b);
    layer0_outputs(10909) <= a and not b;
    layer0_outputs(10910) <= a or b;
    layer0_outputs(10911) <= not a;
    layer0_outputs(10912) <= 1'b1;
    layer0_outputs(10913) <= not (a or b);
    layer0_outputs(10914) <= b;
    layer0_outputs(10915) <= not b or a;
    layer0_outputs(10916) <= not a or b;
    layer0_outputs(10917) <= not a or b;
    layer0_outputs(10918) <= not (a or b);
    layer0_outputs(10919) <= not (a xor b);
    layer0_outputs(10920) <= not a or b;
    layer0_outputs(10921) <= a;
    layer0_outputs(10922) <= a;
    layer0_outputs(10923) <= not a or b;
    layer0_outputs(10924) <= a or b;
    layer0_outputs(10925) <= a xor b;
    layer0_outputs(10926) <= a;
    layer0_outputs(10927) <= b;
    layer0_outputs(10928) <= b and not a;
    layer0_outputs(10929) <= not b or a;
    layer0_outputs(10930) <= not b;
    layer0_outputs(10931) <= a and not b;
    layer0_outputs(10932) <= not a;
    layer0_outputs(10933) <= a;
    layer0_outputs(10934) <= not (a xor b);
    layer0_outputs(10935) <= a or b;
    layer0_outputs(10936) <= not b;
    layer0_outputs(10937) <= not (a xor b);
    layer0_outputs(10938) <= b;
    layer0_outputs(10939) <= not (a or b);
    layer0_outputs(10940) <= not a;
    layer0_outputs(10941) <= a;
    layer0_outputs(10942) <= a xor b;
    layer0_outputs(10943) <= a or b;
    layer0_outputs(10944) <= not b or a;
    layer0_outputs(10945) <= a xor b;
    layer0_outputs(10946) <= a or b;
    layer0_outputs(10947) <= not (a or b);
    layer0_outputs(10948) <= a xor b;
    layer0_outputs(10949) <= not b;
    layer0_outputs(10950) <= not a;
    layer0_outputs(10951) <= b and not a;
    layer0_outputs(10952) <= not b;
    layer0_outputs(10953) <= not (a and b);
    layer0_outputs(10954) <= not a;
    layer0_outputs(10955) <= not (a or b);
    layer0_outputs(10956) <= a or b;
    layer0_outputs(10957) <= not (a or b);
    layer0_outputs(10958) <= a and not b;
    layer0_outputs(10959) <= a and not b;
    layer0_outputs(10960) <= not (a xor b);
    layer0_outputs(10961) <= a or b;
    layer0_outputs(10962) <= a or b;
    layer0_outputs(10963) <= not a;
    layer0_outputs(10964) <= a and b;
    layer0_outputs(10965) <= not a;
    layer0_outputs(10966) <= not a or b;
    layer0_outputs(10967) <= a or b;
    layer0_outputs(10968) <= a or b;
    layer0_outputs(10969) <= not a or b;
    layer0_outputs(10970) <= not b or a;
    layer0_outputs(10971) <= not b or a;
    layer0_outputs(10972) <= not (a xor b);
    layer0_outputs(10973) <= a;
    layer0_outputs(10974) <= a xor b;
    layer0_outputs(10975) <= not a;
    layer0_outputs(10976) <= not (a and b);
    layer0_outputs(10977) <= a;
    layer0_outputs(10978) <= not a;
    layer0_outputs(10979) <= a or b;
    layer0_outputs(10980) <= not b;
    layer0_outputs(10981) <= not (a or b);
    layer0_outputs(10982) <= not (a or b);
    layer0_outputs(10983) <= not (a xor b);
    layer0_outputs(10984) <= not a or b;
    layer0_outputs(10985) <= a;
    layer0_outputs(10986) <= b and not a;
    layer0_outputs(10987) <= not (a or b);
    layer0_outputs(10988) <= not (a or b);
    layer0_outputs(10989) <= 1'b1;
    layer0_outputs(10990) <= a xor b;
    layer0_outputs(10991) <= not a or b;
    layer0_outputs(10992) <= a and b;
    layer0_outputs(10993) <= a or b;
    layer0_outputs(10994) <= a and not b;
    layer0_outputs(10995) <= not a or b;
    layer0_outputs(10996) <= 1'b1;
    layer0_outputs(10997) <= a or b;
    layer0_outputs(10998) <= not (a xor b);
    layer0_outputs(10999) <= a;
    layer0_outputs(11000) <= not b or a;
    layer0_outputs(11001) <= a;
    layer0_outputs(11002) <= not b;
    layer0_outputs(11003) <= not a;
    layer0_outputs(11004) <= not b or a;
    layer0_outputs(11005) <= a and b;
    layer0_outputs(11006) <= not a;
    layer0_outputs(11007) <= a and not b;
    layer0_outputs(11008) <= not b;
    layer0_outputs(11009) <= a;
    layer0_outputs(11010) <= a or b;
    layer0_outputs(11011) <= not a;
    layer0_outputs(11012) <= not (a xor b);
    layer0_outputs(11013) <= a and b;
    layer0_outputs(11014) <= not (a xor b);
    layer0_outputs(11015) <= a xor b;
    layer0_outputs(11016) <= not (a xor b);
    layer0_outputs(11017) <= a or b;
    layer0_outputs(11018) <= not (a xor b);
    layer0_outputs(11019) <= a or b;
    layer0_outputs(11020) <= not a or b;
    layer0_outputs(11021) <= not (a or b);
    layer0_outputs(11022) <= 1'b0;
    layer0_outputs(11023) <= a and not b;
    layer0_outputs(11024) <= not (a or b);
    layer0_outputs(11025) <= not (a xor b);
    layer0_outputs(11026) <= b and not a;
    layer0_outputs(11027) <= not b or a;
    layer0_outputs(11028) <= not a;
    layer0_outputs(11029) <= not (a or b);
    layer0_outputs(11030) <= b;
    layer0_outputs(11031) <= b;
    layer0_outputs(11032) <= b;
    layer0_outputs(11033) <= not (a xor b);
    layer0_outputs(11034) <= a;
    layer0_outputs(11035) <= not b or a;
    layer0_outputs(11036) <= b;
    layer0_outputs(11037) <= 1'b0;
    layer0_outputs(11038) <= a or b;
    layer0_outputs(11039) <= not (a xor b);
    layer0_outputs(11040) <= not a;
    layer0_outputs(11041) <= a xor b;
    layer0_outputs(11042) <= not b;
    layer0_outputs(11043) <= not (a xor b);
    layer0_outputs(11044) <= not a or b;
    layer0_outputs(11045) <= a and not b;
    layer0_outputs(11046) <= a or b;
    layer0_outputs(11047) <= a xor b;
    layer0_outputs(11048) <= not b;
    layer0_outputs(11049) <= a and b;
    layer0_outputs(11050) <= b and not a;
    layer0_outputs(11051) <= a and not b;
    layer0_outputs(11052) <= not b;
    layer0_outputs(11053) <= not b or a;
    layer0_outputs(11054) <= not a or b;
    layer0_outputs(11055) <= not (a xor b);
    layer0_outputs(11056) <= not b or a;
    layer0_outputs(11057) <= b and not a;
    layer0_outputs(11058) <= not a;
    layer0_outputs(11059) <= a and not b;
    layer0_outputs(11060) <= a or b;
    layer0_outputs(11061) <= not (a and b);
    layer0_outputs(11062) <= a xor b;
    layer0_outputs(11063) <= a;
    layer0_outputs(11064) <= a xor b;
    layer0_outputs(11065) <= not (a and b);
    layer0_outputs(11066) <= b and not a;
    layer0_outputs(11067) <= a or b;
    layer0_outputs(11068) <= not (a or b);
    layer0_outputs(11069) <= not a or b;
    layer0_outputs(11070) <= not b;
    layer0_outputs(11071) <= a and b;
    layer0_outputs(11072) <= not (a xor b);
    layer0_outputs(11073) <= a;
    layer0_outputs(11074) <= b and not a;
    layer0_outputs(11075) <= not (a and b);
    layer0_outputs(11076) <= not (a and b);
    layer0_outputs(11077) <= not (a xor b);
    layer0_outputs(11078) <= not (a or b);
    layer0_outputs(11079) <= b and not a;
    layer0_outputs(11080) <= not a;
    layer0_outputs(11081) <= not (a and b);
    layer0_outputs(11082) <= a xor b;
    layer0_outputs(11083) <= 1'b1;
    layer0_outputs(11084) <= not (a xor b);
    layer0_outputs(11085) <= not (a or b);
    layer0_outputs(11086) <= a xor b;
    layer0_outputs(11087) <= 1'b1;
    layer0_outputs(11088) <= not b or a;
    layer0_outputs(11089) <= a and not b;
    layer0_outputs(11090) <= not (a xor b);
    layer0_outputs(11091) <= a or b;
    layer0_outputs(11092) <= a or b;
    layer0_outputs(11093) <= a or b;
    layer0_outputs(11094) <= not b or a;
    layer0_outputs(11095) <= a;
    layer0_outputs(11096) <= a xor b;
    layer0_outputs(11097) <= not (a or b);
    layer0_outputs(11098) <= a;
    layer0_outputs(11099) <= not (a or b);
    layer0_outputs(11100) <= 1'b1;
    layer0_outputs(11101) <= not (a or b);
    layer0_outputs(11102) <= b;
    layer0_outputs(11103) <= not a or b;
    layer0_outputs(11104) <= not b;
    layer0_outputs(11105) <= not a or b;
    layer0_outputs(11106) <= not (a xor b);
    layer0_outputs(11107) <= not (a and b);
    layer0_outputs(11108) <= b;
    layer0_outputs(11109) <= not b;
    layer0_outputs(11110) <= 1'b0;
    layer0_outputs(11111) <= a or b;
    layer0_outputs(11112) <= not (a or b);
    layer0_outputs(11113) <= a and not b;
    layer0_outputs(11114) <= a and b;
    layer0_outputs(11115) <= not a;
    layer0_outputs(11116) <= not b or a;
    layer0_outputs(11117) <= a and b;
    layer0_outputs(11118) <= not a;
    layer0_outputs(11119) <= a;
    layer0_outputs(11120) <= not (a xor b);
    layer0_outputs(11121) <= a;
    layer0_outputs(11122) <= not b or a;
    layer0_outputs(11123) <= not (a and b);
    layer0_outputs(11124) <= a or b;
    layer0_outputs(11125) <= a or b;
    layer0_outputs(11126) <= not a or b;
    layer0_outputs(11127) <= not (a xor b);
    layer0_outputs(11128) <= a xor b;
    layer0_outputs(11129) <= not a or b;
    layer0_outputs(11130) <= a or b;
    layer0_outputs(11131) <= not b or a;
    layer0_outputs(11132) <= not (a or b);
    layer0_outputs(11133) <= not (a or b);
    layer0_outputs(11134) <= not (a or b);
    layer0_outputs(11135) <= a or b;
    layer0_outputs(11136) <= b;
    layer0_outputs(11137) <= a xor b;
    layer0_outputs(11138) <= not b or a;
    layer0_outputs(11139) <= a and b;
    layer0_outputs(11140) <= not a;
    layer0_outputs(11141) <= a and b;
    layer0_outputs(11142) <= a or b;
    layer0_outputs(11143) <= a and not b;
    layer0_outputs(11144) <= not (a or b);
    layer0_outputs(11145) <= not (a and b);
    layer0_outputs(11146) <= b and not a;
    layer0_outputs(11147) <= a xor b;
    layer0_outputs(11148) <= a xor b;
    layer0_outputs(11149) <= not b;
    layer0_outputs(11150) <= not (a xor b);
    layer0_outputs(11151) <= b and not a;
    layer0_outputs(11152) <= not (a xor b);
    layer0_outputs(11153) <= a;
    layer0_outputs(11154) <= not a or b;
    layer0_outputs(11155) <= not (a xor b);
    layer0_outputs(11156) <= not (a or b);
    layer0_outputs(11157) <= not (a or b);
    layer0_outputs(11158) <= b;
    layer0_outputs(11159) <= not (a xor b);
    layer0_outputs(11160) <= not a or b;
    layer0_outputs(11161) <= not b or a;
    layer0_outputs(11162) <= not a;
    layer0_outputs(11163) <= b;
    layer0_outputs(11164) <= a;
    layer0_outputs(11165) <= not a or b;
    layer0_outputs(11166) <= not b or a;
    layer0_outputs(11167) <= not b;
    layer0_outputs(11168) <= not (a or b);
    layer0_outputs(11169) <= not (a and b);
    layer0_outputs(11170) <= a or b;
    layer0_outputs(11171) <= a or b;
    layer0_outputs(11172) <= a and not b;
    layer0_outputs(11173) <= a;
    layer0_outputs(11174) <= a or b;
    layer0_outputs(11175) <= not (a or b);
    layer0_outputs(11176) <= not (a or b);
    layer0_outputs(11177) <= not (a or b);
    layer0_outputs(11178) <= a;
    layer0_outputs(11179) <= a;
    layer0_outputs(11180) <= not (a or b);
    layer0_outputs(11181) <= a;
    layer0_outputs(11182) <= a;
    layer0_outputs(11183) <= a xor b;
    layer0_outputs(11184) <= a xor b;
    layer0_outputs(11185) <= not b or a;
    layer0_outputs(11186) <= a;
    layer0_outputs(11187) <= not (a xor b);
    layer0_outputs(11188) <= a and b;
    layer0_outputs(11189) <= not (a or b);
    layer0_outputs(11190) <= not (a or b);
    layer0_outputs(11191) <= not b;
    layer0_outputs(11192) <= not (a or b);
    layer0_outputs(11193) <= not a;
    layer0_outputs(11194) <= b;
    layer0_outputs(11195) <= not b;
    layer0_outputs(11196) <= not (a or b);
    layer0_outputs(11197) <= not a or b;
    layer0_outputs(11198) <= not (a xor b);
    layer0_outputs(11199) <= a and not b;
    layer0_outputs(11200) <= b;
    layer0_outputs(11201) <= a or b;
    layer0_outputs(11202) <= a;
    layer0_outputs(11203) <= a or b;
    layer0_outputs(11204) <= not a;
    layer0_outputs(11205) <= not (a xor b);
    layer0_outputs(11206) <= a;
    layer0_outputs(11207) <= a or b;
    layer0_outputs(11208) <= not b or a;
    layer0_outputs(11209) <= not (a xor b);
    layer0_outputs(11210) <= a or b;
    layer0_outputs(11211) <= a and not b;
    layer0_outputs(11212) <= not (a or b);
    layer0_outputs(11213) <= a or b;
    layer0_outputs(11214) <= not (a xor b);
    layer0_outputs(11215) <= not b or a;
    layer0_outputs(11216) <= a or b;
    layer0_outputs(11217) <= not (a and b);
    layer0_outputs(11218) <= b and not a;
    layer0_outputs(11219) <= not (a xor b);
    layer0_outputs(11220) <= a xor b;
    layer0_outputs(11221) <= not a or b;
    layer0_outputs(11222) <= not a or b;
    layer0_outputs(11223) <= b;
    layer0_outputs(11224) <= not a;
    layer0_outputs(11225) <= a and not b;
    layer0_outputs(11226) <= b and not a;
    layer0_outputs(11227) <= a;
    layer0_outputs(11228) <= b;
    layer0_outputs(11229) <= not b or a;
    layer0_outputs(11230) <= not a or b;
    layer0_outputs(11231) <= 1'b0;
    layer0_outputs(11232) <= not b or a;
    layer0_outputs(11233) <= a or b;
    layer0_outputs(11234) <= not a or b;
    layer0_outputs(11235) <= b;
    layer0_outputs(11236) <= a and not b;
    layer0_outputs(11237) <= not (a or b);
    layer0_outputs(11238) <= not a;
    layer0_outputs(11239) <= a and b;
    layer0_outputs(11240) <= not b or a;
    layer0_outputs(11241) <= b;
    layer0_outputs(11242) <= 1'b0;
    layer0_outputs(11243) <= not (a xor b);
    layer0_outputs(11244) <= a and not b;
    layer0_outputs(11245) <= a xor b;
    layer0_outputs(11246) <= b;
    layer0_outputs(11247) <= not (a xor b);
    layer0_outputs(11248) <= b;
    layer0_outputs(11249) <= a or b;
    layer0_outputs(11250) <= a or b;
    layer0_outputs(11251) <= not (a or b);
    layer0_outputs(11252) <= b and not a;
    layer0_outputs(11253) <= not a;
    layer0_outputs(11254) <= b and not a;
    layer0_outputs(11255) <= a xor b;
    layer0_outputs(11256) <= 1'b1;
    layer0_outputs(11257) <= a xor b;
    layer0_outputs(11258) <= not b or a;
    layer0_outputs(11259) <= b;
    layer0_outputs(11260) <= a or b;
    layer0_outputs(11261) <= not (a xor b);
    layer0_outputs(11262) <= not a;
    layer0_outputs(11263) <= not b;
    layer0_outputs(11264) <= not (a xor b);
    layer0_outputs(11265) <= a and not b;
    layer0_outputs(11266) <= not b or a;
    layer0_outputs(11267) <= a xor b;
    layer0_outputs(11268) <= a;
    layer0_outputs(11269) <= a or b;
    layer0_outputs(11270) <= not b;
    layer0_outputs(11271) <= b and not a;
    layer0_outputs(11272) <= a xor b;
    layer0_outputs(11273) <= a and b;
    layer0_outputs(11274) <= not (a or b);
    layer0_outputs(11275) <= not (a or b);
    layer0_outputs(11276) <= not b;
    layer0_outputs(11277) <= not (a xor b);
    layer0_outputs(11278) <= 1'b1;
    layer0_outputs(11279) <= a;
    layer0_outputs(11280) <= a or b;
    layer0_outputs(11281) <= not a or b;
    layer0_outputs(11282) <= not (a or b);
    layer0_outputs(11283) <= not a or b;
    layer0_outputs(11284) <= not a;
    layer0_outputs(11285) <= 1'b1;
    layer0_outputs(11286) <= not a;
    layer0_outputs(11287) <= not b or a;
    layer0_outputs(11288) <= not (a xor b);
    layer0_outputs(11289) <= not a;
    layer0_outputs(11290) <= not (a or b);
    layer0_outputs(11291) <= a or b;
    layer0_outputs(11292) <= a or b;
    layer0_outputs(11293) <= a and not b;
    layer0_outputs(11294) <= not b or a;
    layer0_outputs(11295) <= a and not b;
    layer0_outputs(11296) <= a and not b;
    layer0_outputs(11297) <= a or b;
    layer0_outputs(11298) <= not (a and b);
    layer0_outputs(11299) <= not a or b;
    layer0_outputs(11300) <= a;
    layer0_outputs(11301) <= b and not a;
    layer0_outputs(11302) <= a or b;
    layer0_outputs(11303) <= not a or b;
    layer0_outputs(11304) <= a or b;
    layer0_outputs(11305) <= a and not b;
    layer0_outputs(11306) <= 1'b1;
    layer0_outputs(11307) <= a;
    layer0_outputs(11308) <= a xor b;
    layer0_outputs(11309) <= not a or b;
    layer0_outputs(11310) <= not b;
    layer0_outputs(11311) <= a or b;
    layer0_outputs(11312) <= not a or b;
    layer0_outputs(11313) <= b;
    layer0_outputs(11314) <= a and not b;
    layer0_outputs(11315) <= a and not b;
    layer0_outputs(11316) <= a xor b;
    layer0_outputs(11317) <= not a or b;
    layer0_outputs(11318) <= a or b;
    layer0_outputs(11319) <= not b or a;
    layer0_outputs(11320) <= not (a xor b);
    layer0_outputs(11321) <= a or b;
    layer0_outputs(11322) <= a or b;
    layer0_outputs(11323) <= not (a xor b);
    layer0_outputs(11324) <= not b;
    layer0_outputs(11325) <= not (a or b);
    layer0_outputs(11326) <= not b;
    layer0_outputs(11327) <= not a;
    layer0_outputs(11328) <= a;
    layer0_outputs(11329) <= not (a xor b);
    layer0_outputs(11330) <= not (a and b);
    layer0_outputs(11331) <= not a;
    layer0_outputs(11332) <= not b;
    layer0_outputs(11333) <= not b;
    layer0_outputs(11334) <= a xor b;
    layer0_outputs(11335) <= a xor b;
    layer0_outputs(11336) <= a xor b;
    layer0_outputs(11337) <= not a or b;
    layer0_outputs(11338) <= not b or a;
    layer0_outputs(11339) <= a or b;
    layer0_outputs(11340) <= a xor b;
    layer0_outputs(11341) <= a and not b;
    layer0_outputs(11342) <= a or b;
    layer0_outputs(11343) <= 1'b0;
    layer0_outputs(11344) <= b and not a;
    layer0_outputs(11345) <= not b;
    layer0_outputs(11346) <= b and not a;
    layer0_outputs(11347) <= not b;
    layer0_outputs(11348) <= a and not b;
    layer0_outputs(11349) <= a xor b;
    layer0_outputs(11350) <= not b;
    layer0_outputs(11351) <= not (a or b);
    layer0_outputs(11352) <= not (a or b);
    layer0_outputs(11353) <= a or b;
    layer0_outputs(11354) <= not b or a;
    layer0_outputs(11355) <= a xor b;
    layer0_outputs(11356) <= a;
    layer0_outputs(11357) <= 1'b1;
    layer0_outputs(11358) <= a xor b;
    layer0_outputs(11359) <= not b or a;
    layer0_outputs(11360) <= not (a or b);
    layer0_outputs(11361) <= not (a xor b);
    layer0_outputs(11362) <= a and not b;
    layer0_outputs(11363) <= not (a or b);
    layer0_outputs(11364) <= not a or b;
    layer0_outputs(11365) <= not (a and b);
    layer0_outputs(11366) <= not b;
    layer0_outputs(11367) <= a or b;
    layer0_outputs(11368) <= not a;
    layer0_outputs(11369) <= a xor b;
    layer0_outputs(11370) <= not (a or b);
    layer0_outputs(11371) <= not (a or b);
    layer0_outputs(11372) <= not (a xor b);
    layer0_outputs(11373) <= not (a and b);
    layer0_outputs(11374) <= a or b;
    layer0_outputs(11375) <= a;
    layer0_outputs(11376) <= not (a or b);
    layer0_outputs(11377) <= not b or a;
    layer0_outputs(11378) <= a and not b;
    layer0_outputs(11379) <= not (a and b);
    layer0_outputs(11380) <= a xor b;
    layer0_outputs(11381) <= a and b;
    layer0_outputs(11382) <= b;
    layer0_outputs(11383) <= not (a or b);
    layer0_outputs(11384) <= not b;
    layer0_outputs(11385) <= not a or b;
    layer0_outputs(11386) <= not a;
    layer0_outputs(11387) <= b;
    layer0_outputs(11388) <= a;
    layer0_outputs(11389) <= a;
    layer0_outputs(11390) <= not b or a;
    layer0_outputs(11391) <= a and b;
    layer0_outputs(11392) <= not (a or b);
    layer0_outputs(11393) <= not (a or b);
    layer0_outputs(11394) <= not (a or b);
    layer0_outputs(11395) <= b;
    layer0_outputs(11396) <= a or b;
    layer0_outputs(11397) <= a or b;
    layer0_outputs(11398) <= a xor b;
    layer0_outputs(11399) <= not b;
    layer0_outputs(11400) <= not a;
    layer0_outputs(11401) <= not a;
    layer0_outputs(11402) <= not a;
    layer0_outputs(11403) <= not (a or b);
    layer0_outputs(11404) <= not (a and b);
    layer0_outputs(11405) <= b and not a;
    layer0_outputs(11406) <= a xor b;
    layer0_outputs(11407) <= 1'b1;
    layer0_outputs(11408) <= not (a xor b);
    layer0_outputs(11409) <= not a;
    layer0_outputs(11410) <= a and not b;
    layer0_outputs(11411) <= not (a and b);
    layer0_outputs(11412) <= b;
    layer0_outputs(11413) <= b and not a;
    layer0_outputs(11414) <= a xor b;
    layer0_outputs(11415) <= not (a or b);
    layer0_outputs(11416) <= b and not a;
    layer0_outputs(11417) <= b;
    layer0_outputs(11418) <= not b;
    layer0_outputs(11419) <= not a;
    layer0_outputs(11420) <= a xor b;
    layer0_outputs(11421) <= not a;
    layer0_outputs(11422) <= not (a or b);
    layer0_outputs(11423) <= a xor b;
    layer0_outputs(11424) <= a or b;
    layer0_outputs(11425) <= not b;
    layer0_outputs(11426) <= b;
    layer0_outputs(11427) <= a or b;
    layer0_outputs(11428) <= not a;
    layer0_outputs(11429) <= b;
    layer0_outputs(11430) <= not b;
    layer0_outputs(11431) <= not b;
    layer0_outputs(11432) <= a xor b;
    layer0_outputs(11433) <= a;
    layer0_outputs(11434) <= a and b;
    layer0_outputs(11435) <= a;
    layer0_outputs(11436) <= b and not a;
    layer0_outputs(11437) <= not b;
    layer0_outputs(11438) <= not b or a;
    layer0_outputs(11439) <= a xor b;
    layer0_outputs(11440) <= a or b;
    layer0_outputs(11441) <= a xor b;
    layer0_outputs(11442) <= not a or b;
    layer0_outputs(11443) <= b;
    layer0_outputs(11444) <= b and not a;
    layer0_outputs(11445) <= a or b;
    layer0_outputs(11446) <= not a;
    layer0_outputs(11447) <= a xor b;
    layer0_outputs(11448) <= a xor b;
    layer0_outputs(11449) <= not b;
    layer0_outputs(11450) <= b and not a;
    layer0_outputs(11451) <= a;
    layer0_outputs(11452) <= a xor b;
    layer0_outputs(11453) <= 1'b0;
    layer0_outputs(11454) <= b;
    layer0_outputs(11455) <= a or b;
    layer0_outputs(11456) <= not (a or b);
    layer0_outputs(11457) <= not a;
    layer0_outputs(11458) <= not a;
    layer0_outputs(11459) <= a xor b;
    layer0_outputs(11460) <= not (a or b);
    layer0_outputs(11461) <= a or b;
    layer0_outputs(11462) <= a or b;
    layer0_outputs(11463) <= a or b;
    layer0_outputs(11464) <= not (a xor b);
    layer0_outputs(11465) <= b;
    layer0_outputs(11466) <= not a;
    layer0_outputs(11467) <= a or b;
    layer0_outputs(11468) <= not (a or b);
    layer0_outputs(11469) <= not (a xor b);
    layer0_outputs(11470) <= not a or b;
    layer0_outputs(11471) <= not (a xor b);
    layer0_outputs(11472) <= 1'b1;
    layer0_outputs(11473) <= a xor b;
    layer0_outputs(11474) <= not (a xor b);
    layer0_outputs(11475) <= b;
    layer0_outputs(11476) <= a xor b;
    layer0_outputs(11477) <= not a;
    layer0_outputs(11478) <= not (a xor b);
    layer0_outputs(11479) <= not a or b;
    layer0_outputs(11480) <= a;
    layer0_outputs(11481) <= not (a or b);
    layer0_outputs(11482) <= b and not a;
    layer0_outputs(11483) <= a or b;
    layer0_outputs(11484) <= 1'b1;
    layer0_outputs(11485) <= a and b;
    layer0_outputs(11486) <= b and not a;
    layer0_outputs(11487) <= not b;
    layer0_outputs(11488) <= a;
    layer0_outputs(11489) <= a and b;
    layer0_outputs(11490) <= b;
    layer0_outputs(11491) <= a xor b;
    layer0_outputs(11492) <= a or b;
    layer0_outputs(11493) <= not b or a;
    layer0_outputs(11494) <= b and not a;
    layer0_outputs(11495) <= b and not a;
    layer0_outputs(11496) <= a or b;
    layer0_outputs(11497) <= not a or b;
    layer0_outputs(11498) <= b;
    layer0_outputs(11499) <= not (a xor b);
    layer0_outputs(11500) <= not (a xor b);
    layer0_outputs(11501) <= not b or a;
    layer0_outputs(11502) <= not (a or b);
    layer0_outputs(11503) <= not (a or b);
    layer0_outputs(11504) <= not b;
    layer0_outputs(11505) <= a xor b;
    layer0_outputs(11506) <= not a or b;
    layer0_outputs(11507) <= b and not a;
    layer0_outputs(11508) <= not b;
    layer0_outputs(11509) <= a or b;
    layer0_outputs(11510) <= b;
    layer0_outputs(11511) <= a;
    layer0_outputs(11512) <= b;
    layer0_outputs(11513) <= not a or b;
    layer0_outputs(11514) <= a xor b;
    layer0_outputs(11515) <= not (a or b);
    layer0_outputs(11516) <= a or b;
    layer0_outputs(11517) <= not (a xor b);
    layer0_outputs(11518) <= not a or b;
    layer0_outputs(11519) <= b;
    layer0_outputs(11520) <= b;
    layer0_outputs(11521) <= not (a or b);
    layer0_outputs(11522) <= not a;
    layer0_outputs(11523) <= not b or a;
    layer0_outputs(11524) <= not a;
    layer0_outputs(11525) <= not a or b;
    layer0_outputs(11526) <= a xor b;
    layer0_outputs(11527) <= not (a and b);
    layer0_outputs(11528) <= not (a or b);
    layer0_outputs(11529) <= a and b;
    layer0_outputs(11530) <= not (a or b);
    layer0_outputs(11531) <= a or b;
    layer0_outputs(11532) <= a and b;
    layer0_outputs(11533) <= not (a xor b);
    layer0_outputs(11534) <= not (a and b);
    layer0_outputs(11535) <= b;
    layer0_outputs(11536) <= a and not b;
    layer0_outputs(11537) <= not b;
    layer0_outputs(11538) <= a or b;
    layer0_outputs(11539) <= not (a or b);
    layer0_outputs(11540) <= a or b;
    layer0_outputs(11541) <= not b;
    layer0_outputs(11542) <= a xor b;
    layer0_outputs(11543) <= not (a xor b);
    layer0_outputs(11544) <= a and not b;
    layer0_outputs(11545) <= not (a or b);
    layer0_outputs(11546) <= a xor b;
    layer0_outputs(11547) <= not a;
    layer0_outputs(11548) <= not (a or b);
    layer0_outputs(11549) <= 1'b0;
    layer0_outputs(11550) <= b;
    layer0_outputs(11551) <= not (a or b);
    layer0_outputs(11552) <= not a or b;
    layer0_outputs(11553) <= not (a xor b);
    layer0_outputs(11554) <= not (a or b);
    layer0_outputs(11555) <= a xor b;
    layer0_outputs(11556) <= not a;
    layer0_outputs(11557) <= a xor b;
    layer0_outputs(11558) <= a;
    layer0_outputs(11559) <= 1'b0;
    layer0_outputs(11560) <= not (a or b);
    layer0_outputs(11561) <= not b;
    layer0_outputs(11562) <= b;
    layer0_outputs(11563) <= not (a or b);
    layer0_outputs(11564) <= a and not b;
    layer0_outputs(11565) <= not a or b;
    layer0_outputs(11566) <= not (a or b);
    layer0_outputs(11567) <= not b;
    layer0_outputs(11568) <= not (a or b);
    layer0_outputs(11569) <= a;
    layer0_outputs(11570) <= not (a xor b);
    layer0_outputs(11571) <= not (a or b);
    layer0_outputs(11572) <= a;
    layer0_outputs(11573) <= not (a or b);
    layer0_outputs(11574) <= not (a or b);
    layer0_outputs(11575) <= not b;
    layer0_outputs(11576) <= not a or b;
    layer0_outputs(11577) <= a and b;
    layer0_outputs(11578) <= a and b;
    layer0_outputs(11579) <= not (a or b);
    layer0_outputs(11580) <= a or b;
    layer0_outputs(11581) <= not a or b;
    layer0_outputs(11582) <= a xor b;
    layer0_outputs(11583) <= not (a or b);
    layer0_outputs(11584) <= b;
    layer0_outputs(11585) <= not b;
    layer0_outputs(11586) <= b;
    layer0_outputs(11587) <= a and not b;
    layer0_outputs(11588) <= not a;
    layer0_outputs(11589) <= not (a or b);
    layer0_outputs(11590) <= not a or b;
    layer0_outputs(11591) <= not (a and b);
    layer0_outputs(11592) <= a and not b;
    layer0_outputs(11593) <= a and b;
    layer0_outputs(11594) <= a or b;
    layer0_outputs(11595) <= not b;
    layer0_outputs(11596) <= a or b;
    layer0_outputs(11597) <= a and not b;
    layer0_outputs(11598) <= not (a xor b);
    layer0_outputs(11599) <= not (a or b);
    layer0_outputs(11600) <= a and not b;
    layer0_outputs(11601) <= a or b;
    layer0_outputs(11602) <= not (a and b);
    layer0_outputs(11603) <= not (a xor b);
    layer0_outputs(11604) <= a or b;
    layer0_outputs(11605) <= a or b;
    layer0_outputs(11606) <= a and not b;
    layer0_outputs(11607) <= a and not b;
    layer0_outputs(11608) <= 1'b0;
    layer0_outputs(11609) <= a or b;
    layer0_outputs(11610) <= a;
    layer0_outputs(11611) <= a or b;
    layer0_outputs(11612) <= a and not b;
    layer0_outputs(11613) <= not (a xor b);
    layer0_outputs(11614) <= not b;
    layer0_outputs(11615) <= not (a xor b);
    layer0_outputs(11616) <= not (a xor b);
    layer0_outputs(11617) <= not (a xor b);
    layer0_outputs(11618) <= a xor b;
    layer0_outputs(11619) <= not a or b;
    layer0_outputs(11620) <= a or b;
    layer0_outputs(11621) <= a and not b;
    layer0_outputs(11622) <= not (a xor b);
    layer0_outputs(11623) <= b and not a;
    layer0_outputs(11624) <= a xor b;
    layer0_outputs(11625) <= a;
    layer0_outputs(11626) <= a;
    layer0_outputs(11627) <= not a or b;
    layer0_outputs(11628) <= not b;
    layer0_outputs(11629) <= b and not a;
    layer0_outputs(11630) <= not (a or b);
    layer0_outputs(11631) <= a or b;
    layer0_outputs(11632) <= a and not b;
    layer0_outputs(11633) <= not a;
    layer0_outputs(11634) <= a xor b;
    layer0_outputs(11635) <= a or b;
    layer0_outputs(11636) <= not b;
    layer0_outputs(11637) <= a or b;
    layer0_outputs(11638) <= a or b;
    layer0_outputs(11639) <= not a;
    layer0_outputs(11640) <= b;
    layer0_outputs(11641) <= not b;
    layer0_outputs(11642) <= not b or a;
    layer0_outputs(11643) <= a;
    layer0_outputs(11644) <= not a or b;
    layer0_outputs(11645) <= not (a and b);
    layer0_outputs(11646) <= b and not a;
    layer0_outputs(11647) <= b and not a;
    layer0_outputs(11648) <= b and not a;
    layer0_outputs(11649) <= not (a xor b);
    layer0_outputs(11650) <= b and not a;
    layer0_outputs(11651) <= a or b;
    layer0_outputs(11652) <= a xor b;
    layer0_outputs(11653) <= not (a or b);
    layer0_outputs(11654) <= a or b;
    layer0_outputs(11655) <= a or b;
    layer0_outputs(11656) <= a or b;
    layer0_outputs(11657) <= not (a or b);
    layer0_outputs(11658) <= not (a or b);
    layer0_outputs(11659) <= a xor b;
    layer0_outputs(11660) <= b;
    layer0_outputs(11661) <= not a or b;
    layer0_outputs(11662) <= not (a xor b);
    layer0_outputs(11663) <= a and b;
    layer0_outputs(11664) <= not (a or b);
    layer0_outputs(11665) <= not (a and b);
    layer0_outputs(11666) <= not b;
    layer0_outputs(11667) <= not a or b;
    layer0_outputs(11668) <= a or b;
    layer0_outputs(11669) <= not b or a;
    layer0_outputs(11670) <= not b;
    layer0_outputs(11671) <= a xor b;
    layer0_outputs(11672) <= not b or a;
    layer0_outputs(11673) <= not a;
    layer0_outputs(11674) <= a;
    layer0_outputs(11675) <= a or b;
    layer0_outputs(11676) <= a xor b;
    layer0_outputs(11677) <= 1'b0;
    layer0_outputs(11678) <= not (a and b);
    layer0_outputs(11679) <= a xor b;
    layer0_outputs(11680) <= not (a and b);
    layer0_outputs(11681) <= not (a xor b);
    layer0_outputs(11682) <= not (a or b);
    layer0_outputs(11683) <= not (a and b);
    layer0_outputs(11684) <= 1'b0;
    layer0_outputs(11685) <= a;
    layer0_outputs(11686) <= not (a and b);
    layer0_outputs(11687) <= not (a or b);
    layer0_outputs(11688) <= not b;
    layer0_outputs(11689) <= a xor b;
    layer0_outputs(11690) <= a or b;
    layer0_outputs(11691) <= a;
    layer0_outputs(11692) <= b and not a;
    layer0_outputs(11693) <= b;
    layer0_outputs(11694) <= not (a and b);
    layer0_outputs(11695) <= b;
    layer0_outputs(11696) <= a xor b;
    layer0_outputs(11697) <= a or b;
    layer0_outputs(11698) <= not b;
    layer0_outputs(11699) <= not (a xor b);
    layer0_outputs(11700) <= not a;
    layer0_outputs(11701) <= a and b;
    layer0_outputs(11702) <= b;
    layer0_outputs(11703) <= a;
    layer0_outputs(11704) <= b;
    layer0_outputs(11705) <= b and not a;
    layer0_outputs(11706) <= not (a and b);
    layer0_outputs(11707) <= a xor b;
    layer0_outputs(11708) <= a or b;
    layer0_outputs(11709) <= b;
    layer0_outputs(11710) <= a or b;
    layer0_outputs(11711) <= a or b;
    layer0_outputs(11712) <= not (a xor b);
    layer0_outputs(11713) <= not (a and b);
    layer0_outputs(11714) <= not (a or b);
    layer0_outputs(11715) <= not (a xor b);
    layer0_outputs(11716) <= not (a xor b);
    layer0_outputs(11717) <= not a or b;
    layer0_outputs(11718) <= not (a and b);
    layer0_outputs(11719) <= a or b;
    layer0_outputs(11720) <= not (a or b);
    layer0_outputs(11721) <= a xor b;
    layer0_outputs(11722) <= not (a or b);
    layer0_outputs(11723) <= a xor b;
    layer0_outputs(11724) <= a xor b;
    layer0_outputs(11725) <= a and not b;
    layer0_outputs(11726) <= a xor b;
    layer0_outputs(11727) <= not b;
    layer0_outputs(11728) <= a or b;
    layer0_outputs(11729) <= a xor b;
    layer0_outputs(11730) <= not b;
    layer0_outputs(11731) <= 1'b1;
    layer0_outputs(11732) <= b;
    layer0_outputs(11733) <= b;
    layer0_outputs(11734) <= a xor b;
    layer0_outputs(11735) <= not b or a;
    layer0_outputs(11736) <= b and not a;
    layer0_outputs(11737) <= a and not b;
    layer0_outputs(11738) <= not b or a;
    layer0_outputs(11739) <= not (a xor b);
    layer0_outputs(11740) <= not (a or b);
    layer0_outputs(11741) <= a xor b;
    layer0_outputs(11742) <= a or b;
    layer0_outputs(11743) <= not b;
    layer0_outputs(11744) <= a and not b;
    layer0_outputs(11745) <= a xor b;
    layer0_outputs(11746) <= a or b;
    layer0_outputs(11747) <= not (a xor b);
    layer0_outputs(11748) <= not b;
    layer0_outputs(11749) <= not (a xor b);
    layer0_outputs(11750) <= not a or b;
    layer0_outputs(11751) <= a and b;
    layer0_outputs(11752) <= not (a and b);
    layer0_outputs(11753) <= a or b;
    layer0_outputs(11754) <= not (a or b);
    layer0_outputs(11755) <= a or b;
    layer0_outputs(11756) <= a and b;
    layer0_outputs(11757) <= not (a or b);
    layer0_outputs(11758) <= 1'b1;
    layer0_outputs(11759) <= not b or a;
    layer0_outputs(11760) <= b and not a;
    layer0_outputs(11761) <= a;
    layer0_outputs(11762) <= a;
    layer0_outputs(11763) <= b and not a;
    layer0_outputs(11764) <= a and b;
    layer0_outputs(11765) <= not a or b;
    layer0_outputs(11766) <= a xor b;
    layer0_outputs(11767) <= a xor b;
    layer0_outputs(11768) <= b and not a;
    layer0_outputs(11769) <= not (a xor b);
    layer0_outputs(11770) <= not (a xor b);
    layer0_outputs(11771) <= not a or b;
    layer0_outputs(11772) <= not (a or b);
    layer0_outputs(11773) <= 1'b1;
    layer0_outputs(11774) <= a xor b;
    layer0_outputs(11775) <= b;
    layer0_outputs(11776) <= not (a or b);
    layer0_outputs(11777) <= 1'b1;
    layer0_outputs(11778) <= b;
    layer0_outputs(11779) <= not (a xor b);
    layer0_outputs(11780) <= not (a or b);
    layer0_outputs(11781) <= not b;
    layer0_outputs(11782) <= b;
    layer0_outputs(11783) <= b;
    layer0_outputs(11784) <= a xor b;
    layer0_outputs(11785) <= not a or b;
    layer0_outputs(11786) <= not a or b;
    layer0_outputs(11787) <= b and not a;
    layer0_outputs(11788) <= not a;
    layer0_outputs(11789) <= a xor b;
    layer0_outputs(11790) <= not a;
    layer0_outputs(11791) <= not a or b;
    layer0_outputs(11792) <= not a or b;
    layer0_outputs(11793) <= a and not b;
    layer0_outputs(11794) <= not (a xor b);
    layer0_outputs(11795) <= not a;
    layer0_outputs(11796) <= b and not a;
    layer0_outputs(11797) <= a;
    layer0_outputs(11798) <= b;
    layer0_outputs(11799) <= not a;
    layer0_outputs(11800) <= a or b;
    layer0_outputs(11801) <= not a or b;
    layer0_outputs(11802) <= a and not b;
    layer0_outputs(11803) <= a or b;
    layer0_outputs(11804) <= 1'b0;
    layer0_outputs(11805) <= a;
    layer0_outputs(11806) <= not (a xor b);
    layer0_outputs(11807) <= a;
    layer0_outputs(11808) <= a or b;
    layer0_outputs(11809) <= a or b;
    layer0_outputs(11810) <= a or b;
    layer0_outputs(11811) <= a or b;
    layer0_outputs(11812) <= not b;
    layer0_outputs(11813) <= b;
    layer0_outputs(11814) <= not (a and b);
    layer0_outputs(11815) <= a xor b;
    layer0_outputs(11816) <= a or b;
    layer0_outputs(11817) <= not a;
    layer0_outputs(11818) <= not (a or b);
    layer0_outputs(11819) <= not (a xor b);
    layer0_outputs(11820) <= b and not a;
    layer0_outputs(11821) <= a;
    layer0_outputs(11822) <= b;
    layer0_outputs(11823) <= not a;
    layer0_outputs(11824) <= b;
    layer0_outputs(11825) <= a or b;
    layer0_outputs(11826) <= not b or a;
    layer0_outputs(11827) <= b;
    layer0_outputs(11828) <= a and b;
    layer0_outputs(11829) <= not (a or b);
    layer0_outputs(11830) <= b and not a;
    layer0_outputs(11831) <= a or b;
    layer0_outputs(11832) <= not b or a;
    layer0_outputs(11833) <= a and b;
    layer0_outputs(11834) <= not (a xor b);
    layer0_outputs(11835) <= a or b;
    layer0_outputs(11836) <= not (a or b);
    layer0_outputs(11837) <= not (a or b);
    layer0_outputs(11838) <= a and not b;
    layer0_outputs(11839) <= b;
    layer0_outputs(11840) <= a xor b;
    layer0_outputs(11841) <= a;
    layer0_outputs(11842) <= a xor b;
    layer0_outputs(11843) <= not a;
    layer0_outputs(11844) <= a xor b;
    layer0_outputs(11845) <= a and not b;
    layer0_outputs(11846) <= not a or b;
    layer0_outputs(11847) <= a xor b;
    layer0_outputs(11848) <= a;
    layer0_outputs(11849) <= not a or b;
    layer0_outputs(11850) <= not (a or b);
    layer0_outputs(11851) <= not a;
    layer0_outputs(11852) <= not (a or b);
    layer0_outputs(11853) <= a or b;
    layer0_outputs(11854) <= not (a xor b);
    layer0_outputs(11855) <= a and not b;
    layer0_outputs(11856) <= not (a and b);
    layer0_outputs(11857) <= not b;
    layer0_outputs(11858) <= b;
    layer0_outputs(11859) <= b and not a;
    layer0_outputs(11860) <= a and not b;
    layer0_outputs(11861) <= not a or b;
    layer0_outputs(11862) <= not (a xor b);
    layer0_outputs(11863) <= not (a or b);
    layer0_outputs(11864) <= not (a and b);
    layer0_outputs(11865) <= 1'b0;
    layer0_outputs(11866) <= not a;
    layer0_outputs(11867) <= 1'b0;
    layer0_outputs(11868) <= not b or a;
    layer0_outputs(11869) <= a and not b;
    layer0_outputs(11870) <= a xor b;
    layer0_outputs(11871) <= 1'b1;
    layer0_outputs(11872) <= a;
    layer0_outputs(11873) <= a or b;
    layer0_outputs(11874) <= not a;
    layer0_outputs(11875) <= not b;
    layer0_outputs(11876) <= a or b;
    layer0_outputs(11877) <= 1'b0;
    layer0_outputs(11878) <= not a or b;
    layer0_outputs(11879) <= not b or a;
    layer0_outputs(11880) <= not b;
    layer0_outputs(11881) <= b and not a;
    layer0_outputs(11882) <= a or b;
    layer0_outputs(11883) <= not b;
    layer0_outputs(11884) <= a;
    layer0_outputs(11885) <= b and not a;
    layer0_outputs(11886) <= b and not a;
    layer0_outputs(11887) <= b;
    layer0_outputs(11888) <= not (a xor b);
    layer0_outputs(11889) <= a or b;
    layer0_outputs(11890) <= 1'b1;
    layer0_outputs(11891) <= 1'b1;
    layer0_outputs(11892) <= not b or a;
    layer0_outputs(11893) <= a or b;
    layer0_outputs(11894) <= not (a and b);
    layer0_outputs(11895) <= not (a or b);
    layer0_outputs(11896) <= a and b;
    layer0_outputs(11897) <= a xor b;
    layer0_outputs(11898) <= a;
    layer0_outputs(11899) <= b and not a;
    layer0_outputs(11900) <= not (a or b);
    layer0_outputs(11901) <= not b;
    layer0_outputs(11902) <= not b;
    layer0_outputs(11903) <= not b;
    layer0_outputs(11904) <= 1'b1;
    layer0_outputs(11905) <= a xor b;
    layer0_outputs(11906) <= a and not b;
    layer0_outputs(11907) <= not (a and b);
    layer0_outputs(11908) <= a and not b;
    layer0_outputs(11909) <= a or b;
    layer0_outputs(11910) <= a xor b;
    layer0_outputs(11911) <= a or b;
    layer0_outputs(11912) <= a xor b;
    layer0_outputs(11913) <= not (a and b);
    layer0_outputs(11914) <= a or b;
    layer0_outputs(11915) <= a and b;
    layer0_outputs(11916) <= a xor b;
    layer0_outputs(11917) <= not b;
    layer0_outputs(11918) <= not b or a;
    layer0_outputs(11919) <= not (a and b);
    layer0_outputs(11920) <= a or b;
    layer0_outputs(11921) <= a;
    layer0_outputs(11922) <= 1'b1;
    layer0_outputs(11923) <= a and not b;
    layer0_outputs(11924) <= a or b;
    layer0_outputs(11925) <= not (a or b);
    layer0_outputs(11926) <= not (a xor b);
    layer0_outputs(11927) <= b;
    layer0_outputs(11928) <= not (a xor b);
    layer0_outputs(11929) <= a or b;
    layer0_outputs(11930) <= not a or b;
    layer0_outputs(11931) <= a;
    layer0_outputs(11932) <= a xor b;
    layer0_outputs(11933) <= not (a or b);
    layer0_outputs(11934) <= a and not b;
    layer0_outputs(11935) <= 1'b1;
    layer0_outputs(11936) <= b;
    layer0_outputs(11937) <= not a;
    layer0_outputs(11938) <= not (a and b);
    layer0_outputs(11939) <= a and b;
    layer0_outputs(11940) <= not (a or b);
    layer0_outputs(11941) <= not (a or b);
    layer0_outputs(11942) <= a and not b;
    layer0_outputs(11943) <= a and not b;
    layer0_outputs(11944) <= a or b;
    layer0_outputs(11945) <= a xor b;
    layer0_outputs(11946) <= a xor b;
    layer0_outputs(11947) <= not b;
    layer0_outputs(11948) <= not b or a;
    layer0_outputs(11949) <= b;
    layer0_outputs(11950) <= not a;
    layer0_outputs(11951) <= not (a xor b);
    layer0_outputs(11952) <= a;
    layer0_outputs(11953) <= not (a or b);
    layer0_outputs(11954) <= a or b;
    layer0_outputs(11955) <= not a or b;
    layer0_outputs(11956) <= a and b;
    layer0_outputs(11957) <= a xor b;
    layer0_outputs(11958) <= a or b;
    layer0_outputs(11959) <= b;
    layer0_outputs(11960) <= a xor b;
    layer0_outputs(11961) <= not b or a;
    layer0_outputs(11962) <= not a;
    layer0_outputs(11963) <= b;
    layer0_outputs(11964) <= not a;
    layer0_outputs(11965) <= not (a xor b);
    layer0_outputs(11966) <= a and not b;
    layer0_outputs(11967) <= not (a xor b);
    layer0_outputs(11968) <= a;
    layer0_outputs(11969) <= b;
    layer0_outputs(11970) <= a xor b;
    layer0_outputs(11971) <= not a or b;
    layer0_outputs(11972) <= a xor b;
    layer0_outputs(11973) <= a or b;
    layer0_outputs(11974) <= not (a xor b);
    layer0_outputs(11975) <= not (a xor b);
    layer0_outputs(11976) <= a or b;
    layer0_outputs(11977) <= b;
    layer0_outputs(11978) <= a;
    layer0_outputs(11979) <= not a or b;
    layer0_outputs(11980) <= a or b;
    layer0_outputs(11981) <= b;
    layer0_outputs(11982) <= a xor b;
    layer0_outputs(11983) <= not b;
    layer0_outputs(11984) <= not (a xor b);
    layer0_outputs(11985) <= a and not b;
    layer0_outputs(11986) <= not (a xor b);
    layer0_outputs(11987) <= not (a or b);
    layer0_outputs(11988) <= b;
    layer0_outputs(11989) <= b;
    layer0_outputs(11990) <= a xor b;
    layer0_outputs(11991) <= a xor b;
    layer0_outputs(11992) <= a and not b;
    layer0_outputs(11993) <= a or b;
    layer0_outputs(11994) <= b;
    layer0_outputs(11995) <= not b or a;
    layer0_outputs(11996) <= a or b;
    layer0_outputs(11997) <= not a or b;
    layer0_outputs(11998) <= a xor b;
    layer0_outputs(11999) <= not (a xor b);
    layer0_outputs(12000) <= not a;
    layer0_outputs(12001) <= a and not b;
    layer0_outputs(12002) <= a and b;
    layer0_outputs(12003) <= not (a or b);
    layer0_outputs(12004) <= not b;
    layer0_outputs(12005) <= not a;
    layer0_outputs(12006) <= b and not a;
    layer0_outputs(12007) <= not b or a;
    layer0_outputs(12008) <= not b;
    layer0_outputs(12009) <= not a;
    layer0_outputs(12010) <= not b;
    layer0_outputs(12011) <= a;
    layer0_outputs(12012) <= not a or b;
    layer0_outputs(12013) <= a and not b;
    layer0_outputs(12014) <= not a;
    layer0_outputs(12015) <= a and not b;
    layer0_outputs(12016) <= a and not b;
    layer0_outputs(12017) <= not (a xor b);
    layer0_outputs(12018) <= not a or b;
    layer0_outputs(12019) <= not b;
    layer0_outputs(12020) <= b;
    layer0_outputs(12021) <= a or b;
    layer0_outputs(12022) <= not (a or b);
    layer0_outputs(12023) <= 1'b1;
    layer0_outputs(12024) <= b and not a;
    layer0_outputs(12025) <= not b or a;
    layer0_outputs(12026) <= a or b;
    layer0_outputs(12027) <= not a or b;
    layer0_outputs(12028) <= a or b;
    layer0_outputs(12029) <= not b or a;
    layer0_outputs(12030) <= b;
    layer0_outputs(12031) <= a xor b;
    layer0_outputs(12032) <= not b or a;
    layer0_outputs(12033) <= a;
    layer0_outputs(12034) <= not a or b;
    layer0_outputs(12035) <= not (a or b);
    layer0_outputs(12036) <= not (a xor b);
    layer0_outputs(12037) <= b;
    layer0_outputs(12038) <= 1'b1;
    layer0_outputs(12039) <= a;
    layer0_outputs(12040) <= b and not a;
    layer0_outputs(12041) <= a and b;
    layer0_outputs(12042) <= not (a xor b);
    layer0_outputs(12043) <= not (a or b);
    layer0_outputs(12044) <= a and not b;
    layer0_outputs(12045) <= not (a or b);
    layer0_outputs(12046) <= a and not b;
    layer0_outputs(12047) <= not b;
    layer0_outputs(12048) <= not (a or b);
    layer0_outputs(12049) <= a xor b;
    layer0_outputs(12050) <= not (a and b);
    layer0_outputs(12051) <= not (a or b);
    layer0_outputs(12052) <= b;
    layer0_outputs(12053) <= not b;
    layer0_outputs(12054) <= not b;
    layer0_outputs(12055) <= b;
    layer0_outputs(12056) <= a and not b;
    layer0_outputs(12057) <= not b;
    layer0_outputs(12058) <= a;
    layer0_outputs(12059) <= a and not b;
    layer0_outputs(12060) <= a xor b;
    layer0_outputs(12061) <= not (a or b);
    layer0_outputs(12062) <= b;
    layer0_outputs(12063) <= a xor b;
    layer0_outputs(12064) <= b;
    layer0_outputs(12065) <= a xor b;
    layer0_outputs(12066) <= b;
    layer0_outputs(12067) <= not (a xor b);
    layer0_outputs(12068) <= b;
    layer0_outputs(12069) <= 1'b0;
    layer0_outputs(12070) <= a;
    layer0_outputs(12071) <= a or b;
    layer0_outputs(12072) <= not (a or b);
    layer0_outputs(12073) <= not a;
    layer0_outputs(12074) <= not (a xor b);
    layer0_outputs(12075) <= not a or b;
    layer0_outputs(12076) <= not b or a;
    layer0_outputs(12077) <= not (a and b);
    layer0_outputs(12078) <= not (a or b);
    layer0_outputs(12079) <= a or b;
    layer0_outputs(12080) <= b;
    layer0_outputs(12081) <= b and not a;
    layer0_outputs(12082) <= not b;
    layer0_outputs(12083) <= a and not b;
    layer0_outputs(12084) <= not (a xor b);
    layer0_outputs(12085) <= not (a or b);
    layer0_outputs(12086) <= b and not a;
    layer0_outputs(12087) <= 1'b1;
    layer0_outputs(12088) <= 1'b0;
    layer0_outputs(12089) <= a xor b;
    layer0_outputs(12090) <= a xor b;
    layer0_outputs(12091) <= b and not a;
    layer0_outputs(12092) <= a xor b;
    layer0_outputs(12093) <= b and not a;
    layer0_outputs(12094) <= a and b;
    layer0_outputs(12095) <= not a or b;
    layer0_outputs(12096) <= a or b;
    layer0_outputs(12097) <= a;
    layer0_outputs(12098) <= b and not a;
    layer0_outputs(12099) <= not b;
    layer0_outputs(12100) <= 1'b0;
    layer0_outputs(12101) <= not b;
    layer0_outputs(12102) <= not a;
    layer0_outputs(12103) <= b and not a;
    layer0_outputs(12104) <= b and not a;
    layer0_outputs(12105) <= not a;
    layer0_outputs(12106) <= not a;
    layer0_outputs(12107) <= not (a xor b);
    layer0_outputs(12108) <= not a;
    layer0_outputs(12109) <= not (a and b);
    layer0_outputs(12110) <= not b;
    layer0_outputs(12111) <= not a;
    layer0_outputs(12112) <= not (a or b);
    layer0_outputs(12113) <= not b or a;
    layer0_outputs(12114) <= 1'b0;
    layer0_outputs(12115) <= not b;
    layer0_outputs(12116) <= 1'b1;
    layer0_outputs(12117) <= 1'b0;
    layer0_outputs(12118) <= not b or a;
    layer0_outputs(12119) <= a or b;
    layer0_outputs(12120) <= not (a xor b);
    layer0_outputs(12121) <= not b;
    layer0_outputs(12122) <= a or b;
    layer0_outputs(12123) <= b and not a;
    layer0_outputs(12124) <= not b;
    layer0_outputs(12125) <= a;
    layer0_outputs(12126) <= not (a xor b);
    layer0_outputs(12127) <= not (a xor b);
    layer0_outputs(12128) <= b and not a;
    layer0_outputs(12129) <= not a;
    layer0_outputs(12130) <= not b or a;
    layer0_outputs(12131) <= b;
    layer0_outputs(12132) <= not (a and b);
    layer0_outputs(12133) <= not (a or b);
    layer0_outputs(12134) <= 1'b0;
    layer0_outputs(12135) <= a xor b;
    layer0_outputs(12136) <= b;
    layer0_outputs(12137) <= a or b;
    layer0_outputs(12138) <= not a;
    layer0_outputs(12139) <= b and not a;
    layer0_outputs(12140) <= a;
    layer0_outputs(12141) <= not (a or b);
    layer0_outputs(12142) <= a xor b;
    layer0_outputs(12143) <= not a;
    layer0_outputs(12144) <= a or b;
    layer0_outputs(12145) <= not a or b;
    layer0_outputs(12146) <= not b or a;
    layer0_outputs(12147) <= not b;
    layer0_outputs(12148) <= a and not b;
    layer0_outputs(12149) <= a or b;
    layer0_outputs(12150) <= b and not a;
    layer0_outputs(12151) <= not (a xor b);
    layer0_outputs(12152) <= not a or b;
    layer0_outputs(12153) <= not b or a;
    layer0_outputs(12154) <= not b or a;
    layer0_outputs(12155) <= not (a or b);
    layer0_outputs(12156) <= not b;
    layer0_outputs(12157) <= not a or b;
    layer0_outputs(12158) <= not b or a;
    layer0_outputs(12159) <= not a or b;
    layer0_outputs(12160) <= not (a or b);
    layer0_outputs(12161) <= a or b;
    layer0_outputs(12162) <= 1'b1;
    layer0_outputs(12163) <= a or b;
    layer0_outputs(12164) <= b and not a;
    layer0_outputs(12165) <= not (a and b);
    layer0_outputs(12166) <= 1'b1;
    layer0_outputs(12167) <= not (a or b);
    layer0_outputs(12168) <= not b;
    layer0_outputs(12169) <= a;
    layer0_outputs(12170) <= not (a or b);
    layer0_outputs(12171) <= a xor b;
    layer0_outputs(12172) <= not b or a;
    layer0_outputs(12173) <= not (a and b);
    layer0_outputs(12174) <= a and not b;
    layer0_outputs(12175) <= not (a or b);
    layer0_outputs(12176) <= a or b;
    layer0_outputs(12177) <= not b;
    layer0_outputs(12178) <= not (a or b);
    layer0_outputs(12179) <= not a;
    layer0_outputs(12180) <= not (a or b);
    layer0_outputs(12181) <= a xor b;
    layer0_outputs(12182) <= not b or a;
    layer0_outputs(12183) <= a or b;
    layer0_outputs(12184) <= not b or a;
    layer0_outputs(12185) <= not (a xor b);
    layer0_outputs(12186) <= a xor b;
    layer0_outputs(12187) <= not a;
    layer0_outputs(12188) <= a or b;
    layer0_outputs(12189) <= not a;
    layer0_outputs(12190) <= not a;
    layer0_outputs(12191) <= 1'b0;
    layer0_outputs(12192) <= b and not a;
    layer0_outputs(12193) <= a and not b;
    layer0_outputs(12194) <= a;
    layer0_outputs(12195) <= a and not b;
    layer0_outputs(12196) <= not (a or b);
    layer0_outputs(12197) <= a or b;
    layer0_outputs(12198) <= not (a xor b);
    layer0_outputs(12199) <= b and not a;
    layer0_outputs(12200) <= not b or a;
    layer0_outputs(12201) <= not (a or b);
    layer0_outputs(12202) <= not (a xor b);
    layer0_outputs(12203) <= a;
    layer0_outputs(12204) <= not (a xor b);
    layer0_outputs(12205) <= not b;
    layer0_outputs(12206) <= not a or b;
    layer0_outputs(12207) <= a or b;
    layer0_outputs(12208) <= not (a and b);
    layer0_outputs(12209) <= not b;
    layer0_outputs(12210) <= not (a and b);
    layer0_outputs(12211) <= a and not b;
    layer0_outputs(12212) <= not (a xor b);
    layer0_outputs(12213) <= a and b;
    layer0_outputs(12214) <= a and not b;
    layer0_outputs(12215) <= a;
    layer0_outputs(12216) <= not a;
    layer0_outputs(12217) <= a xor b;
    layer0_outputs(12218) <= a;
    layer0_outputs(12219) <= not b;
    layer0_outputs(12220) <= a xor b;
    layer0_outputs(12221) <= a or b;
    layer0_outputs(12222) <= not b;
    layer0_outputs(12223) <= a or b;
    layer0_outputs(12224) <= not b;
    layer0_outputs(12225) <= not b or a;
    layer0_outputs(12226) <= not (a xor b);
    layer0_outputs(12227) <= not (a xor b);
    layer0_outputs(12228) <= a and not b;
    layer0_outputs(12229) <= not (a or b);
    layer0_outputs(12230) <= a xor b;
    layer0_outputs(12231) <= not (a or b);
    layer0_outputs(12232) <= not b or a;
    layer0_outputs(12233) <= a and not b;
    layer0_outputs(12234) <= b and not a;
    layer0_outputs(12235) <= b and not a;
    layer0_outputs(12236) <= 1'b0;
    layer0_outputs(12237) <= not (a or b);
    layer0_outputs(12238) <= a or b;
    layer0_outputs(12239) <= not b or a;
    layer0_outputs(12240) <= not (a or b);
    layer0_outputs(12241) <= a xor b;
    layer0_outputs(12242) <= not b;
    layer0_outputs(12243) <= not b or a;
    layer0_outputs(12244) <= a or b;
    layer0_outputs(12245) <= a;
    layer0_outputs(12246) <= b;
    layer0_outputs(12247) <= a;
    layer0_outputs(12248) <= not a or b;
    layer0_outputs(12249) <= not (a or b);
    layer0_outputs(12250) <= a;
    layer0_outputs(12251) <= not b;
    layer0_outputs(12252) <= a or b;
    layer0_outputs(12253) <= not (a or b);
    layer0_outputs(12254) <= b and not a;
    layer0_outputs(12255) <= not (a xor b);
    layer0_outputs(12256) <= a xor b;
    layer0_outputs(12257) <= not (a or b);
    layer0_outputs(12258) <= not a;
    layer0_outputs(12259) <= not b;
    layer0_outputs(12260) <= not (a xor b);
    layer0_outputs(12261) <= not a;
    layer0_outputs(12262) <= not (a or b);
    layer0_outputs(12263) <= 1'b1;
    layer0_outputs(12264) <= not b;
    layer0_outputs(12265) <= 1'b1;
    layer0_outputs(12266) <= not (a or b);
    layer0_outputs(12267) <= not (a or b);
    layer0_outputs(12268) <= a;
    layer0_outputs(12269) <= a and not b;
    layer0_outputs(12270) <= not b or a;
    layer0_outputs(12271) <= a xor b;
    layer0_outputs(12272) <= not b or a;
    layer0_outputs(12273) <= a;
    layer0_outputs(12274) <= 1'b0;
    layer0_outputs(12275) <= a and not b;
    layer0_outputs(12276) <= not (a or b);
    layer0_outputs(12277) <= a;
    layer0_outputs(12278) <= a or b;
    layer0_outputs(12279) <= not b or a;
    layer0_outputs(12280) <= b;
    layer0_outputs(12281) <= not a or b;
    layer0_outputs(12282) <= not b or a;
    layer0_outputs(12283) <= b and not a;
    layer0_outputs(12284) <= not (a xor b);
    layer0_outputs(12285) <= a or b;
    layer0_outputs(12286) <= not b or a;
    layer0_outputs(12287) <= not (a or b);
    layer0_outputs(12288) <= a xor b;
    layer0_outputs(12289) <= not (a or b);
    layer0_outputs(12290) <= not (a xor b);
    layer0_outputs(12291) <= a and not b;
    layer0_outputs(12292) <= not b;
    layer0_outputs(12293) <= not a or b;
    layer0_outputs(12294) <= a and b;
    layer0_outputs(12295) <= a or b;
    layer0_outputs(12296) <= not (a xor b);
    layer0_outputs(12297) <= a xor b;
    layer0_outputs(12298) <= a xor b;
    layer0_outputs(12299) <= not (a or b);
    layer0_outputs(12300) <= a and b;
    layer0_outputs(12301) <= b;
    layer0_outputs(12302) <= a;
    layer0_outputs(12303) <= a or b;
    layer0_outputs(12304) <= a;
    layer0_outputs(12305) <= not b;
    layer0_outputs(12306) <= a xor b;
    layer0_outputs(12307) <= a and not b;
    layer0_outputs(12308) <= not (a and b);
    layer0_outputs(12309) <= a or b;
    layer0_outputs(12310) <= b;
    layer0_outputs(12311) <= 1'b0;
    layer0_outputs(12312) <= b;
    layer0_outputs(12313) <= a xor b;
    layer0_outputs(12314) <= b and not a;
    layer0_outputs(12315) <= a xor b;
    layer0_outputs(12316) <= not a;
    layer0_outputs(12317) <= not b;
    layer0_outputs(12318) <= a or b;
    layer0_outputs(12319) <= a and not b;
    layer0_outputs(12320) <= not (a or b);
    layer0_outputs(12321) <= a and not b;
    layer0_outputs(12322) <= a;
    layer0_outputs(12323) <= a or b;
    layer0_outputs(12324) <= a xor b;
    layer0_outputs(12325) <= b;
    layer0_outputs(12326) <= not a;
    layer0_outputs(12327) <= a and not b;
    layer0_outputs(12328) <= not a or b;
    layer0_outputs(12329) <= not b or a;
    layer0_outputs(12330) <= not (a and b);
    layer0_outputs(12331) <= a and b;
    layer0_outputs(12332) <= not a;
    layer0_outputs(12333) <= not (a or b);
    layer0_outputs(12334) <= a or b;
    layer0_outputs(12335) <= a xor b;
    layer0_outputs(12336) <= b;
    layer0_outputs(12337) <= a and not b;
    layer0_outputs(12338) <= not (a or b);
    layer0_outputs(12339) <= not b or a;
    layer0_outputs(12340) <= b;
    layer0_outputs(12341) <= not (a and b);
    layer0_outputs(12342) <= 1'b1;
    layer0_outputs(12343) <= not (a and b);
    layer0_outputs(12344) <= not (a or b);
    layer0_outputs(12345) <= a or b;
    layer0_outputs(12346) <= not (a or b);
    layer0_outputs(12347) <= a xor b;
    layer0_outputs(12348) <= b and not a;
    layer0_outputs(12349) <= not b;
    layer0_outputs(12350) <= a and not b;
    layer0_outputs(12351) <= a;
    layer0_outputs(12352) <= not (a xor b);
    layer0_outputs(12353) <= not a or b;
    layer0_outputs(12354) <= 1'b0;
    layer0_outputs(12355) <= 1'b1;
    layer0_outputs(12356) <= not (a and b);
    layer0_outputs(12357) <= a xor b;
    layer0_outputs(12358) <= 1'b0;
    layer0_outputs(12359) <= not (a or b);
    layer0_outputs(12360) <= b and not a;
    layer0_outputs(12361) <= a or b;
    layer0_outputs(12362) <= a or b;
    layer0_outputs(12363) <= not (a or b);
    layer0_outputs(12364) <= not b or a;
    layer0_outputs(12365) <= not a;
    layer0_outputs(12366) <= not a;
    layer0_outputs(12367) <= not b or a;
    layer0_outputs(12368) <= not a or b;
    layer0_outputs(12369) <= a or b;
    layer0_outputs(12370) <= a and not b;
    layer0_outputs(12371) <= a or b;
    layer0_outputs(12372) <= not a;
    layer0_outputs(12373) <= a or b;
    layer0_outputs(12374) <= not (a or b);
    layer0_outputs(12375) <= not a or b;
    layer0_outputs(12376) <= a xor b;
    layer0_outputs(12377) <= b;
    layer0_outputs(12378) <= 1'b1;
    layer0_outputs(12379) <= not b or a;
    layer0_outputs(12380) <= b;
    layer0_outputs(12381) <= not b or a;
    layer0_outputs(12382) <= a xor b;
    layer0_outputs(12383) <= not a or b;
    layer0_outputs(12384) <= b and not a;
    layer0_outputs(12385) <= a and not b;
    layer0_outputs(12386) <= not (a or b);
    layer0_outputs(12387) <= not a;
    layer0_outputs(12388) <= a and not b;
    layer0_outputs(12389) <= not (a xor b);
    layer0_outputs(12390) <= not (a xor b);
    layer0_outputs(12391) <= 1'b1;
    layer0_outputs(12392) <= a xor b;
    layer0_outputs(12393) <= a;
    layer0_outputs(12394) <= b and not a;
    layer0_outputs(12395) <= a or b;
    layer0_outputs(12396) <= not b or a;
    layer0_outputs(12397) <= a and not b;
    layer0_outputs(12398) <= a and not b;
    layer0_outputs(12399) <= not (a or b);
    layer0_outputs(12400) <= not a;
    layer0_outputs(12401) <= not (a xor b);
    layer0_outputs(12402) <= a and not b;
    layer0_outputs(12403) <= a;
    layer0_outputs(12404) <= a and not b;
    layer0_outputs(12405) <= not b;
    layer0_outputs(12406) <= not (a xor b);
    layer0_outputs(12407) <= not (a or b);
    layer0_outputs(12408) <= not b;
    layer0_outputs(12409) <= a;
    layer0_outputs(12410) <= a or b;
    layer0_outputs(12411) <= b and not a;
    layer0_outputs(12412) <= not a or b;
    layer0_outputs(12413) <= not (a or b);
    layer0_outputs(12414) <= b and not a;
    layer0_outputs(12415) <= b;
    layer0_outputs(12416) <= not b;
    layer0_outputs(12417) <= a xor b;
    layer0_outputs(12418) <= a;
    layer0_outputs(12419) <= not a or b;
    layer0_outputs(12420) <= b and not a;
    layer0_outputs(12421) <= not b;
    layer0_outputs(12422) <= 1'b0;
    layer0_outputs(12423) <= a and not b;
    layer0_outputs(12424) <= b and not a;
    layer0_outputs(12425) <= a or b;
    layer0_outputs(12426) <= a;
    layer0_outputs(12427) <= not (a or b);
    layer0_outputs(12428) <= not b or a;
    layer0_outputs(12429) <= b and not a;
    layer0_outputs(12430) <= not (a xor b);
    layer0_outputs(12431) <= not (a xor b);
    layer0_outputs(12432) <= not b;
    layer0_outputs(12433) <= b and not a;
    layer0_outputs(12434) <= b;
    layer0_outputs(12435) <= b and not a;
    layer0_outputs(12436) <= a or b;
    layer0_outputs(12437) <= 1'b1;
    layer0_outputs(12438) <= a;
    layer0_outputs(12439) <= not a or b;
    layer0_outputs(12440) <= not a or b;
    layer0_outputs(12441) <= a and not b;
    layer0_outputs(12442) <= a or b;
    layer0_outputs(12443) <= b;
    layer0_outputs(12444) <= b;
    layer0_outputs(12445) <= a or b;
    layer0_outputs(12446) <= not (a and b);
    layer0_outputs(12447) <= a xor b;
    layer0_outputs(12448) <= a xor b;
    layer0_outputs(12449) <= 1'b1;
    layer0_outputs(12450) <= not (a and b);
    layer0_outputs(12451) <= a and b;
    layer0_outputs(12452) <= not (a or b);
    layer0_outputs(12453) <= not (a and b);
    layer0_outputs(12454) <= a and b;
    layer0_outputs(12455) <= a;
    layer0_outputs(12456) <= b and not a;
    layer0_outputs(12457) <= a xor b;
    layer0_outputs(12458) <= not (a xor b);
    layer0_outputs(12459) <= a;
    layer0_outputs(12460) <= not b;
    layer0_outputs(12461) <= not a;
    layer0_outputs(12462) <= not a;
    layer0_outputs(12463) <= a or b;
    layer0_outputs(12464) <= a and not b;
    layer0_outputs(12465) <= not (a xor b);
    layer0_outputs(12466) <= not b;
    layer0_outputs(12467) <= b;
    layer0_outputs(12468) <= not (a xor b);
    layer0_outputs(12469) <= a xor b;
    layer0_outputs(12470) <= not a or b;
    layer0_outputs(12471) <= not a or b;
    layer0_outputs(12472) <= not b;
    layer0_outputs(12473) <= not (a and b);
    layer0_outputs(12474) <= not (a or b);
    layer0_outputs(12475) <= not a;
    layer0_outputs(12476) <= a and not b;
    layer0_outputs(12477) <= a and not b;
    layer0_outputs(12478) <= 1'b1;
    layer0_outputs(12479) <= not a;
    layer0_outputs(12480) <= not b or a;
    layer0_outputs(12481) <= a or b;
    layer0_outputs(12482) <= b and not a;
    layer0_outputs(12483) <= not (a or b);
    layer0_outputs(12484) <= a and not b;
    layer0_outputs(12485) <= a and b;
    layer0_outputs(12486) <= a;
    layer0_outputs(12487) <= a;
    layer0_outputs(12488) <= not a or b;
    layer0_outputs(12489) <= not b;
    layer0_outputs(12490) <= a or b;
    layer0_outputs(12491) <= 1'b1;
    layer0_outputs(12492) <= a;
    layer0_outputs(12493) <= a xor b;
    layer0_outputs(12494) <= not a or b;
    layer0_outputs(12495) <= not (a or b);
    layer0_outputs(12496) <= a;
    layer0_outputs(12497) <= b and not a;
    layer0_outputs(12498) <= a or b;
    layer0_outputs(12499) <= b;
    layer0_outputs(12500) <= not (a xor b);
    layer0_outputs(12501) <= a xor b;
    layer0_outputs(12502) <= a;
    layer0_outputs(12503) <= not (a or b);
    layer0_outputs(12504) <= a or b;
    layer0_outputs(12505) <= not (a xor b);
    layer0_outputs(12506) <= not b;
    layer0_outputs(12507) <= b and not a;
    layer0_outputs(12508) <= b;
    layer0_outputs(12509) <= b;
    layer0_outputs(12510) <= a or b;
    layer0_outputs(12511) <= a or b;
    layer0_outputs(12512) <= a and not b;
    layer0_outputs(12513) <= b;
    layer0_outputs(12514) <= a and not b;
    layer0_outputs(12515) <= not (a or b);
    layer0_outputs(12516) <= a xor b;
    layer0_outputs(12517) <= not b or a;
    layer0_outputs(12518) <= b;
    layer0_outputs(12519) <= a;
    layer0_outputs(12520) <= a and not b;
    layer0_outputs(12521) <= not a or b;
    layer0_outputs(12522) <= not (a xor b);
    layer0_outputs(12523) <= 1'b1;
    layer0_outputs(12524) <= a;
    layer0_outputs(12525) <= a and not b;
    layer0_outputs(12526) <= a;
    layer0_outputs(12527) <= a xor b;
    layer0_outputs(12528) <= not (a and b);
    layer0_outputs(12529) <= a xor b;
    layer0_outputs(12530) <= a or b;
    layer0_outputs(12531) <= 1'b1;
    layer0_outputs(12532) <= not b;
    layer0_outputs(12533) <= a or b;
    layer0_outputs(12534) <= b and not a;
    layer0_outputs(12535) <= 1'b1;
    layer0_outputs(12536) <= not (a or b);
    layer0_outputs(12537) <= b;
    layer0_outputs(12538) <= a and not b;
    layer0_outputs(12539) <= not b or a;
    layer0_outputs(12540) <= b and not a;
    layer0_outputs(12541) <= not (a or b);
    layer0_outputs(12542) <= not (a xor b);
    layer0_outputs(12543) <= not b;
    layer0_outputs(12544) <= a or b;
    layer0_outputs(12545) <= not a;
    layer0_outputs(12546) <= b and not a;
    layer0_outputs(12547) <= a xor b;
    layer0_outputs(12548) <= a or b;
    layer0_outputs(12549) <= not (a and b);
    layer0_outputs(12550) <= not (a or b);
    layer0_outputs(12551) <= not (a xor b);
    layer0_outputs(12552) <= not b;
    layer0_outputs(12553) <= a xor b;
    layer0_outputs(12554) <= a or b;
    layer0_outputs(12555) <= a or b;
    layer0_outputs(12556) <= a;
    layer0_outputs(12557) <= not (a xor b);
    layer0_outputs(12558) <= not b;
    layer0_outputs(12559) <= a or b;
    layer0_outputs(12560) <= not a;
    layer0_outputs(12561) <= not a;
    layer0_outputs(12562) <= not b or a;
    layer0_outputs(12563) <= a xor b;
    layer0_outputs(12564) <= b and not a;
    layer0_outputs(12565) <= not b or a;
    layer0_outputs(12566) <= not (a and b);
    layer0_outputs(12567) <= not (a xor b);
    layer0_outputs(12568) <= not (a or b);
    layer0_outputs(12569) <= not b or a;
    layer0_outputs(12570) <= not (a and b);
    layer0_outputs(12571) <= a and not b;
    layer0_outputs(12572) <= not (a or b);
    layer0_outputs(12573) <= not b or a;
    layer0_outputs(12574) <= a or b;
    layer0_outputs(12575) <= b;
    layer0_outputs(12576) <= a xor b;
    layer0_outputs(12577) <= not a or b;
    layer0_outputs(12578) <= b and not a;
    layer0_outputs(12579) <= not b or a;
    layer0_outputs(12580) <= a;
    layer0_outputs(12581) <= not a;
    layer0_outputs(12582) <= a and not b;
    layer0_outputs(12583) <= not a;
    layer0_outputs(12584) <= a or b;
    layer0_outputs(12585) <= not b;
    layer0_outputs(12586) <= not (a or b);
    layer0_outputs(12587) <= not b;
    layer0_outputs(12588) <= b and not a;
    layer0_outputs(12589) <= not (a and b);
    layer0_outputs(12590) <= not (a xor b);
    layer0_outputs(12591) <= a or b;
    layer0_outputs(12592) <= not b or a;
    layer0_outputs(12593) <= a or b;
    layer0_outputs(12594) <= not b;
    layer0_outputs(12595) <= not (a or b);
    layer0_outputs(12596) <= not (a xor b);
    layer0_outputs(12597) <= not (a or b);
    layer0_outputs(12598) <= a xor b;
    layer0_outputs(12599) <= not (a or b);
    layer0_outputs(12600) <= not a or b;
    layer0_outputs(12601) <= not a;
    layer0_outputs(12602) <= not (a xor b);
    layer0_outputs(12603) <= 1'b0;
    layer0_outputs(12604) <= a;
    layer0_outputs(12605) <= not (a xor b);
    layer0_outputs(12606) <= b and not a;
    layer0_outputs(12607) <= not a;
    layer0_outputs(12608) <= not b;
    layer0_outputs(12609) <= not b;
    layer0_outputs(12610) <= not b or a;
    layer0_outputs(12611) <= not a;
    layer0_outputs(12612) <= a or b;
    layer0_outputs(12613) <= 1'b1;
    layer0_outputs(12614) <= 1'b0;
    layer0_outputs(12615) <= not b;
    layer0_outputs(12616) <= b and not a;
    layer0_outputs(12617) <= not a or b;
    layer0_outputs(12618) <= b;
    layer0_outputs(12619) <= not (a xor b);
    layer0_outputs(12620) <= a;
    layer0_outputs(12621) <= not b or a;
    layer0_outputs(12622) <= not (a xor b);
    layer0_outputs(12623) <= b;
    layer0_outputs(12624) <= a;
    layer0_outputs(12625) <= a or b;
    layer0_outputs(12626) <= not b;
    layer0_outputs(12627) <= b and not a;
    layer0_outputs(12628) <= b;
    layer0_outputs(12629) <= a xor b;
    layer0_outputs(12630) <= b;
    layer0_outputs(12631) <= not b or a;
    layer0_outputs(12632) <= a or b;
    layer0_outputs(12633) <= a and not b;
    layer0_outputs(12634) <= not b or a;
    layer0_outputs(12635) <= not (a and b);
    layer0_outputs(12636) <= b;
    layer0_outputs(12637) <= not (a xor b);
    layer0_outputs(12638) <= a or b;
    layer0_outputs(12639) <= not b;
    layer0_outputs(12640) <= a xor b;
    layer0_outputs(12641) <= a;
    layer0_outputs(12642) <= not b;
    layer0_outputs(12643) <= b and not a;
    layer0_outputs(12644) <= not (a or b);
    layer0_outputs(12645) <= b and not a;
    layer0_outputs(12646) <= a;
    layer0_outputs(12647) <= not b or a;
    layer0_outputs(12648) <= b;
    layer0_outputs(12649) <= not (a or b);
    layer0_outputs(12650) <= not (a xor b);
    layer0_outputs(12651) <= not a;
    layer0_outputs(12652) <= b and not a;
    layer0_outputs(12653) <= b;
    layer0_outputs(12654) <= not a;
    layer0_outputs(12655) <= not a or b;
    layer0_outputs(12656) <= a or b;
    layer0_outputs(12657) <= not (a or b);
    layer0_outputs(12658) <= not b;
    layer0_outputs(12659) <= a;
    layer0_outputs(12660) <= not b or a;
    layer0_outputs(12661) <= not b or a;
    layer0_outputs(12662) <= a and b;
    layer0_outputs(12663) <= a and b;
    layer0_outputs(12664) <= not (a and b);
    layer0_outputs(12665) <= not (a and b);
    layer0_outputs(12666) <= not a or b;
    layer0_outputs(12667) <= b and not a;
    layer0_outputs(12668) <= b;
    layer0_outputs(12669) <= not a or b;
    layer0_outputs(12670) <= b and not a;
    layer0_outputs(12671) <= not a or b;
    layer0_outputs(12672) <= not b;
    layer0_outputs(12673) <= not (a xor b);
    layer0_outputs(12674) <= a xor b;
    layer0_outputs(12675) <= b and not a;
    layer0_outputs(12676) <= not a or b;
    layer0_outputs(12677) <= a and not b;
    layer0_outputs(12678) <= a or b;
    layer0_outputs(12679) <= 1'b1;
    layer0_outputs(12680) <= b and not a;
    layer0_outputs(12681) <= a and not b;
    layer0_outputs(12682) <= not (a xor b);
    layer0_outputs(12683) <= not b;
    layer0_outputs(12684) <= not a;
    layer0_outputs(12685) <= not a or b;
    layer0_outputs(12686) <= b;
    layer0_outputs(12687) <= not a;
    layer0_outputs(12688) <= not a or b;
    layer0_outputs(12689) <= not b or a;
    layer0_outputs(12690) <= 1'b1;
    layer0_outputs(12691) <= not (a or b);
    layer0_outputs(12692) <= not (a or b);
    layer0_outputs(12693) <= a or b;
    layer0_outputs(12694) <= not a;
    layer0_outputs(12695) <= not b or a;
    layer0_outputs(12696) <= not b;
    layer0_outputs(12697) <= a xor b;
    layer0_outputs(12698) <= not (a or b);
    layer0_outputs(12699) <= a or b;
    layer0_outputs(12700) <= not (a xor b);
    layer0_outputs(12701) <= not (a and b);
    layer0_outputs(12702) <= not b;
    layer0_outputs(12703) <= a xor b;
    layer0_outputs(12704) <= a or b;
    layer0_outputs(12705) <= not b or a;
    layer0_outputs(12706) <= not b or a;
    layer0_outputs(12707) <= a xor b;
    layer0_outputs(12708) <= a or b;
    layer0_outputs(12709) <= b and not a;
    layer0_outputs(12710) <= not a or b;
    layer0_outputs(12711) <= b;
    layer0_outputs(12712) <= not (a xor b);
    layer0_outputs(12713) <= not b;
    layer0_outputs(12714) <= a and b;
    layer0_outputs(12715) <= not (a or b);
    layer0_outputs(12716) <= not b or a;
    layer0_outputs(12717) <= a;
    layer0_outputs(12718) <= not b;
    layer0_outputs(12719) <= a;
    layer0_outputs(12720) <= not (a xor b);
    layer0_outputs(12721) <= b;
    layer0_outputs(12722) <= not (a or b);
    layer0_outputs(12723) <= a xor b;
    layer0_outputs(12724) <= b;
    layer0_outputs(12725) <= not (a or b);
    layer0_outputs(12726) <= not (a or b);
    layer0_outputs(12727) <= a;
    layer0_outputs(12728) <= 1'b1;
    layer0_outputs(12729) <= not (a xor b);
    layer0_outputs(12730) <= not b or a;
    layer0_outputs(12731) <= not (a or b);
    layer0_outputs(12732) <= not (a and b);
    layer0_outputs(12733) <= not (a or b);
    layer0_outputs(12734) <= not b or a;
    layer0_outputs(12735) <= not b or a;
    layer0_outputs(12736) <= b;
    layer0_outputs(12737) <= a;
    layer0_outputs(12738) <= 1'b0;
    layer0_outputs(12739) <= not (a xor b);
    layer0_outputs(12740) <= not (a xor b);
    layer0_outputs(12741) <= not (a or b);
    layer0_outputs(12742) <= a xor b;
    layer0_outputs(12743) <= not (a xor b);
    layer0_outputs(12744) <= b;
    layer0_outputs(12745) <= a and not b;
    layer0_outputs(12746) <= 1'b1;
    layer0_outputs(12747) <= a xor b;
    layer0_outputs(12748) <= 1'b1;
    layer0_outputs(12749) <= 1'b1;
    layer0_outputs(12750) <= a or b;
    layer0_outputs(12751) <= b;
    layer0_outputs(12752) <= b;
    layer0_outputs(12753) <= a;
    layer0_outputs(12754) <= a xor b;
    layer0_outputs(12755) <= not b;
    layer0_outputs(12756) <= not (a or b);
    layer0_outputs(12757) <= not a or b;
    layer0_outputs(12758) <= a xor b;
    layer0_outputs(12759) <= a xor b;
    layer0_outputs(12760) <= a and not b;
    layer0_outputs(12761) <= b;
    layer0_outputs(12762) <= 1'b1;
    layer0_outputs(12763) <= a xor b;
    layer0_outputs(12764) <= b;
    layer0_outputs(12765) <= not a;
    layer0_outputs(12766) <= not (a xor b);
    layer0_outputs(12767) <= a xor b;
    layer0_outputs(12768) <= not b;
    layer0_outputs(12769) <= not b;
    layer0_outputs(12770) <= not a or b;
    layer0_outputs(12771) <= b;
    layer0_outputs(12772) <= a or b;
    layer0_outputs(12773) <= a and b;
    layer0_outputs(12774) <= not (a or b);
    layer0_outputs(12775) <= not a or b;
    layer0_outputs(12776) <= not (a xor b);
    layer0_outputs(12777) <= a xor b;
    layer0_outputs(12778) <= b;
    layer0_outputs(12779) <= not (a or b);
    layer0_outputs(12780) <= not a or b;
    layer0_outputs(12781) <= not (a xor b);
    layer0_outputs(12782) <= 1'b0;
    layer0_outputs(12783) <= a xor b;
    layer0_outputs(12784) <= b;
    layer0_outputs(12785) <= not (a xor b);
    layer0_outputs(12786) <= not b or a;
    layer0_outputs(12787) <= a xor b;
    layer0_outputs(12788) <= not b or a;
    layer0_outputs(12789) <= not b;
    layer0_outputs(12790) <= a;
    layer0_outputs(12791) <= a;
    layer0_outputs(12792) <= not (a xor b);
    layer0_outputs(12793) <= not (a xor b);
    layer0_outputs(12794) <= not (a xor b);
    layer0_outputs(12795) <= a;
    layer0_outputs(12796) <= not (a or b);
    layer0_outputs(12797) <= not a;
    layer0_outputs(12798) <= not (a xor b);
    layer0_outputs(12799) <= not (a or b);
    layer1_outputs(0) <= a or b;
    layer1_outputs(1) <= b and not a;
    layer1_outputs(2) <= b and not a;
    layer1_outputs(3) <= not (a and b);
    layer1_outputs(4) <= not (a xor b);
    layer1_outputs(5) <= not (a xor b);
    layer1_outputs(6) <= 1'b0;
    layer1_outputs(7) <= b;
    layer1_outputs(8) <= not (a or b);
    layer1_outputs(9) <= a xor b;
    layer1_outputs(10) <= not a;
    layer1_outputs(11) <= a and not b;
    layer1_outputs(12) <= b;
    layer1_outputs(13) <= not (a or b);
    layer1_outputs(14) <= not a or b;
    layer1_outputs(15) <= 1'b1;
    layer1_outputs(16) <= not a;
    layer1_outputs(17) <= a and not b;
    layer1_outputs(18) <= not (a xor b);
    layer1_outputs(19) <= a or b;
    layer1_outputs(20) <= a or b;
    layer1_outputs(21) <= not a or b;
    layer1_outputs(22) <= not a;
    layer1_outputs(23) <= a or b;
    layer1_outputs(24) <= b;
    layer1_outputs(25) <= b and not a;
    layer1_outputs(26) <= b;
    layer1_outputs(27) <= 1'b1;
    layer1_outputs(28) <= not (a xor b);
    layer1_outputs(29) <= a xor b;
    layer1_outputs(30) <= b;
    layer1_outputs(31) <= not (a xor b);
    layer1_outputs(32) <= b and not a;
    layer1_outputs(33) <= not a;
    layer1_outputs(34) <= b;
    layer1_outputs(35) <= not b or a;
    layer1_outputs(36) <= not (a or b);
    layer1_outputs(37) <= a and b;
    layer1_outputs(38) <= b and not a;
    layer1_outputs(39) <= not a;
    layer1_outputs(40) <= a or b;
    layer1_outputs(41) <= not a;
    layer1_outputs(42) <= not (a xor b);
    layer1_outputs(43) <= not (a or b);
    layer1_outputs(44) <= a;
    layer1_outputs(45) <= a;
    layer1_outputs(46) <= not (a xor b);
    layer1_outputs(47) <= not (a xor b);
    layer1_outputs(48) <= not b or a;
    layer1_outputs(49) <= not a;
    layer1_outputs(50) <= not a or b;
    layer1_outputs(51) <= a and not b;
    layer1_outputs(52) <= a;
    layer1_outputs(53) <= not (a or b);
    layer1_outputs(54) <= b;
    layer1_outputs(55) <= not b;
    layer1_outputs(56) <= not (a or b);
    layer1_outputs(57) <= not (a xor b);
    layer1_outputs(58) <= not (a xor b);
    layer1_outputs(59) <= a and b;
    layer1_outputs(60) <= a xor b;
    layer1_outputs(61) <= a or b;
    layer1_outputs(62) <= b and not a;
    layer1_outputs(63) <= not a or b;
    layer1_outputs(64) <= a and b;
    layer1_outputs(65) <= a xor b;
    layer1_outputs(66) <= a;
    layer1_outputs(67) <= not a;
    layer1_outputs(68) <= a or b;
    layer1_outputs(69) <= not a or b;
    layer1_outputs(70) <= a;
    layer1_outputs(71) <= a;
    layer1_outputs(72) <= a and not b;
    layer1_outputs(73) <= b;
    layer1_outputs(74) <= not b;
    layer1_outputs(75) <= not b;
    layer1_outputs(76) <= not (a xor b);
    layer1_outputs(77) <= not a;
    layer1_outputs(78) <= b;
    layer1_outputs(79) <= not a;
    layer1_outputs(80) <= not (a xor b);
    layer1_outputs(81) <= not a;
    layer1_outputs(82) <= not (a or b);
    layer1_outputs(83) <= not (a xor b);
    layer1_outputs(84) <= not b or a;
    layer1_outputs(85) <= b and not a;
    layer1_outputs(86) <= not a;
    layer1_outputs(87) <= not a;
    layer1_outputs(88) <= b and not a;
    layer1_outputs(89) <= not a;
    layer1_outputs(90) <= not b or a;
    layer1_outputs(91) <= not b;
    layer1_outputs(92) <= b;
    layer1_outputs(93) <= not b or a;
    layer1_outputs(94) <= not a;
    layer1_outputs(95) <= a;
    layer1_outputs(96) <= b and not a;
    layer1_outputs(97) <= a and b;
    layer1_outputs(98) <= not a or b;
    layer1_outputs(99) <= not a or b;
    layer1_outputs(100) <= a and b;
    layer1_outputs(101) <= not (a and b);
    layer1_outputs(102) <= b;
    layer1_outputs(103) <= not a or b;
    layer1_outputs(104) <= not (a xor b);
    layer1_outputs(105) <= a and not b;
    layer1_outputs(106) <= a;
    layer1_outputs(107) <= not b or a;
    layer1_outputs(108) <= a or b;
    layer1_outputs(109) <= b and not a;
    layer1_outputs(110) <= a xor b;
    layer1_outputs(111) <= not b;
    layer1_outputs(112) <= not b or a;
    layer1_outputs(113) <= not a;
    layer1_outputs(114) <= 1'b1;
    layer1_outputs(115) <= not (a and b);
    layer1_outputs(116) <= 1'b0;
    layer1_outputs(117) <= a and not b;
    layer1_outputs(118) <= b;
    layer1_outputs(119) <= a or b;
    layer1_outputs(120) <= a;
    layer1_outputs(121) <= not b;
    layer1_outputs(122) <= not (a and b);
    layer1_outputs(123) <= 1'b0;
    layer1_outputs(124) <= a and not b;
    layer1_outputs(125) <= not (a or b);
    layer1_outputs(126) <= not b or a;
    layer1_outputs(127) <= 1'b0;
    layer1_outputs(128) <= not a;
    layer1_outputs(129) <= not a or b;
    layer1_outputs(130) <= not b;
    layer1_outputs(131) <= b and not a;
    layer1_outputs(132) <= a and not b;
    layer1_outputs(133) <= not (a and b);
    layer1_outputs(134) <= b and not a;
    layer1_outputs(135) <= b;
    layer1_outputs(136) <= a xor b;
    layer1_outputs(137) <= a or b;
    layer1_outputs(138) <= a and not b;
    layer1_outputs(139) <= a xor b;
    layer1_outputs(140) <= a;
    layer1_outputs(141) <= a or b;
    layer1_outputs(142) <= not b or a;
    layer1_outputs(143) <= not (a xor b);
    layer1_outputs(144) <= not a or b;
    layer1_outputs(145) <= not a;
    layer1_outputs(146) <= a;
    layer1_outputs(147) <= not b or a;
    layer1_outputs(148) <= a and b;
    layer1_outputs(149) <= not (a and b);
    layer1_outputs(150) <= not (a or b);
    layer1_outputs(151) <= b and not a;
    layer1_outputs(152) <= not b;
    layer1_outputs(153) <= a xor b;
    layer1_outputs(154) <= not b;
    layer1_outputs(155) <= not (a or b);
    layer1_outputs(156) <= not a or b;
    layer1_outputs(157) <= a and not b;
    layer1_outputs(158) <= not b;
    layer1_outputs(159) <= not (a xor b);
    layer1_outputs(160) <= a;
    layer1_outputs(161) <= not a;
    layer1_outputs(162) <= not b;
    layer1_outputs(163) <= a;
    layer1_outputs(164) <= b;
    layer1_outputs(165) <= b and not a;
    layer1_outputs(166) <= a xor b;
    layer1_outputs(167) <= not b;
    layer1_outputs(168) <= a xor b;
    layer1_outputs(169) <= a;
    layer1_outputs(170) <= not (a xor b);
    layer1_outputs(171) <= not (a xor b);
    layer1_outputs(172) <= not (a xor b);
    layer1_outputs(173) <= a and not b;
    layer1_outputs(174) <= a and b;
    layer1_outputs(175) <= not b or a;
    layer1_outputs(176) <= a and b;
    layer1_outputs(177) <= not (a or b);
    layer1_outputs(178) <= a and not b;
    layer1_outputs(179) <= not (a or b);
    layer1_outputs(180) <= a;
    layer1_outputs(181) <= a xor b;
    layer1_outputs(182) <= not a;
    layer1_outputs(183) <= a;
    layer1_outputs(184) <= not (a xor b);
    layer1_outputs(185) <= not (a and b);
    layer1_outputs(186) <= not a or b;
    layer1_outputs(187) <= not a;
    layer1_outputs(188) <= not (a or b);
    layer1_outputs(189) <= not (a or b);
    layer1_outputs(190) <= b;
    layer1_outputs(191) <= a or b;
    layer1_outputs(192) <= a xor b;
    layer1_outputs(193) <= b;
    layer1_outputs(194) <= not a or b;
    layer1_outputs(195) <= not b;
    layer1_outputs(196) <= b;
    layer1_outputs(197) <= a or b;
    layer1_outputs(198) <= a and not b;
    layer1_outputs(199) <= a and not b;
    layer1_outputs(200) <= b;
    layer1_outputs(201) <= not b;
    layer1_outputs(202) <= a and b;
    layer1_outputs(203) <= not a;
    layer1_outputs(204) <= b and not a;
    layer1_outputs(205) <= b;
    layer1_outputs(206) <= a xor b;
    layer1_outputs(207) <= a and b;
    layer1_outputs(208) <= a xor b;
    layer1_outputs(209) <= not b;
    layer1_outputs(210) <= b;
    layer1_outputs(211) <= not b;
    layer1_outputs(212) <= not (a or b);
    layer1_outputs(213) <= a and b;
    layer1_outputs(214) <= not (a xor b);
    layer1_outputs(215) <= a;
    layer1_outputs(216) <= not a;
    layer1_outputs(217) <= not b;
    layer1_outputs(218) <= not (a and b);
    layer1_outputs(219) <= b;
    layer1_outputs(220) <= not b or a;
    layer1_outputs(221) <= not (a and b);
    layer1_outputs(222) <= not b;
    layer1_outputs(223) <= not b;
    layer1_outputs(224) <= not b;
    layer1_outputs(225) <= not (a and b);
    layer1_outputs(226) <= a;
    layer1_outputs(227) <= not (a and b);
    layer1_outputs(228) <= a xor b;
    layer1_outputs(229) <= not a or b;
    layer1_outputs(230) <= not (a or b);
    layer1_outputs(231) <= not b;
    layer1_outputs(232) <= b;
    layer1_outputs(233) <= a;
    layer1_outputs(234) <= b;
    layer1_outputs(235) <= not a or b;
    layer1_outputs(236) <= 1'b0;
    layer1_outputs(237) <= not a or b;
    layer1_outputs(238) <= not (a or b);
    layer1_outputs(239) <= not a or b;
    layer1_outputs(240) <= not (a or b);
    layer1_outputs(241) <= not b or a;
    layer1_outputs(242) <= a;
    layer1_outputs(243) <= not a;
    layer1_outputs(244) <= a;
    layer1_outputs(245) <= not b or a;
    layer1_outputs(246) <= b;
    layer1_outputs(247) <= not (a and b);
    layer1_outputs(248) <= b and not a;
    layer1_outputs(249) <= not b;
    layer1_outputs(250) <= b;
    layer1_outputs(251) <= not b;
    layer1_outputs(252) <= a xor b;
    layer1_outputs(253) <= b;
    layer1_outputs(254) <= not (a or b);
    layer1_outputs(255) <= not a;
    layer1_outputs(256) <= not a or b;
    layer1_outputs(257) <= a xor b;
    layer1_outputs(258) <= not (a and b);
    layer1_outputs(259) <= b;
    layer1_outputs(260) <= not b;
    layer1_outputs(261) <= b and not a;
    layer1_outputs(262) <= not (a xor b);
    layer1_outputs(263) <= 1'b0;
    layer1_outputs(264) <= not (a xor b);
    layer1_outputs(265) <= not b or a;
    layer1_outputs(266) <= not a;
    layer1_outputs(267) <= a xor b;
    layer1_outputs(268) <= not b;
    layer1_outputs(269) <= not b;
    layer1_outputs(270) <= not b;
    layer1_outputs(271) <= not b or a;
    layer1_outputs(272) <= not b;
    layer1_outputs(273) <= not (a or b);
    layer1_outputs(274) <= not a or b;
    layer1_outputs(275) <= a or b;
    layer1_outputs(276) <= not (a and b);
    layer1_outputs(277) <= not b;
    layer1_outputs(278) <= a and not b;
    layer1_outputs(279) <= a or b;
    layer1_outputs(280) <= a or b;
    layer1_outputs(281) <= b;
    layer1_outputs(282) <= b and not a;
    layer1_outputs(283) <= not b or a;
    layer1_outputs(284) <= not b or a;
    layer1_outputs(285) <= 1'b0;
    layer1_outputs(286) <= not (a xor b);
    layer1_outputs(287) <= not a or b;
    layer1_outputs(288) <= not (a or b);
    layer1_outputs(289) <= not (a xor b);
    layer1_outputs(290) <= not (a and b);
    layer1_outputs(291) <= not a or b;
    layer1_outputs(292) <= a or b;
    layer1_outputs(293) <= not (a xor b);
    layer1_outputs(294) <= not a;
    layer1_outputs(295) <= not a;
    layer1_outputs(296) <= b;
    layer1_outputs(297) <= a or b;
    layer1_outputs(298) <= not (a or b);
    layer1_outputs(299) <= not a;
    layer1_outputs(300) <= not b;
    layer1_outputs(301) <= not a;
    layer1_outputs(302) <= a or b;
    layer1_outputs(303) <= a xor b;
    layer1_outputs(304) <= not (a or b);
    layer1_outputs(305) <= b and not a;
    layer1_outputs(306) <= a;
    layer1_outputs(307) <= a xor b;
    layer1_outputs(308) <= a;
    layer1_outputs(309) <= a xor b;
    layer1_outputs(310) <= b;
    layer1_outputs(311) <= a;
    layer1_outputs(312) <= not (a and b);
    layer1_outputs(313) <= a and b;
    layer1_outputs(314) <= not a;
    layer1_outputs(315) <= not (a xor b);
    layer1_outputs(316) <= not b;
    layer1_outputs(317) <= 1'b0;
    layer1_outputs(318) <= a;
    layer1_outputs(319) <= not b;
    layer1_outputs(320) <= a or b;
    layer1_outputs(321) <= not a or b;
    layer1_outputs(322) <= not (a xor b);
    layer1_outputs(323) <= a and not b;
    layer1_outputs(324) <= a xor b;
    layer1_outputs(325) <= not (a or b);
    layer1_outputs(326) <= not b or a;
    layer1_outputs(327) <= a and not b;
    layer1_outputs(328) <= b;
    layer1_outputs(329) <= not (a xor b);
    layer1_outputs(330) <= not a;
    layer1_outputs(331) <= not (a xor b);
    layer1_outputs(332) <= a xor b;
    layer1_outputs(333) <= 1'b1;
    layer1_outputs(334) <= not b;
    layer1_outputs(335) <= not (a xor b);
    layer1_outputs(336) <= not (a and b);
    layer1_outputs(337) <= a and b;
    layer1_outputs(338) <= not a;
    layer1_outputs(339) <= b and not a;
    layer1_outputs(340) <= not (a or b);
    layer1_outputs(341) <= a;
    layer1_outputs(342) <= a or b;
    layer1_outputs(343) <= a;
    layer1_outputs(344) <= b;
    layer1_outputs(345) <= a and not b;
    layer1_outputs(346) <= not b;
    layer1_outputs(347) <= a;
    layer1_outputs(348) <= not (a and b);
    layer1_outputs(349) <= a and b;
    layer1_outputs(350) <= a and not b;
    layer1_outputs(351) <= a xor b;
    layer1_outputs(352) <= a or b;
    layer1_outputs(353) <= b;
    layer1_outputs(354) <= not b;
    layer1_outputs(355) <= a;
    layer1_outputs(356) <= a xor b;
    layer1_outputs(357) <= not (a and b);
    layer1_outputs(358) <= not (a and b);
    layer1_outputs(359) <= b and not a;
    layer1_outputs(360) <= b;
    layer1_outputs(361) <= a;
    layer1_outputs(362) <= b and not a;
    layer1_outputs(363) <= b;
    layer1_outputs(364) <= not a;
    layer1_outputs(365) <= not b or a;
    layer1_outputs(366) <= not b;
    layer1_outputs(367) <= not (a xor b);
    layer1_outputs(368) <= not a;
    layer1_outputs(369) <= not a;
    layer1_outputs(370) <= not b;
    layer1_outputs(371) <= not (a xor b);
    layer1_outputs(372) <= not a;
    layer1_outputs(373) <= a and b;
    layer1_outputs(374) <= b;
    layer1_outputs(375) <= not b;
    layer1_outputs(376) <= a xor b;
    layer1_outputs(377) <= a and b;
    layer1_outputs(378) <= a;
    layer1_outputs(379) <= 1'b1;
    layer1_outputs(380) <= a xor b;
    layer1_outputs(381) <= a and not b;
    layer1_outputs(382) <= not (a xor b);
    layer1_outputs(383) <= not a;
    layer1_outputs(384) <= not (a xor b);
    layer1_outputs(385) <= a or b;
    layer1_outputs(386) <= a;
    layer1_outputs(387) <= not b;
    layer1_outputs(388) <= not b or a;
    layer1_outputs(389) <= b;
    layer1_outputs(390) <= not b;
    layer1_outputs(391) <= a or b;
    layer1_outputs(392) <= b and not a;
    layer1_outputs(393) <= not a;
    layer1_outputs(394) <= not b or a;
    layer1_outputs(395) <= not b;
    layer1_outputs(396) <= not (a and b);
    layer1_outputs(397) <= not (a xor b);
    layer1_outputs(398) <= a and not b;
    layer1_outputs(399) <= a and not b;
    layer1_outputs(400) <= not b;
    layer1_outputs(401) <= b and not a;
    layer1_outputs(402) <= a;
    layer1_outputs(403) <= not b;
    layer1_outputs(404) <= b and not a;
    layer1_outputs(405) <= a and b;
    layer1_outputs(406) <= b;
    layer1_outputs(407) <= a and not b;
    layer1_outputs(408) <= a;
    layer1_outputs(409) <= a or b;
    layer1_outputs(410) <= not (a xor b);
    layer1_outputs(411) <= not a or b;
    layer1_outputs(412) <= not a;
    layer1_outputs(413) <= not (a xor b);
    layer1_outputs(414) <= a or b;
    layer1_outputs(415) <= not a;
    layer1_outputs(416) <= not a or b;
    layer1_outputs(417) <= not (a or b);
    layer1_outputs(418) <= not a;
    layer1_outputs(419) <= a;
    layer1_outputs(420) <= b and not a;
    layer1_outputs(421) <= not a;
    layer1_outputs(422) <= not b or a;
    layer1_outputs(423) <= not b;
    layer1_outputs(424) <= b;
    layer1_outputs(425) <= not a or b;
    layer1_outputs(426) <= a;
    layer1_outputs(427) <= a or b;
    layer1_outputs(428) <= not b;
    layer1_outputs(429) <= not (a and b);
    layer1_outputs(430) <= a or b;
    layer1_outputs(431) <= b;
    layer1_outputs(432) <= 1'b0;
    layer1_outputs(433) <= not b;
    layer1_outputs(434) <= not b;
    layer1_outputs(435) <= a xor b;
    layer1_outputs(436) <= a and not b;
    layer1_outputs(437) <= a and b;
    layer1_outputs(438) <= not (a xor b);
    layer1_outputs(439) <= not a;
    layer1_outputs(440) <= not (a xor b);
    layer1_outputs(441) <= a or b;
    layer1_outputs(442) <= not a;
    layer1_outputs(443) <= not b;
    layer1_outputs(444) <= not a;
    layer1_outputs(445) <= not (a xor b);
    layer1_outputs(446) <= not b or a;
    layer1_outputs(447) <= a and b;
    layer1_outputs(448) <= not (a xor b);
    layer1_outputs(449) <= not a;
    layer1_outputs(450) <= b;
    layer1_outputs(451) <= a xor b;
    layer1_outputs(452) <= b;
    layer1_outputs(453) <= not a;
    layer1_outputs(454) <= a;
    layer1_outputs(455) <= not b;
    layer1_outputs(456) <= not (a and b);
    layer1_outputs(457) <= not (a xor b);
    layer1_outputs(458) <= a or b;
    layer1_outputs(459) <= not (a or b);
    layer1_outputs(460) <= a and not b;
    layer1_outputs(461) <= not a;
    layer1_outputs(462) <= not (a and b);
    layer1_outputs(463) <= b;
    layer1_outputs(464) <= b;
    layer1_outputs(465) <= a;
    layer1_outputs(466) <= a or b;
    layer1_outputs(467) <= a and b;
    layer1_outputs(468) <= b;
    layer1_outputs(469) <= a or b;
    layer1_outputs(470) <= a;
    layer1_outputs(471) <= not a or b;
    layer1_outputs(472) <= b;
    layer1_outputs(473) <= a;
    layer1_outputs(474) <= a xor b;
    layer1_outputs(475) <= a xor b;
    layer1_outputs(476) <= not b;
    layer1_outputs(477) <= a xor b;
    layer1_outputs(478) <= not a;
    layer1_outputs(479) <= not (a or b);
    layer1_outputs(480) <= a xor b;
    layer1_outputs(481) <= a xor b;
    layer1_outputs(482) <= b and not a;
    layer1_outputs(483) <= 1'b0;
    layer1_outputs(484) <= b and not a;
    layer1_outputs(485) <= b;
    layer1_outputs(486) <= not (a and b);
    layer1_outputs(487) <= a xor b;
    layer1_outputs(488) <= not b or a;
    layer1_outputs(489) <= a;
    layer1_outputs(490) <= a;
    layer1_outputs(491) <= a xor b;
    layer1_outputs(492) <= not a;
    layer1_outputs(493) <= not b or a;
    layer1_outputs(494) <= a;
    layer1_outputs(495) <= not (a and b);
    layer1_outputs(496) <= a and b;
    layer1_outputs(497) <= b;
    layer1_outputs(498) <= 1'b0;
    layer1_outputs(499) <= not a;
    layer1_outputs(500) <= not a or b;
    layer1_outputs(501) <= a xor b;
    layer1_outputs(502) <= not b or a;
    layer1_outputs(503) <= not (a or b);
    layer1_outputs(504) <= b and not a;
    layer1_outputs(505) <= not (a and b);
    layer1_outputs(506) <= not (a xor b);
    layer1_outputs(507) <= a;
    layer1_outputs(508) <= not b or a;
    layer1_outputs(509) <= not a;
    layer1_outputs(510) <= b;
    layer1_outputs(511) <= a and not b;
    layer1_outputs(512) <= not (a and b);
    layer1_outputs(513) <= a;
    layer1_outputs(514) <= not a;
    layer1_outputs(515) <= a and not b;
    layer1_outputs(516) <= not b or a;
    layer1_outputs(517) <= a xor b;
    layer1_outputs(518) <= not (a and b);
    layer1_outputs(519) <= not (a and b);
    layer1_outputs(520) <= a and not b;
    layer1_outputs(521) <= not a;
    layer1_outputs(522) <= not b or a;
    layer1_outputs(523) <= b;
    layer1_outputs(524) <= a;
    layer1_outputs(525) <= not (a or b);
    layer1_outputs(526) <= not (a xor b);
    layer1_outputs(527) <= b;
    layer1_outputs(528) <= not (a xor b);
    layer1_outputs(529) <= a or b;
    layer1_outputs(530) <= not b or a;
    layer1_outputs(531) <= a and not b;
    layer1_outputs(532) <= a;
    layer1_outputs(533) <= not (a xor b);
    layer1_outputs(534) <= b and not a;
    layer1_outputs(535) <= not a or b;
    layer1_outputs(536) <= not (a xor b);
    layer1_outputs(537) <= not b;
    layer1_outputs(538) <= a and not b;
    layer1_outputs(539) <= a;
    layer1_outputs(540) <= not (a and b);
    layer1_outputs(541) <= b;
    layer1_outputs(542) <= b;
    layer1_outputs(543) <= not b;
    layer1_outputs(544) <= not a;
    layer1_outputs(545) <= b;
    layer1_outputs(546) <= not (a and b);
    layer1_outputs(547) <= a and b;
    layer1_outputs(548) <= a;
    layer1_outputs(549) <= not a or b;
    layer1_outputs(550) <= not b;
    layer1_outputs(551) <= not b;
    layer1_outputs(552) <= a;
    layer1_outputs(553) <= not b;
    layer1_outputs(554) <= a or b;
    layer1_outputs(555) <= a;
    layer1_outputs(556) <= not (a or b);
    layer1_outputs(557) <= a or b;
    layer1_outputs(558) <= not (a xor b);
    layer1_outputs(559) <= not b;
    layer1_outputs(560) <= not a;
    layer1_outputs(561) <= a;
    layer1_outputs(562) <= 1'b0;
    layer1_outputs(563) <= b;
    layer1_outputs(564) <= not a;
    layer1_outputs(565) <= not (a or b);
    layer1_outputs(566) <= not a or b;
    layer1_outputs(567) <= a;
    layer1_outputs(568) <= a;
    layer1_outputs(569) <= a and not b;
    layer1_outputs(570) <= a and b;
    layer1_outputs(571) <= not b or a;
    layer1_outputs(572) <= a and b;
    layer1_outputs(573) <= b;
    layer1_outputs(574) <= not b;
    layer1_outputs(575) <= not a or b;
    layer1_outputs(576) <= a xor b;
    layer1_outputs(577) <= not (a xor b);
    layer1_outputs(578) <= a;
    layer1_outputs(579) <= b and not a;
    layer1_outputs(580) <= not (a xor b);
    layer1_outputs(581) <= not (a or b);
    layer1_outputs(582) <= not (a or b);
    layer1_outputs(583) <= a and b;
    layer1_outputs(584) <= a;
    layer1_outputs(585) <= a and not b;
    layer1_outputs(586) <= not b or a;
    layer1_outputs(587) <= a and not b;
    layer1_outputs(588) <= a;
    layer1_outputs(589) <= a xor b;
    layer1_outputs(590) <= b and not a;
    layer1_outputs(591) <= not a or b;
    layer1_outputs(592) <= not b;
    layer1_outputs(593) <= a or b;
    layer1_outputs(594) <= not a or b;
    layer1_outputs(595) <= not a or b;
    layer1_outputs(596) <= a and b;
    layer1_outputs(597) <= a xor b;
    layer1_outputs(598) <= a;
    layer1_outputs(599) <= not (a xor b);
    layer1_outputs(600) <= a or b;
    layer1_outputs(601) <= not b;
    layer1_outputs(602) <= a;
    layer1_outputs(603) <= not b;
    layer1_outputs(604) <= a and not b;
    layer1_outputs(605) <= not b;
    layer1_outputs(606) <= not b;
    layer1_outputs(607) <= not (a xor b);
    layer1_outputs(608) <= not a;
    layer1_outputs(609) <= not (a and b);
    layer1_outputs(610) <= not (a xor b);
    layer1_outputs(611) <= b;
    layer1_outputs(612) <= b;
    layer1_outputs(613) <= not a;
    layer1_outputs(614) <= a or b;
    layer1_outputs(615) <= b and not a;
    layer1_outputs(616) <= not a or b;
    layer1_outputs(617) <= a or b;
    layer1_outputs(618) <= not (a and b);
    layer1_outputs(619) <= not b or a;
    layer1_outputs(620) <= a and b;
    layer1_outputs(621) <= not b;
    layer1_outputs(622) <= a or b;
    layer1_outputs(623) <= not b or a;
    layer1_outputs(624) <= not (a xor b);
    layer1_outputs(625) <= a or b;
    layer1_outputs(626) <= a xor b;
    layer1_outputs(627) <= not b;
    layer1_outputs(628) <= b and not a;
    layer1_outputs(629) <= a xor b;
    layer1_outputs(630) <= b and not a;
    layer1_outputs(631) <= not a;
    layer1_outputs(632) <= not b;
    layer1_outputs(633) <= a and not b;
    layer1_outputs(634) <= not a;
    layer1_outputs(635) <= b and not a;
    layer1_outputs(636) <= a or b;
    layer1_outputs(637) <= a;
    layer1_outputs(638) <= a xor b;
    layer1_outputs(639) <= b;
    layer1_outputs(640) <= not a or b;
    layer1_outputs(641) <= not b;
    layer1_outputs(642) <= b;
    layer1_outputs(643) <= not b or a;
    layer1_outputs(644) <= b;
    layer1_outputs(645) <= not b or a;
    layer1_outputs(646) <= not a or b;
    layer1_outputs(647) <= not a or b;
    layer1_outputs(648) <= b;
    layer1_outputs(649) <= a;
    layer1_outputs(650) <= not b or a;
    layer1_outputs(651) <= a and b;
    layer1_outputs(652) <= 1'b1;
    layer1_outputs(653) <= a;
    layer1_outputs(654) <= a;
    layer1_outputs(655) <= b;
    layer1_outputs(656) <= b;
    layer1_outputs(657) <= a xor b;
    layer1_outputs(658) <= not a or b;
    layer1_outputs(659) <= a xor b;
    layer1_outputs(660) <= not (a or b);
    layer1_outputs(661) <= b;
    layer1_outputs(662) <= b;
    layer1_outputs(663) <= not a or b;
    layer1_outputs(664) <= not b or a;
    layer1_outputs(665) <= not b;
    layer1_outputs(666) <= a xor b;
    layer1_outputs(667) <= b;
    layer1_outputs(668) <= 1'b0;
    layer1_outputs(669) <= not b;
    layer1_outputs(670) <= not b;
    layer1_outputs(671) <= not (a and b);
    layer1_outputs(672) <= a;
    layer1_outputs(673) <= not a;
    layer1_outputs(674) <= a and not b;
    layer1_outputs(675) <= not a;
    layer1_outputs(676) <= a;
    layer1_outputs(677) <= b and not a;
    layer1_outputs(678) <= not a;
    layer1_outputs(679) <= not b or a;
    layer1_outputs(680) <= a and b;
    layer1_outputs(681) <= not b;
    layer1_outputs(682) <= a xor b;
    layer1_outputs(683) <= not (a or b);
    layer1_outputs(684) <= a or b;
    layer1_outputs(685) <= a or b;
    layer1_outputs(686) <= 1'b0;
    layer1_outputs(687) <= b;
    layer1_outputs(688) <= not b or a;
    layer1_outputs(689) <= not a;
    layer1_outputs(690) <= b;
    layer1_outputs(691) <= a;
    layer1_outputs(692) <= a;
    layer1_outputs(693) <= b;
    layer1_outputs(694) <= b;
    layer1_outputs(695) <= b and not a;
    layer1_outputs(696) <= b and not a;
    layer1_outputs(697) <= not b or a;
    layer1_outputs(698) <= a;
    layer1_outputs(699) <= not a;
    layer1_outputs(700) <= not b;
    layer1_outputs(701) <= a xor b;
    layer1_outputs(702) <= not (a xor b);
    layer1_outputs(703) <= not (a and b);
    layer1_outputs(704) <= a and b;
    layer1_outputs(705) <= b and not a;
    layer1_outputs(706) <= not (a xor b);
    layer1_outputs(707) <= b;
    layer1_outputs(708) <= not b or a;
    layer1_outputs(709) <= 1'b0;
    layer1_outputs(710) <= b;
    layer1_outputs(711) <= a xor b;
    layer1_outputs(712) <= a and b;
    layer1_outputs(713) <= 1'b0;
    layer1_outputs(714) <= b and not a;
    layer1_outputs(715) <= not a;
    layer1_outputs(716) <= not a or b;
    layer1_outputs(717) <= not (a or b);
    layer1_outputs(718) <= not (a xor b);
    layer1_outputs(719) <= not (a xor b);
    layer1_outputs(720) <= not (a xor b);
    layer1_outputs(721) <= not b or a;
    layer1_outputs(722) <= not b or a;
    layer1_outputs(723) <= 1'b1;
    layer1_outputs(724) <= b;
    layer1_outputs(725) <= not (a and b);
    layer1_outputs(726) <= not a;
    layer1_outputs(727) <= not b;
    layer1_outputs(728) <= not (a and b);
    layer1_outputs(729) <= 1'b0;
    layer1_outputs(730) <= b and not a;
    layer1_outputs(731) <= b;
    layer1_outputs(732) <= a or b;
    layer1_outputs(733) <= not a;
    layer1_outputs(734) <= a;
    layer1_outputs(735) <= not b;
    layer1_outputs(736) <= a;
    layer1_outputs(737) <= b;
    layer1_outputs(738) <= a;
    layer1_outputs(739) <= a xor b;
    layer1_outputs(740) <= not a or b;
    layer1_outputs(741) <= b;
    layer1_outputs(742) <= a and not b;
    layer1_outputs(743) <= not (a xor b);
    layer1_outputs(744) <= not (a xor b);
    layer1_outputs(745) <= not b or a;
    layer1_outputs(746) <= a xor b;
    layer1_outputs(747) <= a xor b;
    layer1_outputs(748) <= b;
    layer1_outputs(749) <= not a;
    layer1_outputs(750) <= a xor b;
    layer1_outputs(751) <= b;
    layer1_outputs(752) <= a and not b;
    layer1_outputs(753) <= not b;
    layer1_outputs(754) <= a;
    layer1_outputs(755) <= b;
    layer1_outputs(756) <= not a;
    layer1_outputs(757) <= b and not a;
    layer1_outputs(758) <= a or b;
    layer1_outputs(759) <= not b;
    layer1_outputs(760) <= a;
    layer1_outputs(761) <= b and not a;
    layer1_outputs(762) <= a;
    layer1_outputs(763) <= b;
    layer1_outputs(764) <= not (a or b);
    layer1_outputs(765) <= not a or b;
    layer1_outputs(766) <= not (a and b);
    layer1_outputs(767) <= not b;
    layer1_outputs(768) <= not b or a;
    layer1_outputs(769) <= not (a xor b);
    layer1_outputs(770) <= b and not a;
    layer1_outputs(771) <= not a;
    layer1_outputs(772) <= not b or a;
    layer1_outputs(773) <= 1'b1;
    layer1_outputs(774) <= a or b;
    layer1_outputs(775) <= b and not a;
    layer1_outputs(776) <= not (a xor b);
    layer1_outputs(777) <= b and not a;
    layer1_outputs(778) <= b;
    layer1_outputs(779) <= not a;
    layer1_outputs(780) <= not (a and b);
    layer1_outputs(781) <= a;
    layer1_outputs(782) <= a and b;
    layer1_outputs(783) <= a and b;
    layer1_outputs(784) <= a;
    layer1_outputs(785) <= not b;
    layer1_outputs(786) <= b;
    layer1_outputs(787) <= not a;
    layer1_outputs(788) <= not b;
    layer1_outputs(789) <= b;
    layer1_outputs(790) <= b and not a;
    layer1_outputs(791) <= a xor b;
    layer1_outputs(792) <= not a;
    layer1_outputs(793) <= not a;
    layer1_outputs(794) <= not (a and b);
    layer1_outputs(795) <= not a;
    layer1_outputs(796) <= a and b;
    layer1_outputs(797) <= a and b;
    layer1_outputs(798) <= a and not b;
    layer1_outputs(799) <= a;
    layer1_outputs(800) <= not (a xor b);
    layer1_outputs(801) <= a xor b;
    layer1_outputs(802) <= a xor b;
    layer1_outputs(803) <= not (a or b);
    layer1_outputs(804) <= not (a or b);
    layer1_outputs(805) <= not b;
    layer1_outputs(806) <= not a;
    layer1_outputs(807) <= a or b;
    layer1_outputs(808) <= not a or b;
    layer1_outputs(809) <= a and b;
    layer1_outputs(810) <= a;
    layer1_outputs(811) <= not (a xor b);
    layer1_outputs(812) <= not a;
    layer1_outputs(813) <= b;
    layer1_outputs(814) <= a;
    layer1_outputs(815) <= not b;
    layer1_outputs(816) <= a xor b;
    layer1_outputs(817) <= b;
    layer1_outputs(818) <= not (a xor b);
    layer1_outputs(819) <= not b or a;
    layer1_outputs(820) <= not (a and b);
    layer1_outputs(821) <= not b or a;
    layer1_outputs(822) <= not (a or b);
    layer1_outputs(823) <= a and not b;
    layer1_outputs(824) <= not a or b;
    layer1_outputs(825) <= b;
    layer1_outputs(826) <= not (a xor b);
    layer1_outputs(827) <= not a;
    layer1_outputs(828) <= not b;
    layer1_outputs(829) <= a and b;
    layer1_outputs(830) <= not a;
    layer1_outputs(831) <= 1'b0;
    layer1_outputs(832) <= a or b;
    layer1_outputs(833) <= not a;
    layer1_outputs(834) <= a and not b;
    layer1_outputs(835) <= not a;
    layer1_outputs(836) <= not (a xor b);
    layer1_outputs(837) <= 1'b1;
    layer1_outputs(838) <= not (a or b);
    layer1_outputs(839) <= not (a and b);
    layer1_outputs(840) <= a or b;
    layer1_outputs(841) <= a xor b;
    layer1_outputs(842) <= not b or a;
    layer1_outputs(843) <= not (a and b);
    layer1_outputs(844) <= a and b;
    layer1_outputs(845) <= not b or a;
    layer1_outputs(846) <= a and not b;
    layer1_outputs(847) <= not (a or b);
    layer1_outputs(848) <= a;
    layer1_outputs(849) <= a xor b;
    layer1_outputs(850) <= not a;
    layer1_outputs(851) <= b;
    layer1_outputs(852) <= a xor b;
    layer1_outputs(853) <= b and not a;
    layer1_outputs(854) <= a xor b;
    layer1_outputs(855) <= a and b;
    layer1_outputs(856) <= a or b;
    layer1_outputs(857) <= a xor b;
    layer1_outputs(858) <= a;
    layer1_outputs(859) <= not (a xor b);
    layer1_outputs(860) <= not a;
    layer1_outputs(861) <= a xor b;
    layer1_outputs(862) <= a and b;
    layer1_outputs(863) <= a xor b;
    layer1_outputs(864) <= a and b;
    layer1_outputs(865) <= not a;
    layer1_outputs(866) <= not (a or b);
    layer1_outputs(867) <= a;
    layer1_outputs(868) <= a or b;
    layer1_outputs(869) <= a;
    layer1_outputs(870) <= a;
    layer1_outputs(871) <= b and not a;
    layer1_outputs(872) <= not b or a;
    layer1_outputs(873) <= not (a xor b);
    layer1_outputs(874) <= not (a xor b);
    layer1_outputs(875) <= a;
    layer1_outputs(876) <= a or b;
    layer1_outputs(877) <= not b or a;
    layer1_outputs(878) <= a xor b;
    layer1_outputs(879) <= not (a xor b);
    layer1_outputs(880) <= not b or a;
    layer1_outputs(881) <= not b;
    layer1_outputs(882) <= a;
    layer1_outputs(883) <= a and b;
    layer1_outputs(884) <= a xor b;
    layer1_outputs(885) <= a and b;
    layer1_outputs(886) <= not (a or b);
    layer1_outputs(887) <= not b;
    layer1_outputs(888) <= not (a or b);
    layer1_outputs(889) <= not b;
    layer1_outputs(890) <= not b;
    layer1_outputs(891) <= b;
    layer1_outputs(892) <= a;
    layer1_outputs(893) <= a and b;
    layer1_outputs(894) <= 1'b1;
    layer1_outputs(895) <= a;
    layer1_outputs(896) <= not a or b;
    layer1_outputs(897) <= b;
    layer1_outputs(898) <= not (a and b);
    layer1_outputs(899) <= a and not b;
    layer1_outputs(900) <= a;
    layer1_outputs(901) <= not a;
    layer1_outputs(902) <= not (a xor b);
    layer1_outputs(903) <= not b or a;
    layer1_outputs(904) <= a and not b;
    layer1_outputs(905) <= a and b;
    layer1_outputs(906) <= a;
    layer1_outputs(907) <= b;
    layer1_outputs(908) <= not (a or b);
    layer1_outputs(909) <= not b;
    layer1_outputs(910) <= not b or a;
    layer1_outputs(911) <= b;
    layer1_outputs(912) <= b;
    layer1_outputs(913) <= not b;
    layer1_outputs(914) <= not (a xor b);
    layer1_outputs(915) <= a xor b;
    layer1_outputs(916) <= a;
    layer1_outputs(917) <= b;
    layer1_outputs(918) <= not a;
    layer1_outputs(919) <= b and not a;
    layer1_outputs(920) <= not a;
    layer1_outputs(921) <= b;
    layer1_outputs(922) <= b;
    layer1_outputs(923) <= 1'b0;
    layer1_outputs(924) <= not a;
    layer1_outputs(925) <= a and b;
    layer1_outputs(926) <= not a or b;
    layer1_outputs(927) <= a and not b;
    layer1_outputs(928) <= a and b;
    layer1_outputs(929) <= b;
    layer1_outputs(930) <= a and not b;
    layer1_outputs(931) <= b;
    layer1_outputs(932) <= not a or b;
    layer1_outputs(933) <= b;
    layer1_outputs(934) <= a xor b;
    layer1_outputs(935) <= a;
    layer1_outputs(936) <= b;
    layer1_outputs(937) <= b;
    layer1_outputs(938) <= not (a xor b);
    layer1_outputs(939) <= not a or b;
    layer1_outputs(940) <= a xor b;
    layer1_outputs(941) <= a xor b;
    layer1_outputs(942) <= a xor b;
    layer1_outputs(943) <= 1'b0;
    layer1_outputs(944) <= a or b;
    layer1_outputs(945) <= a and not b;
    layer1_outputs(946) <= not (a or b);
    layer1_outputs(947) <= a;
    layer1_outputs(948) <= not (a and b);
    layer1_outputs(949) <= not (a or b);
    layer1_outputs(950) <= not b or a;
    layer1_outputs(951) <= not b;
    layer1_outputs(952) <= a xor b;
    layer1_outputs(953) <= b;
    layer1_outputs(954) <= not (a or b);
    layer1_outputs(955) <= not (a xor b);
    layer1_outputs(956) <= not b;
    layer1_outputs(957) <= not b;
    layer1_outputs(958) <= a or b;
    layer1_outputs(959) <= not b;
    layer1_outputs(960) <= not (a and b);
    layer1_outputs(961) <= a xor b;
    layer1_outputs(962) <= not b or a;
    layer1_outputs(963) <= not b or a;
    layer1_outputs(964) <= a xor b;
    layer1_outputs(965) <= b;
    layer1_outputs(966) <= not b;
    layer1_outputs(967) <= b and not a;
    layer1_outputs(968) <= a;
    layer1_outputs(969) <= not b;
    layer1_outputs(970) <= not (a and b);
    layer1_outputs(971) <= a;
    layer1_outputs(972) <= not a or b;
    layer1_outputs(973) <= b and not a;
    layer1_outputs(974) <= 1'b1;
    layer1_outputs(975) <= a;
    layer1_outputs(976) <= a and not b;
    layer1_outputs(977) <= not (a xor b);
    layer1_outputs(978) <= not a;
    layer1_outputs(979) <= a;
    layer1_outputs(980) <= a xor b;
    layer1_outputs(981) <= a;
    layer1_outputs(982) <= b and not a;
    layer1_outputs(983) <= a and b;
    layer1_outputs(984) <= a;
    layer1_outputs(985) <= not a;
    layer1_outputs(986) <= not a;
    layer1_outputs(987) <= not (a xor b);
    layer1_outputs(988) <= not (a xor b);
    layer1_outputs(989) <= b and not a;
    layer1_outputs(990) <= b;
    layer1_outputs(991) <= not (a and b);
    layer1_outputs(992) <= a;
    layer1_outputs(993) <= a xor b;
    layer1_outputs(994) <= a or b;
    layer1_outputs(995) <= a and not b;
    layer1_outputs(996) <= b;
    layer1_outputs(997) <= a;
    layer1_outputs(998) <= b and not a;
    layer1_outputs(999) <= not a or b;
    layer1_outputs(1000) <= a and b;
    layer1_outputs(1001) <= a and b;
    layer1_outputs(1002) <= b and not a;
    layer1_outputs(1003) <= not (a xor b);
    layer1_outputs(1004) <= not (a and b);
    layer1_outputs(1005) <= b;
    layer1_outputs(1006) <= not b;
    layer1_outputs(1007) <= not (a xor b);
    layer1_outputs(1008) <= a and not b;
    layer1_outputs(1009) <= not a;
    layer1_outputs(1010) <= not a;
    layer1_outputs(1011) <= not (a or b);
    layer1_outputs(1012) <= not (a and b);
    layer1_outputs(1013) <= not (a xor b);
    layer1_outputs(1014) <= 1'b1;
    layer1_outputs(1015) <= a xor b;
    layer1_outputs(1016) <= not (a xor b);
    layer1_outputs(1017) <= a and b;
    layer1_outputs(1018) <= not (a xor b);
    layer1_outputs(1019) <= b and not a;
    layer1_outputs(1020) <= a;
    layer1_outputs(1021) <= a or b;
    layer1_outputs(1022) <= a or b;
    layer1_outputs(1023) <= a;
    layer1_outputs(1024) <= not (a or b);
    layer1_outputs(1025) <= a;
    layer1_outputs(1026) <= not (a or b);
    layer1_outputs(1027) <= a and b;
    layer1_outputs(1028) <= a and b;
    layer1_outputs(1029) <= not b or a;
    layer1_outputs(1030) <= 1'b1;
    layer1_outputs(1031) <= b and not a;
    layer1_outputs(1032) <= not (a and b);
    layer1_outputs(1033) <= a;
    layer1_outputs(1034) <= not a or b;
    layer1_outputs(1035) <= a or b;
    layer1_outputs(1036) <= not (a xor b);
    layer1_outputs(1037) <= not (a and b);
    layer1_outputs(1038) <= b;
    layer1_outputs(1039) <= not a;
    layer1_outputs(1040) <= not a;
    layer1_outputs(1041) <= not a or b;
    layer1_outputs(1042) <= a or b;
    layer1_outputs(1043) <= not a or b;
    layer1_outputs(1044) <= not (a xor b);
    layer1_outputs(1045) <= not (a xor b);
    layer1_outputs(1046) <= not (a and b);
    layer1_outputs(1047) <= a and b;
    layer1_outputs(1048) <= a or b;
    layer1_outputs(1049) <= a;
    layer1_outputs(1050) <= a or b;
    layer1_outputs(1051) <= not (a xor b);
    layer1_outputs(1052) <= not (a or b);
    layer1_outputs(1053) <= not a;
    layer1_outputs(1054) <= not a;
    layer1_outputs(1055) <= not (a xor b);
    layer1_outputs(1056) <= b and not a;
    layer1_outputs(1057) <= not a;
    layer1_outputs(1058) <= b;
    layer1_outputs(1059) <= a and b;
    layer1_outputs(1060) <= not a;
    layer1_outputs(1061) <= not (a and b);
    layer1_outputs(1062) <= not (a xor b);
    layer1_outputs(1063) <= b and not a;
    layer1_outputs(1064) <= not a or b;
    layer1_outputs(1065) <= 1'b0;
    layer1_outputs(1066) <= not (a and b);
    layer1_outputs(1067) <= not b;
    layer1_outputs(1068) <= a or b;
    layer1_outputs(1069) <= b and not a;
    layer1_outputs(1070) <= not a or b;
    layer1_outputs(1071) <= a;
    layer1_outputs(1072) <= not (a and b);
    layer1_outputs(1073) <= not a;
    layer1_outputs(1074) <= not b or a;
    layer1_outputs(1075) <= not a;
    layer1_outputs(1076) <= a and not b;
    layer1_outputs(1077) <= b;
    layer1_outputs(1078) <= a xor b;
    layer1_outputs(1079) <= not (a xor b);
    layer1_outputs(1080) <= not (a and b);
    layer1_outputs(1081) <= not a;
    layer1_outputs(1082) <= not (a xor b);
    layer1_outputs(1083) <= not b;
    layer1_outputs(1084) <= b and not a;
    layer1_outputs(1085) <= a and not b;
    layer1_outputs(1086) <= a and b;
    layer1_outputs(1087) <= not (a xor b);
    layer1_outputs(1088) <= not a or b;
    layer1_outputs(1089) <= not (a xor b);
    layer1_outputs(1090) <= a xor b;
    layer1_outputs(1091) <= a xor b;
    layer1_outputs(1092) <= not a or b;
    layer1_outputs(1093) <= a and b;
    layer1_outputs(1094) <= not b or a;
    layer1_outputs(1095) <= b and not a;
    layer1_outputs(1096) <= a or b;
    layer1_outputs(1097) <= not b or a;
    layer1_outputs(1098) <= b;
    layer1_outputs(1099) <= a or b;
    layer1_outputs(1100) <= not a;
    layer1_outputs(1101) <= a;
    layer1_outputs(1102) <= not b;
    layer1_outputs(1103) <= b;
    layer1_outputs(1104) <= a and b;
    layer1_outputs(1105) <= b;
    layer1_outputs(1106) <= not (a and b);
    layer1_outputs(1107) <= a or b;
    layer1_outputs(1108) <= not (a xor b);
    layer1_outputs(1109) <= not a;
    layer1_outputs(1110) <= 1'b1;
    layer1_outputs(1111) <= a xor b;
    layer1_outputs(1112) <= not (a xor b);
    layer1_outputs(1113) <= b;
    layer1_outputs(1114) <= not a;
    layer1_outputs(1115) <= not (a xor b);
    layer1_outputs(1116) <= not b or a;
    layer1_outputs(1117) <= a and not b;
    layer1_outputs(1118) <= a and not b;
    layer1_outputs(1119) <= a and not b;
    layer1_outputs(1120) <= not b or a;
    layer1_outputs(1121) <= not a or b;
    layer1_outputs(1122) <= a and b;
    layer1_outputs(1123) <= b;
    layer1_outputs(1124) <= a;
    layer1_outputs(1125) <= 1'b0;
    layer1_outputs(1126) <= b;
    layer1_outputs(1127) <= not b;
    layer1_outputs(1128) <= not (a or b);
    layer1_outputs(1129) <= 1'b1;
    layer1_outputs(1130) <= not (a and b);
    layer1_outputs(1131) <= b;
    layer1_outputs(1132) <= not (a or b);
    layer1_outputs(1133) <= not b or a;
    layer1_outputs(1134) <= not b;
    layer1_outputs(1135) <= not b or a;
    layer1_outputs(1136) <= not b;
    layer1_outputs(1137) <= a and not b;
    layer1_outputs(1138) <= a;
    layer1_outputs(1139) <= not (a or b);
    layer1_outputs(1140) <= b;
    layer1_outputs(1141) <= not b;
    layer1_outputs(1142) <= not (a xor b);
    layer1_outputs(1143) <= a and b;
    layer1_outputs(1144) <= not a;
    layer1_outputs(1145) <= a and not b;
    layer1_outputs(1146) <= a;
    layer1_outputs(1147) <= not b;
    layer1_outputs(1148) <= a and not b;
    layer1_outputs(1149) <= b;
    layer1_outputs(1150) <= not (a xor b);
    layer1_outputs(1151) <= a or b;
    layer1_outputs(1152) <= not (a and b);
    layer1_outputs(1153) <= not a or b;
    layer1_outputs(1154) <= not b or a;
    layer1_outputs(1155) <= not a;
    layer1_outputs(1156) <= a and b;
    layer1_outputs(1157) <= a xor b;
    layer1_outputs(1158) <= not a or b;
    layer1_outputs(1159) <= a;
    layer1_outputs(1160) <= not (a xor b);
    layer1_outputs(1161) <= a and not b;
    layer1_outputs(1162) <= not (a and b);
    layer1_outputs(1163) <= not (a xor b);
    layer1_outputs(1164) <= a and b;
    layer1_outputs(1165) <= not a;
    layer1_outputs(1166) <= not b;
    layer1_outputs(1167) <= not b or a;
    layer1_outputs(1168) <= not (a xor b);
    layer1_outputs(1169) <= not b or a;
    layer1_outputs(1170) <= b;
    layer1_outputs(1171) <= b;
    layer1_outputs(1172) <= a;
    layer1_outputs(1173) <= a xor b;
    layer1_outputs(1174) <= not a;
    layer1_outputs(1175) <= b;
    layer1_outputs(1176) <= not (a xor b);
    layer1_outputs(1177) <= a xor b;
    layer1_outputs(1178) <= not a;
    layer1_outputs(1179) <= not a or b;
    layer1_outputs(1180) <= a xor b;
    layer1_outputs(1181) <= not (a or b);
    layer1_outputs(1182) <= b and not a;
    layer1_outputs(1183) <= a;
    layer1_outputs(1184) <= not a or b;
    layer1_outputs(1185) <= a and b;
    layer1_outputs(1186) <= b;
    layer1_outputs(1187) <= b;
    layer1_outputs(1188) <= not a;
    layer1_outputs(1189) <= not b or a;
    layer1_outputs(1190) <= not (a or b);
    layer1_outputs(1191) <= not (a and b);
    layer1_outputs(1192) <= not a;
    layer1_outputs(1193) <= not b;
    layer1_outputs(1194) <= b and not a;
    layer1_outputs(1195) <= a or b;
    layer1_outputs(1196) <= not (a xor b);
    layer1_outputs(1197) <= not (a and b);
    layer1_outputs(1198) <= not b or a;
    layer1_outputs(1199) <= not a;
    layer1_outputs(1200) <= not b;
    layer1_outputs(1201) <= not (a xor b);
    layer1_outputs(1202) <= a or b;
    layer1_outputs(1203) <= not (a and b);
    layer1_outputs(1204) <= a and b;
    layer1_outputs(1205) <= not b;
    layer1_outputs(1206) <= not (a and b);
    layer1_outputs(1207) <= not (a xor b);
    layer1_outputs(1208) <= not (a or b);
    layer1_outputs(1209) <= b;
    layer1_outputs(1210) <= a xor b;
    layer1_outputs(1211) <= b and not a;
    layer1_outputs(1212) <= a and b;
    layer1_outputs(1213) <= a and not b;
    layer1_outputs(1214) <= a;
    layer1_outputs(1215) <= not b or a;
    layer1_outputs(1216) <= not (a xor b);
    layer1_outputs(1217) <= b and not a;
    layer1_outputs(1218) <= not a or b;
    layer1_outputs(1219) <= not a or b;
    layer1_outputs(1220) <= not (a xor b);
    layer1_outputs(1221) <= b;
    layer1_outputs(1222) <= b and not a;
    layer1_outputs(1223) <= a and not b;
    layer1_outputs(1224) <= not b;
    layer1_outputs(1225) <= a;
    layer1_outputs(1226) <= not (a or b);
    layer1_outputs(1227) <= b;
    layer1_outputs(1228) <= not b or a;
    layer1_outputs(1229) <= a;
    layer1_outputs(1230) <= a;
    layer1_outputs(1231) <= a and b;
    layer1_outputs(1232) <= not (a xor b);
    layer1_outputs(1233) <= a and not b;
    layer1_outputs(1234) <= not (a and b);
    layer1_outputs(1235) <= a and b;
    layer1_outputs(1236) <= a xor b;
    layer1_outputs(1237) <= not a;
    layer1_outputs(1238) <= not a or b;
    layer1_outputs(1239) <= not b;
    layer1_outputs(1240) <= a;
    layer1_outputs(1241) <= a xor b;
    layer1_outputs(1242) <= not b;
    layer1_outputs(1243) <= not b;
    layer1_outputs(1244) <= b and not a;
    layer1_outputs(1245) <= a;
    layer1_outputs(1246) <= a xor b;
    layer1_outputs(1247) <= not b or a;
    layer1_outputs(1248) <= a or b;
    layer1_outputs(1249) <= not b or a;
    layer1_outputs(1250) <= a and not b;
    layer1_outputs(1251) <= not (a and b);
    layer1_outputs(1252) <= a;
    layer1_outputs(1253) <= a xor b;
    layer1_outputs(1254) <= not (a and b);
    layer1_outputs(1255) <= b;
    layer1_outputs(1256) <= a;
    layer1_outputs(1257) <= not (a xor b);
    layer1_outputs(1258) <= a or b;
    layer1_outputs(1259) <= not b or a;
    layer1_outputs(1260) <= not (a xor b);
    layer1_outputs(1261) <= a xor b;
    layer1_outputs(1262) <= a xor b;
    layer1_outputs(1263) <= a and not b;
    layer1_outputs(1264) <= a;
    layer1_outputs(1265) <= not (a xor b);
    layer1_outputs(1266) <= not (a and b);
    layer1_outputs(1267) <= not (a xor b);
    layer1_outputs(1268) <= not a;
    layer1_outputs(1269) <= not a;
    layer1_outputs(1270) <= not a;
    layer1_outputs(1271) <= b;
    layer1_outputs(1272) <= b;
    layer1_outputs(1273) <= a xor b;
    layer1_outputs(1274) <= b;
    layer1_outputs(1275) <= not a or b;
    layer1_outputs(1276) <= a and not b;
    layer1_outputs(1277) <= a;
    layer1_outputs(1278) <= not (a and b);
    layer1_outputs(1279) <= a;
    layer1_outputs(1280) <= b and not a;
    layer1_outputs(1281) <= not a;
    layer1_outputs(1282) <= not (a xor b);
    layer1_outputs(1283) <= b;
    layer1_outputs(1284) <= a and not b;
    layer1_outputs(1285) <= not (a and b);
    layer1_outputs(1286) <= not (a and b);
    layer1_outputs(1287) <= a or b;
    layer1_outputs(1288) <= a and b;
    layer1_outputs(1289) <= a;
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= not (a and b);
    layer1_outputs(1292) <= not a or b;
    layer1_outputs(1293) <= b;
    layer1_outputs(1294) <= not (a and b);
    layer1_outputs(1295) <= a or b;
    layer1_outputs(1296) <= a and not b;
    layer1_outputs(1297) <= b and not a;
    layer1_outputs(1298) <= a and b;
    layer1_outputs(1299) <= not b;
    layer1_outputs(1300) <= a;
    layer1_outputs(1301) <= a xor b;
    layer1_outputs(1302) <= not (a and b);
    layer1_outputs(1303) <= not (a and b);
    layer1_outputs(1304) <= not b or a;
    layer1_outputs(1305) <= a xor b;
    layer1_outputs(1306) <= not b;
    layer1_outputs(1307) <= a;
    layer1_outputs(1308) <= a xor b;
    layer1_outputs(1309) <= b;
    layer1_outputs(1310) <= not b;
    layer1_outputs(1311) <= not (a xor b);
    layer1_outputs(1312) <= a xor b;
    layer1_outputs(1313) <= a;
    layer1_outputs(1314) <= not (a or b);
    layer1_outputs(1315) <= not b;
    layer1_outputs(1316) <= a and b;
    layer1_outputs(1317) <= a and b;
    layer1_outputs(1318) <= not a;
    layer1_outputs(1319) <= not (a and b);
    layer1_outputs(1320) <= not (a and b);
    layer1_outputs(1321) <= not b;
    layer1_outputs(1322) <= b and not a;
    layer1_outputs(1323) <= not b;
    layer1_outputs(1324) <= not (a or b);
    layer1_outputs(1325) <= b;
    layer1_outputs(1326) <= 1'b1;
    layer1_outputs(1327) <= not b;
    layer1_outputs(1328) <= a xor b;
    layer1_outputs(1329) <= not b;
    layer1_outputs(1330) <= a or b;
    layer1_outputs(1331) <= not a;
    layer1_outputs(1332) <= not a;
    layer1_outputs(1333) <= a and b;
    layer1_outputs(1334) <= not (a xor b);
    layer1_outputs(1335) <= b and not a;
    layer1_outputs(1336) <= b;
    layer1_outputs(1337) <= a and not b;
    layer1_outputs(1338) <= not b or a;
    layer1_outputs(1339) <= not (a or b);
    layer1_outputs(1340) <= not a or b;
    layer1_outputs(1341) <= not (a and b);
    layer1_outputs(1342) <= b and not a;
    layer1_outputs(1343) <= not b;
    layer1_outputs(1344) <= a;
    layer1_outputs(1345) <= a;
    layer1_outputs(1346) <= a or b;
    layer1_outputs(1347) <= not a;
    layer1_outputs(1348) <= not (a and b);
    layer1_outputs(1349) <= not (a or b);
    layer1_outputs(1350) <= a or b;
    layer1_outputs(1351) <= not a;
    layer1_outputs(1352) <= not a or b;
    layer1_outputs(1353) <= not b;
    layer1_outputs(1354) <= b and not a;
    layer1_outputs(1355) <= a;
    layer1_outputs(1356) <= a or b;
    layer1_outputs(1357) <= not b;
    layer1_outputs(1358) <= a;
    layer1_outputs(1359) <= a xor b;
    layer1_outputs(1360) <= a or b;
    layer1_outputs(1361) <= a xor b;
    layer1_outputs(1362) <= a and b;
    layer1_outputs(1363) <= b;
    layer1_outputs(1364) <= not b;
    layer1_outputs(1365) <= a and not b;
    layer1_outputs(1366) <= not b or a;
    layer1_outputs(1367) <= not (a or b);
    layer1_outputs(1368) <= not (a and b);
    layer1_outputs(1369) <= not (a or b);
    layer1_outputs(1370) <= not (a xor b);
    layer1_outputs(1371) <= not b;
    layer1_outputs(1372) <= b and not a;
    layer1_outputs(1373) <= not (a xor b);
    layer1_outputs(1374) <= not (a and b);
    layer1_outputs(1375) <= a;
    layer1_outputs(1376) <= a;
    layer1_outputs(1377) <= b;
    layer1_outputs(1378) <= not a;
    layer1_outputs(1379) <= a xor b;
    layer1_outputs(1380) <= a and not b;
    layer1_outputs(1381) <= not b or a;
    layer1_outputs(1382) <= not b;
    layer1_outputs(1383) <= a or b;
    layer1_outputs(1384) <= not (a xor b);
    layer1_outputs(1385) <= not a;
    layer1_outputs(1386) <= a xor b;
    layer1_outputs(1387) <= not b;
    layer1_outputs(1388) <= 1'b0;
    layer1_outputs(1389) <= not (a or b);
    layer1_outputs(1390) <= not b;
    layer1_outputs(1391) <= b and not a;
    layer1_outputs(1392) <= not b or a;
    layer1_outputs(1393) <= a or b;
    layer1_outputs(1394) <= b;
    layer1_outputs(1395) <= not b;
    layer1_outputs(1396) <= not b or a;
    layer1_outputs(1397) <= not a;
    layer1_outputs(1398) <= not b;
    layer1_outputs(1399) <= not (a xor b);
    layer1_outputs(1400) <= not a or b;
    layer1_outputs(1401) <= not b;
    layer1_outputs(1402) <= not b;
    layer1_outputs(1403) <= a or b;
    layer1_outputs(1404) <= not (a xor b);
    layer1_outputs(1405) <= not b;
    layer1_outputs(1406) <= not (a xor b);
    layer1_outputs(1407) <= not (a xor b);
    layer1_outputs(1408) <= not b;
    layer1_outputs(1409) <= a xor b;
    layer1_outputs(1410) <= b;
    layer1_outputs(1411) <= not b;
    layer1_outputs(1412) <= a xor b;
    layer1_outputs(1413) <= a;
    layer1_outputs(1414) <= not (a or b);
    layer1_outputs(1415) <= not (a or b);
    layer1_outputs(1416) <= not (a or b);
    layer1_outputs(1417) <= not a;
    layer1_outputs(1418) <= not a;
    layer1_outputs(1419) <= not a;
    layer1_outputs(1420) <= not a or b;
    layer1_outputs(1421) <= not b;
    layer1_outputs(1422) <= a;
    layer1_outputs(1423) <= b;
    layer1_outputs(1424) <= not a or b;
    layer1_outputs(1425) <= not a;
    layer1_outputs(1426) <= a and not b;
    layer1_outputs(1427) <= b;
    layer1_outputs(1428) <= not (a and b);
    layer1_outputs(1429) <= b;
    layer1_outputs(1430) <= b;
    layer1_outputs(1431) <= not b;
    layer1_outputs(1432) <= not a;
    layer1_outputs(1433) <= not (a and b);
    layer1_outputs(1434) <= a xor b;
    layer1_outputs(1435) <= not a or b;
    layer1_outputs(1436) <= a and b;
    layer1_outputs(1437) <= b;
    layer1_outputs(1438) <= a xor b;
    layer1_outputs(1439) <= not (a xor b);
    layer1_outputs(1440) <= not a or b;
    layer1_outputs(1441) <= a xor b;
    layer1_outputs(1442) <= not b;
    layer1_outputs(1443) <= a and b;
    layer1_outputs(1444) <= b;
    layer1_outputs(1445) <= not a;
    layer1_outputs(1446) <= not (a or b);
    layer1_outputs(1447) <= not (a xor b);
    layer1_outputs(1448) <= not (a xor b);
    layer1_outputs(1449) <= not (a xor b);
    layer1_outputs(1450) <= b;
    layer1_outputs(1451) <= 1'b0;
    layer1_outputs(1452) <= a and not b;
    layer1_outputs(1453) <= b;
    layer1_outputs(1454) <= a;
    layer1_outputs(1455) <= a;
    layer1_outputs(1456) <= a and b;
    layer1_outputs(1457) <= b and not a;
    layer1_outputs(1458) <= not (a and b);
    layer1_outputs(1459) <= a or b;
    layer1_outputs(1460) <= not b or a;
    layer1_outputs(1461) <= a xor b;
    layer1_outputs(1462) <= not a;
    layer1_outputs(1463) <= not (a or b);
    layer1_outputs(1464) <= a or b;
    layer1_outputs(1465) <= b;
    layer1_outputs(1466) <= not a;
    layer1_outputs(1467) <= not b or a;
    layer1_outputs(1468) <= a xor b;
    layer1_outputs(1469) <= not (a and b);
    layer1_outputs(1470) <= not (a and b);
    layer1_outputs(1471) <= not a;
    layer1_outputs(1472) <= a and not b;
    layer1_outputs(1473) <= a xor b;
    layer1_outputs(1474) <= a and b;
    layer1_outputs(1475) <= a xor b;
    layer1_outputs(1476) <= 1'b0;
    layer1_outputs(1477) <= not (a xor b);
    layer1_outputs(1478) <= b and not a;
    layer1_outputs(1479) <= a xor b;
    layer1_outputs(1480) <= a;
    layer1_outputs(1481) <= 1'b1;
    layer1_outputs(1482) <= a and b;
    layer1_outputs(1483) <= not (a xor b);
    layer1_outputs(1484) <= b;
    layer1_outputs(1485) <= not (a and b);
    layer1_outputs(1486) <= not b;
    layer1_outputs(1487) <= a xor b;
    layer1_outputs(1488) <= not b or a;
    layer1_outputs(1489) <= not b or a;
    layer1_outputs(1490) <= not (a and b);
    layer1_outputs(1491) <= not (a xor b);
    layer1_outputs(1492) <= a and not b;
    layer1_outputs(1493) <= not (a or b);
    layer1_outputs(1494) <= not a or b;
    layer1_outputs(1495) <= not (a and b);
    layer1_outputs(1496) <= not (a xor b);
    layer1_outputs(1497) <= not a or b;
    layer1_outputs(1498) <= a and b;
    layer1_outputs(1499) <= a;
    layer1_outputs(1500) <= not b;
    layer1_outputs(1501) <= a;
    layer1_outputs(1502) <= b;
    layer1_outputs(1503) <= not b;
    layer1_outputs(1504) <= a and not b;
    layer1_outputs(1505) <= b;
    layer1_outputs(1506) <= not (a xor b);
    layer1_outputs(1507) <= b;
    layer1_outputs(1508) <= 1'b1;
    layer1_outputs(1509) <= not a;
    layer1_outputs(1510) <= b;
    layer1_outputs(1511) <= not a;
    layer1_outputs(1512) <= not a or b;
    layer1_outputs(1513) <= a xor b;
    layer1_outputs(1514) <= b;
    layer1_outputs(1515) <= a and not b;
    layer1_outputs(1516) <= not a or b;
    layer1_outputs(1517) <= a;
    layer1_outputs(1518) <= not a or b;
    layer1_outputs(1519) <= not a;
    layer1_outputs(1520) <= not a or b;
    layer1_outputs(1521) <= not b;
    layer1_outputs(1522) <= not (a xor b);
    layer1_outputs(1523) <= a;
    layer1_outputs(1524) <= a and not b;
    layer1_outputs(1525) <= not b;
    layer1_outputs(1526) <= a xor b;
    layer1_outputs(1527) <= not (a xor b);
    layer1_outputs(1528) <= not (a and b);
    layer1_outputs(1529) <= a and b;
    layer1_outputs(1530) <= not a or b;
    layer1_outputs(1531) <= b;
    layer1_outputs(1532) <= not b;
    layer1_outputs(1533) <= b;
    layer1_outputs(1534) <= not (a and b);
    layer1_outputs(1535) <= b and not a;
    layer1_outputs(1536) <= not a;
    layer1_outputs(1537) <= b;
    layer1_outputs(1538) <= a;
    layer1_outputs(1539) <= not b;
    layer1_outputs(1540) <= not b or a;
    layer1_outputs(1541) <= a and b;
    layer1_outputs(1542) <= a xor b;
    layer1_outputs(1543) <= b and not a;
    layer1_outputs(1544) <= 1'b1;
    layer1_outputs(1545) <= not (a xor b);
    layer1_outputs(1546) <= a xor b;
    layer1_outputs(1547) <= not a or b;
    layer1_outputs(1548) <= not (a or b);
    layer1_outputs(1549) <= not a;
    layer1_outputs(1550) <= not a or b;
    layer1_outputs(1551) <= not a or b;
    layer1_outputs(1552) <= a;
    layer1_outputs(1553) <= not b;
    layer1_outputs(1554) <= b and not a;
    layer1_outputs(1555) <= b and not a;
    layer1_outputs(1556) <= a xor b;
    layer1_outputs(1557) <= not a;
    layer1_outputs(1558) <= not (a xor b);
    layer1_outputs(1559) <= not a;
    layer1_outputs(1560) <= not a;
    layer1_outputs(1561) <= a;
    layer1_outputs(1562) <= a and b;
    layer1_outputs(1563) <= b;
    layer1_outputs(1564) <= a xor b;
    layer1_outputs(1565) <= not a or b;
    layer1_outputs(1566) <= a and b;
    layer1_outputs(1567) <= a and b;
    layer1_outputs(1568) <= b;
    layer1_outputs(1569) <= not b or a;
    layer1_outputs(1570) <= a and b;
    layer1_outputs(1571) <= a and not b;
    layer1_outputs(1572) <= a xor b;
    layer1_outputs(1573) <= not (a or b);
    layer1_outputs(1574) <= a and not b;
    layer1_outputs(1575) <= a xor b;
    layer1_outputs(1576) <= a;
    layer1_outputs(1577) <= not b or a;
    layer1_outputs(1578) <= a and not b;
    layer1_outputs(1579) <= a and not b;
    layer1_outputs(1580) <= b;
    layer1_outputs(1581) <= not (a or b);
    layer1_outputs(1582) <= not (a or b);
    layer1_outputs(1583) <= not b or a;
    layer1_outputs(1584) <= a and b;
    layer1_outputs(1585) <= a;
    layer1_outputs(1586) <= not a or b;
    layer1_outputs(1587) <= 1'b1;
    layer1_outputs(1588) <= a and b;
    layer1_outputs(1589) <= not (a or b);
    layer1_outputs(1590) <= a and b;
    layer1_outputs(1591) <= b and not a;
    layer1_outputs(1592) <= not b or a;
    layer1_outputs(1593) <= a;
    layer1_outputs(1594) <= b and not a;
    layer1_outputs(1595) <= a;
    layer1_outputs(1596) <= a xor b;
    layer1_outputs(1597) <= not a;
    layer1_outputs(1598) <= b;
    layer1_outputs(1599) <= not a;
    layer1_outputs(1600) <= not (a or b);
    layer1_outputs(1601) <= b;
    layer1_outputs(1602) <= not b or a;
    layer1_outputs(1603) <= not (a xor b);
    layer1_outputs(1604) <= not (a or b);
    layer1_outputs(1605) <= b;
    layer1_outputs(1606) <= not b;
    layer1_outputs(1607) <= a xor b;
    layer1_outputs(1608) <= not b or a;
    layer1_outputs(1609) <= a and b;
    layer1_outputs(1610) <= not (a xor b);
    layer1_outputs(1611) <= not (a xor b);
    layer1_outputs(1612) <= not b or a;
    layer1_outputs(1613) <= not (a xor b);
    layer1_outputs(1614) <= not (a and b);
    layer1_outputs(1615) <= not (a and b);
    layer1_outputs(1616) <= a and not b;
    layer1_outputs(1617) <= not b;
    layer1_outputs(1618) <= b;
    layer1_outputs(1619) <= not (a or b);
    layer1_outputs(1620) <= not b or a;
    layer1_outputs(1621) <= not (a xor b);
    layer1_outputs(1622) <= a and b;
    layer1_outputs(1623) <= not (a and b);
    layer1_outputs(1624) <= a xor b;
    layer1_outputs(1625) <= a;
    layer1_outputs(1626) <= not (a or b);
    layer1_outputs(1627) <= a or b;
    layer1_outputs(1628) <= a and b;
    layer1_outputs(1629) <= not b;
    layer1_outputs(1630) <= a and not b;
    layer1_outputs(1631) <= not (a xor b);
    layer1_outputs(1632) <= not (a and b);
    layer1_outputs(1633) <= a or b;
    layer1_outputs(1634) <= b;
    layer1_outputs(1635) <= a;
    layer1_outputs(1636) <= not (a xor b);
    layer1_outputs(1637) <= not (a or b);
    layer1_outputs(1638) <= a and b;
    layer1_outputs(1639) <= b;
    layer1_outputs(1640) <= b;
    layer1_outputs(1641) <= not a;
    layer1_outputs(1642) <= not b;
    layer1_outputs(1643) <= a or b;
    layer1_outputs(1644) <= not b or a;
    layer1_outputs(1645) <= a;
    layer1_outputs(1646) <= not (a and b);
    layer1_outputs(1647) <= b and not a;
    layer1_outputs(1648) <= a and b;
    layer1_outputs(1649) <= 1'b0;
    layer1_outputs(1650) <= a or b;
    layer1_outputs(1651) <= not (a and b);
    layer1_outputs(1652) <= a or b;
    layer1_outputs(1653) <= not (a or b);
    layer1_outputs(1654) <= a or b;
    layer1_outputs(1655) <= a or b;
    layer1_outputs(1656) <= a;
    layer1_outputs(1657) <= b and not a;
    layer1_outputs(1658) <= 1'b1;
    layer1_outputs(1659) <= not (a and b);
    layer1_outputs(1660) <= b;
    layer1_outputs(1661) <= a xor b;
    layer1_outputs(1662) <= not (a xor b);
    layer1_outputs(1663) <= not (a xor b);
    layer1_outputs(1664) <= not a or b;
    layer1_outputs(1665) <= not a;
    layer1_outputs(1666) <= not (a xor b);
    layer1_outputs(1667) <= 1'b1;
    layer1_outputs(1668) <= not (a and b);
    layer1_outputs(1669) <= not b;
    layer1_outputs(1670) <= not a or b;
    layer1_outputs(1671) <= a xor b;
    layer1_outputs(1672) <= a xor b;
    layer1_outputs(1673) <= not (a or b);
    layer1_outputs(1674) <= b and not a;
    layer1_outputs(1675) <= not a;
    layer1_outputs(1676) <= a or b;
    layer1_outputs(1677) <= b and not a;
    layer1_outputs(1678) <= not (a xor b);
    layer1_outputs(1679) <= b;
    layer1_outputs(1680) <= not (a or b);
    layer1_outputs(1681) <= not b;
    layer1_outputs(1682) <= not (a or b);
    layer1_outputs(1683) <= a;
    layer1_outputs(1684) <= not (a or b);
    layer1_outputs(1685) <= a;
    layer1_outputs(1686) <= not b;
    layer1_outputs(1687) <= a and not b;
    layer1_outputs(1688) <= b;
    layer1_outputs(1689) <= not (a and b);
    layer1_outputs(1690) <= a or b;
    layer1_outputs(1691) <= not (a and b);
    layer1_outputs(1692) <= not (a xor b);
    layer1_outputs(1693) <= not (a or b);
    layer1_outputs(1694) <= a and not b;
    layer1_outputs(1695) <= b and not a;
    layer1_outputs(1696) <= not (a and b);
    layer1_outputs(1697) <= a and not b;
    layer1_outputs(1698) <= not (a or b);
    layer1_outputs(1699) <= b;
    layer1_outputs(1700) <= not b or a;
    layer1_outputs(1701) <= a and b;
    layer1_outputs(1702) <= a and b;
    layer1_outputs(1703) <= a xor b;
    layer1_outputs(1704) <= a;
    layer1_outputs(1705) <= not b or a;
    layer1_outputs(1706) <= not (a xor b);
    layer1_outputs(1707) <= not (a xor b);
    layer1_outputs(1708) <= not a or b;
    layer1_outputs(1709) <= not a;
    layer1_outputs(1710) <= not (a and b);
    layer1_outputs(1711) <= a xor b;
    layer1_outputs(1712) <= b;
    layer1_outputs(1713) <= 1'b0;
    layer1_outputs(1714) <= not b;
    layer1_outputs(1715) <= not b or a;
    layer1_outputs(1716) <= a or b;
    layer1_outputs(1717) <= b;
    layer1_outputs(1718) <= not (a and b);
    layer1_outputs(1719) <= a;
    layer1_outputs(1720) <= not (a or b);
    layer1_outputs(1721) <= not b or a;
    layer1_outputs(1722) <= a or b;
    layer1_outputs(1723) <= b;
    layer1_outputs(1724) <= a xor b;
    layer1_outputs(1725) <= 1'b0;
    layer1_outputs(1726) <= a or b;
    layer1_outputs(1727) <= not a or b;
    layer1_outputs(1728) <= b and not a;
    layer1_outputs(1729) <= a xor b;
    layer1_outputs(1730) <= a and b;
    layer1_outputs(1731) <= not a;
    layer1_outputs(1732) <= not b;
    layer1_outputs(1733) <= a and not b;
    layer1_outputs(1734) <= not b or a;
    layer1_outputs(1735) <= not b;
    layer1_outputs(1736) <= not (a and b);
    layer1_outputs(1737) <= not a;
    layer1_outputs(1738) <= a xor b;
    layer1_outputs(1739) <= a;
    layer1_outputs(1740) <= b;
    layer1_outputs(1741) <= b;
    layer1_outputs(1742) <= a xor b;
    layer1_outputs(1743) <= a and not b;
    layer1_outputs(1744) <= not b;
    layer1_outputs(1745) <= not b;
    layer1_outputs(1746) <= not (a xor b);
    layer1_outputs(1747) <= not a;
    layer1_outputs(1748) <= not b or a;
    layer1_outputs(1749) <= a;
    layer1_outputs(1750) <= a and b;
    layer1_outputs(1751) <= a;
    layer1_outputs(1752) <= not a;
    layer1_outputs(1753) <= b;
    layer1_outputs(1754) <= b and not a;
    layer1_outputs(1755) <= a and b;
    layer1_outputs(1756) <= a or b;
    layer1_outputs(1757) <= b and not a;
    layer1_outputs(1758) <= not a;
    layer1_outputs(1759) <= a;
    layer1_outputs(1760) <= a xor b;
    layer1_outputs(1761) <= not a;
    layer1_outputs(1762) <= not (a xor b);
    layer1_outputs(1763) <= a;
    layer1_outputs(1764) <= not a or b;
    layer1_outputs(1765) <= not b;
    layer1_outputs(1766) <= a;
    layer1_outputs(1767) <= not (a and b);
    layer1_outputs(1768) <= b;
    layer1_outputs(1769) <= b and not a;
    layer1_outputs(1770) <= not (a xor b);
    layer1_outputs(1771) <= b and not a;
    layer1_outputs(1772) <= a;
    layer1_outputs(1773) <= not a;
    layer1_outputs(1774) <= not b;
    layer1_outputs(1775) <= not a;
    layer1_outputs(1776) <= not (a or b);
    layer1_outputs(1777) <= a and not b;
    layer1_outputs(1778) <= a or b;
    layer1_outputs(1779) <= a and b;
    layer1_outputs(1780) <= a and not b;
    layer1_outputs(1781) <= not b or a;
    layer1_outputs(1782) <= b and not a;
    layer1_outputs(1783) <= a xor b;
    layer1_outputs(1784) <= a or b;
    layer1_outputs(1785) <= b and not a;
    layer1_outputs(1786) <= not a or b;
    layer1_outputs(1787) <= not (a and b);
    layer1_outputs(1788) <= not b or a;
    layer1_outputs(1789) <= a and not b;
    layer1_outputs(1790) <= b;
    layer1_outputs(1791) <= not a or b;
    layer1_outputs(1792) <= not (a and b);
    layer1_outputs(1793) <= 1'b1;
    layer1_outputs(1794) <= a and not b;
    layer1_outputs(1795) <= a;
    layer1_outputs(1796) <= b and not a;
    layer1_outputs(1797) <= not b or a;
    layer1_outputs(1798) <= not (a and b);
    layer1_outputs(1799) <= not a or b;
    layer1_outputs(1800) <= 1'b0;
    layer1_outputs(1801) <= not b;
    layer1_outputs(1802) <= b and not a;
    layer1_outputs(1803) <= not (a and b);
    layer1_outputs(1804) <= not a or b;
    layer1_outputs(1805) <= a;
    layer1_outputs(1806) <= not b or a;
    layer1_outputs(1807) <= not a or b;
    layer1_outputs(1808) <= a and b;
    layer1_outputs(1809) <= not b or a;
    layer1_outputs(1810) <= not (a xor b);
    layer1_outputs(1811) <= a xor b;
    layer1_outputs(1812) <= a and not b;
    layer1_outputs(1813) <= a xor b;
    layer1_outputs(1814) <= not (a and b);
    layer1_outputs(1815) <= not (a xor b);
    layer1_outputs(1816) <= b and not a;
    layer1_outputs(1817) <= a or b;
    layer1_outputs(1818) <= not b;
    layer1_outputs(1819) <= a;
    layer1_outputs(1820) <= b;
    layer1_outputs(1821) <= not b or a;
    layer1_outputs(1822) <= not a or b;
    layer1_outputs(1823) <= a and not b;
    layer1_outputs(1824) <= a;
    layer1_outputs(1825) <= not a;
    layer1_outputs(1826) <= not b;
    layer1_outputs(1827) <= not (a and b);
    layer1_outputs(1828) <= not (a xor b);
    layer1_outputs(1829) <= a and b;
    layer1_outputs(1830) <= a or b;
    layer1_outputs(1831) <= not a or b;
    layer1_outputs(1832) <= not b;
    layer1_outputs(1833) <= not (a and b);
    layer1_outputs(1834) <= not b;
    layer1_outputs(1835) <= a and b;
    layer1_outputs(1836) <= not a;
    layer1_outputs(1837) <= not b;
    layer1_outputs(1838) <= not a;
    layer1_outputs(1839) <= not b or a;
    layer1_outputs(1840) <= not a or b;
    layer1_outputs(1841) <= 1'b1;
    layer1_outputs(1842) <= b;
    layer1_outputs(1843) <= a or b;
    layer1_outputs(1844) <= 1'b1;
    layer1_outputs(1845) <= b and not a;
    layer1_outputs(1846) <= b;
    layer1_outputs(1847) <= a and b;
    layer1_outputs(1848) <= not b;
    layer1_outputs(1849) <= a;
    layer1_outputs(1850) <= not (a xor b);
    layer1_outputs(1851) <= not a or b;
    layer1_outputs(1852) <= not a or b;
    layer1_outputs(1853) <= a;
    layer1_outputs(1854) <= a xor b;
    layer1_outputs(1855) <= not b;
    layer1_outputs(1856) <= a or b;
    layer1_outputs(1857) <= b and not a;
    layer1_outputs(1858) <= not a;
    layer1_outputs(1859) <= not (a and b);
    layer1_outputs(1860) <= not a or b;
    layer1_outputs(1861) <= not b or a;
    layer1_outputs(1862) <= not a or b;
    layer1_outputs(1863) <= a and b;
    layer1_outputs(1864) <= not (a or b);
    layer1_outputs(1865) <= not a;
    layer1_outputs(1866) <= not (a xor b);
    layer1_outputs(1867) <= a or b;
    layer1_outputs(1868) <= not b;
    layer1_outputs(1869) <= a or b;
    layer1_outputs(1870) <= not (a xor b);
    layer1_outputs(1871) <= a;
    layer1_outputs(1872) <= b and not a;
    layer1_outputs(1873) <= b;
    layer1_outputs(1874) <= a;
    layer1_outputs(1875) <= not (a or b);
    layer1_outputs(1876) <= not b;
    layer1_outputs(1877) <= not b or a;
    layer1_outputs(1878) <= a and not b;
    layer1_outputs(1879) <= a and not b;
    layer1_outputs(1880) <= not b or a;
    layer1_outputs(1881) <= b;
    layer1_outputs(1882) <= not (a xor b);
    layer1_outputs(1883) <= b;
    layer1_outputs(1884) <= a or b;
    layer1_outputs(1885) <= a;
    layer1_outputs(1886) <= not b or a;
    layer1_outputs(1887) <= not (a or b);
    layer1_outputs(1888) <= a;
    layer1_outputs(1889) <= not (a xor b);
    layer1_outputs(1890) <= not b;
    layer1_outputs(1891) <= b and not a;
    layer1_outputs(1892) <= not (a or b);
    layer1_outputs(1893) <= not b or a;
    layer1_outputs(1894) <= a xor b;
    layer1_outputs(1895) <= not b;
    layer1_outputs(1896) <= a;
    layer1_outputs(1897) <= not (a and b);
    layer1_outputs(1898) <= a;
    layer1_outputs(1899) <= not a;
    layer1_outputs(1900) <= a and b;
    layer1_outputs(1901) <= a;
    layer1_outputs(1902) <= b and not a;
    layer1_outputs(1903) <= not b or a;
    layer1_outputs(1904) <= not (a and b);
    layer1_outputs(1905) <= not b;
    layer1_outputs(1906) <= b;
    layer1_outputs(1907) <= a and b;
    layer1_outputs(1908) <= a xor b;
    layer1_outputs(1909) <= not b;
    layer1_outputs(1910) <= 1'b1;
    layer1_outputs(1911) <= a and not b;
    layer1_outputs(1912) <= not a;
    layer1_outputs(1913) <= not a;
    layer1_outputs(1914) <= a;
    layer1_outputs(1915) <= a;
    layer1_outputs(1916) <= b and not a;
    layer1_outputs(1917) <= not b;
    layer1_outputs(1918) <= a or b;
    layer1_outputs(1919) <= b;
    layer1_outputs(1920) <= not (a xor b);
    layer1_outputs(1921) <= not (a xor b);
    layer1_outputs(1922) <= a and not b;
    layer1_outputs(1923) <= not a;
    layer1_outputs(1924) <= b and not a;
    layer1_outputs(1925) <= not (a and b);
    layer1_outputs(1926) <= a;
    layer1_outputs(1927) <= not (a xor b);
    layer1_outputs(1928) <= not (a or b);
    layer1_outputs(1929) <= not b;
    layer1_outputs(1930) <= not (a and b);
    layer1_outputs(1931) <= not (a and b);
    layer1_outputs(1932) <= a;
    layer1_outputs(1933) <= not b or a;
    layer1_outputs(1934) <= a and not b;
    layer1_outputs(1935) <= a or b;
    layer1_outputs(1936) <= b;
    layer1_outputs(1937) <= a;
    layer1_outputs(1938) <= a and b;
    layer1_outputs(1939) <= a and b;
    layer1_outputs(1940) <= not a or b;
    layer1_outputs(1941) <= not a;
    layer1_outputs(1942) <= not b or a;
    layer1_outputs(1943) <= b and not a;
    layer1_outputs(1944) <= not (a xor b);
    layer1_outputs(1945) <= a or b;
    layer1_outputs(1946) <= not b or a;
    layer1_outputs(1947) <= a and not b;
    layer1_outputs(1948) <= a xor b;
    layer1_outputs(1949) <= b and not a;
    layer1_outputs(1950) <= not (a or b);
    layer1_outputs(1951) <= a and b;
    layer1_outputs(1952) <= b;
    layer1_outputs(1953) <= a xor b;
    layer1_outputs(1954) <= a and b;
    layer1_outputs(1955) <= a and b;
    layer1_outputs(1956) <= not b;
    layer1_outputs(1957) <= b;
    layer1_outputs(1958) <= a;
    layer1_outputs(1959) <= a and b;
    layer1_outputs(1960) <= b and not a;
    layer1_outputs(1961) <= not (a and b);
    layer1_outputs(1962) <= not b or a;
    layer1_outputs(1963) <= not (a and b);
    layer1_outputs(1964) <= not b;
    layer1_outputs(1965) <= a xor b;
    layer1_outputs(1966) <= not (a xor b);
    layer1_outputs(1967) <= a xor b;
    layer1_outputs(1968) <= not b;
    layer1_outputs(1969) <= not b;
    layer1_outputs(1970) <= b;
    layer1_outputs(1971) <= not (a xor b);
    layer1_outputs(1972) <= a;
    layer1_outputs(1973) <= b and not a;
    layer1_outputs(1974) <= not (a xor b);
    layer1_outputs(1975) <= not b;
    layer1_outputs(1976) <= a or b;
    layer1_outputs(1977) <= not (a or b);
    layer1_outputs(1978) <= a and b;
    layer1_outputs(1979) <= not (a xor b);
    layer1_outputs(1980) <= a and not b;
    layer1_outputs(1981) <= not b;
    layer1_outputs(1982) <= a xor b;
    layer1_outputs(1983) <= b;
    layer1_outputs(1984) <= not b or a;
    layer1_outputs(1985) <= not (a xor b);
    layer1_outputs(1986) <= b;
    layer1_outputs(1987) <= a xor b;
    layer1_outputs(1988) <= not b;
    layer1_outputs(1989) <= a xor b;
    layer1_outputs(1990) <= a and not b;
    layer1_outputs(1991) <= b;
    layer1_outputs(1992) <= 1'b1;
    layer1_outputs(1993) <= not b;
    layer1_outputs(1994) <= b;
    layer1_outputs(1995) <= not a or b;
    layer1_outputs(1996) <= a xor b;
    layer1_outputs(1997) <= a or b;
    layer1_outputs(1998) <= not (a xor b);
    layer1_outputs(1999) <= a or b;
    layer1_outputs(2000) <= a and not b;
    layer1_outputs(2001) <= not a;
    layer1_outputs(2002) <= not b or a;
    layer1_outputs(2003) <= not a;
    layer1_outputs(2004) <= a xor b;
    layer1_outputs(2005) <= not b or a;
    layer1_outputs(2006) <= not a;
    layer1_outputs(2007) <= a xor b;
    layer1_outputs(2008) <= not b or a;
    layer1_outputs(2009) <= a and not b;
    layer1_outputs(2010) <= a xor b;
    layer1_outputs(2011) <= a xor b;
    layer1_outputs(2012) <= not a;
    layer1_outputs(2013) <= b;
    layer1_outputs(2014) <= a xor b;
    layer1_outputs(2015) <= a or b;
    layer1_outputs(2016) <= a or b;
    layer1_outputs(2017) <= a;
    layer1_outputs(2018) <= not (a xor b);
    layer1_outputs(2019) <= not b or a;
    layer1_outputs(2020) <= a xor b;
    layer1_outputs(2021) <= not a or b;
    layer1_outputs(2022) <= not b or a;
    layer1_outputs(2023) <= not b;
    layer1_outputs(2024) <= a;
    layer1_outputs(2025) <= a and not b;
    layer1_outputs(2026) <= a and not b;
    layer1_outputs(2027) <= not b;
    layer1_outputs(2028) <= not b;
    layer1_outputs(2029) <= b and not a;
    layer1_outputs(2030) <= not (a xor b);
    layer1_outputs(2031) <= a or b;
    layer1_outputs(2032) <= a xor b;
    layer1_outputs(2033) <= b and not a;
    layer1_outputs(2034) <= not (a or b);
    layer1_outputs(2035) <= not (a and b);
    layer1_outputs(2036) <= not b;
    layer1_outputs(2037) <= a;
    layer1_outputs(2038) <= a xor b;
    layer1_outputs(2039) <= not (a or b);
    layer1_outputs(2040) <= a xor b;
    layer1_outputs(2041) <= a xor b;
    layer1_outputs(2042) <= a;
    layer1_outputs(2043) <= not (a and b);
    layer1_outputs(2044) <= not (a or b);
    layer1_outputs(2045) <= b;
    layer1_outputs(2046) <= a and b;
    layer1_outputs(2047) <= a or b;
    layer1_outputs(2048) <= not (a and b);
    layer1_outputs(2049) <= b;
    layer1_outputs(2050) <= not (a or b);
    layer1_outputs(2051) <= not (a and b);
    layer1_outputs(2052) <= not (a xor b);
    layer1_outputs(2053) <= not b or a;
    layer1_outputs(2054) <= a;
    layer1_outputs(2055) <= not a or b;
    layer1_outputs(2056) <= not b;
    layer1_outputs(2057) <= a xor b;
    layer1_outputs(2058) <= a;
    layer1_outputs(2059) <= a and not b;
    layer1_outputs(2060) <= not a;
    layer1_outputs(2061) <= not a or b;
    layer1_outputs(2062) <= a and b;
    layer1_outputs(2063) <= 1'b0;
    layer1_outputs(2064) <= b and not a;
    layer1_outputs(2065) <= not a;
    layer1_outputs(2066) <= not (a or b);
    layer1_outputs(2067) <= a xor b;
    layer1_outputs(2068) <= b;
    layer1_outputs(2069) <= a and not b;
    layer1_outputs(2070) <= a and b;
    layer1_outputs(2071) <= a and b;
    layer1_outputs(2072) <= not b or a;
    layer1_outputs(2073) <= a or b;
    layer1_outputs(2074) <= not (a xor b);
    layer1_outputs(2075) <= not b;
    layer1_outputs(2076) <= not b;
    layer1_outputs(2077) <= a and not b;
    layer1_outputs(2078) <= a xor b;
    layer1_outputs(2079) <= a and not b;
    layer1_outputs(2080) <= a xor b;
    layer1_outputs(2081) <= not a or b;
    layer1_outputs(2082) <= a and b;
    layer1_outputs(2083) <= b and not a;
    layer1_outputs(2084) <= not a;
    layer1_outputs(2085) <= not (a xor b);
    layer1_outputs(2086) <= a;
    layer1_outputs(2087) <= a or b;
    layer1_outputs(2088) <= a;
    layer1_outputs(2089) <= b;
    layer1_outputs(2090) <= not (a and b);
    layer1_outputs(2091) <= not b;
    layer1_outputs(2092) <= 1'b1;
    layer1_outputs(2093) <= not (a xor b);
    layer1_outputs(2094) <= not (a or b);
    layer1_outputs(2095) <= a xor b;
    layer1_outputs(2096) <= not a or b;
    layer1_outputs(2097) <= not (a or b);
    layer1_outputs(2098) <= not b or a;
    layer1_outputs(2099) <= not b;
    layer1_outputs(2100) <= not b or a;
    layer1_outputs(2101) <= not (a xor b);
    layer1_outputs(2102) <= b and not a;
    layer1_outputs(2103) <= not b;
    layer1_outputs(2104) <= not (a xor b);
    layer1_outputs(2105) <= 1'b0;
    layer1_outputs(2106) <= not (a or b);
    layer1_outputs(2107) <= a;
    layer1_outputs(2108) <= a xor b;
    layer1_outputs(2109) <= a and b;
    layer1_outputs(2110) <= a xor b;
    layer1_outputs(2111) <= not b or a;
    layer1_outputs(2112) <= a xor b;
    layer1_outputs(2113) <= a xor b;
    layer1_outputs(2114) <= not b;
    layer1_outputs(2115) <= a xor b;
    layer1_outputs(2116) <= a;
    layer1_outputs(2117) <= a and not b;
    layer1_outputs(2118) <= a xor b;
    layer1_outputs(2119) <= a xor b;
    layer1_outputs(2120) <= not (a and b);
    layer1_outputs(2121) <= not b or a;
    layer1_outputs(2122) <= not a or b;
    layer1_outputs(2123) <= a and b;
    layer1_outputs(2124) <= 1'b1;
    layer1_outputs(2125) <= not a or b;
    layer1_outputs(2126) <= not (a or b);
    layer1_outputs(2127) <= not a;
    layer1_outputs(2128) <= not b;
    layer1_outputs(2129) <= not (a and b);
    layer1_outputs(2130) <= a or b;
    layer1_outputs(2131) <= not a;
    layer1_outputs(2132) <= a;
    layer1_outputs(2133) <= not a or b;
    layer1_outputs(2134) <= 1'b1;
    layer1_outputs(2135) <= not (a xor b);
    layer1_outputs(2136) <= a and not b;
    layer1_outputs(2137) <= a or b;
    layer1_outputs(2138) <= a or b;
    layer1_outputs(2139) <= a or b;
    layer1_outputs(2140) <= not (a or b);
    layer1_outputs(2141) <= not a or b;
    layer1_outputs(2142) <= a and b;
    layer1_outputs(2143) <= not (a or b);
    layer1_outputs(2144) <= a and not b;
    layer1_outputs(2145) <= a xor b;
    layer1_outputs(2146) <= a xor b;
    layer1_outputs(2147) <= not (a xor b);
    layer1_outputs(2148) <= not a;
    layer1_outputs(2149) <= a xor b;
    layer1_outputs(2150) <= b;
    layer1_outputs(2151) <= a or b;
    layer1_outputs(2152) <= not (a or b);
    layer1_outputs(2153) <= not (a and b);
    layer1_outputs(2154) <= not a;
    layer1_outputs(2155) <= a or b;
    layer1_outputs(2156) <= not (a or b);
    layer1_outputs(2157) <= b and not a;
    layer1_outputs(2158) <= a and not b;
    layer1_outputs(2159) <= a;
    layer1_outputs(2160) <= a xor b;
    layer1_outputs(2161) <= b and not a;
    layer1_outputs(2162) <= not b or a;
    layer1_outputs(2163) <= b and not a;
    layer1_outputs(2164) <= not b or a;
    layer1_outputs(2165) <= not (a and b);
    layer1_outputs(2166) <= a or b;
    layer1_outputs(2167) <= b;
    layer1_outputs(2168) <= a;
    layer1_outputs(2169) <= a and b;
    layer1_outputs(2170) <= a or b;
    layer1_outputs(2171) <= not a;
    layer1_outputs(2172) <= b;
    layer1_outputs(2173) <= not (a and b);
    layer1_outputs(2174) <= a xor b;
    layer1_outputs(2175) <= a xor b;
    layer1_outputs(2176) <= not a;
    layer1_outputs(2177) <= not (a and b);
    layer1_outputs(2178) <= a;
    layer1_outputs(2179) <= a;
    layer1_outputs(2180) <= not (a and b);
    layer1_outputs(2181) <= a xor b;
    layer1_outputs(2182) <= a and b;
    layer1_outputs(2183) <= not (a or b);
    layer1_outputs(2184) <= not a;
    layer1_outputs(2185) <= 1'b0;
    layer1_outputs(2186) <= not (a xor b);
    layer1_outputs(2187) <= a;
    layer1_outputs(2188) <= not (a and b);
    layer1_outputs(2189) <= not a;
    layer1_outputs(2190) <= not a or b;
    layer1_outputs(2191) <= not (a xor b);
    layer1_outputs(2192) <= not b;
    layer1_outputs(2193) <= a;
    layer1_outputs(2194) <= not (a xor b);
    layer1_outputs(2195) <= not (a and b);
    layer1_outputs(2196) <= a xor b;
    layer1_outputs(2197) <= 1'b0;
    layer1_outputs(2198) <= not a;
    layer1_outputs(2199) <= 1'b1;
    layer1_outputs(2200) <= not a;
    layer1_outputs(2201) <= not b;
    layer1_outputs(2202) <= not a or b;
    layer1_outputs(2203) <= a and not b;
    layer1_outputs(2204) <= a;
    layer1_outputs(2205) <= not b;
    layer1_outputs(2206) <= not b;
    layer1_outputs(2207) <= not b;
    layer1_outputs(2208) <= not a;
    layer1_outputs(2209) <= not a;
    layer1_outputs(2210) <= a;
    layer1_outputs(2211) <= a and not b;
    layer1_outputs(2212) <= a and not b;
    layer1_outputs(2213) <= not b;
    layer1_outputs(2214) <= a and b;
    layer1_outputs(2215) <= not (a and b);
    layer1_outputs(2216) <= b;
    layer1_outputs(2217) <= not a;
    layer1_outputs(2218) <= a and b;
    layer1_outputs(2219) <= not b or a;
    layer1_outputs(2220) <= a;
    layer1_outputs(2221) <= not (a xor b);
    layer1_outputs(2222) <= a;
    layer1_outputs(2223) <= a;
    layer1_outputs(2224) <= a;
    layer1_outputs(2225) <= a;
    layer1_outputs(2226) <= not b or a;
    layer1_outputs(2227) <= a;
    layer1_outputs(2228) <= a;
    layer1_outputs(2229) <= a and b;
    layer1_outputs(2230) <= not (a and b);
    layer1_outputs(2231) <= 1'b0;
    layer1_outputs(2232) <= 1'b0;
    layer1_outputs(2233) <= b and not a;
    layer1_outputs(2234) <= not (a xor b);
    layer1_outputs(2235) <= not (a and b);
    layer1_outputs(2236) <= a and b;
    layer1_outputs(2237) <= a or b;
    layer1_outputs(2238) <= a;
    layer1_outputs(2239) <= b and not a;
    layer1_outputs(2240) <= b;
    layer1_outputs(2241) <= not (a or b);
    layer1_outputs(2242) <= a;
    layer1_outputs(2243) <= not a;
    layer1_outputs(2244) <= not (a xor b);
    layer1_outputs(2245) <= not b or a;
    layer1_outputs(2246) <= a;
    layer1_outputs(2247) <= a and b;
    layer1_outputs(2248) <= not a;
    layer1_outputs(2249) <= a and not b;
    layer1_outputs(2250) <= b;
    layer1_outputs(2251) <= not (a xor b);
    layer1_outputs(2252) <= not b or a;
    layer1_outputs(2253) <= a and not b;
    layer1_outputs(2254) <= a or b;
    layer1_outputs(2255) <= b;
    layer1_outputs(2256) <= a xor b;
    layer1_outputs(2257) <= a and b;
    layer1_outputs(2258) <= not a;
    layer1_outputs(2259) <= not (a xor b);
    layer1_outputs(2260) <= not a;
    layer1_outputs(2261) <= a xor b;
    layer1_outputs(2262) <= a xor b;
    layer1_outputs(2263) <= a or b;
    layer1_outputs(2264) <= b and not a;
    layer1_outputs(2265) <= a;
    layer1_outputs(2266) <= b;
    layer1_outputs(2267) <= a and not b;
    layer1_outputs(2268) <= not b;
    layer1_outputs(2269) <= not (a and b);
    layer1_outputs(2270) <= a and b;
    layer1_outputs(2271) <= not a or b;
    layer1_outputs(2272) <= b;
    layer1_outputs(2273) <= a or b;
    layer1_outputs(2274) <= a and not b;
    layer1_outputs(2275) <= b and not a;
    layer1_outputs(2276) <= not b;
    layer1_outputs(2277) <= not (a and b);
    layer1_outputs(2278) <= b;
    layer1_outputs(2279) <= b and not a;
    layer1_outputs(2280) <= b;
    layer1_outputs(2281) <= b and not a;
    layer1_outputs(2282) <= a xor b;
    layer1_outputs(2283) <= not (a and b);
    layer1_outputs(2284) <= a and not b;
    layer1_outputs(2285) <= a xor b;
    layer1_outputs(2286) <= not a;
    layer1_outputs(2287) <= b;
    layer1_outputs(2288) <= not b;
    layer1_outputs(2289) <= not a;
    layer1_outputs(2290) <= a;
    layer1_outputs(2291) <= not a or b;
    layer1_outputs(2292) <= not (a or b);
    layer1_outputs(2293) <= a or b;
    layer1_outputs(2294) <= a xor b;
    layer1_outputs(2295) <= a and not b;
    layer1_outputs(2296) <= b;
    layer1_outputs(2297) <= not b;
    layer1_outputs(2298) <= not (a xor b);
    layer1_outputs(2299) <= not (a xor b);
    layer1_outputs(2300) <= a and not b;
    layer1_outputs(2301) <= not a or b;
    layer1_outputs(2302) <= a;
    layer1_outputs(2303) <= a and not b;
    layer1_outputs(2304) <= a or b;
    layer1_outputs(2305) <= a and b;
    layer1_outputs(2306) <= a xor b;
    layer1_outputs(2307) <= not (a xor b);
    layer1_outputs(2308) <= a xor b;
    layer1_outputs(2309) <= 1'b0;
    layer1_outputs(2310) <= a or b;
    layer1_outputs(2311) <= b;
    layer1_outputs(2312) <= not (a xor b);
    layer1_outputs(2313) <= a and not b;
    layer1_outputs(2314) <= not a;
    layer1_outputs(2315) <= not (a xor b);
    layer1_outputs(2316) <= not a;
    layer1_outputs(2317) <= b;
    layer1_outputs(2318) <= b and not a;
    layer1_outputs(2319) <= b;
    layer1_outputs(2320) <= not b or a;
    layer1_outputs(2321) <= a and b;
    layer1_outputs(2322) <= not a;
    layer1_outputs(2323) <= not (a or b);
    layer1_outputs(2324) <= a or b;
    layer1_outputs(2325) <= a and not b;
    layer1_outputs(2326) <= not (a or b);
    layer1_outputs(2327) <= b;
    layer1_outputs(2328) <= a or b;
    layer1_outputs(2329) <= a xor b;
    layer1_outputs(2330) <= not b;
    layer1_outputs(2331) <= b;
    layer1_outputs(2332) <= a and b;
    layer1_outputs(2333) <= a;
    layer1_outputs(2334) <= a and not b;
    layer1_outputs(2335) <= not a or b;
    layer1_outputs(2336) <= a;
    layer1_outputs(2337) <= not b;
    layer1_outputs(2338) <= b;
    layer1_outputs(2339) <= not b or a;
    layer1_outputs(2340) <= a or b;
    layer1_outputs(2341) <= a xor b;
    layer1_outputs(2342) <= not b or a;
    layer1_outputs(2343) <= 1'b1;
    layer1_outputs(2344) <= a;
    layer1_outputs(2345) <= a and not b;
    layer1_outputs(2346) <= not (a xor b);
    layer1_outputs(2347) <= not (a and b);
    layer1_outputs(2348) <= a;
    layer1_outputs(2349) <= not (a and b);
    layer1_outputs(2350) <= not (a xor b);
    layer1_outputs(2351) <= not (a or b);
    layer1_outputs(2352) <= b and not a;
    layer1_outputs(2353) <= b and not a;
    layer1_outputs(2354) <= not b or a;
    layer1_outputs(2355) <= not (a and b);
    layer1_outputs(2356) <= not (a xor b);
    layer1_outputs(2357) <= b and not a;
    layer1_outputs(2358) <= a and not b;
    layer1_outputs(2359) <= a and not b;
    layer1_outputs(2360) <= not b or a;
    layer1_outputs(2361) <= not a;
    layer1_outputs(2362) <= a;
    layer1_outputs(2363) <= not (a and b);
    layer1_outputs(2364) <= not a or b;
    layer1_outputs(2365) <= 1'b0;
    layer1_outputs(2366) <= not b;
    layer1_outputs(2367) <= a or b;
    layer1_outputs(2368) <= not b;
    layer1_outputs(2369) <= not (a and b);
    layer1_outputs(2370) <= a and b;
    layer1_outputs(2371) <= not (a or b);
    layer1_outputs(2372) <= not a;
    layer1_outputs(2373) <= b and not a;
    layer1_outputs(2374) <= not a;
    layer1_outputs(2375) <= b and not a;
    layer1_outputs(2376) <= not b;
    layer1_outputs(2377) <= not (a xor b);
    layer1_outputs(2378) <= not a;
    layer1_outputs(2379) <= not a;
    layer1_outputs(2380) <= a;
    layer1_outputs(2381) <= not (a xor b);
    layer1_outputs(2382) <= not (a or b);
    layer1_outputs(2383) <= not b or a;
    layer1_outputs(2384) <= b;
    layer1_outputs(2385) <= a or b;
    layer1_outputs(2386) <= not (a or b);
    layer1_outputs(2387) <= a and not b;
    layer1_outputs(2388) <= not a;
    layer1_outputs(2389) <= b;
    layer1_outputs(2390) <= a or b;
    layer1_outputs(2391) <= not a;
    layer1_outputs(2392) <= a;
    layer1_outputs(2393) <= a xor b;
    layer1_outputs(2394) <= b;
    layer1_outputs(2395) <= not a or b;
    layer1_outputs(2396) <= not a;
    layer1_outputs(2397) <= a;
    layer1_outputs(2398) <= not (a or b);
    layer1_outputs(2399) <= a xor b;
    layer1_outputs(2400) <= not (a and b);
    layer1_outputs(2401) <= not a or b;
    layer1_outputs(2402) <= a;
    layer1_outputs(2403) <= a xor b;
    layer1_outputs(2404) <= not b;
    layer1_outputs(2405) <= not (a xor b);
    layer1_outputs(2406) <= 1'b0;
    layer1_outputs(2407) <= not (a xor b);
    layer1_outputs(2408) <= 1'b1;
    layer1_outputs(2409) <= not a;
    layer1_outputs(2410) <= a xor b;
    layer1_outputs(2411) <= a and not b;
    layer1_outputs(2412) <= a xor b;
    layer1_outputs(2413) <= b;
    layer1_outputs(2414) <= a and not b;
    layer1_outputs(2415) <= a and b;
    layer1_outputs(2416) <= not (a or b);
    layer1_outputs(2417) <= not a or b;
    layer1_outputs(2418) <= a;
    layer1_outputs(2419) <= not a;
    layer1_outputs(2420) <= not a;
    layer1_outputs(2421) <= not b or a;
    layer1_outputs(2422) <= a;
    layer1_outputs(2423) <= not b;
    layer1_outputs(2424) <= not b;
    layer1_outputs(2425) <= not (a and b);
    layer1_outputs(2426) <= a;
    layer1_outputs(2427) <= not (a and b);
    layer1_outputs(2428) <= not b;
    layer1_outputs(2429) <= a xor b;
    layer1_outputs(2430) <= not (a xor b);
    layer1_outputs(2431) <= not (a or b);
    layer1_outputs(2432) <= not (a xor b);
    layer1_outputs(2433) <= b and not a;
    layer1_outputs(2434) <= not (a xor b);
    layer1_outputs(2435) <= 1'b1;
    layer1_outputs(2436) <= not (a xor b);
    layer1_outputs(2437) <= 1'b0;
    layer1_outputs(2438) <= a xor b;
    layer1_outputs(2439) <= b;
    layer1_outputs(2440) <= b and not a;
    layer1_outputs(2441) <= a xor b;
    layer1_outputs(2442) <= a xor b;
    layer1_outputs(2443) <= not a;
    layer1_outputs(2444) <= not (a and b);
    layer1_outputs(2445) <= a or b;
    layer1_outputs(2446) <= b;
    layer1_outputs(2447) <= not a;
    layer1_outputs(2448) <= not a;
    layer1_outputs(2449) <= b and not a;
    layer1_outputs(2450) <= not (a and b);
    layer1_outputs(2451) <= not b;
    layer1_outputs(2452) <= b and not a;
    layer1_outputs(2453) <= not b;
    layer1_outputs(2454) <= not (a and b);
    layer1_outputs(2455) <= a and not b;
    layer1_outputs(2456) <= not (a or b);
    layer1_outputs(2457) <= 1'b1;
    layer1_outputs(2458) <= a and not b;
    layer1_outputs(2459) <= not b;
    layer1_outputs(2460) <= a and not b;
    layer1_outputs(2461) <= a xor b;
    layer1_outputs(2462) <= b and not a;
    layer1_outputs(2463) <= not b or a;
    layer1_outputs(2464) <= not a or b;
    layer1_outputs(2465) <= not a or b;
    layer1_outputs(2466) <= b and not a;
    layer1_outputs(2467) <= a;
    layer1_outputs(2468) <= b;
    layer1_outputs(2469) <= a;
    layer1_outputs(2470) <= not (a or b);
    layer1_outputs(2471) <= a;
    layer1_outputs(2472) <= a or b;
    layer1_outputs(2473) <= a;
    layer1_outputs(2474) <= not a or b;
    layer1_outputs(2475) <= b and not a;
    layer1_outputs(2476) <= a xor b;
    layer1_outputs(2477) <= not (a or b);
    layer1_outputs(2478) <= a xor b;
    layer1_outputs(2479) <= not a or b;
    layer1_outputs(2480) <= not (a and b);
    layer1_outputs(2481) <= not (a or b);
    layer1_outputs(2482) <= not (a xor b);
    layer1_outputs(2483) <= a and not b;
    layer1_outputs(2484) <= not a;
    layer1_outputs(2485) <= not (a and b);
    layer1_outputs(2486) <= a or b;
    layer1_outputs(2487) <= not b or a;
    layer1_outputs(2488) <= not b or a;
    layer1_outputs(2489) <= b;
    layer1_outputs(2490) <= not a;
    layer1_outputs(2491) <= a;
    layer1_outputs(2492) <= not a;
    layer1_outputs(2493) <= not b;
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= not b or a;
    layer1_outputs(2496) <= a xor b;
    layer1_outputs(2497) <= not a or b;
    layer1_outputs(2498) <= not b or a;
    layer1_outputs(2499) <= not a;
    layer1_outputs(2500) <= not b or a;
    layer1_outputs(2501) <= b;
    layer1_outputs(2502) <= not b;
    layer1_outputs(2503) <= a;
    layer1_outputs(2504) <= a;
    layer1_outputs(2505) <= a and b;
    layer1_outputs(2506) <= not b or a;
    layer1_outputs(2507) <= not (a and b);
    layer1_outputs(2508) <= not a or b;
    layer1_outputs(2509) <= a and not b;
    layer1_outputs(2510) <= a and not b;
    layer1_outputs(2511) <= not (a xor b);
    layer1_outputs(2512) <= b;
    layer1_outputs(2513) <= 1'b1;
    layer1_outputs(2514) <= b and not a;
    layer1_outputs(2515) <= b and not a;
    layer1_outputs(2516) <= a and b;
    layer1_outputs(2517) <= a and b;
    layer1_outputs(2518) <= a and b;
    layer1_outputs(2519) <= not (a or b);
    layer1_outputs(2520) <= a and not b;
    layer1_outputs(2521) <= a;
    layer1_outputs(2522) <= not b;
    layer1_outputs(2523) <= b and not a;
    layer1_outputs(2524) <= b and not a;
    layer1_outputs(2525) <= not a;
    layer1_outputs(2526) <= b;
    layer1_outputs(2527) <= not a;
    layer1_outputs(2528) <= not a;
    layer1_outputs(2529) <= not a;
    layer1_outputs(2530) <= a;
    layer1_outputs(2531) <= a;
    layer1_outputs(2532) <= b;
    layer1_outputs(2533) <= a xor b;
    layer1_outputs(2534) <= a;
    layer1_outputs(2535) <= a;
    layer1_outputs(2536) <= 1'b1;
    layer1_outputs(2537) <= not b;
    layer1_outputs(2538) <= not b or a;
    layer1_outputs(2539) <= not (a xor b);
    layer1_outputs(2540) <= a or b;
    layer1_outputs(2541) <= a or b;
    layer1_outputs(2542) <= b;
    layer1_outputs(2543) <= b;
    layer1_outputs(2544) <= not a;
    layer1_outputs(2545) <= not a;
    layer1_outputs(2546) <= not b;
    layer1_outputs(2547) <= not a or b;
    layer1_outputs(2548) <= not (a or b);
    layer1_outputs(2549) <= not (a and b);
    layer1_outputs(2550) <= b and not a;
    layer1_outputs(2551) <= not (a or b);
    layer1_outputs(2552) <= not a;
    layer1_outputs(2553) <= not (a xor b);
    layer1_outputs(2554) <= not a or b;
    layer1_outputs(2555) <= 1'b0;
    layer1_outputs(2556) <= not b or a;
    layer1_outputs(2557) <= not b;
    layer1_outputs(2558) <= not (a and b);
    layer1_outputs(2559) <= a or b;
    layer1_outputs(2560) <= b and not a;
    layer1_outputs(2561) <= not (a or b);
    layer1_outputs(2562) <= not a;
    layer1_outputs(2563) <= a;
    layer1_outputs(2564) <= a xor b;
    layer1_outputs(2565) <= not a or b;
    layer1_outputs(2566) <= not b;
    layer1_outputs(2567) <= not b;
    layer1_outputs(2568) <= not (a or b);
    layer1_outputs(2569) <= b and not a;
    layer1_outputs(2570) <= not (a xor b);
    layer1_outputs(2571) <= a or b;
    layer1_outputs(2572) <= not (a and b);
    layer1_outputs(2573) <= b;
    layer1_outputs(2574) <= a;
    layer1_outputs(2575) <= not (a xor b);
    layer1_outputs(2576) <= not (a and b);
    layer1_outputs(2577) <= not b or a;
    layer1_outputs(2578) <= not (a xor b);
    layer1_outputs(2579) <= not b or a;
    layer1_outputs(2580) <= not (a xor b);
    layer1_outputs(2581) <= not a or b;
    layer1_outputs(2582) <= not (a xor b);
    layer1_outputs(2583) <= not a or b;
    layer1_outputs(2584) <= not (a xor b);
    layer1_outputs(2585) <= not b;
    layer1_outputs(2586) <= b;
    layer1_outputs(2587) <= not b or a;
    layer1_outputs(2588) <= not a or b;
    layer1_outputs(2589) <= not a or b;
    layer1_outputs(2590) <= not a;
    layer1_outputs(2591) <= not b or a;
    layer1_outputs(2592) <= a xor b;
    layer1_outputs(2593) <= a and not b;
    layer1_outputs(2594) <= not a or b;
    layer1_outputs(2595) <= b and not a;
    layer1_outputs(2596) <= a or b;
    layer1_outputs(2597) <= a and b;
    layer1_outputs(2598) <= not (a xor b);
    layer1_outputs(2599) <= a xor b;
    layer1_outputs(2600) <= not b;
    layer1_outputs(2601) <= b;
    layer1_outputs(2602) <= b and not a;
    layer1_outputs(2603) <= not a or b;
    layer1_outputs(2604) <= not b;
    layer1_outputs(2605) <= not (a or b);
    layer1_outputs(2606) <= b;
    layer1_outputs(2607) <= b and not a;
    layer1_outputs(2608) <= b and not a;
    layer1_outputs(2609) <= not b;
    layer1_outputs(2610) <= not b or a;
    layer1_outputs(2611) <= a and b;
    layer1_outputs(2612) <= b;
    layer1_outputs(2613) <= not (a or b);
    layer1_outputs(2614) <= not b;
    layer1_outputs(2615) <= b;
    layer1_outputs(2616) <= not b or a;
    layer1_outputs(2617) <= not b or a;
    layer1_outputs(2618) <= b;
    layer1_outputs(2619) <= a;
    layer1_outputs(2620) <= not a;
    layer1_outputs(2621) <= b;
    layer1_outputs(2622) <= a and not b;
    layer1_outputs(2623) <= not (a or b);
    layer1_outputs(2624) <= not a or b;
    layer1_outputs(2625) <= not (a and b);
    layer1_outputs(2626) <= not b;
    layer1_outputs(2627) <= a xor b;
    layer1_outputs(2628) <= not (a or b);
    layer1_outputs(2629) <= not b;
    layer1_outputs(2630) <= not (a xor b);
    layer1_outputs(2631) <= a and b;
    layer1_outputs(2632) <= not (a and b);
    layer1_outputs(2633) <= b and not a;
    layer1_outputs(2634) <= not a or b;
    layer1_outputs(2635) <= a and b;
    layer1_outputs(2636) <= not b;
    layer1_outputs(2637) <= b;
    layer1_outputs(2638) <= b and not a;
    layer1_outputs(2639) <= not (a and b);
    layer1_outputs(2640) <= not (a and b);
    layer1_outputs(2641) <= not b;
    layer1_outputs(2642) <= not (a xor b);
    layer1_outputs(2643) <= not b;
    layer1_outputs(2644) <= not a;
    layer1_outputs(2645) <= b and not a;
    layer1_outputs(2646) <= not a;
    layer1_outputs(2647) <= b and not a;
    layer1_outputs(2648) <= a;
    layer1_outputs(2649) <= not a or b;
    layer1_outputs(2650) <= a or b;
    layer1_outputs(2651) <= not (a and b);
    layer1_outputs(2652) <= a;
    layer1_outputs(2653) <= not a or b;
    layer1_outputs(2654) <= not (a and b);
    layer1_outputs(2655) <= b;
    layer1_outputs(2656) <= not (a xor b);
    layer1_outputs(2657) <= b and not a;
    layer1_outputs(2658) <= 1'b1;
    layer1_outputs(2659) <= not (a and b);
    layer1_outputs(2660) <= not a or b;
    layer1_outputs(2661) <= not b;
    layer1_outputs(2662) <= b and not a;
    layer1_outputs(2663) <= a xor b;
    layer1_outputs(2664) <= not (a xor b);
    layer1_outputs(2665) <= b;
    layer1_outputs(2666) <= not (a and b);
    layer1_outputs(2667) <= not b or a;
    layer1_outputs(2668) <= b and not a;
    layer1_outputs(2669) <= not b;
    layer1_outputs(2670) <= a xor b;
    layer1_outputs(2671) <= not (a and b);
    layer1_outputs(2672) <= a or b;
    layer1_outputs(2673) <= b;
    layer1_outputs(2674) <= not a;
    layer1_outputs(2675) <= not (a xor b);
    layer1_outputs(2676) <= not (a and b);
    layer1_outputs(2677) <= not (a and b);
    layer1_outputs(2678) <= a or b;
    layer1_outputs(2679) <= not a or b;
    layer1_outputs(2680) <= b;
    layer1_outputs(2681) <= a xor b;
    layer1_outputs(2682) <= not b or a;
    layer1_outputs(2683) <= not (a xor b);
    layer1_outputs(2684) <= a or b;
    layer1_outputs(2685) <= not b;
    layer1_outputs(2686) <= not a or b;
    layer1_outputs(2687) <= a xor b;
    layer1_outputs(2688) <= not b or a;
    layer1_outputs(2689) <= not b;
    layer1_outputs(2690) <= not b or a;
    layer1_outputs(2691) <= not a;
    layer1_outputs(2692) <= not b;
    layer1_outputs(2693) <= a;
    layer1_outputs(2694) <= not b or a;
    layer1_outputs(2695) <= not (a xor b);
    layer1_outputs(2696) <= b;
    layer1_outputs(2697) <= a and b;
    layer1_outputs(2698) <= not a;
    layer1_outputs(2699) <= not a or b;
    layer1_outputs(2700) <= not b;
    layer1_outputs(2701) <= not b;
    layer1_outputs(2702) <= a;
    layer1_outputs(2703) <= a;
    layer1_outputs(2704) <= a and not b;
    layer1_outputs(2705) <= not a;
    layer1_outputs(2706) <= b and not a;
    layer1_outputs(2707) <= not (a and b);
    layer1_outputs(2708) <= not (a or b);
    layer1_outputs(2709) <= a xor b;
    layer1_outputs(2710) <= not (a xor b);
    layer1_outputs(2711) <= b;
    layer1_outputs(2712) <= not a;
    layer1_outputs(2713) <= a;
    layer1_outputs(2714) <= a or b;
    layer1_outputs(2715) <= not (a and b);
    layer1_outputs(2716) <= not b;
    layer1_outputs(2717) <= not a or b;
    layer1_outputs(2718) <= not (a and b);
    layer1_outputs(2719) <= not a;
    layer1_outputs(2720) <= not (a and b);
    layer1_outputs(2721) <= not (a and b);
    layer1_outputs(2722) <= not (a or b);
    layer1_outputs(2723) <= a and b;
    layer1_outputs(2724) <= a;
    layer1_outputs(2725) <= b;
    layer1_outputs(2726) <= b;
    layer1_outputs(2727) <= not (a or b);
    layer1_outputs(2728) <= a and not b;
    layer1_outputs(2729) <= not b;
    layer1_outputs(2730) <= a and b;
    layer1_outputs(2731) <= a;
    layer1_outputs(2732) <= a;
    layer1_outputs(2733) <= not b;
    layer1_outputs(2734) <= a or b;
    layer1_outputs(2735) <= a and b;
    layer1_outputs(2736) <= not a or b;
    layer1_outputs(2737) <= not (a and b);
    layer1_outputs(2738) <= b;
    layer1_outputs(2739) <= a and not b;
    layer1_outputs(2740) <= not (a or b);
    layer1_outputs(2741) <= a xor b;
    layer1_outputs(2742) <= a xor b;
    layer1_outputs(2743) <= not (a or b);
    layer1_outputs(2744) <= not a;
    layer1_outputs(2745) <= not a;
    layer1_outputs(2746) <= not a;
    layer1_outputs(2747) <= a;
    layer1_outputs(2748) <= not b;
    layer1_outputs(2749) <= a and not b;
    layer1_outputs(2750) <= not a or b;
    layer1_outputs(2751) <= a and b;
    layer1_outputs(2752) <= a;
    layer1_outputs(2753) <= a xor b;
    layer1_outputs(2754) <= a;
    layer1_outputs(2755) <= not (a and b);
    layer1_outputs(2756) <= b;
    layer1_outputs(2757) <= b and not a;
    layer1_outputs(2758) <= 1'b1;
    layer1_outputs(2759) <= not b;
    layer1_outputs(2760) <= a;
    layer1_outputs(2761) <= not (a or b);
    layer1_outputs(2762) <= not a;
    layer1_outputs(2763) <= a;
    layer1_outputs(2764) <= not (a xor b);
    layer1_outputs(2765) <= b;
    layer1_outputs(2766) <= a or b;
    layer1_outputs(2767) <= not b;
    layer1_outputs(2768) <= b and not a;
    layer1_outputs(2769) <= not b;
    layer1_outputs(2770) <= not a;
    layer1_outputs(2771) <= a;
    layer1_outputs(2772) <= b and not a;
    layer1_outputs(2773) <= a xor b;
    layer1_outputs(2774) <= a;
    layer1_outputs(2775) <= not (a or b);
    layer1_outputs(2776) <= not b;
    layer1_outputs(2777) <= b;
    layer1_outputs(2778) <= b and not a;
    layer1_outputs(2779) <= not a;
    layer1_outputs(2780) <= a;
    layer1_outputs(2781) <= not a or b;
    layer1_outputs(2782) <= a and not b;
    layer1_outputs(2783) <= a;
    layer1_outputs(2784) <= not b;
    layer1_outputs(2785) <= a xor b;
    layer1_outputs(2786) <= not b or a;
    layer1_outputs(2787) <= not b;
    layer1_outputs(2788) <= a xor b;
    layer1_outputs(2789) <= not b;
    layer1_outputs(2790) <= a;
    layer1_outputs(2791) <= b;
    layer1_outputs(2792) <= a and not b;
    layer1_outputs(2793) <= a;
    layer1_outputs(2794) <= a and b;
    layer1_outputs(2795) <= not a or b;
    layer1_outputs(2796) <= not b;
    layer1_outputs(2797) <= a and not b;
    layer1_outputs(2798) <= not a;
    layer1_outputs(2799) <= not (a xor b);
    layer1_outputs(2800) <= not (a or b);
    layer1_outputs(2801) <= not (a and b);
    layer1_outputs(2802) <= b;
    layer1_outputs(2803) <= a and not b;
    layer1_outputs(2804) <= a or b;
    layer1_outputs(2805) <= 1'b1;
    layer1_outputs(2806) <= not a or b;
    layer1_outputs(2807) <= b and not a;
    layer1_outputs(2808) <= b and not a;
    layer1_outputs(2809) <= b;
    layer1_outputs(2810) <= 1'b0;
    layer1_outputs(2811) <= not (a and b);
    layer1_outputs(2812) <= a and not b;
    layer1_outputs(2813) <= a;
    layer1_outputs(2814) <= not b;
    layer1_outputs(2815) <= not a;
    layer1_outputs(2816) <= not a;
    layer1_outputs(2817) <= not (a and b);
    layer1_outputs(2818) <= b and not a;
    layer1_outputs(2819) <= a or b;
    layer1_outputs(2820) <= a;
    layer1_outputs(2821) <= a or b;
    layer1_outputs(2822) <= a;
    layer1_outputs(2823) <= 1'b1;
    layer1_outputs(2824) <= a xor b;
    layer1_outputs(2825) <= not a;
    layer1_outputs(2826) <= a xor b;
    layer1_outputs(2827) <= not b or a;
    layer1_outputs(2828) <= a;
    layer1_outputs(2829) <= a;
    layer1_outputs(2830) <= a and not b;
    layer1_outputs(2831) <= not b or a;
    layer1_outputs(2832) <= not a or b;
    layer1_outputs(2833) <= not (a or b);
    layer1_outputs(2834) <= not (a or b);
    layer1_outputs(2835) <= not b or a;
    layer1_outputs(2836) <= not b;
    layer1_outputs(2837) <= a;
    layer1_outputs(2838) <= a or b;
    layer1_outputs(2839) <= not a;
    layer1_outputs(2840) <= a;
    layer1_outputs(2841) <= not (a xor b);
    layer1_outputs(2842) <= b;
    layer1_outputs(2843) <= not b or a;
    layer1_outputs(2844) <= not (a and b);
    layer1_outputs(2845) <= not b;
    layer1_outputs(2846) <= b and not a;
    layer1_outputs(2847) <= not (a xor b);
    layer1_outputs(2848) <= not (a xor b);
    layer1_outputs(2849) <= not a;
    layer1_outputs(2850) <= not a;
    layer1_outputs(2851) <= b and not a;
    layer1_outputs(2852) <= not b;
    layer1_outputs(2853) <= a and b;
    layer1_outputs(2854) <= not b;
    layer1_outputs(2855) <= b;
    layer1_outputs(2856) <= 1'b1;
    layer1_outputs(2857) <= not b or a;
    layer1_outputs(2858) <= b;
    layer1_outputs(2859) <= a;
    layer1_outputs(2860) <= not (a and b);
    layer1_outputs(2861) <= not (a xor b);
    layer1_outputs(2862) <= not (a or b);
    layer1_outputs(2863) <= a and b;
    layer1_outputs(2864) <= a;
    layer1_outputs(2865) <= a or b;
    layer1_outputs(2866) <= a and not b;
    layer1_outputs(2867) <= not (a or b);
    layer1_outputs(2868) <= not (a or b);
    layer1_outputs(2869) <= b;
    layer1_outputs(2870) <= a and b;
    layer1_outputs(2871) <= a and not b;
    layer1_outputs(2872) <= b;
    layer1_outputs(2873) <= b;
    layer1_outputs(2874) <= a;
    layer1_outputs(2875) <= not (a or b);
    layer1_outputs(2876) <= not (a or b);
    layer1_outputs(2877) <= not b;
    layer1_outputs(2878) <= a or b;
    layer1_outputs(2879) <= a and not b;
    layer1_outputs(2880) <= b;
    layer1_outputs(2881) <= b and not a;
    layer1_outputs(2882) <= a or b;
    layer1_outputs(2883) <= not (a xor b);
    layer1_outputs(2884) <= not b;
    layer1_outputs(2885) <= a xor b;
    layer1_outputs(2886) <= not (a xor b);
    layer1_outputs(2887) <= not (a and b);
    layer1_outputs(2888) <= not (a or b);
    layer1_outputs(2889) <= not (a xor b);
    layer1_outputs(2890) <= a or b;
    layer1_outputs(2891) <= not a or b;
    layer1_outputs(2892) <= b;
    layer1_outputs(2893) <= a xor b;
    layer1_outputs(2894) <= not a;
    layer1_outputs(2895) <= not (a and b);
    layer1_outputs(2896) <= a or b;
    layer1_outputs(2897) <= not (a xor b);
    layer1_outputs(2898) <= a;
    layer1_outputs(2899) <= not (a or b);
    layer1_outputs(2900) <= b;
    layer1_outputs(2901) <= b;
    layer1_outputs(2902) <= not (a xor b);
    layer1_outputs(2903) <= a and not b;
    layer1_outputs(2904) <= a or b;
    layer1_outputs(2905) <= not (a and b);
    layer1_outputs(2906) <= a or b;
    layer1_outputs(2907) <= a xor b;
    layer1_outputs(2908) <= a;
    layer1_outputs(2909) <= b;
    layer1_outputs(2910) <= a;
    layer1_outputs(2911) <= a;
    layer1_outputs(2912) <= not a;
    layer1_outputs(2913) <= 1'b1;
    layer1_outputs(2914) <= not a or b;
    layer1_outputs(2915) <= a and b;
    layer1_outputs(2916) <= a and not b;
    layer1_outputs(2917) <= not b or a;
    layer1_outputs(2918) <= not a or b;
    layer1_outputs(2919) <= a and b;
    layer1_outputs(2920) <= not a;
    layer1_outputs(2921) <= a;
    layer1_outputs(2922) <= not b or a;
    layer1_outputs(2923) <= not (a and b);
    layer1_outputs(2924) <= a xor b;
    layer1_outputs(2925) <= a xor b;
    layer1_outputs(2926) <= not (a xor b);
    layer1_outputs(2927) <= b and not a;
    layer1_outputs(2928) <= not (a or b);
    layer1_outputs(2929) <= not a or b;
    layer1_outputs(2930) <= not a;
    layer1_outputs(2931) <= not a;
    layer1_outputs(2932) <= a;
    layer1_outputs(2933) <= not b or a;
    layer1_outputs(2934) <= a and b;
    layer1_outputs(2935) <= not (a and b);
    layer1_outputs(2936) <= a;
    layer1_outputs(2937) <= not b or a;
    layer1_outputs(2938) <= a or b;
    layer1_outputs(2939) <= not a;
    layer1_outputs(2940) <= 1'b1;
    layer1_outputs(2941) <= a xor b;
    layer1_outputs(2942) <= not b;
    layer1_outputs(2943) <= not b;
    layer1_outputs(2944) <= b;
    layer1_outputs(2945) <= not b;
    layer1_outputs(2946) <= a xor b;
    layer1_outputs(2947) <= a;
    layer1_outputs(2948) <= not b or a;
    layer1_outputs(2949) <= a xor b;
    layer1_outputs(2950) <= a xor b;
    layer1_outputs(2951) <= not (a and b);
    layer1_outputs(2952) <= a;
    layer1_outputs(2953) <= not a or b;
    layer1_outputs(2954) <= not b;
    layer1_outputs(2955) <= b;
    layer1_outputs(2956) <= a and not b;
    layer1_outputs(2957) <= b;
    layer1_outputs(2958) <= not b;
    layer1_outputs(2959) <= a or b;
    layer1_outputs(2960) <= not b or a;
    layer1_outputs(2961) <= a or b;
    layer1_outputs(2962) <= not (a xor b);
    layer1_outputs(2963) <= b;
    layer1_outputs(2964) <= a or b;
    layer1_outputs(2965) <= not a;
    layer1_outputs(2966) <= not b or a;
    layer1_outputs(2967) <= a xor b;
    layer1_outputs(2968) <= not a;
    layer1_outputs(2969) <= a;
    layer1_outputs(2970) <= not (a xor b);
    layer1_outputs(2971) <= not a or b;
    layer1_outputs(2972) <= not a;
    layer1_outputs(2973) <= a or b;
    layer1_outputs(2974) <= not (a or b);
    layer1_outputs(2975) <= a;
    layer1_outputs(2976) <= a or b;
    layer1_outputs(2977) <= a xor b;
    layer1_outputs(2978) <= b;
    layer1_outputs(2979) <= not b;
    layer1_outputs(2980) <= not (a and b);
    layer1_outputs(2981) <= a and not b;
    layer1_outputs(2982) <= not b or a;
    layer1_outputs(2983) <= not a or b;
    layer1_outputs(2984) <= a xor b;
    layer1_outputs(2985) <= not a or b;
    layer1_outputs(2986) <= a and b;
    layer1_outputs(2987) <= a and b;
    layer1_outputs(2988) <= a or b;
    layer1_outputs(2989) <= not (a xor b);
    layer1_outputs(2990) <= b and not a;
    layer1_outputs(2991) <= a or b;
    layer1_outputs(2992) <= not a;
    layer1_outputs(2993) <= not (a xor b);
    layer1_outputs(2994) <= not a;
    layer1_outputs(2995) <= not (a or b);
    layer1_outputs(2996) <= b and not a;
    layer1_outputs(2997) <= b;
    layer1_outputs(2998) <= not b or a;
    layer1_outputs(2999) <= not b or a;
    layer1_outputs(3000) <= a and b;
    layer1_outputs(3001) <= a and b;
    layer1_outputs(3002) <= b and not a;
    layer1_outputs(3003) <= a;
    layer1_outputs(3004) <= not a;
    layer1_outputs(3005) <= not b;
    layer1_outputs(3006) <= 1'b0;
    layer1_outputs(3007) <= not (a xor b);
    layer1_outputs(3008) <= not (a or b);
    layer1_outputs(3009) <= not b;
    layer1_outputs(3010) <= not b;
    layer1_outputs(3011) <= a;
    layer1_outputs(3012) <= not a;
    layer1_outputs(3013) <= not a;
    layer1_outputs(3014) <= a;
    layer1_outputs(3015) <= a or b;
    layer1_outputs(3016) <= a xor b;
    layer1_outputs(3017) <= a and not b;
    layer1_outputs(3018) <= not b;
    layer1_outputs(3019) <= not a;
    layer1_outputs(3020) <= not a or b;
    layer1_outputs(3021) <= not a;
    layer1_outputs(3022) <= not a;
    layer1_outputs(3023) <= not a;
    layer1_outputs(3024) <= not (a xor b);
    layer1_outputs(3025) <= not (a or b);
    layer1_outputs(3026) <= a;
    layer1_outputs(3027) <= a and not b;
    layer1_outputs(3028) <= not a;
    layer1_outputs(3029) <= a xor b;
    layer1_outputs(3030) <= a;
    layer1_outputs(3031) <= a and not b;
    layer1_outputs(3032) <= not (a or b);
    layer1_outputs(3033) <= a xor b;
    layer1_outputs(3034) <= not (a or b);
    layer1_outputs(3035) <= a xor b;
    layer1_outputs(3036) <= not b;
    layer1_outputs(3037) <= a xor b;
    layer1_outputs(3038) <= not (a xor b);
    layer1_outputs(3039) <= a and b;
    layer1_outputs(3040) <= a;
    layer1_outputs(3041) <= a;
    layer1_outputs(3042) <= a or b;
    layer1_outputs(3043) <= a and b;
    layer1_outputs(3044) <= not (a or b);
    layer1_outputs(3045) <= b;
    layer1_outputs(3046) <= not a;
    layer1_outputs(3047) <= not a or b;
    layer1_outputs(3048) <= not (a xor b);
    layer1_outputs(3049) <= a and not b;
    layer1_outputs(3050) <= not (a xor b);
    layer1_outputs(3051) <= not a;
    layer1_outputs(3052) <= not (a or b);
    layer1_outputs(3053) <= a and b;
    layer1_outputs(3054) <= b and not a;
    layer1_outputs(3055) <= not b;
    layer1_outputs(3056) <= not (a or b);
    layer1_outputs(3057) <= not (a xor b);
    layer1_outputs(3058) <= not (a or b);
    layer1_outputs(3059) <= a;
    layer1_outputs(3060) <= a and not b;
    layer1_outputs(3061) <= not (a or b);
    layer1_outputs(3062) <= not (a and b);
    layer1_outputs(3063) <= a;
    layer1_outputs(3064) <= a;
    layer1_outputs(3065) <= not a;
    layer1_outputs(3066) <= a xor b;
    layer1_outputs(3067) <= b;
    layer1_outputs(3068) <= a and b;
    layer1_outputs(3069) <= not a or b;
    layer1_outputs(3070) <= a and b;
    layer1_outputs(3071) <= not (a and b);
    layer1_outputs(3072) <= not (a and b);
    layer1_outputs(3073) <= b;
    layer1_outputs(3074) <= b;
    layer1_outputs(3075) <= a;
    layer1_outputs(3076) <= not b;
    layer1_outputs(3077) <= not (a and b);
    layer1_outputs(3078) <= not b;
    layer1_outputs(3079) <= a;
    layer1_outputs(3080) <= a and b;
    layer1_outputs(3081) <= not (a xor b);
    layer1_outputs(3082) <= a and not b;
    layer1_outputs(3083) <= a;
    layer1_outputs(3084) <= not (a and b);
    layer1_outputs(3085) <= not a;
    layer1_outputs(3086) <= a;
    layer1_outputs(3087) <= a xor b;
    layer1_outputs(3088) <= a and not b;
    layer1_outputs(3089) <= not (a and b);
    layer1_outputs(3090) <= not (a and b);
    layer1_outputs(3091) <= not (a xor b);
    layer1_outputs(3092) <= not b;
    layer1_outputs(3093) <= not (a xor b);
    layer1_outputs(3094) <= not a or b;
    layer1_outputs(3095) <= not a or b;
    layer1_outputs(3096) <= not b;
    layer1_outputs(3097) <= a or b;
    layer1_outputs(3098) <= a xor b;
    layer1_outputs(3099) <= a xor b;
    layer1_outputs(3100) <= not a;
    layer1_outputs(3101) <= not b;
    layer1_outputs(3102) <= a;
    layer1_outputs(3103) <= a;
    layer1_outputs(3104) <= b;
    layer1_outputs(3105) <= a;
    layer1_outputs(3106) <= a and not b;
    layer1_outputs(3107) <= not (a or b);
    layer1_outputs(3108) <= a and b;
    layer1_outputs(3109) <= not (a xor b);
    layer1_outputs(3110) <= not (a and b);
    layer1_outputs(3111) <= not (a or b);
    layer1_outputs(3112) <= not (a xor b);
    layer1_outputs(3113) <= not (a and b);
    layer1_outputs(3114) <= not (a and b);
    layer1_outputs(3115) <= not a or b;
    layer1_outputs(3116) <= not (a xor b);
    layer1_outputs(3117) <= a xor b;
    layer1_outputs(3118) <= not (a and b);
    layer1_outputs(3119) <= not (a and b);
    layer1_outputs(3120) <= not b;
    layer1_outputs(3121) <= not (a or b);
    layer1_outputs(3122) <= 1'b1;
    layer1_outputs(3123) <= not (a and b);
    layer1_outputs(3124) <= not (a or b);
    layer1_outputs(3125) <= not (a xor b);
    layer1_outputs(3126) <= b;
    layer1_outputs(3127) <= not a or b;
    layer1_outputs(3128) <= a and b;
    layer1_outputs(3129) <= not a;
    layer1_outputs(3130) <= not a;
    layer1_outputs(3131) <= a and b;
    layer1_outputs(3132) <= not (a or b);
    layer1_outputs(3133) <= a;
    layer1_outputs(3134) <= not (a xor b);
    layer1_outputs(3135) <= not a;
    layer1_outputs(3136) <= a or b;
    layer1_outputs(3137) <= not b;
    layer1_outputs(3138) <= not a;
    layer1_outputs(3139) <= not (a xor b);
    layer1_outputs(3140) <= not (a or b);
    layer1_outputs(3141) <= not (a and b);
    layer1_outputs(3142) <= a and not b;
    layer1_outputs(3143) <= not a or b;
    layer1_outputs(3144) <= not a;
    layer1_outputs(3145) <= a and not b;
    layer1_outputs(3146) <= a and not b;
    layer1_outputs(3147) <= a or b;
    layer1_outputs(3148) <= not a;
    layer1_outputs(3149) <= not a;
    layer1_outputs(3150) <= a;
    layer1_outputs(3151) <= not a or b;
    layer1_outputs(3152) <= a and not b;
    layer1_outputs(3153) <= not a;
    layer1_outputs(3154) <= a and b;
    layer1_outputs(3155) <= not (a xor b);
    layer1_outputs(3156) <= not b or a;
    layer1_outputs(3157) <= a;
    layer1_outputs(3158) <= a or b;
    layer1_outputs(3159) <= not a;
    layer1_outputs(3160) <= not (a xor b);
    layer1_outputs(3161) <= a;
    layer1_outputs(3162) <= a xor b;
    layer1_outputs(3163) <= not (a and b);
    layer1_outputs(3164) <= not (a or b);
    layer1_outputs(3165) <= not b;
    layer1_outputs(3166) <= a xor b;
    layer1_outputs(3167) <= not (a xor b);
    layer1_outputs(3168) <= a and b;
    layer1_outputs(3169) <= not (a and b);
    layer1_outputs(3170) <= not b;
    layer1_outputs(3171) <= 1'b0;
    layer1_outputs(3172) <= not (a and b);
    layer1_outputs(3173) <= not a or b;
    layer1_outputs(3174) <= not a or b;
    layer1_outputs(3175) <= not (a and b);
    layer1_outputs(3176) <= not (a xor b);
    layer1_outputs(3177) <= not (a and b);
    layer1_outputs(3178) <= b;
    layer1_outputs(3179) <= a;
    layer1_outputs(3180) <= a and b;
    layer1_outputs(3181) <= not a;
    layer1_outputs(3182) <= b;
    layer1_outputs(3183) <= a;
    layer1_outputs(3184) <= not (a or b);
    layer1_outputs(3185) <= not b;
    layer1_outputs(3186) <= 1'b1;
    layer1_outputs(3187) <= not (a or b);
    layer1_outputs(3188) <= not a;
    layer1_outputs(3189) <= not b;
    layer1_outputs(3190) <= not (a xor b);
    layer1_outputs(3191) <= not (a and b);
    layer1_outputs(3192) <= b and not a;
    layer1_outputs(3193) <= b;
    layer1_outputs(3194) <= a xor b;
    layer1_outputs(3195) <= not b or a;
    layer1_outputs(3196) <= not b;
    layer1_outputs(3197) <= not b;
    layer1_outputs(3198) <= b and not a;
    layer1_outputs(3199) <= not a;
    layer1_outputs(3200) <= a and b;
    layer1_outputs(3201) <= not (a and b);
    layer1_outputs(3202) <= not (a or b);
    layer1_outputs(3203) <= not (a or b);
    layer1_outputs(3204) <= not a or b;
    layer1_outputs(3205) <= a;
    layer1_outputs(3206) <= not (a xor b);
    layer1_outputs(3207) <= not a or b;
    layer1_outputs(3208) <= not b;
    layer1_outputs(3209) <= a or b;
    layer1_outputs(3210) <= b and not a;
    layer1_outputs(3211) <= b;
    layer1_outputs(3212) <= not (a xor b);
    layer1_outputs(3213) <= not (a and b);
    layer1_outputs(3214) <= not (a or b);
    layer1_outputs(3215) <= a;
    layer1_outputs(3216) <= not b or a;
    layer1_outputs(3217) <= not a;
    layer1_outputs(3218) <= not a;
    layer1_outputs(3219) <= not (a or b);
    layer1_outputs(3220) <= not (a xor b);
    layer1_outputs(3221) <= not a;
    layer1_outputs(3222) <= 1'b1;
    layer1_outputs(3223) <= not (a and b);
    layer1_outputs(3224) <= a and b;
    layer1_outputs(3225) <= not b or a;
    layer1_outputs(3226) <= a xor b;
    layer1_outputs(3227) <= not a;
    layer1_outputs(3228) <= not (a xor b);
    layer1_outputs(3229) <= a and b;
    layer1_outputs(3230) <= not (a or b);
    layer1_outputs(3231) <= not b;
    layer1_outputs(3232) <= not b or a;
    layer1_outputs(3233) <= a;
    layer1_outputs(3234) <= a or b;
    layer1_outputs(3235) <= not b or a;
    layer1_outputs(3236) <= a or b;
    layer1_outputs(3237) <= a;
    layer1_outputs(3238) <= b;
    layer1_outputs(3239) <= b;
    layer1_outputs(3240) <= not b or a;
    layer1_outputs(3241) <= a;
    layer1_outputs(3242) <= a;
    layer1_outputs(3243) <= a xor b;
    layer1_outputs(3244) <= not a;
    layer1_outputs(3245) <= not a or b;
    layer1_outputs(3246) <= a or b;
    layer1_outputs(3247) <= b;
    layer1_outputs(3248) <= not a;
    layer1_outputs(3249) <= a or b;
    layer1_outputs(3250) <= a and b;
    layer1_outputs(3251) <= not a;
    layer1_outputs(3252) <= not a;
    layer1_outputs(3253) <= not b or a;
    layer1_outputs(3254) <= not a or b;
    layer1_outputs(3255) <= not a or b;
    layer1_outputs(3256) <= a and not b;
    layer1_outputs(3257) <= b and not a;
    layer1_outputs(3258) <= not (a xor b);
    layer1_outputs(3259) <= not (a and b);
    layer1_outputs(3260) <= not a;
    layer1_outputs(3261) <= b;
    layer1_outputs(3262) <= not a;
    layer1_outputs(3263) <= not a;
    layer1_outputs(3264) <= a;
    layer1_outputs(3265) <= b;
    layer1_outputs(3266) <= b;
    layer1_outputs(3267) <= not (a and b);
    layer1_outputs(3268) <= not b or a;
    layer1_outputs(3269) <= b;
    layer1_outputs(3270) <= 1'b0;
    layer1_outputs(3271) <= a or b;
    layer1_outputs(3272) <= not a or b;
    layer1_outputs(3273) <= a and b;
    layer1_outputs(3274) <= not a or b;
    layer1_outputs(3275) <= not b;
    layer1_outputs(3276) <= not a or b;
    layer1_outputs(3277) <= a and not b;
    layer1_outputs(3278) <= a xor b;
    layer1_outputs(3279) <= a and b;
    layer1_outputs(3280) <= b and not a;
    layer1_outputs(3281) <= b;
    layer1_outputs(3282) <= 1'b0;
    layer1_outputs(3283) <= a or b;
    layer1_outputs(3284) <= a and not b;
    layer1_outputs(3285) <= not b;
    layer1_outputs(3286) <= a;
    layer1_outputs(3287) <= not (a or b);
    layer1_outputs(3288) <= a xor b;
    layer1_outputs(3289) <= a xor b;
    layer1_outputs(3290) <= not (a xor b);
    layer1_outputs(3291) <= not b or a;
    layer1_outputs(3292) <= b and not a;
    layer1_outputs(3293) <= not (a xor b);
    layer1_outputs(3294) <= b and not a;
    layer1_outputs(3295) <= a xor b;
    layer1_outputs(3296) <= b;
    layer1_outputs(3297) <= b;
    layer1_outputs(3298) <= not b;
    layer1_outputs(3299) <= a;
    layer1_outputs(3300) <= not b;
    layer1_outputs(3301) <= not a;
    layer1_outputs(3302) <= not b;
    layer1_outputs(3303) <= a;
    layer1_outputs(3304) <= not (a or b);
    layer1_outputs(3305) <= not a;
    layer1_outputs(3306) <= not (a xor b);
    layer1_outputs(3307) <= a or b;
    layer1_outputs(3308) <= not b or a;
    layer1_outputs(3309) <= not (a or b);
    layer1_outputs(3310) <= a;
    layer1_outputs(3311) <= not b;
    layer1_outputs(3312) <= not (a or b);
    layer1_outputs(3313) <= not b;
    layer1_outputs(3314) <= not a;
    layer1_outputs(3315) <= a and b;
    layer1_outputs(3316) <= a and not b;
    layer1_outputs(3317) <= not (a and b);
    layer1_outputs(3318) <= not a or b;
    layer1_outputs(3319) <= not a;
    layer1_outputs(3320) <= not (a and b);
    layer1_outputs(3321) <= not a or b;
    layer1_outputs(3322) <= not a;
    layer1_outputs(3323) <= not (a and b);
    layer1_outputs(3324) <= a or b;
    layer1_outputs(3325) <= not (a xor b);
    layer1_outputs(3326) <= not (a xor b);
    layer1_outputs(3327) <= a and b;
    layer1_outputs(3328) <= a and b;
    layer1_outputs(3329) <= a and not b;
    layer1_outputs(3330) <= a;
    layer1_outputs(3331) <= b and not a;
    layer1_outputs(3332) <= b;
    layer1_outputs(3333) <= b;
    layer1_outputs(3334) <= a;
    layer1_outputs(3335) <= b;
    layer1_outputs(3336) <= 1'b0;
    layer1_outputs(3337) <= not a;
    layer1_outputs(3338) <= b and not a;
    layer1_outputs(3339) <= a and b;
    layer1_outputs(3340) <= not b;
    layer1_outputs(3341) <= a;
    layer1_outputs(3342) <= not b;
    layer1_outputs(3343) <= not (a or b);
    layer1_outputs(3344) <= a;
    layer1_outputs(3345) <= not a;
    layer1_outputs(3346) <= not (a xor b);
    layer1_outputs(3347) <= not a;
    layer1_outputs(3348) <= a;
    layer1_outputs(3349) <= a xor b;
    layer1_outputs(3350) <= a or b;
    layer1_outputs(3351) <= a;
    layer1_outputs(3352) <= a;
    layer1_outputs(3353) <= not a;
    layer1_outputs(3354) <= not b;
    layer1_outputs(3355) <= not b or a;
    layer1_outputs(3356) <= not (a xor b);
    layer1_outputs(3357) <= not b or a;
    layer1_outputs(3358) <= not (a xor b);
    layer1_outputs(3359) <= a;
    layer1_outputs(3360) <= not (a and b);
    layer1_outputs(3361) <= a xor b;
    layer1_outputs(3362) <= a xor b;
    layer1_outputs(3363) <= a xor b;
    layer1_outputs(3364) <= b;
    layer1_outputs(3365) <= not a or b;
    layer1_outputs(3366) <= a and not b;
    layer1_outputs(3367) <= a xor b;
    layer1_outputs(3368) <= a xor b;
    layer1_outputs(3369) <= not a;
    layer1_outputs(3370) <= not b;
    layer1_outputs(3371) <= a or b;
    layer1_outputs(3372) <= not a or b;
    layer1_outputs(3373) <= a;
    layer1_outputs(3374) <= not a or b;
    layer1_outputs(3375) <= a and not b;
    layer1_outputs(3376) <= a and not b;
    layer1_outputs(3377) <= a and not b;
    layer1_outputs(3378) <= not a;
    layer1_outputs(3379) <= a and not b;
    layer1_outputs(3380) <= not (a and b);
    layer1_outputs(3381) <= not (a xor b);
    layer1_outputs(3382) <= b and not a;
    layer1_outputs(3383) <= a;
    layer1_outputs(3384) <= a;
    layer1_outputs(3385) <= not b;
    layer1_outputs(3386) <= a xor b;
    layer1_outputs(3387) <= not a;
    layer1_outputs(3388) <= not b or a;
    layer1_outputs(3389) <= a;
    layer1_outputs(3390) <= not (a or b);
    layer1_outputs(3391) <= not b;
    layer1_outputs(3392) <= not b or a;
    layer1_outputs(3393) <= not (a and b);
    layer1_outputs(3394) <= a;
    layer1_outputs(3395) <= not a;
    layer1_outputs(3396) <= not (a and b);
    layer1_outputs(3397) <= not (a and b);
    layer1_outputs(3398) <= b and not a;
    layer1_outputs(3399) <= a and b;
    layer1_outputs(3400) <= not a or b;
    layer1_outputs(3401) <= not b;
    layer1_outputs(3402) <= b and not a;
    layer1_outputs(3403) <= a and not b;
    layer1_outputs(3404) <= not (a xor b);
    layer1_outputs(3405) <= a xor b;
    layer1_outputs(3406) <= a;
    layer1_outputs(3407) <= not a;
    layer1_outputs(3408) <= a and not b;
    layer1_outputs(3409) <= not (a and b);
    layer1_outputs(3410) <= not (a xor b);
    layer1_outputs(3411) <= not (a xor b);
    layer1_outputs(3412) <= b and not a;
    layer1_outputs(3413) <= 1'b1;
    layer1_outputs(3414) <= a and not b;
    layer1_outputs(3415) <= a;
    layer1_outputs(3416) <= a;
    layer1_outputs(3417) <= b and not a;
    layer1_outputs(3418) <= a and b;
    layer1_outputs(3419) <= b and not a;
    layer1_outputs(3420) <= not b or a;
    layer1_outputs(3421) <= not b or a;
    layer1_outputs(3422) <= not a;
    layer1_outputs(3423) <= 1'b1;
    layer1_outputs(3424) <= not (a xor b);
    layer1_outputs(3425) <= a;
    layer1_outputs(3426) <= a and not b;
    layer1_outputs(3427) <= b and not a;
    layer1_outputs(3428) <= a or b;
    layer1_outputs(3429) <= a;
    layer1_outputs(3430) <= a;
    layer1_outputs(3431) <= not b;
    layer1_outputs(3432) <= b;
    layer1_outputs(3433) <= not (a and b);
    layer1_outputs(3434) <= a and not b;
    layer1_outputs(3435) <= not (a xor b);
    layer1_outputs(3436) <= not b or a;
    layer1_outputs(3437) <= not (a and b);
    layer1_outputs(3438) <= not (a or b);
    layer1_outputs(3439) <= not (a xor b);
    layer1_outputs(3440) <= not (a xor b);
    layer1_outputs(3441) <= not b or a;
    layer1_outputs(3442) <= a xor b;
    layer1_outputs(3443) <= a or b;
    layer1_outputs(3444) <= not a or b;
    layer1_outputs(3445) <= a;
    layer1_outputs(3446) <= a or b;
    layer1_outputs(3447) <= b and not a;
    layer1_outputs(3448) <= a or b;
    layer1_outputs(3449) <= not a or b;
    layer1_outputs(3450) <= not b or a;
    layer1_outputs(3451) <= not (a or b);
    layer1_outputs(3452) <= not a;
    layer1_outputs(3453) <= not (a xor b);
    layer1_outputs(3454) <= not b;
    layer1_outputs(3455) <= a xor b;
    layer1_outputs(3456) <= b and not a;
    layer1_outputs(3457) <= b;
    layer1_outputs(3458) <= not b;
    layer1_outputs(3459) <= not (a xor b);
    layer1_outputs(3460) <= b;
    layer1_outputs(3461) <= a;
    layer1_outputs(3462) <= a xor b;
    layer1_outputs(3463) <= not (a xor b);
    layer1_outputs(3464) <= not (a or b);
    layer1_outputs(3465) <= a and not b;
    layer1_outputs(3466) <= not (a and b);
    layer1_outputs(3467) <= b;
    layer1_outputs(3468) <= not a;
    layer1_outputs(3469) <= not (a xor b);
    layer1_outputs(3470) <= a;
    layer1_outputs(3471) <= not a;
    layer1_outputs(3472) <= a xor b;
    layer1_outputs(3473) <= a xor b;
    layer1_outputs(3474) <= b;
    layer1_outputs(3475) <= a;
    layer1_outputs(3476) <= not a or b;
    layer1_outputs(3477) <= not a;
    layer1_outputs(3478) <= not (a xor b);
    layer1_outputs(3479) <= not a;
    layer1_outputs(3480) <= a xor b;
    layer1_outputs(3481) <= b and not a;
    layer1_outputs(3482) <= a;
    layer1_outputs(3483) <= a and b;
    layer1_outputs(3484) <= a;
    layer1_outputs(3485) <= not a;
    layer1_outputs(3486) <= not (a or b);
    layer1_outputs(3487) <= a xor b;
    layer1_outputs(3488) <= a and not b;
    layer1_outputs(3489) <= not b or a;
    layer1_outputs(3490) <= not b;
    layer1_outputs(3491) <= a or b;
    layer1_outputs(3492) <= a and not b;
    layer1_outputs(3493) <= 1'b0;
    layer1_outputs(3494) <= not a or b;
    layer1_outputs(3495) <= a or b;
    layer1_outputs(3496) <= a or b;
    layer1_outputs(3497) <= b;
    layer1_outputs(3498) <= a xor b;
    layer1_outputs(3499) <= a or b;
    layer1_outputs(3500) <= a and b;
    layer1_outputs(3501) <= a;
    layer1_outputs(3502) <= b;
    layer1_outputs(3503) <= not b or a;
    layer1_outputs(3504) <= a and b;
    layer1_outputs(3505) <= not b;
    layer1_outputs(3506) <= not (a or b);
    layer1_outputs(3507) <= a or b;
    layer1_outputs(3508) <= not b or a;
    layer1_outputs(3509) <= not (a xor b);
    layer1_outputs(3510) <= b;
    layer1_outputs(3511) <= a xor b;
    layer1_outputs(3512) <= not (a or b);
    layer1_outputs(3513) <= a or b;
    layer1_outputs(3514) <= a or b;
    layer1_outputs(3515) <= a and not b;
    layer1_outputs(3516) <= a;
    layer1_outputs(3517) <= b;
    layer1_outputs(3518) <= not (a and b);
    layer1_outputs(3519) <= not (a xor b);
    layer1_outputs(3520) <= not b or a;
    layer1_outputs(3521) <= b;
    layer1_outputs(3522) <= not (a and b);
    layer1_outputs(3523) <= 1'b1;
    layer1_outputs(3524) <= a xor b;
    layer1_outputs(3525) <= not b or a;
    layer1_outputs(3526) <= a;
    layer1_outputs(3527) <= b;
    layer1_outputs(3528) <= a xor b;
    layer1_outputs(3529) <= not (a and b);
    layer1_outputs(3530) <= not b or a;
    layer1_outputs(3531) <= not b or a;
    layer1_outputs(3532) <= b;
    layer1_outputs(3533) <= not (a or b);
    layer1_outputs(3534) <= a and b;
    layer1_outputs(3535) <= not (a and b);
    layer1_outputs(3536) <= a xor b;
    layer1_outputs(3537) <= a or b;
    layer1_outputs(3538) <= a and not b;
    layer1_outputs(3539) <= a;
    layer1_outputs(3540) <= not a;
    layer1_outputs(3541) <= a and not b;
    layer1_outputs(3542) <= a or b;
    layer1_outputs(3543) <= b;
    layer1_outputs(3544) <= not (a or b);
    layer1_outputs(3545) <= not (a xor b);
    layer1_outputs(3546) <= a xor b;
    layer1_outputs(3547) <= not b;
    layer1_outputs(3548) <= a or b;
    layer1_outputs(3549) <= b;
    layer1_outputs(3550) <= a xor b;
    layer1_outputs(3551) <= not a;
    layer1_outputs(3552) <= a and not b;
    layer1_outputs(3553) <= not b;
    layer1_outputs(3554) <= not (a or b);
    layer1_outputs(3555) <= not b;
    layer1_outputs(3556) <= b;
    layer1_outputs(3557) <= a;
    layer1_outputs(3558) <= not a;
    layer1_outputs(3559) <= not (a and b);
    layer1_outputs(3560) <= a and b;
    layer1_outputs(3561) <= not b;
    layer1_outputs(3562) <= a;
    layer1_outputs(3563) <= not (a and b);
    layer1_outputs(3564) <= not b or a;
    layer1_outputs(3565) <= not (a xor b);
    layer1_outputs(3566) <= a and not b;
    layer1_outputs(3567) <= not (a and b);
    layer1_outputs(3568) <= b;
    layer1_outputs(3569) <= b;
    layer1_outputs(3570) <= b;
    layer1_outputs(3571) <= b;
    layer1_outputs(3572) <= not a;
    layer1_outputs(3573) <= not (a or b);
    layer1_outputs(3574) <= b and not a;
    layer1_outputs(3575) <= a xor b;
    layer1_outputs(3576) <= not b;
    layer1_outputs(3577) <= not b;
    layer1_outputs(3578) <= not a;
    layer1_outputs(3579) <= not a;
    layer1_outputs(3580) <= not (a or b);
    layer1_outputs(3581) <= b and not a;
    layer1_outputs(3582) <= not a or b;
    layer1_outputs(3583) <= b and not a;
    layer1_outputs(3584) <= not b;
    layer1_outputs(3585) <= not (a xor b);
    layer1_outputs(3586) <= not b;
    layer1_outputs(3587) <= a xor b;
    layer1_outputs(3588) <= a or b;
    layer1_outputs(3589) <= not b;
    layer1_outputs(3590) <= b and not a;
    layer1_outputs(3591) <= b;
    layer1_outputs(3592) <= not a or b;
    layer1_outputs(3593) <= a xor b;
    layer1_outputs(3594) <= not b;
    layer1_outputs(3595) <= a;
    layer1_outputs(3596) <= not a or b;
    layer1_outputs(3597) <= b;
    layer1_outputs(3598) <= not b or a;
    layer1_outputs(3599) <= not (a xor b);
    layer1_outputs(3600) <= not (a xor b);
    layer1_outputs(3601) <= not (a and b);
    layer1_outputs(3602) <= 1'b1;
    layer1_outputs(3603) <= not b;
    layer1_outputs(3604) <= a or b;
    layer1_outputs(3605) <= not a;
    layer1_outputs(3606) <= a xor b;
    layer1_outputs(3607) <= not (a and b);
    layer1_outputs(3608) <= not b;
    layer1_outputs(3609) <= not b or a;
    layer1_outputs(3610) <= not a;
    layer1_outputs(3611) <= not b;
    layer1_outputs(3612) <= not a;
    layer1_outputs(3613) <= b;
    layer1_outputs(3614) <= not a;
    layer1_outputs(3615) <= not (a and b);
    layer1_outputs(3616) <= not (a or b);
    layer1_outputs(3617) <= not a;
    layer1_outputs(3618) <= a xor b;
    layer1_outputs(3619) <= a xor b;
    layer1_outputs(3620) <= a;
    layer1_outputs(3621) <= b;
    layer1_outputs(3622) <= not a;
    layer1_outputs(3623) <= a;
    layer1_outputs(3624) <= not a;
    layer1_outputs(3625) <= b;
    layer1_outputs(3626) <= not b;
    layer1_outputs(3627) <= not b;
    layer1_outputs(3628) <= not a or b;
    layer1_outputs(3629) <= not b;
    layer1_outputs(3630) <= a and not b;
    layer1_outputs(3631) <= not a or b;
    layer1_outputs(3632) <= b and not a;
    layer1_outputs(3633) <= a;
    layer1_outputs(3634) <= not a;
    layer1_outputs(3635) <= not b;
    layer1_outputs(3636) <= not b;
    layer1_outputs(3637) <= not (a xor b);
    layer1_outputs(3638) <= not (a xor b);
    layer1_outputs(3639) <= not b;
    layer1_outputs(3640) <= a or b;
    layer1_outputs(3641) <= not (a and b);
    layer1_outputs(3642) <= a and not b;
    layer1_outputs(3643) <= not (a or b);
    layer1_outputs(3644) <= not b;
    layer1_outputs(3645) <= not b or a;
    layer1_outputs(3646) <= a xor b;
    layer1_outputs(3647) <= a and not b;
    layer1_outputs(3648) <= not a;
    layer1_outputs(3649) <= not (a and b);
    layer1_outputs(3650) <= not (a or b);
    layer1_outputs(3651) <= not b or a;
    layer1_outputs(3652) <= b;
    layer1_outputs(3653) <= b;
    layer1_outputs(3654) <= a or b;
    layer1_outputs(3655) <= not a or b;
    layer1_outputs(3656) <= a and b;
    layer1_outputs(3657) <= a and b;
    layer1_outputs(3658) <= not b;
    layer1_outputs(3659) <= not b;
    layer1_outputs(3660) <= not a;
    layer1_outputs(3661) <= a and not b;
    layer1_outputs(3662) <= a xor b;
    layer1_outputs(3663) <= b;
    layer1_outputs(3664) <= not b;
    layer1_outputs(3665) <= not (a xor b);
    layer1_outputs(3666) <= a;
    layer1_outputs(3667) <= a or b;
    layer1_outputs(3668) <= a xor b;
    layer1_outputs(3669) <= not (a and b);
    layer1_outputs(3670) <= b and not a;
    layer1_outputs(3671) <= a xor b;
    layer1_outputs(3672) <= a;
    layer1_outputs(3673) <= b and not a;
    layer1_outputs(3674) <= a and not b;
    layer1_outputs(3675) <= a and b;
    layer1_outputs(3676) <= a or b;
    layer1_outputs(3677) <= not b;
    layer1_outputs(3678) <= a xor b;
    layer1_outputs(3679) <= b and not a;
    layer1_outputs(3680) <= b and not a;
    layer1_outputs(3681) <= not b or a;
    layer1_outputs(3682) <= a and b;
    layer1_outputs(3683) <= a and b;
    layer1_outputs(3684) <= a or b;
    layer1_outputs(3685) <= b;
    layer1_outputs(3686) <= 1'b0;
    layer1_outputs(3687) <= not (a xor b);
    layer1_outputs(3688) <= not a;
    layer1_outputs(3689) <= a;
    layer1_outputs(3690) <= not b;
    layer1_outputs(3691) <= not b;
    layer1_outputs(3692) <= a;
    layer1_outputs(3693) <= b;
    layer1_outputs(3694) <= not (a and b);
    layer1_outputs(3695) <= b and not a;
    layer1_outputs(3696) <= a;
    layer1_outputs(3697) <= not b;
    layer1_outputs(3698) <= not (a and b);
    layer1_outputs(3699) <= b and not a;
    layer1_outputs(3700) <= not (a xor b);
    layer1_outputs(3701) <= not a;
    layer1_outputs(3702) <= not b;
    layer1_outputs(3703) <= a xor b;
    layer1_outputs(3704) <= not a;
    layer1_outputs(3705) <= a or b;
    layer1_outputs(3706) <= not (a and b);
    layer1_outputs(3707) <= a or b;
    layer1_outputs(3708) <= a or b;
    layer1_outputs(3709) <= a and not b;
    layer1_outputs(3710) <= not (a xor b);
    layer1_outputs(3711) <= not a or b;
    layer1_outputs(3712) <= a and not b;
    layer1_outputs(3713) <= not b;
    layer1_outputs(3714) <= not b;
    layer1_outputs(3715) <= b;
    layer1_outputs(3716) <= b;
    layer1_outputs(3717) <= not (a or b);
    layer1_outputs(3718) <= b;
    layer1_outputs(3719) <= not a;
    layer1_outputs(3720) <= a and b;
    layer1_outputs(3721) <= a and b;
    layer1_outputs(3722) <= a or b;
    layer1_outputs(3723) <= a and not b;
    layer1_outputs(3724) <= not b or a;
    layer1_outputs(3725) <= a xor b;
    layer1_outputs(3726) <= a and not b;
    layer1_outputs(3727) <= not b;
    layer1_outputs(3728) <= a and b;
    layer1_outputs(3729) <= not a;
    layer1_outputs(3730) <= not b or a;
    layer1_outputs(3731) <= not (a and b);
    layer1_outputs(3732) <= not (a or b);
    layer1_outputs(3733) <= a xor b;
    layer1_outputs(3734) <= not b;
    layer1_outputs(3735) <= not a;
    layer1_outputs(3736) <= b;
    layer1_outputs(3737) <= not b or a;
    layer1_outputs(3738) <= not (a or b);
    layer1_outputs(3739) <= not b or a;
    layer1_outputs(3740) <= a;
    layer1_outputs(3741) <= not b;
    layer1_outputs(3742) <= a and not b;
    layer1_outputs(3743) <= a;
    layer1_outputs(3744) <= not a;
    layer1_outputs(3745) <= a and not b;
    layer1_outputs(3746) <= a and b;
    layer1_outputs(3747) <= not a or b;
    layer1_outputs(3748) <= a or b;
    layer1_outputs(3749) <= not a;
    layer1_outputs(3750) <= a xor b;
    layer1_outputs(3751) <= a xor b;
    layer1_outputs(3752) <= not b;
    layer1_outputs(3753) <= b;
    layer1_outputs(3754) <= not a or b;
    layer1_outputs(3755) <= not a or b;
    layer1_outputs(3756) <= a and b;
    layer1_outputs(3757) <= 1'b0;
    layer1_outputs(3758) <= not a or b;
    layer1_outputs(3759) <= 1'b1;
    layer1_outputs(3760) <= a and b;
    layer1_outputs(3761) <= not b;
    layer1_outputs(3762) <= not b;
    layer1_outputs(3763) <= not a;
    layer1_outputs(3764) <= a and not b;
    layer1_outputs(3765) <= a xor b;
    layer1_outputs(3766) <= a xor b;
    layer1_outputs(3767) <= not (a xor b);
    layer1_outputs(3768) <= a;
    layer1_outputs(3769) <= a and b;
    layer1_outputs(3770) <= b and not a;
    layer1_outputs(3771) <= a or b;
    layer1_outputs(3772) <= a;
    layer1_outputs(3773) <= not b;
    layer1_outputs(3774) <= b and not a;
    layer1_outputs(3775) <= not (a xor b);
    layer1_outputs(3776) <= a or b;
    layer1_outputs(3777) <= a xor b;
    layer1_outputs(3778) <= b;
    layer1_outputs(3779) <= not a or b;
    layer1_outputs(3780) <= b;
    layer1_outputs(3781) <= not (a and b);
    layer1_outputs(3782) <= a or b;
    layer1_outputs(3783) <= not b;
    layer1_outputs(3784) <= not (a xor b);
    layer1_outputs(3785) <= b and not a;
    layer1_outputs(3786) <= a;
    layer1_outputs(3787) <= not a or b;
    layer1_outputs(3788) <= a xor b;
    layer1_outputs(3789) <= not a;
    layer1_outputs(3790) <= a;
    layer1_outputs(3791) <= a xor b;
    layer1_outputs(3792) <= a and b;
    layer1_outputs(3793) <= 1'b1;
    layer1_outputs(3794) <= a xor b;
    layer1_outputs(3795) <= 1'b0;
    layer1_outputs(3796) <= not b or a;
    layer1_outputs(3797) <= b;
    layer1_outputs(3798) <= a;
    layer1_outputs(3799) <= not b or a;
    layer1_outputs(3800) <= not a or b;
    layer1_outputs(3801) <= not a;
    layer1_outputs(3802) <= not (a or b);
    layer1_outputs(3803) <= a;
    layer1_outputs(3804) <= not a;
    layer1_outputs(3805) <= a xor b;
    layer1_outputs(3806) <= b;
    layer1_outputs(3807) <= not a;
    layer1_outputs(3808) <= a;
    layer1_outputs(3809) <= not a;
    layer1_outputs(3810) <= a;
    layer1_outputs(3811) <= a or b;
    layer1_outputs(3812) <= not (a or b);
    layer1_outputs(3813) <= not b or a;
    layer1_outputs(3814) <= not (a xor b);
    layer1_outputs(3815) <= a and b;
    layer1_outputs(3816) <= a and b;
    layer1_outputs(3817) <= b and not a;
    layer1_outputs(3818) <= b;
    layer1_outputs(3819) <= b;
    layer1_outputs(3820) <= b;
    layer1_outputs(3821) <= b;
    layer1_outputs(3822) <= a or b;
    layer1_outputs(3823) <= a;
    layer1_outputs(3824) <= a and b;
    layer1_outputs(3825) <= not (a xor b);
    layer1_outputs(3826) <= not b or a;
    layer1_outputs(3827) <= not (a and b);
    layer1_outputs(3828) <= not (a xor b);
    layer1_outputs(3829) <= a and not b;
    layer1_outputs(3830) <= not (a xor b);
    layer1_outputs(3831) <= not b;
    layer1_outputs(3832) <= a;
    layer1_outputs(3833) <= not (a or b);
    layer1_outputs(3834) <= not b or a;
    layer1_outputs(3835) <= b;
    layer1_outputs(3836) <= b and not a;
    layer1_outputs(3837) <= not a;
    layer1_outputs(3838) <= not (a or b);
    layer1_outputs(3839) <= not a or b;
    layer1_outputs(3840) <= not b or a;
    layer1_outputs(3841) <= a;
    layer1_outputs(3842) <= b and not a;
    layer1_outputs(3843) <= b;
    layer1_outputs(3844) <= a and b;
    layer1_outputs(3845) <= not (a or b);
    layer1_outputs(3846) <= not b or a;
    layer1_outputs(3847) <= not a or b;
    layer1_outputs(3848) <= not b or a;
    layer1_outputs(3849) <= a;
    layer1_outputs(3850) <= not (a xor b);
    layer1_outputs(3851) <= not b or a;
    layer1_outputs(3852) <= not (a xor b);
    layer1_outputs(3853) <= b;
    layer1_outputs(3854) <= a;
    layer1_outputs(3855) <= a;
    layer1_outputs(3856) <= not a or b;
    layer1_outputs(3857) <= b;
    layer1_outputs(3858) <= a or b;
    layer1_outputs(3859) <= b;
    layer1_outputs(3860) <= not b;
    layer1_outputs(3861) <= not a;
    layer1_outputs(3862) <= not (a or b);
    layer1_outputs(3863) <= not b;
    layer1_outputs(3864) <= not b;
    layer1_outputs(3865) <= b;
    layer1_outputs(3866) <= not a;
    layer1_outputs(3867) <= not b or a;
    layer1_outputs(3868) <= not a;
    layer1_outputs(3869) <= not (a and b);
    layer1_outputs(3870) <= not a or b;
    layer1_outputs(3871) <= a or b;
    layer1_outputs(3872) <= a xor b;
    layer1_outputs(3873) <= b;
    layer1_outputs(3874) <= a and b;
    layer1_outputs(3875) <= not a;
    layer1_outputs(3876) <= not (a xor b);
    layer1_outputs(3877) <= a;
    layer1_outputs(3878) <= a and not b;
    layer1_outputs(3879) <= a;
    layer1_outputs(3880) <= a xor b;
    layer1_outputs(3881) <= not (a and b);
    layer1_outputs(3882) <= a and b;
    layer1_outputs(3883) <= not (a xor b);
    layer1_outputs(3884) <= b;
    layer1_outputs(3885) <= b;
    layer1_outputs(3886) <= not a or b;
    layer1_outputs(3887) <= a and b;
    layer1_outputs(3888) <= not (a or b);
    layer1_outputs(3889) <= not b;
    layer1_outputs(3890) <= not a;
    layer1_outputs(3891) <= 1'b1;
    layer1_outputs(3892) <= not a;
    layer1_outputs(3893) <= a or b;
    layer1_outputs(3894) <= not (a or b);
    layer1_outputs(3895) <= not a or b;
    layer1_outputs(3896) <= a and b;
    layer1_outputs(3897) <= not b;
    layer1_outputs(3898) <= a;
    layer1_outputs(3899) <= b;
    layer1_outputs(3900) <= not a;
    layer1_outputs(3901) <= a xor b;
    layer1_outputs(3902) <= not b;
    layer1_outputs(3903) <= b;
    layer1_outputs(3904) <= not (a and b);
    layer1_outputs(3905) <= a;
    layer1_outputs(3906) <= a;
    layer1_outputs(3907) <= a and not b;
    layer1_outputs(3908) <= not b or a;
    layer1_outputs(3909) <= not (a xor b);
    layer1_outputs(3910) <= b;
    layer1_outputs(3911) <= 1'b1;
    layer1_outputs(3912) <= b;
    layer1_outputs(3913) <= not (a or b);
    layer1_outputs(3914) <= not (a xor b);
    layer1_outputs(3915) <= not (a and b);
    layer1_outputs(3916) <= not a;
    layer1_outputs(3917) <= not b;
    layer1_outputs(3918) <= b;
    layer1_outputs(3919) <= not b or a;
    layer1_outputs(3920) <= a and b;
    layer1_outputs(3921) <= a and not b;
    layer1_outputs(3922) <= not (a xor b);
    layer1_outputs(3923) <= not (a xor b);
    layer1_outputs(3924) <= not (a xor b);
    layer1_outputs(3925) <= a and b;
    layer1_outputs(3926) <= not (a and b);
    layer1_outputs(3927) <= b;
    layer1_outputs(3928) <= a and not b;
    layer1_outputs(3929) <= b and not a;
    layer1_outputs(3930) <= not b or a;
    layer1_outputs(3931) <= not (a or b);
    layer1_outputs(3932) <= not (a or b);
    layer1_outputs(3933) <= b and not a;
    layer1_outputs(3934) <= not (a and b);
    layer1_outputs(3935) <= a and b;
    layer1_outputs(3936) <= not a or b;
    layer1_outputs(3937) <= not (a and b);
    layer1_outputs(3938) <= not (a and b);
    layer1_outputs(3939) <= not (a xor b);
    layer1_outputs(3940) <= b;
    layer1_outputs(3941) <= not b;
    layer1_outputs(3942) <= b;
    layer1_outputs(3943) <= a;
    layer1_outputs(3944) <= a and not b;
    layer1_outputs(3945) <= not (a xor b);
    layer1_outputs(3946) <= b;
    layer1_outputs(3947) <= a and not b;
    layer1_outputs(3948) <= not (a xor b);
    layer1_outputs(3949) <= b and not a;
    layer1_outputs(3950) <= a and not b;
    layer1_outputs(3951) <= a xor b;
    layer1_outputs(3952) <= a and b;
    layer1_outputs(3953) <= not b;
    layer1_outputs(3954) <= not b or a;
    layer1_outputs(3955) <= not (a xor b);
    layer1_outputs(3956) <= a;
    layer1_outputs(3957) <= a and b;
    layer1_outputs(3958) <= a or b;
    layer1_outputs(3959) <= not (a xor b);
    layer1_outputs(3960) <= a xor b;
    layer1_outputs(3961) <= a and b;
    layer1_outputs(3962) <= a or b;
    layer1_outputs(3963) <= not b or a;
    layer1_outputs(3964) <= b;
    layer1_outputs(3965) <= a or b;
    layer1_outputs(3966) <= not (a xor b);
    layer1_outputs(3967) <= not b or a;
    layer1_outputs(3968) <= a or b;
    layer1_outputs(3969) <= not b or a;
    layer1_outputs(3970) <= a and b;
    layer1_outputs(3971) <= not b;
    layer1_outputs(3972) <= b;
    layer1_outputs(3973) <= not b or a;
    layer1_outputs(3974) <= a and not b;
    layer1_outputs(3975) <= b;
    layer1_outputs(3976) <= not (a and b);
    layer1_outputs(3977) <= a;
    layer1_outputs(3978) <= not (a and b);
    layer1_outputs(3979) <= a xor b;
    layer1_outputs(3980) <= b;
    layer1_outputs(3981) <= a and b;
    layer1_outputs(3982) <= not a or b;
    layer1_outputs(3983) <= not (a or b);
    layer1_outputs(3984) <= a or b;
    layer1_outputs(3985) <= not a;
    layer1_outputs(3986) <= not b or a;
    layer1_outputs(3987) <= not (a and b);
    layer1_outputs(3988) <= not b;
    layer1_outputs(3989) <= a xor b;
    layer1_outputs(3990) <= a and b;
    layer1_outputs(3991) <= not (a xor b);
    layer1_outputs(3992) <= not (a xor b);
    layer1_outputs(3993) <= not b;
    layer1_outputs(3994) <= b;
    layer1_outputs(3995) <= not (a and b);
    layer1_outputs(3996) <= a or b;
    layer1_outputs(3997) <= not a;
    layer1_outputs(3998) <= not (a and b);
    layer1_outputs(3999) <= not a or b;
    layer1_outputs(4000) <= not b;
    layer1_outputs(4001) <= not b;
    layer1_outputs(4002) <= b;
    layer1_outputs(4003) <= not b;
    layer1_outputs(4004) <= not b or a;
    layer1_outputs(4005) <= a xor b;
    layer1_outputs(4006) <= not a;
    layer1_outputs(4007) <= b and not a;
    layer1_outputs(4008) <= not a;
    layer1_outputs(4009) <= not (a xor b);
    layer1_outputs(4010) <= 1'b0;
    layer1_outputs(4011) <= a;
    layer1_outputs(4012) <= a and not b;
    layer1_outputs(4013) <= not a;
    layer1_outputs(4014) <= not a or b;
    layer1_outputs(4015) <= a and not b;
    layer1_outputs(4016) <= not (a and b);
    layer1_outputs(4017) <= not (a xor b);
    layer1_outputs(4018) <= not (a xor b);
    layer1_outputs(4019) <= not b or a;
    layer1_outputs(4020) <= a and not b;
    layer1_outputs(4021) <= not b or a;
    layer1_outputs(4022) <= b and not a;
    layer1_outputs(4023) <= not (a or b);
    layer1_outputs(4024) <= not b or a;
    layer1_outputs(4025) <= a or b;
    layer1_outputs(4026) <= not b;
    layer1_outputs(4027) <= a or b;
    layer1_outputs(4028) <= not b;
    layer1_outputs(4029) <= b;
    layer1_outputs(4030) <= a xor b;
    layer1_outputs(4031) <= not a or b;
    layer1_outputs(4032) <= not (a or b);
    layer1_outputs(4033) <= a;
    layer1_outputs(4034) <= not a or b;
    layer1_outputs(4035) <= not a;
    layer1_outputs(4036) <= a xor b;
    layer1_outputs(4037) <= b and not a;
    layer1_outputs(4038) <= not a;
    layer1_outputs(4039) <= not b;
    layer1_outputs(4040) <= not b or a;
    layer1_outputs(4041) <= b and not a;
    layer1_outputs(4042) <= not (a and b);
    layer1_outputs(4043) <= b and not a;
    layer1_outputs(4044) <= a and not b;
    layer1_outputs(4045) <= b and not a;
    layer1_outputs(4046) <= a and not b;
    layer1_outputs(4047) <= b and not a;
    layer1_outputs(4048) <= not b or a;
    layer1_outputs(4049) <= a xor b;
    layer1_outputs(4050) <= not (a and b);
    layer1_outputs(4051) <= not (a or b);
    layer1_outputs(4052) <= not (a or b);
    layer1_outputs(4053) <= a;
    layer1_outputs(4054) <= a and not b;
    layer1_outputs(4055) <= not b or a;
    layer1_outputs(4056) <= a;
    layer1_outputs(4057) <= a xor b;
    layer1_outputs(4058) <= a;
    layer1_outputs(4059) <= not a;
    layer1_outputs(4060) <= not (a xor b);
    layer1_outputs(4061) <= not b or a;
    layer1_outputs(4062) <= a xor b;
    layer1_outputs(4063) <= a;
    layer1_outputs(4064) <= b and not a;
    layer1_outputs(4065) <= not a or b;
    layer1_outputs(4066) <= a and b;
    layer1_outputs(4067) <= a or b;
    layer1_outputs(4068) <= not (a or b);
    layer1_outputs(4069) <= not (a and b);
    layer1_outputs(4070) <= not (a or b);
    layer1_outputs(4071) <= b;
    layer1_outputs(4072) <= not (a xor b);
    layer1_outputs(4073) <= a and not b;
    layer1_outputs(4074) <= not a or b;
    layer1_outputs(4075) <= a and not b;
    layer1_outputs(4076) <= a xor b;
    layer1_outputs(4077) <= not a or b;
    layer1_outputs(4078) <= not a;
    layer1_outputs(4079) <= not (a or b);
    layer1_outputs(4080) <= not b;
    layer1_outputs(4081) <= a;
    layer1_outputs(4082) <= a and b;
    layer1_outputs(4083) <= not a;
    layer1_outputs(4084) <= not (a xor b);
    layer1_outputs(4085) <= not a;
    layer1_outputs(4086) <= b;
    layer1_outputs(4087) <= not a or b;
    layer1_outputs(4088) <= not (a and b);
    layer1_outputs(4089) <= not a;
    layer1_outputs(4090) <= not b;
    layer1_outputs(4091) <= not a or b;
    layer1_outputs(4092) <= not a or b;
    layer1_outputs(4093) <= a or b;
    layer1_outputs(4094) <= not (a xor b);
    layer1_outputs(4095) <= a xor b;
    layer1_outputs(4096) <= b and not a;
    layer1_outputs(4097) <= b;
    layer1_outputs(4098) <= b;
    layer1_outputs(4099) <= a xor b;
    layer1_outputs(4100) <= a and not b;
    layer1_outputs(4101) <= not a;
    layer1_outputs(4102) <= a xor b;
    layer1_outputs(4103) <= a and not b;
    layer1_outputs(4104) <= a;
    layer1_outputs(4105) <= not a or b;
    layer1_outputs(4106) <= not (a or b);
    layer1_outputs(4107) <= a xor b;
    layer1_outputs(4108) <= not b or a;
    layer1_outputs(4109) <= a or b;
    layer1_outputs(4110) <= not a or b;
    layer1_outputs(4111) <= not (a or b);
    layer1_outputs(4112) <= a;
    layer1_outputs(4113) <= a;
    layer1_outputs(4114) <= a;
    layer1_outputs(4115) <= b;
    layer1_outputs(4116) <= not b or a;
    layer1_outputs(4117) <= a xor b;
    layer1_outputs(4118) <= a xor b;
    layer1_outputs(4119) <= not b or a;
    layer1_outputs(4120) <= a xor b;
    layer1_outputs(4121) <= a and not b;
    layer1_outputs(4122) <= a;
    layer1_outputs(4123) <= not b or a;
    layer1_outputs(4124) <= not b or a;
    layer1_outputs(4125) <= not (a or b);
    layer1_outputs(4126) <= a and b;
    layer1_outputs(4127) <= not b or a;
    layer1_outputs(4128) <= b and not a;
    layer1_outputs(4129) <= a xor b;
    layer1_outputs(4130) <= not (a or b);
    layer1_outputs(4131) <= not a or b;
    layer1_outputs(4132) <= a and b;
    layer1_outputs(4133) <= not (a xor b);
    layer1_outputs(4134) <= a xor b;
    layer1_outputs(4135) <= a and b;
    layer1_outputs(4136) <= b and not a;
    layer1_outputs(4137) <= a xor b;
    layer1_outputs(4138) <= a or b;
    layer1_outputs(4139) <= a;
    layer1_outputs(4140) <= not b or a;
    layer1_outputs(4141) <= b;
    layer1_outputs(4142) <= not b;
    layer1_outputs(4143) <= a and not b;
    layer1_outputs(4144) <= b and not a;
    layer1_outputs(4145) <= a;
    layer1_outputs(4146) <= b;
    layer1_outputs(4147) <= 1'b0;
    layer1_outputs(4148) <= a xor b;
    layer1_outputs(4149) <= not a;
    layer1_outputs(4150) <= b and not a;
    layer1_outputs(4151) <= not b;
    layer1_outputs(4152) <= a xor b;
    layer1_outputs(4153) <= b and not a;
    layer1_outputs(4154) <= b;
    layer1_outputs(4155) <= not b or a;
    layer1_outputs(4156) <= not (a and b);
    layer1_outputs(4157) <= not b;
    layer1_outputs(4158) <= b;
    layer1_outputs(4159) <= a or b;
    layer1_outputs(4160) <= not b;
    layer1_outputs(4161) <= not b or a;
    layer1_outputs(4162) <= a and not b;
    layer1_outputs(4163) <= not (a xor b);
    layer1_outputs(4164) <= b;
    layer1_outputs(4165) <= not (a or b);
    layer1_outputs(4166) <= not b or a;
    layer1_outputs(4167) <= b and not a;
    layer1_outputs(4168) <= a xor b;
    layer1_outputs(4169) <= not b;
    layer1_outputs(4170) <= not a;
    layer1_outputs(4171) <= not (a or b);
    layer1_outputs(4172) <= b;
    layer1_outputs(4173) <= not a;
    layer1_outputs(4174) <= a;
    layer1_outputs(4175) <= a;
    layer1_outputs(4176) <= not b;
    layer1_outputs(4177) <= a or b;
    layer1_outputs(4178) <= not a or b;
    layer1_outputs(4179) <= not (a xor b);
    layer1_outputs(4180) <= not (a xor b);
    layer1_outputs(4181) <= 1'b0;
    layer1_outputs(4182) <= a xor b;
    layer1_outputs(4183) <= b;
    layer1_outputs(4184) <= not b or a;
    layer1_outputs(4185) <= not (a and b);
    layer1_outputs(4186) <= a xor b;
    layer1_outputs(4187) <= a or b;
    layer1_outputs(4188) <= a and b;
    layer1_outputs(4189) <= a and b;
    layer1_outputs(4190) <= not a;
    layer1_outputs(4191) <= not (a and b);
    layer1_outputs(4192) <= not b;
    layer1_outputs(4193) <= not (a and b);
    layer1_outputs(4194) <= b and not a;
    layer1_outputs(4195) <= not a;
    layer1_outputs(4196) <= not (a or b);
    layer1_outputs(4197) <= not (a or b);
    layer1_outputs(4198) <= a and b;
    layer1_outputs(4199) <= a and not b;
    layer1_outputs(4200) <= a or b;
    layer1_outputs(4201) <= a and not b;
    layer1_outputs(4202) <= not b;
    layer1_outputs(4203) <= a;
    layer1_outputs(4204) <= not b;
    layer1_outputs(4205) <= a;
    layer1_outputs(4206) <= not b or a;
    layer1_outputs(4207) <= not a;
    layer1_outputs(4208) <= a xor b;
    layer1_outputs(4209) <= not a;
    layer1_outputs(4210) <= a and b;
    layer1_outputs(4211) <= not b;
    layer1_outputs(4212) <= not (a and b);
    layer1_outputs(4213) <= not (a and b);
    layer1_outputs(4214) <= not a;
    layer1_outputs(4215) <= not b or a;
    layer1_outputs(4216) <= not a;
    layer1_outputs(4217) <= not (a xor b);
    layer1_outputs(4218) <= a or b;
    layer1_outputs(4219) <= a;
    layer1_outputs(4220) <= not (a xor b);
    layer1_outputs(4221) <= not b;
    layer1_outputs(4222) <= not (a or b);
    layer1_outputs(4223) <= not a;
    layer1_outputs(4224) <= not a or b;
    layer1_outputs(4225) <= not (a and b);
    layer1_outputs(4226) <= a;
    layer1_outputs(4227) <= not (a and b);
    layer1_outputs(4228) <= not b;
    layer1_outputs(4229) <= a xor b;
    layer1_outputs(4230) <= not b;
    layer1_outputs(4231) <= b;
    layer1_outputs(4232) <= not (a xor b);
    layer1_outputs(4233) <= b;
    layer1_outputs(4234) <= a or b;
    layer1_outputs(4235) <= b and not a;
    layer1_outputs(4236) <= a or b;
    layer1_outputs(4237) <= b and not a;
    layer1_outputs(4238) <= a or b;
    layer1_outputs(4239) <= 1'b0;
    layer1_outputs(4240) <= not (a xor b);
    layer1_outputs(4241) <= not b;
    layer1_outputs(4242) <= not (a or b);
    layer1_outputs(4243) <= not b;
    layer1_outputs(4244) <= not b;
    layer1_outputs(4245) <= b;
    layer1_outputs(4246) <= not (a or b);
    layer1_outputs(4247) <= not b or a;
    layer1_outputs(4248) <= not (a xor b);
    layer1_outputs(4249) <= not b;
    layer1_outputs(4250) <= 1'b1;
    layer1_outputs(4251) <= a xor b;
    layer1_outputs(4252) <= a xor b;
    layer1_outputs(4253) <= not b or a;
    layer1_outputs(4254) <= not a;
    layer1_outputs(4255) <= a and not b;
    layer1_outputs(4256) <= a and not b;
    layer1_outputs(4257) <= b;
    layer1_outputs(4258) <= a and b;
    layer1_outputs(4259) <= b;
    layer1_outputs(4260) <= b and not a;
    layer1_outputs(4261) <= b and not a;
    layer1_outputs(4262) <= not b or a;
    layer1_outputs(4263) <= b and not a;
    layer1_outputs(4264) <= not (a xor b);
    layer1_outputs(4265) <= b;
    layer1_outputs(4266) <= not (a xor b);
    layer1_outputs(4267) <= a xor b;
    layer1_outputs(4268) <= a;
    layer1_outputs(4269) <= a or b;
    layer1_outputs(4270) <= a;
    layer1_outputs(4271) <= b and not a;
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= a or b;
    layer1_outputs(4274) <= not b;
    layer1_outputs(4275) <= not b or a;
    layer1_outputs(4276) <= not a;
    layer1_outputs(4277) <= not (a or b);
    layer1_outputs(4278) <= 1'b1;
    layer1_outputs(4279) <= a or b;
    layer1_outputs(4280) <= a;
    layer1_outputs(4281) <= b;
    layer1_outputs(4282) <= not (a or b);
    layer1_outputs(4283) <= a xor b;
    layer1_outputs(4284) <= not a;
    layer1_outputs(4285) <= b;
    layer1_outputs(4286) <= not b;
    layer1_outputs(4287) <= not (a xor b);
    layer1_outputs(4288) <= a and not b;
    layer1_outputs(4289) <= not (a xor b);
    layer1_outputs(4290) <= a xor b;
    layer1_outputs(4291) <= not b;
    layer1_outputs(4292) <= not b or a;
    layer1_outputs(4293) <= b and not a;
    layer1_outputs(4294) <= b;
    layer1_outputs(4295) <= b;
    layer1_outputs(4296) <= a xor b;
    layer1_outputs(4297) <= a or b;
    layer1_outputs(4298) <= not (a and b);
    layer1_outputs(4299) <= a xor b;
    layer1_outputs(4300) <= not a;
    layer1_outputs(4301) <= a and b;
    layer1_outputs(4302) <= not (a xor b);
    layer1_outputs(4303) <= a and not b;
    layer1_outputs(4304) <= not (a xor b);
    layer1_outputs(4305) <= not b or a;
    layer1_outputs(4306) <= not (a xor b);
    layer1_outputs(4307) <= not a or b;
    layer1_outputs(4308) <= not b;
    layer1_outputs(4309) <= not (a and b);
    layer1_outputs(4310) <= not b;
    layer1_outputs(4311) <= not (a and b);
    layer1_outputs(4312) <= a and not b;
    layer1_outputs(4313) <= not (a xor b);
    layer1_outputs(4314) <= not a or b;
    layer1_outputs(4315) <= not a;
    layer1_outputs(4316) <= not a or b;
    layer1_outputs(4317) <= not (a xor b);
    layer1_outputs(4318) <= not (a and b);
    layer1_outputs(4319) <= b;
    layer1_outputs(4320) <= not (a xor b);
    layer1_outputs(4321) <= a and not b;
    layer1_outputs(4322) <= b and not a;
    layer1_outputs(4323) <= b and not a;
    layer1_outputs(4324) <= a;
    layer1_outputs(4325) <= a;
    layer1_outputs(4326) <= a or b;
    layer1_outputs(4327) <= not (a or b);
    layer1_outputs(4328) <= b and not a;
    layer1_outputs(4329) <= a and b;
    layer1_outputs(4330) <= a or b;
    layer1_outputs(4331) <= not (a and b);
    layer1_outputs(4332) <= a or b;
    layer1_outputs(4333) <= not (a xor b);
    layer1_outputs(4334) <= not b;
    layer1_outputs(4335) <= b;
    layer1_outputs(4336) <= a and not b;
    layer1_outputs(4337) <= not b;
    layer1_outputs(4338) <= not (a xor b);
    layer1_outputs(4339) <= not b;
    layer1_outputs(4340) <= a;
    layer1_outputs(4341) <= not (a and b);
    layer1_outputs(4342) <= not b;
    layer1_outputs(4343) <= not a;
    layer1_outputs(4344) <= not (a or b);
    layer1_outputs(4345) <= a xor b;
    layer1_outputs(4346) <= a xor b;
    layer1_outputs(4347) <= a or b;
    layer1_outputs(4348) <= a and not b;
    layer1_outputs(4349) <= a;
    layer1_outputs(4350) <= a and not b;
    layer1_outputs(4351) <= not b;
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= a;
    layer1_outputs(4354) <= b;
    layer1_outputs(4355) <= b;
    layer1_outputs(4356) <= a xor b;
    layer1_outputs(4357) <= not (a or b);
    layer1_outputs(4358) <= b and not a;
    layer1_outputs(4359) <= a xor b;
    layer1_outputs(4360) <= not b;
    layer1_outputs(4361) <= not b;
    layer1_outputs(4362) <= not b;
    layer1_outputs(4363) <= a xor b;
    layer1_outputs(4364) <= b;
    layer1_outputs(4365) <= not (a xor b);
    layer1_outputs(4366) <= not b or a;
    layer1_outputs(4367) <= b and not a;
    layer1_outputs(4368) <= b and not a;
    layer1_outputs(4369) <= a;
    layer1_outputs(4370) <= a xor b;
    layer1_outputs(4371) <= a xor b;
    layer1_outputs(4372) <= not b;
    layer1_outputs(4373) <= a or b;
    layer1_outputs(4374) <= not (a and b);
    layer1_outputs(4375) <= 1'b1;
    layer1_outputs(4376) <= 1'b0;
    layer1_outputs(4377) <= not a or b;
    layer1_outputs(4378) <= not b or a;
    layer1_outputs(4379) <= b;
    layer1_outputs(4380) <= b and not a;
    layer1_outputs(4381) <= a or b;
    layer1_outputs(4382) <= b and not a;
    layer1_outputs(4383) <= not (a xor b);
    layer1_outputs(4384) <= a and b;
    layer1_outputs(4385) <= not (a and b);
    layer1_outputs(4386) <= b;
    layer1_outputs(4387) <= b;
    layer1_outputs(4388) <= not (a and b);
    layer1_outputs(4389) <= a;
    layer1_outputs(4390) <= 1'b1;
    layer1_outputs(4391) <= not a;
    layer1_outputs(4392) <= not (a and b);
    layer1_outputs(4393) <= b and not a;
    layer1_outputs(4394) <= b;
    layer1_outputs(4395) <= b;
    layer1_outputs(4396) <= a or b;
    layer1_outputs(4397) <= a and not b;
    layer1_outputs(4398) <= b and not a;
    layer1_outputs(4399) <= not a;
    layer1_outputs(4400) <= not a;
    layer1_outputs(4401) <= a or b;
    layer1_outputs(4402) <= not a or b;
    layer1_outputs(4403) <= not b or a;
    layer1_outputs(4404) <= not a;
    layer1_outputs(4405) <= b;
    layer1_outputs(4406) <= a;
    layer1_outputs(4407) <= not b or a;
    layer1_outputs(4408) <= not (a or b);
    layer1_outputs(4409) <= a and b;
    layer1_outputs(4410) <= a and b;
    layer1_outputs(4411) <= a and not b;
    layer1_outputs(4412) <= a xor b;
    layer1_outputs(4413) <= not b;
    layer1_outputs(4414) <= not (a and b);
    layer1_outputs(4415) <= a and b;
    layer1_outputs(4416) <= b;
    layer1_outputs(4417) <= a or b;
    layer1_outputs(4418) <= 1'b1;
    layer1_outputs(4419) <= not a or b;
    layer1_outputs(4420) <= not b;
    layer1_outputs(4421) <= a xor b;
    layer1_outputs(4422) <= b and not a;
    layer1_outputs(4423) <= not a;
    layer1_outputs(4424) <= not b;
    layer1_outputs(4425) <= a and b;
    layer1_outputs(4426) <= a and not b;
    layer1_outputs(4427) <= a;
    layer1_outputs(4428) <= not (a and b);
    layer1_outputs(4429) <= b and not a;
    layer1_outputs(4430) <= not b;
    layer1_outputs(4431) <= a and not b;
    layer1_outputs(4432) <= 1'b1;
    layer1_outputs(4433) <= not a or b;
    layer1_outputs(4434) <= not a or b;
    layer1_outputs(4435) <= not (a and b);
    layer1_outputs(4436) <= a;
    layer1_outputs(4437) <= a or b;
    layer1_outputs(4438) <= not (a xor b);
    layer1_outputs(4439) <= not (a xor b);
    layer1_outputs(4440) <= b;
    layer1_outputs(4441) <= b;
    layer1_outputs(4442) <= a and not b;
    layer1_outputs(4443) <= a xor b;
    layer1_outputs(4444) <= not (a and b);
    layer1_outputs(4445) <= b;
    layer1_outputs(4446) <= not (a or b);
    layer1_outputs(4447) <= a and not b;
    layer1_outputs(4448) <= not (a or b);
    layer1_outputs(4449) <= a or b;
    layer1_outputs(4450) <= not a;
    layer1_outputs(4451) <= not (a and b);
    layer1_outputs(4452) <= a xor b;
    layer1_outputs(4453) <= a and b;
    layer1_outputs(4454) <= not a;
    layer1_outputs(4455) <= a or b;
    layer1_outputs(4456) <= not (a xor b);
    layer1_outputs(4457) <= not (a or b);
    layer1_outputs(4458) <= a and not b;
    layer1_outputs(4459) <= b and not a;
    layer1_outputs(4460) <= b and not a;
    layer1_outputs(4461) <= not a or b;
    layer1_outputs(4462) <= b;
    layer1_outputs(4463) <= not (a or b);
    layer1_outputs(4464) <= not b;
    layer1_outputs(4465) <= not (a xor b);
    layer1_outputs(4466) <= a xor b;
    layer1_outputs(4467) <= not a;
    layer1_outputs(4468) <= not (a and b);
    layer1_outputs(4469) <= a;
    layer1_outputs(4470) <= not a or b;
    layer1_outputs(4471) <= not a or b;
    layer1_outputs(4472) <= a and b;
    layer1_outputs(4473) <= b;
    layer1_outputs(4474) <= not b;
    layer1_outputs(4475) <= a or b;
    layer1_outputs(4476) <= not b;
    layer1_outputs(4477) <= a and not b;
    layer1_outputs(4478) <= not b or a;
    layer1_outputs(4479) <= a xor b;
    layer1_outputs(4480) <= not b or a;
    layer1_outputs(4481) <= a xor b;
    layer1_outputs(4482) <= a;
    layer1_outputs(4483) <= not b;
    layer1_outputs(4484) <= a or b;
    layer1_outputs(4485) <= not (a xor b);
    layer1_outputs(4486) <= a xor b;
    layer1_outputs(4487) <= not a or b;
    layer1_outputs(4488) <= not (a xor b);
    layer1_outputs(4489) <= a;
    layer1_outputs(4490) <= a and b;
    layer1_outputs(4491) <= a and b;
    layer1_outputs(4492) <= b;
    layer1_outputs(4493) <= 1'b0;
    layer1_outputs(4494) <= a or b;
    layer1_outputs(4495) <= not b or a;
    layer1_outputs(4496) <= a and b;
    layer1_outputs(4497) <= not b;
    layer1_outputs(4498) <= a;
    layer1_outputs(4499) <= a or b;
    layer1_outputs(4500) <= not b;
    layer1_outputs(4501) <= not b or a;
    layer1_outputs(4502) <= not a;
    layer1_outputs(4503) <= a;
    layer1_outputs(4504) <= not (a or b);
    layer1_outputs(4505) <= a;
    layer1_outputs(4506) <= not (a or b);
    layer1_outputs(4507) <= not a or b;
    layer1_outputs(4508) <= not (a xor b);
    layer1_outputs(4509) <= b and not a;
    layer1_outputs(4510) <= 1'b0;
    layer1_outputs(4511) <= a;
    layer1_outputs(4512) <= not (a and b);
    layer1_outputs(4513) <= a and b;
    layer1_outputs(4514) <= b;
    layer1_outputs(4515) <= a and not b;
    layer1_outputs(4516) <= a xor b;
    layer1_outputs(4517) <= a;
    layer1_outputs(4518) <= a and b;
    layer1_outputs(4519) <= a and not b;
    layer1_outputs(4520) <= a and b;
    layer1_outputs(4521) <= not a;
    layer1_outputs(4522) <= not a;
    layer1_outputs(4523) <= a and b;
    layer1_outputs(4524) <= a;
    layer1_outputs(4525) <= not (a or b);
    layer1_outputs(4526) <= a and b;
    layer1_outputs(4527) <= not b or a;
    layer1_outputs(4528) <= not b;
    layer1_outputs(4529) <= not (a xor b);
    layer1_outputs(4530) <= a and not b;
    layer1_outputs(4531) <= b and not a;
    layer1_outputs(4532) <= not b;
    layer1_outputs(4533) <= not b;
    layer1_outputs(4534) <= a xor b;
    layer1_outputs(4535) <= not b or a;
    layer1_outputs(4536) <= b and not a;
    layer1_outputs(4537) <= not (a and b);
    layer1_outputs(4538) <= not a or b;
    layer1_outputs(4539) <= b;
    layer1_outputs(4540) <= a;
    layer1_outputs(4541) <= not (a xor b);
    layer1_outputs(4542) <= not a;
    layer1_outputs(4543) <= not b;
    layer1_outputs(4544) <= not (a or b);
    layer1_outputs(4545) <= not a or b;
    layer1_outputs(4546) <= b;
    layer1_outputs(4547) <= b;
    layer1_outputs(4548) <= not (a xor b);
    layer1_outputs(4549) <= not a;
    layer1_outputs(4550) <= not a or b;
    layer1_outputs(4551) <= not (a or b);
    layer1_outputs(4552) <= not (a and b);
    layer1_outputs(4553) <= not b or a;
    layer1_outputs(4554) <= not b;
    layer1_outputs(4555) <= not b or a;
    layer1_outputs(4556) <= a and b;
    layer1_outputs(4557) <= a;
    layer1_outputs(4558) <= a and b;
    layer1_outputs(4559) <= not (a xor b);
    layer1_outputs(4560) <= b;
    layer1_outputs(4561) <= a xor b;
    layer1_outputs(4562) <= not (a and b);
    layer1_outputs(4563) <= a or b;
    layer1_outputs(4564) <= 1'b1;
    layer1_outputs(4565) <= not (a xor b);
    layer1_outputs(4566) <= b and not a;
    layer1_outputs(4567) <= not b or a;
    layer1_outputs(4568) <= a or b;
    layer1_outputs(4569) <= not a;
    layer1_outputs(4570) <= b;
    layer1_outputs(4571) <= b and not a;
    layer1_outputs(4572) <= not b or a;
    layer1_outputs(4573) <= not (a and b);
    layer1_outputs(4574) <= b;
    layer1_outputs(4575) <= a and b;
    layer1_outputs(4576) <= not (a and b);
    layer1_outputs(4577) <= not (a and b);
    layer1_outputs(4578) <= not (a and b);
    layer1_outputs(4579) <= not (a xor b);
    layer1_outputs(4580) <= not (a xor b);
    layer1_outputs(4581) <= not a;
    layer1_outputs(4582) <= not (a or b);
    layer1_outputs(4583) <= a and b;
    layer1_outputs(4584) <= not a;
    layer1_outputs(4585) <= not b or a;
    layer1_outputs(4586) <= not a;
    layer1_outputs(4587) <= not (a xor b);
    layer1_outputs(4588) <= b;
    layer1_outputs(4589) <= not (a and b);
    layer1_outputs(4590) <= not b;
    layer1_outputs(4591) <= not (a or b);
    layer1_outputs(4592) <= not b;
    layer1_outputs(4593) <= a or b;
    layer1_outputs(4594) <= b;
    layer1_outputs(4595) <= a;
    layer1_outputs(4596) <= not a;
    layer1_outputs(4597) <= not b;
    layer1_outputs(4598) <= a;
    layer1_outputs(4599) <= not (a xor b);
    layer1_outputs(4600) <= not (a or b);
    layer1_outputs(4601) <= a or b;
    layer1_outputs(4602) <= not a;
    layer1_outputs(4603) <= a;
    layer1_outputs(4604) <= not (a or b);
    layer1_outputs(4605) <= a and not b;
    layer1_outputs(4606) <= b;
    layer1_outputs(4607) <= not (a xor b);
    layer1_outputs(4608) <= not (a xor b);
    layer1_outputs(4609) <= not b;
    layer1_outputs(4610) <= a;
    layer1_outputs(4611) <= a and not b;
    layer1_outputs(4612) <= a xor b;
    layer1_outputs(4613) <= not b or a;
    layer1_outputs(4614) <= not (a and b);
    layer1_outputs(4615) <= b and not a;
    layer1_outputs(4616) <= a and not b;
    layer1_outputs(4617) <= not a;
    layer1_outputs(4618) <= not (a xor b);
    layer1_outputs(4619) <= a or b;
    layer1_outputs(4620) <= not (a and b);
    layer1_outputs(4621) <= a xor b;
    layer1_outputs(4622) <= not a or b;
    layer1_outputs(4623) <= not a;
    layer1_outputs(4624) <= not a or b;
    layer1_outputs(4625) <= b;
    layer1_outputs(4626) <= not (a or b);
    layer1_outputs(4627) <= a and b;
    layer1_outputs(4628) <= b;
    layer1_outputs(4629) <= not b;
    layer1_outputs(4630) <= not (a and b);
    layer1_outputs(4631) <= b;
    layer1_outputs(4632) <= b and not a;
    layer1_outputs(4633) <= not b;
    layer1_outputs(4634) <= not b or a;
    layer1_outputs(4635) <= a and not b;
    layer1_outputs(4636) <= not (a xor b);
    layer1_outputs(4637) <= a and b;
    layer1_outputs(4638) <= a and not b;
    layer1_outputs(4639) <= not a;
    layer1_outputs(4640) <= a xor b;
    layer1_outputs(4641) <= a;
    layer1_outputs(4642) <= a xor b;
    layer1_outputs(4643) <= not a;
    layer1_outputs(4644) <= a xor b;
    layer1_outputs(4645) <= a and not b;
    layer1_outputs(4646) <= not (a and b);
    layer1_outputs(4647) <= a;
    layer1_outputs(4648) <= not (a or b);
    layer1_outputs(4649) <= a and b;
    layer1_outputs(4650) <= a;
    layer1_outputs(4651) <= a and b;
    layer1_outputs(4652) <= not b;
    layer1_outputs(4653) <= b;
    layer1_outputs(4654) <= a;
    layer1_outputs(4655) <= not a;
    layer1_outputs(4656) <= not b;
    layer1_outputs(4657) <= not (a and b);
    layer1_outputs(4658) <= not b;
    layer1_outputs(4659) <= a or b;
    layer1_outputs(4660) <= a and b;
    layer1_outputs(4661) <= a xor b;
    layer1_outputs(4662) <= not b or a;
    layer1_outputs(4663) <= not (a xor b);
    layer1_outputs(4664) <= not (a or b);
    layer1_outputs(4665) <= b;
    layer1_outputs(4666) <= not b;
    layer1_outputs(4667) <= a;
    layer1_outputs(4668) <= not (a and b);
    layer1_outputs(4669) <= not a;
    layer1_outputs(4670) <= a xor b;
    layer1_outputs(4671) <= b and not a;
    layer1_outputs(4672) <= b and not a;
    layer1_outputs(4673) <= a xor b;
    layer1_outputs(4674) <= a xor b;
    layer1_outputs(4675) <= not b;
    layer1_outputs(4676) <= a xor b;
    layer1_outputs(4677) <= not b or a;
    layer1_outputs(4678) <= a or b;
    layer1_outputs(4679) <= a or b;
    layer1_outputs(4680) <= not b;
    layer1_outputs(4681) <= not a;
    layer1_outputs(4682) <= not (a or b);
    layer1_outputs(4683) <= a and b;
    layer1_outputs(4684) <= a;
    layer1_outputs(4685) <= not a;
    layer1_outputs(4686) <= not b;
    layer1_outputs(4687) <= not b;
    layer1_outputs(4688) <= not a or b;
    layer1_outputs(4689) <= a and not b;
    layer1_outputs(4690) <= b;
    layer1_outputs(4691) <= not (a or b);
    layer1_outputs(4692) <= a;
    layer1_outputs(4693) <= b;
    layer1_outputs(4694) <= not a or b;
    layer1_outputs(4695) <= a;
    layer1_outputs(4696) <= a;
    layer1_outputs(4697) <= a or b;
    layer1_outputs(4698) <= not (a or b);
    layer1_outputs(4699) <= a and b;
    layer1_outputs(4700) <= not a or b;
    layer1_outputs(4701) <= not (a xor b);
    layer1_outputs(4702) <= not b;
    layer1_outputs(4703) <= a and b;
    layer1_outputs(4704) <= a and not b;
    layer1_outputs(4705) <= b and not a;
    layer1_outputs(4706) <= not a or b;
    layer1_outputs(4707) <= b;
    layer1_outputs(4708) <= not b or a;
    layer1_outputs(4709) <= not (a and b);
    layer1_outputs(4710) <= a or b;
    layer1_outputs(4711) <= b;
    layer1_outputs(4712) <= a xor b;
    layer1_outputs(4713) <= not a;
    layer1_outputs(4714) <= a and b;
    layer1_outputs(4715) <= not b;
    layer1_outputs(4716) <= not (a or b);
    layer1_outputs(4717) <= not b;
    layer1_outputs(4718) <= a and b;
    layer1_outputs(4719) <= 1'b0;
    layer1_outputs(4720) <= not a;
    layer1_outputs(4721) <= not (a and b);
    layer1_outputs(4722) <= a or b;
    layer1_outputs(4723) <= not (a xor b);
    layer1_outputs(4724) <= not (a and b);
    layer1_outputs(4725) <= a;
    layer1_outputs(4726) <= a or b;
    layer1_outputs(4727) <= b;
    layer1_outputs(4728) <= not a or b;
    layer1_outputs(4729) <= a or b;
    layer1_outputs(4730) <= a and not b;
    layer1_outputs(4731) <= a xor b;
    layer1_outputs(4732) <= not b;
    layer1_outputs(4733) <= a;
    layer1_outputs(4734) <= a xor b;
    layer1_outputs(4735) <= b;
    layer1_outputs(4736) <= b and not a;
    layer1_outputs(4737) <= not a or b;
    layer1_outputs(4738) <= not a;
    layer1_outputs(4739) <= not (a and b);
    layer1_outputs(4740) <= a;
    layer1_outputs(4741) <= a xor b;
    layer1_outputs(4742) <= b;
    layer1_outputs(4743) <= not b or a;
    layer1_outputs(4744) <= not (a xor b);
    layer1_outputs(4745) <= a xor b;
    layer1_outputs(4746) <= a;
    layer1_outputs(4747) <= a xor b;
    layer1_outputs(4748) <= b and not a;
    layer1_outputs(4749) <= a xor b;
    layer1_outputs(4750) <= 1'b0;
    layer1_outputs(4751) <= not b;
    layer1_outputs(4752) <= not a or b;
    layer1_outputs(4753) <= a;
    layer1_outputs(4754) <= b and not a;
    layer1_outputs(4755) <= not b or a;
    layer1_outputs(4756) <= not b;
    layer1_outputs(4757) <= not b;
    layer1_outputs(4758) <= not a;
    layer1_outputs(4759) <= not a or b;
    layer1_outputs(4760) <= not (a xor b);
    layer1_outputs(4761) <= not a or b;
    layer1_outputs(4762) <= a and b;
    layer1_outputs(4763) <= a and not b;
    layer1_outputs(4764) <= not b or a;
    layer1_outputs(4765) <= b;
    layer1_outputs(4766) <= a xor b;
    layer1_outputs(4767) <= a and b;
    layer1_outputs(4768) <= not (a and b);
    layer1_outputs(4769) <= not a;
    layer1_outputs(4770) <= not a;
    layer1_outputs(4771) <= not b or a;
    layer1_outputs(4772) <= b;
    layer1_outputs(4773) <= a or b;
    layer1_outputs(4774) <= b;
    layer1_outputs(4775) <= a;
    layer1_outputs(4776) <= b;
    layer1_outputs(4777) <= not (a xor b);
    layer1_outputs(4778) <= b;
    layer1_outputs(4779) <= a and not b;
    layer1_outputs(4780) <= not b;
    layer1_outputs(4781) <= a;
    layer1_outputs(4782) <= b and not a;
    layer1_outputs(4783) <= not (a and b);
    layer1_outputs(4784) <= not a or b;
    layer1_outputs(4785) <= a and b;
    layer1_outputs(4786) <= not a;
    layer1_outputs(4787) <= not a;
    layer1_outputs(4788) <= a xor b;
    layer1_outputs(4789) <= not (a and b);
    layer1_outputs(4790) <= b;
    layer1_outputs(4791) <= not a;
    layer1_outputs(4792) <= not (a xor b);
    layer1_outputs(4793) <= a and b;
    layer1_outputs(4794) <= not b or a;
    layer1_outputs(4795) <= not a;
    layer1_outputs(4796) <= b and not a;
    layer1_outputs(4797) <= 1'b1;
    layer1_outputs(4798) <= not a;
    layer1_outputs(4799) <= not (a xor b);
    layer1_outputs(4800) <= not a;
    layer1_outputs(4801) <= not b or a;
    layer1_outputs(4802) <= not (a xor b);
    layer1_outputs(4803) <= a;
    layer1_outputs(4804) <= a and not b;
    layer1_outputs(4805) <= 1'b1;
    layer1_outputs(4806) <= a xor b;
    layer1_outputs(4807) <= not a or b;
    layer1_outputs(4808) <= a or b;
    layer1_outputs(4809) <= not (a xor b);
    layer1_outputs(4810) <= a and not b;
    layer1_outputs(4811) <= b;
    layer1_outputs(4812) <= not (a and b);
    layer1_outputs(4813) <= a;
    layer1_outputs(4814) <= a and b;
    layer1_outputs(4815) <= b;
    layer1_outputs(4816) <= b;
    layer1_outputs(4817) <= b;
    layer1_outputs(4818) <= a and b;
    layer1_outputs(4819) <= not b;
    layer1_outputs(4820) <= not a or b;
    layer1_outputs(4821) <= not (a or b);
    layer1_outputs(4822) <= a xor b;
    layer1_outputs(4823) <= b;
    layer1_outputs(4824) <= not (a xor b);
    layer1_outputs(4825) <= a and b;
    layer1_outputs(4826) <= not b or a;
    layer1_outputs(4827) <= not b or a;
    layer1_outputs(4828) <= a and b;
    layer1_outputs(4829) <= a xor b;
    layer1_outputs(4830) <= not (a or b);
    layer1_outputs(4831) <= b;
    layer1_outputs(4832) <= not (a xor b);
    layer1_outputs(4833) <= a and b;
    layer1_outputs(4834) <= not a;
    layer1_outputs(4835) <= not (a xor b);
    layer1_outputs(4836) <= not b;
    layer1_outputs(4837) <= not b;
    layer1_outputs(4838) <= b and not a;
    layer1_outputs(4839) <= not (a xor b);
    layer1_outputs(4840) <= a or b;
    layer1_outputs(4841) <= 1'b1;
    layer1_outputs(4842) <= a and not b;
    layer1_outputs(4843) <= not b;
    layer1_outputs(4844) <= a and b;
    layer1_outputs(4845) <= a;
    layer1_outputs(4846) <= b;
    layer1_outputs(4847) <= not (a and b);
    layer1_outputs(4848) <= a;
    layer1_outputs(4849) <= a xor b;
    layer1_outputs(4850) <= not (a xor b);
    layer1_outputs(4851) <= a xor b;
    layer1_outputs(4852) <= not b;
    layer1_outputs(4853) <= not (a xor b);
    layer1_outputs(4854) <= not (a and b);
    layer1_outputs(4855) <= a or b;
    layer1_outputs(4856) <= a or b;
    layer1_outputs(4857) <= not (a or b);
    layer1_outputs(4858) <= a or b;
    layer1_outputs(4859) <= not a;
    layer1_outputs(4860) <= not b;
    layer1_outputs(4861) <= not (a or b);
    layer1_outputs(4862) <= a;
    layer1_outputs(4863) <= a xor b;
    layer1_outputs(4864) <= not (a and b);
    layer1_outputs(4865) <= a;
    layer1_outputs(4866) <= a;
    layer1_outputs(4867) <= a xor b;
    layer1_outputs(4868) <= a or b;
    layer1_outputs(4869) <= a and b;
    layer1_outputs(4870) <= not (a xor b);
    layer1_outputs(4871) <= not a;
    layer1_outputs(4872) <= not b or a;
    layer1_outputs(4873) <= not (a and b);
    layer1_outputs(4874) <= not a or b;
    layer1_outputs(4875) <= not b;
    layer1_outputs(4876) <= a or b;
    layer1_outputs(4877) <= a and not b;
    layer1_outputs(4878) <= not b or a;
    layer1_outputs(4879) <= a;
    layer1_outputs(4880) <= a;
    layer1_outputs(4881) <= not (a or b);
    layer1_outputs(4882) <= not a;
    layer1_outputs(4883) <= not a or b;
    layer1_outputs(4884) <= not a;
    layer1_outputs(4885) <= not a;
    layer1_outputs(4886) <= not (a or b);
    layer1_outputs(4887) <= not a;
    layer1_outputs(4888) <= a or b;
    layer1_outputs(4889) <= not (a xor b);
    layer1_outputs(4890) <= not (a xor b);
    layer1_outputs(4891) <= a;
    layer1_outputs(4892) <= a xor b;
    layer1_outputs(4893) <= a xor b;
    layer1_outputs(4894) <= a and not b;
    layer1_outputs(4895) <= b and not a;
    layer1_outputs(4896) <= a or b;
    layer1_outputs(4897) <= b and not a;
    layer1_outputs(4898) <= not a;
    layer1_outputs(4899) <= not (a xor b);
    layer1_outputs(4900) <= not a;
    layer1_outputs(4901) <= not (a xor b);
    layer1_outputs(4902) <= a;
    layer1_outputs(4903) <= not (a xor b);
    layer1_outputs(4904) <= a;
    layer1_outputs(4905) <= not (a or b);
    layer1_outputs(4906) <= not (a xor b);
    layer1_outputs(4907) <= b;
    layer1_outputs(4908) <= a and not b;
    layer1_outputs(4909) <= a;
    layer1_outputs(4910) <= not b;
    layer1_outputs(4911) <= not a;
    layer1_outputs(4912) <= not a;
    layer1_outputs(4913) <= b and not a;
    layer1_outputs(4914) <= b and not a;
    layer1_outputs(4915) <= a xor b;
    layer1_outputs(4916) <= b and not a;
    layer1_outputs(4917) <= b;
    layer1_outputs(4918) <= a or b;
    layer1_outputs(4919) <= a;
    layer1_outputs(4920) <= not a;
    layer1_outputs(4921) <= b and not a;
    layer1_outputs(4922) <= b;
    layer1_outputs(4923) <= a or b;
    layer1_outputs(4924) <= not a;
    layer1_outputs(4925) <= not a;
    layer1_outputs(4926) <= b;
    layer1_outputs(4927) <= not (a xor b);
    layer1_outputs(4928) <= not (a xor b);
    layer1_outputs(4929) <= a or b;
    layer1_outputs(4930) <= b and not a;
    layer1_outputs(4931) <= a or b;
    layer1_outputs(4932) <= not (a xor b);
    layer1_outputs(4933) <= not b or a;
    layer1_outputs(4934) <= a;
    layer1_outputs(4935) <= not a or b;
    layer1_outputs(4936) <= a xor b;
    layer1_outputs(4937) <= not a or b;
    layer1_outputs(4938) <= a or b;
    layer1_outputs(4939) <= not b;
    layer1_outputs(4940) <= b and not a;
    layer1_outputs(4941) <= a;
    layer1_outputs(4942) <= b;
    layer1_outputs(4943) <= not (a xor b);
    layer1_outputs(4944) <= b;
    layer1_outputs(4945) <= not a;
    layer1_outputs(4946) <= a;
    layer1_outputs(4947) <= a;
    layer1_outputs(4948) <= not a or b;
    layer1_outputs(4949) <= not (a xor b);
    layer1_outputs(4950) <= b;
    layer1_outputs(4951) <= not b or a;
    layer1_outputs(4952) <= not a;
    layer1_outputs(4953) <= not b;
    layer1_outputs(4954) <= a and b;
    layer1_outputs(4955) <= a and b;
    layer1_outputs(4956) <= a;
    layer1_outputs(4957) <= not (a and b);
    layer1_outputs(4958) <= a and b;
    layer1_outputs(4959) <= not (a or b);
    layer1_outputs(4960) <= not (a and b);
    layer1_outputs(4961) <= not (a and b);
    layer1_outputs(4962) <= a;
    layer1_outputs(4963) <= b;
    layer1_outputs(4964) <= a and not b;
    layer1_outputs(4965) <= not b;
    layer1_outputs(4966) <= a;
    layer1_outputs(4967) <= a and not b;
    layer1_outputs(4968) <= a xor b;
    layer1_outputs(4969) <= not (a or b);
    layer1_outputs(4970) <= a or b;
    layer1_outputs(4971) <= not b;
    layer1_outputs(4972) <= a xor b;
    layer1_outputs(4973) <= not a or b;
    layer1_outputs(4974) <= b and not a;
    layer1_outputs(4975) <= a and not b;
    layer1_outputs(4976) <= b and not a;
    layer1_outputs(4977) <= a;
    layer1_outputs(4978) <= a and not b;
    layer1_outputs(4979) <= not b or a;
    layer1_outputs(4980) <= not (a or b);
    layer1_outputs(4981) <= not b;
    layer1_outputs(4982) <= not a;
    layer1_outputs(4983) <= a;
    layer1_outputs(4984) <= not (a or b);
    layer1_outputs(4985) <= not (a and b);
    layer1_outputs(4986) <= b;
    layer1_outputs(4987) <= not (a or b);
    layer1_outputs(4988) <= a and not b;
    layer1_outputs(4989) <= a and b;
    layer1_outputs(4990) <= not (a xor b);
    layer1_outputs(4991) <= not b;
    layer1_outputs(4992) <= not b;
    layer1_outputs(4993) <= a;
    layer1_outputs(4994) <= not (a xor b);
    layer1_outputs(4995) <= a;
    layer1_outputs(4996) <= a or b;
    layer1_outputs(4997) <= not b;
    layer1_outputs(4998) <= not (a xor b);
    layer1_outputs(4999) <= b;
    layer1_outputs(5000) <= not b or a;
    layer1_outputs(5001) <= b and not a;
    layer1_outputs(5002) <= not (a and b);
    layer1_outputs(5003) <= b and not a;
    layer1_outputs(5004) <= not b;
    layer1_outputs(5005) <= b and not a;
    layer1_outputs(5006) <= a xor b;
    layer1_outputs(5007) <= not (a and b);
    layer1_outputs(5008) <= b;
    layer1_outputs(5009) <= not (a and b);
    layer1_outputs(5010) <= not (a or b);
    layer1_outputs(5011) <= not (a xor b);
    layer1_outputs(5012) <= b;
    layer1_outputs(5013) <= not (a or b);
    layer1_outputs(5014) <= 1'b0;
    layer1_outputs(5015) <= a and not b;
    layer1_outputs(5016) <= 1'b1;
    layer1_outputs(5017) <= b;
    layer1_outputs(5018) <= a or b;
    layer1_outputs(5019) <= not b or a;
    layer1_outputs(5020) <= not (a or b);
    layer1_outputs(5021) <= a;
    layer1_outputs(5022) <= b and not a;
    layer1_outputs(5023) <= a or b;
    layer1_outputs(5024) <= a;
    layer1_outputs(5025) <= a xor b;
    layer1_outputs(5026) <= not b or a;
    layer1_outputs(5027) <= not b or a;
    layer1_outputs(5028) <= not b;
    layer1_outputs(5029) <= not (a and b);
    layer1_outputs(5030) <= not a or b;
    layer1_outputs(5031) <= a xor b;
    layer1_outputs(5032) <= 1'b0;
    layer1_outputs(5033) <= not b;
    layer1_outputs(5034) <= a and b;
    layer1_outputs(5035) <= a;
    layer1_outputs(5036) <= not (a or b);
    layer1_outputs(5037) <= not (a or b);
    layer1_outputs(5038) <= not a or b;
    layer1_outputs(5039) <= a and b;
    layer1_outputs(5040) <= not (a xor b);
    layer1_outputs(5041) <= a and not b;
    layer1_outputs(5042) <= not (a xor b);
    layer1_outputs(5043) <= not a;
    layer1_outputs(5044) <= not a;
    layer1_outputs(5045) <= not b or a;
    layer1_outputs(5046) <= b and not a;
    layer1_outputs(5047) <= not (a xor b);
    layer1_outputs(5048) <= a xor b;
    layer1_outputs(5049) <= not b or a;
    layer1_outputs(5050) <= not a;
    layer1_outputs(5051) <= a and b;
    layer1_outputs(5052) <= a and b;
    layer1_outputs(5053) <= not b;
    layer1_outputs(5054) <= a xor b;
    layer1_outputs(5055) <= not (a and b);
    layer1_outputs(5056) <= a xor b;
    layer1_outputs(5057) <= not a or b;
    layer1_outputs(5058) <= not a;
    layer1_outputs(5059) <= a and not b;
    layer1_outputs(5060) <= not b or a;
    layer1_outputs(5061) <= not b;
    layer1_outputs(5062) <= not b or a;
    layer1_outputs(5063) <= not a;
    layer1_outputs(5064) <= not b;
    layer1_outputs(5065) <= not (a and b);
    layer1_outputs(5066) <= not (a or b);
    layer1_outputs(5067) <= not b or a;
    layer1_outputs(5068) <= a;
    layer1_outputs(5069) <= not b or a;
    layer1_outputs(5070) <= not (a xor b);
    layer1_outputs(5071) <= a and b;
    layer1_outputs(5072) <= a;
    layer1_outputs(5073) <= not b;
    layer1_outputs(5074) <= a;
    layer1_outputs(5075) <= a xor b;
    layer1_outputs(5076) <= not a;
    layer1_outputs(5077) <= a xor b;
    layer1_outputs(5078) <= b and not a;
    layer1_outputs(5079) <= a;
    layer1_outputs(5080) <= a or b;
    layer1_outputs(5081) <= a and not b;
    layer1_outputs(5082) <= not (a xor b);
    layer1_outputs(5083) <= a;
    layer1_outputs(5084) <= a;
    layer1_outputs(5085) <= not (a or b);
    layer1_outputs(5086) <= a or b;
    layer1_outputs(5087) <= b and not a;
    layer1_outputs(5088) <= not a or b;
    layer1_outputs(5089) <= b and not a;
    layer1_outputs(5090) <= 1'b1;
    layer1_outputs(5091) <= not (a xor b);
    layer1_outputs(5092) <= b;
    layer1_outputs(5093) <= a;
    layer1_outputs(5094) <= not a or b;
    layer1_outputs(5095) <= b;
    layer1_outputs(5096) <= a xor b;
    layer1_outputs(5097) <= not a or b;
    layer1_outputs(5098) <= a;
    layer1_outputs(5099) <= a xor b;
    layer1_outputs(5100) <= not (a xor b);
    layer1_outputs(5101) <= a;
    layer1_outputs(5102) <= not (a and b);
    layer1_outputs(5103) <= a and not b;
    layer1_outputs(5104) <= not a;
    layer1_outputs(5105) <= b;
    layer1_outputs(5106) <= a;
    layer1_outputs(5107) <= not (a and b);
    layer1_outputs(5108) <= not b;
    layer1_outputs(5109) <= not b;
    layer1_outputs(5110) <= not b;
    layer1_outputs(5111) <= a xor b;
    layer1_outputs(5112) <= not a or b;
    layer1_outputs(5113) <= a and not b;
    layer1_outputs(5114) <= a and b;
    layer1_outputs(5115) <= not (a and b);
    layer1_outputs(5116) <= b;
    layer1_outputs(5117) <= a or b;
    layer1_outputs(5118) <= not (a xor b);
    layer1_outputs(5119) <= not (a xor b);
    layer1_outputs(5120) <= a xor b;
    layer1_outputs(5121) <= a or b;
    layer1_outputs(5122) <= a xor b;
    layer1_outputs(5123) <= not a or b;
    layer1_outputs(5124) <= not b or a;
    layer1_outputs(5125) <= a or b;
    layer1_outputs(5126) <= b;
    layer1_outputs(5127) <= not (a xor b);
    layer1_outputs(5128) <= not (a and b);
    layer1_outputs(5129) <= not a;
    layer1_outputs(5130) <= a;
    layer1_outputs(5131) <= not a;
    layer1_outputs(5132) <= not a or b;
    layer1_outputs(5133) <= not b;
    layer1_outputs(5134) <= a xor b;
    layer1_outputs(5135) <= b;
    layer1_outputs(5136) <= 1'b1;
    layer1_outputs(5137) <= not a;
    layer1_outputs(5138) <= a xor b;
    layer1_outputs(5139) <= a or b;
    layer1_outputs(5140) <= not b or a;
    layer1_outputs(5141) <= not (a xor b);
    layer1_outputs(5142) <= a;
    layer1_outputs(5143) <= b;
    layer1_outputs(5144) <= a xor b;
    layer1_outputs(5145) <= b;
    layer1_outputs(5146) <= not b or a;
    layer1_outputs(5147) <= a;
    layer1_outputs(5148) <= b;
    layer1_outputs(5149) <= b;
    layer1_outputs(5150) <= a and not b;
    layer1_outputs(5151) <= not a;
    layer1_outputs(5152) <= not (a xor b);
    layer1_outputs(5153) <= not a or b;
    layer1_outputs(5154) <= not (a and b);
    layer1_outputs(5155) <= not (a and b);
    layer1_outputs(5156) <= a xor b;
    layer1_outputs(5157) <= a xor b;
    layer1_outputs(5158) <= a and b;
    layer1_outputs(5159) <= not (a and b);
    layer1_outputs(5160) <= a xor b;
    layer1_outputs(5161) <= not a or b;
    layer1_outputs(5162) <= not a;
    layer1_outputs(5163) <= not b;
    layer1_outputs(5164) <= not b;
    layer1_outputs(5165) <= b;
    layer1_outputs(5166) <= a xor b;
    layer1_outputs(5167) <= not (a and b);
    layer1_outputs(5168) <= 1'b1;
    layer1_outputs(5169) <= not a or b;
    layer1_outputs(5170) <= not (a or b);
    layer1_outputs(5171) <= not (a xor b);
    layer1_outputs(5172) <= not (a xor b);
    layer1_outputs(5173) <= a and not b;
    layer1_outputs(5174) <= b;
    layer1_outputs(5175) <= not b;
    layer1_outputs(5176) <= b;
    layer1_outputs(5177) <= a and not b;
    layer1_outputs(5178) <= not b;
    layer1_outputs(5179) <= not (a or b);
    layer1_outputs(5180) <= a;
    layer1_outputs(5181) <= a or b;
    layer1_outputs(5182) <= not b;
    layer1_outputs(5183) <= not (a or b);
    layer1_outputs(5184) <= b and not a;
    layer1_outputs(5185) <= a or b;
    layer1_outputs(5186) <= b and not a;
    layer1_outputs(5187) <= not (a xor b);
    layer1_outputs(5188) <= b and not a;
    layer1_outputs(5189) <= not (a xor b);
    layer1_outputs(5190) <= b and not a;
    layer1_outputs(5191) <= not b or a;
    layer1_outputs(5192) <= not (a or b);
    layer1_outputs(5193) <= b;
    layer1_outputs(5194) <= a and b;
    layer1_outputs(5195) <= not (a xor b);
    layer1_outputs(5196) <= not a or b;
    layer1_outputs(5197) <= b and not a;
    layer1_outputs(5198) <= 1'b0;
    layer1_outputs(5199) <= not a or b;
    layer1_outputs(5200) <= not (a and b);
    layer1_outputs(5201) <= not a;
    layer1_outputs(5202) <= not (a and b);
    layer1_outputs(5203) <= a and b;
    layer1_outputs(5204) <= not (a and b);
    layer1_outputs(5205) <= a and not b;
    layer1_outputs(5206) <= not b or a;
    layer1_outputs(5207) <= not (a or b);
    layer1_outputs(5208) <= a xor b;
    layer1_outputs(5209) <= a xor b;
    layer1_outputs(5210) <= a;
    layer1_outputs(5211) <= a xor b;
    layer1_outputs(5212) <= a;
    layer1_outputs(5213) <= a;
    layer1_outputs(5214) <= b and not a;
    layer1_outputs(5215) <= a and not b;
    layer1_outputs(5216) <= not b;
    layer1_outputs(5217) <= not b;
    layer1_outputs(5218) <= a and b;
    layer1_outputs(5219) <= not a or b;
    layer1_outputs(5220) <= a or b;
    layer1_outputs(5221) <= not b or a;
    layer1_outputs(5222) <= not (a xor b);
    layer1_outputs(5223) <= a or b;
    layer1_outputs(5224) <= a and b;
    layer1_outputs(5225) <= a and b;
    layer1_outputs(5226) <= 1'b0;
    layer1_outputs(5227) <= a xor b;
    layer1_outputs(5228) <= not a;
    layer1_outputs(5229) <= not a or b;
    layer1_outputs(5230) <= b and not a;
    layer1_outputs(5231) <= not a or b;
    layer1_outputs(5232) <= not b;
    layer1_outputs(5233) <= not (a or b);
    layer1_outputs(5234) <= a or b;
    layer1_outputs(5235) <= a and not b;
    layer1_outputs(5236) <= not a;
    layer1_outputs(5237) <= not b or a;
    layer1_outputs(5238) <= not a;
    layer1_outputs(5239) <= not b or a;
    layer1_outputs(5240) <= not b or a;
    layer1_outputs(5241) <= not a or b;
    layer1_outputs(5242) <= not a or b;
    layer1_outputs(5243) <= a xor b;
    layer1_outputs(5244) <= not a or b;
    layer1_outputs(5245) <= 1'b0;
    layer1_outputs(5246) <= a and not b;
    layer1_outputs(5247) <= a and not b;
    layer1_outputs(5248) <= not a;
    layer1_outputs(5249) <= b and not a;
    layer1_outputs(5250) <= not (a and b);
    layer1_outputs(5251) <= a xor b;
    layer1_outputs(5252) <= not a or b;
    layer1_outputs(5253) <= not a or b;
    layer1_outputs(5254) <= not a;
    layer1_outputs(5255) <= not a;
    layer1_outputs(5256) <= b;
    layer1_outputs(5257) <= not a or b;
    layer1_outputs(5258) <= a xor b;
    layer1_outputs(5259) <= not b;
    layer1_outputs(5260) <= b;
    layer1_outputs(5261) <= a or b;
    layer1_outputs(5262) <= b and not a;
    layer1_outputs(5263) <= not b or a;
    layer1_outputs(5264) <= a xor b;
    layer1_outputs(5265) <= not (a xor b);
    layer1_outputs(5266) <= not (a or b);
    layer1_outputs(5267) <= a;
    layer1_outputs(5268) <= a xor b;
    layer1_outputs(5269) <= a and not b;
    layer1_outputs(5270) <= b;
    layer1_outputs(5271) <= not a;
    layer1_outputs(5272) <= not (a and b);
    layer1_outputs(5273) <= not a or b;
    layer1_outputs(5274) <= a and not b;
    layer1_outputs(5275) <= not (a or b);
    layer1_outputs(5276) <= a and not b;
    layer1_outputs(5277) <= b;
    layer1_outputs(5278) <= not b or a;
    layer1_outputs(5279) <= a;
    layer1_outputs(5280) <= not a;
    layer1_outputs(5281) <= a;
    layer1_outputs(5282) <= not (a and b);
    layer1_outputs(5283) <= a or b;
    layer1_outputs(5284) <= a xor b;
    layer1_outputs(5285) <= not a;
    layer1_outputs(5286) <= not a or b;
    layer1_outputs(5287) <= not b;
    layer1_outputs(5288) <= not a or b;
    layer1_outputs(5289) <= a and not b;
    layer1_outputs(5290) <= not (a or b);
    layer1_outputs(5291) <= a;
    layer1_outputs(5292) <= b and not a;
    layer1_outputs(5293) <= a xor b;
    layer1_outputs(5294) <= not (a xor b);
    layer1_outputs(5295) <= a and b;
    layer1_outputs(5296) <= not b;
    layer1_outputs(5297) <= not (a and b);
    layer1_outputs(5298) <= not a;
    layer1_outputs(5299) <= a xor b;
    layer1_outputs(5300) <= not (a xor b);
    layer1_outputs(5301) <= not a or b;
    layer1_outputs(5302) <= not (a or b);
    layer1_outputs(5303) <= not b;
    layer1_outputs(5304) <= a and b;
    layer1_outputs(5305) <= a xor b;
    layer1_outputs(5306) <= a or b;
    layer1_outputs(5307) <= a;
    layer1_outputs(5308) <= a;
    layer1_outputs(5309) <= a and b;
    layer1_outputs(5310) <= a and b;
    layer1_outputs(5311) <= a and b;
    layer1_outputs(5312) <= not b or a;
    layer1_outputs(5313) <= a and b;
    layer1_outputs(5314) <= a;
    layer1_outputs(5315) <= not (a and b);
    layer1_outputs(5316) <= a or b;
    layer1_outputs(5317) <= a xor b;
    layer1_outputs(5318) <= a and not b;
    layer1_outputs(5319) <= a and b;
    layer1_outputs(5320) <= not a or b;
    layer1_outputs(5321) <= a;
    layer1_outputs(5322) <= a and not b;
    layer1_outputs(5323) <= not b;
    layer1_outputs(5324) <= a and not b;
    layer1_outputs(5325) <= not b;
    layer1_outputs(5326) <= a and not b;
    layer1_outputs(5327) <= b;
    layer1_outputs(5328) <= b;
    layer1_outputs(5329) <= not a or b;
    layer1_outputs(5330) <= not a or b;
    layer1_outputs(5331) <= not b;
    layer1_outputs(5332) <= not a;
    layer1_outputs(5333) <= a and b;
    layer1_outputs(5334) <= a and not b;
    layer1_outputs(5335) <= a;
    layer1_outputs(5336) <= 1'b0;
    layer1_outputs(5337) <= a or b;
    layer1_outputs(5338) <= not (a or b);
    layer1_outputs(5339) <= not a;
    layer1_outputs(5340) <= b;
    layer1_outputs(5341) <= not a;
    layer1_outputs(5342) <= a and not b;
    layer1_outputs(5343) <= not b;
    layer1_outputs(5344) <= not (a and b);
    layer1_outputs(5345) <= not (a or b);
    layer1_outputs(5346) <= a xor b;
    layer1_outputs(5347) <= b and not a;
    layer1_outputs(5348) <= a or b;
    layer1_outputs(5349) <= not a;
    layer1_outputs(5350) <= b;
    layer1_outputs(5351) <= a xor b;
    layer1_outputs(5352) <= not b or a;
    layer1_outputs(5353) <= not (a or b);
    layer1_outputs(5354) <= a or b;
    layer1_outputs(5355) <= not a or b;
    layer1_outputs(5356) <= b and not a;
    layer1_outputs(5357) <= not (a xor b);
    layer1_outputs(5358) <= a;
    layer1_outputs(5359) <= a;
    layer1_outputs(5360) <= a;
    layer1_outputs(5361) <= a and not b;
    layer1_outputs(5362) <= not (a xor b);
    layer1_outputs(5363) <= not a or b;
    layer1_outputs(5364) <= not (a and b);
    layer1_outputs(5365) <= not (a or b);
    layer1_outputs(5366) <= not (a or b);
    layer1_outputs(5367) <= b and not a;
    layer1_outputs(5368) <= a and not b;
    layer1_outputs(5369) <= not a;
    layer1_outputs(5370) <= a and not b;
    layer1_outputs(5371) <= not b;
    layer1_outputs(5372) <= not a or b;
    layer1_outputs(5373) <= not (a xor b);
    layer1_outputs(5374) <= a;
    layer1_outputs(5375) <= b;
    layer1_outputs(5376) <= not a or b;
    layer1_outputs(5377) <= not (a or b);
    layer1_outputs(5378) <= a xor b;
    layer1_outputs(5379) <= not (a or b);
    layer1_outputs(5380) <= not b;
    layer1_outputs(5381) <= a and not b;
    layer1_outputs(5382) <= b;
    layer1_outputs(5383) <= a and not b;
    layer1_outputs(5384) <= b and not a;
    layer1_outputs(5385) <= not a or b;
    layer1_outputs(5386) <= not (a or b);
    layer1_outputs(5387) <= not a;
    layer1_outputs(5388) <= not b or a;
    layer1_outputs(5389) <= a and b;
    layer1_outputs(5390) <= 1'b0;
    layer1_outputs(5391) <= not (a xor b);
    layer1_outputs(5392) <= not a or b;
    layer1_outputs(5393) <= a;
    layer1_outputs(5394) <= a or b;
    layer1_outputs(5395) <= not b;
    layer1_outputs(5396) <= not a or b;
    layer1_outputs(5397) <= not (a xor b);
    layer1_outputs(5398) <= b and not a;
    layer1_outputs(5399) <= a and b;
    layer1_outputs(5400) <= b;
    layer1_outputs(5401) <= not b;
    layer1_outputs(5402) <= not b;
    layer1_outputs(5403) <= not (a or b);
    layer1_outputs(5404) <= not (a xor b);
    layer1_outputs(5405) <= b;
    layer1_outputs(5406) <= a xor b;
    layer1_outputs(5407) <= not b;
    layer1_outputs(5408) <= b;
    layer1_outputs(5409) <= not b or a;
    layer1_outputs(5410) <= not (a or b);
    layer1_outputs(5411) <= a and not b;
    layer1_outputs(5412) <= b;
    layer1_outputs(5413) <= not b or a;
    layer1_outputs(5414) <= not b;
    layer1_outputs(5415) <= a xor b;
    layer1_outputs(5416) <= not (a or b);
    layer1_outputs(5417) <= not b or a;
    layer1_outputs(5418) <= not (a or b);
    layer1_outputs(5419) <= not b or a;
    layer1_outputs(5420) <= b;
    layer1_outputs(5421) <= b;
    layer1_outputs(5422) <= b;
    layer1_outputs(5423) <= not b or a;
    layer1_outputs(5424) <= b;
    layer1_outputs(5425) <= not a;
    layer1_outputs(5426) <= a;
    layer1_outputs(5427) <= b;
    layer1_outputs(5428) <= not (a or b);
    layer1_outputs(5429) <= not a;
    layer1_outputs(5430) <= a and b;
    layer1_outputs(5431) <= not b;
    layer1_outputs(5432) <= not b or a;
    layer1_outputs(5433) <= a or b;
    layer1_outputs(5434) <= not (a xor b);
    layer1_outputs(5435) <= a xor b;
    layer1_outputs(5436) <= b;
    layer1_outputs(5437) <= not b;
    layer1_outputs(5438) <= not b;
    layer1_outputs(5439) <= not (a and b);
    layer1_outputs(5440) <= b;
    layer1_outputs(5441) <= a;
    layer1_outputs(5442) <= a or b;
    layer1_outputs(5443) <= not b or a;
    layer1_outputs(5444) <= a and not b;
    layer1_outputs(5445) <= not (a xor b);
    layer1_outputs(5446) <= not b or a;
    layer1_outputs(5447) <= not (a xor b);
    layer1_outputs(5448) <= not (a xor b);
    layer1_outputs(5449) <= a;
    layer1_outputs(5450) <= 1'b0;
    layer1_outputs(5451) <= not a;
    layer1_outputs(5452) <= not (a or b);
    layer1_outputs(5453) <= a and not b;
    layer1_outputs(5454) <= not (a xor b);
    layer1_outputs(5455) <= b;
    layer1_outputs(5456) <= not (a xor b);
    layer1_outputs(5457) <= not a;
    layer1_outputs(5458) <= a and not b;
    layer1_outputs(5459) <= not a;
    layer1_outputs(5460) <= a or b;
    layer1_outputs(5461) <= not a;
    layer1_outputs(5462) <= a and not b;
    layer1_outputs(5463) <= a xor b;
    layer1_outputs(5464) <= not (a xor b);
    layer1_outputs(5465) <= a xor b;
    layer1_outputs(5466) <= b;
    layer1_outputs(5467) <= not b;
    layer1_outputs(5468) <= a and not b;
    layer1_outputs(5469) <= not (a or b);
    layer1_outputs(5470) <= b and not a;
    layer1_outputs(5471) <= not (a xor b);
    layer1_outputs(5472) <= b and not a;
    layer1_outputs(5473) <= a xor b;
    layer1_outputs(5474) <= a;
    layer1_outputs(5475) <= not (a or b);
    layer1_outputs(5476) <= not a;
    layer1_outputs(5477) <= not a or b;
    layer1_outputs(5478) <= a;
    layer1_outputs(5479) <= not b;
    layer1_outputs(5480) <= not b;
    layer1_outputs(5481) <= not b;
    layer1_outputs(5482) <= a xor b;
    layer1_outputs(5483) <= b and not a;
    layer1_outputs(5484) <= b and not a;
    layer1_outputs(5485) <= not a or b;
    layer1_outputs(5486) <= b;
    layer1_outputs(5487) <= not (a xor b);
    layer1_outputs(5488) <= not (a and b);
    layer1_outputs(5489) <= a and b;
    layer1_outputs(5490) <= not (a and b);
    layer1_outputs(5491) <= not b;
    layer1_outputs(5492) <= not (a xor b);
    layer1_outputs(5493) <= a;
    layer1_outputs(5494) <= not (a and b);
    layer1_outputs(5495) <= a and b;
    layer1_outputs(5496) <= not (a or b);
    layer1_outputs(5497) <= a;
    layer1_outputs(5498) <= b and not a;
    layer1_outputs(5499) <= b;
    layer1_outputs(5500) <= b;
    layer1_outputs(5501) <= b and not a;
    layer1_outputs(5502) <= a;
    layer1_outputs(5503) <= not (a or b);
    layer1_outputs(5504) <= a and not b;
    layer1_outputs(5505) <= a;
    layer1_outputs(5506) <= a xor b;
    layer1_outputs(5507) <= 1'b1;
    layer1_outputs(5508) <= a xor b;
    layer1_outputs(5509) <= a xor b;
    layer1_outputs(5510) <= b;
    layer1_outputs(5511) <= a and not b;
    layer1_outputs(5512) <= not (a xor b);
    layer1_outputs(5513) <= b;
    layer1_outputs(5514) <= not a;
    layer1_outputs(5515) <= a;
    layer1_outputs(5516) <= b and not a;
    layer1_outputs(5517) <= not a;
    layer1_outputs(5518) <= a and b;
    layer1_outputs(5519) <= not (a or b);
    layer1_outputs(5520) <= not b;
    layer1_outputs(5521) <= not a or b;
    layer1_outputs(5522) <= not (a xor b);
    layer1_outputs(5523) <= a or b;
    layer1_outputs(5524) <= b and not a;
    layer1_outputs(5525) <= not (a and b);
    layer1_outputs(5526) <= not (a or b);
    layer1_outputs(5527) <= a;
    layer1_outputs(5528) <= a xor b;
    layer1_outputs(5529) <= b;
    layer1_outputs(5530) <= not a or b;
    layer1_outputs(5531) <= a;
    layer1_outputs(5532) <= a;
    layer1_outputs(5533) <= not (a or b);
    layer1_outputs(5534) <= not (a or b);
    layer1_outputs(5535) <= not a;
    layer1_outputs(5536) <= not (a and b);
    layer1_outputs(5537) <= a xor b;
    layer1_outputs(5538) <= b;
    layer1_outputs(5539) <= not b;
    layer1_outputs(5540) <= not (a or b);
    layer1_outputs(5541) <= not b or a;
    layer1_outputs(5542) <= a or b;
    layer1_outputs(5543) <= a and not b;
    layer1_outputs(5544) <= not (a or b);
    layer1_outputs(5545) <= not (a xor b);
    layer1_outputs(5546) <= a and not b;
    layer1_outputs(5547) <= a and b;
    layer1_outputs(5548) <= not b;
    layer1_outputs(5549) <= a xor b;
    layer1_outputs(5550) <= a or b;
    layer1_outputs(5551) <= a and b;
    layer1_outputs(5552) <= not (a xor b);
    layer1_outputs(5553) <= not (a and b);
    layer1_outputs(5554) <= b and not a;
    layer1_outputs(5555) <= b and not a;
    layer1_outputs(5556) <= not b or a;
    layer1_outputs(5557) <= a and b;
    layer1_outputs(5558) <= not (a xor b);
    layer1_outputs(5559) <= a or b;
    layer1_outputs(5560) <= b;
    layer1_outputs(5561) <= b;
    layer1_outputs(5562) <= a and not b;
    layer1_outputs(5563) <= not a;
    layer1_outputs(5564) <= a and b;
    layer1_outputs(5565) <= not b;
    layer1_outputs(5566) <= not (a xor b);
    layer1_outputs(5567) <= a;
    layer1_outputs(5568) <= a and b;
    layer1_outputs(5569) <= not b;
    layer1_outputs(5570) <= a;
    layer1_outputs(5571) <= a and not b;
    layer1_outputs(5572) <= a;
    layer1_outputs(5573) <= a or b;
    layer1_outputs(5574) <= b;
    layer1_outputs(5575) <= not (a xor b);
    layer1_outputs(5576) <= not (a or b);
    layer1_outputs(5577) <= b and not a;
    layer1_outputs(5578) <= a xor b;
    layer1_outputs(5579) <= not (a xor b);
    layer1_outputs(5580) <= not b or a;
    layer1_outputs(5581) <= a;
    layer1_outputs(5582) <= a and b;
    layer1_outputs(5583) <= not b or a;
    layer1_outputs(5584) <= not b;
    layer1_outputs(5585) <= a and not b;
    layer1_outputs(5586) <= not a;
    layer1_outputs(5587) <= not b or a;
    layer1_outputs(5588) <= a and b;
    layer1_outputs(5589) <= not (a xor b);
    layer1_outputs(5590) <= a and b;
    layer1_outputs(5591) <= not (a and b);
    layer1_outputs(5592) <= a and not b;
    layer1_outputs(5593) <= not (a and b);
    layer1_outputs(5594) <= not b;
    layer1_outputs(5595) <= b;
    layer1_outputs(5596) <= a;
    layer1_outputs(5597) <= b and not a;
    layer1_outputs(5598) <= not a;
    layer1_outputs(5599) <= a;
    layer1_outputs(5600) <= 1'b0;
    layer1_outputs(5601) <= a;
    layer1_outputs(5602) <= not a;
    layer1_outputs(5603) <= a and b;
    layer1_outputs(5604) <= not b;
    layer1_outputs(5605) <= a;
    layer1_outputs(5606) <= not b or a;
    layer1_outputs(5607) <= not a;
    layer1_outputs(5608) <= a and not b;
    layer1_outputs(5609) <= a xor b;
    layer1_outputs(5610) <= not (a xor b);
    layer1_outputs(5611) <= not b or a;
    layer1_outputs(5612) <= b and not a;
    layer1_outputs(5613) <= a;
    layer1_outputs(5614) <= a or b;
    layer1_outputs(5615) <= a and not b;
    layer1_outputs(5616) <= not b;
    layer1_outputs(5617) <= b and not a;
    layer1_outputs(5618) <= b and not a;
    layer1_outputs(5619) <= not a;
    layer1_outputs(5620) <= not a;
    layer1_outputs(5621) <= a and not b;
    layer1_outputs(5622) <= a or b;
    layer1_outputs(5623) <= a or b;
    layer1_outputs(5624) <= a and not b;
    layer1_outputs(5625) <= a;
    layer1_outputs(5626) <= a or b;
    layer1_outputs(5627) <= a and not b;
    layer1_outputs(5628) <= not a;
    layer1_outputs(5629) <= a and b;
    layer1_outputs(5630) <= not (a xor b);
    layer1_outputs(5631) <= not (a or b);
    layer1_outputs(5632) <= a or b;
    layer1_outputs(5633) <= b;
    layer1_outputs(5634) <= a and not b;
    layer1_outputs(5635) <= not a;
    layer1_outputs(5636) <= not a;
    layer1_outputs(5637) <= a;
    layer1_outputs(5638) <= not a;
    layer1_outputs(5639) <= not b or a;
    layer1_outputs(5640) <= a and b;
    layer1_outputs(5641) <= not b;
    layer1_outputs(5642) <= a;
    layer1_outputs(5643) <= a or b;
    layer1_outputs(5644) <= a and not b;
    layer1_outputs(5645) <= b;
    layer1_outputs(5646) <= b;
    layer1_outputs(5647) <= not (a xor b);
    layer1_outputs(5648) <= not b or a;
    layer1_outputs(5649) <= b and not a;
    layer1_outputs(5650) <= a;
    layer1_outputs(5651) <= not (a or b);
    layer1_outputs(5652) <= b;
    layer1_outputs(5653) <= b;
    layer1_outputs(5654) <= b;
    layer1_outputs(5655) <= not (a and b);
    layer1_outputs(5656) <= not a;
    layer1_outputs(5657) <= not (a and b);
    layer1_outputs(5658) <= a or b;
    layer1_outputs(5659) <= a;
    layer1_outputs(5660) <= not a or b;
    layer1_outputs(5661) <= not b;
    layer1_outputs(5662) <= a;
    layer1_outputs(5663) <= not (a xor b);
    layer1_outputs(5664) <= not a or b;
    layer1_outputs(5665) <= a and b;
    layer1_outputs(5666) <= not a;
    layer1_outputs(5667) <= not b;
    layer1_outputs(5668) <= b and not a;
    layer1_outputs(5669) <= not a;
    layer1_outputs(5670) <= not (a and b);
    layer1_outputs(5671) <= a xor b;
    layer1_outputs(5672) <= a and not b;
    layer1_outputs(5673) <= not (a or b);
    layer1_outputs(5674) <= not a or b;
    layer1_outputs(5675) <= a or b;
    layer1_outputs(5676) <= b and not a;
    layer1_outputs(5677) <= 1'b0;
    layer1_outputs(5678) <= not a or b;
    layer1_outputs(5679) <= not a or b;
    layer1_outputs(5680) <= b;
    layer1_outputs(5681) <= not b or a;
    layer1_outputs(5682) <= not (a or b);
    layer1_outputs(5683) <= not a or b;
    layer1_outputs(5684) <= not b;
    layer1_outputs(5685) <= not (a xor b);
    layer1_outputs(5686) <= not (a and b);
    layer1_outputs(5687) <= a and not b;
    layer1_outputs(5688) <= not (a or b);
    layer1_outputs(5689) <= a xor b;
    layer1_outputs(5690) <= a;
    layer1_outputs(5691) <= not b;
    layer1_outputs(5692) <= a;
    layer1_outputs(5693) <= a or b;
    layer1_outputs(5694) <= b and not a;
    layer1_outputs(5695) <= not b;
    layer1_outputs(5696) <= not a;
    layer1_outputs(5697) <= a and not b;
    layer1_outputs(5698) <= a and not b;
    layer1_outputs(5699) <= not (a xor b);
    layer1_outputs(5700) <= a or b;
    layer1_outputs(5701) <= not b;
    layer1_outputs(5702) <= not b;
    layer1_outputs(5703) <= not b;
    layer1_outputs(5704) <= b and not a;
    layer1_outputs(5705) <= not b or a;
    layer1_outputs(5706) <= a and not b;
    layer1_outputs(5707) <= not a;
    layer1_outputs(5708) <= not a or b;
    layer1_outputs(5709) <= a xor b;
    layer1_outputs(5710) <= a and not b;
    layer1_outputs(5711) <= not a;
    layer1_outputs(5712) <= a;
    layer1_outputs(5713) <= a and b;
    layer1_outputs(5714) <= not (a xor b);
    layer1_outputs(5715) <= b;
    layer1_outputs(5716) <= 1'b0;
    layer1_outputs(5717) <= a xor b;
    layer1_outputs(5718) <= not b;
    layer1_outputs(5719) <= a xor b;
    layer1_outputs(5720) <= a or b;
    layer1_outputs(5721) <= a and b;
    layer1_outputs(5722) <= not (a or b);
    layer1_outputs(5723) <= b and not a;
    layer1_outputs(5724) <= not (a xor b);
    layer1_outputs(5725) <= b;
    layer1_outputs(5726) <= a or b;
    layer1_outputs(5727) <= a;
    layer1_outputs(5728) <= not a;
    layer1_outputs(5729) <= b and not a;
    layer1_outputs(5730) <= not (a or b);
    layer1_outputs(5731) <= a;
    layer1_outputs(5732) <= not b or a;
    layer1_outputs(5733) <= a or b;
    layer1_outputs(5734) <= not a or b;
    layer1_outputs(5735) <= not b;
    layer1_outputs(5736) <= not a or b;
    layer1_outputs(5737) <= not b;
    layer1_outputs(5738) <= not (a and b);
    layer1_outputs(5739) <= not (a xor b);
    layer1_outputs(5740) <= not (a and b);
    layer1_outputs(5741) <= a and not b;
    layer1_outputs(5742) <= not a;
    layer1_outputs(5743) <= not (a xor b);
    layer1_outputs(5744) <= a;
    layer1_outputs(5745) <= not (a xor b);
    layer1_outputs(5746) <= not (a and b);
    layer1_outputs(5747) <= not a;
    layer1_outputs(5748) <= a and b;
    layer1_outputs(5749) <= not b or a;
    layer1_outputs(5750) <= not (a xor b);
    layer1_outputs(5751) <= not b or a;
    layer1_outputs(5752) <= a and b;
    layer1_outputs(5753) <= a and b;
    layer1_outputs(5754) <= not a or b;
    layer1_outputs(5755) <= not b;
    layer1_outputs(5756) <= a or b;
    layer1_outputs(5757) <= not (a or b);
    layer1_outputs(5758) <= not b or a;
    layer1_outputs(5759) <= 1'b1;
    layer1_outputs(5760) <= not a;
    layer1_outputs(5761) <= a and not b;
    layer1_outputs(5762) <= b;
    layer1_outputs(5763) <= a;
    layer1_outputs(5764) <= not (a and b);
    layer1_outputs(5765) <= not (a or b);
    layer1_outputs(5766) <= b;
    layer1_outputs(5767) <= a;
    layer1_outputs(5768) <= not b;
    layer1_outputs(5769) <= not (a and b);
    layer1_outputs(5770) <= not a;
    layer1_outputs(5771) <= a;
    layer1_outputs(5772) <= not b;
    layer1_outputs(5773) <= not (a or b);
    layer1_outputs(5774) <= a and not b;
    layer1_outputs(5775) <= a;
    layer1_outputs(5776) <= a;
    layer1_outputs(5777) <= not a;
    layer1_outputs(5778) <= not a;
    layer1_outputs(5779) <= a and not b;
    layer1_outputs(5780) <= a;
    layer1_outputs(5781) <= not (a xor b);
    layer1_outputs(5782) <= a or b;
    layer1_outputs(5783) <= a;
    layer1_outputs(5784) <= a xor b;
    layer1_outputs(5785) <= not a or b;
    layer1_outputs(5786) <= a and not b;
    layer1_outputs(5787) <= b;
    layer1_outputs(5788) <= not a;
    layer1_outputs(5789) <= a and not b;
    layer1_outputs(5790) <= b and not a;
    layer1_outputs(5791) <= not (a xor b);
    layer1_outputs(5792) <= not b or a;
    layer1_outputs(5793) <= not a or b;
    layer1_outputs(5794) <= a xor b;
    layer1_outputs(5795) <= b;
    layer1_outputs(5796) <= b;
    layer1_outputs(5797) <= not b;
    layer1_outputs(5798) <= a and b;
    layer1_outputs(5799) <= a xor b;
    layer1_outputs(5800) <= not (a xor b);
    layer1_outputs(5801) <= a and b;
    layer1_outputs(5802) <= a or b;
    layer1_outputs(5803) <= not (a and b);
    layer1_outputs(5804) <= not (a and b);
    layer1_outputs(5805) <= a;
    layer1_outputs(5806) <= a;
    layer1_outputs(5807) <= not (a xor b);
    layer1_outputs(5808) <= not (a or b);
    layer1_outputs(5809) <= a and not b;
    layer1_outputs(5810) <= b and not a;
    layer1_outputs(5811) <= b;
    layer1_outputs(5812) <= b;
    layer1_outputs(5813) <= a and not b;
    layer1_outputs(5814) <= a and not b;
    layer1_outputs(5815) <= b and not a;
    layer1_outputs(5816) <= not (a and b);
    layer1_outputs(5817) <= a xor b;
    layer1_outputs(5818) <= a xor b;
    layer1_outputs(5819) <= not b;
    layer1_outputs(5820) <= b;
    layer1_outputs(5821) <= not b or a;
    layer1_outputs(5822) <= a or b;
    layer1_outputs(5823) <= not (a and b);
    layer1_outputs(5824) <= not (a or b);
    layer1_outputs(5825) <= not (a and b);
    layer1_outputs(5826) <= not b;
    layer1_outputs(5827) <= a xor b;
    layer1_outputs(5828) <= not (a and b);
    layer1_outputs(5829) <= a and b;
    layer1_outputs(5830) <= a and b;
    layer1_outputs(5831) <= not (a xor b);
    layer1_outputs(5832) <= not b or a;
    layer1_outputs(5833) <= a or b;
    layer1_outputs(5834) <= not (a xor b);
    layer1_outputs(5835) <= not b or a;
    layer1_outputs(5836) <= a and b;
    layer1_outputs(5837) <= not a;
    layer1_outputs(5838) <= a and not b;
    layer1_outputs(5839) <= a and b;
    layer1_outputs(5840) <= a xor b;
    layer1_outputs(5841) <= not a or b;
    layer1_outputs(5842) <= not (a xor b);
    layer1_outputs(5843) <= a xor b;
    layer1_outputs(5844) <= not (a and b);
    layer1_outputs(5845) <= not (a and b);
    layer1_outputs(5846) <= a xor b;
    layer1_outputs(5847) <= not a;
    layer1_outputs(5848) <= not b or a;
    layer1_outputs(5849) <= not (a xor b);
    layer1_outputs(5850) <= not (a and b);
    layer1_outputs(5851) <= not a;
    layer1_outputs(5852) <= b and not a;
    layer1_outputs(5853) <= a;
    layer1_outputs(5854) <= not (a xor b);
    layer1_outputs(5855) <= not b;
    layer1_outputs(5856) <= not b;
    layer1_outputs(5857) <= a;
    layer1_outputs(5858) <= not a;
    layer1_outputs(5859) <= a xor b;
    layer1_outputs(5860) <= a or b;
    layer1_outputs(5861) <= not b or a;
    layer1_outputs(5862) <= a xor b;
    layer1_outputs(5863) <= not a;
    layer1_outputs(5864) <= a;
    layer1_outputs(5865) <= a xor b;
    layer1_outputs(5866) <= a;
    layer1_outputs(5867) <= a;
    layer1_outputs(5868) <= 1'b0;
    layer1_outputs(5869) <= not a or b;
    layer1_outputs(5870) <= a;
    layer1_outputs(5871) <= a and b;
    layer1_outputs(5872) <= a or b;
    layer1_outputs(5873) <= b and not a;
    layer1_outputs(5874) <= a and not b;
    layer1_outputs(5875) <= not (a xor b);
    layer1_outputs(5876) <= a;
    layer1_outputs(5877) <= b and not a;
    layer1_outputs(5878) <= not b;
    layer1_outputs(5879) <= b and not a;
    layer1_outputs(5880) <= a and not b;
    layer1_outputs(5881) <= 1'b0;
    layer1_outputs(5882) <= not (a xor b);
    layer1_outputs(5883) <= not a;
    layer1_outputs(5884) <= b;
    layer1_outputs(5885) <= a and b;
    layer1_outputs(5886) <= not (a xor b);
    layer1_outputs(5887) <= not (a xor b);
    layer1_outputs(5888) <= 1'b1;
    layer1_outputs(5889) <= not a or b;
    layer1_outputs(5890) <= b;
    layer1_outputs(5891) <= not (a xor b);
    layer1_outputs(5892) <= a and not b;
    layer1_outputs(5893) <= not a;
    layer1_outputs(5894) <= 1'b1;
    layer1_outputs(5895) <= a;
    layer1_outputs(5896) <= not a or b;
    layer1_outputs(5897) <= a xor b;
    layer1_outputs(5898) <= not a;
    layer1_outputs(5899) <= a;
    layer1_outputs(5900) <= a;
    layer1_outputs(5901) <= not (a and b);
    layer1_outputs(5902) <= b;
    layer1_outputs(5903) <= not b;
    layer1_outputs(5904) <= not (a or b);
    layer1_outputs(5905) <= not a;
    layer1_outputs(5906) <= a xor b;
    layer1_outputs(5907) <= not a or b;
    layer1_outputs(5908) <= not (a or b);
    layer1_outputs(5909) <= a or b;
    layer1_outputs(5910) <= not a;
    layer1_outputs(5911) <= not a;
    layer1_outputs(5912) <= b and not a;
    layer1_outputs(5913) <= not a;
    layer1_outputs(5914) <= not a;
    layer1_outputs(5915) <= a xor b;
    layer1_outputs(5916) <= b and not a;
    layer1_outputs(5917) <= a or b;
    layer1_outputs(5918) <= a xor b;
    layer1_outputs(5919) <= not b;
    layer1_outputs(5920) <= a xor b;
    layer1_outputs(5921) <= not (a and b);
    layer1_outputs(5922) <= not a;
    layer1_outputs(5923) <= not (a or b);
    layer1_outputs(5924) <= a;
    layer1_outputs(5925) <= not (a xor b);
    layer1_outputs(5926) <= a and not b;
    layer1_outputs(5927) <= not b;
    layer1_outputs(5928) <= not a;
    layer1_outputs(5929) <= a or b;
    layer1_outputs(5930) <= a or b;
    layer1_outputs(5931) <= not (a and b);
    layer1_outputs(5932) <= not (a or b);
    layer1_outputs(5933) <= not (a and b);
    layer1_outputs(5934) <= not (a xor b);
    layer1_outputs(5935) <= a xor b;
    layer1_outputs(5936) <= not (a xor b);
    layer1_outputs(5937) <= a xor b;
    layer1_outputs(5938) <= not b or a;
    layer1_outputs(5939) <= b;
    layer1_outputs(5940) <= not b or a;
    layer1_outputs(5941) <= not a or b;
    layer1_outputs(5942) <= b and not a;
    layer1_outputs(5943) <= not (a or b);
    layer1_outputs(5944) <= not (a or b);
    layer1_outputs(5945) <= b and not a;
    layer1_outputs(5946) <= b and not a;
    layer1_outputs(5947) <= not a;
    layer1_outputs(5948) <= not (a xor b);
    layer1_outputs(5949) <= not a;
    layer1_outputs(5950) <= not b;
    layer1_outputs(5951) <= not a or b;
    layer1_outputs(5952) <= a and not b;
    layer1_outputs(5953) <= a or b;
    layer1_outputs(5954) <= 1'b1;
    layer1_outputs(5955) <= not a or b;
    layer1_outputs(5956) <= b and not a;
    layer1_outputs(5957) <= not a;
    layer1_outputs(5958) <= b;
    layer1_outputs(5959) <= not b or a;
    layer1_outputs(5960) <= a;
    layer1_outputs(5961) <= b;
    layer1_outputs(5962) <= a or b;
    layer1_outputs(5963) <= not b or a;
    layer1_outputs(5964) <= a;
    layer1_outputs(5965) <= not (a xor b);
    layer1_outputs(5966) <= a;
    layer1_outputs(5967) <= a and b;
    layer1_outputs(5968) <= a or b;
    layer1_outputs(5969) <= a;
    layer1_outputs(5970) <= a xor b;
    layer1_outputs(5971) <= not a or b;
    layer1_outputs(5972) <= 1'b0;
    layer1_outputs(5973) <= b;
    layer1_outputs(5974) <= not b or a;
    layer1_outputs(5975) <= a and b;
    layer1_outputs(5976) <= a;
    layer1_outputs(5977) <= not (a xor b);
    layer1_outputs(5978) <= not a or b;
    layer1_outputs(5979) <= not b;
    layer1_outputs(5980) <= not b;
    layer1_outputs(5981) <= not b or a;
    layer1_outputs(5982) <= a;
    layer1_outputs(5983) <= not (a xor b);
    layer1_outputs(5984) <= not b;
    layer1_outputs(5985) <= not a;
    layer1_outputs(5986) <= not b;
    layer1_outputs(5987) <= not (a xor b);
    layer1_outputs(5988) <= a;
    layer1_outputs(5989) <= not (a xor b);
    layer1_outputs(5990) <= a and b;
    layer1_outputs(5991) <= a or b;
    layer1_outputs(5992) <= not (a or b);
    layer1_outputs(5993) <= not a or b;
    layer1_outputs(5994) <= a xor b;
    layer1_outputs(5995) <= not a or b;
    layer1_outputs(5996) <= not (a or b);
    layer1_outputs(5997) <= not (a xor b);
    layer1_outputs(5998) <= not a;
    layer1_outputs(5999) <= not (a or b);
    layer1_outputs(6000) <= not a or b;
    layer1_outputs(6001) <= a and b;
    layer1_outputs(6002) <= b;
    layer1_outputs(6003) <= b and not a;
    layer1_outputs(6004) <= a and b;
    layer1_outputs(6005) <= a or b;
    layer1_outputs(6006) <= not (a or b);
    layer1_outputs(6007) <= not (a xor b);
    layer1_outputs(6008) <= not a;
    layer1_outputs(6009) <= b and not a;
    layer1_outputs(6010) <= not a;
    layer1_outputs(6011) <= not a;
    layer1_outputs(6012) <= not (a xor b);
    layer1_outputs(6013) <= not a;
    layer1_outputs(6014) <= a;
    layer1_outputs(6015) <= not b;
    layer1_outputs(6016) <= a or b;
    layer1_outputs(6017) <= not a;
    layer1_outputs(6018) <= a xor b;
    layer1_outputs(6019) <= a or b;
    layer1_outputs(6020) <= a or b;
    layer1_outputs(6021) <= a;
    layer1_outputs(6022) <= not a;
    layer1_outputs(6023) <= b and not a;
    layer1_outputs(6024) <= b;
    layer1_outputs(6025) <= not a;
    layer1_outputs(6026) <= a and b;
    layer1_outputs(6027) <= not (a xor b);
    layer1_outputs(6028) <= a xor b;
    layer1_outputs(6029) <= b;
    layer1_outputs(6030) <= not b;
    layer1_outputs(6031) <= not (a xor b);
    layer1_outputs(6032) <= a and not b;
    layer1_outputs(6033) <= a xor b;
    layer1_outputs(6034) <= a xor b;
    layer1_outputs(6035) <= not (a and b);
    layer1_outputs(6036) <= b and not a;
    layer1_outputs(6037) <= a or b;
    layer1_outputs(6038) <= a xor b;
    layer1_outputs(6039) <= a;
    layer1_outputs(6040) <= not (a and b);
    layer1_outputs(6041) <= not a;
    layer1_outputs(6042) <= not a or b;
    layer1_outputs(6043) <= a and not b;
    layer1_outputs(6044) <= a;
    layer1_outputs(6045) <= not (a and b);
    layer1_outputs(6046) <= b;
    layer1_outputs(6047) <= a and not b;
    layer1_outputs(6048) <= a xor b;
    layer1_outputs(6049) <= not (a xor b);
    layer1_outputs(6050) <= not a or b;
    layer1_outputs(6051) <= b;
    layer1_outputs(6052) <= a or b;
    layer1_outputs(6053) <= b;
    layer1_outputs(6054) <= not a;
    layer1_outputs(6055) <= a;
    layer1_outputs(6056) <= a and b;
    layer1_outputs(6057) <= not a or b;
    layer1_outputs(6058) <= not a;
    layer1_outputs(6059) <= a and not b;
    layer1_outputs(6060) <= not a;
    layer1_outputs(6061) <= a xor b;
    layer1_outputs(6062) <= not (a or b);
    layer1_outputs(6063) <= not b or a;
    layer1_outputs(6064) <= a and b;
    layer1_outputs(6065) <= a or b;
    layer1_outputs(6066) <= not a or b;
    layer1_outputs(6067) <= not (a or b);
    layer1_outputs(6068) <= b and not a;
    layer1_outputs(6069) <= not (a xor b);
    layer1_outputs(6070) <= a;
    layer1_outputs(6071) <= 1'b1;
    layer1_outputs(6072) <= a xor b;
    layer1_outputs(6073) <= a or b;
    layer1_outputs(6074) <= b;
    layer1_outputs(6075) <= a or b;
    layer1_outputs(6076) <= a or b;
    layer1_outputs(6077) <= not a;
    layer1_outputs(6078) <= not b;
    layer1_outputs(6079) <= a;
    layer1_outputs(6080) <= a and b;
    layer1_outputs(6081) <= not (a xor b);
    layer1_outputs(6082) <= not (a xor b);
    layer1_outputs(6083) <= not b or a;
    layer1_outputs(6084) <= not (a xor b);
    layer1_outputs(6085) <= not (a xor b);
    layer1_outputs(6086) <= not (a or b);
    layer1_outputs(6087) <= not b or a;
    layer1_outputs(6088) <= not (a and b);
    layer1_outputs(6089) <= b;
    layer1_outputs(6090) <= b and not a;
    layer1_outputs(6091) <= a;
    layer1_outputs(6092) <= not (a or b);
    layer1_outputs(6093) <= b;
    layer1_outputs(6094) <= a or b;
    layer1_outputs(6095) <= not a or b;
    layer1_outputs(6096) <= not b;
    layer1_outputs(6097) <= not b or a;
    layer1_outputs(6098) <= not (a xor b);
    layer1_outputs(6099) <= b and not a;
    layer1_outputs(6100) <= 1'b1;
    layer1_outputs(6101) <= b and not a;
    layer1_outputs(6102) <= not b;
    layer1_outputs(6103) <= not b or a;
    layer1_outputs(6104) <= not b or a;
    layer1_outputs(6105) <= b;
    layer1_outputs(6106) <= a and not b;
    layer1_outputs(6107) <= not (a and b);
    layer1_outputs(6108) <= a;
    layer1_outputs(6109) <= not (a xor b);
    layer1_outputs(6110) <= not a or b;
    layer1_outputs(6111) <= b;
    layer1_outputs(6112) <= a and b;
    layer1_outputs(6113) <= not (a or b);
    layer1_outputs(6114) <= 1'b1;
    layer1_outputs(6115) <= b;
    layer1_outputs(6116) <= a xor b;
    layer1_outputs(6117) <= b;
    layer1_outputs(6118) <= not (a and b);
    layer1_outputs(6119) <= b;
    layer1_outputs(6120) <= a xor b;
    layer1_outputs(6121) <= a xor b;
    layer1_outputs(6122) <= not b or a;
    layer1_outputs(6123) <= a and not b;
    layer1_outputs(6124) <= not b;
    layer1_outputs(6125) <= not a;
    layer1_outputs(6126) <= a;
    layer1_outputs(6127) <= not (a and b);
    layer1_outputs(6128) <= a and not b;
    layer1_outputs(6129) <= a or b;
    layer1_outputs(6130) <= not (a and b);
    layer1_outputs(6131) <= not (a or b);
    layer1_outputs(6132) <= not b;
    layer1_outputs(6133) <= a or b;
    layer1_outputs(6134) <= b;
    layer1_outputs(6135) <= a and not b;
    layer1_outputs(6136) <= b;
    layer1_outputs(6137) <= not a;
    layer1_outputs(6138) <= a or b;
    layer1_outputs(6139) <= a;
    layer1_outputs(6140) <= not b or a;
    layer1_outputs(6141) <= b and not a;
    layer1_outputs(6142) <= not (a xor b);
    layer1_outputs(6143) <= a;
    layer1_outputs(6144) <= a or b;
    layer1_outputs(6145) <= a and not b;
    layer1_outputs(6146) <= a and not b;
    layer1_outputs(6147) <= not b or a;
    layer1_outputs(6148) <= not a;
    layer1_outputs(6149) <= b;
    layer1_outputs(6150) <= not (a and b);
    layer1_outputs(6151) <= not b or a;
    layer1_outputs(6152) <= b;
    layer1_outputs(6153) <= not b;
    layer1_outputs(6154) <= b and not a;
    layer1_outputs(6155) <= not (a xor b);
    layer1_outputs(6156) <= not b;
    layer1_outputs(6157) <= not (a and b);
    layer1_outputs(6158) <= b and not a;
    layer1_outputs(6159) <= not b;
    layer1_outputs(6160) <= not b;
    layer1_outputs(6161) <= a xor b;
    layer1_outputs(6162) <= not b;
    layer1_outputs(6163) <= a or b;
    layer1_outputs(6164) <= not a or b;
    layer1_outputs(6165) <= not a or b;
    layer1_outputs(6166) <= a and b;
    layer1_outputs(6167) <= a and not b;
    layer1_outputs(6168) <= a;
    layer1_outputs(6169) <= not b or a;
    layer1_outputs(6170) <= a and b;
    layer1_outputs(6171) <= not b;
    layer1_outputs(6172) <= a and b;
    layer1_outputs(6173) <= not (a or b);
    layer1_outputs(6174) <= not b or a;
    layer1_outputs(6175) <= b;
    layer1_outputs(6176) <= a xor b;
    layer1_outputs(6177) <= b;
    layer1_outputs(6178) <= a and b;
    layer1_outputs(6179) <= not (a or b);
    layer1_outputs(6180) <= not (a and b);
    layer1_outputs(6181) <= a xor b;
    layer1_outputs(6182) <= a xor b;
    layer1_outputs(6183) <= not b;
    layer1_outputs(6184) <= b and not a;
    layer1_outputs(6185) <= a and b;
    layer1_outputs(6186) <= not (a and b);
    layer1_outputs(6187) <= a and b;
    layer1_outputs(6188) <= not a;
    layer1_outputs(6189) <= a;
    layer1_outputs(6190) <= not b or a;
    layer1_outputs(6191) <= a;
    layer1_outputs(6192) <= not a;
    layer1_outputs(6193) <= not a or b;
    layer1_outputs(6194) <= a or b;
    layer1_outputs(6195) <= not (a xor b);
    layer1_outputs(6196) <= not (a or b);
    layer1_outputs(6197) <= b and not a;
    layer1_outputs(6198) <= not b or a;
    layer1_outputs(6199) <= not b;
    layer1_outputs(6200) <= not a;
    layer1_outputs(6201) <= not (a or b);
    layer1_outputs(6202) <= b;
    layer1_outputs(6203) <= not b;
    layer1_outputs(6204) <= b and not a;
    layer1_outputs(6205) <= not (a and b);
    layer1_outputs(6206) <= a xor b;
    layer1_outputs(6207) <= a;
    layer1_outputs(6208) <= b and not a;
    layer1_outputs(6209) <= a;
    layer1_outputs(6210) <= a and not b;
    layer1_outputs(6211) <= not b;
    layer1_outputs(6212) <= not (a or b);
    layer1_outputs(6213) <= not a;
    layer1_outputs(6214) <= not a;
    layer1_outputs(6215) <= not b;
    layer1_outputs(6216) <= not b or a;
    layer1_outputs(6217) <= b and not a;
    layer1_outputs(6218) <= a xor b;
    layer1_outputs(6219) <= a xor b;
    layer1_outputs(6220) <= a;
    layer1_outputs(6221) <= not b or a;
    layer1_outputs(6222) <= a;
    layer1_outputs(6223) <= a xor b;
    layer1_outputs(6224) <= a and b;
    layer1_outputs(6225) <= a and not b;
    layer1_outputs(6226) <= not a;
    layer1_outputs(6227) <= not a;
    layer1_outputs(6228) <= a and b;
    layer1_outputs(6229) <= a;
    layer1_outputs(6230) <= b;
    layer1_outputs(6231) <= a and b;
    layer1_outputs(6232) <= not (a xor b);
    layer1_outputs(6233) <= a;
    layer1_outputs(6234) <= not a or b;
    layer1_outputs(6235) <= a xor b;
    layer1_outputs(6236) <= not (a and b);
    layer1_outputs(6237) <= a;
    layer1_outputs(6238) <= a xor b;
    layer1_outputs(6239) <= not a;
    layer1_outputs(6240) <= not a;
    layer1_outputs(6241) <= 1'b0;
    layer1_outputs(6242) <= b;
    layer1_outputs(6243) <= not b or a;
    layer1_outputs(6244) <= not b;
    layer1_outputs(6245) <= not (a xor b);
    layer1_outputs(6246) <= b;
    layer1_outputs(6247) <= a;
    layer1_outputs(6248) <= not (a and b);
    layer1_outputs(6249) <= not (a xor b);
    layer1_outputs(6250) <= b;
    layer1_outputs(6251) <= a or b;
    layer1_outputs(6252) <= not a;
    layer1_outputs(6253) <= a and not b;
    layer1_outputs(6254) <= not (a xor b);
    layer1_outputs(6255) <= a xor b;
    layer1_outputs(6256) <= b;
    layer1_outputs(6257) <= a;
    layer1_outputs(6258) <= not b or a;
    layer1_outputs(6259) <= not a;
    layer1_outputs(6260) <= not a or b;
    layer1_outputs(6261) <= b;
    layer1_outputs(6262) <= a;
    layer1_outputs(6263) <= a or b;
    layer1_outputs(6264) <= a xor b;
    layer1_outputs(6265) <= a;
    layer1_outputs(6266) <= not b;
    layer1_outputs(6267) <= b;
    layer1_outputs(6268) <= a;
    layer1_outputs(6269) <= b and not a;
    layer1_outputs(6270) <= not b;
    layer1_outputs(6271) <= not a;
    layer1_outputs(6272) <= b;
    layer1_outputs(6273) <= not a;
    layer1_outputs(6274) <= not b;
    layer1_outputs(6275) <= not b or a;
    layer1_outputs(6276) <= b;
    layer1_outputs(6277) <= b;
    layer1_outputs(6278) <= not (a xor b);
    layer1_outputs(6279) <= a and not b;
    layer1_outputs(6280) <= not a;
    layer1_outputs(6281) <= not a;
    layer1_outputs(6282) <= not b;
    layer1_outputs(6283) <= a;
    layer1_outputs(6284) <= a xor b;
    layer1_outputs(6285) <= a and b;
    layer1_outputs(6286) <= not a;
    layer1_outputs(6287) <= not a;
    layer1_outputs(6288) <= not (a or b);
    layer1_outputs(6289) <= not (a and b);
    layer1_outputs(6290) <= a and b;
    layer1_outputs(6291) <= a;
    layer1_outputs(6292) <= not b;
    layer1_outputs(6293) <= b;
    layer1_outputs(6294) <= not a;
    layer1_outputs(6295) <= b and not a;
    layer1_outputs(6296) <= b;
    layer1_outputs(6297) <= not b;
    layer1_outputs(6298) <= not (a and b);
    layer1_outputs(6299) <= not (a or b);
    layer1_outputs(6300) <= not a;
    layer1_outputs(6301) <= not b;
    layer1_outputs(6302) <= a;
    layer1_outputs(6303) <= not a;
    layer1_outputs(6304) <= 1'b0;
    layer1_outputs(6305) <= not (a xor b);
    layer1_outputs(6306) <= a;
    layer1_outputs(6307) <= a xor b;
    layer1_outputs(6308) <= not (a or b);
    layer1_outputs(6309) <= b and not a;
    layer1_outputs(6310) <= not b;
    layer1_outputs(6311) <= b and not a;
    layer1_outputs(6312) <= a or b;
    layer1_outputs(6313) <= b and not a;
    layer1_outputs(6314) <= b;
    layer1_outputs(6315) <= a and b;
    layer1_outputs(6316) <= 1'b1;
    layer1_outputs(6317) <= not (a or b);
    layer1_outputs(6318) <= not a or b;
    layer1_outputs(6319) <= not (a or b);
    layer1_outputs(6320) <= b;
    layer1_outputs(6321) <= a and b;
    layer1_outputs(6322) <= b;
    layer1_outputs(6323) <= b;
    layer1_outputs(6324) <= a;
    layer1_outputs(6325) <= a or b;
    layer1_outputs(6326) <= not b;
    layer1_outputs(6327) <= b and not a;
    layer1_outputs(6328) <= a and not b;
    layer1_outputs(6329) <= not b;
    layer1_outputs(6330) <= not (a xor b);
    layer1_outputs(6331) <= not a or b;
    layer1_outputs(6332) <= not b;
    layer1_outputs(6333) <= a xor b;
    layer1_outputs(6334) <= b and not a;
    layer1_outputs(6335) <= not b or a;
    layer1_outputs(6336) <= not (a xor b);
    layer1_outputs(6337) <= not b;
    layer1_outputs(6338) <= a or b;
    layer1_outputs(6339) <= b and not a;
    layer1_outputs(6340) <= a and not b;
    layer1_outputs(6341) <= not a or b;
    layer1_outputs(6342) <= not (a or b);
    layer1_outputs(6343) <= not a or b;
    layer1_outputs(6344) <= not (a or b);
    layer1_outputs(6345) <= not b or a;
    layer1_outputs(6346) <= not (a and b);
    layer1_outputs(6347) <= a xor b;
    layer1_outputs(6348) <= a and b;
    layer1_outputs(6349) <= b;
    layer1_outputs(6350) <= not a;
    layer1_outputs(6351) <= a;
    layer1_outputs(6352) <= a;
    layer1_outputs(6353) <= not (a xor b);
    layer1_outputs(6354) <= a and not b;
    layer1_outputs(6355) <= a and b;
    layer1_outputs(6356) <= a;
    layer1_outputs(6357) <= a and not b;
    layer1_outputs(6358) <= not (a or b);
    layer1_outputs(6359) <= not (a xor b);
    layer1_outputs(6360) <= 1'b1;
    layer1_outputs(6361) <= a;
    layer1_outputs(6362) <= not a or b;
    layer1_outputs(6363) <= b and not a;
    layer1_outputs(6364) <= not b or a;
    layer1_outputs(6365) <= a xor b;
    layer1_outputs(6366) <= not (a or b);
    layer1_outputs(6367) <= b;
    layer1_outputs(6368) <= not (a and b);
    layer1_outputs(6369) <= a or b;
    layer1_outputs(6370) <= a and not b;
    layer1_outputs(6371) <= not a;
    layer1_outputs(6372) <= a and not b;
    layer1_outputs(6373) <= b;
    layer1_outputs(6374) <= a or b;
    layer1_outputs(6375) <= not a;
    layer1_outputs(6376) <= not (a and b);
    layer1_outputs(6377) <= b;
    layer1_outputs(6378) <= a;
    layer1_outputs(6379) <= not b;
    layer1_outputs(6380) <= b;
    layer1_outputs(6381) <= not b;
    layer1_outputs(6382) <= not (a xor b);
    layer1_outputs(6383) <= b;
    layer1_outputs(6384) <= not (a or b);
    layer1_outputs(6385) <= not a;
    layer1_outputs(6386) <= b;
    layer1_outputs(6387) <= not (a or b);
    layer1_outputs(6388) <= a;
    layer1_outputs(6389) <= not b;
    layer1_outputs(6390) <= a xor b;
    layer1_outputs(6391) <= not b;
    layer1_outputs(6392) <= a xor b;
    layer1_outputs(6393) <= 1'b0;
    layer1_outputs(6394) <= not b;
    layer1_outputs(6395) <= b and not a;
    layer1_outputs(6396) <= 1'b1;
    layer1_outputs(6397) <= b and not a;
    layer1_outputs(6398) <= not (a or b);
    layer1_outputs(6399) <= a xor b;
    layer1_outputs(6400) <= a and b;
    layer1_outputs(6401) <= not a;
    layer1_outputs(6402) <= a and b;
    layer1_outputs(6403) <= b;
    layer1_outputs(6404) <= not (a xor b);
    layer1_outputs(6405) <= not a or b;
    layer1_outputs(6406) <= a;
    layer1_outputs(6407) <= not b or a;
    layer1_outputs(6408) <= not (a xor b);
    layer1_outputs(6409) <= b;
    layer1_outputs(6410) <= not b;
    layer1_outputs(6411) <= not b or a;
    layer1_outputs(6412) <= a and not b;
    layer1_outputs(6413) <= not (a xor b);
    layer1_outputs(6414) <= a;
    layer1_outputs(6415) <= not (a and b);
    layer1_outputs(6416) <= not a;
    layer1_outputs(6417) <= b and not a;
    layer1_outputs(6418) <= a;
    layer1_outputs(6419) <= not (a and b);
    layer1_outputs(6420) <= a xor b;
    layer1_outputs(6421) <= not (a xor b);
    layer1_outputs(6422) <= not (a and b);
    layer1_outputs(6423) <= a and b;
    layer1_outputs(6424) <= 1'b0;
    layer1_outputs(6425) <= not b;
    layer1_outputs(6426) <= not a or b;
    layer1_outputs(6427) <= not b;
    layer1_outputs(6428) <= not a;
    layer1_outputs(6429) <= not a or b;
    layer1_outputs(6430) <= a;
    layer1_outputs(6431) <= not (a and b);
    layer1_outputs(6432) <= not b;
    layer1_outputs(6433) <= a xor b;
    layer1_outputs(6434) <= b;
    layer1_outputs(6435) <= not (a xor b);
    layer1_outputs(6436) <= 1'b0;
    layer1_outputs(6437) <= b and not a;
    layer1_outputs(6438) <= not a;
    layer1_outputs(6439) <= not (a and b);
    layer1_outputs(6440) <= a or b;
    layer1_outputs(6441) <= not a or b;
    layer1_outputs(6442) <= a and not b;
    layer1_outputs(6443) <= b and not a;
    layer1_outputs(6444) <= not (a xor b);
    layer1_outputs(6445) <= not (a or b);
    layer1_outputs(6446) <= not b;
    layer1_outputs(6447) <= a;
    layer1_outputs(6448) <= b;
    layer1_outputs(6449) <= a xor b;
    layer1_outputs(6450) <= not a;
    layer1_outputs(6451) <= a and b;
    layer1_outputs(6452) <= not b or a;
    layer1_outputs(6453) <= a xor b;
    layer1_outputs(6454) <= not b;
    layer1_outputs(6455) <= not (a or b);
    layer1_outputs(6456) <= not (a or b);
    layer1_outputs(6457) <= not (a and b);
    layer1_outputs(6458) <= not b;
    layer1_outputs(6459) <= not a;
    layer1_outputs(6460) <= a;
    layer1_outputs(6461) <= b;
    layer1_outputs(6462) <= not a or b;
    layer1_outputs(6463) <= not a;
    layer1_outputs(6464) <= a or b;
    layer1_outputs(6465) <= not (a and b);
    layer1_outputs(6466) <= not (a or b);
    layer1_outputs(6467) <= 1'b0;
    layer1_outputs(6468) <= a xor b;
    layer1_outputs(6469) <= b and not a;
    layer1_outputs(6470) <= a and b;
    layer1_outputs(6471) <= a and b;
    layer1_outputs(6472) <= not a or b;
    layer1_outputs(6473) <= a xor b;
    layer1_outputs(6474) <= b;
    layer1_outputs(6475) <= a or b;
    layer1_outputs(6476) <= a and not b;
    layer1_outputs(6477) <= not a;
    layer1_outputs(6478) <= a and not b;
    layer1_outputs(6479) <= a xor b;
    layer1_outputs(6480) <= a;
    layer1_outputs(6481) <= a and b;
    layer1_outputs(6482) <= a and not b;
    layer1_outputs(6483) <= a or b;
    layer1_outputs(6484) <= not b or a;
    layer1_outputs(6485) <= a or b;
    layer1_outputs(6486) <= a or b;
    layer1_outputs(6487) <= b and not a;
    layer1_outputs(6488) <= not b;
    layer1_outputs(6489) <= 1'b0;
    layer1_outputs(6490) <= a;
    layer1_outputs(6491) <= not (a or b);
    layer1_outputs(6492) <= not (a xor b);
    layer1_outputs(6493) <= a xor b;
    layer1_outputs(6494) <= not (a xor b);
    layer1_outputs(6495) <= a and b;
    layer1_outputs(6496) <= not a;
    layer1_outputs(6497) <= a xor b;
    layer1_outputs(6498) <= a or b;
    layer1_outputs(6499) <= not a;
    layer1_outputs(6500) <= a or b;
    layer1_outputs(6501) <= not a;
    layer1_outputs(6502) <= not a;
    layer1_outputs(6503) <= 1'b1;
    layer1_outputs(6504) <= not b;
    layer1_outputs(6505) <= not a;
    layer1_outputs(6506) <= b;
    layer1_outputs(6507) <= a xor b;
    layer1_outputs(6508) <= not (a xor b);
    layer1_outputs(6509) <= a and not b;
    layer1_outputs(6510) <= b;
    layer1_outputs(6511) <= a and not b;
    layer1_outputs(6512) <= not b or a;
    layer1_outputs(6513) <= a and not b;
    layer1_outputs(6514) <= not (a and b);
    layer1_outputs(6515) <= b;
    layer1_outputs(6516) <= b;
    layer1_outputs(6517) <= a and b;
    layer1_outputs(6518) <= a and not b;
    layer1_outputs(6519) <= not b;
    layer1_outputs(6520) <= b and not a;
    layer1_outputs(6521) <= a xor b;
    layer1_outputs(6522) <= b and not a;
    layer1_outputs(6523) <= not b;
    layer1_outputs(6524) <= a or b;
    layer1_outputs(6525) <= not b or a;
    layer1_outputs(6526) <= not b or a;
    layer1_outputs(6527) <= a or b;
    layer1_outputs(6528) <= a or b;
    layer1_outputs(6529) <= not b or a;
    layer1_outputs(6530) <= not a;
    layer1_outputs(6531) <= a xor b;
    layer1_outputs(6532) <= not b or a;
    layer1_outputs(6533) <= a or b;
    layer1_outputs(6534) <= a or b;
    layer1_outputs(6535) <= not a;
    layer1_outputs(6536) <= not b;
    layer1_outputs(6537) <= not a or b;
    layer1_outputs(6538) <= a;
    layer1_outputs(6539) <= a or b;
    layer1_outputs(6540) <= a xor b;
    layer1_outputs(6541) <= not b or a;
    layer1_outputs(6542) <= not (a and b);
    layer1_outputs(6543) <= not a or b;
    layer1_outputs(6544) <= not b;
    layer1_outputs(6545) <= not (a or b);
    layer1_outputs(6546) <= not (a and b);
    layer1_outputs(6547) <= a and not b;
    layer1_outputs(6548) <= b;
    layer1_outputs(6549) <= a and b;
    layer1_outputs(6550) <= not a or b;
    layer1_outputs(6551) <= a xor b;
    layer1_outputs(6552) <= not a;
    layer1_outputs(6553) <= not (a xor b);
    layer1_outputs(6554) <= b;
    layer1_outputs(6555) <= not (a xor b);
    layer1_outputs(6556) <= a;
    layer1_outputs(6557) <= a xor b;
    layer1_outputs(6558) <= b and not a;
    layer1_outputs(6559) <= a xor b;
    layer1_outputs(6560) <= a;
    layer1_outputs(6561) <= not b;
    layer1_outputs(6562) <= b and not a;
    layer1_outputs(6563) <= not (a or b);
    layer1_outputs(6564) <= not a;
    layer1_outputs(6565) <= not (a xor b);
    layer1_outputs(6566) <= not (a and b);
    layer1_outputs(6567) <= a and b;
    layer1_outputs(6568) <= not (a or b);
    layer1_outputs(6569) <= a or b;
    layer1_outputs(6570) <= b;
    layer1_outputs(6571) <= a xor b;
    layer1_outputs(6572) <= not (a xor b);
    layer1_outputs(6573) <= b and not a;
    layer1_outputs(6574) <= b and not a;
    layer1_outputs(6575) <= not b or a;
    layer1_outputs(6576) <= not (a and b);
    layer1_outputs(6577) <= 1'b0;
    layer1_outputs(6578) <= not a;
    layer1_outputs(6579) <= b;
    layer1_outputs(6580) <= not b or a;
    layer1_outputs(6581) <= not b;
    layer1_outputs(6582) <= a and b;
    layer1_outputs(6583) <= 1'b0;
    layer1_outputs(6584) <= b;
    layer1_outputs(6585) <= a and b;
    layer1_outputs(6586) <= a and not b;
    layer1_outputs(6587) <= a;
    layer1_outputs(6588) <= a and b;
    layer1_outputs(6589) <= not a;
    layer1_outputs(6590) <= 1'b0;
    layer1_outputs(6591) <= a xor b;
    layer1_outputs(6592) <= a and not b;
    layer1_outputs(6593) <= a and b;
    layer1_outputs(6594) <= a or b;
    layer1_outputs(6595) <= a;
    layer1_outputs(6596) <= not (a and b);
    layer1_outputs(6597) <= not a or b;
    layer1_outputs(6598) <= a or b;
    layer1_outputs(6599) <= a;
    layer1_outputs(6600) <= not (a xor b);
    layer1_outputs(6601) <= b and not a;
    layer1_outputs(6602) <= not a;
    layer1_outputs(6603) <= a or b;
    layer1_outputs(6604) <= not (a or b);
    layer1_outputs(6605) <= a xor b;
    layer1_outputs(6606) <= a;
    layer1_outputs(6607) <= not a or b;
    layer1_outputs(6608) <= b and not a;
    layer1_outputs(6609) <= not (a xor b);
    layer1_outputs(6610) <= not b;
    layer1_outputs(6611) <= not (a and b);
    layer1_outputs(6612) <= a;
    layer1_outputs(6613) <= a and b;
    layer1_outputs(6614) <= a or b;
    layer1_outputs(6615) <= a xor b;
    layer1_outputs(6616) <= b;
    layer1_outputs(6617) <= not b;
    layer1_outputs(6618) <= not (a xor b);
    layer1_outputs(6619) <= a and not b;
    layer1_outputs(6620) <= b;
    layer1_outputs(6621) <= not b or a;
    layer1_outputs(6622) <= b;
    layer1_outputs(6623) <= not (a and b);
    layer1_outputs(6624) <= not a;
    layer1_outputs(6625) <= not (a or b);
    layer1_outputs(6626) <= not b;
    layer1_outputs(6627) <= not (a xor b);
    layer1_outputs(6628) <= a;
    layer1_outputs(6629) <= a and b;
    layer1_outputs(6630) <= not b or a;
    layer1_outputs(6631) <= not a or b;
    layer1_outputs(6632) <= not a or b;
    layer1_outputs(6633) <= not a;
    layer1_outputs(6634) <= b and not a;
    layer1_outputs(6635) <= a;
    layer1_outputs(6636) <= a xor b;
    layer1_outputs(6637) <= a xor b;
    layer1_outputs(6638) <= not b;
    layer1_outputs(6639) <= a xor b;
    layer1_outputs(6640) <= a;
    layer1_outputs(6641) <= a;
    layer1_outputs(6642) <= not b;
    layer1_outputs(6643) <= not (a or b);
    layer1_outputs(6644) <= a xor b;
    layer1_outputs(6645) <= a or b;
    layer1_outputs(6646) <= not (a xor b);
    layer1_outputs(6647) <= a and b;
    layer1_outputs(6648) <= not a;
    layer1_outputs(6649) <= not (a and b);
    layer1_outputs(6650) <= not a or b;
    layer1_outputs(6651) <= b;
    layer1_outputs(6652) <= not b;
    layer1_outputs(6653) <= not (a xor b);
    layer1_outputs(6654) <= not b;
    layer1_outputs(6655) <= a;
    layer1_outputs(6656) <= not b;
    layer1_outputs(6657) <= not (a and b);
    layer1_outputs(6658) <= not b;
    layer1_outputs(6659) <= a;
    layer1_outputs(6660) <= not (a or b);
    layer1_outputs(6661) <= not (a xor b);
    layer1_outputs(6662) <= not (a and b);
    layer1_outputs(6663) <= a;
    layer1_outputs(6664) <= b and not a;
    layer1_outputs(6665) <= a or b;
    layer1_outputs(6666) <= not (a or b);
    layer1_outputs(6667) <= a xor b;
    layer1_outputs(6668) <= not (a or b);
    layer1_outputs(6669) <= a;
    layer1_outputs(6670) <= not (a and b);
    layer1_outputs(6671) <= not b or a;
    layer1_outputs(6672) <= not a or b;
    layer1_outputs(6673) <= b and not a;
    layer1_outputs(6674) <= not b;
    layer1_outputs(6675) <= not (a or b);
    layer1_outputs(6676) <= not b or a;
    layer1_outputs(6677) <= not (a xor b);
    layer1_outputs(6678) <= not (a or b);
    layer1_outputs(6679) <= a xor b;
    layer1_outputs(6680) <= b and not a;
    layer1_outputs(6681) <= a xor b;
    layer1_outputs(6682) <= a;
    layer1_outputs(6683) <= not (a xor b);
    layer1_outputs(6684) <= not (a and b);
    layer1_outputs(6685) <= not (a or b);
    layer1_outputs(6686) <= a xor b;
    layer1_outputs(6687) <= a;
    layer1_outputs(6688) <= a;
    layer1_outputs(6689) <= not b;
    layer1_outputs(6690) <= b and not a;
    layer1_outputs(6691) <= not a;
    layer1_outputs(6692) <= b;
    layer1_outputs(6693) <= not (a or b);
    layer1_outputs(6694) <= a or b;
    layer1_outputs(6695) <= a xor b;
    layer1_outputs(6696) <= not a;
    layer1_outputs(6697) <= a xor b;
    layer1_outputs(6698) <= a and not b;
    layer1_outputs(6699) <= not b;
    layer1_outputs(6700) <= not a;
    layer1_outputs(6701) <= not b;
    layer1_outputs(6702) <= b and not a;
    layer1_outputs(6703) <= a or b;
    layer1_outputs(6704) <= a and b;
    layer1_outputs(6705) <= a or b;
    layer1_outputs(6706) <= b and not a;
    layer1_outputs(6707) <= a and not b;
    layer1_outputs(6708) <= b;
    layer1_outputs(6709) <= b and not a;
    layer1_outputs(6710) <= b;
    layer1_outputs(6711) <= a xor b;
    layer1_outputs(6712) <= not b or a;
    layer1_outputs(6713) <= not (a or b);
    layer1_outputs(6714) <= a xor b;
    layer1_outputs(6715) <= a or b;
    layer1_outputs(6716) <= not a;
    layer1_outputs(6717) <= a xor b;
    layer1_outputs(6718) <= a;
    layer1_outputs(6719) <= b;
    layer1_outputs(6720) <= a xor b;
    layer1_outputs(6721) <= not (a xor b);
    layer1_outputs(6722) <= not a or b;
    layer1_outputs(6723) <= not (a xor b);
    layer1_outputs(6724) <= not a or b;
    layer1_outputs(6725) <= not (a and b);
    layer1_outputs(6726) <= a and not b;
    layer1_outputs(6727) <= a xor b;
    layer1_outputs(6728) <= b;
    layer1_outputs(6729) <= a and b;
    layer1_outputs(6730) <= a;
    layer1_outputs(6731) <= not (a xor b);
    layer1_outputs(6732) <= a xor b;
    layer1_outputs(6733) <= not b;
    layer1_outputs(6734) <= a and not b;
    layer1_outputs(6735) <= not (a or b);
    layer1_outputs(6736) <= not (a xor b);
    layer1_outputs(6737) <= not (a or b);
    layer1_outputs(6738) <= a;
    layer1_outputs(6739) <= not b;
    layer1_outputs(6740) <= b and not a;
    layer1_outputs(6741) <= not b;
    layer1_outputs(6742) <= b;
    layer1_outputs(6743) <= not b;
    layer1_outputs(6744) <= b and not a;
    layer1_outputs(6745) <= not a or b;
    layer1_outputs(6746) <= a or b;
    layer1_outputs(6747) <= not b;
    layer1_outputs(6748) <= not b;
    layer1_outputs(6749) <= not a;
    layer1_outputs(6750) <= a and b;
    layer1_outputs(6751) <= not b;
    layer1_outputs(6752) <= not a or b;
    layer1_outputs(6753) <= not (a and b);
    layer1_outputs(6754) <= not (a xor b);
    layer1_outputs(6755) <= not a;
    layer1_outputs(6756) <= not (a or b);
    layer1_outputs(6757) <= a or b;
    layer1_outputs(6758) <= a;
    layer1_outputs(6759) <= b;
    layer1_outputs(6760) <= not b or a;
    layer1_outputs(6761) <= not b or a;
    layer1_outputs(6762) <= a;
    layer1_outputs(6763) <= not (a and b);
    layer1_outputs(6764) <= not (a or b);
    layer1_outputs(6765) <= a and b;
    layer1_outputs(6766) <= b;
    layer1_outputs(6767) <= a;
    layer1_outputs(6768) <= b;
    layer1_outputs(6769) <= not (a xor b);
    layer1_outputs(6770) <= not a or b;
    layer1_outputs(6771) <= a and not b;
    layer1_outputs(6772) <= a or b;
    layer1_outputs(6773) <= a;
    layer1_outputs(6774) <= not b or a;
    layer1_outputs(6775) <= a;
    layer1_outputs(6776) <= b and not a;
    layer1_outputs(6777) <= a or b;
    layer1_outputs(6778) <= b and not a;
    layer1_outputs(6779) <= b;
    layer1_outputs(6780) <= not b;
    layer1_outputs(6781) <= not (a and b);
    layer1_outputs(6782) <= b and not a;
    layer1_outputs(6783) <= b;
    layer1_outputs(6784) <= a and b;
    layer1_outputs(6785) <= not b;
    layer1_outputs(6786) <= a or b;
    layer1_outputs(6787) <= a;
    layer1_outputs(6788) <= a or b;
    layer1_outputs(6789) <= a and not b;
    layer1_outputs(6790) <= b and not a;
    layer1_outputs(6791) <= not b;
    layer1_outputs(6792) <= not a or b;
    layer1_outputs(6793) <= not a or b;
    layer1_outputs(6794) <= not (a or b);
    layer1_outputs(6795) <= a or b;
    layer1_outputs(6796) <= a and not b;
    layer1_outputs(6797) <= a;
    layer1_outputs(6798) <= a xor b;
    layer1_outputs(6799) <= not a;
    layer1_outputs(6800) <= not (a or b);
    layer1_outputs(6801) <= a or b;
    layer1_outputs(6802) <= not b;
    layer1_outputs(6803) <= not a;
    layer1_outputs(6804) <= a or b;
    layer1_outputs(6805) <= b;
    layer1_outputs(6806) <= b;
    layer1_outputs(6807) <= a or b;
    layer1_outputs(6808) <= not b or a;
    layer1_outputs(6809) <= not b;
    layer1_outputs(6810) <= b;
    layer1_outputs(6811) <= not a;
    layer1_outputs(6812) <= b and not a;
    layer1_outputs(6813) <= not (a xor b);
    layer1_outputs(6814) <= not b;
    layer1_outputs(6815) <= a and not b;
    layer1_outputs(6816) <= a xor b;
    layer1_outputs(6817) <= not (a xor b);
    layer1_outputs(6818) <= a and b;
    layer1_outputs(6819) <= not a or b;
    layer1_outputs(6820) <= not (a or b);
    layer1_outputs(6821) <= a xor b;
    layer1_outputs(6822) <= not a;
    layer1_outputs(6823) <= a;
    layer1_outputs(6824) <= a;
    layer1_outputs(6825) <= 1'b1;
    layer1_outputs(6826) <= not b;
    layer1_outputs(6827) <= not a;
    layer1_outputs(6828) <= not a or b;
    layer1_outputs(6829) <= a;
    layer1_outputs(6830) <= a;
    layer1_outputs(6831) <= a and b;
    layer1_outputs(6832) <= not (a xor b);
    layer1_outputs(6833) <= not b;
    layer1_outputs(6834) <= not (a and b);
    layer1_outputs(6835) <= not a;
    layer1_outputs(6836) <= not a;
    layer1_outputs(6837) <= not b;
    layer1_outputs(6838) <= a or b;
    layer1_outputs(6839) <= not (a or b);
    layer1_outputs(6840) <= not a or b;
    layer1_outputs(6841) <= b and not a;
    layer1_outputs(6842) <= not (a or b);
    layer1_outputs(6843) <= not (a and b);
    layer1_outputs(6844) <= b and not a;
    layer1_outputs(6845) <= b;
    layer1_outputs(6846) <= b;
    layer1_outputs(6847) <= 1'b0;
    layer1_outputs(6848) <= a;
    layer1_outputs(6849) <= a;
    layer1_outputs(6850) <= a and not b;
    layer1_outputs(6851) <= a and not b;
    layer1_outputs(6852) <= not (a xor b);
    layer1_outputs(6853) <= b and not a;
    layer1_outputs(6854) <= not a;
    layer1_outputs(6855) <= not a;
    layer1_outputs(6856) <= not b or a;
    layer1_outputs(6857) <= a and not b;
    layer1_outputs(6858) <= not (a and b);
    layer1_outputs(6859) <= a;
    layer1_outputs(6860) <= not (a and b);
    layer1_outputs(6861) <= a;
    layer1_outputs(6862) <= not b;
    layer1_outputs(6863) <= a or b;
    layer1_outputs(6864) <= not a or b;
    layer1_outputs(6865) <= a;
    layer1_outputs(6866) <= not b;
    layer1_outputs(6867) <= not b;
    layer1_outputs(6868) <= not (a and b);
    layer1_outputs(6869) <= a or b;
    layer1_outputs(6870) <= b and not a;
    layer1_outputs(6871) <= not (a xor b);
    layer1_outputs(6872) <= a;
    layer1_outputs(6873) <= not (a xor b);
    layer1_outputs(6874) <= not a;
    layer1_outputs(6875) <= b;
    layer1_outputs(6876) <= a and b;
    layer1_outputs(6877) <= a and b;
    layer1_outputs(6878) <= not (a and b);
    layer1_outputs(6879) <= a;
    layer1_outputs(6880) <= not b;
    layer1_outputs(6881) <= b;
    layer1_outputs(6882) <= not a;
    layer1_outputs(6883) <= not a or b;
    layer1_outputs(6884) <= not (a or b);
    layer1_outputs(6885) <= not (a or b);
    layer1_outputs(6886) <= b and not a;
    layer1_outputs(6887) <= a or b;
    layer1_outputs(6888) <= b;
    layer1_outputs(6889) <= not (a xor b);
    layer1_outputs(6890) <= a xor b;
    layer1_outputs(6891) <= b and not a;
    layer1_outputs(6892) <= a;
    layer1_outputs(6893) <= not (a xor b);
    layer1_outputs(6894) <= b;
    layer1_outputs(6895) <= not a;
    layer1_outputs(6896) <= not (a xor b);
    layer1_outputs(6897) <= a;
    layer1_outputs(6898) <= not b or a;
    layer1_outputs(6899) <= a xor b;
    layer1_outputs(6900) <= a and b;
    layer1_outputs(6901) <= a or b;
    layer1_outputs(6902) <= not a or b;
    layer1_outputs(6903) <= a and not b;
    layer1_outputs(6904) <= a or b;
    layer1_outputs(6905) <= 1'b1;
    layer1_outputs(6906) <= not b;
    layer1_outputs(6907) <= b;
    layer1_outputs(6908) <= not a;
    layer1_outputs(6909) <= a and not b;
    layer1_outputs(6910) <= not (a xor b);
    layer1_outputs(6911) <= not (a xor b);
    layer1_outputs(6912) <= b and not a;
    layer1_outputs(6913) <= a;
    layer1_outputs(6914) <= not a;
    layer1_outputs(6915) <= a and not b;
    layer1_outputs(6916) <= not (a or b);
    layer1_outputs(6917) <= not (a xor b);
    layer1_outputs(6918) <= not (a xor b);
    layer1_outputs(6919) <= b and not a;
    layer1_outputs(6920) <= a xor b;
    layer1_outputs(6921) <= not a;
    layer1_outputs(6922) <= b;
    layer1_outputs(6923) <= not (a xor b);
    layer1_outputs(6924) <= a and b;
    layer1_outputs(6925) <= not b;
    layer1_outputs(6926) <= not a;
    layer1_outputs(6927) <= not b or a;
    layer1_outputs(6928) <= a or b;
    layer1_outputs(6929) <= not (a and b);
    layer1_outputs(6930) <= a and b;
    layer1_outputs(6931) <= not a;
    layer1_outputs(6932) <= a and not b;
    layer1_outputs(6933) <= not a;
    layer1_outputs(6934) <= a;
    layer1_outputs(6935) <= b and not a;
    layer1_outputs(6936) <= b and not a;
    layer1_outputs(6937) <= a;
    layer1_outputs(6938) <= a;
    layer1_outputs(6939) <= b;
    layer1_outputs(6940) <= a;
    layer1_outputs(6941) <= a;
    layer1_outputs(6942) <= not a;
    layer1_outputs(6943) <= not a or b;
    layer1_outputs(6944) <= not b;
    layer1_outputs(6945) <= a and b;
    layer1_outputs(6946) <= not b or a;
    layer1_outputs(6947) <= a xor b;
    layer1_outputs(6948) <= not (a xor b);
    layer1_outputs(6949) <= not b or a;
    layer1_outputs(6950) <= not a;
    layer1_outputs(6951) <= not a or b;
    layer1_outputs(6952) <= not a or b;
    layer1_outputs(6953) <= a xor b;
    layer1_outputs(6954) <= not (a xor b);
    layer1_outputs(6955) <= not a;
    layer1_outputs(6956) <= not b or a;
    layer1_outputs(6957) <= not (a or b);
    layer1_outputs(6958) <= not (a xor b);
    layer1_outputs(6959) <= a and not b;
    layer1_outputs(6960) <= not b or a;
    layer1_outputs(6961) <= not (a or b);
    layer1_outputs(6962) <= not b or a;
    layer1_outputs(6963) <= a xor b;
    layer1_outputs(6964) <= a and not b;
    layer1_outputs(6965) <= not (a or b);
    layer1_outputs(6966) <= not (a xor b);
    layer1_outputs(6967) <= not (a and b);
    layer1_outputs(6968) <= not a or b;
    layer1_outputs(6969) <= not (a or b);
    layer1_outputs(6970) <= not b or a;
    layer1_outputs(6971) <= not a or b;
    layer1_outputs(6972) <= b and not a;
    layer1_outputs(6973) <= a;
    layer1_outputs(6974) <= not b;
    layer1_outputs(6975) <= 1'b1;
    layer1_outputs(6976) <= 1'b0;
    layer1_outputs(6977) <= b;
    layer1_outputs(6978) <= b and not a;
    layer1_outputs(6979) <= a or b;
    layer1_outputs(6980) <= not (a or b);
    layer1_outputs(6981) <= b and not a;
    layer1_outputs(6982) <= not (a or b);
    layer1_outputs(6983) <= not b;
    layer1_outputs(6984) <= not (a xor b);
    layer1_outputs(6985) <= not b or a;
    layer1_outputs(6986) <= a xor b;
    layer1_outputs(6987) <= a;
    layer1_outputs(6988) <= 1'b0;
    layer1_outputs(6989) <= a and not b;
    layer1_outputs(6990) <= not (a xor b);
    layer1_outputs(6991) <= not a;
    layer1_outputs(6992) <= b and not a;
    layer1_outputs(6993) <= b and not a;
    layer1_outputs(6994) <= b;
    layer1_outputs(6995) <= b and not a;
    layer1_outputs(6996) <= not (a xor b);
    layer1_outputs(6997) <= not a;
    layer1_outputs(6998) <= not (a or b);
    layer1_outputs(6999) <= not a;
    layer1_outputs(7000) <= not a;
    layer1_outputs(7001) <= not b;
    layer1_outputs(7002) <= not (a xor b);
    layer1_outputs(7003) <= not (a xor b);
    layer1_outputs(7004) <= not a;
    layer1_outputs(7005) <= not (a and b);
    layer1_outputs(7006) <= a or b;
    layer1_outputs(7007) <= not a;
    layer1_outputs(7008) <= a xor b;
    layer1_outputs(7009) <= a xor b;
    layer1_outputs(7010) <= not (a or b);
    layer1_outputs(7011) <= not (a xor b);
    layer1_outputs(7012) <= b and not a;
    layer1_outputs(7013) <= not b or a;
    layer1_outputs(7014) <= a or b;
    layer1_outputs(7015) <= a and b;
    layer1_outputs(7016) <= not (a xor b);
    layer1_outputs(7017) <= b and not a;
    layer1_outputs(7018) <= not (a xor b);
    layer1_outputs(7019) <= b and not a;
    layer1_outputs(7020) <= a;
    layer1_outputs(7021) <= not a;
    layer1_outputs(7022) <= not (a and b);
    layer1_outputs(7023) <= a or b;
    layer1_outputs(7024) <= 1'b1;
    layer1_outputs(7025) <= 1'b1;
    layer1_outputs(7026) <= not a;
    layer1_outputs(7027) <= a and not b;
    layer1_outputs(7028) <= b and not a;
    layer1_outputs(7029) <= a xor b;
    layer1_outputs(7030) <= b;
    layer1_outputs(7031) <= not a;
    layer1_outputs(7032) <= a;
    layer1_outputs(7033) <= b and not a;
    layer1_outputs(7034) <= a and not b;
    layer1_outputs(7035) <= not (a xor b);
    layer1_outputs(7036) <= not a or b;
    layer1_outputs(7037) <= a or b;
    layer1_outputs(7038) <= not a;
    layer1_outputs(7039) <= not b;
    layer1_outputs(7040) <= a xor b;
    layer1_outputs(7041) <= not a;
    layer1_outputs(7042) <= not (a xor b);
    layer1_outputs(7043) <= a;
    layer1_outputs(7044) <= a;
    layer1_outputs(7045) <= not (a or b);
    layer1_outputs(7046) <= not (a or b);
    layer1_outputs(7047) <= not b or a;
    layer1_outputs(7048) <= a or b;
    layer1_outputs(7049) <= not a or b;
    layer1_outputs(7050) <= not a;
    layer1_outputs(7051) <= not (a and b);
    layer1_outputs(7052) <= a xor b;
    layer1_outputs(7053) <= not a;
    layer1_outputs(7054) <= not b;
    layer1_outputs(7055) <= b and not a;
    layer1_outputs(7056) <= not (a xor b);
    layer1_outputs(7057) <= a or b;
    layer1_outputs(7058) <= not b;
    layer1_outputs(7059) <= not b;
    layer1_outputs(7060) <= not b;
    layer1_outputs(7061) <= 1'b0;
    layer1_outputs(7062) <= a and b;
    layer1_outputs(7063) <= not b;
    layer1_outputs(7064) <= a and b;
    layer1_outputs(7065) <= a or b;
    layer1_outputs(7066) <= not b or a;
    layer1_outputs(7067) <= not a or b;
    layer1_outputs(7068) <= a xor b;
    layer1_outputs(7069) <= a;
    layer1_outputs(7070) <= a;
    layer1_outputs(7071) <= not (a and b);
    layer1_outputs(7072) <= a and b;
    layer1_outputs(7073) <= a or b;
    layer1_outputs(7074) <= a xor b;
    layer1_outputs(7075) <= not a;
    layer1_outputs(7076) <= not a;
    layer1_outputs(7077) <= a xor b;
    layer1_outputs(7078) <= a;
    layer1_outputs(7079) <= not a;
    layer1_outputs(7080) <= not (a or b);
    layer1_outputs(7081) <= b;
    layer1_outputs(7082) <= not (a or b);
    layer1_outputs(7083) <= not a or b;
    layer1_outputs(7084) <= not (a xor b);
    layer1_outputs(7085) <= b and not a;
    layer1_outputs(7086) <= b and not a;
    layer1_outputs(7087) <= b;
    layer1_outputs(7088) <= a xor b;
    layer1_outputs(7089) <= b and not a;
    layer1_outputs(7090) <= not a;
    layer1_outputs(7091) <= not a or b;
    layer1_outputs(7092) <= not (a and b);
    layer1_outputs(7093) <= not a or b;
    layer1_outputs(7094) <= not b or a;
    layer1_outputs(7095) <= b;
    layer1_outputs(7096) <= a xor b;
    layer1_outputs(7097) <= not b or a;
    layer1_outputs(7098) <= a;
    layer1_outputs(7099) <= b and not a;
    layer1_outputs(7100) <= b and not a;
    layer1_outputs(7101) <= b;
    layer1_outputs(7102) <= not a;
    layer1_outputs(7103) <= a;
    layer1_outputs(7104) <= not a;
    layer1_outputs(7105) <= a and not b;
    layer1_outputs(7106) <= a or b;
    layer1_outputs(7107) <= not (a xor b);
    layer1_outputs(7108) <= not (a and b);
    layer1_outputs(7109) <= not b;
    layer1_outputs(7110) <= a and b;
    layer1_outputs(7111) <= not (a xor b);
    layer1_outputs(7112) <= not (a xor b);
    layer1_outputs(7113) <= b;
    layer1_outputs(7114) <= not (a xor b);
    layer1_outputs(7115) <= not (a or b);
    layer1_outputs(7116) <= not a or b;
    layer1_outputs(7117) <= not b;
    layer1_outputs(7118) <= b and not a;
    layer1_outputs(7119) <= a and not b;
    layer1_outputs(7120) <= a;
    layer1_outputs(7121) <= a or b;
    layer1_outputs(7122) <= not b;
    layer1_outputs(7123) <= not (a or b);
    layer1_outputs(7124) <= b;
    layer1_outputs(7125) <= a or b;
    layer1_outputs(7126) <= a or b;
    layer1_outputs(7127) <= not b;
    layer1_outputs(7128) <= not a;
    layer1_outputs(7129) <= not b;
    layer1_outputs(7130) <= not (a xor b);
    layer1_outputs(7131) <= not a;
    layer1_outputs(7132) <= not (a or b);
    layer1_outputs(7133) <= not a;
    layer1_outputs(7134) <= a xor b;
    layer1_outputs(7135) <= not (a or b);
    layer1_outputs(7136) <= b;
    layer1_outputs(7137) <= b;
    layer1_outputs(7138) <= not a or b;
    layer1_outputs(7139) <= a;
    layer1_outputs(7140) <= a or b;
    layer1_outputs(7141) <= b and not a;
    layer1_outputs(7142) <= not (a or b);
    layer1_outputs(7143) <= not (a and b);
    layer1_outputs(7144) <= not (a xor b);
    layer1_outputs(7145) <= not b;
    layer1_outputs(7146) <= b and not a;
    layer1_outputs(7147) <= not a or b;
    layer1_outputs(7148) <= 1'b1;
    layer1_outputs(7149) <= not (a xor b);
    layer1_outputs(7150) <= not a;
    layer1_outputs(7151) <= a;
    layer1_outputs(7152) <= b;
    layer1_outputs(7153) <= not (a xor b);
    layer1_outputs(7154) <= b;
    layer1_outputs(7155) <= not (a xor b);
    layer1_outputs(7156) <= not a;
    layer1_outputs(7157) <= not a;
    layer1_outputs(7158) <= not a;
    layer1_outputs(7159) <= not a or b;
    layer1_outputs(7160) <= not (a and b);
    layer1_outputs(7161) <= not b;
    layer1_outputs(7162) <= not (a xor b);
    layer1_outputs(7163) <= b and not a;
    layer1_outputs(7164) <= a and b;
    layer1_outputs(7165) <= b and not a;
    layer1_outputs(7166) <= not a or b;
    layer1_outputs(7167) <= not (a and b);
    layer1_outputs(7168) <= a xor b;
    layer1_outputs(7169) <= b and not a;
    layer1_outputs(7170) <= b and not a;
    layer1_outputs(7171) <= a xor b;
    layer1_outputs(7172) <= a or b;
    layer1_outputs(7173) <= not (a xor b);
    layer1_outputs(7174) <= a xor b;
    layer1_outputs(7175) <= a and b;
    layer1_outputs(7176) <= b;
    layer1_outputs(7177) <= not (a xor b);
    layer1_outputs(7178) <= not b;
    layer1_outputs(7179) <= a xor b;
    layer1_outputs(7180) <= b and not a;
    layer1_outputs(7181) <= a or b;
    layer1_outputs(7182) <= a or b;
    layer1_outputs(7183) <= a;
    layer1_outputs(7184) <= b and not a;
    layer1_outputs(7185) <= a or b;
    layer1_outputs(7186) <= a or b;
    layer1_outputs(7187) <= not (a or b);
    layer1_outputs(7188) <= b and not a;
    layer1_outputs(7189) <= a;
    layer1_outputs(7190) <= a;
    layer1_outputs(7191) <= a and not b;
    layer1_outputs(7192) <= a and b;
    layer1_outputs(7193) <= a xor b;
    layer1_outputs(7194) <= not b;
    layer1_outputs(7195) <= b and not a;
    layer1_outputs(7196) <= not b;
    layer1_outputs(7197) <= a;
    layer1_outputs(7198) <= not (a and b);
    layer1_outputs(7199) <= not (a xor b);
    layer1_outputs(7200) <= not b or a;
    layer1_outputs(7201) <= not (a and b);
    layer1_outputs(7202) <= not b;
    layer1_outputs(7203) <= not b or a;
    layer1_outputs(7204) <= a and not b;
    layer1_outputs(7205) <= not (a and b);
    layer1_outputs(7206) <= not a;
    layer1_outputs(7207) <= b;
    layer1_outputs(7208) <= not b;
    layer1_outputs(7209) <= b and not a;
    layer1_outputs(7210) <= a and not b;
    layer1_outputs(7211) <= not b;
    layer1_outputs(7212) <= b;
    layer1_outputs(7213) <= not a or b;
    layer1_outputs(7214) <= b;
    layer1_outputs(7215) <= a and not b;
    layer1_outputs(7216) <= not a or b;
    layer1_outputs(7217) <= a xor b;
    layer1_outputs(7218) <= not b;
    layer1_outputs(7219) <= not (a and b);
    layer1_outputs(7220) <= not a;
    layer1_outputs(7221) <= not a;
    layer1_outputs(7222) <= not a;
    layer1_outputs(7223) <= not (a xor b);
    layer1_outputs(7224) <= not b;
    layer1_outputs(7225) <= a or b;
    layer1_outputs(7226) <= a;
    layer1_outputs(7227) <= not a;
    layer1_outputs(7228) <= a or b;
    layer1_outputs(7229) <= a xor b;
    layer1_outputs(7230) <= a or b;
    layer1_outputs(7231) <= 1'b1;
    layer1_outputs(7232) <= not a or b;
    layer1_outputs(7233) <= not (a or b);
    layer1_outputs(7234) <= not b;
    layer1_outputs(7235) <= b;
    layer1_outputs(7236) <= not b or a;
    layer1_outputs(7237) <= not b;
    layer1_outputs(7238) <= b;
    layer1_outputs(7239) <= a and not b;
    layer1_outputs(7240) <= not a;
    layer1_outputs(7241) <= not (a or b);
    layer1_outputs(7242) <= not (a xor b);
    layer1_outputs(7243) <= not a or b;
    layer1_outputs(7244) <= not b;
    layer1_outputs(7245) <= not a or b;
    layer1_outputs(7246) <= a and b;
    layer1_outputs(7247) <= not a;
    layer1_outputs(7248) <= a xor b;
    layer1_outputs(7249) <= not b;
    layer1_outputs(7250) <= not a;
    layer1_outputs(7251) <= not (a xor b);
    layer1_outputs(7252) <= a;
    layer1_outputs(7253) <= a or b;
    layer1_outputs(7254) <= a or b;
    layer1_outputs(7255) <= a;
    layer1_outputs(7256) <= not (a or b);
    layer1_outputs(7257) <= b and not a;
    layer1_outputs(7258) <= not (a or b);
    layer1_outputs(7259) <= not (a or b);
    layer1_outputs(7260) <= a and b;
    layer1_outputs(7261) <= b;
    layer1_outputs(7262) <= b;
    layer1_outputs(7263) <= b and not a;
    layer1_outputs(7264) <= not (a or b);
    layer1_outputs(7265) <= a or b;
    layer1_outputs(7266) <= not a;
    layer1_outputs(7267) <= 1'b0;
    layer1_outputs(7268) <= a;
    layer1_outputs(7269) <= b;
    layer1_outputs(7270) <= a and not b;
    layer1_outputs(7271) <= a and not b;
    layer1_outputs(7272) <= a xor b;
    layer1_outputs(7273) <= not (a xor b);
    layer1_outputs(7274) <= a;
    layer1_outputs(7275) <= not b;
    layer1_outputs(7276) <= not (a and b);
    layer1_outputs(7277) <= not a;
    layer1_outputs(7278) <= not (a or b);
    layer1_outputs(7279) <= a;
    layer1_outputs(7280) <= not a or b;
    layer1_outputs(7281) <= a and not b;
    layer1_outputs(7282) <= not a;
    layer1_outputs(7283) <= not b;
    layer1_outputs(7284) <= not b;
    layer1_outputs(7285) <= not b;
    layer1_outputs(7286) <= not b or a;
    layer1_outputs(7287) <= a;
    layer1_outputs(7288) <= a xor b;
    layer1_outputs(7289) <= not a or b;
    layer1_outputs(7290) <= not b or a;
    layer1_outputs(7291) <= not (a and b);
    layer1_outputs(7292) <= not a or b;
    layer1_outputs(7293) <= b and not a;
    layer1_outputs(7294) <= not b or a;
    layer1_outputs(7295) <= a and b;
    layer1_outputs(7296) <= b;
    layer1_outputs(7297) <= not a;
    layer1_outputs(7298) <= 1'b0;
    layer1_outputs(7299) <= b;
    layer1_outputs(7300) <= a and not b;
    layer1_outputs(7301) <= not (a xor b);
    layer1_outputs(7302) <= b;
    layer1_outputs(7303) <= a;
    layer1_outputs(7304) <= b;
    layer1_outputs(7305) <= not a or b;
    layer1_outputs(7306) <= b;
    layer1_outputs(7307) <= a;
    layer1_outputs(7308) <= a or b;
    layer1_outputs(7309) <= a xor b;
    layer1_outputs(7310) <= not b;
    layer1_outputs(7311) <= b and not a;
    layer1_outputs(7312) <= not (a and b);
    layer1_outputs(7313) <= not (a xor b);
    layer1_outputs(7314) <= not (a xor b);
    layer1_outputs(7315) <= a xor b;
    layer1_outputs(7316) <= not (a xor b);
    layer1_outputs(7317) <= b;
    layer1_outputs(7318) <= b;
    layer1_outputs(7319) <= not (a or b);
    layer1_outputs(7320) <= not a or b;
    layer1_outputs(7321) <= not a;
    layer1_outputs(7322) <= a;
    layer1_outputs(7323) <= not (a or b);
    layer1_outputs(7324) <= a and b;
    layer1_outputs(7325) <= not b;
    layer1_outputs(7326) <= not b;
    layer1_outputs(7327) <= a;
    layer1_outputs(7328) <= not (a and b);
    layer1_outputs(7329) <= not a or b;
    layer1_outputs(7330) <= not b;
    layer1_outputs(7331) <= not (a and b);
    layer1_outputs(7332) <= b;
    layer1_outputs(7333) <= a and b;
    layer1_outputs(7334) <= not b;
    layer1_outputs(7335) <= not b or a;
    layer1_outputs(7336) <= b and not a;
    layer1_outputs(7337) <= not b or a;
    layer1_outputs(7338) <= b;
    layer1_outputs(7339) <= a and not b;
    layer1_outputs(7340) <= not a;
    layer1_outputs(7341) <= a xor b;
    layer1_outputs(7342) <= a or b;
    layer1_outputs(7343) <= a and not b;
    layer1_outputs(7344) <= a;
    layer1_outputs(7345) <= not a;
    layer1_outputs(7346) <= 1'b1;
    layer1_outputs(7347) <= not (a or b);
    layer1_outputs(7348) <= not (a and b);
    layer1_outputs(7349) <= b;
    layer1_outputs(7350) <= not a or b;
    layer1_outputs(7351) <= b and not a;
    layer1_outputs(7352) <= a xor b;
    layer1_outputs(7353) <= not a;
    layer1_outputs(7354) <= not a;
    layer1_outputs(7355) <= not (a or b);
    layer1_outputs(7356) <= a;
    layer1_outputs(7357) <= a;
    layer1_outputs(7358) <= a or b;
    layer1_outputs(7359) <= b;
    layer1_outputs(7360) <= not b or a;
    layer1_outputs(7361) <= not a;
    layer1_outputs(7362) <= b;
    layer1_outputs(7363) <= b;
    layer1_outputs(7364) <= a and not b;
    layer1_outputs(7365) <= a xor b;
    layer1_outputs(7366) <= not (a or b);
    layer1_outputs(7367) <= a and not b;
    layer1_outputs(7368) <= a and b;
    layer1_outputs(7369) <= a and b;
    layer1_outputs(7370) <= a xor b;
    layer1_outputs(7371) <= not (a and b);
    layer1_outputs(7372) <= a and b;
    layer1_outputs(7373) <= not b;
    layer1_outputs(7374) <= not (a xor b);
    layer1_outputs(7375) <= not a;
    layer1_outputs(7376) <= a and not b;
    layer1_outputs(7377) <= a;
    layer1_outputs(7378) <= not b or a;
    layer1_outputs(7379) <= a;
    layer1_outputs(7380) <= not (a xor b);
    layer1_outputs(7381) <= a xor b;
    layer1_outputs(7382) <= not (a xor b);
    layer1_outputs(7383) <= a;
    layer1_outputs(7384) <= a;
    layer1_outputs(7385) <= a xor b;
    layer1_outputs(7386) <= not a or b;
    layer1_outputs(7387) <= not b or a;
    layer1_outputs(7388) <= not a;
    layer1_outputs(7389) <= not b or a;
    layer1_outputs(7390) <= a;
    layer1_outputs(7391) <= not b;
    layer1_outputs(7392) <= not (a xor b);
    layer1_outputs(7393) <= not a;
    layer1_outputs(7394) <= a;
    layer1_outputs(7395) <= not (a xor b);
    layer1_outputs(7396) <= a xor b;
    layer1_outputs(7397) <= not (a xor b);
    layer1_outputs(7398) <= not (a or b);
    layer1_outputs(7399) <= not (a and b);
    layer1_outputs(7400) <= a;
    layer1_outputs(7401) <= not b;
    layer1_outputs(7402) <= a;
    layer1_outputs(7403) <= b;
    layer1_outputs(7404) <= b and not a;
    layer1_outputs(7405) <= not b or a;
    layer1_outputs(7406) <= a or b;
    layer1_outputs(7407) <= a;
    layer1_outputs(7408) <= not (a and b);
    layer1_outputs(7409) <= b;
    layer1_outputs(7410) <= not a;
    layer1_outputs(7411) <= a;
    layer1_outputs(7412) <= b;
    layer1_outputs(7413) <= a xor b;
    layer1_outputs(7414) <= not b or a;
    layer1_outputs(7415) <= not a;
    layer1_outputs(7416) <= 1'b0;
    layer1_outputs(7417) <= a or b;
    layer1_outputs(7418) <= not b;
    layer1_outputs(7419) <= not a or b;
    layer1_outputs(7420) <= not a;
    layer1_outputs(7421) <= not a;
    layer1_outputs(7422) <= b;
    layer1_outputs(7423) <= b;
    layer1_outputs(7424) <= b and not a;
    layer1_outputs(7425) <= b and not a;
    layer1_outputs(7426) <= b and not a;
    layer1_outputs(7427) <= not (a or b);
    layer1_outputs(7428) <= not (a xor b);
    layer1_outputs(7429) <= b;
    layer1_outputs(7430) <= not (a or b);
    layer1_outputs(7431) <= not (a or b);
    layer1_outputs(7432) <= not b or a;
    layer1_outputs(7433) <= a;
    layer1_outputs(7434) <= a and not b;
    layer1_outputs(7435) <= 1'b1;
    layer1_outputs(7436) <= a or b;
    layer1_outputs(7437) <= not a;
    layer1_outputs(7438) <= a or b;
    layer1_outputs(7439) <= a;
    layer1_outputs(7440) <= a xor b;
    layer1_outputs(7441) <= 1'b0;
    layer1_outputs(7442) <= not b;
    layer1_outputs(7443) <= b;
    layer1_outputs(7444) <= a;
    layer1_outputs(7445) <= not (a and b);
    layer1_outputs(7446) <= a xor b;
    layer1_outputs(7447) <= not a or b;
    layer1_outputs(7448) <= a;
    layer1_outputs(7449) <= a xor b;
    layer1_outputs(7450) <= not (a and b);
    layer1_outputs(7451) <= a and not b;
    layer1_outputs(7452) <= a;
    layer1_outputs(7453) <= 1'b1;
    layer1_outputs(7454) <= not (a or b);
    layer1_outputs(7455) <= a or b;
    layer1_outputs(7456) <= not a or b;
    layer1_outputs(7457) <= not a;
    layer1_outputs(7458) <= not (a or b);
    layer1_outputs(7459) <= not b or a;
    layer1_outputs(7460) <= not (a or b);
    layer1_outputs(7461) <= not a;
    layer1_outputs(7462) <= a or b;
    layer1_outputs(7463) <= not (a and b);
    layer1_outputs(7464) <= a or b;
    layer1_outputs(7465) <= not (a and b);
    layer1_outputs(7466) <= not b;
    layer1_outputs(7467) <= not a;
    layer1_outputs(7468) <= a xor b;
    layer1_outputs(7469) <= b and not a;
    layer1_outputs(7470) <= a and b;
    layer1_outputs(7471) <= not (a or b);
    layer1_outputs(7472) <= not a;
    layer1_outputs(7473) <= b;
    layer1_outputs(7474) <= not (a and b);
    layer1_outputs(7475) <= a xor b;
    layer1_outputs(7476) <= not b or a;
    layer1_outputs(7477) <= not a;
    layer1_outputs(7478) <= not a or b;
    layer1_outputs(7479) <= not (a and b);
    layer1_outputs(7480) <= 1'b1;
    layer1_outputs(7481) <= not (a xor b);
    layer1_outputs(7482) <= not b;
    layer1_outputs(7483) <= a and not b;
    layer1_outputs(7484) <= not a;
    layer1_outputs(7485) <= b;
    layer1_outputs(7486) <= a xor b;
    layer1_outputs(7487) <= not b or a;
    layer1_outputs(7488) <= not b;
    layer1_outputs(7489) <= a;
    layer1_outputs(7490) <= not a;
    layer1_outputs(7491) <= b;
    layer1_outputs(7492) <= a or b;
    layer1_outputs(7493) <= not a;
    layer1_outputs(7494) <= not b or a;
    layer1_outputs(7495) <= not a;
    layer1_outputs(7496) <= b;
    layer1_outputs(7497) <= not (a or b);
    layer1_outputs(7498) <= not a;
    layer1_outputs(7499) <= b;
    layer1_outputs(7500) <= not a;
    layer1_outputs(7501) <= a and not b;
    layer1_outputs(7502) <= a and b;
    layer1_outputs(7503) <= a;
    layer1_outputs(7504) <= not a;
    layer1_outputs(7505) <= a and b;
    layer1_outputs(7506) <= not b or a;
    layer1_outputs(7507) <= not (a xor b);
    layer1_outputs(7508) <= not (a or b);
    layer1_outputs(7509) <= not b;
    layer1_outputs(7510) <= not (a and b);
    layer1_outputs(7511) <= 1'b1;
    layer1_outputs(7512) <= b and not a;
    layer1_outputs(7513) <= not a;
    layer1_outputs(7514) <= not a;
    layer1_outputs(7515) <= not b;
    layer1_outputs(7516) <= a xor b;
    layer1_outputs(7517) <= not a or b;
    layer1_outputs(7518) <= not (a or b);
    layer1_outputs(7519) <= a and b;
    layer1_outputs(7520) <= a and b;
    layer1_outputs(7521) <= a;
    layer1_outputs(7522) <= not (a or b);
    layer1_outputs(7523) <= not (a xor b);
    layer1_outputs(7524) <= 1'b0;
    layer1_outputs(7525) <= 1'b1;
    layer1_outputs(7526) <= not a;
    layer1_outputs(7527) <= not b;
    layer1_outputs(7528) <= b and not a;
    layer1_outputs(7529) <= not b or a;
    layer1_outputs(7530) <= not a;
    layer1_outputs(7531) <= not (a or b);
    layer1_outputs(7532) <= not a;
    layer1_outputs(7533) <= b and not a;
    layer1_outputs(7534) <= not b;
    layer1_outputs(7535) <= not a or b;
    layer1_outputs(7536) <= not (a or b);
    layer1_outputs(7537) <= not (a and b);
    layer1_outputs(7538) <= not a;
    layer1_outputs(7539) <= a and b;
    layer1_outputs(7540) <= a;
    layer1_outputs(7541) <= a and b;
    layer1_outputs(7542) <= not b or a;
    layer1_outputs(7543) <= not (a xor b);
    layer1_outputs(7544) <= not a or b;
    layer1_outputs(7545) <= b and not a;
    layer1_outputs(7546) <= not b or a;
    layer1_outputs(7547) <= not b;
    layer1_outputs(7548) <= not a;
    layer1_outputs(7549) <= a xor b;
    layer1_outputs(7550) <= not b;
    layer1_outputs(7551) <= b;
    layer1_outputs(7552) <= a and not b;
    layer1_outputs(7553) <= a or b;
    layer1_outputs(7554) <= b and not a;
    layer1_outputs(7555) <= a;
    layer1_outputs(7556) <= not (a or b);
    layer1_outputs(7557) <= a xor b;
    layer1_outputs(7558) <= not a;
    layer1_outputs(7559) <= not (a and b);
    layer1_outputs(7560) <= b;
    layer1_outputs(7561) <= a;
    layer1_outputs(7562) <= not a;
    layer1_outputs(7563) <= a and not b;
    layer1_outputs(7564) <= a xor b;
    layer1_outputs(7565) <= not (a and b);
    layer1_outputs(7566) <= a and b;
    layer1_outputs(7567) <= 1'b0;
    layer1_outputs(7568) <= b;
    layer1_outputs(7569) <= not (a xor b);
    layer1_outputs(7570) <= a or b;
    layer1_outputs(7571) <= a;
    layer1_outputs(7572) <= a;
    layer1_outputs(7573) <= a xor b;
    layer1_outputs(7574) <= not (a or b);
    layer1_outputs(7575) <= not b or a;
    layer1_outputs(7576) <= not a;
    layer1_outputs(7577) <= a;
    layer1_outputs(7578) <= not b or a;
    layer1_outputs(7579) <= not (a and b);
    layer1_outputs(7580) <= not a or b;
    layer1_outputs(7581) <= a xor b;
    layer1_outputs(7582) <= a xor b;
    layer1_outputs(7583) <= b and not a;
    layer1_outputs(7584) <= not a or b;
    layer1_outputs(7585) <= a and not b;
    layer1_outputs(7586) <= b and not a;
    layer1_outputs(7587) <= not b or a;
    layer1_outputs(7588) <= not b;
    layer1_outputs(7589) <= not a or b;
    layer1_outputs(7590) <= a and not b;
    layer1_outputs(7591) <= not (a or b);
    layer1_outputs(7592) <= not a;
    layer1_outputs(7593) <= b;
    layer1_outputs(7594) <= not (a xor b);
    layer1_outputs(7595) <= a;
    layer1_outputs(7596) <= a or b;
    layer1_outputs(7597) <= a or b;
    layer1_outputs(7598) <= not (a or b);
    layer1_outputs(7599) <= not b;
    layer1_outputs(7600) <= b;
    layer1_outputs(7601) <= a xor b;
    layer1_outputs(7602) <= not a or b;
    layer1_outputs(7603) <= b;
    layer1_outputs(7604) <= not a or b;
    layer1_outputs(7605) <= a xor b;
    layer1_outputs(7606) <= not a or b;
    layer1_outputs(7607) <= a or b;
    layer1_outputs(7608) <= not b;
    layer1_outputs(7609) <= not (a and b);
    layer1_outputs(7610) <= a;
    layer1_outputs(7611) <= not b or a;
    layer1_outputs(7612) <= not a;
    layer1_outputs(7613) <= not (a or b);
    layer1_outputs(7614) <= not (a or b);
    layer1_outputs(7615) <= a xor b;
    layer1_outputs(7616) <= not a or b;
    layer1_outputs(7617) <= b;
    layer1_outputs(7618) <= a;
    layer1_outputs(7619) <= not b;
    layer1_outputs(7620) <= a xor b;
    layer1_outputs(7621) <= not b or a;
    layer1_outputs(7622) <= not a or b;
    layer1_outputs(7623) <= b;
    layer1_outputs(7624) <= b and not a;
    layer1_outputs(7625) <= b and not a;
    layer1_outputs(7626) <= a and b;
    layer1_outputs(7627) <= not b;
    layer1_outputs(7628) <= a xor b;
    layer1_outputs(7629) <= not (a or b);
    layer1_outputs(7630) <= not b;
    layer1_outputs(7631) <= a and not b;
    layer1_outputs(7632) <= not (a and b);
    layer1_outputs(7633) <= b;
    layer1_outputs(7634) <= not a or b;
    layer1_outputs(7635) <= a;
    layer1_outputs(7636) <= not (a and b);
    layer1_outputs(7637) <= not (a or b);
    layer1_outputs(7638) <= a and b;
    layer1_outputs(7639) <= not (a or b);
    layer1_outputs(7640) <= not b;
    layer1_outputs(7641) <= not a or b;
    layer1_outputs(7642) <= not a;
    layer1_outputs(7643) <= a and not b;
    layer1_outputs(7644) <= b;
    layer1_outputs(7645) <= not a;
    layer1_outputs(7646) <= a;
    layer1_outputs(7647) <= not b or a;
    layer1_outputs(7648) <= not a;
    layer1_outputs(7649) <= b;
    layer1_outputs(7650) <= b and not a;
    layer1_outputs(7651) <= a xor b;
    layer1_outputs(7652) <= not (a and b);
    layer1_outputs(7653) <= a and b;
    layer1_outputs(7654) <= a;
    layer1_outputs(7655) <= a or b;
    layer1_outputs(7656) <= not a;
    layer1_outputs(7657) <= not b;
    layer1_outputs(7658) <= b and not a;
    layer1_outputs(7659) <= not b;
    layer1_outputs(7660) <= not (a xor b);
    layer1_outputs(7661) <= b;
    layer1_outputs(7662) <= not a;
    layer1_outputs(7663) <= 1'b0;
    layer1_outputs(7664) <= not a or b;
    layer1_outputs(7665) <= not a;
    layer1_outputs(7666) <= not (a or b);
    layer1_outputs(7667) <= a xor b;
    layer1_outputs(7668) <= b;
    layer1_outputs(7669) <= not b;
    layer1_outputs(7670) <= b;
    layer1_outputs(7671) <= b and not a;
    layer1_outputs(7672) <= a xor b;
    layer1_outputs(7673) <= b;
    layer1_outputs(7674) <= b and not a;
    layer1_outputs(7675) <= not a;
    layer1_outputs(7676) <= 1'b1;
    layer1_outputs(7677) <= not (a or b);
    layer1_outputs(7678) <= not a or b;
    layer1_outputs(7679) <= a;
    layer1_outputs(7680) <= a;
    layer1_outputs(7681) <= not a;
    layer1_outputs(7682) <= b;
    layer1_outputs(7683) <= not b;
    layer1_outputs(7684) <= not b;
    layer1_outputs(7685) <= b;
    layer1_outputs(7686) <= 1'b1;
    layer1_outputs(7687) <= a;
    layer1_outputs(7688) <= a xor b;
    layer1_outputs(7689) <= b and not a;
    layer1_outputs(7690) <= b;
    layer1_outputs(7691) <= not a;
    layer1_outputs(7692) <= not (a and b);
    layer1_outputs(7693) <= a xor b;
    layer1_outputs(7694) <= a and not b;
    layer1_outputs(7695) <= a xor b;
    layer1_outputs(7696) <= not b;
    layer1_outputs(7697) <= b and not a;
    layer1_outputs(7698) <= a and not b;
    layer1_outputs(7699) <= not (a xor b);
    layer1_outputs(7700) <= a xor b;
    layer1_outputs(7701) <= a or b;
    layer1_outputs(7702) <= a xor b;
    layer1_outputs(7703) <= a;
    layer1_outputs(7704) <= a;
    layer1_outputs(7705) <= not b or a;
    layer1_outputs(7706) <= a and not b;
    layer1_outputs(7707) <= not a or b;
    layer1_outputs(7708) <= not b;
    layer1_outputs(7709) <= not b;
    layer1_outputs(7710) <= b and not a;
    layer1_outputs(7711) <= a xor b;
    layer1_outputs(7712) <= not b;
    layer1_outputs(7713) <= not (a xor b);
    layer1_outputs(7714) <= not (a and b);
    layer1_outputs(7715) <= not (a xor b);
    layer1_outputs(7716) <= b;
    layer1_outputs(7717) <= not (a and b);
    layer1_outputs(7718) <= not (a or b);
    layer1_outputs(7719) <= a xor b;
    layer1_outputs(7720) <= a xor b;
    layer1_outputs(7721) <= not (a xor b);
    layer1_outputs(7722) <= a;
    layer1_outputs(7723) <= a and b;
    layer1_outputs(7724) <= not b or a;
    layer1_outputs(7725) <= b and not a;
    layer1_outputs(7726) <= a and not b;
    layer1_outputs(7727) <= a xor b;
    layer1_outputs(7728) <= not (a or b);
    layer1_outputs(7729) <= b;
    layer1_outputs(7730) <= not a or b;
    layer1_outputs(7731) <= not a;
    layer1_outputs(7732) <= not (a xor b);
    layer1_outputs(7733) <= not (a and b);
    layer1_outputs(7734) <= not a or b;
    layer1_outputs(7735) <= not a;
    layer1_outputs(7736) <= not (a or b);
    layer1_outputs(7737) <= a xor b;
    layer1_outputs(7738) <= not b;
    layer1_outputs(7739) <= not a or b;
    layer1_outputs(7740) <= not b;
    layer1_outputs(7741) <= not a or b;
    layer1_outputs(7742) <= a or b;
    layer1_outputs(7743) <= a and not b;
    layer1_outputs(7744) <= not (a or b);
    layer1_outputs(7745) <= not (a and b);
    layer1_outputs(7746) <= a and not b;
    layer1_outputs(7747) <= a and b;
    layer1_outputs(7748) <= a and not b;
    layer1_outputs(7749) <= not (a or b);
    layer1_outputs(7750) <= a;
    layer1_outputs(7751) <= not b;
    layer1_outputs(7752) <= b and not a;
    layer1_outputs(7753) <= b;
    layer1_outputs(7754) <= not (a or b);
    layer1_outputs(7755) <= not (a or b);
    layer1_outputs(7756) <= a xor b;
    layer1_outputs(7757) <= a;
    layer1_outputs(7758) <= not a;
    layer1_outputs(7759) <= not a or b;
    layer1_outputs(7760) <= not a or b;
    layer1_outputs(7761) <= a xor b;
    layer1_outputs(7762) <= a and b;
    layer1_outputs(7763) <= a and b;
    layer1_outputs(7764) <= not (a and b);
    layer1_outputs(7765) <= a and b;
    layer1_outputs(7766) <= not (a xor b);
    layer1_outputs(7767) <= not b or a;
    layer1_outputs(7768) <= a;
    layer1_outputs(7769) <= not a;
    layer1_outputs(7770) <= not (a xor b);
    layer1_outputs(7771) <= not (a xor b);
    layer1_outputs(7772) <= not (a xor b);
    layer1_outputs(7773) <= a or b;
    layer1_outputs(7774) <= not b;
    layer1_outputs(7775) <= not (a xor b);
    layer1_outputs(7776) <= a;
    layer1_outputs(7777) <= not (a xor b);
    layer1_outputs(7778) <= not (a and b);
    layer1_outputs(7779) <= b;
    layer1_outputs(7780) <= not a;
    layer1_outputs(7781) <= a or b;
    layer1_outputs(7782) <= b;
    layer1_outputs(7783) <= b;
    layer1_outputs(7784) <= not (a xor b);
    layer1_outputs(7785) <= not a or b;
    layer1_outputs(7786) <= a;
    layer1_outputs(7787) <= not (a or b);
    layer1_outputs(7788) <= 1'b1;
    layer1_outputs(7789) <= not b;
    layer1_outputs(7790) <= a and b;
    layer1_outputs(7791) <= a xor b;
    layer1_outputs(7792) <= not a;
    layer1_outputs(7793) <= a or b;
    layer1_outputs(7794) <= b;
    layer1_outputs(7795) <= a or b;
    layer1_outputs(7796) <= not (a or b);
    layer1_outputs(7797) <= not (a and b);
    layer1_outputs(7798) <= not (a xor b);
    layer1_outputs(7799) <= b and not a;
    layer1_outputs(7800) <= a xor b;
    layer1_outputs(7801) <= not b;
    layer1_outputs(7802) <= a xor b;
    layer1_outputs(7803) <= b;
    layer1_outputs(7804) <= a and b;
    layer1_outputs(7805) <= a and not b;
    layer1_outputs(7806) <= b and not a;
    layer1_outputs(7807) <= a;
    layer1_outputs(7808) <= not a;
    layer1_outputs(7809) <= 1'b0;
    layer1_outputs(7810) <= not b;
    layer1_outputs(7811) <= not (a or b);
    layer1_outputs(7812) <= a or b;
    layer1_outputs(7813) <= a and b;
    layer1_outputs(7814) <= not (a or b);
    layer1_outputs(7815) <= b and not a;
    layer1_outputs(7816) <= not b;
    layer1_outputs(7817) <= not a;
    layer1_outputs(7818) <= b;
    layer1_outputs(7819) <= not a or b;
    layer1_outputs(7820) <= a xor b;
    layer1_outputs(7821) <= not b or a;
    layer1_outputs(7822) <= not (a xor b);
    layer1_outputs(7823) <= b;
    layer1_outputs(7824) <= b and not a;
    layer1_outputs(7825) <= a and b;
    layer1_outputs(7826) <= b;
    layer1_outputs(7827) <= not b;
    layer1_outputs(7828) <= not (a and b);
    layer1_outputs(7829) <= a or b;
    layer1_outputs(7830) <= not a;
    layer1_outputs(7831) <= not (a or b);
    layer1_outputs(7832) <= a xor b;
    layer1_outputs(7833) <= not a;
    layer1_outputs(7834) <= not (a and b);
    layer1_outputs(7835) <= a or b;
    layer1_outputs(7836) <= b and not a;
    layer1_outputs(7837) <= not b;
    layer1_outputs(7838) <= b and not a;
    layer1_outputs(7839) <= a or b;
    layer1_outputs(7840) <= a;
    layer1_outputs(7841) <= a and not b;
    layer1_outputs(7842) <= b and not a;
    layer1_outputs(7843) <= not a or b;
    layer1_outputs(7844) <= a;
    layer1_outputs(7845) <= not (a xor b);
    layer1_outputs(7846) <= b;
    layer1_outputs(7847) <= not a or b;
    layer1_outputs(7848) <= a and b;
    layer1_outputs(7849) <= not b;
    layer1_outputs(7850) <= a and not b;
    layer1_outputs(7851) <= not b;
    layer1_outputs(7852) <= not a;
    layer1_outputs(7853) <= a and b;
    layer1_outputs(7854) <= a xor b;
    layer1_outputs(7855) <= not (a and b);
    layer1_outputs(7856) <= not a;
    layer1_outputs(7857) <= a and not b;
    layer1_outputs(7858) <= a and not b;
    layer1_outputs(7859) <= b and not a;
    layer1_outputs(7860) <= a and not b;
    layer1_outputs(7861) <= a xor b;
    layer1_outputs(7862) <= not (a and b);
    layer1_outputs(7863) <= not a or b;
    layer1_outputs(7864) <= a or b;
    layer1_outputs(7865) <= not (a or b);
    layer1_outputs(7866) <= not a or b;
    layer1_outputs(7867) <= a and not b;
    layer1_outputs(7868) <= not (a xor b);
    layer1_outputs(7869) <= a and b;
    layer1_outputs(7870) <= not (a xor b);
    layer1_outputs(7871) <= a;
    layer1_outputs(7872) <= a and not b;
    layer1_outputs(7873) <= a and b;
    layer1_outputs(7874) <= not (a or b);
    layer1_outputs(7875) <= not a;
    layer1_outputs(7876) <= a and not b;
    layer1_outputs(7877) <= not a or b;
    layer1_outputs(7878) <= a;
    layer1_outputs(7879) <= a or b;
    layer1_outputs(7880) <= b;
    layer1_outputs(7881) <= a;
    layer1_outputs(7882) <= a xor b;
    layer1_outputs(7883) <= a;
    layer1_outputs(7884) <= a and not b;
    layer1_outputs(7885) <= a xor b;
    layer1_outputs(7886) <= a xor b;
    layer1_outputs(7887) <= not a;
    layer1_outputs(7888) <= b;
    layer1_outputs(7889) <= a;
    layer1_outputs(7890) <= a xor b;
    layer1_outputs(7891) <= not a or b;
    layer1_outputs(7892) <= not b or a;
    layer1_outputs(7893) <= not (a xor b);
    layer1_outputs(7894) <= a and not b;
    layer1_outputs(7895) <= not b or a;
    layer1_outputs(7896) <= not b or a;
    layer1_outputs(7897) <= a and b;
    layer1_outputs(7898) <= b and not a;
    layer1_outputs(7899) <= not (a xor b);
    layer1_outputs(7900) <= b and not a;
    layer1_outputs(7901) <= not (a xor b);
    layer1_outputs(7902) <= a or b;
    layer1_outputs(7903) <= not (a xor b);
    layer1_outputs(7904) <= a;
    layer1_outputs(7905) <= not a or b;
    layer1_outputs(7906) <= not (a and b);
    layer1_outputs(7907) <= a and not b;
    layer1_outputs(7908) <= not b or a;
    layer1_outputs(7909) <= not a or b;
    layer1_outputs(7910) <= b;
    layer1_outputs(7911) <= a xor b;
    layer1_outputs(7912) <= not (a xor b);
    layer1_outputs(7913) <= not (a or b);
    layer1_outputs(7914) <= not (a xor b);
    layer1_outputs(7915) <= not a or b;
    layer1_outputs(7916) <= a;
    layer1_outputs(7917) <= not (a and b);
    layer1_outputs(7918) <= not (a or b);
    layer1_outputs(7919) <= a;
    layer1_outputs(7920) <= not (a xor b);
    layer1_outputs(7921) <= a;
    layer1_outputs(7922) <= not b or a;
    layer1_outputs(7923) <= not (a xor b);
    layer1_outputs(7924) <= a or b;
    layer1_outputs(7925) <= not a;
    layer1_outputs(7926) <= not (a or b);
    layer1_outputs(7927) <= not b;
    layer1_outputs(7928) <= not (a xor b);
    layer1_outputs(7929) <= 1'b0;
    layer1_outputs(7930) <= a xor b;
    layer1_outputs(7931) <= not a;
    layer1_outputs(7932) <= b and not a;
    layer1_outputs(7933) <= not (a xor b);
    layer1_outputs(7934) <= a;
    layer1_outputs(7935) <= not b;
    layer1_outputs(7936) <= not b;
    layer1_outputs(7937) <= not a or b;
    layer1_outputs(7938) <= not (a xor b);
    layer1_outputs(7939) <= not (a and b);
    layer1_outputs(7940) <= not (a xor b);
    layer1_outputs(7941) <= not b;
    layer1_outputs(7942) <= not (a xor b);
    layer1_outputs(7943) <= a;
    layer1_outputs(7944) <= not b;
    layer1_outputs(7945) <= a or b;
    layer1_outputs(7946) <= b;
    layer1_outputs(7947) <= b;
    layer1_outputs(7948) <= a;
    layer1_outputs(7949) <= a xor b;
    layer1_outputs(7950) <= not (a or b);
    layer1_outputs(7951) <= not a;
    layer1_outputs(7952) <= not a or b;
    layer1_outputs(7953) <= a or b;
    layer1_outputs(7954) <= not b or a;
    layer1_outputs(7955) <= not b;
    layer1_outputs(7956) <= not a or b;
    layer1_outputs(7957) <= a and b;
    layer1_outputs(7958) <= a or b;
    layer1_outputs(7959) <= b;
    layer1_outputs(7960) <= a xor b;
    layer1_outputs(7961) <= a;
    layer1_outputs(7962) <= not b or a;
    layer1_outputs(7963) <= a;
    layer1_outputs(7964) <= not a;
    layer1_outputs(7965) <= a and b;
    layer1_outputs(7966) <= not a or b;
    layer1_outputs(7967) <= not b;
    layer1_outputs(7968) <= not b or a;
    layer1_outputs(7969) <= not (a xor b);
    layer1_outputs(7970) <= not (a and b);
    layer1_outputs(7971) <= b and not a;
    layer1_outputs(7972) <= not a;
    layer1_outputs(7973) <= a;
    layer1_outputs(7974) <= not b;
    layer1_outputs(7975) <= a and not b;
    layer1_outputs(7976) <= not (a and b);
    layer1_outputs(7977) <= not b;
    layer1_outputs(7978) <= a;
    layer1_outputs(7979) <= a;
    layer1_outputs(7980) <= a;
    layer1_outputs(7981) <= not b or a;
    layer1_outputs(7982) <= a;
    layer1_outputs(7983) <= 1'b0;
    layer1_outputs(7984) <= not a or b;
    layer1_outputs(7985) <= not b;
    layer1_outputs(7986) <= not (a or b);
    layer1_outputs(7987) <= b and not a;
    layer1_outputs(7988) <= not (a xor b);
    layer1_outputs(7989) <= a;
    layer1_outputs(7990) <= a and b;
    layer1_outputs(7991) <= b;
    layer1_outputs(7992) <= b;
    layer1_outputs(7993) <= not b;
    layer1_outputs(7994) <= a xor b;
    layer1_outputs(7995) <= not a;
    layer1_outputs(7996) <= b;
    layer1_outputs(7997) <= not a;
    layer1_outputs(7998) <= not b or a;
    layer1_outputs(7999) <= a and b;
    layer1_outputs(8000) <= not a;
    layer1_outputs(8001) <= not (a xor b);
    layer1_outputs(8002) <= not b or a;
    layer1_outputs(8003) <= not (a xor b);
    layer1_outputs(8004) <= a and not b;
    layer1_outputs(8005) <= not b;
    layer1_outputs(8006) <= not a or b;
    layer1_outputs(8007) <= a and b;
    layer1_outputs(8008) <= a or b;
    layer1_outputs(8009) <= not a or b;
    layer1_outputs(8010) <= not a;
    layer1_outputs(8011) <= 1'b1;
    layer1_outputs(8012) <= not (a xor b);
    layer1_outputs(8013) <= not b;
    layer1_outputs(8014) <= a;
    layer1_outputs(8015) <= not b;
    layer1_outputs(8016) <= not a or b;
    layer1_outputs(8017) <= a;
    layer1_outputs(8018) <= not b or a;
    layer1_outputs(8019) <= not a;
    layer1_outputs(8020) <= b and not a;
    layer1_outputs(8021) <= not b or a;
    layer1_outputs(8022) <= b;
    layer1_outputs(8023) <= b;
    layer1_outputs(8024) <= not (a or b);
    layer1_outputs(8025) <= a and not b;
    layer1_outputs(8026) <= b;
    layer1_outputs(8027) <= a xor b;
    layer1_outputs(8028) <= not a;
    layer1_outputs(8029) <= not b;
    layer1_outputs(8030) <= a and not b;
    layer1_outputs(8031) <= 1'b0;
    layer1_outputs(8032) <= a xor b;
    layer1_outputs(8033) <= not b or a;
    layer1_outputs(8034) <= 1'b0;
    layer1_outputs(8035) <= b and not a;
    layer1_outputs(8036) <= b;
    layer1_outputs(8037) <= not a;
    layer1_outputs(8038) <= a;
    layer1_outputs(8039) <= not a or b;
    layer1_outputs(8040) <= a and b;
    layer1_outputs(8041) <= a and not b;
    layer1_outputs(8042) <= a and b;
    layer1_outputs(8043) <= not b;
    layer1_outputs(8044) <= a xor b;
    layer1_outputs(8045) <= b and not a;
    layer1_outputs(8046) <= not a;
    layer1_outputs(8047) <= 1'b1;
    layer1_outputs(8048) <= a or b;
    layer1_outputs(8049) <= not a or b;
    layer1_outputs(8050) <= not a or b;
    layer1_outputs(8051) <= a xor b;
    layer1_outputs(8052) <= a xor b;
    layer1_outputs(8053) <= a xor b;
    layer1_outputs(8054) <= a xor b;
    layer1_outputs(8055) <= not a;
    layer1_outputs(8056) <= not (a and b);
    layer1_outputs(8057) <= a xor b;
    layer1_outputs(8058) <= not b;
    layer1_outputs(8059) <= b;
    layer1_outputs(8060) <= a and not b;
    layer1_outputs(8061) <= not a;
    layer1_outputs(8062) <= b;
    layer1_outputs(8063) <= a and b;
    layer1_outputs(8064) <= not (a xor b);
    layer1_outputs(8065) <= a;
    layer1_outputs(8066) <= a;
    layer1_outputs(8067) <= b and not a;
    layer1_outputs(8068) <= a or b;
    layer1_outputs(8069) <= 1'b0;
    layer1_outputs(8070) <= a;
    layer1_outputs(8071) <= b;
    layer1_outputs(8072) <= not (a xor b);
    layer1_outputs(8073) <= a xor b;
    layer1_outputs(8074) <= a;
    layer1_outputs(8075) <= not b;
    layer1_outputs(8076) <= a;
    layer1_outputs(8077) <= a xor b;
    layer1_outputs(8078) <= not b or a;
    layer1_outputs(8079) <= a xor b;
    layer1_outputs(8080) <= not b or a;
    layer1_outputs(8081) <= not b or a;
    layer1_outputs(8082) <= not b or a;
    layer1_outputs(8083) <= a;
    layer1_outputs(8084) <= a;
    layer1_outputs(8085) <= not b;
    layer1_outputs(8086) <= not a;
    layer1_outputs(8087) <= a and b;
    layer1_outputs(8088) <= not (a and b);
    layer1_outputs(8089) <= b;
    layer1_outputs(8090) <= a;
    layer1_outputs(8091) <= a or b;
    layer1_outputs(8092) <= not a;
    layer1_outputs(8093) <= a and not b;
    layer1_outputs(8094) <= a or b;
    layer1_outputs(8095) <= not b or a;
    layer1_outputs(8096) <= not a or b;
    layer1_outputs(8097) <= not a;
    layer1_outputs(8098) <= not (a or b);
    layer1_outputs(8099) <= not b or a;
    layer1_outputs(8100) <= not a or b;
    layer1_outputs(8101) <= b and not a;
    layer1_outputs(8102) <= not (a xor b);
    layer1_outputs(8103) <= not (a and b);
    layer1_outputs(8104) <= not (a or b);
    layer1_outputs(8105) <= a;
    layer1_outputs(8106) <= not a;
    layer1_outputs(8107) <= not b or a;
    layer1_outputs(8108) <= not a or b;
    layer1_outputs(8109) <= a or b;
    layer1_outputs(8110) <= not b;
    layer1_outputs(8111) <= not b;
    layer1_outputs(8112) <= a and b;
    layer1_outputs(8113) <= not a;
    layer1_outputs(8114) <= not b or a;
    layer1_outputs(8115) <= b;
    layer1_outputs(8116) <= not a;
    layer1_outputs(8117) <= not a;
    layer1_outputs(8118) <= not b;
    layer1_outputs(8119) <= a xor b;
    layer1_outputs(8120) <= a xor b;
    layer1_outputs(8121) <= a;
    layer1_outputs(8122) <= a or b;
    layer1_outputs(8123) <= a or b;
    layer1_outputs(8124) <= a and not b;
    layer1_outputs(8125) <= b;
    layer1_outputs(8126) <= not b or a;
    layer1_outputs(8127) <= a or b;
    layer1_outputs(8128) <= not (a or b);
    layer1_outputs(8129) <= not a;
    layer1_outputs(8130) <= not a;
    layer1_outputs(8131) <= a xor b;
    layer1_outputs(8132) <= b;
    layer1_outputs(8133) <= a xor b;
    layer1_outputs(8134) <= not (a or b);
    layer1_outputs(8135) <= b;
    layer1_outputs(8136) <= not a or b;
    layer1_outputs(8137) <= a xor b;
    layer1_outputs(8138) <= b;
    layer1_outputs(8139) <= a xor b;
    layer1_outputs(8140) <= not a or b;
    layer1_outputs(8141) <= a or b;
    layer1_outputs(8142) <= a and b;
    layer1_outputs(8143) <= a;
    layer1_outputs(8144) <= not b or a;
    layer1_outputs(8145) <= b;
    layer1_outputs(8146) <= not b or a;
    layer1_outputs(8147) <= a;
    layer1_outputs(8148) <= not b or a;
    layer1_outputs(8149) <= not (a and b);
    layer1_outputs(8150) <= not (a xor b);
    layer1_outputs(8151) <= a;
    layer1_outputs(8152) <= a xor b;
    layer1_outputs(8153) <= a;
    layer1_outputs(8154) <= b;
    layer1_outputs(8155) <= not a;
    layer1_outputs(8156) <= b and not a;
    layer1_outputs(8157) <= not b;
    layer1_outputs(8158) <= b and not a;
    layer1_outputs(8159) <= not a or b;
    layer1_outputs(8160) <= not (a or b);
    layer1_outputs(8161) <= not (a xor b);
    layer1_outputs(8162) <= 1'b1;
    layer1_outputs(8163) <= b;
    layer1_outputs(8164) <= a;
    layer1_outputs(8165) <= not (a and b);
    layer1_outputs(8166) <= not b or a;
    layer1_outputs(8167) <= not a;
    layer1_outputs(8168) <= not b;
    layer1_outputs(8169) <= not a;
    layer1_outputs(8170) <= not (a or b);
    layer1_outputs(8171) <= b;
    layer1_outputs(8172) <= not b;
    layer1_outputs(8173) <= not a;
    layer1_outputs(8174) <= not b;
    layer1_outputs(8175) <= not a;
    layer1_outputs(8176) <= a xor b;
    layer1_outputs(8177) <= b;
    layer1_outputs(8178) <= b;
    layer1_outputs(8179) <= b;
    layer1_outputs(8180) <= b;
    layer1_outputs(8181) <= b;
    layer1_outputs(8182) <= not (a or b);
    layer1_outputs(8183) <= not a;
    layer1_outputs(8184) <= a and b;
    layer1_outputs(8185) <= b and not a;
    layer1_outputs(8186) <= not a or b;
    layer1_outputs(8187) <= not b;
    layer1_outputs(8188) <= not b or a;
    layer1_outputs(8189) <= not (a xor b);
    layer1_outputs(8190) <= b;
    layer1_outputs(8191) <= 1'b0;
    layer1_outputs(8192) <= not (a and b);
    layer1_outputs(8193) <= not a or b;
    layer1_outputs(8194) <= a and not b;
    layer1_outputs(8195) <= a and not b;
    layer1_outputs(8196) <= not b;
    layer1_outputs(8197) <= not (a xor b);
    layer1_outputs(8198) <= not a or b;
    layer1_outputs(8199) <= b;
    layer1_outputs(8200) <= b;
    layer1_outputs(8201) <= a;
    layer1_outputs(8202) <= a;
    layer1_outputs(8203) <= a and not b;
    layer1_outputs(8204) <= a and not b;
    layer1_outputs(8205) <= a;
    layer1_outputs(8206) <= a xor b;
    layer1_outputs(8207) <= not a or b;
    layer1_outputs(8208) <= 1'b0;
    layer1_outputs(8209) <= a or b;
    layer1_outputs(8210) <= not b;
    layer1_outputs(8211) <= a and not b;
    layer1_outputs(8212) <= not (a or b);
    layer1_outputs(8213) <= not (a or b);
    layer1_outputs(8214) <= b;
    layer1_outputs(8215) <= not b;
    layer1_outputs(8216) <= a and not b;
    layer1_outputs(8217) <= not (a or b);
    layer1_outputs(8218) <= 1'b0;
    layer1_outputs(8219) <= not (a or b);
    layer1_outputs(8220) <= not (a and b);
    layer1_outputs(8221) <= a and b;
    layer1_outputs(8222) <= not (a and b);
    layer1_outputs(8223) <= b and not a;
    layer1_outputs(8224) <= not (a or b);
    layer1_outputs(8225) <= a or b;
    layer1_outputs(8226) <= not b or a;
    layer1_outputs(8227) <= a xor b;
    layer1_outputs(8228) <= a xor b;
    layer1_outputs(8229) <= not (a xor b);
    layer1_outputs(8230) <= not b;
    layer1_outputs(8231) <= not b;
    layer1_outputs(8232) <= a xor b;
    layer1_outputs(8233) <= a and not b;
    layer1_outputs(8234) <= not b;
    layer1_outputs(8235) <= a and b;
    layer1_outputs(8236) <= not b or a;
    layer1_outputs(8237) <= a and b;
    layer1_outputs(8238) <= not b;
    layer1_outputs(8239) <= not (a and b);
    layer1_outputs(8240) <= not (a xor b);
    layer1_outputs(8241) <= not a;
    layer1_outputs(8242) <= a and not b;
    layer1_outputs(8243) <= a xor b;
    layer1_outputs(8244) <= a;
    layer1_outputs(8245) <= not (a xor b);
    layer1_outputs(8246) <= not b;
    layer1_outputs(8247) <= a and b;
    layer1_outputs(8248) <= not (a xor b);
    layer1_outputs(8249) <= not b;
    layer1_outputs(8250) <= a and b;
    layer1_outputs(8251) <= not (a or b);
    layer1_outputs(8252) <= b and not a;
    layer1_outputs(8253) <= not (a xor b);
    layer1_outputs(8254) <= b;
    layer1_outputs(8255) <= a or b;
    layer1_outputs(8256) <= a xor b;
    layer1_outputs(8257) <= a xor b;
    layer1_outputs(8258) <= b and not a;
    layer1_outputs(8259) <= a;
    layer1_outputs(8260) <= b;
    layer1_outputs(8261) <= not a or b;
    layer1_outputs(8262) <= a xor b;
    layer1_outputs(8263) <= a or b;
    layer1_outputs(8264) <= not (a or b);
    layer1_outputs(8265) <= a or b;
    layer1_outputs(8266) <= a xor b;
    layer1_outputs(8267) <= a and b;
    layer1_outputs(8268) <= not a or b;
    layer1_outputs(8269) <= not a;
    layer1_outputs(8270) <= a;
    layer1_outputs(8271) <= b;
    layer1_outputs(8272) <= a;
    layer1_outputs(8273) <= a xor b;
    layer1_outputs(8274) <= a and b;
    layer1_outputs(8275) <= not a;
    layer1_outputs(8276) <= a and not b;
    layer1_outputs(8277) <= a;
    layer1_outputs(8278) <= a and not b;
    layer1_outputs(8279) <= b and not a;
    layer1_outputs(8280) <= a and b;
    layer1_outputs(8281) <= b;
    layer1_outputs(8282) <= not a or b;
    layer1_outputs(8283) <= b and not a;
    layer1_outputs(8284) <= b and not a;
    layer1_outputs(8285) <= not a;
    layer1_outputs(8286) <= a xor b;
    layer1_outputs(8287) <= a and not b;
    layer1_outputs(8288) <= a or b;
    layer1_outputs(8289) <= not b;
    layer1_outputs(8290) <= a and not b;
    layer1_outputs(8291) <= b;
    layer1_outputs(8292) <= b;
    layer1_outputs(8293) <= b;
    layer1_outputs(8294) <= not a;
    layer1_outputs(8295) <= not (a or b);
    layer1_outputs(8296) <= not b or a;
    layer1_outputs(8297) <= a or b;
    layer1_outputs(8298) <= a and b;
    layer1_outputs(8299) <= a and b;
    layer1_outputs(8300) <= a and b;
    layer1_outputs(8301) <= not a or b;
    layer1_outputs(8302) <= a xor b;
    layer1_outputs(8303) <= not (a and b);
    layer1_outputs(8304) <= not b;
    layer1_outputs(8305) <= not (a or b);
    layer1_outputs(8306) <= not b or a;
    layer1_outputs(8307) <= b and not a;
    layer1_outputs(8308) <= b and not a;
    layer1_outputs(8309) <= a xor b;
    layer1_outputs(8310) <= b;
    layer1_outputs(8311) <= not (a and b);
    layer1_outputs(8312) <= b;
    layer1_outputs(8313) <= not a or b;
    layer1_outputs(8314) <= a xor b;
    layer1_outputs(8315) <= b and not a;
    layer1_outputs(8316) <= not a;
    layer1_outputs(8317) <= not a or b;
    layer1_outputs(8318) <= a xor b;
    layer1_outputs(8319) <= not b;
    layer1_outputs(8320) <= a xor b;
    layer1_outputs(8321) <= a and not b;
    layer1_outputs(8322) <= not (a or b);
    layer1_outputs(8323) <= a or b;
    layer1_outputs(8324) <= 1'b1;
    layer1_outputs(8325) <= not b or a;
    layer1_outputs(8326) <= a xor b;
    layer1_outputs(8327) <= not b;
    layer1_outputs(8328) <= not (a xor b);
    layer1_outputs(8329) <= b and not a;
    layer1_outputs(8330) <= b;
    layer1_outputs(8331) <= b;
    layer1_outputs(8332) <= a or b;
    layer1_outputs(8333) <= not (a and b);
    layer1_outputs(8334) <= a or b;
    layer1_outputs(8335) <= not a;
    layer1_outputs(8336) <= a or b;
    layer1_outputs(8337) <= b and not a;
    layer1_outputs(8338) <= a;
    layer1_outputs(8339) <= not b;
    layer1_outputs(8340) <= not (a and b);
    layer1_outputs(8341) <= a and not b;
    layer1_outputs(8342) <= a;
    layer1_outputs(8343) <= not (a xor b);
    layer1_outputs(8344) <= not a or b;
    layer1_outputs(8345) <= b;
    layer1_outputs(8346) <= a or b;
    layer1_outputs(8347) <= a and b;
    layer1_outputs(8348) <= not (a or b);
    layer1_outputs(8349) <= a;
    layer1_outputs(8350) <= not a or b;
    layer1_outputs(8351) <= a and not b;
    layer1_outputs(8352) <= 1'b1;
    layer1_outputs(8353) <= a and b;
    layer1_outputs(8354) <= not a or b;
    layer1_outputs(8355) <= a and b;
    layer1_outputs(8356) <= a xor b;
    layer1_outputs(8357) <= a;
    layer1_outputs(8358) <= a xor b;
    layer1_outputs(8359) <= not a or b;
    layer1_outputs(8360) <= b;
    layer1_outputs(8361) <= not a;
    layer1_outputs(8362) <= not a;
    layer1_outputs(8363) <= b and not a;
    layer1_outputs(8364) <= a and not b;
    layer1_outputs(8365) <= not (a xor b);
    layer1_outputs(8366) <= not (a xor b);
    layer1_outputs(8367) <= not (a xor b);
    layer1_outputs(8368) <= a or b;
    layer1_outputs(8369) <= not b;
    layer1_outputs(8370) <= not b or a;
    layer1_outputs(8371) <= not (a or b);
    layer1_outputs(8372) <= b and not a;
    layer1_outputs(8373) <= not b;
    layer1_outputs(8374) <= a xor b;
    layer1_outputs(8375) <= 1'b0;
    layer1_outputs(8376) <= not (a and b);
    layer1_outputs(8377) <= a or b;
    layer1_outputs(8378) <= not (a xor b);
    layer1_outputs(8379) <= not (a and b);
    layer1_outputs(8380) <= b and not a;
    layer1_outputs(8381) <= not b or a;
    layer1_outputs(8382) <= not (a xor b);
    layer1_outputs(8383) <= a and b;
    layer1_outputs(8384) <= not (a and b);
    layer1_outputs(8385) <= a xor b;
    layer1_outputs(8386) <= not b;
    layer1_outputs(8387) <= not b;
    layer1_outputs(8388) <= not (a or b);
    layer1_outputs(8389) <= a and not b;
    layer1_outputs(8390) <= b;
    layer1_outputs(8391) <= 1'b1;
    layer1_outputs(8392) <= a or b;
    layer1_outputs(8393) <= a or b;
    layer1_outputs(8394) <= a xor b;
    layer1_outputs(8395) <= b and not a;
    layer1_outputs(8396) <= not b;
    layer1_outputs(8397) <= not a;
    layer1_outputs(8398) <= not (a and b);
    layer1_outputs(8399) <= a and not b;
    layer1_outputs(8400) <= a or b;
    layer1_outputs(8401) <= not b;
    layer1_outputs(8402) <= a and b;
    layer1_outputs(8403) <= a;
    layer1_outputs(8404) <= not (a and b);
    layer1_outputs(8405) <= a;
    layer1_outputs(8406) <= not (a xor b);
    layer1_outputs(8407) <= a;
    layer1_outputs(8408) <= not a or b;
    layer1_outputs(8409) <= not (a and b);
    layer1_outputs(8410) <= not a;
    layer1_outputs(8411) <= a xor b;
    layer1_outputs(8412) <= not (a xor b);
    layer1_outputs(8413) <= a xor b;
    layer1_outputs(8414) <= a;
    layer1_outputs(8415) <= not (a xor b);
    layer1_outputs(8416) <= not a or b;
    layer1_outputs(8417) <= 1'b1;
    layer1_outputs(8418) <= a and b;
    layer1_outputs(8419) <= 1'b1;
    layer1_outputs(8420) <= b;
    layer1_outputs(8421) <= not b or a;
    layer1_outputs(8422) <= not b or a;
    layer1_outputs(8423) <= a;
    layer1_outputs(8424) <= b;
    layer1_outputs(8425) <= a;
    layer1_outputs(8426) <= b;
    layer1_outputs(8427) <= not b;
    layer1_outputs(8428) <= not (a and b);
    layer1_outputs(8429) <= not (a or b);
    layer1_outputs(8430) <= not (a xor b);
    layer1_outputs(8431) <= not b or a;
    layer1_outputs(8432) <= not (a and b);
    layer1_outputs(8433) <= not b;
    layer1_outputs(8434) <= not (a and b);
    layer1_outputs(8435) <= a or b;
    layer1_outputs(8436) <= not b or a;
    layer1_outputs(8437) <= b;
    layer1_outputs(8438) <= not (a or b);
    layer1_outputs(8439) <= b and not a;
    layer1_outputs(8440) <= a;
    layer1_outputs(8441) <= b;
    layer1_outputs(8442) <= a and b;
    layer1_outputs(8443) <= a xor b;
    layer1_outputs(8444) <= not b;
    layer1_outputs(8445) <= b and not a;
    layer1_outputs(8446) <= not a or b;
    layer1_outputs(8447) <= not b or a;
    layer1_outputs(8448) <= not (a and b);
    layer1_outputs(8449) <= a or b;
    layer1_outputs(8450) <= b;
    layer1_outputs(8451) <= not b or a;
    layer1_outputs(8452) <= a or b;
    layer1_outputs(8453) <= not b;
    layer1_outputs(8454) <= a xor b;
    layer1_outputs(8455) <= b and not a;
    layer1_outputs(8456) <= not b;
    layer1_outputs(8457) <= b and not a;
    layer1_outputs(8458) <= not (a or b);
    layer1_outputs(8459) <= a;
    layer1_outputs(8460) <= not a;
    layer1_outputs(8461) <= not a;
    layer1_outputs(8462) <= not (a xor b);
    layer1_outputs(8463) <= a xor b;
    layer1_outputs(8464) <= not (a xor b);
    layer1_outputs(8465) <= not (a and b);
    layer1_outputs(8466) <= b;
    layer1_outputs(8467) <= not a;
    layer1_outputs(8468) <= not a;
    layer1_outputs(8469) <= a;
    layer1_outputs(8470) <= a;
    layer1_outputs(8471) <= a;
    layer1_outputs(8472) <= not b or a;
    layer1_outputs(8473) <= a or b;
    layer1_outputs(8474) <= not (a xor b);
    layer1_outputs(8475) <= a and not b;
    layer1_outputs(8476) <= not a or b;
    layer1_outputs(8477) <= b;
    layer1_outputs(8478) <= a;
    layer1_outputs(8479) <= a xor b;
    layer1_outputs(8480) <= a and not b;
    layer1_outputs(8481) <= not a;
    layer1_outputs(8482) <= a;
    layer1_outputs(8483) <= b;
    layer1_outputs(8484) <= not (a and b);
    layer1_outputs(8485) <= not (a or b);
    layer1_outputs(8486) <= not b or a;
    layer1_outputs(8487) <= a and b;
    layer1_outputs(8488) <= a;
    layer1_outputs(8489) <= not b or a;
    layer1_outputs(8490) <= not (a and b);
    layer1_outputs(8491) <= a and not b;
    layer1_outputs(8492) <= not a;
    layer1_outputs(8493) <= b and not a;
    layer1_outputs(8494) <= not (a or b);
    layer1_outputs(8495) <= not b or a;
    layer1_outputs(8496) <= not (a xor b);
    layer1_outputs(8497) <= a;
    layer1_outputs(8498) <= not (a xor b);
    layer1_outputs(8499) <= not b or a;
    layer1_outputs(8500) <= a xor b;
    layer1_outputs(8501) <= a or b;
    layer1_outputs(8502) <= a or b;
    layer1_outputs(8503) <= not b;
    layer1_outputs(8504) <= not b or a;
    layer1_outputs(8505) <= a;
    layer1_outputs(8506) <= not (a xor b);
    layer1_outputs(8507) <= not b;
    layer1_outputs(8508) <= not (a xor b);
    layer1_outputs(8509) <= not a;
    layer1_outputs(8510) <= not (a xor b);
    layer1_outputs(8511) <= not (a or b);
    layer1_outputs(8512) <= not (a or b);
    layer1_outputs(8513) <= a;
    layer1_outputs(8514) <= a xor b;
    layer1_outputs(8515) <= not b or a;
    layer1_outputs(8516) <= not a;
    layer1_outputs(8517) <= not a;
    layer1_outputs(8518) <= not (a or b);
    layer1_outputs(8519) <= a;
    layer1_outputs(8520) <= not b;
    layer1_outputs(8521) <= not b or a;
    layer1_outputs(8522) <= not b or a;
    layer1_outputs(8523) <= a xor b;
    layer1_outputs(8524) <= a xor b;
    layer1_outputs(8525) <= not b or a;
    layer1_outputs(8526) <= not a or b;
    layer1_outputs(8527) <= not a;
    layer1_outputs(8528) <= not a;
    layer1_outputs(8529) <= not b or a;
    layer1_outputs(8530) <= b;
    layer1_outputs(8531) <= a xor b;
    layer1_outputs(8532) <= a;
    layer1_outputs(8533) <= not b;
    layer1_outputs(8534) <= not (a and b);
    layer1_outputs(8535) <= a and not b;
    layer1_outputs(8536) <= not a;
    layer1_outputs(8537) <= a xor b;
    layer1_outputs(8538) <= not b or a;
    layer1_outputs(8539) <= not a;
    layer1_outputs(8540) <= a;
    layer1_outputs(8541) <= b;
    layer1_outputs(8542) <= not b or a;
    layer1_outputs(8543) <= a;
    layer1_outputs(8544) <= not a;
    layer1_outputs(8545) <= not a;
    layer1_outputs(8546) <= a;
    layer1_outputs(8547) <= a and not b;
    layer1_outputs(8548) <= a xor b;
    layer1_outputs(8549) <= not b;
    layer1_outputs(8550) <= a and b;
    layer1_outputs(8551) <= a or b;
    layer1_outputs(8552) <= a xor b;
    layer1_outputs(8553) <= not (a xor b);
    layer1_outputs(8554) <= a and not b;
    layer1_outputs(8555) <= a;
    layer1_outputs(8556) <= a and b;
    layer1_outputs(8557) <= 1'b1;
    layer1_outputs(8558) <= not (a or b);
    layer1_outputs(8559) <= not b;
    layer1_outputs(8560) <= not (a xor b);
    layer1_outputs(8561) <= b;
    layer1_outputs(8562) <= a;
    layer1_outputs(8563) <= not (a and b);
    layer1_outputs(8564) <= not (a xor b);
    layer1_outputs(8565) <= not b or a;
    layer1_outputs(8566) <= not b or a;
    layer1_outputs(8567) <= not (a xor b);
    layer1_outputs(8568) <= a xor b;
    layer1_outputs(8569) <= not (a xor b);
    layer1_outputs(8570) <= not a or b;
    layer1_outputs(8571) <= a and b;
    layer1_outputs(8572) <= a or b;
    layer1_outputs(8573) <= a xor b;
    layer1_outputs(8574) <= not b;
    layer1_outputs(8575) <= a and not b;
    layer1_outputs(8576) <= b and not a;
    layer1_outputs(8577) <= not a or b;
    layer1_outputs(8578) <= not (a and b);
    layer1_outputs(8579) <= a xor b;
    layer1_outputs(8580) <= not b or a;
    layer1_outputs(8581) <= b;
    layer1_outputs(8582) <= a and b;
    layer1_outputs(8583) <= not a;
    layer1_outputs(8584) <= a xor b;
    layer1_outputs(8585) <= a and b;
    layer1_outputs(8586) <= not a;
    layer1_outputs(8587) <= a xor b;
    layer1_outputs(8588) <= not (a xor b);
    layer1_outputs(8589) <= not b or a;
    layer1_outputs(8590) <= not b;
    layer1_outputs(8591) <= a and b;
    layer1_outputs(8592) <= not b or a;
    layer1_outputs(8593) <= a or b;
    layer1_outputs(8594) <= a and b;
    layer1_outputs(8595) <= not b;
    layer1_outputs(8596) <= not a or b;
    layer1_outputs(8597) <= a and not b;
    layer1_outputs(8598) <= not a or b;
    layer1_outputs(8599) <= a or b;
    layer1_outputs(8600) <= not a or b;
    layer1_outputs(8601) <= not a;
    layer1_outputs(8602) <= not (a xor b);
    layer1_outputs(8603) <= a and not b;
    layer1_outputs(8604) <= not (a and b);
    layer1_outputs(8605) <= not (a xor b);
    layer1_outputs(8606) <= a xor b;
    layer1_outputs(8607) <= a or b;
    layer1_outputs(8608) <= 1'b1;
    layer1_outputs(8609) <= not b or a;
    layer1_outputs(8610) <= not b or a;
    layer1_outputs(8611) <= b and not a;
    layer1_outputs(8612) <= not a;
    layer1_outputs(8613) <= a or b;
    layer1_outputs(8614) <= a;
    layer1_outputs(8615) <= not b or a;
    layer1_outputs(8616) <= a xor b;
    layer1_outputs(8617) <= a xor b;
    layer1_outputs(8618) <= not (a and b);
    layer1_outputs(8619) <= b;
    layer1_outputs(8620) <= not a;
    layer1_outputs(8621) <= a xor b;
    layer1_outputs(8622) <= a and not b;
    layer1_outputs(8623) <= not b;
    layer1_outputs(8624) <= not a or b;
    layer1_outputs(8625) <= not (a or b);
    layer1_outputs(8626) <= not a;
    layer1_outputs(8627) <= not b;
    layer1_outputs(8628) <= not a;
    layer1_outputs(8629) <= not a;
    layer1_outputs(8630) <= 1'b1;
    layer1_outputs(8631) <= a;
    layer1_outputs(8632) <= not b;
    layer1_outputs(8633) <= a or b;
    layer1_outputs(8634) <= a xor b;
    layer1_outputs(8635) <= not a or b;
    layer1_outputs(8636) <= not a or b;
    layer1_outputs(8637) <= not (a and b);
    layer1_outputs(8638) <= a or b;
    layer1_outputs(8639) <= 1'b1;
    layer1_outputs(8640) <= a xor b;
    layer1_outputs(8641) <= not (a or b);
    layer1_outputs(8642) <= b;
    layer1_outputs(8643) <= a xor b;
    layer1_outputs(8644) <= a xor b;
    layer1_outputs(8645) <= not b;
    layer1_outputs(8646) <= not a;
    layer1_outputs(8647) <= a;
    layer1_outputs(8648) <= not b or a;
    layer1_outputs(8649) <= not b or a;
    layer1_outputs(8650) <= not a or b;
    layer1_outputs(8651) <= not a or b;
    layer1_outputs(8652) <= not (a xor b);
    layer1_outputs(8653) <= not a;
    layer1_outputs(8654) <= not a;
    layer1_outputs(8655) <= a or b;
    layer1_outputs(8656) <= not b;
    layer1_outputs(8657) <= a;
    layer1_outputs(8658) <= not a;
    layer1_outputs(8659) <= not (a xor b);
    layer1_outputs(8660) <= a and b;
    layer1_outputs(8661) <= a;
    layer1_outputs(8662) <= b;
    layer1_outputs(8663) <= not a;
    layer1_outputs(8664) <= a;
    layer1_outputs(8665) <= a xor b;
    layer1_outputs(8666) <= not a or b;
    layer1_outputs(8667) <= not (a and b);
    layer1_outputs(8668) <= not a;
    layer1_outputs(8669) <= not a or b;
    layer1_outputs(8670) <= not a;
    layer1_outputs(8671) <= not a;
    layer1_outputs(8672) <= not b;
    layer1_outputs(8673) <= a or b;
    layer1_outputs(8674) <= not (a and b);
    layer1_outputs(8675) <= not (a or b);
    layer1_outputs(8676) <= a xor b;
    layer1_outputs(8677) <= a and not b;
    layer1_outputs(8678) <= a and not b;
    layer1_outputs(8679) <= b;
    layer1_outputs(8680) <= a;
    layer1_outputs(8681) <= not (a and b);
    layer1_outputs(8682) <= not b;
    layer1_outputs(8683) <= a or b;
    layer1_outputs(8684) <= a and b;
    layer1_outputs(8685) <= not a or b;
    layer1_outputs(8686) <= not b;
    layer1_outputs(8687) <= not (a xor b);
    layer1_outputs(8688) <= a xor b;
    layer1_outputs(8689) <= a;
    layer1_outputs(8690) <= not (a or b);
    layer1_outputs(8691) <= a and b;
    layer1_outputs(8692) <= not (a xor b);
    layer1_outputs(8693) <= not (a xor b);
    layer1_outputs(8694) <= not (a and b);
    layer1_outputs(8695) <= not (a and b);
    layer1_outputs(8696) <= b;
    layer1_outputs(8697) <= not (a xor b);
    layer1_outputs(8698) <= not b or a;
    layer1_outputs(8699) <= a and b;
    layer1_outputs(8700) <= not b or a;
    layer1_outputs(8701) <= not b;
    layer1_outputs(8702) <= a and not b;
    layer1_outputs(8703) <= not b;
    layer1_outputs(8704) <= not b;
    layer1_outputs(8705) <= a and b;
    layer1_outputs(8706) <= b;
    layer1_outputs(8707) <= b and not a;
    layer1_outputs(8708) <= not a;
    layer1_outputs(8709) <= not (a and b);
    layer1_outputs(8710) <= not b;
    layer1_outputs(8711) <= a or b;
    layer1_outputs(8712) <= a xor b;
    layer1_outputs(8713) <= not b;
    layer1_outputs(8714) <= a and not b;
    layer1_outputs(8715) <= a and not b;
    layer1_outputs(8716) <= b and not a;
    layer1_outputs(8717) <= a xor b;
    layer1_outputs(8718) <= not a or b;
    layer1_outputs(8719) <= not b or a;
    layer1_outputs(8720) <= b;
    layer1_outputs(8721) <= not a or b;
    layer1_outputs(8722) <= a and b;
    layer1_outputs(8723) <= 1'b1;
    layer1_outputs(8724) <= a or b;
    layer1_outputs(8725) <= a;
    layer1_outputs(8726) <= not b;
    layer1_outputs(8727) <= not (a or b);
    layer1_outputs(8728) <= b and not a;
    layer1_outputs(8729) <= a or b;
    layer1_outputs(8730) <= not (a or b);
    layer1_outputs(8731) <= not (a or b);
    layer1_outputs(8732) <= b and not a;
    layer1_outputs(8733) <= a and b;
    layer1_outputs(8734) <= b;
    layer1_outputs(8735) <= a xor b;
    layer1_outputs(8736) <= not (a and b);
    layer1_outputs(8737) <= a;
    layer1_outputs(8738) <= a and b;
    layer1_outputs(8739) <= not a;
    layer1_outputs(8740) <= not b;
    layer1_outputs(8741) <= not (a xor b);
    layer1_outputs(8742) <= a and b;
    layer1_outputs(8743) <= not (a xor b);
    layer1_outputs(8744) <= a or b;
    layer1_outputs(8745) <= a or b;
    layer1_outputs(8746) <= not (a and b);
    layer1_outputs(8747) <= not a;
    layer1_outputs(8748) <= a and not b;
    layer1_outputs(8749) <= not a or b;
    layer1_outputs(8750) <= not a;
    layer1_outputs(8751) <= a and b;
    layer1_outputs(8752) <= a and not b;
    layer1_outputs(8753) <= a xor b;
    layer1_outputs(8754) <= a xor b;
    layer1_outputs(8755) <= not a or b;
    layer1_outputs(8756) <= b and not a;
    layer1_outputs(8757) <= not a;
    layer1_outputs(8758) <= not b;
    layer1_outputs(8759) <= not (a xor b);
    layer1_outputs(8760) <= not b;
    layer1_outputs(8761) <= a or b;
    layer1_outputs(8762) <= a and not b;
    layer1_outputs(8763) <= not b;
    layer1_outputs(8764) <= a xor b;
    layer1_outputs(8765) <= a;
    layer1_outputs(8766) <= not (a or b);
    layer1_outputs(8767) <= b and not a;
    layer1_outputs(8768) <= a or b;
    layer1_outputs(8769) <= a or b;
    layer1_outputs(8770) <= not (a xor b);
    layer1_outputs(8771) <= not a or b;
    layer1_outputs(8772) <= not (a and b);
    layer1_outputs(8773) <= not (a xor b);
    layer1_outputs(8774) <= not (a or b);
    layer1_outputs(8775) <= not (a xor b);
    layer1_outputs(8776) <= not (a or b);
    layer1_outputs(8777) <= b and not a;
    layer1_outputs(8778) <= 1'b0;
    layer1_outputs(8779) <= not (a xor b);
    layer1_outputs(8780) <= not (a xor b);
    layer1_outputs(8781) <= a xor b;
    layer1_outputs(8782) <= a xor b;
    layer1_outputs(8783) <= not (a xor b);
    layer1_outputs(8784) <= not (a and b);
    layer1_outputs(8785) <= not b;
    layer1_outputs(8786) <= not a;
    layer1_outputs(8787) <= not (a xor b);
    layer1_outputs(8788) <= not a;
    layer1_outputs(8789) <= b and not a;
    layer1_outputs(8790) <= not a;
    layer1_outputs(8791) <= a;
    layer1_outputs(8792) <= a xor b;
    layer1_outputs(8793) <= not b;
    layer1_outputs(8794) <= not a or b;
    layer1_outputs(8795) <= a xor b;
    layer1_outputs(8796) <= a and not b;
    layer1_outputs(8797) <= not (a xor b);
    layer1_outputs(8798) <= not (a xor b);
    layer1_outputs(8799) <= 1'b1;
    layer1_outputs(8800) <= not (a xor b);
    layer1_outputs(8801) <= a or b;
    layer1_outputs(8802) <= not b or a;
    layer1_outputs(8803) <= not (a and b);
    layer1_outputs(8804) <= 1'b0;
    layer1_outputs(8805) <= a xor b;
    layer1_outputs(8806) <= a xor b;
    layer1_outputs(8807) <= not a;
    layer1_outputs(8808) <= b and not a;
    layer1_outputs(8809) <= a and not b;
    layer1_outputs(8810) <= not b;
    layer1_outputs(8811) <= not a;
    layer1_outputs(8812) <= a xor b;
    layer1_outputs(8813) <= a;
    layer1_outputs(8814) <= not a;
    layer1_outputs(8815) <= a or b;
    layer1_outputs(8816) <= a or b;
    layer1_outputs(8817) <= b and not a;
    layer1_outputs(8818) <= a and not b;
    layer1_outputs(8819) <= not a;
    layer1_outputs(8820) <= not (a xor b);
    layer1_outputs(8821) <= a and not b;
    layer1_outputs(8822) <= not (a or b);
    layer1_outputs(8823) <= a and b;
    layer1_outputs(8824) <= a and not b;
    layer1_outputs(8825) <= a or b;
    layer1_outputs(8826) <= b and not a;
    layer1_outputs(8827) <= a;
    layer1_outputs(8828) <= b;
    layer1_outputs(8829) <= not (a xor b);
    layer1_outputs(8830) <= b and not a;
    layer1_outputs(8831) <= b and not a;
    layer1_outputs(8832) <= a and not b;
    layer1_outputs(8833) <= not (a xor b);
    layer1_outputs(8834) <= not (a xor b);
    layer1_outputs(8835) <= a;
    layer1_outputs(8836) <= not (a xor b);
    layer1_outputs(8837) <= not a or b;
    layer1_outputs(8838) <= not (a or b);
    layer1_outputs(8839) <= not (a or b);
    layer1_outputs(8840) <= b;
    layer1_outputs(8841) <= a or b;
    layer1_outputs(8842) <= not a or b;
    layer1_outputs(8843) <= a and not b;
    layer1_outputs(8844) <= a and not b;
    layer1_outputs(8845) <= not b;
    layer1_outputs(8846) <= not (a or b);
    layer1_outputs(8847) <= not (a or b);
    layer1_outputs(8848) <= b and not a;
    layer1_outputs(8849) <= not (a and b);
    layer1_outputs(8850) <= not (a xor b);
    layer1_outputs(8851) <= not (a and b);
    layer1_outputs(8852) <= b;
    layer1_outputs(8853) <= a xor b;
    layer1_outputs(8854) <= not a or b;
    layer1_outputs(8855) <= not b or a;
    layer1_outputs(8856) <= a and b;
    layer1_outputs(8857) <= b;
    layer1_outputs(8858) <= not (a xor b);
    layer1_outputs(8859) <= a and b;
    layer1_outputs(8860) <= a;
    layer1_outputs(8861) <= not a or b;
    layer1_outputs(8862) <= a;
    layer1_outputs(8863) <= a;
    layer1_outputs(8864) <= a or b;
    layer1_outputs(8865) <= not b;
    layer1_outputs(8866) <= a;
    layer1_outputs(8867) <= not a;
    layer1_outputs(8868) <= a or b;
    layer1_outputs(8869) <= a and b;
    layer1_outputs(8870) <= not a;
    layer1_outputs(8871) <= not (a and b);
    layer1_outputs(8872) <= not a;
    layer1_outputs(8873) <= 1'b1;
    layer1_outputs(8874) <= a or b;
    layer1_outputs(8875) <= a and not b;
    layer1_outputs(8876) <= a xor b;
    layer1_outputs(8877) <= b;
    layer1_outputs(8878) <= b;
    layer1_outputs(8879) <= b and not a;
    layer1_outputs(8880) <= not (a and b);
    layer1_outputs(8881) <= a and b;
    layer1_outputs(8882) <= not a;
    layer1_outputs(8883) <= not (a xor b);
    layer1_outputs(8884) <= 1'b0;
    layer1_outputs(8885) <= b and not a;
    layer1_outputs(8886) <= not a or b;
    layer1_outputs(8887) <= not a or b;
    layer1_outputs(8888) <= not a;
    layer1_outputs(8889) <= b;
    layer1_outputs(8890) <= a xor b;
    layer1_outputs(8891) <= b;
    layer1_outputs(8892) <= not (a or b);
    layer1_outputs(8893) <= not a;
    layer1_outputs(8894) <= not (a or b);
    layer1_outputs(8895) <= a and b;
    layer1_outputs(8896) <= a or b;
    layer1_outputs(8897) <= not (a or b);
    layer1_outputs(8898) <= a;
    layer1_outputs(8899) <= not (a or b);
    layer1_outputs(8900) <= not a or b;
    layer1_outputs(8901) <= not a;
    layer1_outputs(8902) <= a xor b;
    layer1_outputs(8903) <= not a or b;
    layer1_outputs(8904) <= a xor b;
    layer1_outputs(8905) <= a and not b;
    layer1_outputs(8906) <= not a or b;
    layer1_outputs(8907) <= a and not b;
    layer1_outputs(8908) <= not b;
    layer1_outputs(8909) <= not a;
    layer1_outputs(8910) <= a xor b;
    layer1_outputs(8911) <= not a or b;
    layer1_outputs(8912) <= a and b;
    layer1_outputs(8913) <= 1'b1;
    layer1_outputs(8914) <= not (a and b);
    layer1_outputs(8915) <= b;
    layer1_outputs(8916) <= a and not b;
    layer1_outputs(8917) <= a and b;
    layer1_outputs(8918) <= a and not b;
    layer1_outputs(8919) <= not a;
    layer1_outputs(8920) <= 1'b0;
    layer1_outputs(8921) <= a;
    layer1_outputs(8922) <= a xor b;
    layer1_outputs(8923) <= a and b;
    layer1_outputs(8924) <= a xor b;
    layer1_outputs(8925) <= a and not b;
    layer1_outputs(8926) <= not b or a;
    layer1_outputs(8927) <= not b or a;
    layer1_outputs(8928) <= b;
    layer1_outputs(8929) <= not (a and b);
    layer1_outputs(8930) <= a xor b;
    layer1_outputs(8931) <= not b;
    layer1_outputs(8932) <= not b;
    layer1_outputs(8933) <= a;
    layer1_outputs(8934) <= a xor b;
    layer1_outputs(8935) <= not (a or b);
    layer1_outputs(8936) <= b;
    layer1_outputs(8937) <= not a;
    layer1_outputs(8938) <= not b or a;
    layer1_outputs(8939) <= a;
    layer1_outputs(8940) <= b;
    layer1_outputs(8941) <= not a;
    layer1_outputs(8942) <= a or b;
    layer1_outputs(8943) <= a or b;
    layer1_outputs(8944) <= a;
    layer1_outputs(8945) <= not (a xor b);
    layer1_outputs(8946) <= not (a xor b);
    layer1_outputs(8947) <= not (a and b);
    layer1_outputs(8948) <= b;
    layer1_outputs(8949) <= a;
    layer1_outputs(8950) <= a or b;
    layer1_outputs(8951) <= a and b;
    layer1_outputs(8952) <= not (a xor b);
    layer1_outputs(8953) <= not (a xor b);
    layer1_outputs(8954) <= b and not a;
    layer1_outputs(8955) <= 1'b1;
    layer1_outputs(8956) <= b and not a;
    layer1_outputs(8957) <= not a;
    layer1_outputs(8958) <= not a or b;
    layer1_outputs(8959) <= a;
    layer1_outputs(8960) <= not a or b;
    layer1_outputs(8961) <= a and not b;
    layer1_outputs(8962) <= not a or b;
    layer1_outputs(8963) <= a and b;
    layer1_outputs(8964) <= b;
    layer1_outputs(8965) <= b and not a;
    layer1_outputs(8966) <= not a;
    layer1_outputs(8967) <= not a;
    layer1_outputs(8968) <= not b;
    layer1_outputs(8969) <= not (a xor b);
    layer1_outputs(8970) <= not b or a;
    layer1_outputs(8971) <= not a;
    layer1_outputs(8972) <= not a;
    layer1_outputs(8973) <= not a;
    layer1_outputs(8974) <= not a or b;
    layer1_outputs(8975) <= not b;
    layer1_outputs(8976) <= a and not b;
    layer1_outputs(8977) <= not a;
    layer1_outputs(8978) <= not a;
    layer1_outputs(8979) <= b;
    layer1_outputs(8980) <= not b;
    layer1_outputs(8981) <= not b;
    layer1_outputs(8982) <= a xor b;
    layer1_outputs(8983) <= not b or a;
    layer1_outputs(8984) <= not (a or b);
    layer1_outputs(8985) <= not (a or b);
    layer1_outputs(8986) <= a and not b;
    layer1_outputs(8987) <= not (a xor b);
    layer1_outputs(8988) <= b;
    layer1_outputs(8989) <= not a;
    layer1_outputs(8990) <= b and not a;
    layer1_outputs(8991) <= not a;
    layer1_outputs(8992) <= a;
    layer1_outputs(8993) <= a and b;
    layer1_outputs(8994) <= not (a or b);
    layer1_outputs(8995) <= not (a or b);
    layer1_outputs(8996) <= not (a and b);
    layer1_outputs(8997) <= not (a xor b);
    layer1_outputs(8998) <= a xor b;
    layer1_outputs(8999) <= b;
    layer1_outputs(9000) <= a or b;
    layer1_outputs(9001) <= a;
    layer1_outputs(9002) <= not a;
    layer1_outputs(9003) <= not (a xor b);
    layer1_outputs(9004) <= not a;
    layer1_outputs(9005) <= not (a xor b);
    layer1_outputs(9006) <= not (a xor b);
    layer1_outputs(9007) <= not (a or b);
    layer1_outputs(9008) <= a;
    layer1_outputs(9009) <= a;
    layer1_outputs(9010) <= a;
    layer1_outputs(9011) <= a and b;
    layer1_outputs(9012) <= not (a and b);
    layer1_outputs(9013) <= b and not a;
    layer1_outputs(9014) <= a and b;
    layer1_outputs(9015) <= not b;
    layer1_outputs(9016) <= not (a xor b);
    layer1_outputs(9017) <= a;
    layer1_outputs(9018) <= a xor b;
    layer1_outputs(9019) <= a and b;
    layer1_outputs(9020) <= not a or b;
    layer1_outputs(9021) <= not b;
    layer1_outputs(9022) <= not (a or b);
    layer1_outputs(9023) <= b;
    layer1_outputs(9024) <= not (a and b);
    layer1_outputs(9025) <= not (a xor b);
    layer1_outputs(9026) <= not (a xor b);
    layer1_outputs(9027) <= a xor b;
    layer1_outputs(9028) <= b;
    layer1_outputs(9029) <= a and not b;
    layer1_outputs(9030) <= b and not a;
    layer1_outputs(9031) <= not b;
    layer1_outputs(9032) <= b;
    layer1_outputs(9033) <= not b;
    layer1_outputs(9034) <= a or b;
    layer1_outputs(9035) <= not b;
    layer1_outputs(9036) <= a xor b;
    layer1_outputs(9037) <= not a or b;
    layer1_outputs(9038) <= not (a or b);
    layer1_outputs(9039) <= not a;
    layer1_outputs(9040) <= a xor b;
    layer1_outputs(9041) <= not a;
    layer1_outputs(9042) <= a xor b;
    layer1_outputs(9043) <= a;
    layer1_outputs(9044) <= not (a and b);
    layer1_outputs(9045) <= not b;
    layer1_outputs(9046) <= b;
    layer1_outputs(9047) <= not a or b;
    layer1_outputs(9048) <= a and not b;
    layer1_outputs(9049) <= not (a and b);
    layer1_outputs(9050) <= not b;
    layer1_outputs(9051) <= a xor b;
    layer1_outputs(9052) <= not (a and b);
    layer1_outputs(9053) <= not a;
    layer1_outputs(9054) <= not b;
    layer1_outputs(9055) <= not (a and b);
    layer1_outputs(9056) <= not b or a;
    layer1_outputs(9057) <= b;
    layer1_outputs(9058) <= not a;
    layer1_outputs(9059) <= not (a xor b);
    layer1_outputs(9060) <= not (a xor b);
    layer1_outputs(9061) <= not (a xor b);
    layer1_outputs(9062) <= a and b;
    layer1_outputs(9063) <= not a;
    layer1_outputs(9064) <= b;
    layer1_outputs(9065) <= b and not a;
    layer1_outputs(9066) <= not a;
    layer1_outputs(9067) <= not a;
    layer1_outputs(9068) <= b and not a;
    layer1_outputs(9069) <= not (a and b);
    layer1_outputs(9070) <= not b;
    layer1_outputs(9071) <= b and not a;
    layer1_outputs(9072) <= b;
    layer1_outputs(9073) <= b and not a;
    layer1_outputs(9074) <= b;
    layer1_outputs(9075) <= not b;
    layer1_outputs(9076) <= a;
    layer1_outputs(9077) <= not b;
    layer1_outputs(9078) <= not (a or b);
    layer1_outputs(9079) <= not (a or b);
    layer1_outputs(9080) <= not a;
    layer1_outputs(9081) <= a and b;
    layer1_outputs(9082) <= b;
    layer1_outputs(9083) <= not a;
    layer1_outputs(9084) <= a xor b;
    layer1_outputs(9085) <= not (a or b);
    layer1_outputs(9086) <= not b;
    layer1_outputs(9087) <= b and not a;
    layer1_outputs(9088) <= a;
    layer1_outputs(9089) <= b;
    layer1_outputs(9090) <= b and not a;
    layer1_outputs(9091) <= not (a and b);
    layer1_outputs(9092) <= not b;
    layer1_outputs(9093) <= not (a or b);
    layer1_outputs(9094) <= not b or a;
    layer1_outputs(9095) <= b;
    layer1_outputs(9096) <= a;
    layer1_outputs(9097) <= 1'b1;
    layer1_outputs(9098) <= not b;
    layer1_outputs(9099) <= not (a or b);
    layer1_outputs(9100) <= not (a xor b);
    layer1_outputs(9101) <= not a;
    layer1_outputs(9102) <= not b or a;
    layer1_outputs(9103) <= b;
    layer1_outputs(9104) <= 1'b0;
    layer1_outputs(9105) <= not a or b;
    layer1_outputs(9106) <= b;
    layer1_outputs(9107) <= not b;
    layer1_outputs(9108) <= not (a or b);
    layer1_outputs(9109) <= not (a xor b);
    layer1_outputs(9110) <= a or b;
    layer1_outputs(9111) <= a xor b;
    layer1_outputs(9112) <= a and not b;
    layer1_outputs(9113) <= not b or a;
    layer1_outputs(9114) <= not b or a;
    layer1_outputs(9115) <= not b;
    layer1_outputs(9116) <= b and not a;
    layer1_outputs(9117) <= not (a or b);
    layer1_outputs(9118) <= not b;
    layer1_outputs(9119) <= a;
    layer1_outputs(9120) <= not a or b;
    layer1_outputs(9121) <= not b;
    layer1_outputs(9122) <= not (a xor b);
    layer1_outputs(9123) <= not a;
    layer1_outputs(9124) <= a xor b;
    layer1_outputs(9125) <= 1'b0;
    layer1_outputs(9126) <= not (a xor b);
    layer1_outputs(9127) <= not (a xor b);
    layer1_outputs(9128) <= b;
    layer1_outputs(9129) <= a and b;
    layer1_outputs(9130) <= not (a and b);
    layer1_outputs(9131) <= not a;
    layer1_outputs(9132) <= a or b;
    layer1_outputs(9133) <= b;
    layer1_outputs(9134) <= 1'b1;
    layer1_outputs(9135) <= a and b;
    layer1_outputs(9136) <= b;
    layer1_outputs(9137) <= b and not a;
    layer1_outputs(9138) <= not b;
    layer1_outputs(9139) <= a xor b;
    layer1_outputs(9140) <= a or b;
    layer1_outputs(9141) <= b;
    layer1_outputs(9142) <= a xor b;
    layer1_outputs(9143) <= not (a and b);
    layer1_outputs(9144) <= not (a and b);
    layer1_outputs(9145) <= not (a or b);
    layer1_outputs(9146) <= not b;
    layer1_outputs(9147) <= a xor b;
    layer1_outputs(9148) <= not b;
    layer1_outputs(9149) <= a and b;
    layer1_outputs(9150) <= a or b;
    layer1_outputs(9151) <= not b;
    layer1_outputs(9152) <= not (a and b);
    layer1_outputs(9153) <= not a or b;
    layer1_outputs(9154) <= not b;
    layer1_outputs(9155) <= not (a xor b);
    layer1_outputs(9156) <= not a or b;
    layer1_outputs(9157) <= not (a or b);
    layer1_outputs(9158) <= not b;
    layer1_outputs(9159) <= not b or a;
    layer1_outputs(9160) <= not a;
    layer1_outputs(9161) <= not a or b;
    layer1_outputs(9162) <= b;
    layer1_outputs(9163) <= a;
    layer1_outputs(9164) <= not (a xor b);
    layer1_outputs(9165) <= not b or a;
    layer1_outputs(9166) <= b;
    layer1_outputs(9167) <= not b;
    layer1_outputs(9168) <= not a or b;
    layer1_outputs(9169) <= a xor b;
    layer1_outputs(9170) <= a and not b;
    layer1_outputs(9171) <= a or b;
    layer1_outputs(9172) <= a xor b;
    layer1_outputs(9173) <= a;
    layer1_outputs(9174) <= not a or b;
    layer1_outputs(9175) <= not b or a;
    layer1_outputs(9176) <= a or b;
    layer1_outputs(9177) <= b and not a;
    layer1_outputs(9178) <= b;
    layer1_outputs(9179) <= not (a xor b);
    layer1_outputs(9180) <= not b or a;
    layer1_outputs(9181) <= not (a and b);
    layer1_outputs(9182) <= not a;
    layer1_outputs(9183) <= a and not b;
    layer1_outputs(9184) <= a and b;
    layer1_outputs(9185) <= a;
    layer1_outputs(9186) <= a;
    layer1_outputs(9187) <= a;
    layer1_outputs(9188) <= b and not a;
    layer1_outputs(9189) <= not (a xor b);
    layer1_outputs(9190) <= a and b;
    layer1_outputs(9191) <= b;
    layer1_outputs(9192) <= not (a and b);
    layer1_outputs(9193) <= not (a or b);
    layer1_outputs(9194) <= not b or a;
    layer1_outputs(9195) <= b;
    layer1_outputs(9196) <= a;
    layer1_outputs(9197) <= not (a and b);
    layer1_outputs(9198) <= b;
    layer1_outputs(9199) <= b and not a;
    layer1_outputs(9200) <= a xor b;
    layer1_outputs(9201) <= b;
    layer1_outputs(9202) <= not (a or b);
    layer1_outputs(9203) <= a and b;
    layer1_outputs(9204) <= a xor b;
    layer1_outputs(9205) <= a;
    layer1_outputs(9206) <= not a;
    layer1_outputs(9207) <= not (a or b);
    layer1_outputs(9208) <= not b;
    layer1_outputs(9209) <= a;
    layer1_outputs(9210) <= 1'b1;
    layer1_outputs(9211) <= not a or b;
    layer1_outputs(9212) <= not (a or b);
    layer1_outputs(9213) <= not a;
    layer1_outputs(9214) <= a;
    layer1_outputs(9215) <= a or b;
    layer1_outputs(9216) <= not a;
    layer1_outputs(9217) <= not (a and b);
    layer1_outputs(9218) <= a or b;
    layer1_outputs(9219) <= not b or a;
    layer1_outputs(9220) <= not a or b;
    layer1_outputs(9221) <= a;
    layer1_outputs(9222) <= a;
    layer1_outputs(9223) <= a;
    layer1_outputs(9224) <= a and b;
    layer1_outputs(9225) <= not a;
    layer1_outputs(9226) <= a;
    layer1_outputs(9227) <= b and not a;
    layer1_outputs(9228) <= not a;
    layer1_outputs(9229) <= a xor b;
    layer1_outputs(9230) <= not (a and b);
    layer1_outputs(9231) <= a;
    layer1_outputs(9232) <= b;
    layer1_outputs(9233) <= a and not b;
    layer1_outputs(9234) <= not a;
    layer1_outputs(9235) <= not (a and b);
    layer1_outputs(9236) <= a or b;
    layer1_outputs(9237) <= a or b;
    layer1_outputs(9238) <= not (a and b);
    layer1_outputs(9239) <= not (a and b);
    layer1_outputs(9240) <= a and b;
    layer1_outputs(9241) <= a or b;
    layer1_outputs(9242) <= not a;
    layer1_outputs(9243) <= a xor b;
    layer1_outputs(9244) <= b and not a;
    layer1_outputs(9245) <= a xor b;
    layer1_outputs(9246) <= a xor b;
    layer1_outputs(9247) <= a and not b;
    layer1_outputs(9248) <= not b;
    layer1_outputs(9249) <= a;
    layer1_outputs(9250) <= 1'b0;
    layer1_outputs(9251) <= not (a xor b);
    layer1_outputs(9252) <= a xor b;
    layer1_outputs(9253) <= a and not b;
    layer1_outputs(9254) <= b;
    layer1_outputs(9255) <= b;
    layer1_outputs(9256) <= 1'b0;
    layer1_outputs(9257) <= not b or a;
    layer1_outputs(9258) <= 1'b0;
    layer1_outputs(9259) <= not a;
    layer1_outputs(9260) <= not b;
    layer1_outputs(9261) <= a xor b;
    layer1_outputs(9262) <= a and not b;
    layer1_outputs(9263) <= not (a or b);
    layer1_outputs(9264) <= a xor b;
    layer1_outputs(9265) <= not a;
    layer1_outputs(9266) <= not (a or b);
    layer1_outputs(9267) <= not a;
    layer1_outputs(9268) <= not a or b;
    layer1_outputs(9269) <= not a;
    layer1_outputs(9270) <= b and not a;
    layer1_outputs(9271) <= 1'b1;
    layer1_outputs(9272) <= not a;
    layer1_outputs(9273) <= a and b;
    layer1_outputs(9274) <= not (a or b);
    layer1_outputs(9275) <= a and b;
    layer1_outputs(9276) <= a and b;
    layer1_outputs(9277) <= not a;
    layer1_outputs(9278) <= not (a xor b);
    layer1_outputs(9279) <= a xor b;
    layer1_outputs(9280) <= 1'b1;
    layer1_outputs(9281) <= not (a or b);
    layer1_outputs(9282) <= not (a and b);
    layer1_outputs(9283) <= not b;
    layer1_outputs(9284) <= not (a xor b);
    layer1_outputs(9285) <= not b or a;
    layer1_outputs(9286) <= a xor b;
    layer1_outputs(9287) <= 1'b0;
    layer1_outputs(9288) <= not a or b;
    layer1_outputs(9289) <= not a;
    layer1_outputs(9290) <= b and not a;
    layer1_outputs(9291) <= not (a or b);
    layer1_outputs(9292) <= 1'b0;
    layer1_outputs(9293) <= not (a xor b);
    layer1_outputs(9294) <= not (a xor b);
    layer1_outputs(9295) <= a and not b;
    layer1_outputs(9296) <= not b;
    layer1_outputs(9297) <= not (a xor b);
    layer1_outputs(9298) <= not (a xor b);
    layer1_outputs(9299) <= not (a or b);
    layer1_outputs(9300) <= not b;
    layer1_outputs(9301) <= not a;
    layer1_outputs(9302) <= b and not a;
    layer1_outputs(9303) <= not a or b;
    layer1_outputs(9304) <= b and not a;
    layer1_outputs(9305) <= b;
    layer1_outputs(9306) <= not (a xor b);
    layer1_outputs(9307) <= not (a and b);
    layer1_outputs(9308) <= a and not b;
    layer1_outputs(9309) <= not a;
    layer1_outputs(9310) <= not a or b;
    layer1_outputs(9311) <= a and b;
    layer1_outputs(9312) <= a or b;
    layer1_outputs(9313) <= not b or a;
    layer1_outputs(9314) <= not (a xor b);
    layer1_outputs(9315) <= not (a or b);
    layer1_outputs(9316) <= a and b;
    layer1_outputs(9317) <= b and not a;
    layer1_outputs(9318) <= not b or a;
    layer1_outputs(9319) <= a xor b;
    layer1_outputs(9320) <= not a or b;
    layer1_outputs(9321) <= a and not b;
    layer1_outputs(9322) <= 1'b0;
    layer1_outputs(9323) <= not a or b;
    layer1_outputs(9324) <= not (a xor b);
    layer1_outputs(9325) <= not (a and b);
    layer1_outputs(9326) <= not a or b;
    layer1_outputs(9327) <= not (a xor b);
    layer1_outputs(9328) <= a or b;
    layer1_outputs(9329) <= not a;
    layer1_outputs(9330) <= not a or b;
    layer1_outputs(9331) <= b and not a;
    layer1_outputs(9332) <= b and not a;
    layer1_outputs(9333) <= b;
    layer1_outputs(9334) <= not a or b;
    layer1_outputs(9335) <= not a;
    layer1_outputs(9336) <= a xor b;
    layer1_outputs(9337) <= not a;
    layer1_outputs(9338) <= not (a and b);
    layer1_outputs(9339) <= a xor b;
    layer1_outputs(9340) <= b;
    layer1_outputs(9341) <= b;
    layer1_outputs(9342) <= a and b;
    layer1_outputs(9343) <= a and not b;
    layer1_outputs(9344) <= a or b;
    layer1_outputs(9345) <= a;
    layer1_outputs(9346) <= not (a and b);
    layer1_outputs(9347) <= not (a xor b);
    layer1_outputs(9348) <= not b;
    layer1_outputs(9349) <= a;
    layer1_outputs(9350) <= not b or a;
    layer1_outputs(9351) <= not a;
    layer1_outputs(9352) <= a or b;
    layer1_outputs(9353) <= not a;
    layer1_outputs(9354) <= not (a xor b);
    layer1_outputs(9355) <= a xor b;
    layer1_outputs(9356) <= a xor b;
    layer1_outputs(9357) <= b and not a;
    layer1_outputs(9358) <= not b;
    layer1_outputs(9359) <= a xor b;
    layer1_outputs(9360) <= not b or a;
    layer1_outputs(9361) <= 1'b0;
    layer1_outputs(9362) <= a xor b;
    layer1_outputs(9363) <= b;
    layer1_outputs(9364) <= a xor b;
    layer1_outputs(9365) <= not a or b;
    layer1_outputs(9366) <= not (a and b);
    layer1_outputs(9367) <= b;
    layer1_outputs(9368) <= not (a xor b);
    layer1_outputs(9369) <= a;
    layer1_outputs(9370) <= not b;
    layer1_outputs(9371) <= a xor b;
    layer1_outputs(9372) <= a and b;
    layer1_outputs(9373) <= a xor b;
    layer1_outputs(9374) <= a xor b;
    layer1_outputs(9375) <= b;
    layer1_outputs(9376) <= not (a xor b);
    layer1_outputs(9377) <= not a;
    layer1_outputs(9378) <= not (a or b);
    layer1_outputs(9379) <= not a or b;
    layer1_outputs(9380) <= a and not b;
    layer1_outputs(9381) <= a and b;
    layer1_outputs(9382) <= not b;
    layer1_outputs(9383) <= b;
    layer1_outputs(9384) <= a and b;
    layer1_outputs(9385) <= a xor b;
    layer1_outputs(9386) <= not a or b;
    layer1_outputs(9387) <= not b or a;
    layer1_outputs(9388) <= a and b;
    layer1_outputs(9389) <= not a or b;
    layer1_outputs(9390) <= not b;
    layer1_outputs(9391) <= not (a or b);
    layer1_outputs(9392) <= not a;
    layer1_outputs(9393) <= b;
    layer1_outputs(9394) <= not b or a;
    layer1_outputs(9395) <= a xor b;
    layer1_outputs(9396) <= not a;
    layer1_outputs(9397) <= not (a xor b);
    layer1_outputs(9398) <= not a;
    layer1_outputs(9399) <= not (a or b);
    layer1_outputs(9400) <= a;
    layer1_outputs(9401) <= a xor b;
    layer1_outputs(9402) <= a xor b;
    layer1_outputs(9403) <= a and b;
    layer1_outputs(9404) <= not b;
    layer1_outputs(9405) <= not a;
    layer1_outputs(9406) <= a and b;
    layer1_outputs(9407) <= not a;
    layer1_outputs(9408) <= not (a or b);
    layer1_outputs(9409) <= b and not a;
    layer1_outputs(9410) <= b;
    layer1_outputs(9411) <= not a;
    layer1_outputs(9412) <= not (a xor b);
    layer1_outputs(9413) <= not a;
    layer1_outputs(9414) <= a and b;
    layer1_outputs(9415) <= not a;
    layer1_outputs(9416) <= a and not b;
    layer1_outputs(9417) <= not b or a;
    layer1_outputs(9418) <= a and not b;
    layer1_outputs(9419) <= a or b;
    layer1_outputs(9420) <= a or b;
    layer1_outputs(9421) <= a and b;
    layer1_outputs(9422) <= not a;
    layer1_outputs(9423) <= a;
    layer1_outputs(9424) <= not a or b;
    layer1_outputs(9425) <= not b or a;
    layer1_outputs(9426) <= a xor b;
    layer1_outputs(9427) <= a or b;
    layer1_outputs(9428) <= not b or a;
    layer1_outputs(9429) <= not b;
    layer1_outputs(9430) <= a;
    layer1_outputs(9431) <= not (a or b);
    layer1_outputs(9432) <= b and not a;
    layer1_outputs(9433) <= a xor b;
    layer1_outputs(9434) <= 1'b1;
    layer1_outputs(9435) <= a xor b;
    layer1_outputs(9436) <= not a;
    layer1_outputs(9437) <= b and not a;
    layer1_outputs(9438) <= not b;
    layer1_outputs(9439) <= not b or a;
    layer1_outputs(9440) <= a;
    layer1_outputs(9441) <= b;
    layer1_outputs(9442) <= not b or a;
    layer1_outputs(9443) <= not (a xor b);
    layer1_outputs(9444) <= not a;
    layer1_outputs(9445) <= a;
    layer1_outputs(9446) <= not (a and b);
    layer1_outputs(9447) <= a and b;
    layer1_outputs(9448) <= a xor b;
    layer1_outputs(9449) <= not (a or b);
    layer1_outputs(9450) <= a and b;
    layer1_outputs(9451) <= not (a or b);
    layer1_outputs(9452) <= not b or a;
    layer1_outputs(9453) <= b and not a;
    layer1_outputs(9454) <= b and not a;
    layer1_outputs(9455) <= a xor b;
    layer1_outputs(9456) <= a and b;
    layer1_outputs(9457) <= not b or a;
    layer1_outputs(9458) <= not (a and b);
    layer1_outputs(9459) <= not a;
    layer1_outputs(9460) <= a or b;
    layer1_outputs(9461) <= not b;
    layer1_outputs(9462) <= a and not b;
    layer1_outputs(9463) <= 1'b0;
    layer1_outputs(9464) <= not (a and b);
    layer1_outputs(9465) <= not (a or b);
    layer1_outputs(9466) <= not (a or b);
    layer1_outputs(9467) <= not (a and b);
    layer1_outputs(9468) <= a or b;
    layer1_outputs(9469) <= not (a and b);
    layer1_outputs(9470) <= a;
    layer1_outputs(9471) <= 1'b0;
    layer1_outputs(9472) <= a;
    layer1_outputs(9473) <= a;
    layer1_outputs(9474) <= 1'b1;
    layer1_outputs(9475) <= not b;
    layer1_outputs(9476) <= not b;
    layer1_outputs(9477) <= b;
    layer1_outputs(9478) <= not b;
    layer1_outputs(9479) <= not (a or b);
    layer1_outputs(9480) <= not b or a;
    layer1_outputs(9481) <= a xor b;
    layer1_outputs(9482) <= not a or b;
    layer1_outputs(9483) <= a;
    layer1_outputs(9484) <= not a;
    layer1_outputs(9485) <= a xor b;
    layer1_outputs(9486) <= not (a or b);
    layer1_outputs(9487) <= not (a xor b);
    layer1_outputs(9488) <= b;
    layer1_outputs(9489) <= a and not b;
    layer1_outputs(9490) <= a;
    layer1_outputs(9491) <= a;
    layer1_outputs(9492) <= not (a xor b);
    layer1_outputs(9493) <= b;
    layer1_outputs(9494) <= not a;
    layer1_outputs(9495) <= a and not b;
    layer1_outputs(9496) <= not b;
    layer1_outputs(9497) <= a or b;
    layer1_outputs(9498) <= not (a and b);
    layer1_outputs(9499) <= not a;
    layer1_outputs(9500) <= a xor b;
    layer1_outputs(9501) <= a and not b;
    layer1_outputs(9502) <= a xor b;
    layer1_outputs(9503) <= not b or a;
    layer1_outputs(9504) <= a and not b;
    layer1_outputs(9505) <= b;
    layer1_outputs(9506) <= a;
    layer1_outputs(9507) <= not a or b;
    layer1_outputs(9508) <= not b;
    layer1_outputs(9509) <= b and not a;
    layer1_outputs(9510) <= not (a or b);
    layer1_outputs(9511) <= b;
    layer1_outputs(9512) <= not (a and b);
    layer1_outputs(9513) <= b;
    layer1_outputs(9514) <= not a;
    layer1_outputs(9515) <= not a or b;
    layer1_outputs(9516) <= not (a and b);
    layer1_outputs(9517) <= a xor b;
    layer1_outputs(9518) <= a or b;
    layer1_outputs(9519) <= not b;
    layer1_outputs(9520) <= a;
    layer1_outputs(9521) <= a;
    layer1_outputs(9522) <= not (a or b);
    layer1_outputs(9523) <= a or b;
    layer1_outputs(9524) <= not a;
    layer1_outputs(9525) <= not (a xor b);
    layer1_outputs(9526) <= b;
    layer1_outputs(9527) <= a or b;
    layer1_outputs(9528) <= not b;
    layer1_outputs(9529) <= not a;
    layer1_outputs(9530) <= b and not a;
    layer1_outputs(9531) <= a;
    layer1_outputs(9532) <= a or b;
    layer1_outputs(9533) <= b;
    layer1_outputs(9534) <= not a;
    layer1_outputs(9535) <= not (a or b);
    layer1_outputs(9536) <= a and b;
    layer1_outputs(9537) <= not a;
    layer1_outputs(9538) <= a or b;
    layer1_outputs(9539) <= a xor b;
    layer1_outputs(9540) <= not (a or b);
    layer1_outputs(9541) <= a and not b;
    layer1_outputs(9542) <= not (a xor b);
    layer1_outputs(9543) <= b and not a;
    layer1_outputs(9544) <= a xor b;
    layer1_outputs(9545) <= 1'b1;
    layer1_outputs(9546) <= a or b;
    layer1_outputs(9547) <= a;
    layer1_outputs(9548) <= a;
    layer1_outputs(9549) <= not b or a;
    layer1_outputs(9550) <= not a or b;
    layer1_outputs(9551) <= not a;
    layer1_outputs(9552) <= not (a xor b);
    layer1_outputs(9553) <= a and not b;
    layer1_outputs(9554) <= a and b;
    layer1_outputs(9555) <= not (a xor b);
    layer1_outputs(9556) <= b and not a;
    layer1_outputs(9557) <= a xor b;
    layer1_outputs(9558) <= a;
    layer1_outputs(9559) <= not (a xor b);
    layer1_outputs(9560) <= b;
    layer1_outputs(9561) <= not b or a;
    layer1_outputs(9562) <= not (a and b);
    layer1_outputs(9563) <= not (a xor b);
    layer1_outputs(9564) <= not (a xor b);
    layer1_outputs(9565) <= not b or a;
    layer1_outputs(9566) <= b and not a;
    layer1_outputs(9567) <= a;
    layer1_outputs(9568) <= not b;
    layer1_outputs(9569) <= a xor b;
    layer1_outputs(9570) <= a xor b;
    layer1_outputs(9571) <= not a;
    layer1_outputs(9572) <= a or b;
    layer1_outputs(9573) <= not (a or b);
    layer1_outputs(9574) <= b;
    layer1_outputs(9575) <= not (a and b);
    layer1_outputs(9576) <= not b;
    layer1_outputs(9577) <= a and b;
    layer1_outputs(9578) <= b;
    layer1_outputs(9579) <= a and not b;
    layer1_outputs(9580) <= b;
    layer1_outputs(9581) <= not (a or b);
    layer1_outputs(9582) <= not b or a;
    layer1_outputs(9583) <= not a;
    layer1_outputs(9584) <= not (a xor b);
    layer1_outputs(9585) <= 1'b1;
    layer1_outputs(9586) <= not (a xor b);
    layer1_outputs(9587) <= not (a and b);
    layer1_outputs(9588) <= a and not b;
    layer1_outputs(9589) <= not a or b;
    layer1_outputs(9590) <= not b or a;
    layer1_outputs(9591) <= a or b;
    layer1_outputs(9592) <= not (a and b);
    layer1_outputs(9593) <= a;
    layer1_outputs(9594) <= not a or b;
    layer1_outputs(9595) <= not b;
    layer1_outputs(9596) <= a xor b;
    layer1_outputs(9597) <= a or b;
    layer1_outputs(9598) <= 1'b1;
    layer1_outputs(9599) <= not (a and b);
    layer1_outputs(9600) <= not a or b;
    layer1_outputs(9601) <= b;
    layer1_outputs(9602) <= not b or a;
    layer1_outputs(9603) <= not b;
    layer1_outputs(9604) <= b;
    layer1_outputs(9605) <= not (a xor b);
    layer1_outputs(9606) <= not (a or b);
    layer1_outputs(9607) <= a;
    layer1_outputs(9608) <= not (a and b);
    layer1_outputs(9609) <= not (a xor b);
    layer1_outputs(9610) <= b;
    layer1_outputs(9611) <= not b or a;
    layer1_outputs(9612) <= a or b;
    layer1_outputs(9613) <= not (a xor b);
    layer1_outputs(9614) <= not b or a;
    layer1_outputs(9615) <= not (a or b);
    layer1_outputs(9616) <= not a;
    layer1_outputs(9617) <= not (a or b);
    layer1_outputs(9618) <= 1'b1;
    layer1_outputs(9619) <= not (a xor b);
    layer1_outputs(9620) <= a and not b;
    layer1_outputs(9621) <= b;
    layer1_outputs(9622) <= not a;
    layer1_outputs(9623) <= a;
    layer1_outputs(9624) <= a and not b;
    layer1_outputs(9625) <= a;
    layer1_outputs(9626) <= a xor b;
    layer1_outputs(9627) <= b;
    layer1_outputs(9628) <= a or b;
    layer1_outputs(9629) <= not a;
    layer1_outputs(9630) <= not a or b;
    layer1_outputs(9631) <= b;
    layer1_outputs(9632) <= b;
    layer1_outputs(9633) <= not (a xor b);
    layer1_outputs(9634) <= a and not b;
    layer1_outputs(9635) <= not b;
    layer1_outputs(9636) <= not b;
    layer1_outputs(9637) <= a and not b;
    layer1_outputs(9638) <= not (a or b);
    layer1_outputs(9639) <= b;
    layer1_outputs(9640) <= a;
    layer1_outputs(9641) <= a and not b;
    layer1_outputs(9642) <= b and not a;
    layer1_outputs(9643) <= a and b;
    layer1_outputs(9644) <= b;
    layer1_outputs(9645) <= not b;
    layer1_outputs(9646) <= not (a and b);
    layer1_outputs(9647) <= not b;
    layer1_outputs(9648) <= a xor b;
    layer1_outputs(9649) <= not (a xor b);
    layer1_outputs(9650) <= 1'b0;
    layer1_outputs(9651) <= not (a xor b);
    layer1_outputs(9652) <= a or b;
    layer1_outputs(9653) <= 1'b1;
    layer1_outputs(9654) <= b;
    layer1_outputs(9655) <= a or b;
    layer1_outputs(9656) <= not b or a;
    layer1_outputs(9657) <= not (a and b);
    layer1_outputs(9658) <= a and b;
    layer1_outputs(9659) <= a xor b;
    layer1_outputs(9660) <= a and not b;
    layer1_outputs(9661) <= a and b;
    layer1_outputs(9662) <= a;
    layer1_outputs(9663) <= not (a xor b);
    layer1_outputs(9664) <= not a or b;
    layer1_outputs(9665) <= b and not a;
    layer1_outputs(9666) <= not (a or b);
    layer1_outputs(9667) <= not a or b;
    layer1_outputs(9668) <= not (a or b);
    layer1_outputs(9669) <= b and not a;
    layer1_outputs(9670) <= not (a and b);
    layer1_outputs(9671) <= not (a and b);
    layer1_outputs(9672) <= a and not b;
    layer1_outputs(9673) <= not a;
    layer1_outputs(9674) <= not a;
    layer1_outputs(9675) <= not b;
    layer1_outputs(9676) <= b and not a;
    layer1_outputs(9677) <= not b or a;
    layer1_outputs(9678) <= a and b;
    layer1_outputs(9679) <= b and not a;
    layer1_outputs(9680) <= not (a and b);
    layer1_outputs(9681) <= not b or a;
    layer1_outputs(9682) <= a or b;
    layer1_outputs(9683) <= not (a xor b);
    layer1_outputs(9684) <= a;
    layer1_outputs(9685) <= not (a or b);
    layer1_outputs(9686) <= not (a xor b);
    layer1_outputs(9687) <= not b;
    layer1_outputs(9688) <= not a or b;
    layer1_outputs(9689) <= not (a or b);
    layer1_outputs(9690) <= a;
    layer1_outputs(9691) <= a;
    layer1_outputs(9692) <= not a;
    layer1_outputs(9693) <= b;
    layer1_outputs(9694) <= b and not a;
    layer1_outputs(9695) <= not (a xor b);
    layer1_outputs(9696) <= a or b;
    layer1_outputs(9697) <= not (a xor b);
    layer1_outputs(9698) <= not a;
    layer1_outputs(9699) <= not (a xor b);
    layer1_outputs(9700) <= 1'b0;
    layer1_outputs(9701) <= not (a or b);
    layer1_outputs(9702) <= a or b;
    layer1_outputs(9703) <= a;
    layer1_outputs(9704) <= a or b;
    layer1_outputs(9705) <= not a;
    layer1_outputs(9706) <= not a;
    layer1_outputs(9707) <= a and not b;
    layer1_outputs(9708) <= not (a xor b);
    layer1_outputs(9709) <= a xor b;
    layer1_outputs(9710) <= a xor b;
    layer1_outputs(9711) <= not b;
    layer1_outputs(9712) <= not (a and b);
    layer1_outputs(9713) <= not a;
    layer1_outputs(9714) <= a;
    layer1_outputs(9715) <= a or b;
    layer1_outputs(9716) <= b and not a;
    layer1_outputs(9717) <= b;
    layer1_outputs(9718) <= not (a xor b);
    layer1_outputs(9719) <= b;
    layer1_outputs(9720) <= not (a and b);
    layer1_outputs(9721) <= not (a and b);
    layer1_outputs(9722) <= not a or b;
    layer1_outputs(9723) <= not a;
    layer1_outputs(9724) <= 1'b1;
    layer1_outputs(9725) <= not (a or b);
    layer1_outputs(9726) <= a and not b;
    layer1_outputs(9727) <= a xor b;
    layer1_outputs(9728) <= not b or a;
    layer1_outputs(9729) <= not (a or b);
    layer1_outputs(9730) <= not b;
    layer1_outputs(9731) <= not a;
    layer1_outputs(9732) <= not (a and b);
    layer1_outputs(9733) <= not b;
    layer1_outputs(9734) <= not (a and b);
    layer1_outputs(9735) <= not b;
    layer1_outputs(9736) <= a and b;
    layer1_outputs(9737) <= a and not b;
    layer1_outputs(9738) <= 1'b0;
    layer1_outputs(9739) <= not b or a;
    layer1_outputs(9740) <= not (a xor b);
    layer1_outputs(9741) <= not a;
    layer1_outputs(9742) <= a;
    layer1_outputs(9743) <= not a;
    layer1_outputs(9744) <= a and not b;
    layer1_outputs(9745) <= 1'b0;
    layer1_outputs(9746) <= b;
    layer1_outputs(9747) <= not a or b;
    layer1_outputs(9748) <= b and not a;
    layer1_outputs(9749) <= b;
    layer1_outputs(9750) <= not b or a;
    layer1_outputs(9751) <= a and not b;
    layer1_outputs(9752) <= b and not a;
    layer1_outputs(9753) <= a xor b;
    layer1_outputs(9754) <= not a;
    layer1_outputs(9755) <= b and not a;
    layer1_outputs(9756) <= not (a and b);
    layer1_outputs(9757) <= not a or b;
    layer1_outputs(9758) <= a and b;
    layer1_outputs(9759) <= not b;
    layer1_outputs(9760) <= a and b;
    layer1_outputs(9761) <= b and not a;
    layer1_outputs(9762) <= b and not a;
    layer1_outputs(9763) <= a;
    layer1_outputs(9764) <= a and b;
    layer1_outputs(9765) <= b;
    layer1_outputs(9766) <= not (a xor b);
    layer1_outputs(9767) <= not (a and b);
    layer1_outputs(9768) <= not (a and b);
    layer1_outputs(9769) <= not b;
    layer1_outputs(9770) <= b;
    layer1_outputs(9771) <= not (a xor b);
    layer1_outputs(9772) <= not b;
    layer1_outputs(9773) <= a xor b;
    layer1_outputs(9774) <= not (a or b);
    layer1_outputs(9775) <= a and not b;
    layer1_outputs(9776) <= a;
    layer1_outputs(9777) <= not (a or b);
    layer1_outputs(9778) <= not (a xor b);
    layer1_outputs(9779) <= a and not b;
    layer1_outputs(9780) <= not a or b;
    layer1_outputs(9781) <= b and not a;
    layer1_outputs(9782) <= a or b;
    layer1_outputs(9783) <= a xor b;
    layer1_outputs(9784) <= a;
    layer1_outputs(9785) <= not a or b;
    layer1_outputs(9786) <= not b or a;
    layer1_outputs(9787) <= not a or b;
    layer1_outputs(9788) <= not (a or b);
    layer1_outputs(9789) <= not (a xor b);
    layer1_outputs(9790) <= a and b;
    layer1_outputs(9791) <= not (a or b);
    layer1_outputs(9792) <= not a;
    layer1_outputs(9793) <= a and not b;
    layer1_outputs(9794) <= a xor b;
    layer1_outputs(9795) <= not (a xor b);
    layer1_outputs(9796) <= not b or a;
    layer1_outputs(9797) <= not a;
    layer1_outputs(9798) <= a and not b;
    layer1_outputs(9799) <= not (a xor b);
    layer1_outputs(9800) <= not a;
    layer1_outputs(9801) <= a;
    layer1_outputs(9802) <= not (a or b);
    layer1_outputs(9803) <= not (a xor b);
    layer1_outputs(9804) <= not a;
    layer1_outputs(9805) <= a and not b;
    layer1_outputs(9806) <= not a or b;
    layer1_outputs(9807) <= a and not b;
    layer1_outputs(9808) <= b and not a;
    layer1_outputs(9809) <= b;
    layer1_outputs(9810) <= a or b;
    layer1_outputs(9811) <= not b;
    layer1_outputs(9812) <= b and not a;
    layer1_outputs(9813) <= a or b;
    layer1_outputs(9814) <= not (a xor b);
    layer1_outputs(9815) <= not (a xor b);
    layer1_outputs(9816) <= a and b;
    layer1_outputs(9817) <= b;
    layer1_outputs(9818) <= a xor b;
    layer1_outputs(9819) <= a or b;
    layer1_outputs(9820) <= b;
    layer1_outputs(9821) <= not a;
    layer1_outputs(9822) <= a or b;
    layer1_outputs(9823) <= b and not a;
    layer1_outputs(9824) <= not (a or b);
    layer1_outputs(9825) <= not (a or b);
    layer1_outputs(9826) <= a xor b;
    layer1_outputs(9827) <= not (a or b);
    layer1_outputs(9828) <= a or b;
    layer1_outputs(9829) <= b and not a;
    layer1_outputs(9830) <= a xor b;
    layer1_outputs(9831) <= not a or b;
    layer1_outputs(9832) <= b and not a;
    layer1_outputs(9833) <= not (a xor b);
    layer1_outputs(9834) <= b and not a;
    layer1_outputs(9835) <= a;
    layer1_outputs(9836) <= not a or b;
    layer1_outputs(9837) <= not b;
    layer1_outputs(9838) <= a and b;
    layer1_outputs(9839) <= a and not b;
    layer1_outputs(9840) <= a;
    layer1_outputs(9841) <= a;
    layer1_outputs(9842) <= not a;
    layer1_outputs(9843) <= a and not b;
    layer1_outputs(9844) <= not (a or b);
    layer1_outputs(9845) <= not a;
    layer1_outputs(9846) <= b;
    layer1_outputs(9847) <= not b;
    layer1_outputs(9848) <= not a or b;
    layer1_outputs(9849) <= not b or a;
    layer1_outputs(9850) <= not b;
    layer1_outputs(9851) <= a and b;
    layer1_outputs(9852) <= b;
    layer1_outputs(9853) <= not a or b;
    layer1_outputs(9854) <= a;
    layer1_outputs(9855) <= a;
    layer1_outputs(9856) <= not (a and b);
    layer1_outputs(9857) <= a;
    layer1_outputs(9858) <= not (a and b);
    layer1_outputs(9859) <= not (a or b);
    layer1_outputs(9860) <= not (a and b);
    layer1_outputs(9861) <= a;
    layer1_outputs(9862) <= not b or a;
    layer1_outputs(9863) <= a and b;
    layer1_outputs(9864) <= not (a or b);
    layer1_outputs(9865) <= 1'b0;
    layer1_outputs(9866) <= not a;
    layer1_outputs(9867) <= b;
    layer1_outputs(9868) <= not (a and b);
    layer1_outputs(9869) <= not b;
    layer1_outputs(9870) <= a and b;
    layer1_outputs(9871) <= a;
    layer1_outputs(9872) <= not (a or b);
    layer1_outputs(9873) <= a;
    layer1_outputs(9874) <= b;
    layer1_outputs(9875) <= b;
    layer1_outputs(9876) <= b and not a;
    layer1_outputs(9877) <= not (a and b);
    layer1_outputs(9878) <= b;
    layer1_outputs(9879) <= not b or a;
    layer1_outputs(9880) <= a and b;
    layer1_outputs(9881) <= not (a xor b);
    layer1_outputs(9882) <= b and not a;
    layer1_outputs(9883) <= not b or a;
    layer1_outputs(9884) <= b;
    layer1_outputs(9885) <= not b or a;
    layer1_outputs(9886) <= a;
    layer1_outputs(9887) <= a;
    layer1_outputs(9888) <= not a;
    layer1_outputs(9889) <= b;
    layer1_outputs(9890) <= b;
    layer1_outputs(9891) <= not (a and b);
    layer1_outputs(9892) <= not a or b;
    layer1_outputs(9893) <= a;
    layer1_outputs(9894) <= not (a or b);
    layer1_outputs(9895) <= a xor b;
    layer1_outputs(9896) <= not (a xor b);
    layer1_outputs(9897) <= a;
    layer1_outputs(9898) <= not (a and b);
    layer1_outputs(9899) <= not b;
    layer1_outputs(9900) <= not a;
    layer1_outputs(9901) <= not b or a;
    layer1_outputs(9902) <= a and not b;
    layer1_outputs(9903) <= not (a and b);
    layer1_outputs(9904) <= a or b;
    layer1_outputs(9905) <= a xor b;
    layer1_outputs(9906) <= b and not a;
    layer1_outputs(9907) <= not b;
    layer1_outputs(9908) <= b and not a;
    layer1_outputs(9909) <= b;
    layer1_outputs(9910) <= not a;
    layer1_outputs(9911) <= a xor b;
    layer1_outputs(9912) <= b;
    layer1_outputs(9913) <= not (a and b);
    layer1_outputs(9914) <= a or b;
    layer1_outputs(9915) <= not a;
    layer1_outputs(9916) <= not (a xor b);
    layer1_outputs(9917) <= a or b;
    layer1_outputs(9918) <= not b;
    layer1_outputs(9919) <= a or b;
    layer1_outputs(9920) <= not (a xor b);
    layer1_outputs(9921) <= not b or a;
    layer1_outputs(9922) <= a xor b;
    layer1_outputs(9923) <= not b;
    layer1_outputs(9924) <= a;
    layer1_outputs(9925) <= not (a or b);
    layer1_outputs(9926) <= b and not a;
    layer1_outputs(9927) <= a xor b;
    layer1_outputs(9928) <= a xor b;
    layer1_outputs(9929) <= b;
    layer1_outputs(9930) <= not (a or b);
    layer1_outputs(9931) <= not b;
    layer1_outputs(9932) <= not b or a;
    layer1_outputs(9933) <= a xor b;
    layer1_outputs(9934) <= not a;
    layer1_outputs(9935) <= a and not b;
    layer1_outputs(9936) <= 1'b1;
    layer1_outputs(9937) <= not a or b;
    layer1_outputs(9938) <= not b;
    layer1_outputs(9939) <= b;
    layer1_outputs(9940) <= not (a xor b);
    layer1_outputs(9941) <= not (a xor b);
    layer1_outputs(9942) <= a xor b;
    layer1_outputs(9943) <= a or b;
    layer1_outputs(9944) <= not b;
    layer1_outputs(9945) <= not (a xor b);
    layer1_outputs(9946) <= a;
    layer1_outputs(9947) <= a and not b;
    layer1_outputs(9948) <= 1'b0;
    layer1_outputs(9949) <= not b or a;
    layer1_outputs(9950) <= b;
    layer1_outputs(9951) <= not b or a;
    layer1_outputs(9952) <= a xor b;
    layer1_outputs(9953) <= not a or b;
    layer1_outputs(9954) <= b and not a;
    layer1_outputs(9955) <= a and b;
    layer1_outputs(9956) <= a and b;
    layer1_outputs(9957) <= not b;
    layer1_outputs(9958) <= not (a or b);
    layer1_outputs(9959) <= not b;
    layer1_outputs(9960) <= a;
    layer1_outputs(9961) <= a xor b;
    layer1_outputs(9962) <= not (a xor b);
    layer1_outputs(9963) <= not a;
    layer1_outputs(9964) <= a or b;
    layer1_outputs(9965) <= a and b;
    layer1_outputs(9966) <= a xor b;
    layer1_outputs(9967) <= not b;
    layer1_outputs(9968) <= a xor b;
    layer1_outputs(9969) <= a xor b;
    layer1_outputs(9970) <= b;
    layer1_outputs(9971) <= not b;
    layer1_outputs(9972) <= not b or a;
    layer1_outputs(9973) <= b;
    layer1_outputs(9974) <= not a or b;
    layer1_outputs(9975) <= a xor b;
    layer1_outputs(9976) <= a or b;
    layer1_outputs(9977) <= 1'b1;
    layer1_outputs(9978) <= b;
    layer1_outputs(9979) <= a and b;
    layer1_outputs(9980) <= not b or a;
    layer1_outputs(9981) <= not (a and b);
    layer1_outputs(9982) <= a or b;
    layer1_outputs(9983) <= not a;
    layer1_outputs(9984) <= not a;
    layer1_outputs(9985) <= not (a or b);
    layer1_outputs(9986) <= not (a and b);
    layer1_outputs(9987) <= not (a or b);
    layer1_outputs(9988) <= a xor b;
    layer1_outputs(9989) <= not a;
    layer1_outputs(9990) <= b;
    layer1_outputs(9991) <= a or b;
    layer1_outputs(9992) <= not a;
    layer1_outputs(9993) <= not b;
    layer1_outputs(9994) <= not a;
    layer1_outputs(9995) <= b and not a;
    layer1_outputs(9996) <= a or b;
    layer1_outputs(9997) <= b and not a;
    layer1_outputs(9998) <= not a or b;
    layer1_outputs(9999) <= a;
    layer1_outputs(10000) <= not b;
    layer1_outputs(10001) <= a and not b;
    layer1_outputs(10002) <= not b;
    layer1_outputs(10003) <= b and not a;
    layer1_outputs(10004) <= b;
    layer1_outputs(10005) <= a and b;
    layer1_outputs(10006) <= a or b;
    layer1_outputs(10007) <= a xor b;
    layer1_outputs(10008) <= not (a xor b);
    layer1_outputs(10009) <= a and b;
    layer1_outputs(10010) <= a xor b;
    layer1_outputs(10011) <= a and not b;
    layer1_outputs(10012) <= not b or a;
    layer1_outputs(10013) <= not (a and b);
    layer1_outputs(10014) <= b;
    layer1_outputs(10015) <= not a;
    layer1_outputs(10016) <= 1'b0;
    layer1_outputs(10017) <= not b or a;
    layer1_outputs(10018) <= b and not a;
    layer1_outputs(10019) <= not (a and b);
    layer1_outputs(10020) <= not (a xor b);
    layer1_outputs(10021) <= a xor b;
    layer1_outputs(10022) <= a;
    layer1_outputs(10023) <= a and b;
    layer1_outputs(10024) <= not b;
    layer1_outputs(10025) <= not (a or b);
    layer1_outputs(10026) <= a xor b;
    layer1_outputs(10027) <= b and not a;
    layer1_outputs(10028) <= b and not a;
    layer1_outputs(10029) <= not (a or b);
    layer1_outputs(10030) <= not (a xor b);
    layer1_outputs(10031) <= not a;
    layer1_outputs(10032) <= a and b;
    layer1_outputs(10033) <= not (a xor b);
    layer1_outputs(10034) <= not b or a;
    layer1_outputs(10035) <= b;
    layer1_outputs(10036) <= not b or a;
    layer1_outputs(10037) <= not (a xor b);
    layer1_outputs(10038) <= a xor b;
    layer1_outputs(10039) <= a and not b;
    layer1_outputs(10040) <= b;
    layer1_outputs(10041) <= a xor b;
    layer1_outputs(10042) <= not (a xor b);
    layer1_outputs(10043) <= b;
    layer1_outputs(10044) <= not a;
    layer1_outputs(10045) <= a and not b;
    layer1_outputs(10046) <= a;
    layer1_outputs(10047) <= not a or b;
    layer1_outputs(10048) <= not (a and b);
    layer1_outputs(10049) <= not (a and b);
    layer1_outputs(10050) <= not b;
    layer1_outputs(10051) <= not b;
    layer1_outputs(10052) <= not a or b;
    layer1_outputs(10053) <= not (a and b);
    layer1_outputs(10054) <= b;
    layer1_outputs(10055) <= b and not a;
    layer1_outputs(10056) <= a;
    layer1_outputs(10057) <= 1'b0;
    layer1_outputs(10058) <= not (a or b);
    layer1_outputs(10059) <= not a or b;
    layer1_outputs(10060) <= not b or a;
    layer1_outputs(10061) <= not b;
    layer1_outputs(10062) <= not (a or b);
    layer1_outputs(10063) <= a xor b;
    layer1_outputs(10064) <= a and b;
    layer1_outputs(10065) <= a;
    layer1_outputs(10066) <= not b;
    layer1_outputs(10067) <= not (a and b);
    layer1_outputs(10068) <= a xor b;
    layer1_outputs(10069) <= not b;
    layer1_outputs(10070) <= not a;
    layer1_outputs(10071) <= a and not b;
    layer1_outputs(10072) <= a;
    layer1_outputs(10073) <= a and not b;
    layer1_outputs(10074) <= a and b;
    layer1_outputs(10075) <= not (a or b);
    layer1_outputs(10076) <= not b or a;
    layer1_outputs(10077) <= a;
    layer1_outputs(10078) <= a and b;
    layer1_outputs(10079) <= not a;
    layer1_outputs(10080) <= not a or b;
    layer1_outputs(10081) <= not a;
    layer1_outputs(10082) <= not b;
    layer1_outputs(10083) <= not (a or b);
    layer1_outputs(10084) <= not (a xor b);
    layer1_outputs(10085) <= a;
    layer1_outputs(10086) <= a;
    layer1_outputs(10087) <= a and not b;
    layer1_outputs(10088) <= not b;
    layer1_outputs(10089) <= not (a or b);
    layer1_outputs(10090) <= not (a xor b);
    layer1_outputs(10091) <= not a;
    layer1_outputs(10092) <= a and not b;
    layer1_outputs(10093) <= not a or b;
    layer1_outputs(10094) <= not a;
    layer1_outputs(10095) <= b;
    layer1_outputs(10096) <= a or b;
    layer1_outputs(10097) <= not b;
    layer1_outputs(10098) <= not b or a;
    layer1_outputs(10099) <= not a;
    layer1_outputs(10100) <= a and not b;
    layer1_outputs(10101) <= not (a or b);
    layer1_outputs(10102) <= not b or a;
    layer1_outputs(10103) <= not b;
    layer1_outputs(10104) <= b;
    layer1_outputs(10105) <= not a;
    layer1_outputs(10106) <= not (a and b);
    layer1_outputs(10107) <= a;
    layer1_outputs(10108) <= not b;
    layer1_outputs(10109) <= b and not a;
    layer1_outputs(10110) <= not (a and b);
    layer1_outputs(10111) <= not b;
    layer1_outputs(10112) <= not a;
    layer1_outputs(10113) <= not a;
    layer1_outputs(10114) <= not b;
    layer1_outputs(10115) <= not a or b;
    layer1_outputs(10116) <= not b or a;
    layer1_outputs(10117) <= not (a and b);
    layer1_outputs(10118) <= 1'b1;
    layer1_outputs(10119) <= a;
    layer1_outputs(10120) <= b;
    layer1_outputs(10121) <= not b;
    layer1_outputs(10122) <= a;
    layer1_outputs(10123) <= b and not a;
    layer1_outputs(10124) <= not b;
    layer1_outputs(10125) <= 1'b0;
    layer1_outputs(10126) <= not b;
    layer1_outputs(10127) <= not (a xor b);
    layer1_outputs(10128) <= not (a xor b);
    layer1_outputs(10129) <= a xor b;
    layer1_outputs(10130) <= not a;
    layer1_outputs(10131) <= a and b;
    layer1_outputs(10132) <= b;
    layer1_outputs(10133) <= a;
    layer1_outputs(10134) <= a;
    layer1_outputs(10135) <= a;
    layer1_outputs(10136) <= a or b;
    layer1_outputs(10137) <= a and not b;
    layer1_outputs(10138) <= 1'b1;
    layer1_outputs(10139) <= a and not b;
    layer1_outputs(10140) <= not b;
    layer1_outputs(10141) <= not a or b;
    layer1_outputs(10142) <= not (a or b);
    layer1_outputs(10143) <= not b or a;
    layer1_outputs(10144) <= not b;
    layer1_outputs(10145) <= a;
    layer1_outputs(10146) <= a or b;
    layer1_outputs(10147) <= not (a and b);
    layer1_outputs(10148) <= not b;
    layer1_outputs(10149) <= not b or a;
    layer1_outputs(10150) <= 1'b0;
    layer1_outputs(10151) <= b;
    layer1_outputs(10152) <= a;
    layer1_outputs(10153) <= not a or b;
    layer1_outputs(10154) <= a;
    layer1_outputs(10155) <= a xor b;
    layer1_outputs(10156) <= not b;
    layer1_outputs(10157) <= a xor b;
    layer1_outputs(10158) <= not b or a;
    layer1_outputs(10159) <= a and not b;
    layer1_outputs(10160) <= a xor b;
    layer1_outputs(10161) <= not (a or b);
    layer1_outputs(10162) <= b;
    layer1_outputs(10163) <= not (a xor b);
    layer1_outputs(10164) <= not a;
    layer1_outputs(10165) <= not (a xor b);
    layer1_outputs(10166) <= a xor b;
    layer1_outputs(10167) <= a and b;
    layer1_outputs(10168) <= not (a xor b);
    layer1_outputs(10169) <= not a;
    layer1_outputs(10170) <= b and not a;
    layer1_outputs(10171) <= b and not a;
    layer1_outputs(10172) <= a;
    layer1_outputs(10173) <= a and b;
    layer1_outputs(10174) <= a xor b;
    layer1_outputs(10175) <= a;
    layer1_outputs(10176) <= not (a and b);
    layer1_outputs(10177) <= not (a and b);
    layer1_outputs(10178) <= not (a and b);
    layer1_outputs(10179) <= b;
    layer1_outputs(10180) <= not b;
    layer1_outputs(10181) <= a;
    layer1_outputs(10182) <= a or b;
    layer1_outputs(10183) <= not a;
    layer1_outputs(10184) <= not (a or b);
    layer1_outputs(10185) <= not (a xor b);
    layer1_outputs(10186) <= 1'b1;
    layer1_outputs(10187) <= b;
    layer1_outputs(10188) <= b;
    layer1_outputs(10189) <= not b or a;
    layer1_outputs(10190) <= a and not b;
    layer1_outputs(10191) <= not (a and b);
    layer1_outputs(10192) <= b and not a;
    layer1_outputs(10193) <= not b;
    layer1_outputs(10194) <= not a or b;
    layer1_outputs(10195) <= not a;
    layer1_outputs(10196) <= b;
    layer1_outputs(10197) <= not a or b;
    layer1_outputs(10198) <= b;
    layer1_outputs(10199) <= a or b;
    layer1_outputs(10200) <= a xor b;
    layer1_outputs(10201) <= b;
    layer1_outputs(10202) <= a;
    layer1_outputs(10203) <= a;
    layer1_outputs(10204) <= a or b;
    layer1_outputs(10205) <= b;
    layer1_outputs(10206) <= b and not a;
    layer1_outputs(10207) <= a and b;
    layer1_outputs(10208) <= a and not b;
    layer1_outputs(10209) <= b and not a;
    layer1_outputs(10210) <= not a or b;
    layer1_outputs(10211) <= a;
    layer1_outputs(10212) <= b;
    layer1_outputs(10213) <= a and not b;
    layer1_outputs(10214) <= not b;
    layer1_outputs(10215) <= not a;
    layer1_outputs(10216) <= not (a and b);
    layer1_outputs(10217) <= a;
    layer1_outputs(10218) <= not a or b;
    layer1_outputs(10219) <= not (a or b);
    layer1_outputs(10220) <= a or b;
    layer1_outputs(10221) <= not (a and b);
    layer1_outputs(10222) <= a or b;
    layer1_outputs(10223) <= b;
    layer1_outputs(10224) <= not a;
    layer1_outputs(10225) <= not (a or b);
    layer1_outputs(10226) <= not (a xor b);
    layer1_outputs(10227) <= a;
    layer1_outputs(10228) <= not a or b;
    layer1_outputs(10229) <= a;
    layer1_outputs(10230) <= a or b;
    layer1_outputs(10231) <= not (a xor b);
    layer1_outputs(10232) <= b;
    layer1_outputs(10233) <= not (a and b);
    layer1_outputs(10234) <= a or b;
    layer1_outputs(10235) <= not a;
    layer1_outputs(10236) <= not (a xor b);
    layer1_outputs(10237) <= not b or a;
    layer1_outputs(10238) <= not (a xor b);
    layer1_outputs(10239) <= a or b;
    layer1_outputs(10240) <= a and b;
    layer1_outputs(10241) <= not (a xor b);
    layer1_outputs(10242) <= not b or a;
    layer1_outputs(10243) <= not b or a;
    layer1_outputs(10244) <= not (a xor b);
    layer1_outputs(10245) <= a and b;
    layer1_outputs(10246) <= a or b;
    layer1_outputs(10247) <= not b;
    layer1_outputs(10248) <= a and b;
    layer1_outputs(10249) <= b and not a;
    layer1_outputs(10250) <= a and b;
    layer1_outputs(10251) <= a xor b;
    layer1_outputs(10252) <= not a or b;
    layer1_outputs(10253) <= not (a and b);
    layer1_outputs(10254) <= not (a and b);
    layer1_outputs(10255) <= not a;
    layer1_outputs(10256) <= a or b;
    layer1_outputs(10257) <= b;
    layer1_outputs(10258) <= not a or b;
    layer1_outputs(10259) <= not b;
    layer1_outputs(10260) <= 1'b1;
    layer1_outputs(10261) <= not b;
    layer1_outputs(10262) <= not a or b;
    layer1_outputs(10263) <= a;
    layer1_outputs(10264) <= a;
    layer1_outputs(10265) <= b and not a;
    layer1_outputs(10266) <= a;
    layer1_outputs(10267) <= a;
    layer1_outputs(10268) <= a;
    layer1_outputs(10269) <= a and not b;
    layer1_outputs(10270) <= b;
    layer1_outputs(10271) <= not (a or b);
    layer1_outputs(10272) <= a or b;
    layer1_outputs(10273) <= not a;
    layer1_outputs(10274) <= not a;
    layer1_outputs(10275) <= a and b;
    layer1_outputs(10276) <= not b or a;
    layer1_outputs(10277) <= not b;
    layer1_outputs(10278) <= not (a or b);
    layer1_outputs(10279) <= a and b;
    layer1_outputs(10280) <= not a;
    layer1_outputs(10281) <= not b;
    layer1_outputs(10282) <= b and not a;
    layer1_outputs(10283) <= a and not b;
    layer1_outputs(10284) <= a;
    layer1_outputs(10285) <= a or b;
    layer1_outputs(10286) <= a or b;
    layer1_outputs(10287) <= not b;
    layer1_outputs(10288) <= not a or b;
    layer1_outputs(10289) <= a xor b;
    layer1_outputs(10290) <= not a;
    layer1_outputs(10291) <= not (a and b);
    layer1_outputs(10292) <= not b;
    layer1_outputs(10293) <= b;
    layer1_outputs(10294) <= not (a xor b);
    layer1_outputs(10295) <= not b;
    layer1_outputs(10296) <= not b or a;
    layer1_outputs(10297) <= a xor b;
    layer1_outputs(10298) <= not a;
    layer1_outputs(10299) <= not (a and b);
    layer1_outputs(10300) <= b;
    layer1_outputs(10301) <= not a;
    layer1_outputs(10302) <= a or b;
    layer1_outputs(10303) <= b;
    layer1_outputs(10304) <= a xor b;
    layer1_outputs(10305) <= not a or b;
    layer1_outputs(10306) <= not b;
    layer1_outputs(10307) <= not a;
    layer1_outputs(10308) <= not b;
    layer1_outputs(10309) <= a and not b;
    layer1_outputs(10310) <= a and b;
    layer1_outputs(10311) <= a and not b;
    layer1_outputs(10312) <= not b;
    layer1_outputs(10313) <= not a or b;
    layer1_outputs(10314) <= not (a xor b);
    layer1_outputs(10315) <= a;
    layer1_outputs(10316) <= not (a and b);
    layer1_outputs(10317) <= not (a xor b);
    layer1_outputs(10318) <= not (a or b);
    layer1_outputs(10319) <= a xor b;
    layer1_outputs(10320) <= a;
    layer1_outputs(10321) <= b;
    layer1_outputs(10322) <= a xor b;
    layer1_outputs(10323) <= a;
    layer1_outputs(10324) <= not b;
    layer1_outputs(10325) <= not b or a;
    layer1_outputs(10326) <= not a;
    layer1_outputs(10327) <= not b or a;
    layer1_outputs(10328) <= not b or a;
    layer1_outputs(10329) <= not (a xor b);
    layer1_outputs(10330) <= a or b;
    layer1_outputs(10331) <= not a;
    layer1_outputs(10332) <= a xor b;
    layer1_outputs(10333) <= not a;
    layer1_outputs(10334) <= b;
    layer1_outputs(10335) <= not (a or b);
    layer1_outputs(10336) <= not (a xor b);
    layer1_outputs(10337) <= not (a xor b);
    layer1_outputs(10338) <= not a;
    layer1_outputs(10339) <= not b;
    layer1_outputs(10340) <= not (a and b);
    layer1_outputs(10341) <= not (a or b);
    layer1_outputs(10342) <= a;
    layer1_outputs(10343) <= not (a xor b);
    layer1_outputs(10344) <= not b;
    layer1_outputs(10345) <= not b;
    layer1_outputs(10346) <= a xor b;
    layer1_outputs(10347) <= not (a or b);
    layer1_outputs(10348) <= a and not b;
    layer1_outputs(10349) <= b and not a;
    layer1_outputs(10350) <= b;
    layer1_outputs(10351) <= a and b;
    layer1_outputs(10352) <= not (a xor b);
    layer1_outputs(10353) <= not a or b;
    layer1_outputs(10354) <= not a or b;
    layer1_outputs(10355) <= not (a and b);
    layer1_outputs(10356) <= not (a or b);
    layer1_outputs(10357) <= not a or b;
    layer1_outputs(10358) <= a and not b;
    layer1_outputs(10359) <= a;
    layer1_outputs(10360) <= not b or a;
    layer1_outputs(10361) <= not a or b;
    layer1_outputs(10362) <= 1'b1;
    layer1_outputs(10363) <= not (a xor b);
    layer1_outputs(10364) <= not (a xor b);
    layer1_outputs(10365) <= not b or a;
    layer1_outputs(10366) <= not (a or b);
    layer1_outputs(10367) <= a xor b;
    layer1_outputs(10368) <= a or b;
    layer1_outputs(10369) <= not (a xor b);
    layer1_outputs(10370) <= a;
    layer1_outputs(10371) <= not (a xor b);
    layer1_outputs(10372) <= a and not b;
    layer1_outputs(10373) <= not a or b;
    layer1_outputs(10374) <= 1'b1;
    layer1_outputs(10375) <= not (a xor b);
    layer1_outputs(10376) <= not a;
    layer1_outputs(10377) <= a or b;
    layer1_outputs(10378) <= a xor b;
    layer1_outputs(10379) <= not (a or b);
    layer1_outputs(10380) <= not (a and b);
    layer1_outputs(10381) <= a and not b;
    layer1_outputs(10382) <= not a;
    layer1_outputs(10383) <= a xor b;
    layer1_outputs(10384) <= b;
    layer1_outputs(10385) <= not b or a;
    layer1_outputs(10386) <= a and not b;
    layer1_outputs(10387) <= not (a or b);
    layer1_outputs(10388) <= a;
    layer1_outputs(10389) <= a or b;
    layer1_outputs(10390) <= b and not a;
    layer1_outputs(10391) <= not (a xor b);
    layer1_outputs(10392) <= b;
    layer1_outputs(10393) <= not (a and b);
    layer1_outputs(10394) <= not (a or b);
    layer1_outputs(10395) <= not a;
    layer1_outputs(10396) <= not a or b;
    layer1_outputs(10397) <= not (a xor b);
    layer1_outputs(10398) <= a and not b;
    layer1_outputs(10399) <= a or b;
    layer1_outputs(10400) <= b and not a;
    layer1_outputs(10401) <= a and not b;
    layer1_outputs(10402) <= a or b;
    layer1_outputs(10403) <= not (a or b);
    layer1_outputs(10404) <= not b;
    layer1_outputs(10405) <= b and not a;
    layer1_outputs(10406) <= not a or b;
    layer1_outputs(10407) <= not (a and b);
    layer1_outputs(10408) <= b;
    layer1_outputs(10409) <= not (a and b);
    layer1_outputs(10410) <= a and not b;
    layer1_outputs(10411) <= a and b;
    layer1_outputs(10412) <= a and not b;
    layer1_outputs(10413) <= b and not a;
    layer1_outputs(10414) <= a or b;
    layer1_outputs(10415) <= a and not b;
    layer1_outputs(10416) <= a and b;
    layer1_outputs(10417) <= a;
    layer1_outputs(10418) <= not b;
    layer1_outputs(10419) <= a;
    layer1_outputs(10420) <= not (a and b);
    layer1_outputs(10421) <= not a;
    layer1_outputs(10422) <= b and not a;
    layer1_outputs(10423) <= not (a or b);
    layer1_outputs(10424) <= b;
    layer1_outputs(10425) <= not (a or b);
    layer1_outputs(10426) <= not b;
    layer1_outputs(10427) <= a;
    layer1_outputs(10428) <= not (a xor b);
    layer1_outputs(10429) <= not a;
    layer1_outputs(10430) <= 1'b1;
    layer1_outputs(10431) <= not (a or b);
    layer1_outputs(10432) <= not a;
    layer1_outputs(10433) <= not (a and b);
    layer1_outputs(10434) <= a or b;
    layer1_outputs(10435) <= not (a and b);
    layer1_outputs(10436) <= not (a or b);
    layer1_outputs(10437) <= a;
    layer1_outputs(10438) <= 1'b0;
    layer1_outputs(10439) <= b;
    layer1_outputs(10440) <= a xor b;
    layer1_outputs(10441) <= a or b;
    layer1_outputs(10442) <= not (a or b);
    layer1_outputs(10443) <= b;
    layer1_outputs(10444) <= not a or b;
    layer1_outputs(10445) <= a or b;
    layer1_outputs(10446) <= not b or a;
    layer1_outputs(10447) <= a and not b;
    layer1_outputs(10448) <= b;
    layer1_outputs(10449) <= not b or a;
    layer1_outputs(10450) <= a or b;
    layer1_outputs(10451) <= a xor b;
    layer1_outputs(10452) <= not a;
    layer1_outputs(10453) <= 1'b1;
    layer1_outputs(10454) <= not a or b;
    layer1_outputs(10455) <= not a;
    layer1_outputs(10456) <= b;
    layer1_outputs(10457) <= not a;
    layer1_outputs(10458) <= a xor b;
    layer1_outputs(10459) <= a and b;
    layer1_outputs(10460) <= not a or b;
    layer1_outputs(10461) <= not b or a;
    layer1_outputs(10462) <= not b or a;
    layer1_outputs(10463) <= not b;
    layer1_outputs(10464) <= a and b;
    layer1_outputs(10465) <= not b;
    layer1_outputs(10466) <= not (a or b);
    layer1_outputs(10467) <= a and not b;
    layer1_outputs(10468) <= b;
    layer1_outputs(10469) <= not b or a;
    layer1_outputs(10470) <= a and not b;
    layer1_outputs(10471) <= not (a xor b);
    layer1_outputs(10472) <= a and b;
    layer1_outputs(10473) <= a xor b;
    layer1_outputs(10474) <= a xor b;
    layer1_outputs(10475) <= not a or b;
    layer1_outputs(10476) <= not b;
    layer1_outputs(10477) <= not a;
    layer1_outputs(10478) <= b and not a;
    layer1_outputs(10479) <= a xor b;
    layer1_outputs(10480) <= not a;
    layer1_outputs(10481) <= a xor b;
    layer1_outputs(10482) <= b and not a;
    layer1_outputs(10483) <= not (a or b);
    layer1_outputs(10484) <= a xor b;
    layer1_outputs(10485) <= a xor b;
    layer1_outputs(10486) <= a or b;
    layer1_outputs(10487) <= not b;
    layer1_outputs(10488) <= a or b;
    layer1_outputs(10489) <= not a;
    layer1_outputs(10490) <= not a or b;
    layer1_outputs(10491) <= not a;
    layer1_outputs(10492) <= a or b;
    layer1_outputs(10493) <= not a;
    layer1_outputs(10494) <= a xor b;
    layer1_outputs(10495) <= 1'b1;
    layer1_outputs(10496) <= not (a or b);
    layer1_outputs(10497) <= b;
    layer1_outputs(10498) <= a or b;
    layer1_outputs(10499) <= b;
    layer1_outputs(10500) <= b and not a;
    layer1_outputs(10501) <= a;
    layer1_outputs(10502) <= b and not a;
    layer1_outputs(10503) <= not b or a;
    layer1_outputs(10504) <= not a or b;
    layer1_outputs(10505) <= a or b;
    layer1_outputs(10506) <= a and not b;
    layer1_outputs(10507) <= a or b;
    layer1_outputs(10508) <= not a or b;
    layer1_outputs(10509) <= a and b;
    layer1_outputs(10510) <= b;
    layer1_outputs(10511) <= not (a xor b);
    layer1_outputs(10512) <= not a;
    layer1_outputs(10513) <= not b;
    layer1_outputs(10514) <= a xor b;
    layer1_outputs(10515) <= not (a xor b);
    layer1_outputs(10516) <= not a;
    layer1_outputs(10517) <= a and not b;
    layer1_outputs(10518) <= b;
    layer1_outputs(10519) <= a;
    layer1_outputs(10520) <= not a;
    layer1_outputs(10521) <= a xor b;
    layer1_outputs(10522) <= not a or b;
    layer1_outputs(10523) <= not (a xor b);
    layer1_outputs(10524) <= a xor b;
    layer1_outputs(10525) <= not (a and b);
    layer1_outputs(10526) <= not a or b;
    layer1_outputs(10527) <= not b or a;
    layer1_outputs(10528) <= b and not a;
    layer1_outputs(10529) <= b;
    layer1_outputs(10530) <= not a;
    layer1_outputs(10531) <= b;
    layer1_outputs(10532) <= b;
    layer1_outputs(10533) <= not a;
    layer1_outputs(10534) <= a;
    layer1_outputs(10535) <= not (a xor b);
    layer1_outputs(10536) <= not a;
    layer1_outputs(10537) <= not b;
    layer1_outputs(10538) <= not b;
    layer1_outputs(10539) <= a and not b;
    layer1_outputs(10540) <= not a;
    layer1_outputs(10541) <= not (a xor b);
    layer1_outputs(10542) <= a and not b;
    layer1_outputs(10543) <= not b or a;
    layer1_outputs(10544) <= not (a or b);
    layer1_outputs(10545) <= not a;
    layer1_outputs(10546) <= a;
    layer1_outputs(10547) <= b;
    layer1_outputs(10548) <= not b;
    layer1_outputs(10549) <= not (a or b);
    layer1_outputs(10550) <= a;
    layer1_outputs(10551) <= a or b;
    layer1_outputs(10552) <= not b or a;
    layer1_outputs(10553) <= not (a and b);
    layer1_outputs(10554) <= a and not b;
    layer1_outputs(10555) <= 1'b1;
    layer1_outputs(10556) <= a or b;
    layer1_outputs(10557) <= not a;
    layer1_outputs(10558) <= not (a xor b);
    layer1_outputs(10559) <= not b;
    layer1_outputs(10560) <= b;
    layer1_outputs(10561) <= not a or b;
    layer1_outputs(10562) <= a xor b;
    layer1_outputs(10563) <= not a;
    layer1_outputs(10564) <= not (a or b);
    layer1_outputs(10565) <= a and b;
    layer1_outputs(10566) <= not b;
    layer1_outputs(10567) <= a or b;
    layer1_outputs(10568) <= a;
    layer1_outputs(10569) <= not b or a;
    layer1_outputs(10570) <= a;
    layer1_outputs(10571) <= a and b;
    layer1_outputs(10572) <= not (a or b);
    layer1_outputs(10573) <= a;
    layer1_outputs(10574) <= not b or a;
    layer1_outputs(10575) <= a and b;
    layer1_outputs(10576) <= b;
    layer1_outputs(10577) <= not (a xor b);
    layer1_outputs(10578) <= not a;
    layer1_outputs(10579) <= not a or b;
    layer1_outputs(10580) <= not b or a;
    layer1_outputs(10581) <= not b;
    layer1_outputs(10582) <= a xor b;
    layer1_outputs(10583) <= not (a and b);
    layer1_outputs(10584) <= a and not b;
    layer1_outputs(10585) <= a and not b;
    layer1_outputs(10586) <= a or b;
    layer1_outputs(10587) <= not b or a;
    layer1_outputs(10588) <= a xor b;
    layer1_outputs(10589) <= not (a and b);
    layer1_outputs(10590) <= not b;
    layer1_outputs(10591) <= b;
    layer1_outputs(10592) <= not (a xor b);
    layer1_outputs(10593) <= not (a xor b);
    layer1_outputs(10594) <= not a or b;
    layer1_outputs(10595) <= not b or a;
    layer1_outputs(10596) <= b;
    layer1_outputs(10597) <= not b or a;
    layer1_outputs(10598) <= b;
    layer1_outputs(10599) <= b;
    layer1_outputs(10600) <= a xor b;
    layer1_outputs(10601) <= not a;
    layer1_outputs(10602) <= a or b;
    layer1_outputs(10603) <= a and not b;
    layer1_outputs(10604) <= not a;
    layer1_outputs(10605) <= a and b;
    layer1_outputs(10606) <= not a or b;
    layer1_outputs(10607) <= not b;
    layer1_outputs(10608) <= a xor b;
    layer1_outputs(10609) <= not (a or b);
    layer1_outputs(10610) <= a and b;
    layer1_outputs(10611) <= not b or a;
    layer1_outputs(10612) <= a and b;
    layer1_outputs(10613) <= a and b;
    layer1_outputs(10614) <= not b;
    layer1_outputs(10615) <= a xor b;
    layer1_outputs(10616) <= a xor b;
    layer1_outputs(10617) <= a and not b;
    layer1_outputs(10618) <= b;
    layer1_outputs(10619) <= not (a or b);
    layer1_outputs(10620) <= not (a or b);
    layer1_outputs(10621) <= not a or b;
    layer1_outputs(10622) <= a xor b;
    layer1_outputs(10623) <= a;
    layer1_outputs(10624) <= not b;
    layer1_outputs(10625) <= a or b;
    layer1_outputs(10626) <= b;
    layer1_outputs(10627) <= a or b;
    layer1_outputs(10628) <= a and b;
    layer1_outputs(10629) <= not (a xor b);
    layer1_outputs(10630) <= not b;
    layer1_outputs(10631) <= not (a and b);
    layer1_outputs(10632) <= a and not b;
    layer1_outputs(10633) <= a or b;
    layer1_outputs(10634) <= 1'b1;
    layer1_outputs(10635) <= not (a xor b);
    layer1_outputs(10636) <= b and not a;
    layer1_outputs(10637) <= not (a xor b);
    layer1_outputs(10638) <= b and not a;
    layer1_outputs(10639) <= 1'b1;
    layer1_outputs(10640) <= not (a xor b);
    layer1_outputs(10641) <= not (a xor b);
    layer1_outputs(10642) <= not b;
    layer1_outputs(10643) <= a xor b;
    layer1_outputs(10644) <= b and not a;
    layer1_outputs(10645) <= not b;
    layer1_outputs(10646) <= a and not b;
    layer1_outputs(10647) <= b;
    layer1_outputs(10648) <= b;
    layer1_outputs(10649) <= not (a and b);
    layer1_outputs(10650) <= not (a or b);
    layer1_outputs(10651) <= not (a xor b);
    layer1_outputs(10652) <= a or b;
    layer1_outputs(10653) <= not b;
    layer1_outputs(10654) <= a or b;
    layer1_outputs(10655) <= not b or a;
    layer1_outputs(10656) <= not a;
    layer1_outputs(10657) <= not (a xor b);
    layer1_outputs(10658) <= 1'b1;
    layer1_outputs(10659) <= b;
    layer1_outputs(10660) <= not a;
    layer1_outputs(10661) <= not (a xor b);
    layer1_outputs(10662) <= not a;
    layer1_outputs(10663) <= not b or a;
    layer1_outputs(10664) <= not (a and b);
    layer1_outputs(10665) <= a or b;
    layer1_outputs(10666) <= a and b;
    layer1_outputs(10667) <= not b or a;
    layer1_outputs(10668) <= a or b;
    layer1_outputs(10669) <= not a or b;
    layer1_outputs(10670) <= a and b;
    layer1_outputs(10671) <= a;
    layer1_outputs(10672) <= a or b;
    layer1_outputs(10673) <= not b or a;
    layer1_outputs(10674) <= a;
    layer1_outputs(10675) <= not b;
    layer1_outputs(10676) <= not b;
    layer1_outputs(10677) <= not (a and b);
    layer1_outputs(10678) <= a and not b;
    layer1_outputs(10679) <= not a;
    layer1_outputs(10680) <= a;
    layer1_outputs(10681) <= a and not b;
    layer1_outputs(10682) <= not b;
    layer1_outputs(10683) <= a and b;
    layer1_outputs(10684) <= not b;
    layer1_outputs(10685) <= b and not a;
    layer1_outputs(10686) <= not (a or b);
    layer1_outputs(10687) <= not a or b;
    layer1_outputs(10688) <= a;
    layer1_outputs(10689) <= not a;
    layer1_outputs(10690) <= a xor b;
    layer1_outputs(10691) <= a and b;
    layer1_outputs(10692) <= a xor b;
    layer1_outputs(10693) <= not b;
    layer1_outputs(10694) <= b and not a;
    layer1_outputs(10695) <= not (a xor b);
    layer1_outputs(10696) <= b;
    layer1_outputs(10697) <= not (a or b);
    layer1_outputs(10698) <= not b or a;
    layer1_outputs(10699) <= not a;
    layer1_outputs(10700) <= not a or b;
    layer1_outputs(10701) <= not (a xor b);
    layer1_outputs(10702) <= a;
    layer1_outputs(10703) <= not a or b;
    layer1_outputs(10704) <= not a or b;
    layer1_outputs(10705) <= not a or b;
    layer1_outputs(10706) <= not (a and b);
    layer1_outputs(10707) <= not a;
    layer1_outputs(10708) <= b and not a;
    layer1_outputs(10709) <= b;
    layer1_outputs(10710) <= not b or a;
    layer1_outputs(10711) <= not (a or b);
    layer1_outputs(10712) <= b;
    layer1_outputs(10713) <= b;
    layer1_outputs(10714) <= a and b;
    layer1_outputs(10715) <= not (a or b);
    layer1_outputs(10716) <= not b;
    layer1_outputs(10717) <= a and not b;
    layer1_outputs(10718) <= not a;
    layer1_outputs(10719) <= b;
    layer1_outputs(10720) <= not b;
    layer1_outputs(10721) <= 1'b1;
    layer1_outputs(10722) <= not a;
    layer1_outputs(10723) <= not a or b;
    layer1_outputs(10724) <= a and b;
    layer1_outputs(10725) <= b;
    layer1_outputs(10726) <= a or b;
    layer1_outputs(10727) <= b and not a;
    layer1_outputs(10728) <= not (a xor b);
    layer1_outputs(10729) <= a xor b;
    layer1_outputs(10730) <= not b;
    layer1_outputs(10731) <= b and not a;
    layer1_outputs(10732) <= a xor b;
    layer1_outputs(10733) <= not (a or b);
    layer1_outputs(10734) <= not a or b;
    layer1_outputs(10735) <= not (a and b);
    layer1_outputs(10736) <= not (a xor b);
    layer1_outputs(10737) <= a or b;
    layer1_outputs(10738) <= a and b;
    layer1_outputs(10739) <= not b;
    layer1_outputs(10740) <= b;
    layer1_outputs(10741) <= not a;
    layer1_outputs(10742) <= not a or b;
    layer1_outputs(10743) <= a or b;
    layer1_outputs(10744) <= not b;
    layer1_outputs(10745) <= a and not b;
    layer1_outputs(10746) <= b and not a;
    layer1_outputs(10747) <= b;
    layer1_outputs(10748) <= 1'b0;
    layer1_outputs(10749) <= not b or a;
    layer1_outputs(10750) <= not (a and b);
    layer1_outputs(10751) <= a and not b;
    layer1_outputs(10752) <= not (a or b);
    layer1_outputs(10753) <= not b or a;
    layer1_outputs(10754) <= not b or a;
    layer1_outputs(10755) <= not (a xor b);
    layer1_outputs(10756) <= a;
    layer1_outputs(10757) <= a and b;
    layer1_outputs(10758) <= a and not b;
    layer1_outputs(10759) <= a and b;
    layer1_outputs(10760) <= not a or b;
    layer1_outputs(10761) <= a xor b;
    layer1_outputs(10762) <= not b;
    layer1_outputs(10763) <= not a;
    layer1_outputs(10764) <= not a or b;
    layer1_outputs(10765) <= a and b;
    layer1_outputs(10766) <= a and not b;
    layer1_outputs(10767) <= not (a or b);
    layer1_outputs(10768) <= not b or a;
    layer1_outputs(10769) <= not b or a;
    layer1_outputs(10770) <= a or b;
    layer1_outputs(10771) <= not (a and b);
    layer1_outputs(10772) <= not (a or b);
    layer1_outputs(10773) <= 1'b1;
    layer1_outputs(10774) <= b;
    layer1_outputs(10775) <= not b;
    layer1_outputs(10776) <= a;
    layer1_outputs(10777) <= a xor b;
    layer1_outputs(10778) <= not a;
    layer1_outputs(10779) <= not a;
    layer1_outputs(10780) <= not (a and b);
    layer1_outputs(10781) <= a and b;
    layer1_outputs(10782) <= a and b;
    layer1_outputs(10783) <= not a;
    layer1_outputs(10784) <= not a;
    layer1_outputs(10785) <= a xor b;
    layer1_outputs(10786) <= a or b;
    layer1_outputs(10787) <= not a;
    layer1_outputs(10788) <= not a;
    layer1_outputs(10789) <= b and not a;
    layer1_outputs(10790) <= a and b;
    layer1_outputs(10791) <= b;
    layer1_outputs(10792) <= a or b;
    layer1_outputs(10793) <= not (a xor b);
    layer1_outputs(10794) <= a and b;
    layer1_outputs(10795) <= a and b;
    layer1_outputs(10796) <= b;
    layer1_outputs(10797) <= not (a and b);
    layer1_outputs(10798) <= a xor b;
    layer1_outputs(10799) <= not (a and b);
    layer1_outputs(10800) <= a xor b;
    layer1_outputs(10801) <= a and not b;
    layer1_outputs(10802) <= a and b;
    layer1_outputs(10803) <= b;
    layer1_outputs(10804) <= a xor b;
    layer1_outputs(10805) <= not (a and b);
    layer1_outputs(10806) <= b;
    layer1_outputs(10807) <= not (a or b);
    layer1_outputs(10808) <= b and not a;
    layer1_outputs(10809) <= not (a or b);
    layer1_outputs(10810) <= b and not a;
    layer1_outputs(10811) <= not a or b;
    layer1_outputs(10812) <= b and not a;
    layer1_outputs(10813) <= not a;
    layer1_outputs(10814) <= a or b;
    layer1_outputs(10815) <= b and not a;
    layer1_outputs(10816) <= not (a and b);
    layer1_outputs(10817) <= not b or a;
    layer1_outputs(10818) <= not a;
    layer1_outputs(10819) <= not (a or b);
    layer1_outputs(10820) <= not (a and b);
    layer1_outputs(10821) <= 1'b0;
    layer1_outputs(10822) <= not (a xor b);
    layer1_outputs(10823) <= a and not b;
    layer1_outputs(10824) <= not (a or b);
    layer1_outputs(10825) <= b;
    layer1_outputs(10826) <= a;
    layer1_outputs(10827) <= b and not a;
    layer1_outputs(10828) <= a and not b;
    layer1_outputs(10829) <= b and not a;
    layer1_outputs(10830) <= a or b;
    layer1_outputs(10831) <= a xor b;
    layer1_outputs(10832) <= not (a or b);
    layer1_outputs(10833) <= b;
    layer1_outputs(10834) <= a or b;
    layer1_outputs(10835) <= not (a and b);
    layer1_outputs(10836) <= not a;
    layer1_outputs(10837) <= not a or b;
    layer1_outputs(10838) <= a and b;
    layer1_outputs(10839) <= b;
    layer1_outputs(10840) <= not a;
    layer1_outputs(10841) <= not b or a;
    layer1_outputs(10842) <= not a;
    layer1_outputs(10843) <= b;
    layer1_outputs(10844) <= a or b;
    layer1_outputs(10845) <= a and not b;
    layer1_outputs(10846) <= not a or b;
    layer1_outputs(10847) <= not a;
    layer1_outputs(10848) <= not a or b;
    layer1_outputs(10849) <= a or b;
    layer1_outputs(10850) <= not (a xor b);
    layer1_outputs(10851) <= a xor b;
    layer1_outputs(10852) <= not a;
    layer1_outputs(10853) <= b and not a;
    layer1_outputs(10854) <= not b or a;
    layer1_outputs(10855) <= a and b;
    layer1_outputs(10856) <= a and b;
    layer1_outputs(10857) <= a and not b;
    layer1_outputs(10858) <= not b;
    layer1_outputs(10859) <= b and not a;
    layer1_outputs(10860) <= not a or b;
    layer1_outputs(10861) <= a or b;
    layer1_outputs(10862) <= not a;
    layer1_outputs(10863) <= b and not a;
    layer1_outputs(10864) <= not b;
    layer1_outputs(10865) <= not (a xor b);
    layer1_outputs(10866) <= not b;
    layer1_outputs(10867) <= a or b;
    layer1_outputs(10868) <= a and b;
    layer1_outputs(10869) <= b;
    layer1_outputs(10870) <= a and b;
    layer1_outputs(10871) <= b;
    layer1_outputs(10872) <= not a;
    layer1_outputs(10873) <= not (a and b);
    layer1_outputs(10874) <= a and not b;
    layer1_outputs(10875) <= not (a and b);
    layer1_outputs(10876) <= not a;
    layer1_outputs(10877) <= a and not b;
    layer1_outputs(10878) <= b and not a;
    layer1_outputs(10879) <= not a or b;
    layer1_outputs(10880) <= not a or b;
    layer1_outputs(10881) <= b;
    layer1_outputs(10882) <= not b;
    layer1_outputs(10883) <= a;
    layer1_outputs(10884) <= not b or a;
    layer1_outputs(10885) <= not a;
    layer1_outputs(10886) <= b and not a;
    layer1_outputs(10887) <= a and b;
    layer1_outputs(10888) <= not a;
    layer1_outputs(10889) <= not a;
    layer1_outputs(10890) <= a;
    layer1_outputs(10891) <= a;
    layer1_outputs(10892) <= b;
    layer1_outputs(10893) <= a and not b;
    layer1_outputs(10894) <= not (a and b);
    layer1_outputs(10895) <= 1'b0;
    layer1_outputs(10896) <= not b;
    layer1_outputs(10897) <= a;
    layer1_outputs(10898) <= not (a and b);
    layer1_outputs(10899) <= not b or a;
    layer1_outputs(10900) <= not a;
    layer1_outputs(10901) <= not a or b;
    layer1_outputs(10902) <= not (a xor b);
    layer1_outputs(10903) <= not (a xor b);
    layer1_outputs(10904) <= a xor b;
    layer1_outputs(10905) <= not a;
    layer1_outputs(10906) <= not (a or b);
    layer1_outputs(10907) <= not b or a;
    layer1_outputs(10908) <= not a;
    layer1_outputs(10909) <= a xor b;
    layer1_outputs(10910) <= 1'b1;
    layer1_outputs(10911) <= not a;
    layer1_outputs(10912) <= not (a and b);
    layer1_outputs(10913) <= not a or b;
    layer1_outputs(10914) <= a;
    layer1_outputs(10915) <= not b or a;
    layer1_outputs(10916) <= not b;
    layer1_outputs(10917) <= b and not a;
    layer1_outputs(10918) <= not b;
    layer1_outputs(10919) <= a and b;
    layer1_outputs(10920) <= not (a xor b);
    layer1_outputs(10921) <= b;
    layer1_outputs(10922) <= 1'b1;
    layer1_outputs(10923) <= a;
    layer1_outputs(10924) <= not (a xor b);
    layer1_outputs(10925) <= not b or a;
    layer1_outputs(10926) <= a and not b;
    layer1_outputs(10927) <= not b;
    layer1_outputs(10928) <= a or b;
    layer1_outputs(10929) <= a;
    layer1_outputs(10930) <= a;
    layer1_outputs(10931) <= a xor b;
    layer1_outputs(10932) <= not (a and b);
    layer1_outputs(10933) <= not a or b;
    layer1_outputs(10934) <= not b or a;
    layer1_outputs(10935) <= not (a xor b);
    layer1_outputs(10936) <= 1'b0;
    layer1_outputs(10937) <= not b;
    layer1_outputs(10938) <= a or b;
    layer1_outputs(10939) <= not (a or b);
    layer1_outputs(10940) <= not (a and b);
    layer1_outputs(10941) <= a or b;
    layer1_outputs(10942) <= a;
    layer1_outputs(10943) <= not a;
    layer1_outputs(10944) <= b;
    layer1_outputs(10945) <= a or b;
    layer1_outputs(10946) <= not a or b;
    layer1_outputs(10947) <= not b or a;
    layer1_outputs(10948) <= not (a or b);
    layer1_outputs(10949) <= a and b;
    layer1_outputs(10950) <= not b;
    layer1_outputs(10951) <= a xor b;
    layer1_outputs(10952) <= a and b;
    layer1_outputs(10953) <= not (a and b);
    layer1_outputs(10954) <= 1'b0;
    layer1_outputs(10955) <= 1'b1;
    layer1_outputs(10956) <= not (a or b);
    layer1_outputs(10957) <= a or b;
    layer1_outputs(10958) <= a or b;
    layer1_outputs(10959) <= not a;
    layer1_outputs(10960) <= b;
    layer1_outputs(10961) <= not a;
    layer1_outputs(10962) <= not b;
    layer1_outputs(10963) <= not b or a;
    layer1_outputs(10964) <= b;
    layer1_outputs(10965) <= not b;
    layer1_outputs(10966) <= not (a xor b);
    layer1_outputs(10967) <= a xor b;
    layer1_outputs(10968) <= not a or b;
    layer1_outputs(10969) <= not (a or b);
    layer1_outputs(10970) <= not a;
    layer1_outputs(10971) <= b and not a;
    layer1_outputs(10972) <= a;
    layer1_outputs(10973) <= not (a or b);
    layer1_outputs(10974) <= a;
    layer1_outputs(10975) <= b and not a;
    layer1_outputs(10976) <= b and not a;
    layer1_outputs(10977) <= not a or b;
    layer1_outputs(10978) <= a xor b;
    layer1_outputs(10979) <= not b or a;
    layer1_outputs(10980) <= a or b;
    layer1_outputs(10981) <= not a or b;
    layer1_outputs(10982) <= a or b;
    layer1_outputs(10983) <= not (a xor b);
    layer1_outputs(10984) <= b and not a;
    layer1_outputs(10985) <= a or b;
    layer1_outputs(10986) <= a and b;
    layer1_outputs(10987) <= not (a and b);
    layer1_outputs(10988) <= a;
    layer1_outputs(10989) <= a xor b;
    layer1_outputs(10990) <= b;
    layer1_outputs(10991) <= not a or b;
    layer1_outputs(10992) <= not (a xor b);
    layer1_outputs(10993) <= not a;
    layer1_outputs(10994) <= b and not a;
    layer1_outputs(10995) <= not b;
    layer1_outputs(10996) <= a;
    layer1_outputs(10997) <= a;
    layer1_outputs(10998) <= a or b;
    layer1_outputs(10999) <= a and not b;
    layer1_outputs(11000) <= b and not a;
    layer1_outputs(11001) <= b and not a;
    layer1_outputs(11002) <= not b or a;
    layer1_outputs(11003) <= b;
    layer1_outputs(11004) <= not (a xor b);
    layer1_outputs(11005) <= a and not b;
    layer1_outputs(11006) <= a or b;
    layer1_outputs(11007) <= not b;
    layer1_outputs(11008) <= not b;
    layer1_outputs(11009) <= not a;
    layer1_outputs(11010) <= not (a xor b);
    layer1_outputs(11011) <= not a or b;
    layer1_outputs(11012) <= b;
    layer1_outputs(11013) <= not b;
    layer1_outputs(11014) <= not b;
    layer1_outputs(11015) <= 1'b1;
    layer1_outputs(11016) <= a and b;
    layer1_outputs(11017) <= a and b;
    layer1_outputs(11018) <= a;
    layer1_outputs(11019) <= not a or b;
    layer1_outputs(11020) <= a or b;
    layer1_outputs(11021) <= not (a and b);
    layer1_outputs(11022) <= a xor b;
    layer1_outputs(11023) <= not (a or b);
    layer1_outputs(11024) <= a and b;
    layer1_outputs(11025) <= not b or a;
    layer1_outputs(11026) <= not (a xor b);
    layer1_outputs(11027) <= b;
    layer1_outputs(11028) <= not b;
    layer1_outputs(11029) <= not (a xor b);
    layer1_outputs(11030) <= a and not b;
    layer1_outputs(11031) <= not b;
    layer1_outputs(11032) <= not a;
    layer1_outputs(11033) <= a or b;
    layer1_outputs(11034) <= not a or b;
    layer1_outputs(11035) <= a and b;
    layer1_outputs(11036) <= not (a xor b);
    layer1_outputs(11037) <= a xor b;
    layer1_outputs(11038) <= a and b;
    layer1_outputs(11039) <= b;
    layer1_outputs(11040) <= not a;
    layer1_outputs(11041) <= not (a and b);
    layer1_outputs(11042) <= not a;
    layer1_outputs(11043) <= a;
    layer1_outputs(11044) <= a and b;
    layer1_outputs(11045) <= not b;
    layer1_outputs(11046) <= not a or b;
    layer1_outputs(11047) <= b;
    layer1_outputs(11048) <= not (a and b);
    layer1_outputs(11049) <= a and b;
    layer1_outputs(11050) <= not b;
    layer1_outputs(11051) <= not (a and b);
    layer1_outputs(11052) <= b and not a;
    layer1_outputs(11053) <= not (a and b);
    layer1_outputs(11054) <= not (a xor b);
    layer1_outputs(11055) <= b and not a;
    layer1_outputs(11056) <= b;
    layer1_outputs(11057) <= not (a xor b);
    layer1_outputs(11058) <= b and not a;
    layer1_outputs(11059) <= not (a and b);
    layer1_outputs(11060) <= b and not a;
    layer1_outputs(11061) <= a or b;
    layer1_outputs(11062) <= not a or b;
    layer1_outputs(11063) <= b and not a;
    layer1_outputs(11064) <= not a;
    layer1_outputs(11065) <= not a;
    layer1_outputs(11066) <= 1'b0;
    layer1_outputs(11067) <= not (a and b);
    layer1_outputs(11068) <= a and not b;
    layer1_outputs(11069) <= a and not b;
    layer1_outputs(11070) <= not a;
    layer1_outputs(11071) <= not (a or b);
    layer1_outputs(11072) <= a;
    layer1_outputs(11073) <= b;
    layer1_outputs(11074) <= not a or b;
    layer1_outputs(11075) <= not b or a;
    layer1_outputs(11076) <= not (a xor b);
    layer1_outputs(11077) <= not b or a;
    layer1_outputs(11078) <= not a or b;
    layer1_outputs(11079) <= not (a or b);
    layer1_outputs(11080) <= 1'b1;
    layer1_outputs(11081) <= 1'b1;
    layer1_outputs(11082) <= b;
    layer1_outputs(11083) <= not (a and b);
    layer1_outputs(11084) <= b and not a;
    layer1_outputs(11085) <= a and b;
    layer1_outputs(11086) <= not a or b;
    layer1_outputs(11087) <= not a or b;
    layer1_outputs(11088) <= a and b;
    layer1_outputs(11089) <= a or b;
    layer1_outputs(11090) <= a and not b;
    layer1_outputs(11091) <= a xor b;
    layer1_outputs(11092) <= a;
    layer1_outputs(11093) <= a or b;
    layer1_outputs(11094) <= b and not a;
    layer1_outputs(11095) <= not a or b;
    layer1_outputs(11096) <= a;
    layer1_outputs(11097) <= not (a or b);
    layer1_outputs(11098) <= not b or a;
    layer1_outputs(11099) <= not a;
    layer1_outputs(11100) <= a;
    layer1_outputs(11101) <= a and b;
    layer1_outputs(11102) <= not b;
    layer1_outputs(11103) <= a;
    layer1_outputs(11104) <= not a or b;
    layer1_outputs(11105) <= not a or b;
    layer1_outputs(11106) <= a;
    layer1_outputs(11107) <= a or b;
    layer1_outputs(11108) <= b;
    layer1_outputs(11109) <= b and not a;
    layer1_outputs(11110) <= not a or b;
    layer1_outputs(11111) <= not (a and b);
    layer1_outputs(11112) <= not (a and b);
    layer1_outputs(11113) <= not a;
    layer1_outputs(11114) <= not (a or b);
    layer1_outputs(11115) <= not b;
    layer1_outputs(11116) <= a and b;
    layer1_outputs(11117) <= a xor b;
    layer1_outputs(11118) <= a or b;
    layer1_outputs(11119) <= not b or a;
    layer1_outputs(11120) <= not (a xor b);
    layer1_outputs(11121) <= a;
    layer1_outputs(11122) <= not a;
    layer1_outputs(11123) <= b;
    layer1_outputs(11124) <= b;
    layer1_outputs(11125) <= not b;
    layer1_outputs(11126) <= not (a or b);
    layer1_outputs(11127) <= a and b;
    layer1_outputs(11128) <= 1'b1;
    layer1_outputs(11129) <= b;
    layer1_outputs(11130) <= a;
    layer1_outputs(11131) <= not b or a;
    layer1_outputs(11132) <= a and not b;
    layer1_outputs(11133) <= not (a xor b);
    layer1_outputs(11134) <= not (a xor b);
    layer1_outputs(11135) <= a xor b;
    layer1_outputs(11136) <= a and not b;
    layer1_outputs(11137) <= not a;
    layer1_outputs(11138) <= not b or a;
    layer1_outputs(11139) <= a xor b;
    layer1_outputs(11140) <= not b or a;
    layer1_outputs(11141) <= not a;
    layer1_outputs(11142) <= a;
    layer1_outputs(11143) <= not (a xor b);
    layer1_outputs(11144) <= not b;
    layer1_outputs(11145) <= b;
    layer1_outputs(11146) <= b and not a;
    layer1_outputs(11147) <= not (a or b);
    layer1_outputs(11148) <= not a or b;
    layer1_outputs(11149) <= a or b;
    layer1_outputs(11150) <= not a or b;
    layer1_outputs(11151) <= a xor b;
    layer1_outputs(11152) <= not a or b;
    layer1_outputs(11153) <= a or b;
    layer1_outputs(11154) <= a xor b;
    layer1_outputs(11155) <= not (a xor b);
    layer1_outputs(11156) <= b;
    layer1_outputs(11157) <= 1'b0;
    layer1_outputs(11158) <= a xor b;
    layer1_outputs(11159) <= not (a and b);
    layer1_outputs(11160) <= a and not b;
    layer1_outputs(11161) <= a;
    layer1_outputs(11162) <= not b or a;
    layer1_outputs(11163) <= not (a or b);
    layer1_outputs(11164) <= not a;
    layer1_outputs(11165) <= not a;
    layer1_outputs(11166) <= a xor b;
    layer1_outputs(11167) <= 1'b1;
    layer1_outputs(11168) <= not b or a;
    layer1_outputs(11169) <= a;
    layer1_outputs(11170) <= not b;
    layer1_outputs(11171) <= not b;
    layer1_outputs(11172) <= not b;
    layer1_outputs(11173) <= not a;
    layer1_outputs(11174) <= b;
    layer1_outputs(11175) <= 1'b0;
    layer1_outputs(11176) <= a xor b;
    layer1_outputs(11177) <= a and not b;
    layer1_outputs(11178) <= not (a xor b);
    layer1_outputs(11179) <= a xor b;
    layer1_outputs(11180) <= a xor b;
    layer1_outputs(11181) <= b and not a;
    layer1_outputs(11182) <= a;
    layer1_outputs(11183) <= not (a or b);
    layer1_outputs(11184) <= a xor b;
    layer1_outputs(11185) <= a;
    layer1_outputs(11186) <= not a or b;
    layer1_outputs(11187) <= not (a xor b);
    layer1_outputs(11188) <= a and not b;
    layer1_outputs(11189) <= a or b;
    layer1_outputs(11190) <= b;
    layer1_outputs(11191) <= a and b;
    layer1_outputs(11192) <= not a;
    layer1_outputs(11193) <= a or b;
    layer1_outputs(11194) <= a xor b;
    layer1_outputs(11195) <= not a or b;
    layer1_outputs(11196) <= b and not a;
    layer1_outputs(11197) <= a and b;
    layer1_outputs(11198) <= not b;
    layer1_outputs(11199) <= not b;
    layer1_outputs(11200) <= 1'b0;
    layer1_outputs(11201) <= a xor b;
    layer1_outputs(11202) <= a;
    layer1_outputs(11203) <= a and not b;
    layer1_outputs(11204) <= not a;
    layer1_outputs(11205) <= not (a or b);
    layer1_outputs(11206) <= a or b;
    layer1_outputs(11207) <= a and not b;
    layer1_outputs(11208) <= not b or a;
    layer1_outputs(11209) <= not a or b;
    layer1_outputs(11210) <= a;
    layer1_outputs(11211) <= a;
    layer1_outputs(11212) <= a;
    layer1_outputs(11213) <= not b;
    layer1_outputs(11214) <= not b or a;
    layer1_outputs(11215) <= not (a or b);
    layer1_outputs(11216) <= 1'b1;
    layer1_outputs(11217) <= not a;
    layer1_outputs(11218) <= not (a xor b);
    layer1_outputs(11219) <= a or b;
    layer1_outputs(11220) <= not (a and b);
    layer1_outputs(11221) <= not (a or b);
    layer1_outputs(11222) <= not b;
    layer1_outputs(11223) <= not (a or b);
    layer1_outputs(11224) <= not b or a;
    layer1_outputs(11225) <= a xor b;
    layer1_outputs(11226) <= not (a or b);
    layer1_outputs(11227) <= not (a or b);
    layer1_outputs(11228) <= not a;
    layer1_outputs(11229) <= not a;
    layer1_outputs(11230) <= a xor b;
    layer1_outputs(11231) <= a;
    layer1_outputs(11232) <= b and not a;
    layer1_outputs(11233) <= a or b;
    layer1_outputs(11234) <= not b;
    layer1_outputs(11235) <= not a or b;
    layer1_outputs(11236) <= a or b;
    layer1_outputs(11237) <= a or b;
    layer1_outputs(11238) <= not (a xor b);
    layer1_outputs(11239) <= b;
    layer1_outputs(11240) <= not a;
    layer1_outputs(11241) <= not (a and b);
    layer1_outputs(11242) <= not a;
    layer1_outputs(11243) <= a or b;
    layer1_outputs(11244) <= not a;
    layer1_outputs(11245) <= not b;
    layer1_outputs(11246) <= not (a and b);
    layer1_outputs(11247) <= a xor b;
    layer1_outputs(11248) <= a or b;
    layer1_outputs(11249) <= not a;
    layer1_outputs(11250) <= not a;
    layer1_outputs(11251) <= not (a and b);
    layer1_outputs(11252) <= a or b;
    layer1_outputs(11253) <= not (a or b);
    layer1_outputs(11254) <= a or b;
    layer1_outputs(11255) <= not (a xor b);
    layer1_outputs(11256) <= b;
    layer1_outputs(11257) <= not (a xor b);
    layer1_outputs(11258) <= not (a xor b);
    layer1_outputs(11259) <= a or b;
    layer1_outputs(11260) <= b and not a;
    layer1_outputs(11261) <= a;
    layer1_outputs(11262) <= not a;
    layer1_outputs(11263) <= not a or b;
    layer1_outputs(11264) <= not (a or b);
    layer1_outputs(11265) <= a and not b;
    layer1_outputs(11266) <= not a or b;
    layer1_outputs(11267) <= not (a and b);
    layer1_outputs(11268) <= a or b;
    layer1_outputs(11269) <= not a;
    layer1_outputs(11270) <= a;
    layer1_outputs(11271) <= not (a and b);
    layer1_outputs(11272) <= not b;
    layer1_outputs(11273) <= a xor b;
    layer1_outputs(11274) <= not (a or b);
    layer1_outputs(11275) <= not b;
    layer1_outputs(11276) <= 1'b0;
    layer1_outputs(11277) <= a and b;
    layer1_outputs(11278) <= not a or b;
    layer1_outputs(11279) <= a or b;
    layer1_outputs(11280) <= b and not a;
    layer1_outputs(11281) <= not a or b;
    layer1_outputs(11282) <= not a;
    layer1_outputs(11283) <= not (a and b);
    layer1_outputs(11284) <= 1'b0;
    layer1_outputs(11285) <= not a;
    layer1_outputs(11286) <= a;
    layer1_outputs(11287) <= not (a and b);
    layer1_outputs(11288) <= not (a and b);
    layer1_outputs(11289) <= not b;
    layer1_outputs(11290) <= not (a and b);
    layer1_outputs(11291) <= not b or a;
    layer1_outputs(11292) <= a xor b;
    layer1_outputs(11293) <= not (a or b);
    layer1_outputs(11294) <= a;
    layer1_outputs(11295) <= not b;
    layer1_outputs(11296) <= b;
    layer1_outputs(11297) <= a;
    layer1_outputs(11298) <= a and not b;
    layer1_outputs(11299) <= a or b;
    layer1_outputs(11300) <= a and not b;
    layer1_outputs(11301) <= a or b;
    layer1_outputs(11302) <= not (a xor b);
    layer1_outputs(11303) <= not (a xor b);
    layer1_outputs(11304) <= not a;
    layer1_outputs(11305) <= not (a xor b);
    layer1_outputs(11306) <= not b;
    layer1_outputs(11307) <= a and b;
    layer1_outputs(11308) <= not (a or b);
    layer1_outputs(11309) <= not a;
    layer1_outputs(11310) <= a and b;
    layer1_outputs(11311) <= a or b;
    layer1_outputs(11312) <= not (a and b);
    layer1_outputs(11313) <= not b or a;
    layer1_outputs(11314) <= a or b;
    layer1_outputs(11315) <= a xor b;
    layer1_outputs(11316) <= a;
    layer1_outputs(11317) <= b and not a;
    layer1_outputs(11318) <= a and b;
    layer1_outputs(11319) <= a xor b;
    layer1_outputs(11320) <= not a;
    layer1_outputs(11321) <= b and not a;
    layer1_outputs(11322) <= not b;
    layer1_outputs(11323) <= not a;
    layer1_outputs(11324) <= not a;
    layer1_outputs(11325) <= not (a xor b);
    layer1_outputs(11326) <= a and b;
    layer1_outputs(11327) <= a xor b;
    layer1_outputs(11328) <= not (a xor b);
    layer1_outputs(11329) <= not b;
    layer1_outputs(11330) <= b and not a;
    layer1_outputs(11331) <= not b;
    layer1_outputs(11332) <= not b;
    layer1_outputs(11333) <= not (a or b);
    layer1_outputs(11334) <= b;
    layer1_outputs(11335) <= a and b;
    layer1_outputs(11336) <= b;
    layer1_outputs(11337) <= a and b;
    layer1_outputs(11338) <= b and not a;
    layer1_outputs(11339) <= not a or b;
    layer1_outputs(11340) <= not (a and b);
    layer1_outputs(11341) <= a xor b;
    layer1_outputs(11342) <= not (a and b);
    layer1_outputs(11343) <= b;
    layer1_outputs(11344) <= a and b;
    layer1_outputs(11345) <= not a or b;
    layer1_outputs(11346) <= not b or a;
    layer1_outputs(11347) <= a;
    layer1_outputs(11348) <= a xor b;
    layer1_outputs(11349) <= b and not a;
    layer1_outputs(11350) <= a xor b;
    layer1_outputs(11351) <= not (a or b);
    layer1_outputs(11352) <= a and b;
    layer1_outputs(11353) <= not (a or b);
    layer1_outputs(11354) <= not (a and b);
    layer1_outputs(11355) <= not b;
    layer1_outputs(11356) <= a;
    layer1_outputs(11357) <= not a;
    layer1_outputs(11358) <= b and not a;
    layer1_outputs(11359) <= not (a and b);
    layer1_outputs(11360) <= a or b;
    layer1_outputs(11361) <= not b;
    layer1_outputs(11362) <= b and not a;
    layer1_outputs(11363) <= not (a and b);
    layer1_outputs(11364) <= a xor b;
    layer1_outputs(11365) <= a and b;
    layer1_outputs(11366) <= a and b;
    layer1_outputs(11367) <= a or b;
    layer1_outputs(11368) <= a and not b;
    layer1_outputs(11369) <= b;
    layer1_outputs(11370) <= b and not a;
    layer1_outputs(11371) <= not (a and b);
    layer1_outputs(11372) <= a;
    layer1_outputs(11373) <= a;
    layer1_outputs(11374) <= not (a or b);
    layer1_outputs(11375) <= not a or b;
    layer1_outputs(11376) <= not (a and b);
    layer1_outputs(11377) <= a and not b;
    layer1_outputs(11378) <= a and not b;
    layer1_outputs(11379) <= not (a and b);
    layer1_outputs(11380) <= b and not a;
    layer1_outputs(11381) <= not a;
    layer1_outputs(11382) <= b;
    layer1_outputs(11383) <= a;
    layer1_outputs(11384) <= not a;
    layer1_outputs(11385) <= not (a xor b);
    layer1_outputs(11386) <= not b;
    layer1_outputs(11387) <= not (a or b);
    layer1_outputs(11388) <= a and not b;
    layer1_outputs(11389) <= not b or a;
    layer1_outputs(11390) <= not a or b;
    layer1_outputs(11391) <= a or b;
    layer1_outputs(11392) <= b and not a;
    layer1_outputs(11393) <= not a or b;
    layer1_outputs(11394) <= not (a xor b);
    layer1_outputs(11395) <= not b or a;
    layer1_outputs(11396) <= not (a and b);
    layer1_outputs(11397) <= a and b;
    layer1_outputs(11398) <= b and not a;
    layer1_outputs(11399) <= not a;
    layer1_outputs(11400) <= b and not a;
    layer1_outputs(11401) <= b;
    layer1_outputs(11402) <= not a;
    layer1_outputs(11403) <= a xor b;
    layer1_outputs(11404) <= a xor b;
    layer1_outputs(11405) <= not a or b;
    layer1_outputs(11406) <= b;
    layer1_outputs(11407) <= not a;
    layer1_outputs(11408) <= not a;
    layer1_outputs(11409) <= a and not b;
    layer1_outputs(11410) <= a and b;
    layer1_outputs(11411) <= not a or b;
    layer1_outputs(11412) <= b;
    layer1_outputs(11413) <= not b;
    layer1_outputs(11414) <= a and b;
    layer1_outputs(11415) <= not (a or b);
    layer1_outputs(11416) <= not (a xor b);
    layer1_outputs(11417) <= b;
    layer1_outputs(11418) <= a or b;
    layer1_outputs(11419) <= not b;
    layer1_outputs(11420) <= not a or b;
    layer1_outputs(11421) <= a xor b;
    layer1_outputs(11422) <= a and not b;
    layer1_outputs(11423) <= not (a and b);
    layer1_outputs(11424) <= a;
    layer1_outputs(11425) <= not (a xor b);
    layer1_outputs(11426) <= a xor b;
    layer1_outputs(11427) <= a;
    layer1_outputs(11428) <= not b;
    layer1_outputs(11429) <= not (a xor b);
    layer1_outputs(11430) <= not b or a;
    layer1_outputs(11431) <= a and b;
    layer1_outputs(11432) <= not (a or b);
    layer1_outputs(11433) <= not (a and b);
    layer1_outputs(11434) <= a xor b;
    layer1_outputs(11435) <= b;
    layer1_outputs(11436) <= not a;
    layer1_outputs(11437) <= not (a and b);
    layer1_outputs(11438) <= not b;
    layer1_outputs(11439) <= b;
    layer1_outputs(11440) <= a xor b;
    layer1_outputs(11441) <= not (a xor b);
    layer1_outputs(11442) <= a and not b;
    layer1_outputs(11443) <= not b;
    layer1_outputs(11444) <= a or b;
    layer1_outputs(11445) <= a;
    layer1_outputs(11446) <= not a or b;
    layer1_outputs(11447) <= not a or b;
    layer1_outputs(11448) <= not (a and b);
    layer1_outputs(11449) <= a;
    layer1_outputs(11450) <= not a;
    layer1_outputs(11451) <= a and not b;
    layer1_outputs(11452) <= a;
    layer1_outputs(11453) <= not b or a;
    layer1_outputs(11454) <= 1'b1;
    layer1_outputs(11455) <= a;
    layer1_outputs(11456) <= not a or b;
    layer1_outputs(11457) <= a;
    layer1_outputs(11458) <= not (a or b);
    layer1_outputs(11459) <= b;
    layer1_outputs(11460) <= not (a and b);
    layer1_outputs(11461) <= not (a xor b);
    layer1_outputs(11462) <= not b or a;
    layer1_outputs(11463) <= not a or b;
    layer1_outputs(11464) <= not a;
    layer1_outputs(11465) <= a and not b;
    layer1_outputs(11466) <= b and not a;
    layer1_outputs(11467) <= a;
    layer1_outputs(11468) <= not b;
    layer1_outputs(11469) <= not (a and b);
    layer1_outputs(11470) <= not a;
    layer1_outputs(11471) <= not b;
    layer1_outputs(11472) <= not (a and b);
    layer1_outputs(11473) <= not b or a;
    layer1_outputs(11474) <= not b;
    layer1_outputs(11475) <= not b;
    layer1_outputs(11476) <= not (a xor b);
    layer1_outputs(11477) <= not b;
    layer1_outputs(11478) <= a or b;
    layer1_outputs(11479) <= a;
    layer1_outputs(11480) <= not b or a;
    layer1_outputs(11481) <= not a;
    layer1_outputs(11482) <= not b or a;
    layer1_outputs(11483) <= a and b;
    layer1_outputs(11484) <= a and b;
    layer1_outputs(11485) <= a;
    layer1_outputs(11486) <= a and not b;
    layer1_outputs(11487) <= b and not a;
    layer1_outputs(11488) <= not (a xor b);
    layer1_outputs(11489) <= b;
    layer1_outputs(11490) <= not a;
    layer1_outputs(11491) <= a xor b;
    layer1_outputs(11492) <= not b;
    layer1_outputs(11493) <= not a;
    layer1_outputs(11494) <= not a or b;
    layer1_outputs(11495) <= not (a and b);
    layer1_outputs(11496) <= b and not a;
    layer1_outputs(11497) <= a and not b;
    layer1_outputs(11498) <= b and not a;
    layer1_outputs(11499) <= b;
    layer1_outputs(11500) <= a;
    layer1_outputs(11501) <= a and b;
    layer1_outputs(11502) <= not a;
    layer1_outputs(11503) <= b and not a;
    layer1_outputs(11504) <= not a;
    layer1_outputs(11505) <= not (a xor b);
    layer1_outputs(11506) <= b;
    layer1_outputs(11507) <= a xor b;
    layer1_outputs(11508) <= b and not a;
    layer1_outputs(11509) <= not b or a;
    layer1_outputs(11510) <= not a;
    layer1_outputs(11511) <= b;
    layer1_outputs(11512) <= a and b;
    layer1_outputs(11513) <= a xor b;
    layer1_outputs(11514) <= a xor b;
    layer1_outputs(11515) <= a and not b;
    layer1_outputs(11516) <= a xor b;
    layer1_outputs(11517) <= b;
    layer1_outputs(11518) <= not (a xor b);
    layer1_outputs(11519) <= a and b;
    layer1_outputs(11520) <= not (a xor b);
    layer1_outputs(11521) <= a and b;
    layer1_outputs(11522) <= not (a or b);
    layer1_outputs(11523) <= a or b;
    layer1_outputs(11524) <= a and not b;
    layer1_outputs(11525) <= a;
    layer1_outputs(11526) <= b;
    layer1_outputs(11527) <= a;
    layer1_outputs(11528) <= not a;
    layer1_outputs(11529) <= not (a xor b);
    layer1_outputs(11530) <= b;
    layer1_outputs(11531) <= a and not b;
    layer1_outputs(11532) <= b;
    layer1_outputs(11533) <= b and not a;
    layer1_outputs(11534) <= not a or b;
    layer1_outputs(11535) <= a or b;
    layer1_outputs(11536) <= not a or b;
    layer1_outputs(11537) <= not (a xor b);
    layer1_outputs(11538) <= a;
    layer1_outputs(11539) <= a and not b;
    layer1_outputs(11540) <= not b or a;
    layer1_outputs(11541) <= b;
    layer1_outputs(11542) <= not b;
    layer1_outputs(11543) <= b;
    layer1_outputs(11544) <= not (a xor b);
    layer1_outputs(11545) <= a;
    layer1_outputs(11546) <= a;
    layer1_outputs(11547) <= a and b;
    layer1_outputs(11548) <= a or b;
    layer1_outputs(11549) <= not b;
    layer1_outputs(11550) <= not a;
    layer1_outputs(11551) <= not b;
    layer1_outputs(11552) <= not (a and b);
    layer1_outputs(11553) <= not a;
    layer1_outputs(11554) <= b;
    layer1_outputs(11555) <= a xor b;
    layer1_outputs(11556) <= b;
    layer1_outputs(11557) <= 1'b0;
    layer1_outputs(11558) <= b and not a;
    layer1_outputs(11559) <= b and not a;
    layer1_outputs(11560) <= not b;
    layer1_outputs(11561) <= a and not b;
    layer1_outputs(11562) <= a or b;
    layer1_outputs(11563) <= b;
    layer1_outputs(11564) <= a;
    layer1_outputs(11565) <= b;
    layer1_outputs(11566) <= a or b;
    layer1_outputs(11567) <= not (a or b);
    layer1_outputs(11568) <= not b or a;
    layer1_outputs(11569) <= a;
    layer1_outputs(11570) <= a;
    layer1_outputs(11571) <= not b;
    layer1_outputs(11572) <= not b or a;
    layer1_outputs(11573) <= a or b;
    layer1_outputs(11574) <= not (a xor b);
    layer1_outputs(11575) <= not (a or b);
    layer1_outputs(11576) <= not (a and b);
    layer1_outputs(11577) <= not (a xor b);
    layer1_outputs(11578) <= a;
    layer1_outputs(11579) <= b and not a;
    layer1_outputs(11580) <= not b or a;
    layer1_outputs(11581) <= not a;
    layer1_outputs(11582) <= b;
    layer1_outputs(11583) <= not b;
    layer1_outputs(11584) <= not b;
    layer1_outputs(11585) <= a and b;
    layer1_outputs(11586) <= b;
    layer1_outputs(11587) <= a;
    layer1_outputs(11588) <= not a or b;
    layer1_outputs(11589) <= not a or b;
    layer1_outputs(11590) <= a and b;
    layer1_outputs(11591) <= not a or b;
    layer1_outputs(11592) <= b;
    layer1_outputs(11593) <= b and not a;
    layer1_outputs(11594) <= a or b;
    layer1_outputs(11595) <= b and not a;
    layer1_outputs(11596) <= not (a and b);
    layer1_outputs(11597) <= a;
    layer1_outputs(11598) <= not b;
    layer1_outputs(11599) <= not (a or b);
    layer1_outputs(11600) <= not b;
    layer1_outputs(11601) <= not b;
    layer1_outputs(11602) <= not (a or b);
    layer1_outputs(11603) <= not (a and b);
    layer1_outputs(11604) <= not b;
    layer1_outputs(11605) <= a and b;
    layer1_outputs(11606) <= 1'b0;
    layer1_outputs(11607) <= not (a or b);
    layer1_outputs(11608) <= a;
    layer1_outputs(11609) <= not b;
    layer1_outputs(11610) <= a or b;
    layer1_outputs(11611) <= not a;
    layer1_outputs(11612) <= not (a xor b);
    layer1_outputs(11613) <= not a or b;
    layer1_outputs(11614) <= not (a or b);
    layer1_outputs(11615) <= not a or b;
    layer1_outputs(11616) <= b and not a;
    layer1_outputs(11617) <= not b or a;
    layer1_outputs(11618) <= not a;
    layer1_outputs(11619) <= a and not b;
    layer1_outputs(11620) <= not (a xor b);
    layer1_outputs(11621) <= a xor b;
    layer1_outputs(11622) <= not (a xor b);
    layer1_outputs(11623) <= a;
    layer1_outputs(11624) <= not (a xor b);
    layer1_outputs(11625) <= b;
    layer1_outputs(11626) <= b;
    layer1_outputs(11627) <= not b;
    layer1_outputs(11628) <= not a;
    layer1_outputs(11629) <= not (a xor b);
    layer1_outputs(11630) <= a and b;
    layer1_outputs(11631) <= a;
    layer1_outputs(11632) <= b and not a;
    layer1_outputs(11633) <= a;
    layer1_outputs(11634) <= a xor b;
    layer1_outputs(11635) <= not (a and b);
    layer1_outputs(11636) <= not a;
    layer1_outputs(11637) <= not a;
    layer1_outputs(11638) <= 1'b0;
    layer1_outputs(11639) <= not b;
    layer1_outputs(11640) <= not b or a;
    layer1_outputs(11641) <= not a;
    layer1_outputs(11642) <= not (a xor b);
    layer1_outputs(11643) <= not (a xor b);
    layer1_outputs(11644) <= not b or a;
    layer1_outputs(11645) <= a and not b;
    layer1_outputs(11646) <= a and not b;
    layer1_outputs(11647) <= a or b;
    layer1_outputs(11648) <= a and not b;
    layer1_outputs(11649) <= a and not b;
    layer1_outputs(11650) <= not a;
    layer1_outputs(11651) <= b and not a;
    layer1_outputs(11652) <= b;
    layer1_outputs(11653) <= not a or b;
    layer1_outputs(11654) <= b;
    layer1_outputs(11655) <= 1'b0;
    layer1_outputs(11656) <= b;
    layer1_outputs(11657) <= a;
    layer1_outputs(11658) <= not b or a;
    layer1_outputs(11659) <= not (a xor b);
    layer1_outputs(11660) <= a or b;
    layer1_outputs(11661) <= a;
    layer1_outputs(11662) <= not a;
    layer1_outputs(11663) <= not (a or b);
    layer1_outputs(11664) <= b and not a;
    layer1_outputs(11665) <= a or b;
    layer1_outputs(11666) <= b and not a;
    layer1_outputs(11667) <= not (a xor b);
    layer1_outputs(11668) <= a;
    layer1_outputs(11669) <= b;
    layer1_outputs(11670) <= a xor b;
    layer1_outputs(11671) <= not a;
    layer1_outputs(11672) <= not (a xor b);
    layer1_outputs(11673) <= a xor b;
    layer1_outputs(11674) <= not (a xor b);
    layer1_outputs(11675) <= b;
    layer1_outputs(11676) <= a xor b;
    layer1_outputs(11677) <= a or b;
    layer1_outputs(11678) <= b;
    layer1_outputs(11679) <= a and not b;
    layer1_outputs(11680) <= a;
    layer1_outputs(11681) <= not a or b;
    layer1_outputs(11682) <= a and b;
    layer1_outputs(11683) <= a xor b;
    layer1_outputs(11684) <= not a;
    layer1_outputs(11685) <= not (a xor b);
    layer1_outputs(11686) <= a and not b;
    layer1_outputs(11687) <= b;
    layer1_outputs(11688) <= not a or b;
    layer1_outputs(11689) <= 1'b1;
    layer1_outputs(11690) <= not (a xor b);
    layer1_outputs(11691) <= not b;
    layer1_outputs(11692) <= a and not b;
    layer1_outputs(11693) <= a and b;
    layer1_outputs(11694) <= 1'b1;
    layer1_outputs(11695) <= not a;
    layer1_outputs(11696) <= not (a xor b);
    layer1_outputs(11697) <= b;
    layer1_outputs(11698) <= a or b;
    layer1_outputs(11699) <= not (a and b);
    layer1_outputs(11700) <= a xor b;
    layer1_outputs(11701) <= not (a or b);
    layer1_outputs(11702) <= not a;
    layer1_outputs(11703) <= not (a or b);
    layer1_outputs(11704) <= not b;
    layer1_outputs(11705) <= not b or a;
    layer1_outputs(11706) <= not b or a;
    layer1_outputs(11707) <= b;
    layer1_outputs(11708) <= not (a or b);
    layer1_outputs(11709) <= a or b;
    layer1_outputs(11710) <= b;
    layer1_outputs(11711) <= a and not b;
    layer1_outputs(11712) <= not (a xor b);
    layer1_outputs(11713) <= not a;
    layer1_outputs(11714) <= not (a or b);
    layer1_outputs(11715) <= a;
    layer1_outputs(11716) <= a;
    layer1_outputs(11717) <= not a or b;
    layer1_outputs(11718) <= b and not a;
    layer1_outputs(11719) <= not b;
    layer1_outputs(11720) <= not b or a;
    layer1_outputs(11721) <= a or b;
    layer1_outputs(11722) <= not (a and b);
    layer1_outputs(11723) <= not b;
    layer1_outputs(11724) <= 1'b1;
    layer1_outputs(11725) <= not (a xor b);
    layer1_outputs(11726) <= a or b;
    layer1_outputs(11727) <= not a or b;
    layer1_outputs(11728) <= a xor b;
    layer1_outputs(11729) <= not (a and b);
    layer1_outputs(11730) <= a xor b;
    layer1_outputs(11731) <= not (a and b);
    layer1_outputs(11732) <= a and b;
    layer1_outputs(11733) <= not a;
    layer1_outputs(11734) <= not (a or b);
    layer1_outputs(11735) <= b;
    layer1_outputs(11736) <= b;
    layer1_outputs(11737) <= not a;
    layer1_outputs(11738) <= not a;
    layer1_outputs(11739) <= not a or b;
    layer1_outputs(11740) <= not a;
    layer1_outputs(11741) <= a and b;
    layer1_outputs(11742) <= not b;
    layer1_outputs(11743) <= b;
    layer1_outputs(11744) <= not b;
    layer1_outputs(11745) <= not b;
    layer1_outputs(11746) <= not b;
    layer1_outputs(11747) <= b;
    layer1_outputs(11748) <= not (a or b);
    layer1_outputs(11749) <= not (a xor b);
    layer1_outputs(11750) <= not a;
    layer1_outputs(11751) <= b and not a;
    layer1_outputs(11752) <= not (a xor b);
    layer1_outputs(11753) <= not a or b;
    layer1_outputs(11754) <= a and not b;
    layer1_outputs(11755) <= not (a xor b);
    layer1_outputs(11756) <= a;
    layer1_outputs(11757) <= a;
    layer1_outputs(11758) <= not a;
    layer1_outputs(11759) <= a and not b;
    layer1_outputs(11760) <= b;
    layer1_outputs(11761) <= not (a or b);
    layer1_outputs(11762) <= a and not b;
    layer1_outputs(11763) <= not b;
    layer1_outputs(11764) <= a and not b;
    layer1_outputs(11765) <= not a or b;
    layer1_outputs(11766) <= a xor b;
    layer1_outputs(11767) <= b;
    layer1_outputs(11768) <= a xor b;
    layer1_outputs(11769) <= a xor b;
    layer1_outputs(11770) <= not (a and b);
    layer1_outputs(11771) <= not b;
    layer1_outputs(11772) <= a and not b;
    layer1_outputs(11773) <= a and b;
    layer1_outputs(11774) <= not b or a;
    layer1_outputs(11775) <= a;
    layer1_outputs(11776) <= not a or b;
    layer1_outputs(11777) <= not (a and b);
    layer1_outputs(11778) <= a;
    layer1_outputs(11779) <= not a or b;
    layer1_outputs(11780) <= b;
    layer1_outputs(11781) <= not (a or b);
    layer1_outputs(11782) <= not b or a;
    layer1_outputs(11783) <= b and not a;
    layer1_outputs(11784) <= a or b;
    layer1_outputs(11785) <= not b or a;
    layer1_outputs(11786) <= not a;
    layer1_outputs(11787) <= b and not a;
    layer1_outputs(11788) <= not a;
    layer1_outputs(11789) <= not (a and b);
    layer1_outputs(11790) <= not (a xor b);
    layer1_outputs(11791) <= a or b;
    layer1_outputs(11792) <= a xor b;
    layer1_outputs(11793) <= a;
    layer1_outputs(11794) <= not (a and b);
    layer1_outputs(11795) <= not a or b;
    layer1_outputs(11796) <= a xor b;
    layer1_outputs(11797) <= a and b;
    layer1_outputs(11798) <= not a;
    layer1_outputs(11799) <= not (a or b);
    layer1_outputs(11800) <= not a;
    layer1_outputs(11801) <= not b or a;
    layer1_outputs(11802) <= not (a and b);
    layer1_outputs(11803) <= b and not a;
    layer1_outputs(11804) <= a and not b;
    layer1_outputs(11805) <= not a or b;
    layer1_outputs(11806) <= a and not b;
    layer1_outputs(11807) <= 1'b1;
    layer1_outputs(11808) <= not b;
    layer1_outputs(11809) <= not (a or b);
    layer1_outputs(11810) <= not (a and b);
    layer1_outputs(11811) <= not a or b;
    layer1_outputs(11812) <= not a;
    layer1_outputs(11813) <= a and not b;
    layer1_outputs(11814) <= a;
    layer1_outputs(11815) <= a xor b;
    layer1_outputs(11816) <= a or b;
    layer1_outputs(11817) <= not b;
    layer1_outputs(11818) <= not (a and b);
    layer1_outputs(11819) <= a and b;
    layer1_outputs(11820) <= b and not a;
    layer1_outputs(11821) <= not a;
    layer1_outputs(11822) <= b;
    layer1_outputs(11823) <= a or b;
    layer1_outputs(11824) <= a and not b;
    layer1_outputs(11825) <= a or b;
    layer1_outputs(11826) <= a or b;
    layer1_outputs(11827) <= b and not a;
    layer1_outputs(11828) <= a and not b;
    layer1_outputs(11829) <= not (a xor b);
    layer1_outputs(11830) <= b;
    layer1_outputs(11831) <= b;
    layer1_outputs(11832) <= a and b;
    layer1_outputs(11833) <= not (a xor b);
    layer1_outputs(11834) <= b;
    layer1_outputs(11835) <= not a;
    layer1_outputs(11836) <= not b;
    layer1_outputs(11837) <= not a;
    layer1_outputs(11838) <= a and b;
    layer1_outputs(11839) <= a or b;
    layer1_outputs(11840) <= a and b;
    layer1_outputs(11841) <= not a;
    layer1_outputs(11842) <= not b or a;
    layer1_outputs(11843) <= not (a and b);
    layer1_outputs(11844) <= not a or b;
    layer1_outputs(11845) <= b;
    layer1_outputs(11846) <= not b;
    layer1_outputs(11847) <= b and not a;
    layer1_outputs(11848) <= not (a xor b);
    layer1_outputs(11849) <= a and not b;
    layer1_outputs(11850) <= not (a or b);
    layer1_outputs(11851) <= b and not a;
    layer1_outputs(11852) <= a and not b;
    layer1_outputs(11853) <= not (a and b);
    layer1_outputs(11854) <= not b;
    layer1_outputs(11855) <= not (a or b);
    layer1_outputs(11856) <= not (a or b);
    layer1_outputs(11857) <= not b;
    layer1_outputs(11858) <= not (a and b);
    layer1_outputs(11859) <= not (a xor b);
    layer1_outputs(11860) <= b and not a;
    layer1_outputs(11861) <= a and not b;
    layer1_outputs(11862) <= not (a xor b);
    layer1_outputs(11863) <= a or b;
    layer1_outputs(11864) <= not a or b;
    layer1_outputs(11865) <= b and not a;
    layer1_outputs(11866) <= b and not a;
    layer1_outputs(11867) <= not (a and b);
    layer1_outputs(11868) <= a;
    layer1_outputs(11869) <= a;
    layer1_outputs(11870) <= not (a or b);
    layer1_outputs(11871) <= a xor b;
    layer1_outputs(11872) <= not (a xor b);
    layer1_outputs(11873) <= b;
    layer1_outputs(11874) <= a;
    layer1_outputs(11875) <= b;
    layer1_outputs(11876) <= b and not a;
    layer1_outputs(11877) <= not b or a;
    layer1_outputs(11878) <= not (a and b);
    layer1_outputs(11879) <= b and not a;
    layer1_outputs(11880) <= not a;
    layer1_outputs(11881) <= a or b;
    layer1_outputs(11882) <= a and b;
    layer1_outputs(11883) <= not (a xor b);
    layer1_outputs(11884) <= a;
    layer1_outputs(11885) <= a;
    layer1_outputs(11886) <= a xor b;
    layer1_outputs(11887) <= a;
    layer1_outputs(11888) <= not b;
    layer1_outputs(11889) <= 1'b1;
    layer1_outputs(11890) <= not b;
    layer1_outputs(11891) <= not (a and b);
    layer1_outputs(11892) <= b;
    layer1_outputs(11893) <= a xor b;
    layer1_outputs(11894) <= not a or b;
    layer1_outputs(11895) <= a and not b;
    layer1_outputs(11896) <= a;
    layer1_outputs(11897) <= a and b;
    layer1_outputs(11898) <= a;
    layer1_outputs(11899) <= not a;
    layer1_outputs(11900) <= not (a and b);
    layer1_outputs(11901) <= a and b;
    layer1_outputs(11902) <= a and b;
    layer1_outputs(11903) <= a;
    layer1_outputs(11904) <= a and not b;
    layer1_outputs(11905) <= not a;
    layer1_outputs(11906) <= b;
    layer1_outputs(11907) <= a and not b;
    layer1_outputs(11908) <= a and b;
    layer1_outputs(11909) <= not a;
    layer1_outputs(11910) <= not (a and b);
    layer1_outputs(11911) <= not (a and b);
    layer1_outputs(11912) <= not a or b;
    layer1_outputs(11913) <= b;
    layer1_outputs(11914) <= a and b;
    layer1_outputs(11915) <= not (a xor b);
    layer1_outputs(11916) <= b and not a;
    layer1_outputs(11917) <= b;
    layer1_outputs(11918) <= a or b;
    layer1_outputs(11919) <= not (a and b);
    layer1_outputs(11920) <= 1'b1;
    layer1_outputs(11921) <= a or b;
    layer1_outputs(11922) <= not (a and b);
    layer1_outputs(11923) <= a xor b;
    layer1_outputs(11924) <= a and not b;
    layer1_outputs(11925) <= 1'b1;
    layer1_outputs(11926) <= a or b;
    layer1_outputs(11927) <= not b;
    layer1_outputs(11928) <= not b;
    layer1_outputs(11929) <= a or b;
    layer1_outputs(11930) <= a;
    layer1_outputs(11931) <= a;
    layer1_outputs(11932) <= a and not b;
    layer1_outputs(11933) <= not b;
    layer1_outputs(11934) <= b;
    layer1_outputs(11935) <= not b or a;
    layer1_outputs(11936) <= 1'b1;
    layer1_outputs(11937) <= a and b;
    layer1_outputs(11938) <= b and not a;
    layer1_outputs(11939) <= a or b;
    layer1_outputs(11940) <= a and b;
    layer1_outputs(11941) <= not b;
    layer1_outputs(11942) <= not (a and b);
    layer1_outputs(11943) <= a xor b;
    layer1_outputs(11944) <= not b;
    layer1_outputs(11945) <= not b;
    layer1_outputs(11946) <= not b or a;
    layer1_outputs(11947) <= not a;
    layer1_outputs(11948) <= not a;
    layer1_outputs(11949) <= not (a or b);
    layer1_outputs(11950) <= not a;
    layer1_outputs(11951) <= 1'b0;
    layer1_outputs(11952) <= not (a and b);
    layer1_outputs(11953) <= a and not b;
    layer1_outputs(11954) <= 1'b0;
    layer1_outputs(11955) <= b and not a;
    layer1_outputs(11956) <= b;
    layer1_outputs(11957) <= not (a or b);
    layer1_outputs(11958) <= b;
    layer1_outputs(11959) <= a;
    layer1_outputs(11960) <= a and not b;
    layer1_outputs(11961) <= 1'b1;
    layer1_outputs(11962) <= a and not b;
    layer1_outputs(11963) <= a;
    layer1_outputs(11964) <= a;
    layer1_outputs(11965) <= a and not b;
    layer1_outputs(11966) <= a and b;
    layer1_outputs(11967) <= not b;
    layer1_outputs(11968) <= a xor b;
    layer1_outputs(11969) <= not (a xor b);
    layer1_outputs(11970) <= not a;
    layer1_outputs(11971) <= not (a or b);
    layer1_outputs(11972) <= not b;
    layer1_outputs(11973) <= a xor b;
    layer1_outputs(11974) <= b;
    layer1_outputs(11975) <= a;
    layer1_outputs(11976) <= not (a and b);
    layer1_outputs(11977) <= not (a xor b);
    layer1_outputs(11978) <= 1'b0;
    layer1_outputs(11979) <= not (a and b);
    layer1_outputs(11980) <= a;
    layer1_outputs(11981) <= b;
    layer1_outputs(11982) <= b and not a;
    layer1_outputs(11983) <= a xor b;
    layer1_outputs(11984) <= not (a xor b);
    layer1_outputs(11985) <= not b or a;
    layer1_outputs(11986) <= not a;
    layer1_outputs(11987) <= b;
    layer1_outputs(11988) <= b;
    layer1_outputs(11989) <= a;
    layer1_outputs(11990) <= b and not a;
    layer1_outputs(11991) <= not (a xor b);
    layer1_outputs(11992) <= a;
    layer1_outputs(11993) <= not (a xor b);
    layer1_outputs(11994) <= not (a xor b);
    layer1_outputs(11995) <= not a;
    layer1_outputs(11996) <= not b;
    layer1_outputs(11997) <= not (a and b);
    layer1_outputs(11998) <= 1'b1;
    layer1_outputs(11999) <= not (a and b);
    layer1_outputs(12000) <= not b;
    layer1_outputs(12001) <= not (a or b);
    layer1_outputs(12002) <= a and b;
    layer1_outputs(12003) <= not (a and b);
    layer1_outputs(12004) <= a xor b;
    layer1_outputs(12005) <= a or b;
    layer1_outputs(12006) <= 1'b0;
    layer1_outputs(12007) <= not (a or b);
    layer1_outputs(12008) <= not (a xor b);
    layer1_outputs(12009) <= a xor b;
    layer1_outputs(12010) <= not b;
    layer1_outputs(12011) <= not (a or b);
    layer1_outputs(12012) <= b and not a;
    layer1_outputs(12013) <= 1'b1;
    layer1_outputs(12014) <= not a;
    layer1_outputs(12015) <= a xor b;
    layer1_outputs(12016) <= a and b;
    layer1_outputs(12017) <= a;
    layer1_outputs(12018) <= not a;
    layer1_outputs(12019) <= a xor b;
    layer1_outputs(12020) <= not a;
    layer1_outputs(12021) <= a xor b;
    layer1_outputs(12022) <= not (a or b);
    layer1_outputs(12023) <= not b or a;
    layer1_outputs(12024) <= b;
    layer1_outputs(12025) <= not (a or b);
    layer1_outputs(12026) <= a or b;
    layer1_outputs(12027) <= not a or b;
    layer1_outputs(12028) <= a xor b;
    layer1_outputs(12029) <= a;
    layer1_outputs(12030) <= not b or a;
    layer1_outputs(12031) <= b;
    layer1_outputs(12032) <= a;
    layer1_outputs(12033) <= not a;
    layer1_outputs(12034) <= not (a xor b);
    layer1_outputs(12035) <= not b;
    layer1_outputs(12036) <= a or b;
    layer1_outputs(12037) <= not a or b;
    layer1_outputs(12038) <= b and not a;
    layer1_outputs(12039) <= a;
    layer1_outputs(12040) <= not (a xor b);
    layer1_outputs(12041) <= not (a or b);
    layer1_outputs(12042) <= a or b;
    layer1_outputs(12043) <= not b or a;
    layer1_outputs(12044) <= b;
    layer1_outputs(12045) <= a and not b;
    layer1_outputs(12046) <= a xor b;
    layer1_outputs(12047) <= not (a xor b);
    layer1_outputs(12048) <= b and not a;
    layer1_outputs(12049) <= not a;
    layer1_outputs(12050) <= a xor b;
    layer1_outputs(12051) <= a;
    layer1_outputs(12052) <= not a;
    layer1_outputs(12053) <= not (a and b);
    layer1_outputs(12054) <= a or b;
    layer1_outputs(12055) <= 1'b0;
    layer1_outputs(12056) <= a;
    layer1_outputs(12057) <= not (a and b);
    layer1_outputs(12058) <= not (a and b);
    layer1_outputs(12059) <= b;
    layer1_outputs(12060) <= not (a xor b);
    layer1_outputs(12061) <= not (a or b);
    layer1_outputs(12062) <= not (a and b);
    layer1_outputs(12063) <= not (a xor b);
    layer1_outputs(12064) <= b and not a;
    layer1_outputs(12065) <= a and not b;
    layer1_outputs(12066) <= not a;
    layer1_outputs(12067) <= b and not a;
    layer1_outputs(12068) <= not a or b;
    layer1_outputs(12069) <= a;
    layer1_outputs(12070) <= a and b;
    layer1_outputs(12071) <= a and b;
    layer1_outputs(12072) <= not b or a;
    layer1_outputs(12073) <= not a or b;
    layer1_outputs(12074) <= b;
    layer1_outputs(12075) <= a or b;
    layer1_outputs(12076) <= not a;
    layer1_outputs(12077) <= b;
    layer1_outputs(12078) <= not a;
    layer1_outputs(12079) <= a and b;
    layer1_outputs(12080) <= not b or a;
    layer1_outputs(12081) <= not a;
    layer1_outputs(12082) <= not a or b;
    layer1_outputs(12083) <= not b or a;
    layer1_outputs(12084) <= a and b;
    layer1_outputs(12085) <= b;
    layer1_outputs(12086) <= not b;
    layer1_outputs(12087) <= b;
    layer1_outputs(12088) <= not (a and b);
    layer1_outputs(12089) <= a and b;
    layer1_outputs(12090) <= a;
    layer1_outputs(12091) <= not b;
    layer1_outputs(12092) <= b and not a;
    layer1_outputs(12093) <= a or b;
    layer1_outputs(12094) <= not (a or b);
    layer1_outputs(12095) <= not (a and b);
    layer1_outputs(12096) <= not (a or b);
    layer1_outputs(12097) <= not a;
    layer1_outputs(12098) <= b and not a;
    layer1_outputs(12099) <= b;
    layer1_outputs(12100) <= not b;
    layer1_outputs(12101) <= not a;
    layer1_outputs(12102) <= a or b;
    layer1_outputs(12103) <= a and b;
    layer1_outputs(12104) <= not (a xor b);
    layer1_outputs(12105) <= b;
    layer1_outputs(12106) <= not (a or b);
    layer1_outputs(12107) <= not (a or b);
    layer1_outputs(12108) <= a;
    layer1_outputs(12109) <= not a;
    layer1_outputs(12110) <= not (a xor b);
    layer1_outputs(12111) <= b;
    layer1_outputs(12112) <= not (a xor b);
    layer1_outputs(12113) <= a and b;
    layer1_outputs(12114) <= a xor b;
    layer1_outputs(12115) <= not b or a;
    layer1_outputs(12116) <= not (a xor b);
    layer1_outputs(12117) <= a and b;
    layer1_outputs(12118) <= not a;
    layer1_outputs(12119) <= a xor b;
    layer1_outputs(12120) <= b and not a;
    layer1_outputs(12121) <= not (a or b);
    layer1_outputs(12122) <= not (a xor b);
    layer1_outputs(12123) <= not (a xor b);
    layer1_outputs(12124) <= not a;
    layer1_outputs(12125) <= not a;
    layer1_outputs(12126) <= 1'b0;
    layer1_outputs(12127) <= a and b;
    layer1_outputs(12128) <= not (a and b);
    layer1_outputs(12129) <= b and not a;
    layer1_outputs(12130) <= not a;
    layer1_outputs(12131) <= a and not b;
    layer1_outputs(12132) <= b and not a;
    layer1_outputs(12133) <= not b or a;
    layer1_outputs(12134) <= b and not a;
    layer1_outputs(12135) <= not b or a;
    layer1_outputs(12136) <= 1'b1;
    layer1_outputs(12137) <= a and b;
    layer1_outputs(12138) <= b;
    layer1_outputs(12139) <= a xor b;
    layer1_outputs(12140) <= a or b;
    layer1_outputs(12141) <= not a;
    layer1_outputs(12142) <= a xor b;
    layer1_outputs(12143) <= not b;
    layer1_outputs(12144) <= b;
    layer1_outputs(12145) <= not b or a;
    layer1_outputs(12146) <= not b;
    layer1_outputs(12147) <= not (a and b);
    layer1_outputs(12148) <= a or b;
    layer1_outputs(12149) <= not a or b;
    layer1_outputs(12150) <= not (a xor b);
    layer1_outputs(12151) <= not b;
    layer1_outputs(12152) <= not b;
    layer1_outputs(12153) <= not b or a;
    layer1_outputs(12154) <= a and b;
    layer1_outputs(12155) <= b and not a;
    layer1_outputs(12156) <= not a or b;
    layer1_outputs(12157) <= not (a or b);
    layer1_outputs(12158) <= not b;
    layer1_outputs(12159) <= not (a and b);
    layer1_outputs(12160) <= a xor b;
    layer1_outputs(12161) <= a;
    layer1_outputs(12162) <= not a;
    layer1_outputs(12163) <= not a;
    layer1_outputs(12164) <= b and not a;
    layer1_outputs(12165) <= not b;
    layer1_outputs(12166) <= a;
    layer1_outputs(12167) <= b and not a;
    layer1_outputs(12168) <= not (a xor b);
    layer1_outputs(12169) <= not (a and b);
    layer1_outputs(12170) <= a and not b;
    layer1_outputs(12171) <= b and not a;
    layer1_outputs(12172) <= not b or a;
    layer1_outputs(12173) <= not b or a;
    layer1_outputs(12174) <= b;
    layer1_outputs(12175) <= not a or b;
    layer1_outputs(12176) <= a xor b;
    layer1_outputs(12177) <= not a;
    layer1_outputs(12178) <= not a;
    layer1_outputs(12179) <= a and not b;
    layer1_outputs(12180) <= b and not a;
    layer1_outputs(12181) <= b;
    layer1_outputs(12182) <= a and not b;
    layer1_outputs(12183) <= not a;
    layer1_outputs(12184) <= not a;
    layer1_outputs(12185) <= a and not b;
    layer1_outputs(12186) <= a and b;
    layer1_outputs(12187) <= not (a or b);
    layer1_outputs(12188) <= b;
    layer1_outputs(12189) <= not (a or b);
    layer1_outputs(12190) <= not b;
    layer1_outputs(12191) <= not (a and b);
    layer1_outputs(12192) <= a and not b;
    layer1_outputs(12193) <= a;
    layer1_outputs(12194) <= b;
    layer1_outputs(12195) <= not b;
    layer1_outputs(12196) <= a and b;
    layer1_outputs(12197) <= 1'b0;
    layer1_outputs(12198) <= not b or a;
    layer1_outputs(12199) <= a;
    layer1_outputs(12200) <= a and b;
    layer1_outputs(12201) <= not a or b;
    layer1_outputs(12202) <= b;
    layer1_outputs(12203) <= not (a and b);
    layer1_outputs(12204) <= not (a xor b);
    layer1_outputs(12205) <= a xor b;
    layer1_outputs(12206) <= not a or b;
    layer1_outputs(12207) <= b;
    layer1_outputs(12208) <= not a;
    layer1_outputs(12209) <= b and not a;
    layer1_outputs(12210) <= not b or a;
    layer1_outputs(12211) <= a or b;
    layer1_outputs(12212) <= a;
    layer1_outputs(12213) <= not (a xor b);
    layer1_outputs(12214) <= a or b;
    layer1_outputs(12215) <= not (a xor b);
    layer1_outputs(12216) <= not a or b;
    layer1_outputs(12217) <= not a or b;
    layer1_outputs(12218) <= not a;
    layer1_outputs(12219) <= a;
    layer1_outputs(12220) <= not b;
    layer1_outputs(12221) <= not b;
    layer1_outputs(12222) <= a xor b;
    layer1_outputs(12223) <= not b;
    layer1_outputs(12224) <= not b or a;
    layer1_outputs(12225) <= a;
    layer1_outputs(12226) <= a;
    layer1_outputs(12227) <= a and b;
    layer1_outputs(12228) <= a and b;
    layer1_outputs(12229) <= a or b;
    layer1_outputs(12230) <= not (a xor b);
    layer1_outputs(12231) <= not a;
    layer1_outputs(12232) <= not (a and b);
    layer1_outputs(12233) <= not b;
    layer1_outputs(12234) <= a and not b;
    layer1_outputs(12235) <= not a;
    layer1_outputs(12236) <= b and not a;
    layer1_outputs(12237) <= b;
    layer1_outputs(12238) <= not b or a;
    layer1_outputs(12239) <= not b;
    layer1_outputs(12240) <= not (a or b);
    layer1_outputs(12241) <= not (a and b);
    layer1_outputs(12242) <= not (a or b);
    layer1_outputs(12243) <= not a;
    layer1_outputs(12244) <= a and b;
    layer1_outputs(12245) <= a and b;
    layer1_outputs(12246) <= b and not a;
    layer1_outputs(12247) <= not a or b;
    layer1_outputs(12248) <= a;
    layer1_outputs(12249) <= b;
    layer1_outputs(12250) <= b;
    layer1_outputs(12251) <= not a or b;
    layer1_outputs(12252) <= a xor b;
    layer1_outputs(12253) <= a or b;
    layer1_outputs(12254) <= not (a xor b);
    layer1_outputs(12255) <= b;
    layer1_outputs(12256) <= a xor b;
    layer1_outputs(12257) <= not a;
    layer1_outputs(12258) <= b and not a;
    layer1_outputs(12259) <= a;
    layer1_outputs(12260) <= a xor b;
    layer1_outputs(12261) <= not (a xor b);
    layer1_outputs(12262) <= not (a or b);
    layer1_outputs(12263) <= b;
    layer1_outputs(12264) <= b;
    layer1_outputs(12265) <= b;
    layer1_outputs(12266) <= a and b;
    layer1_outputs(12267) <= a or b;
    layer1_outputs(12268) <= not (a xor b);
    layer1_outputs(12269) <= b;
    layer1_outputs(12270) <= a and b;
    layer1_outputs(12271) <= b and not a;
    layer1_outputs(12272) <= a or b;
    layer1_outputs(12273) <= not a;
    layer1_outputs(12274) <= a xor b;
    layer1_outputs(12275) <= not (a xor b);
    layer1_outputs(12276) <= not (a and b);
    layer1_outputs(12277) <= not a;
    layer1_outputs(12278) <= not (a or b);
    layer1_outputs(12279) <= b;
    layer1_outputs(12280) <= not (a and b);
    layer1_outputs(12281) <= not (a or b);
    layer1_outputs(12282) <= a or b;
    layer1_outputs(12283) <= not a;
    layer1_outputs(12284) <= b and not a;
    layer1_outputs(12285) <= not b;
    layer1_outputs(12286) <= a and b;
    layer1_outputs(12287) <= a or b;
    layer1_outputs(12288) <= b;
    layer1_outputs(12289) <= not b or a;
    layer1_outputs(12290) <= not (a xor b);
    layer1_outputs(12291) <= not b or a;
    layer1_outputs(12292) <= a;
    layer1_outputs(12293) <= a or b;
    layer1_outputs(12294) <= not a or b;
    layer1_outputs(12295) <= a and b;
    layer1_outputs(12296) <= not (a and b);
    layer1_outputs(12297) <= b;
    layer1_outputs(12298) <= not (a xor b);
    layer1_outputs(12299) <= b and not a;
    layer1_outputs(12300) <= a;
    layer1_outputs(12301) <= not a;
    layer1_outputs(12302) <= not b or a;
    layer1_outputs(12303) <= a and b;
    layer1_outputs(12304) <= a or b;
    layer1_outputs(12305) <= not a;
    layer1_outputs(12306) <= a or b;
    layer1_outputs(12307) <= a and b;
    layer1_outputs(12308) <= a or b;
    layer1_outputs(12309) <= b and not a;
    layer1_outputs(12310) <= not (a or b);
    layer1_outputs(12311) <= a and not b;
    layer1_outputs(12312) <= b;
    layer1_outputs(12313) <= a xor b;
    layer1_outputs(12314) <= not (a and b);
    layer1_outputs(12315) <= b;
    layer1_outputs(12316) <= not b or a;
    layer1_outputs(12317) <= not a or b;
    layer1_outputs(12318) <= a or b;
    layer1_outputs(12319) <= a and b;
    layer1_outputs(12320) <= not b or a;
    layer1_outputs(12321) <= not (a xor b);
    layer1_outputs(12322) <= not (a and b);
    layer1_outputs(12323) <= not a;
    layer1_outputs(12324) <= a and b;
    layer1_outputs(12325) <= not (a and b);
    layer1_outputs(12326) <= not a or b;
    layer1_outputs(12327) <= a;
    layer1_outputs(12328) <= 1'b1;
    layer1_outputs(12329) <= a;
    layer1_outputs(12330) <= a and b;
    layer1_outputs(12331) <= not a;
    layer1_outputs(12332) <= not b or a;
    layer1_outputs(12333) <= not b or a;
    layer1_outputs(12334) <= not (a or b);
    layer1_outputs(12335) <= b and not a;
    layer1_outputs(12336) <= a and b;
    layer1_outputs(12337) <= a;
    layer1_outputs(12338) <= not (a and b);
    layer1_outputs(12339) <= not (a xor b);
    layer1_outputs(12340) <= a and not b;
    layer1_outputs(12341) <= 1'b1;
    layer1_outputs(12342) <= not a;
    layer1_outputs(12343) <= not (a and b);
    layer1_outputs(12344) <= not a;
    layer1_outputs(12345) <= b and not a;
    layer1_outputs(12346) <= a xor b;
    layer1_outputs(12347) <= not (a and b);
    layer1_outputs(12348) <= a and not b;
    layer1_outputs(12349) <= not b or a;
    layer1_outputs(12350) <= not a;
    layer1_outputs(12351) <= not b;
    layer1_outputs(12352) <= not b or a;
    layer1_outputs(12353) <= a or b;
    layer1_outputs(12354) <= a and not b;
    layer1_outputs(12355) <= b;
    layer1_outputs(12356) <= a or b;
    layer1_outputs(12357) <= b;
    layer1_outputs(12358) <= not a or b;
    layer1_outputs(12359) <= not (a and b);
    layer1_outputs(12360) <= 1'b0;
    layer1_outputs(12361) <= not (a or b);
    layer1_outputs(12362) <= a xor b;
    layer1_outputs(12363) <= not b;
    layer1_outputs(12364) <= not a or b;
    layer1_outputs(12365) <= not b;
    layer1_outputs(12366) <= not a;
    layer1_outputs(12367) <= not a;
    layer1_outputs(12368) <= not b;
    layer1_outputs(12369) <= not (a or b);
    layer1_outputs(12370) <= a xor b;
    layer1_outputs(12371) <= not (a and b);
    layer1_outputs(12372) <= not b;
    layer1_outputs(12373) <= a xor b;
    layer1_outputs(12374) <= not a;
    layer1_outputs(12375) <= a and b;
    layer1_outputs(12376) <= b and not a;
    layer1_outputs(12377) <= b;
    layer1_outputs(12378) <= not (a and b);
    layer1_outputs(12379) <= not a or b;
    layer1_outputs(12380) <= not b or a;
    layer1_outputs(12381) <= a and not b;
    layer1_outputs(12382) <= not (a xor b);
    layer1_outputs(12383) <= not (a or b);
    layer1_outputs(12384) <= not b or a;
    layer1_outputs(12385) <= a;
    layer1_outputs(12386) <= b;
    layer1_outputs(12387) <= a or b;
    layer1_outputs(12388) <= a and not b;
    layer1_outputs(12389) <= not b or a;
    layer1_outputs(12390) <= b;
    layer1_outputs(12391) <= b and not a;
    layer1_outputs(12392) <= not b;
    layer1_outputs(12393) <= b and not a;
    layer1_outputs(12394) <= b;
    layer1_outputs(12395) <= not (a and b);
    layer1_outputs(12396) <= a or b;
    layer1_outputs(12397) <= not (a xor b);
    layer1_outputs(12398) <= not b;
    layer1_outputs(12399) <= not a or b;
    layer1_outputs(12400) <= a;
    layer1_outputs(12401) <= b;
    layer1_outputs(12402) <= not (a or b);
    layer1_outputs(12403) <= not (a xor b);
    layer1_outputs(12404) <= a and not b;
    layer1_outputs(12405) <= not (a xor b);
    layer1_outputs(12406) <= not b;
    layer1_outputs(12407) <= not a or b;
    layer1_outputs(12408) <= not b or a;
    layer1_outputs(12409) <= not (a xor b);
    layer1_outputs(12410) <= not a or b;
    layer1_outputs(12411) <= a or b;
    layer1_outputs(12412) <= not b or a;
    layer1_outputs(12413) <= not a;
    layer1_outputs(12414) <= not (a or b);
    layer1_outputs(12415) <= b and not a;
    layer1_outputs(12416) <= b and not a;
    layer1_outputs(12417) <= not a;
    layer1_outputs(12418) <= a xor b;
    layer1_outputs(12419) <= not (a xor b);
    layer1_outputs(12420) <= a;
    layer1_outputs(12421) <= a;
    layer1_outputs(12422) <= a and b;
    layer1_outputs(12423) <= not (a xor b);
    layer1_outputs(12424) <= a;
    layer1_outputs(12425) <= a and b;
    layer1_outputs(12426) <= not a;
    layer1_outputs(12427) <= not a;
    layer1_outputs(12428) <= not a or b;
    layer1_outputs(12429) <= b;
    layer1_outputs(12430) <= not b;
    layer1_outputs(12431) <= not (a and b);
    layer1_outputs(12432) <= a or b;
    layer1_outputs(12433) <= not (a or b);
    layer1_outputs(12434) <= not a;
    layer1_outputs(12435) <= a;
    layer1_outputs(12436) <= not a or b;
    layer1_outputs(12437) <= a and b;
    layer1_outputs(12438) <= a;
    layer1_outputs(12439) <= a or b;
    layer1_outputs(12440) <= not a or b;
    layer1_outputs(12441) <= b and not a;
    layer1_outputs(12442) <= not b;
    layer1_outputs(12443) <= a;
    layer1_outputs(12444) <= a or b;
    layer1_outputs(12445) <= not (a or b);
    layer1_outputs(12446) <= a or b;
    layer1_outputs(12447) <= not b;
    layer1_outputs(12448) <= not (a xor b);
    layer1_outputs(12449) <= not (a and b);
    layer1_outputs(12450) <= b;
    layer1_outputs(12451) <= a xor b;
    layer1_outputs(12452) <= a and not b;
    layer1_outputs(12453) <= not b or a;
    layer1_outputs(12454) <= a;
    layer1_outputs(12455) <= a xor b;
    layer1_outputs(12456) <= not b;
    layer1_outputs(12457) <= not (a xor b);
    layer1_outputs(12458) <= a and b;
    layer1_outputs(12459) <= not b;
    layer1_outputs(12460) <= b and not a;
    layer1_outputs(12461) <= a;
    layer1_outputs(12462) <= not a;
    layer1_outputs(12463) <= not b or a;
    layer1_outputs(12464) <= not a or b;
    layer1_outputs(12465) <= not (a xor b);
    layer1_outputs(12466) <= b;
    layer1_outputs(12467) <= not a or b;
    layer1_outputs(12468) <= not (a xor b);
    layer1_outputs(12469) <= a xor b;
    layer1_outputs(12470) <= not (a xor b);
    layer1_outputs(12471) <= a or b;
    layer1_outputs(12472) <= a;
    layer1_outputs(12473) <= not b;
    layer1_outputs(12474) <= not (a or b);
    layer1_outputs(12475) <= a or b;
    layer1_outputs(12476) <= b;
    layer1_outputs(12477) <= not (a or b);
    layer1_outputs(12478) <= a or b;
    layer1_outputs(12479) <= not a or b;
    layer1_outputs(12480) <= not (a xor b);
    layer1_outputs(12481) <= not b or a;
    layer1_outputs(12482) <= b and not a;
    layer1_outputs(12483) <= not (a or b);
    layer1_outputs(12484) <= a xor b;
    layer1_outputs(12485) <= b;
    layer1_outputs(12486) <= a;
    layer1_outputs(12487) <= b;
    layer1_outputs(12488) <= a and b;
    layer1_outputs(12489) <= a xor b;
    layer1_outputs(12490) <= a;
    layer1_outputs(12491) <= a;
    layer1_outputs(12492) <= 1'b1;
    layer1_outputs(12493) <= a;
    layer1_outputs(12494) <= not (a xor b);
    layer1_outputs(12495) <= a and b;
    layer1_outputs(12496) <= not a or b;
    layer1_outputs(12497) <= not (a xor b);
    layer1_outputs(12498) <= a or b;
    layer1_outputs(12499) <= a xor b;
    layer1_outputs(12500) <= not b;
    layer1_outputs(12501) <= not b or a;
    layer1_outputs(12502) <= a or b;
    layer1_outputs(12503) <= not b;
    layer1_outputs(12504) <= a and b;
    layer1_outputs(12505) <= not (a xor b);
    layer1_outputs(12506) <= not a;
    layer1_outputs(12507) <= not b;
    layer1_outputs(12508) <= not b or a;
    layer1_outputs(12509) <= not a or b;
    layer1_outputs(12510) <= a;
    layer1_outputs(12511) <= not b or a;
    layer1_outputs(12512) <= not (a or b);
    layer1_outputs(12513) <= not a or b;
    layer1_outputs(12514) <= a and b;
    layer1_outputs(12515) <= a;
    layer1_outputs(12516) <= a and not b;
    layer1_outputs(12517) <= b and not a;
    layer1_outputs(12518) <= b;
    layer1_outputs(12519) <= not b;
    layer1_outputs(12520) <= a and b;
    layer1_outputs(12521) <= a;
    layer1_outputs(12522) <= not b;
    layer1_outputs(12523) <= not a or b;
    layer1_outputs(12524) <= a and b;
    layer1_outputs(12525) <= not (a xor b);
    layer1_outputs(12526) <= not a;
    layer1_outputs(12527) <= 1'b0;
    layer1_outputs(12528) <= not b or a;
    layer1_outputs(12529) <= not (a xor b);
    layer1_outputs(12530) <= not a or b;
    layer1_outputs(12531) <= not a;
    layer1_outputs(12532) <= a;
    layer1_outputs(12533) <= b and not a;
    layer1_outputs(12534) <= not a or b;
    layer1_outputs(12535) <= not b;
    layer1_outputs(12536) <= not (a or b);
    layer1_outputs(12537) <= not (a and b);
    layer1_outputs(12538) <= a xor b;
    layer1_outputs(12539) <= a and b;
    layer1_outputs(12540) <= not b;
    layer1_outputs(12541) <= not a or b;
    layer1_outputs(12542) <= b and not a;
    layer1_outputs(12543) <= not (a and b);
    layer1_outputs(12544) <= not (a xor b);
    layer1_outputs(12545) <= a;
    layer1_outputs(12546) <= a and not b;
    layer1_outputs(12547) <= not a;
    layer1_outputs(12548) <= a and not b;
    layer1_outputs(12549) <= not a or b;
    layer1_outputs(12550) <= a xor b;
    layer1_outputs(12551) <= b and not a;
    layer1_outputs(12552) <= a xor b;
    layer1_outputs(12553) <= not (a xor b);
    layer1_outputs(12554) <= not (a xor b);
    layer1_outputs(12555) <= not (a or b);
    layer1_outputs(12556) <= not a;
    layer1_outputs(12557) <= not a or b;
    layer1_outputs(12558) <= not b;
    layer1_outputs(12559) <= b;
    layer1_outputs(12560) <= b;
    layer1_outputs(12561) <= not a;
    layer1_outputs(12562) <= not (a or b);
    layer1_outputs(12563) <= not a;
    layer1_outputs(12564) <= a;
    layer1_outputs(12565) <= not b;
    layer1_outputs(12566) <= a;
    layer1_outputs(12567) <= not b or a;
    layer1_outputs(12568) <= b and not a;
    layer1_outputs(12569) <= a and b;
    layer1_outputs(12570) <= not b or a;
    layer1_outputs(12571) <= a;
    layer1_outputs(12572) <= a;
    layer1_outputs(12573) <= a xor b;
    layer1_outputs(12574) <= not a or b;
    layer1_outputs(12575) <= b;
    layer1_outputs(12576) <= not a;
    layer1_outputs(12577) <= not b;
    layer1_outputs(12578) <= b;
    layer1_outputs(12579) <= not (a xor b);
    layer1_outputs(12580) <= b and not a;
    layer1_outputs(12581) <= a or b;
    layer1_outputs(12582) <= a or b;
    layer1_outputs(12583) <= a;
    layer1_outputs(12584) <= not (a xor b);
    layer1_outputs(12585) <= a and not b;
    layer1_outputs(12586) <= a or b;
    layer1_outputs(12587) <= a;
    layer1_outputs(12588) <= a and not b;
    layer1_outputs(12589) <= not b or a;
    layer1_outputs(12590) <= a;
    layer1_outputs(12591) <= not b;
    layer1_outputs(12592) <= a xor b;
    layer1_outputs(12593) <= b;
    layer1_outputs(12594) <= not a;
    layer1_outputs(12595) <= b;
    layer1_outputs(12596) <= a or b;
    layer1_outputs(12597) <= not (a xor b);
    layer1_outputs(12598) <= not b or a;
    layer1_outputs(12599) <= not a;
    layer1_outputs(12600) <= b and not a;
    layer1_outputs(12601) <= b;
    layer1_outputs(12602) <= not a or b;
    layer1_outputs(12603) <= a and b;
    layer1_outputs(12604) <= 1'b1;
    layer1_outputs(12605) <= not a;
    layer1_outputs(12606) <= a and not b;
    layer1_outputs(12607) <= b;
    layer1_outputs(12608) <= not a;
    layer1_outputs(12609) <= a;
    layer1_outputs(12610) <= not a;
    layer1_outputs(12611) <= a;
    layer1_outputs(12612) <= a;
    layer1_outputs(12613) <= not (a xor b);
    layer1_outputs(12614) <= not a;
    layer1_outputs(12615) <= a and b;
    layer1_outputs(12616) <= not (a xor b);
    layer1_outputs(12617) <= b and not a;
    layer1_outputs(12618) <= not (a or b);
    layer1_outputs(12619) <= not b or a;
    layer1_outputs(12620) <= b and not a;
    layer1_outputs(12621) <= a and b;
    layer1_outputs(12622) <= not b or a;
    layer1_outputs(12623) <= not b;
    layer1_outputs(12624) <= not (a xor b);
    layer1_outputs(12625) <= not a or b;
    layer1_outputs(12626) <= a and b;
    layer1_outputs(12627) <= not a;
    layer1_outputs(12628) <= not (a xor b);
    layer1_outputs(12629) <= b;
    layer1_outputs(12630) <= not a;
    layer1_outputs(12631) <= not (a or b);
    layer1_outputs(12632) <= not b;
    layer1_outputs(12633) <= not b;
    layer1_outputs(12634) <= a or b;
    layer1_outputs(12635) <= not b;
    layer1_outputs(12636) <= not a or b;
    layer1_outputs(12637) <= a xor b;
    layer1_outputs(12638) <= not b or a;
    layer1_outputs(12639) <= a and not b;
    layer1_outputs(12640) <= not (a xor b);
    layer1_outputs(12641) <= not a or b;
    layer1_outputs(12642) <= not a or b;
    layer1_outputs(12643) <= not (a or b);
    layer1_outputs(12644) <= not a;
    layer1_outputs(12645) <= b and not a;
    layer1_outputs(12646) <= b;
    layer1_outputs(12647) <= b;
    layer1_outputs(12648) <= not (a or b);
    layer1_outputs(12649) <= 1'b0;
    layer1_outputs(12650) <= b and not a;
    layer1_outputs(12651) <= a and not b;
    layer1_outputs(12652) <= not (a or b);
    layer1_outputs(12653) <= a xor b;
    layer1_outputs(12654) <= not (a or b);
    layer1_outputs(12655) <= not (a and b);
    layer1_outputs(12656) <= b;
    layer1_outputs(12657) <= a and b;
    layer1_outputs(12658) <= not (a or b);
    layer1_outputs(12659) <= not a or b;
    layer1_outputs(12660) <= not a;
    layer1_outputs(12661) <= not a;
    layer1_outputs(12662) <= a;
    layer1_outputs(12663) <= not (a or b);
    layer1_outputs(12664) <= not (a or b);
    layer1_outputs(12665) <= not b or a;
    layer1_outputs(12666) <= b;
    layer1_outputs(12667) <= not (a xor b);
    layer1_outputs(12668) <= a and b;
    layer1_outputs(12669) <= not (a xor b);
    layer1_outputs(12670) <= a and not b;
    layer1_outputs(12671) <= a and not b;
    layer1_outputs(12672) <= a;
    layer1_outputs(12673) <= not (a xor b);
    layer1_outputs(12674) <= not (a or b);
    layer1_outputs(12675) <= b;
    layer1_outputs(12676) <= a;
    layer1_outputs(12677) <= not a;
    layer1_outputs(12678) <= not b;
    layer1_outputs(12679) <= b and not a;
    layer1_outputs(12680) <= not b;
    layer1_outputs(12681) <= a xor b;
    layer1_outputs(12682) <= b;
    layer1_outputs(12683) <= a;
    layer1_outputs(12684) <= a xor b;
    layer1_outputs(12685) <= not b;
    layer1_outputs(12686) <= not b;
    layer1_outputs(12687) <= not (a xor b);
    layer1_outputs(12688) <= b;
    layer1_outputs(12689) <= not (a or b);
    layer1_outputs(12690) <= a xor b;
    layer1_outputs(12691) <= a xor b;
    layer1_outputs(12692) <= not b;
    layer1_outputs(12693) <= not b or a;
    layer1_outputs(12694) <= a;
    layer1_outputs(12695) <= not b or a;
    layer1_outputs(12696) <= not (a or b);
    layer1_outputs(12697) <= a xor b;
    layer1_outputs(12698) <= a xor b;
    layer1_outputs(12699) <= a xor b;
    layer1_outputs(12700) <= not (a xor b);
    layer1_outputs(12701) <= b and not a;
    layer1_outputs(12702) <= not (a xor b);
    layer1_outputs(12703) <= a xor b;
    layer1_outputs(12704) <= not a;
    layer1_outputs(12705) <= b;
    layer1_outputs(12706) <= not (a xor b);
    layer1_outputs(12707) <= not b or a;
    layer1_outputs(12708) <= not b or a;
    layer1_outputs(12709) <= b;
    layer1_outputs(12710) <= a and b;
    layer1_outputs(12711) <= a and not b;
    layer1_outputs(12712) <= not (a xor b);
    layer1_outputs(12713) <= not b;
    layer1_outputs(12714) <= not a or b;
    layer1_outputs(12715) <= not (a and b);
    layer1_outputs(12716) <= a or b;
    layer1_outputs(12717) <= not (a xor b);
    layer1_outputs(12718) <= a xor b;
    layer1_outputs(12719) <= not (a xor b);
    layer1_outputs(12720) <= b;
    layer1_outputs(12721) <= b and not a;
    layer1_outputs(12722) <= not a;
    layer1_outputs(12723) <= a;
    layer1_outputs(12724) <= a and b;
    layer1_outputs(12725) <= a and b;
    layer1_outputs(12726) <= a;
    layer1_outputs(12727) <= a;
    layer1_outputs(12728) <= not (a and b);
    layer1_outputs(12729) <= not (a or b);
    layer1_outputs(12730) <= not (a xor b);
    layer1_outputs(12731) <= not a or b;
    layer1_outputs(12732) <= b;
    layer1_outputs(12733) <= not a or b;
    layer1_outputs(12734) <= a or b;
    layer1_outputs(12735) <= a or b;
    layer1_outputs(12736) <= not (a xor b);
    layer1_outputs(12737) <= a;
    layer1_outputs(12738) <= not (a and b);
    layer1_outputs(12739) <= 1'b0;
    layer1_outputs(12740) <= 1'b0;
    layer1_outputs(12741) <= a xor b;
    layer1_outputs(12742) <= not (a and b);
    layer1_outputs(12743) <= b;
    layer1_outputs(12744) <= not (a or b);
    layer1_outputs(12745) <= not b or a;
    layer1_outputs(12746) <= a xor b;
    layer1_outputs(12747) <= a and b;
    layer1_outputs(12748) <= not a;
    layer1_outputs(12749) <= not (a or b);
    layer1_outputs(12750) <= a;
    layer1_outputs(12751) <= not b;
    layer1_outputs(12752) <= b;
    layer1_outputs(12753) <= a or b;
    layer1_outputs(12754) <= not a;
    layer1_outputs(12755) <= a and b;
    layer1_outputs(12756) <= a and not b;
    layer1_outputs(12757) <= not (a and b);
    layer1_outputs(12758) <= not (a or b);
    layer1_outputs(12759) <= not (a or b);
    layer1_outputs(12760) <= not (a or b);
    layer1_outputs(12761) <= a xor b;
    layer1_outputs(12762) <= not (a xor b);
    layer1_outputs(12763) <= a and b;
    layer1_outputs(12764) <= a and b;
    layer1_outputs(12765) <= b;
    layer1_outputs(12766) <= not a;
    layer1_outputs(12767) <= not (a or b);
    layer1_outputs(12768) <= not (a or b);
    layer1_outputs(12769) <= not b;
    layer1_outputs(12770) <= not a or b;
    layer1_outputs(12771) <= a or b;
    layer1_outputs(12772) <= a and b;
    layer1_outputs(12773) <= not b or a;
    layer1_outputs(12774) <= not a or b;
    layer1_outputs(12775) <= not a;
    layer1_outputs(12776) <= a and not b;
    layer1_outputs(12777) <= not (a or b);
    layer1_outputs(12778) <= a or b;
    layer1_outputs(12779) <= not a or b;
    layer1_outputs(12780) <= not a or b;
    layer1_outputs(12781) <= a and not b;
    layer1_outputs(12782) <= not b or a;
    layer1_outputs(12783) <= a;
    layer1_outputs(12784) <= not b;
    layer1_outputs(12785) <= not (a and b);
    layer1_outputs(12786) <= a xor b;
    layer1_outputs(12787) <= a;
    layer1_outputs(12788) <= not (a xor b);
    layer1_outputs(12789) <= not a or b;
    layer1_outputs(12790) <= b and not a;
    layer1_outputs(12791) <= a and not b;
    layer1_outputs(12792) <= a and not b;
    layer1_outputs(12793) <= a;
    layer1_outputs(12794) <= a xor b;
    layer1_outputs(12795) <= a and not b;
    layer1_outputs(12796) <= not (a xor b);
    layer1_outputs(12797) <= not (a xor b);
    layer1_outputs(12798) <= a and b;
    layer1_outputs(12799) <= a xor b;
    layer2_outputs(0) <= b;
    layer2_outputs(1) <= not (a or b);
    layer2_outputs(2) <= a;
    layer2_outputs(3) <= a xor b;
    layer2_outputs(4) <= not a;
    layer2_outputs(5) <= not b;
    layer2_outputs(6) <= not a or b;
    layer2_outputs(7) <= not (a and b);
    layer2_outputs(8) <= b and not a;
    layer2_outputs(9) <= not (a and b);
    layer2_outputs(10) <= b;
    layer2_outputs(11) <= a xor b;
    layer2_outputs(12) <= not a;
    layer2_outputs(13) <= a;
    layer2_outputs(14) <= b;
    layer2_outputs(15) <= not (a xor b);
    layer2_outputs(16) <= not a or b;
    layer2_outputs(17) <= b;
    layer2_outputs(18) <= a or b;
    layer2_outputs(19) <= a;
    layer2_outputs(20) <= not (a xor b);
    layer2_outputs(21) <= a;
    layer2_outputs(22) <= not a;
    layer2_outputs(23) <= a and b;
    layer2_outputs(24) <= not (a or b);
    layer2_outputs(25) <= a;
    layer2_outputs(26) <= not (a xor b);
    layer2_outputs(27) <= not a or b;
    layer2_outputs(28) <= a and b;
    layer2_outputs(29) <= not b or a;
    layer2_outputs(30) <= b and not a;
    layer2_outputs(31) <= not a;
    layer2_outputs(32) <= not a;
    layer2_outputs(33) <= not (a xor b);
    layer2_outputs(34) <= a xor b;
    layer2_outputs(35) <= not (a and b);
    layer2_outputs(36) <= a xor b;
    layer2_outputs(37) <= b;
    layer2_outputs(38) <= not (a or b);
    layer2_outputs(39) <= a and not b;
    layer2_outputs(40) <= b;
    layer2_outputs(41) <= a;
    layer2_outputs(42) <= a;
    layer2_outputs(43) <= not b;
    layer2_outputs(44) <= b;
    layer2_outputs(45) <= not b or a;
    layer2_outputs(46) <= a and not b;
    layer2_outputs(47) <= b;
    layer2_outputs(48) <= not (a and b);
    layer2_outputs(49) <= a;
    layer2_outputs(50) <= b;
    layer2_outputs(51) <= a xor b;
    layer2_outputs(52) <= 1'b1;
    layer2_outputs(53) <= not (a and b);
    layer2_outputs(54) <= not b or a;
    layer2_outputs(55) <= a;
    layer2_outputs(56) <= not (a or b);
    layer2_outputs(57) <= a or b;
    layer2_outputs(58) <= a xor b;
    layer2_outputs(59) <= not b or a;
    layer2_outputs(60) <= a;
    layer2_outputs(61) <= not (a or b);
    layer2_outputs(62) <= a and b;
    layer2_outputs(63) <= not b;
    layer2_outputs(64) <= a and b;
    layer2_outputs(65) <= not (a xor b);
    layer2_outputs(66) <= not b;
    layer2_outputs(67) <= b;
    layer2_outputs(68) <= not b or a;
    layer2_outputs(69) <= a and b;
    layer2_outputs(70) <= b;
    layer2_outputs(71) <= a;
    layer2_outputs(72) <= a xor b;
    layer2_outputs(73) <= not (a xor b);
    layer2_outputs(74) <= not (a or b);
    layer2_outputs(75) <= b;
    layer2_outputs(76) <= not a or b;
    layer2_outputs(77) <= not b;
    layer2_outputs(78) <= a and b;
    layer2_outputs(79) <= not (a xor b);
    layer2_outputs(80) <= not a or b;
    layer2_outputs(81) <= b;
    layer2_outputs(82) <= not a or b;
    layer2_outputs(83) <= a xor b;
    layer2_outputs(84) <= not b;
    layer2_outputs(85) <= a and not b;
    layer2_outputs(86) <= not (a xor b);
    layer2_outputs(87) <= not b;
    layer2_outputs(88) <= not a or b;
    layer2_outputs(89) <= a and b;
    layer2_outputs(90) <= not b;
    layer2_outputs(91) <= a or b;
    layer2_outputs(92) <= b;
    layer2_outputs(93) <= not b or a;
    layer2_outputs(94) <= a and not b;
    layer2_outputs(95) <= a and not b;
    layer2_outputs(96) <= not b;
    layer2_outputs(97) <= b;
    layer2_outputs(98) <= a xor b;
    layer2_outputs(99) <= not b;
    layer2_outputs(100) <= not b;
    layer2_outputs(101) <= not (a and b);
    layer2_outputs(102) <= not (a xor b);
    layer2_outputs(103) <= a xor b;
    layer2_outputs(104) <= not b;
    layer2_outputs(105) <= a or b;
    layer2_outputs(106) <= not a;
    layer2_outputs(107) <= a and not b;
    layer2_outputs(108) <= not (a xor b);
    layer2_outputs(109) <= not a;
    layer2_outputs(110) <= not (a or b);
    layer2_outputs(111) <= not b;
    layer2_outputs(112) <= b;
    layer2_outputs(113) <= not a;
    layer2_outputs(114) <= not b;
    layer2_outputs(115) <= not b;
    layer2_outputs(116) <= not a;
    layer2_outputs(117) <= not a;
    layer2_outputs(118) <= a xor b;
    layer2_outputs(119) <= a;
    layer2_outputs(120) <= not b or a;
    layer2_outputs(121) <= a or b;
    layer2_outputs(122) <= not (a and b);
    layer2_outputs(123) <= a xor b;
    layer2_outputs(124) <= a;
    layer2_outputs(125) <= a;
    layer2_outputs(126) <= not (a xor b);
    layer2_outputs(127) <= not (a xor b);
    layer2_outputs(128) <= a and b;
    layer2_outputs(129) <= not (a and b);
    layer2_outputs(130) <= not b;
    layer2_outputs(131) <= a and b;
    layer2_outputs(132) <= b and not a;
    layer2_outputs(133) <= a and b;
    layer2_outputs(134) <= not b;
    layer2_outputs(135) <= not (a and b);
    layer2_outputs(136) <= a or b;
    layer2_outputs(137) <= not a or b;
    layer2_outputs(138) <= a and not b;
    layer2_outputs(139) <= a;
    layer2_outputs(140) <= not (a or b);
    layer2_outputs(141) <= a xor b;
    layer2_outputs(142) <= not b;
    layer2_outputs(143) <= a;
    layer2_outputs(144) <= a xor b;
    layer2_outputs(145) <= not b;
    layer2_outputs(146) <= not (a xor b);
    layer2_outputs(147) <= not b or a;
    layer2_outputs(148) <= not (a xor b);
    layer2_outputs(149) <= b and not a;
    layer2_outputs(150) <= not (a or b);
    layer2_outputs(151) <= not b or a;
    layer2_outputs(152) <= not b or a;
    layer2_outputs(153) <= not a;
    layer2_outputs(154) <= b;
    layer2_outputs(155) <= not b;
    layer2_outputs(156) <= b and not a;
    layer2_outputs(157) <= not (a or b);
    layer2_outputs(158) <= not b or a;
    layer2_outputs(159) <= not (a and b);
    layer2_outputs(160) <= not (a xor b);
    layer2_outputs(161) <= b and not a;
    layer2_outputs(162) <= not (a xor b);
    layer2_outputs(163) <= not (a xor b);
    layer2_outputs(164) <= not b or a;
    layer2_outputs(165) <= a xor b;
    layer2_outputs(166) <= a or b;
    layer2_outputs(167) <= not (a or b);
    layer2_outputs(168) <= a;
    layer2_outputs(169) <= not a or b;
    layer2_outputs(170) <= a;
    layer2_outputs(171) <= not a;
    layer2_outputs(172) <= not a;
    layer2_outputs(173) <= not b;
    layer2_outputs(174) <= a;
    layer2_outputs(175) <= not (a or b);
    layer2_outputs(176) <= a xor b;
    layer2_outputs(177) <= not a;
    layer2_outputs(178) <= not b;
    layer2_outputs(179) <= a xor b;
    layer2_outputs(180) <= not b or a;
    layer2_outputs(181) <= not a;
    layer2_outputs(182) <= not b;
    layer2_outputs(183) <= not b;
    layer2_outputs(184) <= not (a and b);
    layer2_outputs(185) <= b and not a;
    layer2_outputs(186) <= a and not b;
    layer2_outputs(187) <= not a;
    layer2_outputs(188) <= not (a and b);
    layer2_outputs(189) <= not (a xor b);
    layer2_outputs(190) <= not (a xor b);
    layer2_outputs(191) <= b and not a;
    layer2_outputs(192) <= not a;
    layer2_outputs(193) <= not (a and b);
    layer2_outputs(194) <= a;
    layer2_outputs(195) <= not (a xor b);
    layer2_outputs(196) <= not (a xor b);
    layer2_outputs(197) <= b;
    layer2_outputs(198) <= not a;
    layer2_outputs(199) <= not a or b;
    layer2_outputs(200) <= b and not a;
    layer2_outputs(201) <= not b;
    layer2_outputs(202) <= a and not b;
    layer2_outputs(203) <= not (a or b);
    layer2_outputs(204) <= not (a xor b);
    layer2_outputs(205) <= not b;
    layer2_outputs(206) <= a;
    layer2_outputs(207) <= not (a and b);
    layer2_outputs(208) <= a;
    layer2_outputs(209) <= a xor b;
    layer2_outputs(210) <= b and not a;
    layer2_outputs(211) <= not (a or b);
    layer2_outputs(212) <= not b or a;
    layer2_outputs(213) <= a;
    layer2_outputs(214) <= not (a xor b);
    layer2_outputs(215) <= not b;
    layer2_outputs(216) <= a and not b;
    layer2_outputs(217) <= a xor b;
    layer2_outputs(218) <= not b;
    layer2_outputs(219) <= not (a and b);
    layer2_outputs(220) <= a and not b;
    layer2_outputs(221) <= not a or b;
    layer2_outputs(222) <= a xor b;
    layer2_outputs(223) <= not (a xor b);
    layer2_outputs(224) <= not a;
    layer2_outputs(225) <= not a;
    layer2_outputs(226) <= b;
    layer2_outputs(227) <= not (a xor b);
    layer2_outputs(228) <= a;
    layer2_outputs(229) <= a;
    layer2_outputs(230) <= a;
    layer2_outputs(231) <= not a;
    layer2_outputs(232) <= not (a xor b);
    layer2_outputs(233) <= not (a xor b);
    layer2_outputs(234) <= not b;
    layer2_outputs(235) <= not b;
    layer2_outputs(236) <= not (a xor b);
    layer2_outputs(237) <= a or b;
    layer2_outputs(238) <= not b;
    layer2_outputs(239) <= not b;
    layer2_outputs(240) <= not a;
    layer2_outputs(241) <= not b or a;
    layer2_outputs(242) <= not (a xor b);
    layer2_outputs(243) <= 1'b1;
    layer2_outputs(244) <= not b;
    layer2_outputs(245) <= a;
    layer2_outputs(246) <= not a;
    layer2_outputs(247) <= a and not b;
    layer2_outputs(248) <= a and not b;
    layer2_outputs(249) <= a xor b;
    layer2_outputs(250) <= not (a xor b);
    layer2_outputs(251) <= a and b;
    layer2_outputs(252) <= a xor b;
    layer2_outputs(253) <= not a or b;
    layer2_outputs(254) <= b;
    layer2_outputs(255) <= a xor b;
    layer2_outputs(256) <= a xor b;
    layer2_outputs(257) <= not a;
    layer2_outputs(258) <= a;
    layer2_outputs(259) <= a xor b;
    layer2_outputs(260) <= b;
    layer2_outputs(261) <= b;
    layer2_outputs(262) <= a and b;
    layer2_outputs(263) <= not (a xor b);
    layer2_outputs(264) <= not a or b;
    layer2_outputs(265) <= a and not b;
    layer2_outputs(266) <= a;
    layer2_outputs(267) <= not b;
    layer2_outputs(268) <= not (a xor b);
    layer2_outputs(269) <= a and not b;
    layer2_outputs(270) <= a;
    layer2_outputs(271) <= not (a xor b);
    layer2_outputs(272) <= not b;
    layer2_outputs(273) <= not (a xor b);
    layer2_outputs(274) <= 1'b0;
    layer2_outputs(275) <= a;
    layer2_outputs(276) <= a xor b;
    layer2_outputs(277) <= b;
    layer2_outputs(278) <= not b or a;
    layer2_outputs(279) <= not (a or b);
    layer2_outputs(280) <= not b or a;
    layer2_outputs(281) <= not (a and b);
    layer2_outputs(282) <= not a;
    layer2_outputs(283) <= not b or a;
    layer2_outputs(284) <= not (a xor b);
    layer2_outputs(285) <= a or b;
    layer2_outputs(286) <= b;
    layer2_outputs(287) <= not b or a;
    layer2_outputs(288) <= not b or a;
    layer2_outputs(289) <= a;
    layer2_outputs(290) <= a;
    layer2_outputs(291) <= not (a xor b);
    layer2_outputs(292) <= b;
    layer2_outputs(293) <= not b;
    layer2_outputs(294) <= not (a or b);
    layer2_outputs(295) <= b;
    layer2_outputs(296) <= not (a or b);
    layer2_outputs(297) <= not a or b;
    layer2_outputs(298) <= a and not b;
    layer2_outputs(299) <= b;
    layer2_outputs(300) <= not a;
    layer2_outputs(301) <= not a or b;
    layer2_outputs(302) <= not (a and b);
    layer2_outputs(303) <= not b;
    layer2_outputs(304) <= not (a xor b);
    layer2_outputs(305) <= not (a or b);
    layer2_outputs(306) <= not a or b;
    layer2_outputs(307) <= b;
    layer2_outputs(308) <= not b or a;
    layer2_outputs(309) <= a;
    layer2_outputs(310) <= not (a xor b);
    layer2_outputs(311) <= not (a and b);
    layer2_outputs(312) <= a or b;
    layer2_outputs(313) <= not a or b;
    layer2_outputs(314) <= a;
    layer2_outputs(315) <= a and b;
    layer2_outputs(316) <= not a or b;
    layer2_outputs(317) <= a and b;
    layer2_outputs(318) <= not b;
    layer2_outputs(319) <= a;
    layer2_outputs(320) <= not b or a;
    layer2_outputs(321) <= not a;
    layer2_outputs(322) <= a;
    layer2_outputs(323) <= b and not a;
    layer2_outputs(324) <= a;
    layer2_outputs(325) <= not (a and b);
    layer2_outputs(326) <= not a;
    layer2_outputs(327) <= a xor b;
    layer2_outputs(328) <= a;
    layer2_outputs(329) <= not (a xor b);
    layer2_outputs(330) <= not a;
    layer2_outputs(331) <= not a;
    layer2_outputs(332) <= not b;
    layer2_outputs(333) <= a;
    layer2_outputs(334) <= not a or b;
    layer2_outputs(335) <= a and not b;
    layer2_outputs(336) <= b and not a;
    layer2_outputs(337) <= a xor b;
    layer2_outputs(338) <= b;
    layer2_outputs(339) <= not b;
    layer2_outputs(340) <= not a;
    layer2_outputs(341) <= a and b;
    layer2_outputs(342) <= not (a xor b);
    layer2_outputs(343) <= a and b;
    layer2_outputs(344) <= a and b;
    layer2_outputs(345) <= not b or a;
    layer2_outputs(346) <= b;
    layer2_outputs(347) <= not b or a;
    layer2_outputs(348) <= b;
    layer2_outputs(349) <= b;
    layer2_outputs(350) <= not (a and b);
    layer2_outputs(351) <= not b;
    layer2_outputs(352) <= a;
    layer2_outputs(353) <= a and not b;
    layer2_outputs(354) <= 1'b1;
    layer2_outputs(355) <= not b or a;
    layer2_outputs(356) <= not b;
    layer2_outputs(357) <= b and not a;
    layer2_outputs(358) <= not a;
    layer2_outputs(359) <= not a;
    layer2_outputs(360) <= a and b;
    layer2_outputs(361) <= b;
    layer2_outputs(362) <= a xor b;
    layer2_outputs(363) <= not a;
    layer2_outputs(364) <= not b;
    layer2_outputs(365) <= not b or a;
    layer2_outputs(366) <= a xor b;
    layer2_outputs(367) <= not a or b;
    layer2_outputs(368) <= a and b;
    layer2_outputs(369) <= a and not b;
    layer2_outputs(370) <= a;
    layer2_outputs(371) <= a or b;
    layer2_outputs(372) <= b;
    layer2_outputs(373) <= b;
    layer2_outputs(374) <= not (a xor b);
    layer2_outputs(375) <= not b;
    layer2_outputs(376) <= a xor b;
    layer2_outputs(377) <= not a or b;
    layer2_outputs(378) <= not (a or b);
    layer2_outputs(379) <= b and not a;
    layer2_outputs(380) <= not b;
    layer2_outputs(381) <= a;
    layer2_outputs(382) <= a;
    layer2_outputs(383) <= b and not a;
    layer2_outputs(384) <= a and b;
    layer2_outputs(385) <= not b;
    layer2_outputs(386) <= not b;
    layer2_outputs(387) <= a xor b;
    layer2_outputs(388) <= a and not b;
    layer2_outputs(389) <= not b;
    layer2_outputs(390) <= b and not a;
    layer2_outputs(391) <= not b;
    layer2_outputs(392) <= a;
    layer2_outputs(393) <= not a;
    layer2_outputs(394) <= not (a xor b);
    layer2_outputs(395) <= not b;
    layer2_outputs(396) <= not (a or b);
    layer2_outputs(397) <= not (a xor b);
    layer2_outputs(398) <= a and not b;
    layer2_outputs(399) <= not b;
    layer2_outputs(400) <= a;
    layer2_outputs(401) <= not a;
    layer2_outputs(402) <= b and not a;
    layer2_outputs(403) <= not a;
    layer2_outputs(404) <= not (a xor b);
    layer2_outputs(405) <= not a or b;
    layer2_outputs(406) <= b and not a;
    layer2_outputs(407) <= not (a or b);
    layer2_outputs(408) <= not (a or b);
    layer2_outputs(409) <= b and not a;
    layer2_outputs(410) <= not b;
    layer2_outputs(411) <= a;
    layer2_outputs(412) <= not (a or b);
    layer2_outputs(413) <= b;
    layer2_outputs(414) <= b;
    layer2_outputs(415) <= not b;
    layer2_outputs(416) <= a and b;
    layer2_outputs(417) <= not (a xor b);
    layer2_outputs(418) <= b;
    layer2_outputs(419) <= not a or b;
    layer2_outputs(420) <= a;
    layer2_outputs(421) <= a;
    layer2_outputs(422) <= a or b;
    layer2_outputs(423) <= not a;
    layer2_outputs(424) <= not b;
    layer2_outputs(425) <= not a;
    layer2_outputs(426) <= not (a xor b);
    layer2_outputs(427) <= b and not a;
    layer2_outputs(428) <= not b;
    layer2_outputs(429) <= a and b;
    layer2_outputs(430) <= a xor b;
    layer2_outputs(431) <= not a or b;
    layer2_outputs(432) <= not a or b;
    layer2_outputs(433) <= b and not a;
    layer2_outputs(434) <= a or b;
    layer2_outputs(435) <= not b;
    layer2_outputs(436) <= a;
    layer2_outputs(437) <= a;
    layer2_outputs(438) <= a xor b;
    layer2_outputs(439) <= a xor b;
    layer2_outputs(440) <= not (a xor b);
    layer2_outputs(441) <= not (a and b);
    layer2_outputs(442) <= b;
    layer2_outputs(443) <= not (a or b);
    layer2_outputs(444) <= not a;
    layer2_outputs(445) <= a or b;
    layer2_outputs(446) <= a and not b;
    layer2_outputs(447) <= a or b;
    layer2_outputs(448) <= not (a xor b);
    layer2_outputs(449) <= 1'b1;
    layer2_outputs(450) <= b;
    layer2_outputs(451) <= b;
    layer2_outputs(452) <= a and not b;
    layer2_outputs(453) <= a;
    layer2_outputs(454) <= a xor b;
    layer2_outputs(455) <= not (a and b);
    layer2_outputs(456) <= a and not b;
    layer2_outputs(457) <= not a;
    layer2_outputs(458) <= not a or b;
    layer2_outputs(459) <= not a;
    layer2_outputs(460) <= b and not a;
    layer2_outputs(461) <= a or b;
    layer2_outputs(462) <= not a;
    layer2_outputs(463) <= not b;
    layer2_outputs(464) <= a and not b;
    layer2_outputs(465) <= b and not a;
    layer2_outputs(466) <= not b;
    layer2_outputs(467) <= a xor b;
    layer2_outputs(468) <= b;
    layer2_outputs(469) <= not a;
    layer2_outputs(470) <= a;
    layer2_outputs(471) <= b;
    layer2_outputs(472) <= not b or a;
    layer2_outputs(473) <= not (a or b);
    layer2_outputs(474) <= not a or b;
    layer2_outputs(475) <= b;
    layer2_outputs(476) <= b;
    layer2_outputs(477) <= not (a or b);
    layer2_outputs(478) <= a;
    layer2_outputs(479) <= a;
    layer2_outputs(480) <= not a;
    layer2_outputs(481) <= b and not a;
    layer2_outputs(482) <= not b;
    layer2_outputs(483) <= a;
    layer2_outputs(484) <= not a;
    layer2_outputs(485) <= a or b;
    layer2_outputs(486) <= b;
    layer2_outputs(487) <= 1'b1;
    layer2_outputs(488) <= a or b;
    layer2_outputs(489) <= b;
    layer2_outputs(490) <= a xor b;
    layer2_outputs(491) <= not (a or b);
    layer2_outputs(492) <= a and b;
    layer2_outputs(493) <= 1'b1;
    layer2_outputs(494) <= not (a and b);
    layer2_outputs(495) <= a;
    layer2_outputs(496) <= not (a xor b);
    layer2_outputs(497) <= not (a xor b);
    layer2_outputs(498) <= a;
    layer2_outputs(499) <= a and b;
    layer2_outputs(500) <= b;
    layer2_outputs(501) <= not a;
    layer2_outputs(502) <= a or b;
    layer2_outputs(503) <= not (a or b);
    layer2_outputs(504) <= b;
    layer2_outputs(505) <= not a;
    layer2_outputs(506) <= a and not b;
    layer2_outputs(507) <= not a or b;
    layer2_outputs(508) <= not (a and b);
    layer2_outputs(509) <= a or b;
    layer2_outputs(510) <= a xor b;
    layer2_outputs(511) <= not a;
    layer2_outputs(512) <= a;
    layer2_outputs(513) <= 1'b0;
    layer2_outputs(514) <= not (a xor b);
    layer2_outputs(515) <= a xor b;
    layer2_outputs(516) <= b and not a;
    layer2_outputs(517) <= a xor b;
    layer2_outputs(518) <= not a;
    layer2_outputs(519) <= not b;
    layer2_outputs(520) <= a;
    layer2_outputs(521) <= not (a xor b);
    layer2_outputs(522) <= a;
    layer2_outputs(523) <= not b or a;
    layer2_outputs(524) <= a xor b;
    layer2_outputs(525) <= a xor b;
    layer2_outputs(526) <= not b or a;
    layer2_outputs(527) <= a and not b;
    layer2_outputs(528) <= a xor b;
    layer2_outputs(529) <= not b;
    layer2_outputs(530) <= b;
    layer2_outputs(531) <= b;
    layer2_outputs(532) <= not (a and b);
    layer2_outputs(533) <= 1'b1;
    layer2_outputs(534) <= a xor b;
    layer2_outputs(535) <= not (a xor b);
    layer2_outputs(536) <= not (a xor b);
    layer2_outputs(537) <= a;
    layer2_outputs(538) <= not a;
    layer2_outputs(539) <= not (a xor b);
    layer2_outputs(540) <= a;
    layer2_outputs(541) <= 1'b1;
    layer2_outputs(542) <= b;
    layer2_outputs(543) <= a xor b;
    layer2_outputs(544) <= b;
    layer2_outputs(545) <= not (a xor b);
    layer2_outputs(546) <= a;
    layer2_outputs(547) <= b;
    layer2_outputs(548) <= b;
    layer2_outputs(549) <= not (a or b);
    layer2_outputs(550) <= a;
    layer2_outputs(551) <= not b;
    layer2_outputs(552) <= not a;
    layer2_outputs(553) <= a xor b;
    layer2_outputs(554) <= b;
    layer2_outputs(555) <= not a or b;
    layer2_outputs(556) <= not b or a;
    layer2_outputs(557) <= b;
    layer2_outputs(558) <= a;
    layer2_outputs(559) <= not a;
    layer2_outputs(560) <= not a;
    layer2_outputs(561) <= a;
    layer2_outputs(562) <= not a or b;
    layer2_outputs(563) <= b;
    layer2_outputs(564) <= not b or a;
    layer2_outputs(565) <= not b;
    layer2_outputs(566) <= not (a xor b);
    layer2_outputs(567) <= a xor b;
    layer2_outputs(568) <= not b;
    layer2_outputs(569) <= a xor b;
    layer2_outputs(570) <= a xor b;
    layer2_outputs(571) <= not a;
    layer2_outputs(572) <= b and not a;
    layer2_outputs(573) <= not b;
    layer2_outputs(574) <= not b;
    layer2_outputs(575) <= not (a and b);
    layer2_outputs(576) <= not a;
    layer2_outputs(577) <= b;
    layer2_outputs(578) <= not b;
    layer2_outputs(579) <= not b;
    layer2_outputs(580) <= a xor b;
    layer2_outputs(581) <= a;
    layer2_outputs(582) <= a;
    layer2_outputs(583) <= not a;
    layer2_outputs(584) <= not (a xor b);
    layer2_outputs(585) <= not a or b;
    layer2_outputs(586) <= a xor b;
    layer2_outputs(587) <= not a;
    layer2_outputs(588) <= a and not b;
    layer2_outputs(589) <= a and b;
    layer2_outputs(590) <= not a;
    layer2_outputs(591) <= a xor b;
    layer2_outputs(592) <= not a;
    layer2_outputs(593) <= not a or b;
    layer2_outputs(594) <= b;
    layer2_outputs(595) <= not (a xor b);
    layer2_outputs(596) <= a or b;
    layer2_outputs(597) <= a and not b;
    layer2_outputs(598) <= a xor b;
    layer2_outputs(599) <= b and not a;
    layer2_outputs(600) <= not (a or b);
    layer2_outputs(601) <= not b or a;
    layer2_outputs(602) <= a;
    layer2_outputs(603) <= a;
    layer2_outputs(604) <= not (a or b);
    layer2_outputs(605) <= not a or b;
    layer2_outputs(606) <= not b;
    layer2_outputs(607) <= not (a xor b);
    layer2_outputs(608) <= not (a and b);
    layer2_outputs(609) <= not a;
    layer2_outputs(610) <= a and not b;
    layer2_outputs(611) <= not b;
    layer2_outputs(612) <= a and b;
    layer2_outputs(613) <= b and not a;
    layer2_outputs(614) <= a or b;
    layer2_outputs(615) <= b;
    layer2_outputs(616) <= a or b;
    layer2_outputs(617) <= not b;
    layer2_outputs(618) <= b;
    layer2_outputs(619) <= a;
    layer2_outputs(620) <= not a;
    layer2_outputs(621) <= b and not a;
    layer2_outputs(622) <= a xor b;
    layer2_outputs(623) <= a and b;
    layer2_outputs(624) <= not b;
    layer2_outputs(625) <= b;
    layer2_outputs(626) <= a and b;
    layer2_outputs(627) <= not b;
    layer2_outputs(628) <= a;
    layer2_outputs(629) <= not b;
    layer2_outputs(630) <= not b;
    layer2_outputs(631) <= not (a and b);
    layer2_outputs(632) <= b;
    layer2_outputs(633) <= not a;
    layer2_outputs(634) <= b;
    layer2_outputs(635) <= a;
    layer2_outputs(636) <= not a;
    layer2_outputs(637) <= a xor b;
    layer2_outputs(638) <= not a;
    layer2_outputs(639) <= not b;
    layer2_outputs(640) <= a;
    layer2_outputs(641) <= not (a and b);
    layer2_outputs(642) <= not b or a;
    layer2_outputs(643) <= not (a xor b);
    layer2_outputs(644) <= a and not b;
    layer2_outputs(645) <= not (a or b);
    layer2_outputs(646) <= not b or a;
    layer2_outputs(647) <= b;
    layer2_outputs(648) <= a and b;
    layer2_outputs(649) <= 1'b0;
    layer2_outputs(650) <= not b;
    layer2_outputs(651) <= a xor b;
    layer2_outputs(652) <= 1'b1;
    layer2_outputs(653) <= not b;
    layer2_outputs(654) <= b;
    layer2_outputs(655) <= a and b;
    layer2_outputs(656) <= not b or a;
    layer2_outputs(657) <= not a;
    layer2_outputs(658) <= not (a xor b);
    layer2_outputs(659) <= a and not b;
    layer2_outputs(660) <= b and not a;
    layer2_outputs(661) <= not (a xor b);
    layer2_outputs(662) <= a xor b;
    layer2_outputs(663) <= not (a or b);
    layer2_outputs(664) <= a or b;
    layer2_outputs(665) <= not (a xor b);
    layer2_outputs(666) <= a and b;
    layer2_outputs(667) <= not b or a;
    layer2_outputs(668) <= a and not b;
    layer2_outputs(669) <= a;
    layer2_outputs(670) <= a;
    layer2_outputs(671) <= not (a or b);
    layer2_outputs(672) <= not (a xor b);
    layer2_outputs(673) <= not b or a;
    layer2_outputs(674) <= not a;
    layer2_outputs(675) <= a;
    layer2_outputs(676) <= a;
    layer2_outputs(677) <= b;
    layer2_outputs(678) <= a xor b;
    layer2_outputs(679) <= not b;
    layer2_outputs(680) <= a xor b;
    layer2_outputs(681) <= a and b;
    layer2_outputs(682) <= not a;
    layer2_outputs(683) <= not (a xor b);
    layer2_outputs(684) <= a xor b;
    layer2_outputs(685) <= not (a and b);
    layer2_outputs(686) <= not b;
    layer2_outputs(687) <= not b or a;
    layer2_outputs(688) <= a or b;
    layer2_outputs(689) <= not (a xor b);
    layer2_outputs(690) <= not a;
    layer2_outputs(691) <= a;
    layer2_outputs(692) <= b;
    layer2_outputs(693) <= not b;
    layer2_outputs(694) <= a and b;
    layer2_outputs(695) <= a xor b;
    layer2_outputs(696) <= a and not b;
    layer2_outputs(697) <= not a;
    layer2_outputs(698) <= not b or a;
    layer2_outputs(699) <= b;
    layer2_outputs(700) <= b;
    layer2_outputs(701) <= not a;
    layer2_outputs(702) <= not a;
    layer2_outputs(703) <= a;
    layer2_outputs(704) <= b;
    layer2_outputs(705) <= not a or b;
    layer2_outputs(706) <= not (a or b);
    layer2_outputs(707) <= a and b;
    layer2_outputs(708) <= not b;
    layer2_outputs(709) <= not a or b;
    layer2_outputs(710) <= not (a xor b);
    layer2_outputs(711) <= not (a xor b);
    layer2_outputs(712) <= b;
    layer2_outputs(713) <= not (a xor b);
    layer2_outputs(714) <= a and b;
    layer2_outputs(715) <= a or b;
    layer2_outputs(716) <= a and not b;
    layer2_outputs(717) <= a or b;
    layer2_outputs(718) <= a xor b;
    layer2_outputs(719) <= a or b;
    layer2_outputs(720) <= a xor b;
    layer2_outputs(721) <= not a;
    layer2_outputs(722) <= b;
    layer2_outputs(723) <= not a;
    layer2_outputs(724) <= a xor b;
    layer2_outputs(725) <= not (a or b);
    layer2_outputs(726) <= not (a xor b);
    layer2_outputs(727) <= not (a xor b);
    layer2_outputs(728) <= not b or a;
    layer2_outputs(729) <= not (a xor b);
    layer2_outputs(730) <= a;
    layer2_outputs(731) <= b;
    layer2_outputs(732) <= not b;
    layer2_outputs(733) <= not b or a;
    layer2_outputs(734) <= b;
    layer2_outputs(735) <= not a or b;
    layer2_outputs(736) <= not (a xor b);
    layer2_outputs(737) <= b;
    layer2_outputs(738) <= a xor b;
    layer2_outputs(739) <= not (a or b);
    layer2_outputs(740) <= not b or a;
    layer2_outputs(741) <= b;
    layer2_outputs(742) <= a or b;
    layer2_outputs(743) <= a;
    layer2_outputs(744) <= not b or a;
    layer2_outputs(745) <= a and b;
    layer2_outputs(746) <= not (a xor b);
    layer2_outputs(747) <= a and not b;
    layer2_outputs(748) <= a and b;
    layer2_outputs(749) <= a;
    layer2_outputs(750) <= not (a or b);
    layer2_outputs(751) <= not a;
    layer2_outputs(752) <= a and not b;
    layer2_outputs(753) <= not a;
    layer2_outputs(754) <= not a;
    layer2_outputs(755) <= not (a xor b);
    layer2_outputs(756) <= not b;
    layer2_outputs(757) <= a xor b;
    layer2_outputs(758) <= a;
    layer2_outputs(759) <= not a or b;
    layer2_outputs(760) <= a and not b;
    layer2_outputs(761) <= a and b;
    layer2_outputs(762) <= b;
    layer2_outputs(763) <= not (a xor b);
    layer2_outputs(764) <= b;
    layer2_outputs(765) <= a and b;
    layer2_outputs(766) <= not a;
    layer2_outputs(767) <= a and b;
    layer2_outputs(768) <= not a;
    layer2_outputs(769) <= not a or b;
    layer2_outputs(770) <= b and not a;
    layer2_outputs(771) <= not b;
    layer2_outputs(772) <= 1'b0;
    layer2_outputs(773) <= 1'b0;
    layer2_outputs(774) <= not b;
    layer2_outputs(775) <= not a;
    layer2_outputs(776) <= not b or a;
    layer2_outputs(777) <= a;
    layer2_outputs(778) <= a xor b;
    layer2_outputs(779) <= a or b;
    layer2_outputs(780) <= b;
    layer2_outputs(781) <= not (a xor b);
    layer2_outputs(782) <= b;
    layer2_outputs(783) <= a xor b;
    layer2_outputs(784) <= not (a xor b);
    layer2_outputs(785) <= b;
    layer2_outputs(786) <= a;
    layer2_outputs(787) <= not a or b;
    layer2_outputs(788) <= a xor b;
    layer2_outputs(789) <= not b;
    layer2_outputs(790) <= a;
    layer2_outputs(791) <= not b;
    layer2_outputs(792) <= a and not b;
    layer2_outputs(793) <= a xor b;
    layer2_outputs(794) <= a xor b;
    layer2_outputs(795) <= a xor b;
    layer2_outputs(796) <= not (a or b);
    layer2_outputs(797) <= not a;
    layer2_outputs(798) <= not b;
    layer2_outputs(799) <= a or b;
    layer2_outputs(800) <= a;
    layer2_outputs(801) <= a xor b;
    layer2_outputs(802) <= a and b;
    layer2_outputs(803) <= not b;
    layer2_outputs(804) <= not (a and b);
    layer2_outputs(805) <= a and b;
    layer2_outputs(806) <= b and not a;
    layer2_outputs(807) <= b;
    layer2_outputs(808) <= a and b;
    layer2_outputs(809) <= b;
    layer2_outputs(810) <= a;
    layer2_outputs(811) <= not b;
    layer2_outputs(812) <= a or b;
    layer2_outputs(813) <= a xor b;
    layer2_outputs(814) <= not a or b;
    layer2_outputs(815) <= a xor b;
    layer2_outputs(816) <= not b;
    layer2_outputs(817) <= a xor b;
    layer2_outputs(818) <= a;
    layer2_outputs(819) <= a and not b;
    layer2_outputs(820) <= b;
    layer2_outputs(821) <= b;
    layer2_outputs(822) <= b;
    layer2_outputs(823) <= b and not a;
    layer2_outputs(824) <= not b;
    layer2_outputs(825) <= not a;
    layer2_outputs(826) <= a xor b;
    layer2_outputs(827) <= b and not a;
    layer2_outputs(828) <= not b;
    layer2_outputs(829) <= b and not a;
    layer2_outputs(830) <= not a or b;
    layer2_outputs(831) <= a xor b;
    layer2_outputs(832) <= a and b;
    layer2_outputs(833) <= not b;
    layer2_outputs(834) <= not (a xor b);
    layer2_outputs(835) <= a;
    layer2_outputs(836) <= not (a and b);
    layer2_outputs(837) <= not (a or b);
    layer2_outputs(838) <= a and b;
    layer2_outputs(839) <= a;
    layer2_outputs(840) <= not (a xor b);
    layer2_outputs(841) <= a;
    layer2_outputs(842) <= not a;
    layer2_outputs(843) <= not (a and b);
    layer2_outputs(844) <= not b;
    layer2_outputs(845) <= a and b;
    layer2_outputs(846) <= not b;
    layer2_outputs(847) <= not a or b;
    layer2_outputs(848) <= not (a or b);
    layer2_outputs(849) <= b;
    layer2_outputs(850) <= not b or a;
    layer2_outputs(851) <= not (a xor b);
    layer2_outputs(852) <= b and not a;
    layer2_outputs(853) <= not b;
    layer2_outputs(854) <= not (a or b);
    layer2_outputs(855) <= a xor b;
    layer2_outputs(856) <= a;
    layer2_outputs(857) <= a xor b;
    layer2_outputs(858) <= not a;
    layer2_outputs(859) <= b;
    layer2_outputs(860) <= a;
    layer2_outputs(861) <= not (a xor b);
    layer2_outputs(862) <= not b or a;
    layer2_outputs(863) <= not a;
    layer2_outputs(864) <= not a or b;
    layer2_outputs(865) <= a;
    layer2_outputs(866) <= not b or a;
    layer2_outputs(867) <= a and not b;
    layer2_outputs(868) <= not b or a;
    layer2_outputs(869) <= b;
    layer2_outputs(870) <= not a;
    layer2_outputs(871) <= b;
    layer2_outputs(872) <= b;
    layer2_outputs(873) <= a xor b;
    layer2_outputs(874) <= not b;
    layer2_outputs(875) <= not b;
    layer2_outputs(876) <= a or b;
    layer2_outputs(877) <= a and not b;
    layer2_outputs(878) <= not (a xor b);
    layer2_outputs(879) <= not b;
    layer2_outputs(880) <= a xor b;
    layer2_outputs(881) <= b;
    layer2_outputs(882) <= a xor b;
    layer2_outputs(883) <= b and not a;
    layer2_outputs(884) <= not b;
    layer2_outputs(885) <= a;
    layer2_outputs(886) <= b;
    layer2_outputs(887) <= a xor b;
    layer2_outputs(888) <= not a;
    layer2_outputs(889) <= a xor b;
    layer2_outputs(890) <= a and b;
    layer2_outputs(891) <= not (a and b);
    layer2_outputs(892) <= a and not b;
    layer2_outputs(893) <= not b or a;
    layer2_outputs(894) <= a and b;
    layer2_outputs(895) <= b;
    layer2_outputs(896) <= a and not b;
    layer2_outputs(897) <= a and not b;
    layer2_outputs(898) <= not (a or b);
    layer2_outputs(899) <= a;
    layer2_outputs(900) <= b;
    layer2_outputs(901) <= not a;
    layer2_outputs(902) <= b;
    layer2_outputs(903) <= not b or a;
    layer2_outputs(904) <= not (a xor b);
    layer2_outputs(905) <= a;
    layer2_outputs(906) <= b;
    layer2_outputs(907) <= b;
    layer2_outputs(908) <= a;
    layer2_outputs(909) <= b;
    layer2_outputs(910) <= b and not a;
    layer2_outputs(911) <= a or b;
    layer2_outputs(912) <= not b or a;
    layer2_outputs(913) <= not a or b;
    layer2_outputs(914) <= a;
    layer2_outputs(915) <= not a;
    layer2_outputs(916) <= not a or b;
    layer2_outputs(917) <= not (a xor b);
    layer2_outputs(918) <= not (a xor b);
    layer2_outputs(919) <= a and b;
    layer2_outputs(920) <= not (a xor b);
    layer2_outputs(921) <= a;
    layer2_outputs(922) <= not b;
    layer2_outputs(923) <= a;
    layer2_outputs(924) <= a xor b;
    layer2_outputs(925) <= not a;
    layer2_outputs(926) <= a or b;
    layer2_outputs(927) <= 1'b1;
    layer2_outputs(928) <= b;
    layer2_outputs(929) <= not (a xor b);
    layer2_outputs(930) <= not (a or b);
    layer2_outputs(931) <= not a;
    layer2_outputs(932) <= not (a xor b);
    layer2_outputs(933) <= a;
    layer2_outputs(934) <= not b or a;
    layer2_outputs(935) <= not b;
    layer2_outputs(936) <= a and b;
    layer2_outputs(937) <= a xor b;
    layer2_outputs(938) <= not b;
    layer2_outputs(939) <= not b;
    layer2_outputs(940) <= a;
    layer2_outputs(941) <= not (a xor b);
    layer2_outputs(942) <= a xor b;
    layer2_outputs(943) <= a;
    layer2_outputs(944) <= not b;
    layer2_outputs(945) <= not (a and b);
    layer2_outputs(946) <= a and b;
    layer2_outputs(947) <= not a or b;
    layer2_outputs(948) <= not (a xor b);
    layer2_outputs(949) <= b and not a;
    layer2_outputs(950) <= not a or b;
    layer2_outputs(951) <= not (a or b);
    layer2_outputs(952) <= not a;
    layer2_outputs(953) <= not a;
    layer2_outputs(954) <= b and not a;
    layer2_outputs(955) <= not b or a;
    layer2_outputs(956) <= a;
    layer2_outputs(957) <= not a;
    layer2_outputs(958) <= not a or b;
    layer2_outputs(959) <= a;
    layer2_outputs(960) <= a xor b;
    layer2_outputs(961) <= not a;
    layer2_outputs(962) <= b;
    layer2_outputs(963) <= not b;
    layer2_outputs(964) <= a;
    layer2_outputs(965) <= not (a or b);
    layer2_outputs(966) <= not b;
    layer2_outputs(967) <= a;
    layer2_outputs(968) <= not b or a;
    layer2_outputs(969) <= a or b;
    layer2_outputs(970) <= not (a xor b);
    layer2_outputs(971) <= not b;
    layer2_outputs(972) <= not a;
    layer2_outputs(973) <= not a;
    layer2_outputs(974) <= b;
    layer2_outputs(975) <= a or b;
    layer2_outputs(976) <= not a;
    layer2_outputs(977) <= not b;
    layer2_outputs(978) <= b;
    layer2_outputs(979) <= b;
    layer2_outputs(980) <= not a;
    layer2_outputs(981) <= a xor b;
    layer2_outputs(982) <= not (a and b);
    layer2_outputs(983) <= not (a or b);
    layer2_outputs(984) <= not (a xor b);
    layer2_outputs(985) <= not b;
    layer2_outputs(986) <= not (a or b);
    layer2_outputs(987) <= not b;
    layer2_outputs(988) <= not b;
    layer2_outputs(989) <= a xor b;
    layer2_outputs(990) <= not (a xor b);
    layer2_outputs(991) <= not a;
    layer2_outputs(992) <= b and not a;
    layer2_outputs(993) <= a or b;
    layer2_outputs(994) <= b;
    layer2_outputs(995) <= not (a or b);
    layer2_outputs(996) <= b and not a;
    layer2_outputs(997) <= not (a xor b);
    layer2_outputs(998) <= a or b;
    layer2_outputs(999) <= a or b;
    layer2_outputs(1000) <= b and not a;
    layer2_outputs(1001) <= not (a xor b);
    layer2_outputs(1002) <= not (a or b);
    layer2_outputs(1003) <= a;
    layer2_outputs(1004) <= a xor b;
    layer2_outputs(1005) <= not (a xor b);
    layer2_outputs(1006) <= b;
    layer2_outputs(1007) <= a and b;
    layer2_outputs(1008) <= a or b;
    layer2_outputs(1009) <= not (a or b);
    layer2_outputs(1010) <= not a;
    layer2_outputs(1011) <= not b;
    layer2_outputs(1012) <= b and not a;
    layer2_outputs(1013) <= not a;
    layer2_outputs(1014) <= a and b;
    layer2_outputs(1015) <= a or b;
    layer2_outputs(1016) <= a or b;
    layer2_outputs(1017) <= not (a xor b);
    layer2_outputs(1018) <= a and b;
    layer2_outputs(1019) <= not a or b;
    layer2_outputs(1020) <= not b or a;
    layer2_outputs(1021) <= a or b;
    layer2_outputs(1022) <= a;
    layer2_outputs(1023) <= not (a or b);
    layer2_outputs(1024) <= a;
    layer2_outputs(1025) <= not a or b;
    layer2_outputs(1026) <= not b;
    layer2_outputs(1027) <= not (a xor b);
    layer2_outputs(1028) <= b;
    layer2_outputs(1029) <= b;
    layer2_outputs(1030) <= a;
    layer2_outputs(1031) <= not b;
    layer2_outputs(1032) <= a and not b;
    layer2_outputs(1033) <= not b or a;
    layer2_outputs(1034) <= b;
    layer2_outputs(1035) <= a and b;
    layer2_outputs(1036) <= not (a or b);
    layer2_outputs(1037) <= not (a xor b);
    layer2_outputs(1038) <= b;
    layer2_outputs(1039) <= b;
    layer2_outputs(1040) <= a;
    layer2_outputs(1041) <= not (a or b);
    layer2_outputs(1042) <= a;
    layer2_outputs(1043) <= a;
    layer2_outputs(1044) <= not b;
    layer2_outputs(1045) <= not (a xor b);
    layer2_outputs(1046) <= b;
    layer2_outputs(1047) <= b and not a;
    layer2_outputs(1048) <= not (a xor b);
    layer2_outputs(1049) <= not (a xor b);
    layer2_outputs(1050) <= not (a and b);
    layer2_outputs(1051) <= not b;
    layer2_outputs(1052) <= not a or b;
    layer2_outputs(1053) <= not b;
    layer2_outputs(1054) <= not (a and b);
    layer2_outputs(1055) <= a;
    layer2_outputs(1056) <= b;
    layer2_outputs(1057) <= not (a xor b);
    layer2_outputs(1058) <= b;
    layer2_outputs(1059) <= a and b;
    layer2_outputs(1060) <= not b;
    layer2_outputs(1061) <= a;
    layer2_outputs(1062) <= b and not a;
    layer2_outputs(1063) <= not a or b;
    layer2_outputs(1064) <= not b;
    layer2_outputs(1065) <= a or b;
    layer2_outputs(1066) <= not (a xor b);
    layer2_outputs(1067) <= not b;
    layer2_outputs(1068) <= a xor b;
    layer2_outputs(1069) <= not (a xor b);
    layer2_outputs(1070) <= not a or b;
    layer2_outputs(1071) <= not (a xor b);
    layer2_outputs(1072) <= a and not b;
    layer2_outputs(1073) <= b;
    layer2_outputs(1074) <= not b;
    layer2_outputs(1075) <= not (a xor b);
    layer2_outputs(1076) <= b and not a;
    layer2_outputs(1077) <= not (a and b);
    layer2_outputs(1078) <= not b;
    layer2_outputs(1079) <= b;
    layer2_outputs(1080) <= not b;
    layer2_outputs(1081) <= not (a xor b);
    layer2_outputs(1082) <= not (a xor b);
    layer2_outputs(1083) <= not (a xor b);
    layer2_outputs(1084) <= not (a xor b);
    layer2_outputs(1085) <= a;
    layer2_outputs(1086) <= not (a xor b);
    layer2_outputs(1087) <= not (a and b);
    layer2_outputs(1088) <= not a or b;
    layer2_outputs(1089) <= b;
    layer2_outputs(1090) <= a;
    layer2_outputs(1091) <= a xor b;
    layer2_outputs(1092) <= not (a xor b);
    layer2_outputs(1093) <= a or b;
    layer2_outputs(1094) <= not (a xor b);
    layer2_outputs(1095) <= b and not a;
    layer2_outputs(1096) <= a;
    layer2_outputs(1097) <= a xor b;
    layer2_outputs(1098) <= not a;
    layer2_outputs(1099) <= not a;
    layer2_outputs(1100) <= not a or b;
    layer2_outputs(1101) <= a or b;
    layer2_outputs(1102) <= b and not a;
    layer2_outputs(1103) <= not (a xor b);
    layer2_outputs(1104) <= not a;
    layer2_outputs(1105) <= b;
    layer2_outputs(1106) <= a or b;
    layer2_outputs(1107) <= not b or a;
    layer2_outputs(1108) <= 1'b0;
    layer2_outputs(1109) <= a or b;
    layer2_outputs(1110) <= a;
    layer2_outputs(1111) <= b and not a;
    layer2_outputs(1112) <= 1'b1;
    layer2_outputs(1113) <= a;
    layer2_outputs(1114) <= not (a or b);
    layer2_outputs(1115) <= not b;
    layer2_outputs(1116) <= b;
    layer2_outputs(1117) <= a;
    layer2_outputs(1118) <= not a or b;
    layer2_outputs(1119) <= not b;
    layer2_outputs(1120) <= not a;
    layer2_outputs(1121) <= a and b;
    layer2_outputs(1122) <= a or b;
    layer2_outputs(1123) <= not b;
    layer2_outputs(1124) <= not (a or b);
    layer2_outputs(1125) <= not a or b;
    layer2_outputs(1126) <= not b;
    layer2_outputs(1127) <= b;
    layer2_outputs(1128) <= a and b;
    layer2_outputs(1129) <= a xor b;
    layer2_outputs(1130) <= a;
    layer2_outputs(1131) <= a xor b;
    layer2_outputs(1132) <= not b;
    layer2_outputs(1133) <= not b or a;
    layer2_outputs(1134) <= a xor b;
    layer2_outputs(1135) <= a xor b;
    layer2_outputs(1136) <= not (a xor b);
    layer2_outputs(1137) <= not (a or b);
    layer2_outputs(1138) <= not (a or b);
    layer2_outputs(1139) <= a;
    layer2_outputs(1140) <= not b;
    layer2_outputs(1141) <= not a or b;
    layer2_outputs(1142) <= not (a xor b);
    layer2_outputs(1143) <= a or b;
    layer2_outputs(1144) <= not (a or b);
    layer2_outputs(1145) <= not b;
    layer2_outputs(1146) <= not b;
    layer2_outputs(1147) <= b;
    layer2_outputs(1148) <= not (a and b);
    layer2_outputs(1149) <= not a or b;
    layer2_outputs(1150) <= a or b;
    layer2_outputs(1151) <= b and not a;
    layer2_outputs(1152) <= not (a xor b);
    layer2_outputs(1153) <= not a or b;
    layer2_outputs(1154) <= a and b;
    layer2_outputs(1155) <= b and not a;
    layer2_outputs(1156) <= not (a and b);
    layer2_outputs(1157) <= a;
    layer2_outputs(1158) <= a;
    layer2_outputs(1159) <= a xor b;
    layer2_outputs(1160) <= not (a xor b);
    layer2_outputs(1161) <= not b;
    layer2_outputs(1162) <= b;
    layer2_outputs(1163) <= a and not b;
    layer2_outputs(1164) <= not a;
    layer2_outputs(1165) <= not a or b;
    layer2_outputs(1166) <= a;
    layer2_outputs(1167) <= not (a and b);
    layer2_outputs(1168) <= a;
    layer2_outputs(1169) <= a xor b;
    layer2_outputs(1170) <= not a;
    layer2_outputs(1171) <= not b;
    layer2_outputs(1172) <= a or b;
    layer2_outputs(1173) <= not (a and b);
    layer2_outputs(1174) <= a;
    layer2_outputs(1175) <= not (a and b);
    layer2_outputs(1176) <= a xor b;
    layer2_outputs(1177) <= a and b;
    layer2_outputs(1178) <= not b or a;
    layer2_outputs(1179) <= not a or b;
    layer2_outputs(1180) <= not (a or b);
    layer2_outputs(1181) <= not a or b;
    layer2_outputs(1182) <= a xor b;
    layer2_outputs(1183) <= b;
    layer2_outputs(1184) <= not b;
    layer2_outputs(1185) <= not a;
    layer2_outputs(1186) <= a and not b;
    layer2_outputs(1187) <= b;
    layer2_outputs(1188) <= a and not b;
    layer2_outputs(1189) <= a or b;
    layer2_outputs(1190) <= not b or a;
    layer2_outputs(1191) <= not b;
    layer2_outputs(1192) <= a xor b;
    layer2_outputs(1193) <= not a or b;
    layer2_outputs(1194) <= not (a and b);
    layer2_outputs(1195) <= not a;
    layer2_outputs(1196) <= b and not a;
    layer2_outputs(1197) <= not (a and b);
    layer2_outputs(1198) <= a;
    layer2_outputs(1199) <= a and not b;
    layer2_outputs(1200) <= b;
    layer2_outputs(1201) <= not a or b;
    layer2_outputs(1202) <= a;
    layer2_outputs(1203) <= not b;
    layer2_outputs(1204) <= a xor b;
    layer2_outputs(1205) <= not (a or b);
    layer2_outputs(1206) <= not (a and b);
    layer2_outputs(1207) <= a;
    layer2_outputs(1208) <= a xor b;
    layer2_outputs(1209) <= b and not a;
    layer2_outputs(1210) <= not a;
    layer2_outputs(1211) <= not b or a;
    layer2_outputs(1212) <= a;
    layer2_outputs(1213) <= a xor b;
    layer2_outputs(1214) <= not (a xor b);
    layer2_outputs(1215) <= a xor b;
    layer2_outputs(1216) <= not b;
    layer2_outputs(1217) <= not a;
    layer2_outputs(1218) <= a and not b;
    layer2_outputs(1219) <= b and not a;
    layer2_outputs(1220) <= a xor b;
    layer2_outputs(1221) <= a and not b;
    layer2_outputs(1222) <= a;
    layer2_outputs(1223) <= a xor b;
    layer2_outputs(1224) <= not a;
    layer2_outputs(1225) <= a xor b;
    layer2_outputs(1226) <= not a;
    layer2_outputs(1227) <= 1'b0;
    layer2_outputs(1228) <= not b;
    layer2_outputs(1229) <= not a;
    layer2_outputs(1230) <= a and not b;
    layer2_outputs(1231) <= a;
    layer2_outputs(1232) <= a or b;
    layer2_outputs(1233) <= a and b;
    layer2_outputs(1234) <= not (a xor b);
    layer2_outputs(1235) <= not b;
    layer2_outputs(1236) <= not b or a;
    layer2_outputs(1237) <= a and b;
    layer2_outputs(1238) <= a;
    layer2_outputs(1239) <= a;
    layer2_outputs(1240) <= b;
    layer2_outputs(1241) <= not b or a;
    layer2_outputs(1242) <= a or b;
    layer2_outputs(1243) <= a and not b;
    layer2_outputs(1244) <= a and b;
    layer2_outputs(1245) <= not (a xor b);
    layer2_outputs(1246) <= a;
    layer2_outputs(1247) <= a and not b;
    layer2_outputs(1248) <= a;
    layer2_outputs(1249) <= a and not b;
    layer2_outputs(1250) <= not a;
    layer2_outputs(1251) <= a;
    layer2_outputs(1252) <= not a;
    layer2_outputs(1253) <= not (a xor b);
    layer2_outputs(1254) <= not a;
    layer2_outputs(1255) <= a;
    layer2_outputs(1256) <= a xor b;
    layer2_outputs(1257) <= a xor b;
    layer2_outputs(1258) <= a;
    layer2_outputs(1259) <= not b or a;
    layer2_outputs(1260) <= a xor b;
    layer2_outputs(1261) <= not (a or b);
    layer2_outputs(1262) <= a or b;
    layer2_outputs(1263) <= a and b;
    layer2_outputs(1264) <= not b;
    layer2_outputs(1265) <= a or b;
    layer2_outputs(1266) <= b;
    layer2_outputs(1267) <= b;
    layer2_outputs(1268) <= a and not b;
    layer2_outputs(1269) <= not a;
    layer2_outputs(1270) <= a xor b;
    layer2_outputs(1271) <= a and not b;
    layer2_outputs(1272) <= b and not a;
    layer2_outputs(1273) <= b;
    layer2_outputs(1274) <= not a;
    layer2_outputs(1275) <= not b;
    layer2_outputs(1276) <= not b;
    layer2_outputs(1277) <= a xor b;
    layer2_outputs(1278) <= a or b;
    layer2_outputs(1279) <= not a;
    layer2_outputs(1280) <= not b;
    layer2_outputs(1281) <= b and not a;
    layer2_outputs(1282) <= not (a xor b);
    layer2_outputs(1283) <= not a;
    layer2_outputs(1284) <= a and not b;
    layer2_outputs(1285) <= b and not a;
    layer2_outputs(1286) <= b;
    layer2_outputs(1287) <= b;
    layer2_outputs(1288) <= not b;
    layer2_outputs(1289) <= b;
    layer2_outputs(1290) <= b;
    layer2_outputs(1291) <= not (a xor b);
    layer2_outputs(1292) <= not (a xor b);
    layer2_outputs(1293) <= not b;
    layer2_outputs(1294) <= not b;
    layer2_outputs(1295) <= b;
    layer2_outputs(1296) <= b and not a;
    layer2_outputs(1297) <= not (a xor b);
    layer2_outputs(1298) <= not b;
    layer2_outputs(1299) <= not b or a;
    layer2_outputs(1300) <= b;
    layer2_outputs(1301) <= not (a xor b);
    layer2_outputs(1302) <= not a;
    layer2_outputs(1303) <= not (a xor b);
    layer2_outputs(1304) <= not b;
    layer2_outputs(1305) <= not b;
    layer2_outputs(1306) <= not (a xor b);
    layer2_outputs(1307) <= a xor b;
    layer2_outputs(1308) <= not b or a;
    layer2_outputs(1309) <= not (a xor b);
    layer2_outputs(1310) <= not b;
    layer2_outputs(1311) <= not (a xor b);
    layer2_outputs(1312) <= a xor b;
    layer2_outputs(1313) <= a or b;
    layer2_outputs(1314) <= b;
    layer2_outputs(1315) <= not b or a;
    layer2_outputs(1316) <= b;
    layer2_outputs(1317) <= not (a xor b);
    layer2_outputs(1318) <= a and not b;
    layer2_outputs(1319) <= not b;
    layer2_outputs(1320) <= a and b;
    layer2_outputs(1321) <= a and not b;
    layer2_outputs(1322) <= a or b;
    layer2_outputs(1323) <= a;
    layer2_outputs(1324) <= a xor b;
    layer2_outputs(1325) <= a xor b;
    layer2_outputs(1326) <= not (a or b);
    layer2_outputs(1327) <= a;
    layer2_outputs(1328) <= b;
    layer2_outputs(1329) <= b;
    layer2_outputs(1330) <= not b;
    layer2_outputs(1331) <= a and b;
    layer2_outputs(1332) <= not (a and b);
    layer2_outputs(1333) <= not (a xor b);
    layer2_outputs(1334) <= not a;
    layer2_outputs(1335) <= a;
    layer2_outputs(1336) <= 1'b0;
    layer2_outputs(1337) <= not a or b;
    layer2_outputs(1338) <= not (a or b);
    layer2_outputs(1339) <= not a;
    layer2_outputs(1340) <= a and b;
    layer2_outputs(1341) <= a xor b;
    layer2_outputs(1342) <= not a;
    layer2_outputs(1343) <= a or b;
    layer2_outputs(1344) <= not a or b;
    layer2_outputs(1345) <= b;
    layer2_outputs(1346) <= not (a xor b);
    layer2_outputs(1347) <= not a or b;
    layer2_outputs(1348) <= a or b;
    layer2_outputs(1349) <= a xor b;
    layer2_outputs(1350) <= a xor b;
    layer2_outputs(1351) <= b;
    layer2_outputs(1352) <= b;
    layer2_outputs(1353) <= not a;
    layer2_outputs(1354) <= 1'b1;
    layer2_outputs(1355) <= not b;
    layer2_outputs(1356) <= a or b;
    layer2_outputs(1357) <= a;
    layer2_outputs(1358) <= b and not a;
    layer2_outputs(1359) <= not a;
    layer2_outputs(1360) <= a and b;
    layer2_outputs(1361) <= a and b;
    layer2_outputs(1362) <= a;
    layer2_outputs(1363) <= b and not a;
    layer2_outputs(1364) <= not b or a;
    layer2_outputs(1365) <= a or b;
    layer2_outputs(1366) <= not b or a;
    layer2_outputs(1367) <= not b or a;
    layer2_outputs(1368) <= not (a xor b);
    layer2_outputs(1369) <= a and b;
    layer2_outputs(1370) <= not (a xor b);
    layer2_outputs(1371) <= a or b;
    layer2_outputs(1372) <= a or b;
    layer2_outputs(1373) <= a xor b;
    layer2_outputs(1374) <= not b or a;
    layer2_outputs(1375) <= not (a and b);
    layer2_outputs(1376) <= not a or b;
    layer2_outputs(1377) <= a;
    layer2_outputs(1378) <= b;
    layer2_outputs(1379) <= a;
    layer2_outputs(1380) <= a;
    layer2_outputs(1381) <= a and b;
    layer2_outputs(1382) <= not (a xor b);
    layer2_outputs(1383) <= not a;
    layer2_outputs(1384) <= b;
    layer2_outputs(1385) <= b and not a;
    layer2_outputs(1386) <= a and b;
    layer2_outputs(1387) <= not b or a;
    layer2_outputs(1388) <= a or b;
    layer2_outputs(1389) <= a and not b;
    layer2_outputs(1390) <= not a or b;
    layer2_outputs(1391) <= not (a or b);
    layer2_outputs(1392) <= a;
    layer2_outputs(1393) <= not (a or b);
    layer2_outputs(1394) <= not (a xor b);
    layer2_outputs(1395) <= a or b;
    layer2_outputs(1396) <= not a or b;
    layer2_outputs(1397) <= a xor b;
    layer2_outputs(1398) <= a and b;
    layer2_outputs(1399) <= a;
    layer2_outputs(1400) <= a or b;
    layer2_outputs(1401) <= a or b;
    layer2_outputs(1402) <= b;
    layer2_outputs(1403) <= b;
    layer2_outputs(1404) <= not (a and b);
    layer2_outputs(1405) <= not b;
    layer2_outputs(1406) <= not b;
    layer2_outputs(1407) <= not a;
    layer2_outputs(1408) <= not (a xor b);
    layer2_outputs(1409) <= not a;
    layer2_outputs(1410) <= not b;
    layer2_outputs(1411) <= b;
    layer2_outputs(1412) <= a and b;
    layer2_outputs(1413) <= not b;
    layer2_outputs(1414) <= not a;
    layer2_outputs(1415) <= not a or b;
    layer2_outputs(1416) <= not (a or b);
    layer2_outputs(1417) <= not a or b;
    layer2_outputs(1418) <= a;
    layer2_outputs(1419) <= a;
    layer2_outputs(1420) <= not (a xor b);
    layer2_outputs(1421) <= not a or b;
    layer2_outputs(1422) <= a xor b;
    layer2_outputs(1423) <= b;
    layer2_outputs(1424) <= not a;
    layer2_outputs(1425) <= not a or b;
    layer2_outputs(1426) <= not b or a;
    layer2_outputs(1427) <= not b or a;
    layer2_outputs(1428) <= not a or b;
    layer2_outputs(1429) <= not a;
    layer2_outputs(1430) <= not (a or b);
    layer2_outputs(1431) <= not a or b;
    layer2_outputs(1432) <= a;
    layer2_outputs(1433) <= not a or b;
    layer2_outputs(1434) <= a;
    layer2_outputs(1435) <= not (a xor b);
    layer2_outputs(1436) <= not (a or b);
    layer2_outputs(1437) <= b and not a;
    layer2_outputs(1438) <= a xor b;
    layer2_outputs(1439) <= not a;
    layer2_outputs(1440) <= not b;
    layer2_outputs(1441) <= b;
    layer2_outputs(1442) <= a or b;
    layer2_outputs(1443) <= not (a xor b);
    layer2_outputs(1444) <= b;
    layer2_outputs(1445) <= not a;
    layer2_outputs(1446) <= not (a and b);
    layer2_outputs(1447) <= not (a xor b);
    layer2_outputs(1448) <= not (a and b);
    layer2_outputs(1449) <= a or b;
    layer2_outputs(1450) <= b and not a;
    layer2_outputs(1451) <= not (a or b);
    layer2_outputs(1452) <= a;
    layer2_outputs(1453) <= b;
    layer2_outputs(1454) <= a or b;
    layer2_outputs(1455) <= not (a or b);
    layer2_outputs(1456) <= not b;
    layer2_outputs(1457) <= not (a or b);
    layer2_outputs(1458) <= b;
    layer2_outputs(1459) <= not b or a;
    layer2_outputs(1460) <= a xor b;
    layer2_outputs(1461) <= a;
    layer2_outputs(1462) <= not (a and b);
    layer2_outputs(1463) <= a xor b;
    layer2_outputs(1464) <= a xor b;
    layer2_outputs(1465) <= a xor b;
    layer2_outputs(1466) <= b and not a;
    layer2_outputs(1467) <= a xor b;
    layer2_outputs(1468) <= a;
    layer2_outputs(1469) <= not (a xor b);
    layer2_outputs(1470) <= not (a xor b);
    layer2_outputs(1471) <= not (a or b);
    layer2_outputs(1472) <= a and not b;
    layer2_outputs(1473) <= not (a and b);
    layer2_outputs(1474) <= not b;
    layer2_outputs(1475) <= not (a or b);
    layer2_outputs(1476) <= b and not a;
    layer2_outputs(1477) <= not (a and b);
    layer2_outputs(1478) <= b;
    layer2_outputs(1479) <= not a or b;
    layer2_outputs(1480) <= a or b;
    layer2_outputs(1481) <= a;
    layer2_outputs(1482) <= not (a and b);
    layer2_outputs(1483) <= not (a xor b);
    layer2_outputs(1484) <= not (a and b);
    layer2_outputs(1485) <= not a or b;
    layer2_outputs(1486) <= b;
    layer2_outputs(1487) <= not (a xor b);
    layer2_outputs(1488) <= a and b;
    layer2_outputs(1489) <= a and b;
    layer2_outputs(1490) <= a;
    layer2_outputs(1491) <= a and b;
    layer2_outputs(1492) <= a and b;
    layer2_outputs(1493) <= not a or b;
    layer2_outputs(1494) <= not a;
    layer2_outputs(1495) <= not a;
    layer2_outputs(1496) <= b and not a;
    layer2_outputs(1497) <= not b;
    layer2_outputs(1498) <= not b;
    layer2_outputs(1499) <= not b or a;
    layer2_outputs(1500) <= b;
    layer2_outputs(1501) <= a;
    layer2_outputs(1502) <= a;
    layer2_outputs(1503) <= not (a xor b);
    layer2_outputs(1504) <= not b;
    layer2_outputs(1505) <= not (a or b);
    layer2_outputs(1506) <= not b;
    layer2_outputs(1507) <= not (a xor b);
    layer2_outputs(1508) <= not a;
    layer2_outputs(1509) <= not a;
    layer2_outputs(1510) <= not a or b;
    layer2_outputs(1511) <= a or b;
    layer2_outputs(1512) <= a and not b;
    layer2_outputs(1513) <= a or b;
    layer2_outputs(1514) <= a xor b;
    layer2_outputs(1515) <= a;
    layer2_outputs(1516) <= a;
    layer2_outputs(1517) <= not b;
    layer2_outputs(1518) <= not b or a;
    layer2_outputs(1519) <= a;
    layer2_outputs(1520) <= not a;
    layer2_outputs(1521) <= b;
    layer2_outputs(1522) <= b;
    layer2_outputs(1523) <= a xor b;
    layer2_outputs(1524) <= b;
    layer2_outputs(1525) <= not a or b;
    layer2_outputs(1526) <= not a;
    layer2_outputs(1527) <= a and not b;
    layer2_outputs(1528) <= not a;
    layer2_outputs(1529) <= not (a and b);
    layer2_outputs(1530) <= not a;
    layer2_outputs(1531) <= b;
    layer2_outputs(1532) <= b;
    layer2_outputs(1533) <= a xor b;
    layer2_outputs(1534) <= not a;
    layer2_outputs(1535) <= a and b;
    layer2_outputs(1536) <= not (a xor b);
    layer2_outputs(1537) <= not (a xor b);
    layer2_outputs(1538) <= not a;
    layer2_outputs(1539) <= a xor b;
    layer2_outputs(1540) <= not a;
    layer2_outputs(1541) <= b and not a;
    layer2_outputs(1542) <= a xor b;
    layer2_outputs(1543) <= b;
    layer2_outputs(1544) <= not (a xor b);
    layer2_outputs(1545) <= a and not b;
    layer2_outputs(1546) <= not (a or b);
    layer2_outputs(1547) <= not b or a;
    layer2_outputs(1548) <= a;
    layer2_outputs(1549) <= not b;
    layer2_outputs(1550) <= a or b;
    layer2_outputs(1551) <= a xor b;
    layer2_outputs(1552) <= not (a xor b);
    layer2_outputs(1553) <= not (a xor b);
    layer2_outputs(1554) <= a and b;
    layer2_outputs(1555) <= not b or a;
    layer2_outputs(1556) <= b;
    layer2_outputs(1557) <= a xor b;
    layer2_outputs(1558) <= b;
    layer2_outputs(1559) <= not a;
    layer2_outputs(1560) <= a xor b;
    layer2_outputs(1561) <= not (a xor b);
    layer2_outputs(1562) <= b and not a;
    layer2_outputs(1563) <= b;
    layer2_outputs(1564) <= a or b;
    layer2_outputs(1565) <= not (a and b);
    layer2_outputs(1566) <= b and not a;
    layer2_outputs(1567) <= not a or b;
    layer2_outputs(1568) <= not (a xor b);
    layer2_outputs(1569) <= not a or b;
    layer2_outputs(1570) <= a or b;
    layer2_outputs(1571) <= not a;
    layer2_outputs(1572) <= not a;
    layer2_outputs(1573) <= not (a xor b);
    layer2_outputs(1574) <= a xor b;
    layer2_outputs(1575) <= a and not b;
    layer2_outputs(1576) <= not b or a;
    layer2_outputs(1577) <= a and not b;
    layer2_outputs(1578) <= a and b;
    layer2_outputs(1579) <= not b;
    layer2_outputs(1580) <= b and not a;
    layer2_outputs(1581) <= not b;
    layer2_outputs(1582) <= a xor b;
    layer2_outputs(1583) <= a xor b;
    layer2_outputs(1584) <= not (a and b);
    layer2_outputs(1585) <= a xor b;
    layer2_outputs(1586) <= not b or a;
    layer2_outputs(1587) <= not (a and b);
    layer2_outputs(1588) <= a xor b;
    layer2_outputs(1589) <= a or b;
    layer2_outputs(1590) <= b;
    layer2_outputs(1591) <= a;
    layer2_outputs(1592) <= a;
    layer2_outputs(1593) <= not (a xor b);
    layer2_outputs(1594) <= a;
    layer2_outputs(1595) <= b;
    layer2_outputs(1596) <= a xor b;
    layer2_outputs(1597) <= b and not a;
    layer2_outputs(1598) <= a or b;
    layer2_outputs(1599) <= a or b;
    layer2_outputs(1600) <= b;
    layer2_outputs(1601) <= not b;
    layer2_outputs(1602) <= a xor b;
    layer2_outputs(1603) <= not (a xor b);
    layer2_outputs(1604) <= not b;
    layer2_outputs(1605) <= not a;
    layer2_outputs(1606) <= a;
    layer2_outputs(1607) <= not a;
    layer2_outputs(1608) <= not a;
    layer2_outputs(1609) <= a and b;
    layer2_outputs(1610) <= not (a xor b);
    layer2_outputs(1611) <= b;
    layer2_outputs(1612) <= not b or a;
    layer2_outputs(1613) <= a;
    layer2_outputs(1614) <= a;
    layer2_outputs(1615) <= not b or a;
    layer2_outputs(1616) <= b;
    layer2_outputs(1617) <= not a;
    layer2_outputs(1618) <= not a;
    layer2_outputs(1619) <= not a;
    layer2_outputs(1620) <= not (a xor b);
    layer2_outputs(1621) <= not b;
    layer2_outputs(1622) <= a xor b;
    layer2_outputs(1623) <= a;
    layer2_outputs(1624) <= not (a and b);
    layer2_outputs(1625) <= not (a or b);
    layer2_outputs(1626) <= not b;
    layer2_outputs(1627) <= b;
    layer2_outputs(1628) <= a and not b;
    layer2_outputs(1629) <= not b;
    layer2_outputs(1630) <= not (a and b);
    layer2_outputs(1631) <= not a;
    layer2_outputs(1632) <= not a;
    layer2_outputs(1633) <= not (a and b);
    layer2_outputs(1634) <= not a or b;
    layer2_outputs(1635) <= not b;
    layer2_outputs(1636) <= not a;
    layer2_outputs(1637) <= a xor b;
    layer2_outputs(1638) <= a and b;
    layer2_outputs(1639) <= not b;
    layer2_outputs(1640) <= not b;
    layer2_outputs(1641) <= not (a and b);
    layer2_outputs(1642) <= not b or a;
    layer2_outputs(1643) <= not (a or b);
    layer2_outputs(1644) <= not (a xor b);
    layer2_outputs(1645) <= a xor b;
    layer2_outputs(1646) <= not a;
    layer2_outputs(1647) <= b;
    layer2_outputs(1648) <= b and not a;
    layer2_outputs(1649) <= a xor b;
    layer2_outputs(1650) <= a;
    layer2_outputs(1651) <= b and not a;
    layer2_outputs(1652) <= not a;
    layer2_outputs(1653) <= a xor b;
    layer2_outputs(1654) <= not b or a;
    layer2_outputs(1655) <= a xor b;
    layer2_outputs(1656) <= not b or a;
    layer2_outputs(1657) <= a and not b;
    layer2_outputs(1658) <= a or b;
    layer2_outputs(1659) <= not a or b;
    layer2_outputs(1660) <= not a;
    layer2_outputs(1661) <= a or b;
    layer2_outputs(1662) <= not a;
    layer2_outputs(1663) <= a and not b;
    layer2_outputs(1664) <= not a;
    layer2_outputs(1665) <= a and b;
    layer2_outputs(1666) <= a xor b;
    layer2_outputs(1667) <= a xor b;
    layer2_outputs(1668) <= not a or b;
    layer2_outputs(1669) <= not a;
    layer2_outputs(1670) <= not b or a;
    layer2_outputs(1671) <= not (a xor b);
    layer2_outputs(1672) <= not b;
    layer2_outputs(1673) <= not b;
    layer2_outputs(1674) <= a xor b;
    layer2_outputs(1675) <= b and not a;
    layer2_outputs(1676) <= not (a xor b);
    layer2_outputs(1677) <= not b;
    layer2_outputs(1678) <= b;
    layer2_outputs(1679) <= not b or a;
    layer2_outputs(1680) <= not a or b;
    layer2_outputs(1681) <= not b or a;
    layer2_outputs(1682) <= b;
    layer2_outputs(1683) <= not a;
    layer2_outputs(1684) <= not a;
    layer2_outputs(1685) <= not b;
    layer2_outputs(1686) <= b;
    layer2_outputs(1687) <= 1'b1;
    layer2_outputs(1688) <= not a;
    layer2_outputs(1689) <= a xor b;
    layer2_outputs(1690) <= a or b;
    layer2_outputs(1691) <= not b;
    layer2_outputs(1692) <= not a or b;
    layer2_outputs(1693) <= a;
    layer2_outputs(1694) <= a;
    layer2_outputs(1695) <= a xor b;
    layer2_outputs(1696) <= not (a or b);
    layer2_outputs(1697) <= not b;
    layer2_outputs(1698) <= not b;
    layer2_outputs(1699) <= not b or a;
    layer2_outputs(1700) <= b and not a;
    layer2_outputs(1701) <= 1'b0;
    layer2_outputs(1702) <= b;
    layer2_outputs(1703) <= not a;
    layer2_outputs(1704) <= not b;
    layer2_outputs(1705) <= not b;
    layer2_outputs(1706) <= b;
    layer2_outputs(1707) <= a xor b;
    layer2_outputs(1708) <= not (a xor b);
    layer2_outputs(1709) <= a or b;
    layer2_outputs(1710) <= a or b;
    layer2_outputs(1711) <= not a;
    layer2_outputs(1712) <= a and b;
    layer2_outputs(1713) <= not a or b;
    layer2_outputs(1714) <= a;
    layer2_outputs(1715) <= not (a or b);
    layer2_outputs(1716) <= a and not b;
    layer2_outputs(1717) <= a xor b;
    layer2_outputs(1718) <= not a;
    layer2_outputs(1719) <= not a or b;
    layer2_outputs(1720) <= a xor b;
    layer2_outputs(1721) <= b;
    layer2_outputs(1722) <= a and b;
    layer2_outputs(1723) <= a xor b;
    layer2_outputs(1724) <= not b;
    layer2_outputs(1725) <= not b;
    layer2_outputs(1726) <= not (a xor b);
    layer2_outputs(1727) <= not a;
    layer2_outputs(1728) <= a xor b;
    layer2_outputs(1729) <= not (a xor b);
    layer2_outputs(1730) <= a xor b;
    layer2_outputs(1731) <= not (a or b);
    layer2_outputs(1732) <= a xor b;
    layer2_outputs(1733) <= not (a xor b);
    layer2_outputs(1734) <= not b or a;
    layer2_outputs(1735) <= not (a and b);
    layer2_outputs(1736) <= a xor b;
    layer2_outputs(1737) <= a;
    layer2_outputs(1738) <= a;
    layer2_outputs(1739) <= not (a xor b);
    layer2_outputs(1740) <= not (a or b);
    layer2_outputs(1741) <= not (a and b);
    layer2_outputs(1742) <= a and not b;
    layer2_outputs(1743) <= not b or a;
    layer2_outputs(1744) <= not a;
    layer2_outputs(1745) <= a xor b;
    layer2_outputs(1746) <= b;
    layer2_outputs(1747) <= a;
    layer2_outputs(1748) <= a xor b;
    layer2_outputs(1749) <= not b;
    layer2_outputs(1750) <= b;
    layer2_outputs(1751) <= b;
    layer2_outputs(1752) <= b;
    layer2_outputs(1753) <= not a or b;
    layer2_outputs(1754) <= b;
    layer2_outputs(1755) <= not b;
    layer2_outputs(1756) <= not b;
    layer2_outputs(1757) <= a xor b;
    layer2_outputs(1758) <= not (a xor b);
    layer2_outputs(1759) <= not (a xor b);
    layer2_outputs(1760) <= a or b;
    layer2_outputs(1761) <= not b;
    layer2_outputs(1762) <= a;
    layer2_outputs(1763) <= not b;
    layer2_outputs(1764) <= not (a xor b);
    layer2_outputs(1765) <= not a;
    layer2_outputs(1766) <= not a;
    layer2_outputs(1767) <= a xor b;
    layer2_outputs(1768) <= not (a xor b);
    layer2_outputs(1769) <= a xor b;
    layer2_outputs(1770) <= b;
    layer2_outputs(1771) <= b and not a;
    layer2_outputs(1772) <= not a or b;
    layer2_outputs(1773) <= not b;
    layer2_outputs(1774) <= not b or a;
    layer2_outputs(1775) <= a and not b;
    layer2_outputs(1776) <= a or b;
    layer2_outputs(1777) <= a xor b;
    layer2_outputs(1778) <= not (a and b);
    layer2_outputs(1779) <= a xor b;
    layer2_outputs(1780) <= a;
    layer2_outputs(1781) <= not a;
    layer2_outputs(1782) <= a xor b;
    layer2_outputs(1783) <= not (a and b);
    layer2_outputs(1784) <= not b or a;
    layer2_outputs(1785) <= not b;
    layer2_outputs(1786) <= a xor b;
    layer2_outputs(1787) <= a xor b;
    layer2_outputs(1788) <= not (a xor b);
    layer2_outputs(1789) <= b and not a;
    layer2_outputs(1790) <= a xor b;
    layer2_outputs(1791) <= a or b;
    layer2_outputs(1792) <= not (a or b);
    layer2_outputs(1793) <= not (a xor b);
    layer2_outputs(1794) <= not (a or b);
    layer2_outputs(1795) <= b and not a;
    layer2_outputs(1796) <= a;
    layer2_outputs(1797) <= not (a and b);
    layer2_outputs(1798) <= not b;
    layer2_outputs(1799) <= not (a xor b);
    layer2_outputs(1800) <= not a;
    layer2_outputs(1801) <= a or b;
    layer2_outputs(1802) <= a or b;
    layer2_outputs(1803) <= a;
    layer2_outputs(1804) <= not (a and b);
    layer2_outputs(1805) <= a xor b;
    layer2_outputs(1806) <= a xor b;
    layer2_outputs(1807) <= not b;
    layer2_outputs(1808) <= not a;
    layer2_outputs(1809) <= not a;
    layer2_outputs(1810) <= not (a xor b);
    layer2_outputs(1811) <= not b or a;
    layer2_outputs(1812) <= not a or b;
    layer2_outputs(1813) <= a or b;
    layer2_outputs(1814) <= b;
    layer2_outputs(1815) <= not (a xor b);
    layer2_outputs(1816) <= a and not b;
    layer2_outputs(1817) <= not b;
    layer2_outputs(1818) <= not a or b;
    layer2_outputs(1819) <= not b or a;
    layer2_outputs(1820) <= not b;
    layer2_outputs(1821) <= a xor b;
    layer2_outputs(1822) <= not b or a;
    layer2_outputs(1823) <= b;
    layer2_outputs(1824) <= not b or a;
    layer2_outputs(1825) <= a and not b;
    layer2_outputs(1826) <= not a;
    layer2_outputs(1827) <= not (a xor b);
    layer2_outputs(1828) <= not b;
    layer2_outputs(1829) <= a or b;
    layer2_outputs(1830) <= a or b;
    layer2_outputs(1831) <= a xor b;
    layer2_outputs(1832) <= not b or a;
    layer2_outputs(1833) <= not (a xor b);
    layer2_outputs(1834) <= b;
    layer2_outputs(1835) <= not b;
    layer2_outputs(1836) <= a and b;
    layer2_outputs(1837) <= not (a or b);
    layer2_outputs(1838) <= not a;
    layer2_outputs(1839) <= not (a xor b);
    layer2_outputs(1840) <= not (a or b);
    layer2_outputs(1841) <= b;
    layer2_outputs(1842) <= not (a or b);
    layer2_outputs(1843) <= not (a xor b);
    layer2_outputs(1844) <= a;
    layer2_outputs(1845) <= not (a xor b);
    layer2_outputs(1846) <= a and b;
    layer2_outputs(1847) <= not (a xor b);
    layer2_outputs(1848) <= a and not b;
    layer2_outputs(1849) <= not (a and b);
    layer2_outputs(1850) <= b and not a;
    layer2_outputs(1851) <= not (a xor b);
    layer2_outputs(1852) <= a and not b;
    layer2_outputs(1853) <= a and not b;
    layer2_outputs(1854) <= a or b;
    layer2_outputs(1855) <= a or b;
    layer2_outputs(1856) <= not (a xor b);
    layer2_outputs(1857) <= not (a or b);
    layer2_outputs(1858) <= a and not b;
    layer2_outputs(1859) <= b and not a;
    layer2_outputs(1860) <= not (a xor b);
    layer2_outputs(1861) <= not (a xor b);
    layer2_outputs(1862) <= not a;
    layer2_outputs(1863) <= not b;
    layer2_outputs(1864) <= b;
    layer2_outputs(1865) <= not b or a;
    layer2_outputs(1866) <= not b or a;
    layer2_outputs(1867) <= a and b;
    layer2_outputs(1868) <= not a;
    layer2_outputs(1869) <= a and b;
    layer2_outputs(1870) <= 1'b0;
    layer2_outputs(1871) <= a or b;
    layer2_outputs(1872) <= b;
    layer2_outputs(1873) <= not b or a;
    layer2_outputs(1874) <= not b;
    layer2_outputs(1875) <= not b;
    layer2_outputs(1876) <= not a or b;
    layer2_outputs(1877) <= a or b;
    layer2_outputs(1878) <= not b;
    layer2_outputs(1879) <= a;
    layer2_outputs(1880) <= not (a xor b);
    layer2_outputs(1881) <= not b;
    layer2_outputs(1882) <= a xor b;
    layer2_outputs(1883) <= not (a xor b);
    layer2_outputs(1884) <= a xor b;
    layer2_outputs(1885) <= a and not b;
    layer2_outputs(1886) <= not a;
    layer2_outputs(1887) <= not b;
    layer2_outputs(1888) <= not a or b;
    layer2_outputs(1889) <= not (a xor b);
    layer2_outputs(1890) <= a xor b;
    layer2_outputs(1891) <= not (a xor b);
    layer2_outputs(1892) <= a xor b;
    layer2_outputs(1893) <= b and not a;
    layer2_outputs(1894) <= not b;
    layer2_outputs(1895) <= a;
    layer2_outputs(1896) <= a xor b;
    layer2_outputs(1897) <= not (a or b);
    layer2_outputs(1898) <= not (a or b);
    layer2_outputs(1899) <= a and not b;
    layer2_outputs(1900) <= not b or a;
    layer2_outputs(1901) <= a xor b;
    layer2_outputs(1902) <= not a or b;
    layer2_outputs(1903) <= not a;
    layer2_outputs(1904) <= a and not b;
    layer2_outputs(1905) <= not b or a;
    layer2_outputs(1906) <= not b;
    layer2_outputs(1907) <= a xor b;
    layer2_outputs(1908) <= not a;
    layer2_outputs(1909) <= b and not a;
    layer2_outputs(1910) <= a and b;
    layer2_outputs(1911) <= a and not b;
    layer2_outputs(1912) <= a and b;
    layer2_outputs(1913) <= not b;
    layer2_outputs(1914) <= a;
    layer2_outputs(1915) <= not a;
    layer2_outputs(1916) <= b and not a;
    layer2_outputs(1917) <= b;
    layer2_outputs(1918) <= b;
    layer2_outputs(1919) <= not (a xor b);
    layer2_outputs(1920) <= not a or b;
    layer2_outputs(1921) <= not b or a;
    layer2_outputs(1922) <= not a;
    layer2_outputs(1923) <= not (a or b);
    layer2_outputs(1924) <= b;
    layer2_outputs(1925) <= not a or b;
    layer2_outputs(1926) <= not b or a;
    layer2_outputs(1927) <= not a;
    layer2_outputs(1928) <= a and not b;
    layer2_outputs(1929) <= a;
    layer2_outputs(1930) <= not (a and b);
    layer2_outputs(1931) <= not (a xor b);
    layer2_outputs(1932) <= not a or b;
    layer2_outputs(1933) <= not a;
    layer2_outputs(1934) <= not a;
    layer2_outputs(1935) <= not (a and b);
    layer2_outputs(1936) <= not a;
    layer2_outputs(1937) <= b;
    layer2_outputs(1938) <= not (a xor b);
    layer2_outputs(1939) <= b;
    layer2_outputs(1940) <= a xor b;
    layer2_outputs(1941) <= a xor b;
    layer2_outputs(1942) <= not (a or b);
    layer2_outputs(1943) <= b and not a;
    layer2_outputs(1944) <= not a or b;
    layer2_outputs(1945) <= b;
    layer2_outputs(1946) <= a and b;
    layer2_outputs(1947) <= not b or a;
    layer2_outputs(1948) <= not (a xor b);
    layer2_outputs(1949) <= b;
    layer2_outputs(1950) <= not (a or b);
    layer2_outputs(1951) <= not b or a;
    layer2_outputs(1952) <= not (a xor b);
    layer2_outputs(1953) <= not (a or b);
    layer2_outputs(1954) <= a xor b;
    layer2_outputs(1955) <= not (a or b);
    layer2_outputs(1956) <= b;
    layer2_outputs(1957) <= not (a xor b);
    layer2_outputs(1958) <= a xor b;
    layer2_outputs(1959) <= not (a or b);
    layer2_outputs(1960) <= a;
    layer2_outputs(1961) <= a;
    layer2_outputs(1962) <= a and not b;
    layer2_outputs(1963) <= a and b;
    layer2_outputs(1964) <= not (a and b);
    layer2_outputs(1965) <= not (a or b);
    layer2_outputs(1966) <= not (a and b);
    layer2_outputs(1967) <= a xor b;
    layer2_outputs(1968) <= a xor b;
    layer2_outputs(1969) <= not (a xor b);
    layer2_outputs(1970) <= a and not b;
    layer2_outputs(1971) <= b;
    layer2_outputs(1972) <= not (a or b);
    layer2_outputs(1973) <= not b;
    layer2_outputs(1974) <= a or b;
    layer2_outputs(1975) <= b;
    layer2_outputs(1976) <= a xor b;
    layer2_outputs(1977) <= not (a or b);
    layer2_outputs(1978) <= a;
    layer2_outputs(1979) <= not (a xor b);
    layer2_outputs(1980) <= not a;
    layer2_outputs(1981) <= a and not b;
    layer2_outputs(1982) <= not a;
    layer2_outputs(1983) <= b;
    layer2_outputs(1984) <= a and not b;
    layer2_outputs(1985) <= a and not b;
    layer2_outputs(1986) <= not b;
    layer2_outputs(1987) <= a;
    layer2_outputs(1988) <= not a or b;
    layer2_outputs(1989) <= not (a xor b);
    layer2_outputs(1990) <= a and b;
    layer2_outputs(1991) <= not a;
    layer2_outputs(1992) <= a;
    layer2_outputs(1993) <= not a;
    layer2_outputs(1994) <= a and not b;
    layer2_outputs(1995) <= not a or b;
    layer2_outputs(1996) <= not a or b;
    layer2_outputs(1997) <= a and b;
    layer2_outputs(1998) <= a or b;
    layer2_outputs(1999) <= not (a or b);
    layer2_outputs(2000) <= a xor b;
    layer2_outputs(2001) <= a xor b;
    layer2_outputs(2002) <= not b or a;
    layer2_outputs(2003) <= a;
    layer2_outputs(2004) <= a and b;
    layer2_outputs(2005) <= not b;
    layer2_outputs(2006) <= not b;
    layer2_outputs(2007) <= not (a xor b);
    layer2_outputs(2008) <= a xor b;
    layer2_outputs(2009) <= not a;
    layer2_outputs(2010) <= a or b;
    layer2_outputs(2011) <= a xor b;
    layer2_outputs(2012) <= not b;
    layer2_outputs(2013) <= a xor b;
    layer2_outputs(2014) <= not b;
    layer2_outputs(2015) <= a or b;
    layer2_outputs(2016) <= b and not a;
    layer2_outputs(2017) <= not (a xor b);
    layer2_outputs(2018) <= not (a and b);
    layer2_outputs(2019) <= a xor b;
    layer2_outputs(2020) <= a xor b;
    layer2_outputs(2021) <= not b;
    layer2_outputs(2022) <= not b;
    layer2_outputs(2023) <= not a or b;
    layer2_outputs(2024) <= not (a xor b);
    layer2_outputs(2025) <= b and not a;
    layer2_outputs(2026) <= not (a xor b);
    layer2_outputs(2027) <= b and not a;
    layer2_outputs(2028) <= not b;
    layer2_outputs(2029) <= not (a and b);
    layer2_outputs(2030) <= 1'b1;
    layer2_outputs(2031) <= a;
    layer2_outputs(2032) <= b and not a;
    layer2_outputs(2033) <= not a;
    layer2_outputs(2034) <= not b;
    layer2_outputs(2035) <= not b;
    layer2_outputs(2036) <= not a;
    layer2_outputs(2037) <= not (a or b);
    layer2_outputs(2038) <= not b;
    layer2_outputs(2039) <= a xor b;
    layer2_outputs(2040) <= b;
    layer2_outputs(2041) <= a and b;
    layer2_outputs(2042) <= not a;
    layer2_outputs(2043) <= a xor b;
    layer2_outputs(2044) <= b and not a;
    layer2_outputs(2045) <= not a or b;
    layer2_outputs(2046) <= not (a xor b);
    layer2_outputs(2047) <= a xor b;
    layer2_outputs(2048) <= a or b;
    layer2_outputs(2049) <= a xor b;
    layer2_outputs(2050) <= a xor b;
    layer2_outputs(2051) <= a and b;
    layer2_outputs(2052) <= not b or a;
    layer2_outputs(2053) <= b;
    layer2_outputs(2054) <= a xor b;
    layer2_outputs(2055) <= not b or a;
    layer2_outputs(2056) <= not (a xor b);
    layer2_outputs(2057) <= not a;
    layer2_outputs(2058) <= not b;
    layer2_outputs(2059) <= not a;
    layer2_outputs(2060) <= not (a xor b);
    layer2_outputs(2061) <= not b or a;
    layer2_outputs(2062) <= a or b;
    layer2_outputs(2063) <= a or b;
    layer2_outputs(2064) <= a xor b;
    layer2_outputs(2065) <= not (a and b);
    layer2_outputs(2066) <= b and not a;
    layer2_outputs(2067) <= a xor b;
    layer2_outputs(2068) <= not a or b;
    layer2_outputs(2069) <= a;
    layer2_outputs(2070) <= a;
    layer2_outputs(2071) <= a xor b;
    layer2_outputs(2072) <= 1'b1;
    layer2_outputs(2073) <= not b;
    layer2_outputs(2074) <= b;
    layer2_outputs(2075) <= a xor b;
    layer2_outputs(2076) <= not (a xor b);
    layer2_outputs(2077) <= a and b;
    layer2_outputs(2078) <= not (a xor b);
    layer2_outputs(2079) <= not (a xor b);
    layer2_outputs(2080) <= a xor b;
    layer2_outputs(2081) <= a;
    layer2_outputs(2082) <= a;
    layer2_outputs(2083) <= not (a xor b);
    layer2_outputs(2084) <= b;
    layer2_outputs(2085) <= a and not b;
    layer2_outputs(2086) <= b;
    layer2_outputs(2087) <= not (a or b);
    layer2_outputs(2088) <= not (a xor b);
    layer2_outputs(2089) <= a xor b;
    layer2_outputs(2090) <= a or b;
    layer2_outputs(2091) <= a and b;
    layer2_outputs(2092) <= not (a or b);
    layer2_outputs(2093) <= a and b;
    layer2_outputs(2094) <= not a;
    layer2_outputs(2095) <= a;
    layer2_outputs(2096) <= a;
    layer2_outputs(2097) <= a and b;
    layer2_outputs(2098) <= a or b;
    layer2_outputs(2099) <= not (a and b);
    layer2_outputs(2100) <= not (a xor b);
    layer2_outputs(2101) <= not (a and b);
    layer2_outputs(2102) <= not a;
    layer2_outputs(2103) <= a xor b;
    layer2_outputs(2104) <= not b or a;
    layer2_outputs(2105) <= not a or b;
    layer2_outputs(2106) <= not b;
    layer2_outputs(2107) <= not b;
    layer2_outputs(2108) <= not b;
    layer2_outputs(2109) <= not a;
    layer2_outputs(2110) <= b and not a;
    layer2_outputs(2111) <= not b;
    layer2_outputs(2112) <= b;
    layer2_outputs(2113) <= a and not b;
    layer2_outputs(2114) <= not a or b;
    layer2_outputs(2115) <= a xor b;
    layer2_outputs(2116) <= not a;
    layer2_outputs(2117) <= a;
    layer2_outputs(2118) <= b;
    layer2_outputs(2119) <= not a;
    layer2_outputs(2120) <= a and b;
    layer2_outputs(2121) <= not a or b;
    layer2_outputs(2122) <= not a;
    layer2_outputs(2123) <= not b or a;
    layer2_outputs(2124) <= a;
    layer2_outputs(2125) <= a and b;
    layer2_outputs(2126) <= not a;
    layer2_outputs(2127) <= a or b;
    layer2_outputs(2128) <= a;
    layer2_outputs(2129) <= not a or b;
    layer2_outputs(2130) <= not a;
    layer2_outputs(2131) <= not a or b;
    layer2_outputs(2132) <= not (a and b);
    layer2_outputs(2133) <= not b;
    layer2_outputs(2134) <= a or b;
    layer2_outputs(2135) <= not a;
    layer2_outputs(2136) <= a xor b;
    layer2_outputs(2137) <= not a or b;
    layer2_outputs(2138) <= b;
    layer2_outputs(2139) <= a and b;
    layer2_outputs(2140) <= a and not b;
    layer2_outputs(2141) <= 1'b0;
    layer2_outputs(2142) <= b and not a;
    layer2_outputs(2143) <= a;
    layer2_outputs(2144) <= not (a or b);
    layer2_outputs(2145) <= b;
    layer2_outputs(2146) <= a;
    layer2_outputs(2147) <= not (a xor b);
    layer2_outputs(2148) <= b and not a;
    layer2_outputs(2149) <= not (a xor b);
    layer2_outputs(2150) <= a xor b;
    layer2_outputs(2151) <= b;
    layer2_outputs(2152) <= not b;
    layer2_outputs(2153) <= not (a or b);
    layer2_outputs(2154) <= a xor b;
    layer2_outputs(2155) <= not (a xor b);
    layer2_outputs(2156) <= not b or a;
    layer2_outputs(2157) <= not b or a;
    layer2_outputs(2158) <= not (a xor b);
    layer2_outputs(2159) <= a and not b;
    layer2_outputs(2160) <= not (a and b);
    layer2_outputs(2161) <= b and not a;
    layer2_outputs(2162) <= not b or a;
    layer2_outputs(2163) <= a;
    layer2_outputs(2164) <= a;
    layer2_outputs(2165) <= b;
    layer2_outputs(2166) <= a xor b;
    layer2_outputs(2167) <= b;
    layer2_outputs(2168) <= not (a and b);
    layer2_outputs(2169) <= not b or a;
    layer2_outputs(2170) <= not a;
    layer2_outputs(2171) <= a and b;
    layer2_outputs(2172) <= not b;
    layer2_outputs(2173) <= not a;
    layer2_outputs(2174) <= b;
    layer2_outputs(2175) <= a xor b;
    layer2_outputs(2176) <= b and not a;
    layer2_outputs(2177) <= b and not a;
    layer2_outputs(2178) <= b;
    layer2_outputs(2179) <= not b or a;
    layer2_outputs(2180) <= not (a and b);
    layer2_outputs(2181) <= a or b;
    layer2_outputs(2182) <= a or b;
    layer2_outputs(2183) <= not b;
    layer2_outputs(2184) <= a or b;
    layer2_outputs(2185) <= not (a xor b);
    layer2_outputs(2186) <= not (a and b);
    layer2_outputs(2187) <= not (a or b);
    layer2_outputs(2188) <= b;
    layer2_outputs(2189) <= a and not b;
    layer2_outputs(2190) <= not b;
    layer2_outputs(2191) <= b and not a;
    layer2_outputs(2192) <= b and not a;
    layer2_outputs(2193) <= not (a and b);
    layer2_outputs(2194) <= b;
    layer2_outputs(2195) <= not b or a;
    layer2_outputs(2196) <= b and not a;
    layer2_outputs(2197) <= b and not a;
    layer2_outputs(2198) <= a and b;
    layer2_outputs(2199) <= not (a xor b);
    layer2_outputs(2200) <= a and b;
    layer2_outputs(2201) <= a xor b;
    layer2_outputs(2202) <= a and b;
    layer2_outputs(2203) <= not b or a;
    layer2_outputs(2204) <= not (a or b);
    layer2_outputs(2205) <= a;
    layer2_outputs(2206) <= not (a or b);
    layer2_outputs(2207) <= a;
    layer2_outputs(2208) <= not b;
    layer2_outputs(2209) <= a;
    layer2_outputs(2210) <= b and not a;
    layer2_outputs(2211) <= a xor b;
    layer2_outputs(2212) <= a and b;
    layer2_outputs(2213) <= not b;
    layer2_outputs(2214) <= not a or b;
    layer2_outputs(2215) <= not b or a;
    layer2_outputs(2216) <= b and not a;
    layer2_outputs(2217) <= not a;
    layer2_outputs(2218) <= not (a xor b);
    layer2_outputs(2219) <= a xor b;
    layer2_outputs(2220) <= b;
    layer2_outputs(2221) <= not (a and b);
    layer2_outputs(2222) <= a;
    layer2_outputs(2223) <= not a or b;
    layer2_outputs(2224) <= not b;
    layer2_outputs(2225) <= a;
    layer2_outputs(2226) <= a;
    layer2_outputs(2227) <= b;
    layer2_outputs(2228) <= not (a or b);
    layer2_outputs(2229) <= not b;
    layer2_outputs(2230) <= b;
    layer2_outputs(2231) <= not a or b;
    layer2_outputs(2232) <= not b;
    layer2_outputs(2233) <= not (a xor b);
    layer2_outputs(2234) <= b;
    layer2_outputs(2235) <= not (a xor b);
    layer2_outputs(2236) <= not a;
    layer2_outputs(2237) <= not (a and b);
    layer2_outputs(2238) <= b;
    layer2_outputs(2239) <= not (a or b);
    layer2_outputs(2240) <= not (a xor b);
    layer2_outputs(2241) <= not (a and b);
    layer2_outputs(2242) <= not (a xor b);
    layer2_outputs(2243) <= not (a and b);
    layer2_outputs(2244) <= a xor b;
    layer2_outputs(2245) <= not a or b;
    layer2_outputs(2246) <= a and b;
    layer2_outputs(2247) <= not a;
    layer2_outputs(2248) <= not a;
    layer2_outputs(2249) <= not b;
    layer2_outputs(2250) <= not b or a;
    layer2_outputs(2251) <= not (a xor b);
    layer2_outputs(2252) <= not a;
    layer2_outputs(2253) <= not b;
    layer2_outputs(2254) <= a;
    layer2_outputs(2255) <= b;
    layer2_outputs(2256) <= b and not a;
    layer2_outputs(2257) <= not (a xor b);
    layer2_outputs(2258) <= a and not b;
    layer2_outputs(2259) <= not b;
    layer2_outputs(2260) <= b;
    layer2_outputs(2261) <= not a or b;
    layer2_outputs(2262) <= not b;
    layer2_outputs(2263) <= not (a xor b);
    layer2_outputs(2264) <= not a;
    layer2_outputs(2265) <= not a or b;
    layer2_outputs(2266) <= not a;
    layer2_outputs(2267) <= b;
    layer2_outputs(2268) <= not b or a;
    layer2_outputs(2269) <= not b or a;
    layer2_outputs(2270) <= not b;
    layer2_outputs(2271) <= not (a and b);
    layer2_outputs(2272) <= not (a xor b);
    layer2_outputs(2273) <= a xor b;
    layer2_outputs(2274) <= a xor b;
    layer2_outputs(2275) <= not a;
    layer2_outputs(2276) <= not a or b;
    layer2_outputs(2277) <= not b or a;
    layer2_outputs(2278) <= a and not b;
    layer2_outputs(2279) <= a;
    layer2_outputs(2280) <= not (a and b);
    layer2_outputs(2281) <= a;
    layer2_outputs(2282) <= a and not b;
    layer2_outputs(2283) <= not b;
    layer2_outputs(2284) <= not (a or b);
    layer2_outputs(2285) <= not (a or b);
    layer2_outputs(2286) <= a or b;
    layer2_outputs(2287) <= a xor b;
    layer2_outputs(2288) <= a and not b;
    layer2_outputs(2289) <= not b;
    layer2_outputs(2290) <= not (a xor b);
    layer2_outputs(2291) <= not (a or b);
    layer2_outputs(2292) <= a and not b;
    layer2_outputs(2293) <= b and not a;
    layer2_outputs(2294) <= not (a and b);
    layer2_outputs(2295) <= a;
    layer2_outputs(2296) <= not b or a;
    layer2_outputs(2297) <= not (a and b);
    layer2_outputs(2298) <= b;
    layer2_outputs(2299) <= a;
    layer2_outputs(2300) <= a xor b;
    layer2_outputs(2301) <= b and not a;
    layer2_outputs(2302) <= a;
    layer2_outputs(2303) <= b;
    layer2_outputs(2304) <= b and not a;
    layer2_outputs(2305) <= not a;
    layer2_outputs(2306) <= not b;
    layer2_outputs(2307) <= not (a xor b);
    layer2_outputs(2308) <= a xor b;
    layer2_outputs(2309) <= b and not a;
    layer2_outputs(2310) <= a xor b;
    layer2_outputs(2311) <= a or b;
    layer2_outputs(2312) <= b;
    layer2_outputs(2313) <= not a or b;
    layer2_outputs(2314) <= not b;
    layer2_outputs(2315) <= not (a xor b);
    layer2_outputs(2316) <= not (a xor b);
    layer2_outputs(2317) <= b;
    layer2_outputs(2318) <= not (a or b);
    layer2_outputs(2319) <= not b;
    layer2_outputs(2320) <= not b;
    layer2_outputs(2321) <= not b;
    layer2_outputs(2322) <= b;
    layer2_outputs(2323) <= a and not b;
    layer2_outputs(2324) <= a xor b;
    layer2_outputs(2325) <= a and b;
    layer2_outputs(2326) <= not b or a;
    layer2_outputs(2327) <= a;
    layer2_outputs(2328) <= not (a or b);
    layer2_outputs(2329) <= a;
    layer2_outputs(2330) <= b;
    layer2_outputs(2331) <= a;
    layer2_outputs(2332) <= a;
    layer2_outputs(2333) <= a;
    layer2_outputs(2334) <= not b or a;
    layer2_outputs(2335) <= not a or b;
    layer2_outputs(2336) <= b;
    layer2_outputs(2337) <= not (a and b);
    layer2_outputs(2338) <= a xor b;
    layer2_outputs(2339) <= not (a and b);
    layer2_outputs(2340) <= not a;
    layer2_outputs(2341) <= not (a or b);
    layer2_outputs(2342) <= not (a and b);
    layer2_outputs(2343) <= b and not a;
    layer2_outputs(2344) <= not b;
    layer2_outputs(2345) <= a xor b;
    layer2_outputs(2346) <= a;
    layer2_outputs(2347) <= a and not b;
    layer2_outputs(2348) <= not (a xor b);
    layer2_outputs(2349) <= b;
    layer2_outputs(2350) <= not b;
    layer2_outputs(2351) <= a;
    layer2_outputs(2352) <= not (a xor b);
    layer2_outputs(2353) <= not b;
    layer2_outputs(2354) <= a xor b;
    layer2_outputs(2355) <= not b or a;
    layer2_outputs(2356) <= a or b;
    layer2_outputs(2357) <= a or b;
    layer2_outputs(2358) <= a;
    layer2_outputs(2359) <= b;
    layer2_outputs(2360) <= not a;
    layer2_outputs(2361) <= a and b;
    layer2_outputs(2362) <= not b or a;
    layer2_outputs(2363) <= 1'b1;
    layer2_outputs(2364) <= not (a or b);
    layer2_outputs(2365) <= not (a or b);
    layer2_outputs(2366) <= not b or a;
    layer2_outputs(2367) <= not a;
    layer2_outputs(2368) <= a xor b;
    layer2_outputs(2369) <= not a;
    layer2_outputs(2370) <= b and not a;
    layer2_outputs(2371) <= b;
    layer2_outputs(2372) <= b and not a;
    layer2_outputs(2373) <= a and b;
    layer2_outputs(2374) <= not (a xor b);
    layer2_outputs(2375) <= b;
    layer2_outputs(2376) <= a xor b;
    layer2_outputs(2377) <= a;
    layer2_outputs(2378) <= not b;
    layer2_outputs(2379) <= b;
    layer2_outputs(2380) <= not b;
    layer2_outputs(2381) <= not (a and b);
    layer2_outputs(2382) <= b;
    layer2_outputs(2383) <= a and b;
    layer2_outputs(2384) <= not a or b;
    layer2_outputs(2385) <= a and not b;
    layer2_outputs(2386) <= a xor b;
    layer2_outputs(2387) <= not a;
    layer2_outputs(2388) <= not a or b;
    layer2_outputs(2389) <= b;
    layer2_outputs(2390) <= not b or a;
    layer2_outputs(2391) <= b;
    layer2_outputs(2392) <= not (a and b);
    layer2_outputs(2393) <= not (a and b);
    layer2_outputs(2394) <= a xor b;
    layer2_outputs(2395) <= a;
    layer2_outputs(2396) <= not (a or b);
    layer2_outputs(2397) <= not b;
    layer2_outputs(2398) <= not (a xor b);
    layer2_outputs(2399) <= a;
    layer2_outputs(2400) <= a;
    layer2_outputs(2401) <= not (a xor b);
    layer2_outputs(2402) <= not (a and b);
    layer2_outputs(2403) <= not (a xor b);
    layer2_outputs(2404) <= b;
    layer2_outputs(2405) <= not a;
    layer2_outputs(2406) <= a or b;
    layer2_outputs(2407) <= b;
    layer2_outputs(2408) <= b;
    layer2_outputs(2409) <= a xor b;
    layer2_outputs(2410) <= not b or a;
    layer2_outputs(2411) <= b;
    layer2_outputs(2412) <= not (a and b);
    layer2_outputs(2413) <= not b;
    layer2_outputs(2414) <= a and not b;
    layer2_outputs(2415) <= not b;
    layer2_outputs(2416) <= not b;
    layer2_outputs(2417) <= a or b;
    layer2_outputs(2418) <= a;
    layer2_outputs(2419) <= not a or b;
    layer2_outputs(2420) <= not b or a;
    layer2_outputs(2421) <= not b;
    layer2_outputs(2422) <= a and b;
    layer2_outputs(2423) <= a or b;
    layer2_outputs(2424) <= not a or b;
    layer2_outputs(2425) <= not (a or b);
    layer2_outputs(2426) <= b and not a;
    layer2_outputs(2427) <= b;
    layer2_outputs(2428) <= not a;
    layer2_outputs(2429) <= a xor b;
    layer2_outputs(2430) <= a xor b;
    layer2_outputs(2431) <= not b;
    layer2_outputs(2432) <= a and b;
    layer2_outputs(2433) <= not (a xor b);
    layer2_outputs(2434) <= a and b;
    layer2_outputs(2435) <= not (a xor b);
    layer2_outputs(2436) <= not a;
    layer2_outputs(2437) <= not a;
    layer2_outputs(2438) <= a and b;
    layer2_outputs(2439) <= not b;
    layer2_outputs(2440) <= b;
    layer2_outputs(2441) <= not a;
    layer2_outputs(2442) <= not b;
    layer2_outputs(2443) <= a and b;
    layer2_outputs(2444) <= not a;
    layer2_outputs(2445) <= not a;
    layer2_outputs(2446) <= a;
    layer2_outputs(2447) <= b;
    layer2_outputs(2448) <= not (a xor b);
    layer2_outputs(2449) <= a and not b;
    layer2_outputs(2450) <= a;
    layer2_outputs(2451) <= a;
    layer2_outputs(2452) <= not (a xor b);
    layer2_outputs(2453) <= b;
    layer2_outputs(2454) <= not (a xor b);
    layer2_outputs(2455) <= not (a or b);
    layer2_outputs(2456) <= not a;
    layer2_outputs(2457) <= a and b;
    layer2_outputs(2458) <= not b or a;
    layer2_outputs(2459) <= not a;
    layer2_outputs(2460) <= b;
    layer2_outputs(2461) <= not (a xor b);
    layer2_outputs(2462) <= not b;
    layer2_outputs(2463) <= b and not a;
    layer2_outputs(2464) <= a;
    layer2_outputs(2465) <= b;
    layer2_outputs(2466) <= a and b;
    layer2_outputs(2467) <= a xor b;
    layer2_outputs(2468) <= a xor b;
    layer2_outputs(2469) <= not a;
    layer2_outputs(2470) <= not a;
    layer2_outputs(2471) <= b and not a;
    layer2_outputs(2472) <= b;
    layer2_outputs(2473) <= not (a xor b);
    layer2_outputs(2474) <= not a;
    layer2_outputs(2475) <= b;
    layer2_outputs(2476) <= a and not b;
    layer2_outputs(2477) <= a;
    layer2_outputs(2478) <= not b;
    layer2_outputs(2479) <= not a;
    layer2_outputs(2480) <= not (a xor b);
    layer2_outputs(2481) <= a xor b;
    layer2_outputs(2482) <= a;
    layer2_outputs(2483) <= a and not b;
    layer2_outputs(2484) <= a xor b;
    layer2_outputs(2485) <= a xor b;
    layer2_outputs(2486) <= not a or b;
    layer2_outputs(2487) <= not (a xor b);
    layer2_outputs(2488) <= not (a xor b);
    layer2_outputs(2489) <= not (a xor b);
    layer2_outputs(2490) <= not (a xor b);
    layer2_outputs(2491) <= a xor b;
    layer2_outputs(2492) <= a;
    layer2_outputs(2493) <= not (a xor b);
    layer2_outputs(2494) <= a;
    layer2_outputs(2495) <= not (a and b);
    layer2_outputs(2496) <= a xor b;
    layer2_outputs(2497) <= not a or b;
    layer2_outputs(2498) <= a and not b;
    layer2_outputs(2499) <= a xor b;
    layer2_outputs(2500) <= a;
    layer2_outputs(2501) <= not a;
    layer2_outputs(2502) <= a xor b;
    layer2_outputs(2503) <= b and not a;
    layer2_outputs(2504) <= a xor b;
    layer2_outputs(2505) <= not a;
    layer2_outputs(2506) <= b and not a;
    layer2_outputs(2507) <= not b;
    layer2_outputs(2508) <= not b or a;
    layer2_outputs(2509) <= not b;
    layer2_outputs(2510) <= not (a xor b);
    layer2_outputs(2511) <= not (a xor b);
    layer2_outputs(2512) <= b;
    layer2_outputs(2513) <= not (a and b);
    layer2_outputs(2514) <= b;
    layer2_outputs(2515) <= not a;
    layer2_outputs(2516) <= not a;
    layer2_outputs(2517) <= not a;
    layer2_outputs(2518) <= not b or a;
    layer2_outputs(2519) <= not a;
    layer2_outputs(2520) <= not (a or b);
    layer2_outputs(2521) <= a or b;
    layer2_outputs(2522) <= not a or b;
    layer2_outputs(2523) <= a;
    layer2_outputs(2524) <= a xor b;
    layer2_outputs(2525) <= not a or b;
    layer2_outputs(2526) <= not a;
    layer2_outputs(2527) <= b;
    layer2_outputs(2528) <= 1'b1;
    layer2_outputs(2529) <= a and not b;
    layer2_outputs(2530) <= not (a xor b);
    layer2_outputs(2531) <= not (a and b);
    layer2_outputs(2532) <= not a;
    layer2_outputs(2533) <= a;
    layer2_outputs(2534) <= b and not a;
    layer2_outputs(2535) <= b and not a;
    layer2_outputs(2536) <= a and b;
    layer2_outputs(2537) <= a and not b;
    layer2_outputs(2538) <= not b;
    layer2_outputs(2539) <= not (a and b);
    layer2_outputs(2540) <= a;
    layer2_outputs(2541) <= not (a and b);
    layer2_outputs(2542) <= not b;
    layer2_outputs(2543) <= a xor b;
    layer2_outputs(2544) <= not (a xor b);
    layer2_outputs(2545) <= a and not b;
    layer2_outputs(2546) <= not a;
    layer2_outputs(2547) <= not a;
    layer2_outputs(2548) <= a;
    layer2_outputs(2549) <= not a;
    layer2_outputs(2550) <= not (a and b);
    layer2_outputs(2551) <= a;
    layer2_outputs(2552) <= a xor b;
    layer2_outputs(2553) <= a;
    layer2_outputs(2554) <= a xor b;
    layer2_outputs(2555) <= a;
    layer2_outputs(2556) <= not a;
    layer2_outputs(2557) <= a xor b;
    layer2_outputs(2558) <= not (a and b);
    layer2_outputs(2559) <= b;
    layer2_outputs(2560) <= not b;
    layer2_outputs(2561) <= a;
    layer2_outputs(2562) <= a xor b;
    layer2_outputs(2563) <= not (a or b);
    layer2_outputs(2564) <= not a or b;
    layer2_outputs(2565) <= not b or a;
    layer2_outputs(2566) <= not a;
    layer2_outputs(2567) <= not (a xor b);
    layer2_outputs(2568) <= a;
    layer2_outputs(2569) <= not a or b;
    layer2_outputs(2570) <= b;
    layer2_outputs(2571) <= b;
    layer2_outputs(2572) <= not (a or b);
    layer2_outputs(2573) <= not a;
    layer2_outputs(2574) <= b;
    layer2_outputs(2575) <= not a or b;
    layer2_outputs(2576) <= not (a or b);
    layer2_outputs(2577) <= not (a and b);
    layer2_outputs(2578) <= b and not a;
    layer2_outputs(2579) <= a;
    layer2_outputs(2580) <= b;
    layer2_outputs(2581) <= b;
    layer2_outputs(2582) <= not b;
    layer2_outputs(2583) <= not (a and b);
    layer2_outputs(2584) <= b and not a;
    layer2_outputs(2585) <= not (a and b);
    layer2_outputs(2586) <= a;
    layer2_outputs(2587) <= not b;
    layer2_outputs(2588) <= a;
    layer2_outputs(2589) <= not (a or b);
    layer2_outputs(2590) <= a;
    layer2_outputs(2591) <= not (a and b);
    layer2_outputs(2592) <= a;
    layer2_outputs(2593) <= not a;
    layer2_outputs(2594) <= a;
    layer2_outputs(2595) <= b;
    layer2_outputs(2596) <= not b;
    layer2_outputs(2597) <= not a;
    layer2_outputs(2598) <= not a;
    layer2_outputs(2599) <= not (a xor b);
    layer2_outputs(2600) <= b and not a;
    layer2_outputs(2601) <= not b;
    layer2_outputs(2602) <= not b or a;
    layer2_outputs(2603) <= not a;
    layer2_outputs(2604) <= b;
    layer2_outputs(2605) <= not b;
    layer2_outputs(2606) <= a;
    layer2_outputs(2607) <= b and not a;
    layer2_outputs(2608) <= a xor b;
    layer2_outputs(2609) <= a and not b;
    layer2_outputs(2610) <= not b;
    layer2_outputs(2611) <= b;
    layer2_outputs(2612) <= not (a xor b);
    layer2_outputs(2613) <= not a or b;
    layer2_outputs(2614) <= not b or a;
    layer2_outputs(2615) <= not (a xor b);
    layer2_outputs(2616) <= b;
    layer2_outputs(2617) <= not a or b;
    layer2_outputs(2618) <= b;
    layer2_outputs(2619) <= a;
    layer2_outputs(2620) <= not b;
    layer2_outputs(2621) <= a;
    layer2_outputs(2622) <= not a or b;
    layer2_outputs(2623) <= a;
    layer2_outputs(2624) <= not a;
    layer2_outputs(2625) <= a xor b;
    layer2_outputs(2626) <= not a;
    layer2_outputs(2627) <= not (a xor b);
    layer2_outputs(2628) <= b;
    layer2_outputs(2629) <= not (a xor b);
    layer2_outputs(2630) <= a;
    layer2_outputs(2631) <= not (a and b);
    layer2_outputs(2632) <= a;
    layer2_outputs(2633) <= a xor b;
    layer2_outputs(2634) <= not (a xor b);
    layer2_outputs(2635) <= not (a xor b);
    layer2_outputs(2636) <= not a;
    layer2_outputs(2637) <= not a;
    layer2_outputs(2638) <= not b or a;
    layer2_outputs(2639) <= a;
    layer2_outputs(2640) <= a xor b;
    layer2_outputs(2641) <= a and not b;
    layer2_outputs(2642) <= b;
    layer2_outputs(2643) <= not b;
    layer2_outputs(2644) <= b;
    layer2_outputs(2645) <= not (a or b);
    layer2_outputs(2646) <= b;
    layer2_outputs(2647) <= b and not a;
    layer2_outputs(2648) <= b and not a;
    layer2_outputs(2649) <= b;
    layer2_outputs(2650) <= not b;
    layer2_outputs(2651) <= not (a xor b);
    layer2_outputs(2652) <= not b or a;
    layer2_outputs(2653) <= not (a xor b);
    layer2_outputs(2654) <= not (a and b);
    layer2_outputs(2655) <= not (a or b);
    layer2_outputs(2656) <= a;
    layer2_outputs(2657) <= not (a xor b);
    layer2_outputs(2658) <= not a or b;
    layer2_outputs(2659) <= not b;
    layer2_outputs(2660) <= a;
    layer2_outputs(2661) <= a;
    layer2_outputs(2662) <= not (a and b);
    layer2_outputs(2663) <= a or b;
    layer2_outputs(2664) <= b and not a;
    layer2_outputs(2665) <= not (a or b);
    layer2_outputs(2666) <= not (a xor b);
    layer2_outputs(2667) <= a and b;
    layer2_outputs(2668) <= not a;
    layer2_outputs(2669) <= a xor b;
    layer2_outputs(2670) <= b and not a;
    layer2_outputs(2671) <= b;
    layer2_outputs(2672) <= a xor b;
    layer2_outputs(2673) <= not b;
    layer2_outputs(2674) <= b and not a;
    layer2_outputs(2675) <= a and b;
    layer2_outputs(2676) <= not (a xor b);
    layer2_outputs(2677) <= not a;
    layer2_outputs(2678) <= a;
    layer2_outputs(2679) <= not (a and b);
    layer2_outputs(2680) <= a;
    layer2_outputs(2681) <= not a;
    layer2_outputs(2682) <= not a;
    layer2_outputs(2683) <= not (a or b);
    layer2_outputs(2684) <= a and not b;
    layer2_outputs(2685) <= a;
    layer2_outputs(2686) <= not a;
    layer2_outputs(2687) <= b;
    layer2_outputs(2688) <= a xor b;
    layer2_outputs(2689) <= a xor b;
    layer2_outputs(2690) <= a or b;
    layer2_outputs(2691) <= a;
    layer2_outputs(2692) <= b;
    layer2_outputs(2693) <= not (a and b);
    layer2_outputs(2694) <= a and not b;
    layer2_outputs(2695) <= not (a or b);
    layer2_outputs(2696) <= not b or a;
    layer2_outputs(2697) <= a;
    layer2_outputs(2698) <= not b;
    layer2_outputs(2699) <= a xor b;
    layer2_outputs(2700) <= a;
    layer2_outputs(2701) <= not (a or b);
    layer2_outputs(2702) <= not b;
    layer2_outputs(2703) <= a;
    layer2_outputs(2704) <= b and not a;
    layer2_outputs(2705) <= a xor b;
    layer2_outputs(2706) <= not (a and b);
    layer2_outputs(2707) <= a xor b;
    layer2_outputs(2708) <= not (a xor b);
    layer2_outputs(2709) <= b;
    layer2_outputs(2710) <= not (a and b);
    layer2_outputs(2711) <= not (a or b);
    layer2_outputs(2712) <= not (a xor b);
    layer2_outputs(2713) <= not b or a;
    layer2_outputs(2714) <= a or b;
    layer2_outputs(2715) <= a xor b;
    layer2_outputs(2716) <= b and not a;
    layer2_outputs(2717) <= a and b;
    layer2_outputs(2718) <= a and not b;
    layer2_outputs(2719) <= not (a and b);
    layer2_outputs(2720) <= b and not a;
    layer2_outputs(2721) <= 1'b1;
    layer2_outputs(2722) <= b;
    layer2_outputs(2723) <= not a;
    layer2_outputs(2724) <= not b;
    layer2_outputs(2725) <= a;
    layer2_outputs(2726) <= not a;
    layer2_outputs(2727) <= a and not b;
    layer2_outputs(2728) <= not (a and b);
    layer2_outputs(2729) <= not (a xor b);
    layer2_outputs(2730) <= a and not b;
    layer2_outputs(2731) <= a xor b;
    layer2_outputs(2732) <= not b or a;
    layer2_outputs(2733) <= not (a and b);
    layer2_outputs(2734) <= a xor b;
    layer2_outputs(2735) <= a;
    layer2_outputs(2736) <= not a;
    layer2_outputs(2737) <= not (a or b);
    layer2_outputs(2738) <= a or b;
    layer2_outputs(2739) <= b;
    layer2_outputs(2740) <= a xor b;
    layer2_outputs(2741) <= a xor b;
    layer2_outputs(2742) <= not a;
    layer2_outputs(2743) <= b;
    layer2_outputs(2744) <= not (a xor b);
    layer2_outputs(2745) <= not (a xor b);
    layer2_outputs(2746) <= not (a xor b);
    layer2_outputs(2747) <= not (a xor b);
    layer2_outputs(2748) <= not (a xor b);
    layer2_outputs(2749) <= a;
    layer2_outputs(2750) <= not a;
    layer2_outputs(2751) <= a or b;
    layer2_outputs(2752) <= 1'b1;
    layer2_outputs(2753) <= not b;
    layer2_outputs(2754) <= b and not a;
    layer2_outputs(2755) <= not b;
    layer2_outputs(2756) <= not a or b;
    layer2_outputs(2757) <= a xor b;
    layer2_outputs(2758) <= not a or b;
    layer2_outputs(2759) <= not b;
    layer2_outputs(2760) <= not b or a;
    layer2_outputs(2761) <= a and not b;
    layer2_outputs(2762) <= not a or b;
    layer2_outputs(2763) <= not b;
    layer2_outputs(2764) <= not b;
    layer2_outputs(2765) <= not a or b;
    layer2_outputs(2766) <= a;
    layer2_outputs(2767) <= a;
    layer2_outputs(2768) <= b;
    layer2_outputs(2769) <= a;
    layer2_outputs(2770) <= not b;
    layer2_outputs(2771) <= not (a xor b);
    layer2_outputs(2772) <= b;
    layer2_outputs(2773) <= not b;
    layer2_outputs(2774) <= a xor b;
    layer2_outputs(2775) <= not a or b;
    layer2_outputs(2776) <= b;
    layer2_outputs(2777) <= a;
    layer2_outputs(2778) <= a xor b;
    layer2_outputs(2779) <= not a;
    layer2_outputs(2780) <= b;
    layer2_outputs(2781) <= b;
    layer2_outputs(2782) <= a xor b;
    layer2_outputs(2783) <= a xor b;
    layer2_outputs(2784) <= a and not b;
    layer2_outputs(2785) <= 1'b0;
    layer2_outputs(2786) <= a xor b;
    layer2_outputs(2787) <= a xor b;
    layer2_outputs(2788) <= a xor b;
    layer2_outputs(2789) <= a and not b;
    layer2_outputs(2790) <= not (a or b);
    layer2_outputs(2791) <= not a or b;
    layer2_outputs(2792) <= not (a xor b);
    layer2_outputs(2793) <= not a;
    layer2_outputs(2794) <= a or b;
    layer2_outputs(2795) <= a xor b;
    layer2_outputs(2796) <= b and not a;
    layer2_outputs(2797) <= a xor b;
    layer2_outputs(2798) <= not a;
    layer2_outputs(2799) <= not a;
    layer2_outputs(2800) <= a;
    layer2_outputs(2801) <= b;
    layer2_outputs(2802) <= not (a xor b);
    layer2_outputs(2803) <= not (a xor b);
    layer2_outputs(2804) <= a;
    layer2_outputs(2805) <= not a;
    layer2_outputs(2806) <= not b;
    layer2_outputs(2807) <= a xor b;
    layer2_outputs(2808) <= a or b;
    layer2_outputs(2809) <= not a or b;
    layer2_outputs(2810) <= not (a and b);
    layer2_outputs(2811) <= a xor b;
    layer2_outputs(2812) <= a and b;
    layer2_outputs(2813) <= b;
    layer2_outputs(2814) <= a;
    layer2_outputs(2815) <= not b;
    layer2_outputs(2816) <= b;
    layer2_outputs(2817) <= a;
    layer2_outputs(2818) <= b and not a;
    layer2_outputs(2819) <= b;
    layer2_outputs(2820) <= a and b;
    layer2_outputs(2821) <= a and not b;
    layer2_outputs(2822) <= a xor b;
    layer2_outputs(2823) <= not b or a;
    layer2_outputs(2824) <= b;
    layer2_outputs(2825) <= not (a xor b);
    layer2_outputs(2826) <= a and not b;
    layer2_outputs(2827) <= b;
    layer2_outputs(2828) <= a and b;
    layer2_outputs(2829) <= not b;
    layer2_outputs(2830) <= not (a and b);
    layer2_outputs(2831) <= not (a and b);
    layer2_outputs(2832) <= not (a xor b);
    layer2_outputs(2833) <= not a;
    layer2_outputs(2834) <= not a or b;
    layer2_outputs(2835) <= not (a xor b);
    layer2_outputs(2836) <= not a or b;
    layer2_outputs(2837) <= a xor b;
    layer2_outputs(2838) <= a or b;
    layer2_outputs(2839) <= a;
    layer2_outputs(2840) <= not a;
    layer2_outputs(2841) <= 1'b1;
    layer2_outputs(2842) <= not a or b;
    layer2_outputs(2843) <= a;
    layer2_outputs(2844) <= a xor b;
    layer2_outputs(2845) <= a xor b;
    layer2_outputs(2846) <= a or b;
    layer2_outputs(2847) <= a xor b;
    layer2_outputs(2848) <= not (a and b);
    layer2_outputs(2849) <= a xor b;
    layer2_outputs(2850) <= b;
    layer2_outputs(2851) <= a;
    layer2_outputs(2852) <= a;
    layer2_outputs(2853) <= not b;
    layer2_outputs(2854) <= b;
    layer2_outputs(2855) <= not a or b;
    layer2_outputs(2856) <= not a or b;
    layer2_outputs(2857) <= not (a or b);
    layer2_outputs(2858) <= a;
    layer2_outputs(2859) <= b;
    layer2_outputs(2860) <= b;
    layer2_outputs(2861) <= a and b;
    layer2_outputs(2862) <= a and not b;
    layer2_outputs(2863) <= a xor b;
    layer2_outputs(2864) <= b and not a;
    layer2_outputs(2865) <= not a or b;
    layer2_outputs(2866) <= not (a or b);
    layer2_outputs(2867) <= not (a or b);
    layer2_outputs(2868) <= not (a xor b);
    layer2_outputs(2869) <= a and b;
    layer2_outputs(2870) <= not a;
    layer2_outputs(2871) <= a or b;
    layer2_outputs(2872) <= not b;
    layer2_outputs(2873) <= b and not a;
    layer2_outputs(2874) <= a or b;
    layer2_outputs(2875) <= a or b;
    layer2_outputs(2876) <= not b or a;
    layer2_outputs(2877) <= not b;
    layer2_outputs(2878) <= a xor b;
    layer2_outputs(2879) <= 1'b1;
    layer2_outputs(2880) <= not a;
    layer2_outputs(2881) <= not (a xor b);
    layer2_outputs(2882) <= not (a or b);
    layer2_outputs(2883) <= a;
    layer2_outputs(2884) <= a;
    layer2_outputs(2885) <= a;
    layer2_outputs(2886) <= not a;
    layer2_outputs(2887) <= b;
    layer2_outputs(2888) <= not (a or b);
    layer2_outputs(2889) <= b;
    layer2_outputs(2890) <= not (a and b);
    layer2_outputs(2891) <= a xor b;
    layer2_outputs(2892) <= not (a and b);
    layer2_outputs(2893) <= not (a or b);
    layer2_outputs(2894) <= a;
    layer2_outputs(2895) <= not a;
    layer2_outputs(2896) <= a xor b;
    layer2_outputs(2897) <= b and not a;
    layer2_outputs(2898) <= a xor b;
    layer2_outputs(2899) <= a xor b;
    layer2_outputs(2900) <= not a;
    layer2_outputs(2901) <= not a or b;
    layer2_outputs(2902) <= not b;
    layer2_outputs(2903) <= b;
    layer2_outputs(2904) <= not a;
    layer2_outputs(2905) <= not a or b;
    layer2_outputs(2906) <= a xor b;
    layer2_outputs(2907) <= a and b;
    layer2_outputs(2908) <= a and b;
    layer2_outputs(2909) <= not (a or b);
    layer2_outputs(2910) <= a;
    layer2_outputs(2911) <= not (a or b);
    layer2_outputs(2912) <= not a or b;
    layer2_outputs(2913) <= b;
    layer2_outputs(2914) <= not a;
    layer2_outputs(2915) <= not a;
    layer2_outputs(2916) <= not b;
    layer2_outputs(2917) <= a xor b;
    layer2_outputs(2918) <= not (a and b);
    layer2_outputs(2919) <= b;
    layer2_outputs(2920) <= a xor b;
    layer2_outputs(2921) <= not (a or b);
    layer2_outputs(2922) <= not (a xor b);
    layer2_outputs(2923) <= not b;
    layer2_outputs(2924) <= a;
    layer2_outputs(2925) <= b;
    layer2_outputs(2926) <= not b;
    layer2_outputs(2927) <= not a or b;
    layer2_outputs(2928) <= not (a or b);
    layer2_outputs(2929) <= not (a and b);
    layer2_outputs(2930) <= not a or b;
    layer2_outputs(2931) <= not a;
    layer2_outputs(2932) <= a;
    layer2_outputs(2933) <= not (a xor b);
    layer2_outputs(2934) <= a and b;
    layer2_outputs(2935) <= a xor b;
    layer2_outputs(2936) <= a and b;
    layer2_outputs(2937) <= not b or a;
    layer2_outputs(2938) <= not (a or b);
    layer2_outputs(2939) <= b;
    layer2_outputs(2940) <= not (a or b);
    layer2_outputs(2941) <= not b or a;
    layer2_outputs(2942) <= not b or a;
    layer2_outputs(2943) <= not a;
    layer2_outputs(2944) <= b;
    layer2_outputs(2945) <= not (a xor b);
    layer2_outputs(2946) <= not (a or b);
    layer2_outputs(2947) <= not (a xor b);
    layer2_outputs(2948) <= not a;
    layer2_outputs(2949) <= not b;
    layer2_outputs(2950) <= not b;
    layer2_outputs(2951) <= not a;
    layer2_outputs(2952) <= a;
    layer2_outputs(2953) <= not b;
    layer2_outputs(2954) <= b and not a;
    layer2_outputs(2955) <= not a;
    layer2_outputs(2956) <= a xor b;
    layer2_outputs(2957) <= a;
    layer2_outputs(2958) <= a or b;
    layer2_outputs(2959) <= b;
    layer2_outputs(2960) <= a xor b;
    layer2_outputs(2961) <= not b or a;
    layer2_outputs(2962) <= not (a xor b);
    layer2_outputs(2963) <= a xor b;
    layer2_outputs(2964) <= a xor b;
    layer2_outputs(2965) <= b;
    layer2_outputs(2966) <= not (a and b);
    layer2_outputs(2967) <= not (a xor b);
    layer2_outputs(2968) <= not b;
    layer2_outputs(2969) <= not b or a;
    layer2_outputs(2970) <= a xor b;
    layer2_outputs(2971) <= not a or b;
    layer2_outputs(2972) <= b;
    layer2_outputs(2973) <= a and not b;
    layer2_outputs(2974) <= not (a and b);
    layer2_outputs(2975) <= not b;
    layer2_outputs(2976) <= not (a and b);
    layer2_outputs(2977) <= not (a xor b);
    layer2_outputs(2978) <= a;
    layer2_outputs(2979) <= a xor b;
    layer2_outputs(2980) <= not (a xor b);
    layer2_outputs(2981) <= not (a xor b);
    layer2_outputs(2982) <= a;
    layer2_outputs(2983) <= not b;
    layer2_outputs(2984) <= not (a and b);
    layer2_outputs(2985) <= b;
    layer2_outputs(2986) <= not b or a;
    layer2_outputs(2987) <= not (a or b);
    layer2_outputs(2988) <= a and not b;
    layer2_outputs(2989) <= a or b;
    layer2_outputs(2990) <= a and b;
    layer2_outputs(2991) <= b;
    layer2_outputs(2992) <= a and b;
    layer2_outputs(2993) <= b;
    layer2_outputs(2994) <= not b;
    layer2_outputs(2995) <= not a or b;
    layer2_outputs(2996) <= not a;
    layer2_outputs(2997) <= b;
    layer2_outputs(2998) <= a;
    layer2_outputs(2999) <= not a;
    layer2_outputs(3000) <= a and not b;
    layer2_outputs(3001) <= not b or a;
    layer2_outputs(3002) <= a xor b;
    layer2_outputs(3003) <= a and b;
    layer2_outputs(3004) <= not a or b;
    layer2_outputs(3005) <= a or b;
    layer2_outputs(3006) <= not b;
    layer2_outputs(3007) <= not (a and b);
    layer2_outputs(3008) <= b and not a;
    layer2_outputs(3009) <= a;
    layer2_outputs(3010) <= a xor b;
    layer2_outputs(3011) <= a;
    layer2_outputs(3012) <= a and not b;
    layer2_outputs(3013) <= b;
    layer2_outputs(3014) <= b;
    layer2_outputs(3015) <= b;
    layer2_outputs(3016) <= not a;
    layer2_outputs(3017) <= not b or a;
    layer2_outputs(3018) <= a or b;
    layer2_outputs(3019) <= not a or b;
    layer2_outputs(3020) <= b;
    layer2_outputs(3021) <= a xor b;
    layer2_outputs(3022) <= not (a and b);
    layer2_outputs(3023) <= not b or a;
    layer2_outputs(3024) <= not (a and b);
    layer2_outputs(3025) <= not a;
    layer2_outputs(3026) <= a and b;
    layer2_outputs(3027) <= b;
    layer2_outputs(3028) <= not a;
    layer2_outputs(3029) <= not (a xor b);
    layer2_outputs(3030) <= a;
    layer2_outputs(3031) <= not a;
    layer2_outputs(3032) <= not (a xor b);
    layer2_outputs(3033) <= not b or a;
    layer2_outputs(3034) <= not b;
    layer2_outputs(3035) <= not (a and b);
    layer2_outputs(3036) <= a and b;
    layer2_outputs(3037) <= not a;
    layer2_outputs(3038) <= b;
    layer2_outputs(3039) <= b;
    layer2_outputs(3040) <= a and b;
    layer2_outputs(3041) <= not b;
    layer2_outputs(3042) <= not a;
    layer2_outputs(3043) <= a;
    layer2_outputs(3044) <= a xor b;
    layer2_outputs(3045) <= a;
    layer2_outputs(3046) <= a;
    layer2_outputs(3047) <= a;
    layer2_outputs(3048) <= not b or a;
    layer2_outputs(3049) <= a;
    layer2_outputs(3050) <= not (a xor b);
    layer2_outputs(3051) <= not (a and b);
    layer2_outputs(3052) <= not b or a;
    layer2_outputs(3053) <= a;
    layer2_outputs(3054) <= not (a or b);
    layer2_outputs(3055) <= a or b;
    layer2_outputs(3056) <= b and not a;
    layer2_outputs(3057) <= a xor b;
    layer2_outputs(3058) <= a and not b;
    layer2_outputs(3059) <= not a;
    layer2_outputs(3060) <= not b;
    layer2_outputs(3061) <= not (a and b);
    layer2_outputs(3062) <= a;
    layer2_outputs(3063) <= not a;
    layer2_outputs(3064) <= a xor b;
    layer2_outputs(3065) <= a or b;
    layer2_outputs(3066) <= not a;
    layer2_outputs(3067) <= a or b;
    layer2_outputs(3068) <= a;
    layer2_outputs(3069) <= not b or a;
    layer2_outputs(3070) <= a xor b;
    layer2_outputs(3071) <= not (a and b);
    layer2_outputs(3072) <= a xor b;
    layer2_outputs(3073) <= not a;
    layer2_outputs(3074) <= not (a and b);
    layer2_outputs(3075) <= not b or a;
    layer2_outputs(3076) <= not a;
    layer2_outputs(3077) <= not (a and b);
    layer2_outputs(3078) <= a and b;
    layer2_outputs(3079) <= not b or a;
    layer2_outputs(3080) <= a xor b;
    layer2_outputs(3081) <= b and not a;
    layer2_outputs(3082) <= not b;
    layer2_outputs(3083) <= not b;
    layer2_outputs(3084) <= a;
    layer2_outputs(3085) <= a;
    layer2_outputs(3086) <= a;
    layer2_outputs(3087) <= not b;
    layer2_outputs(3088) <= not b;
    layer2_outputs(3089) <= a;
    layer2_outputs(3090) <= a;
    layer2_outputs(3091) <= a xor b;
    layer2_outputs(3092) <= not a;
    layer2_outputs(3093) <= not a;
    layer2_outputs(3094) <= a;
    layer2_outputs(3095) <= not a or b;
    layer2_outputs(3096) <= not b or a;
    layer2_outputs(3097) <= not b;
    layer2_outputs(3098) <= not a;
    layer2_outputs(3099) <= not a or b;
    layer2_outputs(3100) <= not (a or b);
    layer2_outputs(3101) <= not (a and b);
    layer2_outputs(3102) <= a xor b;
    layer2_outputs(3103) <= not (a and b);
    layer2_outputs(3104) <= a;
    layer2_outputs(3105) <= a xor b;
    layer2_outputs(3106) <= not a;
    layer2_outputs(3107) <= not (a xor b);
    layer2_outputs(3108) <= not b;
    layer2_outputs(3109) <= a xor b;
    layer2_outputs(3110) <= not b;
    layer2_outputs(3111) <= b;
    layer2_outputs(3112) <= a;
    layer2_outputs(3113) <= b;
    layer2_outputs(3114) <= not a or b;
    layer2_outputs(3115) <= not (a or b);
    layer2_outputs(3116) <= not (a or b);
    layer2_outputs(3117) <= not (a xor b);
    layer2_outputs(3118) <= a xor b;
    layer2_outputs(3119) <= b and not a;
    layer2_outputs(3120) <= not (a and b);
    layer2_outputs(3121) <= not (a xor b);
    layer2_outputs(3122) <= not (a or b);
    layer2_outputs(3123) <= b;
    layer2_outputs(3124) <= a xor b;
    layer2_outputs(3125) <= a and not b;
    layer2_outputs(3126) <= not b;
    layer2_outputs(3127) <= a;
    layer2_outputs(3128) <= not b;
    layer2_outputs(3129) <= not (a or b);
    layer2_outputs(3130) <= a;
    layer2_outputs(3131) <= b;
    layer2_outputs(3132) <= b;
    layer2_outputs(3133) <= not (a xor b);
    layer2_outputs(3134) <= not a;
    layer2_outputs(3135) <= not (a xor b);
    layer2_outputs(3136) <= a xor b;
    layer2_outputs(3137) <= not b or a;
    layer2_outputs(3138) <= not (a and b);
    layer2_outputs(3139) <= a;
    layer2_outputs(3140) <= not a;
    layer2_outputs(3141) <= a or b;
    layer2_outputs(3142) <= not (a xor b);
    layer2_outputs(3143) <= b;
    layer2_outputs(3144) <= a xor b;
    layer2_outputs(3145) <= not b;
    layer2_outputs(3146) <= a xor b;
    layer2_outputs(3147) <= not a;
    layer2_outputs(3148) <= a;
    layer2_outputs(3149) <= not (a xor b);
    layer2_outputs(3150) <= a xor b;
    layer2_outputs(3151) <= not (a and b);
    layer2_outputs(3152) <= not b;
    layer2_outputs(3153) <= not (a or b);
    layer2_outputs(3154) <= a or b;
    layer2_outputs(3155) <= not (a xor b);
    layer2_outputs(3156) <= a;
    layer2_outputs(3157) <= a and b;
    layer2_outputs(3158) <= a xor b;
    layer2_outputs(3159) <= a;
    layer2_outputs(3160) <= not (a xor b);
    layer2_outputs(3161) <= not (a or b);
    layer2_outputs(3162) <= a and not b;
    layer2_outputs(3163) <= not (a or b);
    layer2_outputs(3164) <= a or b;
    layer2_outputs(3165) <= b;
    layer2_outputs(3166) <= not b;
    layer2_outputs(3167) <= not a or b;
    layer2_outputs(3168) <= not a;
    layer2_outputs(3169) <= not (a and b);
    layer2_outputs(3170) <= not (a xor b);
    layer2_outputs(3171) <= a xor b;
    layer2_outputs(3172) <= a xor b;
    layer2_outputs(3173) <= a or b;
    layer2_outputs(3174) <= not (a xor b);
    layer2_outputs(3175) <= b;
    layer2_outputs(3176) <= a or b;
    layer2_outputs(3177) <= b;
    layer2_outputs(3178) <= not b;
    layer2_outputs(3179) <= a xor b;
    layer2_outputs(3180) <= b and not a;
    layer2_outputs(3181) <= not b;
    layer2_outputs(3182) <= not (a xor b);
    layer2_outputs(3183) <= b;
    layer2_outputs(3184) <= b and not a;
    layer2_outputs(3185) <= not a;
    layer2_outputs(3186) <= not a or b;
    layer2_outputs(3187) <= b;
    layer2_outputs(3188) <= not (a and b);
    layer2_outputs(3189) <= a;
    layer2_outputs(3190) <= a or b;
    layer2_outputs(3191) <= a and b;
    layer2_outputs(3192) <= a xor b;
    layer2_outputs(3193) <= not (a and b);
    layer2_outputs(3194) <= not a;
    layer2_outputs(3195) <= a and b;
    layer2_outputs(3196) <= b;
    layer2_outputs(3197) <= not a or b;
    layer2_outputs(3198) <= not (a xor b);
    layer2_outputs(3199) <= a and b;
    layer2_outputs(3200) <= b;
    layer2_outputs(3201) <= not b;
    layer2_outputs(3202) <= not a;
    layer2_outputs(3203) <= not b or a;
    layer2_outputs(3204) <= a and not b;
    layer2_outputs(3205) <= not (a and b);
    layer2_outputs(3206) <= a and b;
    layer2_outputs(3207) <= 1'b1;
    layer2_outputs(3208) <= not a or b;
    layer2_outputs(3209) <= not a or b;
    layer2_outputs(3210) <= not (a xor b);
    layer2_outputs(3211) <= a;
    layer2_outputs(3212) <= not a;
    layer2_outputs(3213) <= a or b;
    layer2_outputs(3214) <= a or b;
    layer2_outputs(3215) <= not (a xor b);
    layer2_outputs(3216) <= a xor b;
    layer2_outputs(3217) <= a and b;
    layer2_outputs(3218) <= not b;
    layer2_outputs(3219) <= a;
    layer2_outputs(3220) <= a;
    layer2_outputs(3221) <= a;
    layer2_outputs(3222) <= b and not a;
    layer2_outputs(3223) <= not a or b;
    layer2_outputs(3224) <= a xor b;
    layer2_outputs(3225) <= not a or b;
    layer2_outputs(3226) <= not b;
    layer2_outputs(3227) <= a and b;
    layer2_outputs(3228) <= not (a xor b);
    layer2_outputs(3229) <= b;
    layer2_outputs(3230) <= 1'b0;
    layer2_outputs(3231) <= b;
    layer2_outputs(3232) <= b and not a;
    layer2_outputs(3233) <= not a;
    layer2_outputs(3234) <= not (a or b);
    layer2_outputs(3235) <= a and b;
    layer2_outputs(3236) <= not a or b;
    layer2_outputs(3237) <= not b or a;
    layer2_outputs(3238) <= not (a or b);
    layer2_outputs(3239) <= a;
    layer2_outputs(3240) <= a xor b;
    layer2_outputs(3241) <= not a;
    layer2_outputs(3242) <= not b or a;
    layer2_outputs(3243) <= a;
    layer2_outputs(3244) <= not (a or b);
    layer2_outputs(3245) <= not a or b;
    layer2_outputs(3246) <= not b;
    layer2_outputs(3247) <= a or b;
    layer2_outputs(3248) <= b;
    layer2_outputs(3249) <= b;
    layer2_outputs(3250) <= a and not b;
    layer2_outputs(3251) <= a or b;
    layer2_outputs(3252) <= not b;
    layer2_outputs(3253) <= not a or b;
    layer2_outputs(3254) <= not b;
    layer2_outputs(3255) <= not (a and b);
    layer2_outputs(3256) <= b;
    layer2_outputs(3257) <= not (a and b);
    layer2_outputs(3258) <= a and not b;
    layer2_outputs(3259) <= not a or b;
    layer2_outputs(3260) <= a;
    layer2_outputs(3261) <= not b or a;
    layer2_outputs(3262) <= a xor b;
    layer2_outputs(3263) <= not a;
    layer2_outputs(3264) <= b;
    layer2_outputs(3265) <= not a;
    layer2_outputs(3266) <= a and not b;
    layer2_outputs(3267) <= a;
    layer2_outputs(3268) <= a xor b;
    layer2_outputs(3269) <= a xor b;
    layer2_outputs(3270) <= not (a xor b);
    layer2_outputs(3271) <= a;
    layer2_outputs(3272) <= not (a xor b);
    layer2_outputs(3273) <= a and b;
    layer2_outputs(3274) <= a xor b;
    layer2_outputs(3275) <= not a;
    layer2_outputs(3276) <= b;
    layer2_outputs(3277) <= not (a or b);
    layer2_outputs(3278) <= a;
    layer2_outputs(3279) <= not b or a;
    layer2_outputs(3280) <= b and not a;
    layer2_outputs(3281) <= a and not b;
    layer2_outputs(3282) <= not (a or b);
    layer2_outputs(3283) <= not b;
    layer2_outputs(3284) <= not (a or b);
    layer2_outputs(3285) <= a;
    layer2_outputs(3286) <= b and not a;
    layer2_outputs(3287) <= not a;
    layer2_outputs(3288) <= b;
    layer2_outputs(3289) <= not (a and b);
    layer2_outputs(3290) <= not a;
    layer2_outputs(3291) <= not (a xor b);
    layer2_outputs(3292) <= not (a xor b);
    layer2_outputs(3293) <= not b or a;
    layer2_outputs(3294) <= a xor b;
    layer2_outputs(3295) <= not b;
    layer2_outputs(3296) <= a xor b;
    layer2_outputs(3297) <= not (a xor b);
    layer2_outputs(3298) <= b;
    layer2_outputs(3299) <= not b;
    layer2_outputs(3300) <= not a;
    layer2_outputs(3301) <= a xor b;
    layer2_outputs(3302) <= not (a xor b);
    layer2_outputs(3303) <= not a;
    layer2_outputs(3304) <= a and not b;
    layer2_outputs(3305) <= a and not b;
    layer2_outputs(3306) <= a and b;
    layer2_outputs(3307) <= not b;
    layer2_outputs(3308) <= a and b;
    layer2_outputs(3309) <= a or b;
    layer2_outputs(3310) <= not a;
    layer2_outputs(3311) <= not a;
    layer2_outputs(3312) <= not a;
    layer2_outputs(3313) <= a and not b;
    layer2_outputs(3314) <= not (a xor b);
    layer2_outputs(3315) <= not (a or b);
    layer2_outputs(3316) <= not a or b;
    layer2_outputs(3317) <= a xor b;
    layer2_outputs(3318) <= not a or b;
    layer2_outputs(3319) <= not (a and b);
    layer2_outputs(3320) <= a and b;
    layer2_outputs(3321) <= not a;
    layer2_outputs(3322) <= not (a or b);
    layer2_outputs(3323) <= not a or b;
    layer2_outputs(3324) <= a xor b;
    layer2_outputs(3325) <= a or b;
    layer2_outputs(3326) <= not (a xor b);
    layer2_outputs(3327) <= a xor b;
    layer2_outputs(3328) <= b;
    layer2_outputs(3329) <= a and not b;
    layer2_outputs(3330) <= not b or a;
    layer2_outputs(3331) <= not (a or b);
    layer2_outputs(3332) <= a and not b;
    layer2_outputs(3333) <= not b;
    layer2_outputs(3334) <= a and not b;
    layer2_outputs(3335) <= not a or b;
    layer2_outputs(3336) <= 1'b0;
    layer2_outputs(3337) <= not a or b;
    layer2_outputs(3338) <= not b;
    layer2_outputs(3339) <= not a;
    layer2_outputs(3340) <= a and not b;
    layer2_outputs(3341) <= not a;
    layer2_outputs(3342) <= a xor b;
    layer2_outputs(3343) <= not b;
    layer2_outputs(3344) <= not b;
    layer2_outputs(3345) <= a xor b;
    layer2_outputs(3346) <= b and not a;
    layer2_outputs(3347) <= not b or a;
    layer2_outputs(3348) <= not b;
    layer2_outputs(3349) <= b;
    layer2_outputs(3350) <= not b;
    layer2_outputs(3351) <= not b or a;
    layer2_outputs(3352) <= not (a and b);
    layer2_outputs(3353) <= not (a and b);
    layer2_outputs(3354) <= b and not a;
    layer2_outputs(3355) <= a;
    layer2_outputs(3356) <= a and b;
    layer2_outputs(3357) <= a and not b;
    layer2_outputs(3358) <= not a;
    layer2_outputs(3359) <= a xor b;
    layer2_outputs(3360) <= not a;
    layer2_outputs(3361) <= not a;
    layer2_outputs(3362) <= a xor b;
    layer2_outputs(3363) <= not a or b;
    layer2_outputs(3364) <= not a or b;
    layer2_outputs(3365) <= not b;
    layer2_outputs(3366) <= not a;
    layer2_outputs(3367) <= not a or b;
    layer2_outputs(3368) <= not (a xor b);
    layer2_outputs(3369) <= not a;
    layer2_outputs(3370) <= not a;
    layer2_outputs(3371) <= a;
    layer2_outputs(3372) <= not b;
    layer2_outputs(3373) <= not (a or b);
    layer2_outputs(3374) <= not b or a;
    layer2_outputs(3375) <= not a;
    layer2_outputs(3376) <= not b or a;
    layer2_outputs(3377) <= not a;
    layer2_outputs(3378) <= not a;
    layer2_outputs(3379) <= b and not a;
    layer2_outputs(3380) <= a xor b;
    layer2_outputs(3381) <= b and not a;
    layer2_outputs(3382) <= b and not a;
    layer2_outputs(3383) <= not b;
    layer2_outputs(3384) <= not b;
    layer2_outputs(3385) <= a;
    layer2_outputs(3386) <= a xor b;
    layer2_outputs(3387) <= a;
    layer2_outputs(3388) <= not b;
    layer2_outputs(3389) <= a or b;
    layer2_outputs(3390) <= not a;
    layer2_outputs(3391) <= not b;
    layer2_outputs(3392) <= a;
    layer2_outputs(3393) <= a;
    layer2_outputs(3394) <= a and not b;
    layer2_outputs(3395) <= a and b;
    layer2_outputs(3396) <= not b;
    layer2_outputs(3397) <= a or b;
    layer2_outputs(3398) <= a xor b;
    layer2_outputs(3399) <= a;
    layer2_outputs(3400) <= not a or b;
    layer2_outputs(3401) <= a or b;
    layer2_outputs(3402) <= a;
    layer2_outputs(3403) <= not a or b;
    layer2_outputs(3404) <= b;
    layer2_outputs(3405) <= not (a xor b);
    layer2_outputs(3406) <= a xor b;
    layer2_outputs(3407) <= b and not a;
    layer2_outputs(3408) <= not a;
    layer2_outputs(3409) <= a and not b;
    layer2_outputs(3410) <= not b;
    layer2_outputs(3411) <= a xor b;
    layer2_outputs(3412) <= a;
    layer2_outputs(3413) <= not a;
    layer2_outputs(3414) <= not (a xor b);
    layer2_outputs(3415) <= b;
    layer2_outputs(3416) <= not (a xor b);
    layer2_outputs(3417) <= a and b;
    layer2_outputs(3418) <= a xor b;
    layer2_outputs(3419) <= b and not a;
    layer2_outputs(3420) <= a xor b;
    layer2_outputs(3421) <= not (a or b);
    layer2_outputs(3422) <= not b or a;
    layer2_outputs(3423) <= not (a or b);
    layer2_outputs(3424) <= b and not a;
    layer2_outputs(3425) <= a;
    layer2_outputs(3426) <= not b;
    layer2_outputs(3427) <= b;
    layer2_outputs(3428) <= b;
    layer2_outputs(3429) <= a and b;
    layer2_outputs(3430) <= a;
    layer2_outputs(3431) <= b;
    layer2_outputs(3432) <= not (a xor b);
    layer2_outputs(3433) <= b and not a;
    layer2_outputs(3434) <= not b or a;
    layer2_outputs(3435) <= not a;
    layer2_outputs(3436) <= not (a xor b);
    layer2_outputs(3437) <= b and not a;
    layer2_outputs(3438) <= not (a xor b);
    layer2_outputs(3439) <= b;
    layer2_outputs(3440) <= b and not a;
    layer2_outputs(3441) <= b;
    layer2_outputs(3442) <= b and not a;
    layer2_outputs(3443) <= not a;
    layer2_outputs(3444) <= a and b;
    layer2_outputs(3445) <= b;
    layer2_outputs(3446) <= a xor b;
    layer2_outputs(3447) <= not b or a;
    layer2_outputs(3448) <= a xor b;
    layer2_outputs(3449) <= not a;
    layer2_outputs(3450) <= a;
    layer2_outputs(3451) <= not (a xor b);
    layer2_outputs(3452) <= a xor b;
    layer2_outputs(3453) <= not b;
    layer2_outputs(3454) <= not (a and b);
    layer2_outputs(3455) <= a and not b;
    layer2_outputs(3456) <= a;
    layer2_outputs(3457) <= not b or a;
    layer2_outputs(3458) <= not a or b;
    layer2_outputs(3459) <= a and b;
    layer2_outputs(3460) <= not b or a;
    layer2_outputs(3461) <= a xor b;
    layer2_outputs(3462) <= a;
    layer2_outputs(3463) <= not a or b;
    layer2_outputs(3464) <= a xor b;
    layer2_outputs(3465) <= a;
    layer2_outputs(3466) <= not a;
    layer2_outputs(3467) <= a and b;
    layer2_outputs(3468) <= not b;
    layer2_outputs(3469) <= a or b;
    layer2_outputs(3470) <= not (a xor b);
    layer2_outputs(3471) <= b;
    layer2_outputs(3472) <= not b;
    layer2_outputs(3473) <= a;
    layer2_outputs(3474) <= b and not a;
    layer2_outputs(3475) <= not b;
    layer2_outputs(3476) <= not b or a;
    layer2_outputs(3477) <= a and not b;
    layer2_outputs(3478) <= not (a xor b);
    layer2_outputs(3479) <= not b or a;
    layer2_outputs(3480) <= a xor b;
    layer2_outputs(3481) <= a xor b;
    layer2_outputs(3482) <= not (a xor b);
    layer2_outputs(3483) <= a or b;
    layer2_outputs(3484) <= not (a xor b);
    layer2_outputs(3485) <= a xor b;
    layer2_outputs(3486) <= a;
    layer2_outputs(3487) <= b;
    layer2_outputs(3488) <= b;
    layer2_outputs(3489) <= not (a and b);
    layer2_outputs(3490) <= not b or a;
    layer2_outputs(3491) <= not a or b;
    layer2_outputs(3492) <= not a;
    layer2_outputs(3493) <= not (a xor b);
    layer2_outputs(3494) <= not b or a;
    layer2_outputs(3495) <= not (a and b);
    layer2_outputs(3496) <= b and not a;
    layer2_outputs(3497) <= a or b;
    layer2_outputs(3498) <= b and not a;
    layer2_outputs(3499) <= not b or a;
    layer2_outputs(3500) <= not (a xor b);
    layer2_outputs(3501) <= not (a xor b);
    layer2_outputs(3502) <= not (a and b);
    layer2_outputs(3503) <= b and not a;
    layer2_outputs(3504) <= a;
    layer2_outputs(3505) <= b;
    layer2_outputs(3506) <= a and not b;
    layer2_outputs(3507) <= b;
    layer2_outputs(3508) <= a and b;
    layer2_outputs(3509) <= not (a or b);
    layer2_outputs(3510) <= b;
    layer2_outputs(3511) <= b and not a;
    layer2_outputs(3512) <= 1'b0;
    layer2_outputs(3513) <= not (a xor b);
    layer2_outputs(3514) <= not b;
    layer2_outputs(3515) <= a or b;
    layer2_outputs(3516) <= not (a and b);
    layer2_outputs(3517) <= a and not b;
    layer2_outputs(3518) <= not (a or b);
    layer2_outputs(3519) <= b;
    layer2_outputs(3520) <= a;
    layer2_outputs(3521) <= not b;
    layer2_outputs(3522) <= not a or b;
    layer2_outputs(3523) <= not a;
    layer2_outputs(3524) <= not a or b;
    layer2_outputs(3525) <= a xor b;
    layer2_outputs(3526) <= a xor b;
    layer2_outputs(3527) <= not b;
    layer2_outputs(3528) <= b and not a;
    layer2_outputs(3529) <= a;
    layer2_outputs(3530) <= not (a and b);
    layer2_outputs(3531) <= b and not a;
    layer2_outputs(3532) <= not (a or b);
    layer2_outputs(3533) <= not b or a;
    layer2_outputs(3534) <= a;
    layer2_outputs(3535) <= not (a xor b);
    layer2_outputs(3536) <= a xor b;
    layer2_outputs(3537) <= a or b;
    layer2_outputs(3538) <= not (a or b);
    layer2_outputs(3539) <= a or b;
    layer2_outputs(3540) <= not (a xor b);
    layer2_outputs(3541) <= not (a xor b);
    layer2_outputs(3542) <= b;
    layer2_outputs(3543) <= a;
    layer2_outputs(3544) <= a;
    layer2_outputs(3545) <= not (a xor b);
    layer2_outputs(3546) <= not a;
    layer2_outputs(3547) <= a xor b;
    layer2_outputs(3548) <= not b;
    layer2_outputs(3549) <= not (a xor b);
    layer2_outputs(3550) <= not (a or b);
    layer2_outputs(3551) <= a and b;
    layer2_outputs(3552) <= not b;
    layer2_outputs(3553) <= a xor b;
    layer2_outputs(3554) <= a;
    layer2_outputs(3555) <= b;
    layer2_outputs(3556) <= a and b;
    layer2_outputs(3557) <= a and b;
    layer2_outputs(3558) <= not b or a;
    layer2_outputs(3559) <= not (a xor b);
    layer2_outputs(3560) <= not (a xor b);
    layer2_outputs(3561) <= a;
    layer2_outputs(3562) <= not b or a;
    layer2_outputs(3563) <= not a or b;
    layer2_outputs(3564) <= not (a xor b);
    layer2_outputs(3565) <= a xor b;
    layer2_outputs(3566) <= a;
    layer2_outputs(3567) <= a xor b;
    layer2_outputs(3568) <= a and b;
    layer2_outputs(3569) <= not b;
    layer2_outputs(3570) <= not b;
    layer2_outputs(3571) <= b;
    layer2_outputs(3572) <= b;
    layer2_outputs(3573) <= a xor b;
    layer2_outputs(3574) <= not a;
    layer2_outputs(3575) <= not a;
    layer2_outputs(3576) <= a;
    layer2_outputs(3577) <= not (a xor b);
    layer2_outputs(3578) <= not a or b;
    layer2_outputs(3579) <= a xor b;
    layer2_outputs(3580) <= a and not b;
    layer2_outputs(3581) <= b;
    layer2_outputs(3582) <= not a or b;
    layer2_outputs(3583) <= not (a and b);
    layer2_outputs(3584) <= a and b;
    layer2_outputs(3585) <= not a;
    layer2_outputs(3586) <= not (a xor b);
    layer2_outputs(3587) <= a xor b;
    layer2_outputs(3588) <= not a or b;
    layer2_outputs(3589) <= b;
    layer2_outputs(3590) <= b;
    layer2_outputs(3591) <= not a;
    layer2_outputs(3592) <= a;
    layer2_outputs(3593) <= a or b;
    layer2_outputs(3594) <= not (a xor b);
    layer2_outputs(3595) <= not (a xor b);
    layer2_outputs(3596) <= a;
    layer2_outputs(3597) <= not (a xor b);
    layer2_outputs(3598) <= b and not a;
    layer2_outputs(3599) <= b and not a;
    layer2_outputs(3600) <= not b;
    layer2_outputs(3601) <= b and not a;
    layer2_outputs(3602) <= not b or a;
    layer2_outputs(3603) <= not (a or b);
    layer2_outputs(3604) <= a or b;
    layer2_outputs(3605) <= a and b;
    layer2_outputs(3606) <= not (a or b);
    layer2_outputs(3607) <= a;
    layer2_outputs(3608) <= not a;
    layer2_outputs(3609) <= not b;
    layer2_outputs(3610) <= not a or b;
    layer2_outputs(3611) <= a;
    layer2_outputs(3612) <= b;
    layer2_outputs(3613) <= not b;
    layer2_outputs(3614) <= not b;
    layer2_outputs(3615) <= a and b;
    layer2_outputs(3616) <= a xor b;
    layer2_outputs(3617) <= b;
    layer2_outputs(3618) <= b;
    layer2_outputs(3619) <= not b or a;
    layer2_outputs(3620) <= b and not a;
    layer2_outputs(3621) <= not (a xor b);
    layer2_outputs(3622) <= b and not a;
    layer2_outputs(3623) <= a;
    layer2_outputs(3624) <= b;
    layer2_outputs(3625) <= not a;
    layer2_outputs(3626) <= a;
    layer2_outputs(3627) <= not (a xor b);
    layer2_outputs(3628) <= not a;
    layer2_outputs(3629) <= not a;
    layer2_outputs(3630) <= not a or b;
    layer2_outputs(3631) <= not b;
    layer2_outputs(3632) <= a xor b;
    layer2_outputs(3633) <= a and not b;
    layer2_outputs(3634) <= a;
    layer2_outputs(3635) <= not b;
    layer2_outputs(3636) <= not a or b;
    layer2_outputs(3637) <= not b;
    layer2_outputs(3638) <= not a;
    layer2_outputs(3639) <= a and not b;
    layer2_outputs(3640) <= not b;
    layer2_outputs(3641) <= a and b;
    layer2_outputs(3642) <= not a or b;
    layer2_outputs(3643) <= b;
    layer2_outputs(3644) <= not a;
    layer2_outputs(3645) <= not a;
    layer2_outputs(3646) <= a and not b;
    layer2_outputs(3647) <= not a;
    layer2_outputs(3648) <= b;
    layer2_outputs(3649) <= not b or a;
    layer2_outputs(3650) <= b;
    layer2_outputs(3651) <= a;
    layer2_outputs(3652) <= not a or b;
    layer2_outputs(3653) <= not (a and b);
    layer2_outputs(3654) <= not (a and b);
    layer2_outputs(3655) <= a xor b;
    layer2_outputs(3656) <= a and not b;
    layer2_outputs(3657) <= a;
    layer2_outputs(3658) <= b;
    layer2_outputs(3659) <= not (a or b);
    layer2_outputs(3660) <= b;
    layer2_outputs(3661) <= a xor b;
    layer2_outputs(3662) <= b;
    layer2_outputs(3663) <= not b or a;
    layer2_outputs(3664) <= a xor b;
    layer2_outputs(3665) <= not (a xor b);
    layer2_outputs(3666) <= not (a xor b);
    layer2_outputs(3667) <= not b or a;
    layer2_outputs(3668) <= a or b;
    layer2_outputs(3669) <= b;
    layer2_outputs(3670) <= a or b;
    layer2_outputs(3671) <= b;
    layer2_outputs(3672) <= not a;
    layer2_outputs(3673) <= a;
    layer2_outputs(3674) <= not b;
    layer2_outputs(3675) <= b;
    layer2_outputs(3676) <= not (a or b);
    layer2_outputs(3677) <= a and not b;
    layer2_outputs(3678) <= a and not b;
    layer2_outputs(3679) <= a and not b;
    layer2_outputs(3680) <= not a;
    layer2_outputs(3681) <= not a;
    layer2_outputs(3682) <= not b;
    layer2_outputs(3683) <= b and not a;
    layer2_outputs(3684) <= not b or a;
    layer2_outputs(3685) <= a;
    layer2_outputs(3686) <= not b or a;
    layer2_outputs(3687) <= a and b;
    layer2_outputs(3688) <= b;
    layer2_outputs(3689) <= not b or a;
    layer2_outputs(3690) <= not a;
    layer2_outputs(3691) <= not (a xor b);
    layer2_outputs(3692) <= not b or a;
    layer2_outputs(3693) <= a;
    layer2_outputs(3694) <= a xor b;
    layer2_outputs(3695) <= b and not a;
    layer2_outputs(3696) <= a and not b;
    layer2_outputs(3697) <= not a or b;
    layer2_outputs(3698) <= not a or b;
    layer2_outputs(3699) <= not (a xor b);
    layer2_outputs(3700) <= not (a xor b);
    layer2_outputs(3701) <= a and not b;
    layer2_outputs(3702) <= a or b;
    layer2_outputs(3703) <= b;
    layer2_outputs(3704) <= a and not b;
    layer2_outputs(3705) <= not (a xor b);
    layer2_outputs(3706) <= not a;
    layer2_outputs(3707) <= a xor b;
    layer2_outputs(3708) <= b;
    layer2_outputs(3709) <= not b;
    layer2_outputs(3710) <= not (a xor b);
    layer2_outputs(3711) <= a;
    layer2_outputs(3712) <= a xor b;
    layer2_outputs(3713) <= b;
    layer2_outputs(3714) <= not a or b;
    layer2_outputs(3715) <= b and not a;
    layer2_outputs(3716) <= not b;
    layer2_outputs(3717) <= b;
    layer2_outputs(3718) <= not (a xor b);
    layer2_outputs(3719) <= not (a and b);
    layer2_outputs(3720) <= a xor b;
    layer2_outputs(3721) <= not (a xor b);
    layer2_outputs(3722) <= b;
    layer2_outputs(3723) <= not b;
    layer2_outputs(3724) <= b;
    layer2_outputs(3725) <= a and b;
    layer2_outputs(3726) <= not b;
    layer2_outputs(3727) <= b;
    layer2_outputs(3728) <= a and not b;
    layer2_outputs(3729) <= a and b;
    layer2_outputs(3730) <= a xor b;
    layer2_outputs(3731) <= a and b;
    layer2_outputs(3732) <= a xor b;
    layer2_outputs(3733) <= not b;
    layer2_outputs(3734) <= a;
    layer2_outputs(3735) <= not b;
    layer2_outputs(3736) <= b;
    layer2_outputs(3737) <= b;
    layer2_outputs(3738) <= not (a xor b);
    layer2_outputs(3739) <= a;
    layer2_outputs(3740) <= not a or b;
    layer2_outputs(3741) <= not a;
    layer2_outputs(3742) <= a xor b;
    layer2_outputs(3743) <= a xor b;
    layer2_outputs(3744) <= not (a xor b);
    layer2_outputs(3745) <= not b;
    layer2_outputs(3746) <= a or b;
    layer2_outputs(3747) <= not b;
    layer2_outputs(3748) <= not b;
    layer2_outputs(3749) <= not a;
    layer2_outputs(3750) <= not a or b;
    layer2_outputs(3751) <= not (a and b);
    layer2_outputs(3752) <= not b or a;
    layer2_outputs(3753) <= a xor b;
    layer2_outputs(3754) <= not a;
    layer2_outputs(3755) <= b;
    layer2_outputs(3756) <= not b;
    layer2_outputs(3757) <= not a;
    layer2_outputs(3758) <= not (a or b);
    layer2_outputs(3759) <= not (a or b);
    layer2_outputs(3760) <= not (a xor b);
    layer2_outputs(3761) <= a and b;
    layer2_outputs(3762) <= a and not b;
    layer2_outputs(3763) <= a or b;
    layer2_outputs(3764) <= a;
    layer2_outputs(3765) <= a;
    layer2_outputs(3766) <= b and not a;
    layer2_outputs(3767) <= a xor b;
    layer2_outputs(3768) <= not (a and b);
    layer2_outputs(3769) <= b and not a;
    layer2_outputs(3770) <= not b;
    layer2_outputs(3771) <= not a;
    layer2_outputs(3772) <= not (a xor b);
    layer2_outputs(3773) <= not b or a;
    layer2_outputs(3774) <= not a;
    layer2_outputs(3775) <= not b;
    layer2_outputs(3776) <= not b or a;
    layer2_outputs(3777) <= a and b;
    layer2_outputs(3778) <= not (a and b);
    layer2_outputs(3779) <= not b or a;
    layer2_outputs(3780) <= not (a xor b);
    layer2_outputs(3781) <= not (a xor b);
    layer2_outputs(3782) <= a;
    layer2_outputs(3783) <= a xor b;
    layer2_outputs(3784) <= a and not b;
    layer2_outputs(3785) <= a xor b;
    layer2_outputs(3786) <= a;
    layer2_outputs(3787) <= a xor b;
    layer2_outputs(3788) <= b;
    layer2_outputs(3789) <= b;
    layer2_outputs(3790) <= a xor b;
    layer2_outputs(3791) <= b;
    layer2_outputs(3792) <= not b;
    layer2_outputs(3793) <= a;
    layer2_outputs(3794) <= not (a xor b);
    layer2_outputs(3795) <= not a;
    layer2_outputs(3796) <= a;
    layer2_outputs(3797) <= not b;
    layer2_outputs(3798) <= not (a xor b);
    layer2_outputs(3799) <= a or b;
    layer2_outputs(3800) <= not b;
    layer2_outputs(3801) <= a;
    layer2_outputs(3802) <= not b;
    layer2_outputs(3803) <= not (a and b);
    layer2_outputs(3804) <= not a or b;
    layer2_outputs(3805) <= not b or a;
    layer2_outputs(3806) <= not b or a;
    layer2_outputs(3807) <= b;
    layer2_outputs(3808) <= a;
    layer2_outputs(3809) <= a or b;
    layer2_outputs(3810) <= not b;
    layer2_outputs(3811) <= a and not b;
    layer2_outputs(3812) <= not a;
    layer2_outputs(3813) <= not b or a;
    layer2_outputs(3814) <= not (a and b);
    layer2_outputs(3815) <= a;
    layer2_outputs(3816) <= not (a xor b);
    layer2_outputs(3817) <= b and not a;
    layer2_outputs(3818) <= a xor b;
    layer2_outputs(3819) <= not a or b;
    layer2_outputs(3820) <= not a;
    layer2_outputs(3821) <= not b;
    layer2_outputs(3822) <= not a;
    layer2_outputs(3823) <= b;
    layer2_outputs(3824) <= not (a and b);
    layer2_outputs(3825) <= a and b;
    layer2_outputs(3826) <= not a or b;
    layer2_outputs(3827) <= not (a xor b);
    layer2_outputs(3828) <= b;
    layer2_outputs(3829) <= a;
    layer2_outputs(3830) <= a and not b;
    layer2_outputs(3831) <= a xor b;
    layer2_outputs(3832) <= a xor b;
    layer2_outputs(3833) <= not b;
    layer2_outputs(3834) <= not (a xor b);
    layer2_outputs(3835) <= a;
    layer2_outputs(3836) <= a or b;
    layer2_outputs(3837) <= a xor b;
    layer2_outputs(3838) <= a xor b;
    layer2_outputs(3839) <= not b;
    layer2_outputs(3840) <= not b;
    layer2_outputs(3841) <= not a;
    layer2_outputs(3842) <= not b or a;
    layer2_outputs(3843) <= a or b;
    layer2_outputs(3844) <= not a or b;
    layer2_outputs(3845) <= a and b;
    layer2_outputs(3846) <= not (a and b);
    layer2_outputs(3847) <= a or b;
    layer2_outputs(3848) <= a;
    layer2_outputs(3849) <= not (a xor b);
    layer2_outputs(3850) <= not a;
    layer2_outputs(3851) <= a;
    layer2_outputs(3852) <= a xor b;
    layer2_outputs(3853) <= not b;
    layer2_outputs(3854) <= not b;
    layer2_outputs(3855) <= not a;
    layer2_outputs(3856) <= b and not a;
    layer2_outputs(3857) <= not (a and b);
    layer2_outputs(3858) <= not b;
    layer2_outputs(3859) <= not (a xor b);
    layer2_outputs(3860) <= not a;
    layer2_outputs(3861) <= b and not a;
    layer2_outputs(3862) <= a and b;
    layer2_outputs(3863) <= not b or a;
    layer2_outputs(3864) <= not b;
    layer2_outputs(3865) <= not (a or b);
    layer2_outputs(3866) <= not b;
    layer2_outputs(3867) <= b;
    layer2_outputs(3868) <= not a;
    layer2_outputs(3869) <= not b;
    layer2_outputs(3870) <= a xor b;
    layer2_outputs(3871) <= b;
    layer2_outputs(3872) <= a and b;
    layer2_outputs(3873) <= not (a xor b);
    layer2_outputs(3874) <= not (a xor b);
    layer2_outputs(3875) <= not b;
    layer2_outputs(3876) <= a or b;
    layer2_outputs(3877) <= not (a xor b);
    layer2_outputs(3878) <= not b or a;
    layer2_outputs(3879) <= a and b;
    layer2_outputs(3880) <= not a;
    layer2_outputs(3881) <= not a;
    layer2_outputs(3882) <= b and not a;
    layer2_outputs(3883) <= not a or b;
    layer2_outputs(3884) <= a xor b;
    layer2_outputs(3885) <= a xor b;
    layer2_outputs(3886) <= not a;
    layer2_outputs(3887) <= b;
    layer2_outputs(3888) <= a xor b;
    layer2_outputs(3889) <= not a;
    layer2_outputs(3890) <= b;
    layer2_outputs(3891) <= a;
    layer2_outputs(3892) <= a or b;
    layer2_outputs(3893) <= not b;
    layer2_outputs(3894) <= not (a xor b);
    layer2_outputs(3895) <= a or b;
    layer2_outputs(3896) <= not b or a;
    layer2_outputs(3897) <= a xor b;
    layer2_outputs(3898) <= a xor b;
    layer2_outputs(3899) <= not a or b;
    layer2_outputs(3900) <= a;
    layer2_outputs(3901) <= not (a xor b);
    layer2_outputs(3902) <= not b;
    layer2_outputs(3903) <= not (a xor b);
    layer2_outputs(3904) <= a;
    layer2_outputs(3905) <= not b;
    layer2_outputs(3906) <= not a;
    layer2_outputs(3907) <= not b;
    layer2_outputs(3908) <= b;
    layer2_outputs(3909) <= not (a or b);
    layer2_outputs(3910) <= a and b;
    layer2_outputs(3911) <= not (a xor b);
    layer2_outputs(3912) <= a;
    layer2_outputs(3913) <= not a;
    layer2_outputs(3914) <= a;
    layer2_outputs(3915) <= not b;
    layer2_outputs(3916) <= not (a and b);
    layer2_outputs(3917) <= a;
    layer2_outputs(3918) <= not (a and b);
    layer2_outputs(3919) <= not (a and b);
    layer2_outputs(3920) <= a;
    layer2_outputs(3921) <= not a;
    layer2_outputs(3922) <= not b;
    layer2_outputs(3923) <= not (a xor b);
    layer2_outputs(3924) <= not (a xor b);
    layer2_outputs(3925) <= not a;
    layer2_outputs(3926) <= not (a xor b);
    layer2_outputs(3927) <= not (a xor b);
    layer2_outputs(3928) <= not b;
    layer2_outputs(3929) <= a and b;
    layer2_outputs(3930) <= not b;
    layer2_outputs(3931) <= not (a xor b);
    layer2_outputs(3932) <= b;
    layer2_outputs(3933) <= not b;
    layer2_outputs(3934) <= b and not a;
    layer2_outputs(3935) <= not a;
    layer2_outputs(3936) <= not (a or b);
    layer2_outputs(3937) <= a;
    layer2_outputs(3938) <= not b or a;
    layer2_outputs(3939) <= not (a or b);
    layer2_outputs(3940) <= a or b;
    layer2_outputs(3941) <= 1'b1;
    layer2_outputs(3942) <= not b;
    layer2_outputs(3943) <= b;
    layer2_outputs(3944) <= not (a xor b);
    layer2_outputs(3945) <= a xor b;
    layer2_outputs(3946) <= not b or a;
    layer2_outputs(3947) <= a;
    layer2_outputs(3948) <= a and b;
    layer2_outputs(3949) <= not (a xor b);
    layer2_outputs(3950) <= not (a xor b);
    layer2_outputs(3951) <= not (a xor b);
    layer2_outputs(3952) <= b;
    layer2_outputs(3953) <= not (a or b);
    layer2_outputs(3954) <= not a or b;
    layer2_outputs(3955) <= not b or a;
    layer2_outputs(3956) <= a and b;
    layer2_outputs(3957) <= not b;
    layer2_outputs(3958) <= not b or a;
    layer2_outputs(3959) <= a and not b;
    layer2_outputs(3960) <= b;
    layer2_outputs(3961) <= not (a xor b);
    layer2_outputs(3962) <= a and b;
    layer2_outputs(3963) <= not a;
    layer2_outputs(3964) <= not (a xor b);
    layer2_outputs(3965) <= a or b;
    layer2_outputs(3966) <= b and not a;
    layer2_outputs(3967) <= b;
    layer2_outputs(3968) <= not (a xor b);
    layer2_outputs(3969) <= a and b;
    layer2_outputs(3970) <= b and not a;
    layer2_outputs(3971) <= a;
    layer2_outputs(3972) <= b;
    layer2_outputs(3973) <= not (a or b);
    layer2_outputs(3974) <= not a;
    layer2_outputs(3975) <= a;
    layer2_outputs(3976) <= a xor b;
    layer2_outputs(3977) <= not (a and b);
    layer2_outputs(3978) <= not b;
    layer2_outputs(3979) <= a and b;
    layer2_outputs(3980) <= b;
    layer2_outputs(3981) <= not b;
    layer2_outputs(3982) <= not (a or b);
    layer2_outputs(3983) <= a xor b;
    layer2_outputs(3984) <= not (a and b);
    layer2_outputs(3985) <= not a;
    layer2_outputs(3986) <= a xor b;
    layer2_outputs(3987) <= not b;
    layer2_outputs(3988) <= a xor b;
    layer2_outputs(3989) <= a and b;
    layer2_outputs(3990) <= not b;
    layer2_outputs(3991) <= not (a or b);
    layer2_outputs(3992) <= not b or a;
    layer2_outputs(3993) <= not (a xor b);
    layer2_outputs(3994) <= not a;
    layer2_outputs(3995) <= a and b;
    layer2_outputs(3996) <= not b or a;
    layer2_outputs(3997) <= not (a or b);
    layer2_outputs(3998) <= a or b;
    layer2_outputs(3999) <= b and not a;
    layer2_outputs(4000) <= not b;
    layer2_outputs(4001) <= a and not b;
    layer2_outputs(4002) <= not b;
    layer2_outputs(4003) <= not b or a;
    layer2_outputs(4004) <= not b or a;
    layer2_outputs(4005) <= not a;
    layer2_outputs(4006) <= a xor b;
    layer2_outputs(4007) <= not (a or b);
    layer2_outputs(4008) <= not b or a;
    layer2_outputs(4009) <= not (a or b);
    layer2_outputs(4010) <= not b;
    layer2_outputs(4011) <= not b;
    layer2_outputs(4012) <= a and not b;
    layer2_outputs(4013) <= not a;
    layer2_outputs(4014) <= not (a and b);
    layer2_outputs(4015) <= b;
    layer2_outputs(4016) <= a and b;
    layer2_outputs(4017) <= a xor b;
    layer2_outputs(4018) <= not b;
    layer2_outputs(4019) <= not (a xor b);
    layer2_outputs(4020) <= not (a and b);
    layer2_outputs(4021) <= b and not a;
    layer2_outputs(4022) <= not b;
    layer2_outputs(4023) <= a xor b;
    layer2_outputs(4024) <= not b;
    layer2_outputs(4025) <= a and b;
    layer2_outputs(4026) <= not b;
    layer2_outputs(4027) <= b and not a;
    layer2_outputs(4028) <= b and not a;
    layer2_outputs(4029) <= not (a xor b);
    layer2_outputs(4030) <= a xor b;
    layer2_outputs(4031) <= a and not b;
    layer2_outputs(4032) <= a xor b;
    layer2_outputs(4033) <= a and not b;
    layer2_outputs(4034) <= not b;
    layer2_outputs(4035) <= not (a and b);
    layer2_outputs(4036) <= b and not a;
    layer2_outputs(4037) <= not (a and b);
    layer2_outputs(4038) <= not b;
    layer2_outputs(4039) <= not b;
    layer2_outputs(4040) <= not a;
    layer2_outputs(4041) <= b;
    layer2_outputs(4042) <= a or b;
    layer2_outputs(4043) <= not a;
    layer2_outputs(4044) <= a or b;
    layer2_outputs(4045) <= not b;
    layer2_outputs(4046) <= not b;
    layer2_outputs(4047) <= a;
    layer2_outputs(4048) <= b;
    layer2_outputs(4049) <= not (a or b);
    layer2_outputs(4050) <= not (a and b);
    layer2_outputs(4051) <= b and not a;
    layer2_outputs(4052) <= not b;
    layer2_outputs(4053) <= b;
    layer2_outputs(4054) <= a;
    layer2_outputs(4055) <= a and b;
    layer2_outputs(4056) <= a and not b;
    layer2_outputs(4057) <= a;
    layer2_outputs(4058) <= not (a xor b);
    layer2_outputs(4059) <= not b or a;
    layer2_outputs(4060) <= a and b;
    layer2_outputs(4061) <= a;
    layer2_outputs(4062) <= a and not b;
    layer2_outputs(4063) <= not b or a;
    layer2_outputs(4064) <= b;
    layer2_outputs(4065) <= not b or a;
    layer2_outputs(4066) <= a xor b;
    layer2_outputs(4067) <= a;
    layer2_outputs(4068) <= b and not a;
    layer2_outputs(4069) <= not a;
    layer2_outputs(4070) <= not (a xor b);
    layer2_outputs(4071) <= not (a or b);
    layer2_outputs(4072) <= not (a xor b);
    layer2_outputs(4073) <= b;
    layer2_outputs(4074) <= b;
    layer2_outputs(4075) <= not (a xor b);
    layer2_outputs(4076) <= not a;
    layer2_outputs(4077) <= a and b;
    layer2_outputs(4078) <= not b or a;
    layer2_outputs(4079) <= a and not b;
    layer2_outputs(4080) <= b and not a;
    layer2_outputs(4081) <= a or b;
    layer2_outputs(4082) <= not (a xor b);
    layer2_outputs(4083) <= b;
    layer2_outputs(4084) <= b and not a;
    layer2_outputs(4085) <= a or b;
    layer2_outputs(4086) <= not (a and b);
    layer2_outputs(4087) <= a and b;
    layer2_outputs(4088) <= not a;
    layer2_outputs(4089) <= b;
    layer2_outputs(4090) <= a xor b;
    layer2_outputs(4091) <= not (a and b);
    layer2_outputs(4092) <= not b;
    layer2_outputs(4093) <= not a;
    layer2_outputs(4094) <= 1'b0;
    layer2_outputs(4095) <= a;
    layer2_outputs(4096) <= b;
    layer2_outputs(4097) <= a xor b;
    layer2_outputs(4098) <= b;
    layer2_outputs(4099) <= b and not a;
    layer2_outputs(4100) <= not a;
    layer2_outputs(4101) <= a and not b;
    layer2_outputs(4102) <= not b or a;
    layer2_outputs(4103) <= not a;
    layer2_outputs(4104) <= b and not a;
    layer2_outputs(4105) <= b;
    layer2_outputs(4106) <= a;
    layer2_outputs(4107) <= a xor b;
    layer2_outputs(4108) <= not b;
    layer2_outputs(4109) <= not (a or b);
    layer2_outputs(4110) <= not a;
    layer2_outputs(4111) <= not (a xor b);
    layer2_outputs(4112) <= not b;
    layer2_outputs(4113) <= not b;
    layer2_outputs(4114) <= not (a or b);
    layer2_outputs(4115) <= a and b;
    layer2_outputs(4116) <= a and not b;
    layer2_outputs(4117) <= a xor b;
    layer2_outputs(4118) <= a;
    layer2_outputs(4119) <= not b;
    layer2_outputs(4120) <= b;
    layer2_outputs(4121) <= not a;
    layer2_outputs(4122) <= not a;
    layer2_outputs(4123) <= a and b;
    layer2_outputs(4124) <= a and not b;
    layer2_outputs(4125) <= a and not b;
    layer2_outputs(4126) <= b and not a;
    layer2_outputs(4127) <= not a;
    layer2_outputs(4128) <= not b;
    layer2_outputs(4129) <= not a;
    layer2_outputs(4130) <= b;
    layer2_outputs(4131) <= not b;
    layer2_outputs(4132) <= not b;
    layer2_outputs(4133) <= not a;
    layer2_outputs(4134) <= not (a and b);
    layer2_outputs(4135) <= a xor b;
    layer2_outputs(4136) <= not (a xor b);
    layer2_outputs(4137) <= a;
    layer2_outputs(4138) <= a xor b;
    layer2_outputs(4139) <= b;
    layer2_outputs(4140) <= not a;
    layer2_outputs(4141) <= a xor b;
    layer2_outputs(4142) <= not (a xor b);
    layer2_outputs(4143) <= a or b;
    layer2_outputs(4144) <= a xor b;
    layer2_outputs(4145) <= b and not a;
    layer2_outputs(4146) <= not (a xor b);
    layer2_outputs(4147) <= not (a xor b);
    layer2_outputs(4148) <= not a or b;
    layer2_outputs(4149) <= a;
    layer2_outputs(4150) <= 1'b1;
    layer2_outputs(4151) <= a and not b;
    layer2_outputs(4152) <= a xor b;
    layer2_outputs(4153) <= a;
    layer2_outputs(4154) <= a or b;
    layer2_outputs(4155) <= not a;
    layer2_outputs(4156) <= b;
    layer2_outputs(4157) <= not b;
    layer2_outputs(4158) <= a and not b;
    layer2_outputs(4159) <= b and not a;
    layer2_outputs(4160) <= not b;
    layer2_outputs(4161) <= not a;
    layer2_outputs(4162) <= b;
    layer2_outputs(4163) <= not (a or b);
    layer2_outputs(4164) <= not (a or b);
    layer2_outputs(4165) <= b;
    layer2_outputs(4166) <= b;
    layer2_outputs(4167) <= not a or b;
    layer2_outputs(4168) <= a xor b;
    layer2_outputs(4169) <= a and b;
    layer2_outputs(4170) <= b and not a;
    layer2_outputs(4171) <= not (a or b);
    layer2_outputs(4172) <= b;
    layer2_outputs(4173) <= b;
    layer2_outputs(4174) <= b;
    layer2_outputs(4175) <= not (a or b);
    layer2_outputs(4176) <= not a;
    layer2_outputs(4177) <= b;
    layer2_outputs(4178) <= not (a and b);
    layer2_outputs(4179) <= not a or b;
    layer2_outputs(4180) <= not b;
    layer2_outputs(4181) <= not b;
    layer2_outputs(4182) <= b;
    layer2_outputs(4183) <= not (a and b);
    layer2_outputs(4184) <= a xor b;
    layer2_outputs(4185) <= not b or a;
    layer2_outputs(4186) <= a;
    layer2_outputs(4187) <= b;
    layer2_outputs(4188) <= not b or a;
    layer2_outputs(4189) <= not a or b;
    layer2_outputs(4190) <= b;
    layer2_outputs(4191) <= not (a and b);
    layer2_outputs(4192) <= a or b;
    layer2_outputs(4193) <= a xor b;
    layer2_outputs(4194) <= a xor b;
    layer2_outputs(4195) <= a;
    layer2_outputs(4196) <= not b or a;
    layer2_outputs(4197) <= a and not b;
    layer2_outputs(4198) <= a or b;
    layer2_outputs(4199) <= a xor b;
    layer2_outputs(4200) <= b;
    layer2_outputs(4201) <= not a;
    layer2_outputs(4202) <= a and b;
    layer2_outputs(4203) <= b and not a;
    layer2_outputs(4204) <= not a;
    layer2_outputs(4205) <= a xor b;
    layer2_outputs(4206) <= not a;
    layer2_outputs(4207) <= b;
    layer2_outputs(4208) <= b;
    layer2_outputs(4209) <= not (a or b);
    layer2_outputs(4210) <= a xor b;
    layer2_outputs(4211) <= a and b;
    layer2_outputs(4212) <= a;
    layer2_outputs(4213) <= a and b;
    layer2_outputs(4214) <= not (a xor b);
    layer2_outputs(4215) <= not b;
    layer2_outputs(4216) <= b and not a;
    layer2_outputs(4217) <= not b;
    layer2_outputs(4218) <= not a or b;
    layer2_outputs(4219) <= a and b;
    layer2_outputs(4220) <= a and not b;
    layer2_outputs(4221) <= not (a and b);
    layer2_outputs(4222) <= a xor b;
    layer2_outputs(4223) <= a and not b;
    layer2_outputs(4224) <= not (a and b);
    layer2_outputs(4225) <= not (a xor b);
    layer2_outputs(4226) <= b;
    layer2_outputs(4227) <= a;
    layer2_outputs(4228) <= a and b;
    layer2_outputs(4229) <= not a;
    layer2_outputs(4230) <= b;
    layer2_outputs(4231) <= a or b;
    layer2_outputs(4232) <= a and not b;
    layer2_outputs(4233) <= not (a xor b);
    layer2_outputs(4234) <= not (a and b);
    layer2_outputs(4235) <= not (a xor b);
    layer2_outputs(4236) <= b;
    layer2_outputs(4237) <= not b;
    layer2_outputs(4238) <= b;
    layer2_outputs(4239) <= not a or b;
    layer2_outputs(4240) <= not (a or b);
    layer2_outputs(4241) <= a xor b;
    layer2_outputs(4242) <= a;
    layer2_outputs(4243) <= a;
    layer2_outputs(4244) <= a and b;
    layer2_outputs(4245) <= not (a xor b);
    layer2_outputs(4246) <= not b or a;
    layer2_outputs(4247) <= a;
    layer2_outputs(4248) <= b and not a;
    layer2_outputs(4249) <= a;
    layer2_outputs(4250) <= not (a xor b);
    layer2_outputs(4251) <= a xor b;
    layer2_outputs(4252) <= a;
    layer2_outputs(4253) <= 1'b0;
    layer2_outputs(4254) <= not (a and b);
    layer2_outputs(4255) <= a;
    layer2_outputs(4256) <= not a;
    layer2_outputs(4257) <= a xor b;
    layer2_outputs(4258) <= a or b;
    layer2_outputs(4259) <= a or b;
    layer2_outputs(4260) <= not a or b;
    layer2_outputs(4261) <= a;
    layer2_outputs(4262) <= a and b;
    layer2_outputs(4263) <= b and not a;
    layer2_outputs(4264) <= a or b;
    layer2_outputs(4265) <= b;
    layer2_outputs(4266) <= b;
    layer2_outputs(4267) <= not (a xor b);
    layer2_outputs(4268) <= a and b;
    layer2_outputs(4269) <= not b;
    layer2_outputs(4270) <= a or b;
    layer2_outputs(4271) <= not b;
    layer2_outputs(4272) <= not a;
    layer2_outputs(4273) <= not a or b;
    layer2_outputs(4274) <= not b or a;
    layer2_outputs(4275) <= b;
    layer2_outputs(4276) <= a and b;
    layer2_outputs(4277) <= a and b;
    layer2_outputs(4278) <= not b or a;
    layer2_outputs(4279) <= not (a xor b);
    layer2_outputs(4280) <= a xor b;
    layer2_outputs(4281) <= not (a or b);
    layer2_outputs(4282) <= not a or b;
    layer2_outputs(4283) <= a;
    layer2_outputs(4284) <= a;
    layer2_outputs(4285) <= a and b;
    layer2_outputs(4286) <= a and not b;
    layer2_outputs(4287) <= not b;
    layer2_outputs(4288) <= a and b;
    layer2_outputs(4289) <= a and not b;
    layer2_outputs(4290) <= 1'b1;
    layer2_outputs(4291) <= not a or b;
    layer2_outputs(4292) <= not a;
    layer2_outputs(4293) <= not (a and b);
    layer2_outputs(4294) <= not b;
    layer2_outputs(4295) <= a xor b;
    layer2_outputs(4296) <= a and not b;
    layer2_outputs(4297) <= not (a and b);
    layer2_outputs(4298) <= not a;
    layer2_outputs(4299) <= not (a xor b);
    layer2_outputs(4300) <= a;
    layer2_outputs(4301) <= not b;
    layer2_outputs(4302) <= b and not a;
    layer2_outputs(4303) <= a xor b;
    layer2_outputs(4304) <= a xor b;
    layer2_outputs(4305) <= not b;
    layer2_outputs(4306) <= not b;
    layer2_outputs(4307) <= a;
    layer2_outputs(4308) <= not b;
    layer2_outputs(4309) <= not b;
    layer2_outputs(4310) <= not a or b;
    layer2_outputs(4311) <= a and b;
    layer2_outputs(4312) <= b;
    layer2_outputs(4313) <= not a;
    layer2_outputs(4314) <= a or b;
    layer2_outputs(4315) <= not a;
    layer2_outputs(4316) <= a xor b;
    layer2_outputs(4317) <= a xor b;
    layer2_outputs(4318) <= a xor b;
    layer2_outputs(4319) <= a and b;
    layer2_outputs(4320) <= not (a or b);
    layer2_outputs(4321) <= not b or a;
    layer2_outputs(4322) <= not (a and b);
    layer2_outputs(4323) <= not b;
    layer2_outputs(4324) <= b;
    layer2_outputs(4325) <= a;
    layer2_outputs(4326) <= a xor b;
    layer2_outputs(4327) <= not a;
    layer2_outputs(4328) <= a and not b;
    layer2_outputs(4329) <= not (a and b);
    layer2_outputs(4330) <= a;
    layer2_outputs(4331) <= a and b;
    layer2_outputs(4332) <= not b;
    layer2_outputs(4333) <= a;
    layer2_outputs(4334) <= not b or a;
    layer2_outputs(4335) <= not a or b;
    layer2_outputs(4336) <= a;
    layer2_outputs(4337) <= a and b;
    layer2_outputs(4338) <= a;
    layer2_outputs(4339) <= not (a xor b);
    layer2_outputs(4340) <= not b;
    layer2_outputs(4341) <= not (a xor b);
    layer2_outputs(4342) <= a xor b;
    layer2_outputs(4343) <= not b;
    layer2_outputs(4344) <= not a or b;
    layer2_outputs(4345) <= not b;
    layer2_outputs(4346) <= a or b;
    layer2_outputs(4347) <= not a;
    layer2_outputs(4348) <= a and not b;
    layer2_outputs(4349) <= a;
    layer2_outputs(4350) <= b;
    layer2_outputs(4351) <= not a;
    layer2_outputs(4352) <= a and not b;
    layer2_outputs(4353) <= a;
    layer2_outputs(4354) <= a and not b;
    layer2_outputs(4355) <= a;
    layer2_outputs(4356) <= not b;
    layer2_outputs(4357) <= not b;
    layer2_outputs(4358) <= not b;
    layer2_outputs(4359) <= not a or b;
    layer2_outputs(4360) <= not b;
    layer2_outputs(4361) <= a and b;
    layer2_outputs(4362) <= not b or a;
    layer2_outputs(4363) <= a xor b;
    layer2_outputs(4364) <= a and not b;
    layer2_outputs(4365) <= a;
    layer2_outputs(4366) <= 1'b1;
    layer2_outputs(4367) <= b;
    layer2_outputs(4368) <= not b;
    layer2_outputs(4369) <= not b;
    layer2_outputs(4370) <= not a or b;
    layer2_outputs(4371) <= not a or b;
    layer2_outputs(4372) <= not a or b;
    layer2_outputs(4373) <= a;
    layer2_outputs(4374) <= not (a and b);
    layer2_outputs(4375) <= a and b;
    layer2_outputs(4376) <= a and b;
    layer2_outputs(4377) <= a and not b;
    layer2_outputs(4378) <= a;
    layer2_outputs(4379) <= a;
    layer2_outputs(4380) <= not b or a;
    layer2_outputs(4381) <= not (a xor b);
    layer2_outputs(4382) <= b and not a;
    layer2_outputs(4383) <= not (a xor b);
    layer2_outputs(4384) <= a;
    layer2_outputs(4385) <= not b;
    layer2_outputs(4386) <= a;
    layer2_outputs(4387) <= not a;
    layer2_outputs(4388) <= b;
    layer2_outputs(4389) <= a and b;
    layer2_outputs(4390) <= a;
    layer2_outputs(4391) <= b and not a;
    layer2_outputs(4392) <= not (a xor b);
    layer2_outputs(4393) <= not b;
    layer2_outputs(4394) <= not (a xor b);
    layer2_outputs(4395) <= b;
    layer2_outputs(4396) <= a;
    layer2_outputs(4397) <= a or b;
    layer2_outputs(4398) <= a;
    layer2_outputs(4399) <= b;
    layer2_outputs(4400) <= a and b;
    layer2_outputs(4401) <= a xor b;
    layer2_outputs(4402) <= a xor b;
    layer2_outputs(4403) <= not (a xor b);
    layer2_outputs(4404) <= not (a and b);
    layer2_outputs(4405) <= not b or a;
    layer2_outputs(4406) <= a;
    layer2_outputs(4407) <= not b;
    layer2_outputs(4408) <= not (a xor b);
    layer2_outputs(4409) <= not a;
    layer2_outputs(4410) <= a xor b;
    layer2_outputs(4411) <= not b;
    layer2_outputs(4412) <= b and not a;
    layer2_outputs(4413) <= a xor b;
    layer2_outputs(4414) <= not a;
    layer2_outputs(4415) <= not a;
    layer2_outputs(4416) <= a;
    layer2_outputs(4417) <= a xor b;
    layer2_outputs(4418) <= not b or a;
    layer2_outputs(4419) <= b;
    layer2_outputs(4420) <= b;
    layer2_outputs(4421) <= not a;
    layer2_outputs(4422) <= not b;
    layer2_outputs(4423) <= b and not a;
    layer2_outputs(4424) <= not a or b;
    layer2_outputs(4425) <= a or b;
    layer2_outputs(4426) <= not a;
    layer2_outputs(4427) <= b;
    layer2_outputs(4428) <= not (a or b);
    layer2_outputs(4429) <= not (a and b);
    layer2_outputs(4430) <= b;
    layer2_outputs(4431) <= a;
    layer2_outputs(4432) <= a;
    layer2_outputs(4433) <= b;
    layer2_outputs(4434) <= not (a and b);
    layer2_outputs(4435) <= b;
    layer2_outputs(4436) <= a;
    layer2_outputs(4437) <= not (a xor b);
    layer2_outputs(4438) <= not a;
    layer2_outputs(4439) <= b and not a;
    layer2_outputs(4440) <= not b or a;
    layer2_outputs(4441) <= b;
    layer2_outputs(4442) <= not (a or b);
    layer2_outputs(4443) <= b;
    layer2_outputs(4444) <= not (a or b);
    layer2_outputs(4445) <= a xor b;
    layer2_outputs(4446) <= b;
    layer2_outputs(4447) <= not b or a;
    layer2_outputs(4448) <= not b;
    layer2_outputs(4449) <= not b;
    layer2_outputs(4450) <= a or b;
    layer2_outputs(4451) <= not a;
    layer2_outputs(4452) <= not a;
    layer2_outputs(4453) <= not a;
    layer2_outputs(4454) <= a;
    layer2_outputs(4455) <= a;
    layer2_outputs(4456) <= a;
    layer2_outputs(4457) <= b;
    layer2_outputs(4458) <= not b or a;
    layer2_outputs(4459) <= 1'b0;
    layer2_outputs(4460) <= not b;
    layer2_outputs(4461) <= not b or a;
    layer2_outputs(4462) <= not a;
    layer2_outputs(4463) <= not b;
    layer2_outputs(4464) <= a;
    layer2_outputs(4465) <= a xor b;
    layer2_outputs(4466) <= not (a and b);
    layer2_outputs(4467) <= not (a xor b);
    layer2_outputs(4468) <= not a or b;
    layer2_outputs(4469) <= not a;
    layer2_outputs(4470) <= not b;
    layer2_outputs(4471) <= a or b;
    layer2_outputs(4472) <= not a;
    layer2_outputs(4473) <= a xor b;
    layer2_outputs(4474) <= b;
    layer2_outputs(4475) <= not (a or b);
    layer2_outputs(4476) <= a and b;
    layer2_outputs(4477) <= not (a xor b);
    layer2_outputs(4478) <= not a or b;
    layer2_outputs(4479) <= a;
    layer2_outputs(4480) <= b and not a;
    layer2_outputs(4481) <= not b;
    layer2_outputs(4482) <= b;
    layer2_outputs(4483) <= b and not a;
    layer2_outputs(4484) <= not (a and b);
    layer2_outputs(4485) <= not (a or b);
    layer2_outputs(4486) <= not b or a;
    layer2_outputs(4487) <= a and b;
    layer2_outputs(4488) <= not a;
    layer2_outputs(4489) <= b;
    layer2_outputs(4490) <= not a;
    layer2_outputs(4491) <= not a or b;
    layer2_outputs(4492) <= a;
    layer2_outputs(4493) <= not (a and b);
    layer2_outputs(4494) <= a and not b;
    layer2_outputs(4495) <= b;
    layer2_outputs(4496) <= not b;
    layer2_outputs(4497) <= not (a xor b);
    layer2_outputs(4498) <= a and b;
    layer2_outputs(4499) <= a or b;
    layer2_outputs(4500) <= not a or b;
    layer2_outputs(4501) <= not a;
    layer2_outputs(4502) <= not a;
    layer2_outputs(4503) <= not a or b;
    layer2_outputs(4504) <= not (a xor b);
    layer2_outputs(4505) <= not (a xor b);
    layer2_outputs(4506) <= b;
    layer2_outputs(4507) <= not a;
    layer2_outputs(4508) <= not a;
    layer2_outputs(4509) <= not a;
    layer2_outputs(4510) <= a;
    layer2_outputs(4511) <= not (a and b);
    layer2_outputs(4512) <= a xor b;
    layer2_outputs(4513) <= a and not b;
    layer2_outputs(4514) <= a xor b;
    layer2_outputs(4515) <= not b or a;
    layer2_outputs(4516) <= not a;
    layer2_outputs(4517) <= a or b;
    layer2_outputs(4518) <= not b or a;
    layer2_outputs(4519) <= a xor b;
    layer2_outputs(4520) <= a and not b;
    layer2_outputs(4521) <= not a;
    layer2_outputs(4522) <= a and b;
    layer2_outputs(4523) <= a;
    layer2_outputs(4524) <= not b or a;
    layer2_outputs(4525) <= not a;
    layer2_outputs(4526) <= a;
    layer2_outputs(4527) <= a;
    layer2_outputs(4528) <= b;
    layer2_outputs(4529) <= b;
    layer2_outputs(4530) <= not a;
    layer2_outputs(4531) <= not (a xor b);
    layer2_outputs(4532) <= b;
    layer2_outputs(4533) <= a and not b;
    layer2_outputs(4534) <= b;
    layer2_outputs(4535) <= not a;
    layer2_outputs(4536) <= not (a or b);
    layer2_outputs(4537) <= a and b;
    layer2_outputs(4538) <= not (a and b);
    layer2_outputs(4539) <= not a or b;
    layer2_outputs(4540) <= not b;
    layer2_outputs(4541) <= not b;
    layer2_outputs(4542) <= a and b;
    layer2_outputs(4543) <= not b;
    layer2_outputs(4544) <= a xor b;
    layer2_outputs(4545) <= b;
    layer2_outputs(4546) <= not (a xor b);
    layer2_outputs(4547) <= a xor b;
    layer2_outputs(4548) <= not b;
    layer2_outputs(4549) <= not a or b;
    layer2_outputs(4550) <= not (a xor b);
    layer2_outputs(4551) <= not a;
    layer2_outputs(4552) <= not a;
    layer2_outputs(4553) <= not b;
    layer2_outputs(4554) <= b;
    layer2_outputs(4555) <= not (a or b);
    layer2_outputs(4556) <= a and not b;
    layer2_outputs(4557) <= b;
    layer2_outputs(4558) <= not b;
    layer2_outputs(4559) <= a;
    layer2_outputs(4560) <= a and not b;
    layer2_outputs(4561) <= not (a xor b);
    layer2_outputs(4562) <= a;
    layer2_outputs(4563) <= not (a and b);
    layer2_outputs(4564) <= not b or a;
    layer2_outputs(4565) <= a or b;
    layer2_outputs(4566) <= not b;
    layer2_outputs(4567) <= a xor b;
    layer2_outputs(4568) <= not a;
    layer2_outputs(4569) <= not (a xor b);
    layer2_outputs(4570) <= b;
    layer2_outputs(4571) <= b and not a;
    layer2_outputs(4572) <= not a;
    layer2_outputs(4573) <= not b;
    layer2_outputs(4574) <= a xor b;
    layer2_outputs(4575) <= not b or a;
    layer2_outputs(4576) <= a;
    layer2_outputs(4577) <= not (a and b);
    layer2_outputs(4578) <= not b;
    layer2_outputs(4579) <= not a;
    layer2_outputs(4580) <= not a;
    layer2_outputs(4581) <= not (a and b);
    layer2_outputs(4582) <= not b;
    layer2_outputs(4583) <= a and not b;
    layer2_outputs(4584) <= not (a and b);
    layer2_outputs(4585) <= b;
    layer2_outputs(4586) <= not (a xor b);
    layer2_outputs(4587) <= not a;
    layer2_outputs(4588) <= a xor b;
    layer2_outputs(4589) <= not a;
    layer2_outputs(4590) <= not b;
    layer2_outputs(4591) <= a and b;
    layer2_outputs(4592) <= not a or b;
    layer2_outputs(4593) <= a xor b;
    layer2_outputs(4594) <= not b or a;
    layer2_outputs(4595) <= a or b;
    layer2_outputs(4596) <= not b or a;
    layer2_outputs(4597) <= not a;
    layer2_outputs(4598) <= not a;
    layer2_outputs(4599) <= not (a xor b);
    layer2_outputs(4600) <= not (a or b);
    layer2_outputs(4601) <= a;
    layer2_outputs(4602) <= a;
    layer2_outputs(4603) <= a or b;
    layer2_outputs(4604) <= not a;
    layer2_outputs(4605) <= a and not b;
    layer2_outputs(4606) <= a;
    layer2_outputs(4607) <= not (a and b);
    layer2_outputs(4608) <= a and not b;
    layer2_outputs(4609) <= not b;
    layer2_outputs(4610) <= a;
    layer2_outputs(4611) <= not (a xor b);
    layer2_outputs(4612) <= not (a xor b);
    layer2_outputs(4613) <= a;
    layer2_outputs(4614) <= not a;
    layer2_outputs(4615) <= a;
    layer2_outputs(4616) <= a or b;
    layer2_outputs(4617) <= a;
    layer2_outputs(4618) <= a xor b;
    layer2_outputs(4619) <= not b;
    layer2_outputs(4620) <= b;
    layer2_outputs(4621) <= a;
    layer2_outputs(4622) <= b and not a;
    layer2_outputs(4623) <= not (a and b);
    layer2_outputs(4624) <= not (a or b);
    layer2_outputs(4625) <= not (a and b);
    layer2_outputs(4626) <= b;
    layer2_outputs(4627) <= not (a or b);
    layer2_outputs(4628) <= a and not b;
    layer2_outputs(4629) <= not (a and b);
    layer2_outputs(4630) <= not (a and b);
    layer2_outputs(4631) <= a or b;
    layer2_outputs(4632) <= not a;
    layer2_outputs(4633) <= a or b;
    layer2_outputs(4634) <= not a;
    layer2_outputs(4635) <= a;
    layer2_outputs(4636) <= b;
    layer2_outputs(4637) <= not b or a;
    layer2_outputs(4638) <= b and not a;
    layer2_outputs(4639) <= a xor b;
    layer2_outputs(4640) <= a or b;
    layer2_outputs(4641) <= not (a and b);
    layer2_outputs(4642) <= a or b;
    layer2_outputs(4643) <= a xor b;
    layer2_outputs(4644) <= not a;
    layer2_outputs(4645) <= a xor b;
    layer2_outputs(4646) <= b and not a;
    layer2_outputs(4647) <= not b or a;
    layer2_outputs(4648) <= b;
    layer2_outputs(4649) <= a and b;
    layer2_outputs(4650) <= b;
    layer2_outputs(4651) <= b;
    layer2_outputs(4652) <= b and not a;
    layer2_outputs(4653) <= not (a xor b);
    layer2_outputs(4654) <= not b;
    layer2_outputs(4655) <= not (a or b);
    layer2_outputs(4656) <= not b;
    layer2_outputs(4657) <= not b;
    layer2_outputs(4658) <= a and b;
    layer2_outputs(4659) <= not a;
    layer2_outputs(4660) <= not (a or b);
    layer2_outputs(4661) <= not b or a;
    layer2_outputs(4662) <= not (a xor b);
    layer2_outputs(4663) <= not a;
    layer2_outputs(4664) <= a and not b;
    layer2_outputs(4665) <= b;
    layer2_outputs(4666) <= not (a or b);
    layer2_outputs(4667) <= a xor b;
    layer2_outputs(4668) <= not (a xor b);
    layer2_outputs(4669) <= b and not a;
    layer2_outputs(4670) <= a;
    layer2_outputs(4671) <= a;
    layer2_outputs(4672) <= not b;
    layer2_outputs(4673) <= b;
    layer2_outputs(4674) <= a xor b;
    layer2_outputs(4675) <= a or b;
    layer2_outputs(4676) <= a xor b;
    layer2_outputs(4677) <= a and b;
    layer2_outputs(4678) <= not b or a;
    layer2_outputs(4679) <= not b;
    layer2_outputs(4680) <= a and b;
    layer2_outputs(4681) <= a and not b;
    layer2_outputs(4682) <= a or b;
    layer2_outputs(4683) <= b and not a;
    layer2_outputs(4684) <= a and not b;
    layer2_outputs(4685) <= not (a xor b);
    layer2_outputs(4686) <= not (a xor b);
    layer2_outputs(4687) <= not b;
    layer2_outputs(4688) <= not (a xor b);
    layer2_outputs(4689) <= a;
    layer2_outputs(4690) <= a and not b;
    layer2_outputs(4691) <= a and not b;
    layer2_outputs(4692) <= not b;
    layer2_outputs(4693) <= a xor b;
    layer2_outputs(4694) <= b;
    layer2_outputs(4695) <= not (a xor b);
    layer2_outputs(4696) <= a and not b;
    layer2_outputs(4697) <= not b;
    layer2_outputs(4698) <= not b or a;
    layer2_outputs(4699) <= a and b;
    layer2_outputs(4700) <= not (a xor b);
    layer2_outputs(4701) <= not a;
    layer2_outputs(4702) <= a or b;
    layer2_outputs(4703) <= a;
    layer2_outputs(4704) <= not b;
    layer2_outputs(4705) <= not a;
    layer2_outputs(4706) <= not b;
    layer2_outputs(4707) <= a xor b;
    layer2_outputs(4708) <= not b;
    layer2_outputs(4709) <= b;
    layer2_outputs(4710) <= b;
    layer2_outputs(4711) <= 1'b0;
    layer2_outputs(4712) <= b;
    layer2_outputs(4713) <= a;
    layer2_outputs(4714) <= b and not a;
    layer2_outputs(4715) <= b;
    layer2_outputs(4716) <= not a;
    layer2_outputs(4717) <= not (a or b);
    layer2_outputs(4718) <= a;
    layer2_outputs(4719) <= not a or b;
    layer2_outputs(4720) <= a xor b;
    layer2_outputs(4721) <= not (a or b);
    layer2_outputs(4722) <= a and b;
    layer2_outputs(4723) <= b and not a;
    layer2_outputs(4724) <= a and b;
    layer2_outputs(4725) <= not (a and b);
    layer2_outputs(4726) <= not (a or b);
    layer2_outputs(4727) <= not b;
    layer2_outputs(4728) <= not b;
    layer2_outputs(4729) <= a;
    layer2_outputs(4730) <= a and not b;
    layer2_outputs(4731) <= b and not a;
    layer2_outputs(4732) <= not b;
    layer2_outputs(4733) <= not a;
    layer2_outputs(4734) <= a and not b;
    layer2_outputs(4735) <= b and not a;
    layer2_outputs(4736) <= not b;
    layer2_outputs(4737) <= not (a and b);
    layer2_outputs(4738) <= b and not a;
    layer2_outputs(4739) <= a or b;
    layer2_outputs(4740) <= not (a or b);
    layer2_outputs(4741) <= not a;
    layer2_outputs(4742) <= not (a xor b);
    layer2_outputs(4743) <= not b;
    layer2_outputs(4744) <= not (a xor b);
    layer2_outputs(4745) <= not a;
    layer2_outputs(4746) <= b;
    layer2_outputs(4747) <= not (a xor b);
    layer2_outputs(4748) <= a or b;
    layer2_outputs(4749) <= b;
    layer2_outputs(4750) <= a xor b;
    layer2_outputs(4751) <= not b;
    layer2_outputs(4752) <= not a;
    layer2_outputs(4753) <= not b or a;
    layer2_outputs(4754) <= not b;
    layer2_outputs(4755) <= not (a xor b);
    layer2_outputs(4756) <= not a;
    layer2_outputs(4757) <= a xor b;
    layer2_outputs(4758) <= not (a or b);
    layer2_outputs(4759) <= not a;
    layer2_outputs(4760) <= not b;
    layer2_outputs(4761) <= a;
    layer2_outputs(4762) <= a and b;
    layer2_outputs(4763) <= b;
    layer2_outputs(4764) <= not b;
    layer2_outputs(4765) <= a xor b;
    layer2_outputs(4766) <= not b;
    layer2_outputs(4767) <= a;
    layer2_outputs(4768) <= not a or b;
    layer2_outputs(4769) <= not b or a;
    layer2_outputs(4770) <= not (a xor b);
    layer2_outputs(4771) <= not (a xor b);
    layer2_outputs(4772) <= not (a and b);
    layer2_outputs(4773) <= not b or a;
    layer2_outputs(4774) <= a;
    layer2_outputs(4775) <= a;
    layer2_outputs(4776) <= a and not b;
    layer2_outputs(4777) <= not b or a;
    layer2_outputs(4778) <= a xor b;
    layer2_outputs(4779) <= not a;
    layer2_outputs(4780) <= a and b;
    layer2_outputs(4781) <= a and not b;
    layer2_outputs(4782) <= not a;
    layer2_outputs(4783) <= not (a xor b);
    layer2_outputs(4784) <= a xor b;
    layer2_outputs(4785) <= not a;
    layer2_outputs(4786) <= not b;
    layer2_outputs(4787) <= a and not b;
    layer2_outputs(4788) <= a or b;
    layer2_outputs(4789) <= b and not a;
    layer2_outputs(4790) <= not (a and b);
    layer2_outputs(4791) <= b;
    layer2_outputs(4792) <= a and not b;
    layer2_outputs(4793) <= not (a and b);
    layer2_outputs(4794) <= a and b;
    layer2_outputs(4795) <= b;
    layer2_outputs(4796) <= a;
    layer2_outputs(4797) <= b;
    layer2_outputs(4798) <= not a or b;
    layer2_outputs(4799) <= a;
    layer2_outputs(4800) <= not b;
    layer2_outputs(4801) <= a;
    layer2_outputs(4802) <= not a;
    layer2_outputs(4803) <= b and not a;
    layer2_outputs(4804) <= not (a or b);
    layer2_outputs(4805) <= not a;
    layer2_outputs(4806) <= not (a xor b);
    layer2_outputs(4807) <= not a;
    layer2_outputs(4808) <= not a;
    layer2_outputs(4809) <= not (a xor b);
    layer2_outputs(4810) <= a or b;
    layer2_outputs(4811) <= b;
    layer2_outputs(4812) <= not b;
    layer2_outputs(4813) <= not a;
    layer2_outputs(4814) <= not (a xor b);
    layer2_outputs(4815) <= a;
    layer2_outputs(4816) <= not b or a;
    layer2_outputs(4817) <= not (a xor b);
    layer2_outputs(4818) <= not b;
    layer2_outputs(4819) <= b and not a;
    layer2_outputs(4820) <= not a;
    layer2_outputs(4821) <= b and not a;
    layer2_outputs(4822) <= a;
    layer2_outputs(4823) <= not b or a;
    layer2_outputs(4824) <= a;
    layer2_outputs(4825) <= not b or a;
    layer2_outputs(4826) <= a;
    layer2_outputs(4827) <= not a or b;
    layer2_outputs(4828) <= not b;
    layer2_outputs(4829) <= a or b;
    layer2_outputs(4830) <= not b;
    layer2_outputs(4831) <= not (a xor b);
    layer2_outputs(4832) <= not a or b;
    layer2_outputs(4833) <= not b;
    layer2_outputs(4834) <= not (a xor b);
    layer2_outputs(4835) <= a;
    layer2_outputs(4836) <= not (a or b);
    layer2_outputs(4837) <= a xor b;
    layer2_outputs(4838) <= not b;
    layer2_outputs(4839) <= not b;
    layer2_outputs(4840) <= not b or a;
    layer2_outputs(4841) <= a and not b;
    layer2_outputs(4842) <= not (a and b);
    layer2_outputs(4843) <= b and not a;
    layer2_outputs(4844) <= a;
    layer2_outputs(4845) <= not b;
    layer2_outputs(4846) <= not (a xor b);
    layer2_outputs(4847) <= b and not a;
    layer2_outputs(4848) <= a;
    layer2_outputs(4849) <= a xor b;
    layer2_outputs(4850) <= b;
    layer2_outputs(4851) <= b and not a;
    layer2_outputs(4852) <= a and b;
    layer2_outputs(4853) <= not (a or b);
    layer2_outputs(4854) <= not b;
    layer2_outputs(4855) <= a;
    layer2_outputs(4856) <= not a;
    layer2_outputs(4857) <= a;
    layer2_outputs(4858) <= a xor b;
    layer2_outputs(4859) <= not (a and b);
    layer2_outputs(4860) <= not b;
    layer2_outputs(4861) <= b;
    layer2_outputs(4862) <= not (a and b);
    layer2_outputs(4863) <= not b;
    layer2_outputs(4864) <= not b;
    layer2_outputs(4865) <= not b;
    layer2_outputs(4866) <= b and not a;
    layer2_outputs(4867) <= a;
    layer2_outputs(4868) <= a and not b;
    layer2_outputs(4869) <= not b;
    layer2_outputs(4870) <= b;
    layer2_outputs(4871) <= not a;
    layer2_outputs(4872) <= not (a xor b);
    layer2_outputs(4873) <= not a or b;
    layer2_outputs(4874) <= a xor b;
    layer2_outputs(4875) <= not a;
    layer2_outputs(4876) <= 1'b0;
    layer2_outputs(4877) <= a xor b;
    layer2_outputs(4878) <= not a;
    layer2_outputs(4879) <= not b;
    layer2_outputs(4880) <= a xor b;
    layer2_outputs(4881) <= not a or b;
    layer2_outputs(4882) <= not (a xor b);
    layer2_outputs(4883) <= a xor b;
    layer2_outputs(4884) <= not b;
    layer2_outputs(4885) <= a xor b;
    layer2_outputs(4886) <= b;
    layer2_outputs(4887) <= not (a xor b);
    layer2_outputs(4888) <= not b or a;
    layer2_outputs(4889) <= not (a xor b);
    layer2_outputs(4890) <= not b;
    layer2_outputs(4891) <= b;
    layer2_outputs(4892) <= not b or a;
    layer2_outputs(4893) <= not (a or b);
    layer2_outputs(4894) <= not (a and b);
    layer2_outputs(4895) <= a and b;
    layer2_outputs(4896) <= not (a or b);
    layer2_outputs(4897) <= not b;
    layer2_outputs(4898) <= a;
    layer2_outputs(4899) <= a or b;
    layer2_outputs(4900) <= not a;
    layer2_outputs(4901) <= not b;
    layer2_outputs(4902) <= not a or b;
    layer2_outputs(4903) <= not (a or b);
    layer2_outputs(4904) <= not b;
    layer2_outputs(4905) <= a or b;
    layer2_outputs(4906) <= a and b;
    layer2_outputs(4907) <= not a;
    layer2_outputs(4908) <= not a;
    layer2_outputs(4909) <= not (a or b);
    layer2_outputs(4910) <= a xor b;
    layer2_outputs(4911) <= a xor b;
    layer2_outputs(4912) <= not (a xor b);
    layer2_outputs(4913) <= b;
    layer2_outputs(4914) <= a xor b;
    layer2_outputs(4915) <= b;
    layer2_outputs(4916) <= a;
    layer2_outputs(4917) <= a or b;
    layer2_outputs(4918) <= not (a xor b);
    layer2_outputs(4919) <= a and not b;
    layer2_outputs(4920) <= a;
    layer2_outputs(4921) <= a xor b;
    layer2_outputs(4922) <= not (a xor b);
    layer2_outputs(4923) <= b;
    layer2_outputs(4924) <= a xor b;
    layer2_outputs(4925) <= b;
    layer2_outputs(4926) <= not a;
    layer2_outputs(4927) <= a xor b;
    layer2_outputs(4928) <= not (a xor b);
    layer2_outputs(4929) <= b;
    layer2_outputs(4930) <= not b or a;
    layer2_outputs(4931) <= a xor b;
    layer2_outputs(4932) <= b;
    layer2_outputs(4933) <= not (a or b);
    layer2_outputs(4934) <= a;
    layer2_outputs(4935) <= a xor b;
    layer2_outputs(4936) <= not (a xor b);
    layer2_outputs(4937) <= a xor b;
    layer2_outputs(4938) <= not a or b;
    layer2_outputs(4939) <= b;
    layer2_outputs(4940) <= not (a xor b);
    layer2_outputs(4941) <= not b or a;
    layer2_outputs(4942) <= a xor b;
    layer2_outputs(4943) <= not (a or b);
    layer2_outputs(4944) <= not a;
    layer2_outputs(4945) <= a and not b;
    layer2_outputs(4946) <= not (a or b);
    layer2_outputs(4947) <= a and b;
    layer2_outputs(4948) <= a;
    layer2_outputs(4949) <= b and not a;
    layer2_outputs(4950) <= b;
    layer2_outputs(4951) <= not (a xor b);
    layer2_outputs(4952) <= b and not a;
    layer2_outputs(4953) <= not a;
    layer2_outputs(4954) <= a and not b;
    layer2_outputs(4955) <= b and not a;
    layer2_outputs(4956) <= not (a xor b);
    layer2_outputs(4957) <= a xor b;
    layer2_outputs(4958) <= not (a xor b);
    layer2_outputs(4959) <= a;
    layer2_outputs(4960) <= not (a or b);
    layer2_outputs(4961) <= not a;
    layer2_outputs(4962) <= not a;
    layer2_outputs(4963) <= not (a xor b);
    layer2_outputs(4964) <= b;
    layer2_outputs(4965) <= b and not a;
    layer2_outputs(4966) <= not (a and b);
    layer2_outputs(4967) <= b;
    layer2_outputs(4968) <= not (a and b);
    layer2_outputs(4969) <= b;
    layer2_outputs(4970) <= not a;
    layer2_outputs(4971) <= not a;
    layer2_outputs(4972) <= b and not a;
    layer2_outputs(4973) <= a or b;
    layer2_outputs(4974) <= b;
    layer2_outputs(4975) <= a and not b;
    layer2_outputs(4976) <= not a or b;
    layer2_outputs(4977) <= not b;
    layer2_outputs(4978) <= not b or a;
    layer2_outputs(4979) <= not b;
    layer2_outputs(4980) <= not b;
    layer2_outputs(4981) <= a;
    layer2_outputs(4982) <= b;
    layer2_outputs(4983) <= not b or a;
    layer2_outputs(4984) <= b and not a;
    layer2_outputs(4985) <= not a or b;
    layer2_outputs(4986) <= b;
    layer2_outputs(4987) <= a and not b;
    layer2_outputs(4988) <= b;
    layer2_outputs(4989) <= not a;
    layer2_outputs(4990) <= not b or a;
    layer2_outputs(4991) <= not (a and b);
    layer2_outputs(4992) <= b;
    layer2_outputs(4993) <= not b or a;
    layer2_outputs(4994) <= a;
    layer2_outputs(4995) <= not (a or b);
    layer2_outputs(4996) <= not (a or b);
    layer2_outputs(4997) <= a and not b;
    layer2_outputs(4998) <= not (a and b);
    layer2_outputs(4999) <= not (a and b);
    layer2_outputs(5000) <= not b;
    layer2_outputs(5001) <= a;
    layer2_outputs(5002) <= not b;
    layer2_outputs(5003) <= not (a xor b);
    layer2_outputs(5004) <= not (a xor b);
    layer2_outputs(5005) <= b;
    layer2_outputs(5006) <= not b or a;
    layer2_outputs(5007) <= a and b;
    layer2_outputs(5008) <= b;
    layer2_outputs(5009) <= not a;
    layer2_outputs(5010) <= b and not a;
    layer2_outputs(5011) <= not b or a;
    layer2_outputs(5012) <= not b or a;
    layer2_outputs(5013) <= a and not b;
    layer2_outputs(5014) <= a xor b;
    layer2_outputs(5015) <= not b or a;
    layer2_outputs(5016) <= a;
    layer2_outputs(5017) <= b;
    layer2_outputs(5018) <= a or b;
    layer2_outputs(5019) <= a;
    layer2_outputs(5020) <= not b or a;
    layer2_outputs(5021) <= b and not a;
    layer2_outputs(5022) <= not a or b;
    layer2_outputs(5023) <= b;
    layer2_outputs(5024) <= a;
    layer2_outputs(5025) <= b;
    layer2_outputs(5026) <= not a;
    layer2_outputs(5027) <= a and not b;
    layer2_outputs(5028) <= b;
    layer2_outputs(5029) <= a;
    layer2_outputs(5030) <= a or b;
    layer2_outputs(5031) <= b;
    layer2_outputs(5032) <= b;
    layer2_outputs(5033) <= a and not b;
    layer2_outputs(5034) <= not b or a;
    layer2_outputs(5035) <= not b;
    layer2_outputs(5036) <= b;
    layer2_outputs(5037) <= a and not b;
    layer2_outputs(5038) <= a and not b;
    layer2_outputs(5039) <= b and not a;
    layer2_outputs(5040) <= not b;
    layer2_outputs(5041) <= not b;
    layer2_outputs(5042) <= b;
    layer2_outputs(5043) <= b;
    layer2_outputs(5044) <= not b or a;
    layer2_outputs(5045) <= a xor b;
    layer2_outputs(5046) <= not (a and b);
    layer2_outputs(5047) <= not a;
    layer2_outputs(5048) <= not a;
    layer2_outputs(5049) <= a xor b;
    layer2_outputs(5050) <= not a or b;
    layer2_outputs(5051) <= a xor b;
    layer2_outputs(5052) <= b;
    layer2_outputs(5053) <= b;
    layer2_outputs(5054) <= a xor b;
    layer2_outputs(5055) <= a xor b;
    layer2_outputs(5056) <= not (a xor b);
    layer2_outputs(5057) <= b;
    layer2_outputs(5058) <= a;
    layer2_outputs(5059) <= not b;
    layer2_outputs(5060) <= not b;
    layer2_outputs(5061) <= not a;
    layer2_outputs(5062) <= b and not a;
    layer2_outputs(5063) <= a;
    layer2_outputs(5064) <= a or b;
    layer2_outputs(5065) <= b and not a;
    layer2_outputs(5066) <= a xor b;
    layer2_outputs(5067) <= a and b;
    layer2_outputs(5068) <= not a or b;
    layer2_outputs(5069) <= not (a xor b);
    layer2_outputs(5070) <= not (a xor b);
    layer2_outputs(5071) <= not (a and b);
    layer2_outputs(5072) <= not b;
    layer2_outputs(5073) <= b;
    layer2_outputs(5074) <= b;
    layer2_outputs(5075) <= b and not a;
    layer2_outputs(5076) <= b and not a;
    layer2_outputs(5077) <= not (a and b);
    layer2_outputs(5078) <= 1'b0;
    layer2_outputs(5079) <= a;
    layer2_outputs(5080) <= not b;
    layer2_outputs(5081) <= not a or b;
    layer2_outputs(5082) <= a xor b;
    layer2_outputs(5083) <= not b;
    layer2_outputs(5084) <= a;
    layer2_outputs(5085) <= a xor b;
    layer2_outputs(5086) <= a or b;
    layer2_outputs(5087) <= not (a xor b);
    layer2_outputs(5088) <= not b;
    layer2_outputs(5089) <= not (a xor b);
    layer2_outputs(5090) <= not a;
    layer2_outputs(5091) <= b and not a;
    layer2_outputs(5092) <= a xor b;
    layer2_outputs(5093) <= a and not b;
    layer2_outputs(5094) <= not (a and b);
    layer2_outputs(5095) <= a;
    layer2_outputs(5096) <= a and not b;
    layer2_outputs(5097) <= not (a and b);
    layer2_outputs(5098) <= a or b;
    layer2_outputs(5099) <= not b;
    layer2_outputs(5100) <= b and not a;
    layer2_outputs(5101) <= a and b;
    layer2_outputs(5102) <= b;
    layer2_outputs(5103) <= not (a xor b);
    layer2_outputs(5104) <= a xor b;
    layer2_outputs(5105) <= b;
    layer2_outputs(5106) <= not a;
    layer2_outputs(5107) <= b;
    layer2_outputs(5108) <= a or b;
    layer2_outputs(5109) <= not a;
    layer2_outputs(5110) <= not (a and b);
    layer2_outputs(5111) <= not a or b;
    layer2_outputs(5112) <= not a or b;
    layer2_outputs(5113) <= not (a or b);
    layer2_outputs(5114) <= a and b;
    layer2_outputs(5115) <= not a;
    layer2_outputs(5116) <= not b or a;
    layer2_outputs(5117) <= a and b;
    layer2_outputs(5118) <= not b;
    layer2_outputs(5119) <= not a;
    layer2_outputs(5120) <= a and b;
    layer2_outputs(5121) <= not b;
    layer2_outputs(5122) <= not (a xor b);
    layer2_outputs(5123) <= not (a xor b);
    layer2_outputs(5124) <= not b;
    layer2_outputs(5125) <= b;
    layer2_outputs(5126) <= b and not a;
    layer2_outputs(5127) <= not b;
    layer2_outputs(5128) <= not (a xor b);
    layer2_outputs(5129) <= not a or b;
    layer2_outputs(5130) <= not (a xor b);
    layer2_outputs(5131) <= a or b;
    layer2_outputs(5132) <= not b;
    layer2_outputs(5133) <= not a or b;
    layer2_outputs(5134) <= not (a xor b);
    layer2_outputs(5135) <= not b or a;
    layer2_outputs(5136) <= a;
    layer2_outputs(5137) <= not (a or b);
    layer2_outputs(5138) <= not a;
    layer2_outputs(5139) <= not (a and b);
    layer2_outputs(5140) <= not (a xor b);
    layer2_outputs(5141) <= b and not a;
    layer2_outputs(5142) <= a and not b;
    layer2_outputs(5143) <= not a;
    layer2_outputs(5144) <= not b;
    layer2_outputs(5145) <= not (a and b);
    layer2_outputs(5146) <= a;
    layer2_outputs(5147) <= not (a or b);
    layer2_outputs(5148) <= not (a or b);
    layer2_outputs(5149) <= not (a xor b);
    layer2_outputs(5150) <= not b or a;
    layer2_outputs(5151) <= b;
    layer2_outputs(5152) <= not a or b;
    layer2_outputs(5153) <= b;
    layer2_outputs(5154) <= b and not a;
    layer2_outputs(5155) <= a xor b;
    layer2_outputs(5156) <= not (a or b);
    layer2_outputs(5157) <= b and not a;
    layer2_outputs(5158) <= a;
    layer2_outputs(5159) <= a xor b;
    layer2_outputs(5160) <= not a or b;
    layer2_outputs(5161) <= b;
    layer2_outputs(5162) <= a xor b;
    layer2_outputs(5163) <= not (a and b);
    layer2_outputs(5164) <= a or b;
    layer2_outputs(5165) <= not a;
    layer2_outputs(5166) <= not a or b;
    layer2_outputs(5167) <= b;
    layer2_outputs(5168) <= not b;
    layer2_outputs(5169) <= a or b;
    layer2_outputs(5170) <= b;
    layer2_outputs(5171) <= not (a xor b);
    layer2_outputs(5172) <= not b;
    layer2_outputs(5173) <= a xor b;
    layer2_outputs(5174) <= not b;
    layer2_outputs(5175) <= not (a xor b);
    layer2_outputs(5176) <= not (a xor b);
    layer2_outputs(5177) <= not (a xor b);
    layer2_outputs(5178) <= b;
    layer2_outputs(5179) <= a and not b;
    layer2_outputs(5180) <= a and not b;
    layer2_outputs(5181) <= b;
    layer2_outputs(5182) <= not (a xor b);
    layer2_outputs(5183) <= a or b;
    layer2_outputs(5184) <= not a;
    layer2_outputs(5185) <= not a;
    layer2_outputs(5186) <= b;
    layer2_outputs(5187) <= a;
    layer2_outputs(5188) <= a xor b;
    layer2_outputs(5189) <= not b;
    layer2_outputs(5190) <= not (a xor b);
    layer2_outputs(5191) <= not a;
    layer2_outputs(5192) <= a;
    layer2_outputs(5193) <= not a or b;
    layer2_outputs(5194) <= a and not b;
    layer2_outputs(5195) <= a or b;
    layer2_outputs(5196) <= a or b;
    layer2_outputs(5197) <= not a;
    layer2_outputs(5198) <= a xor b;
    layer2_outputs(5199) <= a;
    layer2_outputs(5200) <= not b;
    layer2_outputs(5201) <= not (a and b);
    layer2_outputs(5202) <= not (a or b);
    layer2_outputs(5203) <= not a or b;
    layer2_outputs(5204) <= not a;
    layer2_outputs(5205) <= not (a or b);
    layer2_outputs(5206) <= not a;
    layer2_outputs(5207) <= not (a xor b);
    layer2_outputs(5208) <= not b or a;
    layer2_outputs(5209) <= a;
    layer2_outputs(5210) <= a;
    layer2_outputs(5211) <= a xor b;
    layer2_outputs(5212) <= a and not b;
    layer2_outputs(5213) <= not (a xor b);
    layer2_outputs(5214) <= not (a xor b);
    layer2_outputs(5215) <= b and not a;
    layer2_outputs(5216) <= not a or b;
    layer2_outputs(5217) <= not (a and b);
    layer2_outputs(5218) <= not b;
    layer2_outputs(5219) <= not a;
    layer2_outputs(5220) <= not b or a;
    layer2_outputs(5221) <= a xor b;
    layer2_outputs(5222) <= a and not b;
    layer2_outputs(5223) <= a;
    layer2_outputs(5224) <= a or b;
    layer2_outputs(5225) <= not a;
    layer2_outputs(5226) <= a xor b;
    layer2_outputs(5227) <= not (a xor b);
    layer2_outputs(5228) <= not (a xor b);
    layer2_outputs(5229) <= a or b;
    layer2_outputs(5230) <= a and b;
    layer2_outputs(5231) <= a and b;
    layer2_outputs(5232) <= a and not b;
    layer2_outputs(5233) <= a and not b;
    layer2_outputs(5234) <= not (a xor b);
    layer2_outputs(5235) <= a or b;
    layer2_outputs(5236) <= not a or b;
    layer2_outputs(5237) <= not a;
    layer2_outputs(5238) <= not a;
    layer2_outputs(5239) <= not (a and b);
    layer2_outputs(5240) <= not (a or b);
    layer2_outputs(5241) <= not a;
    layer2_outputs(5242) <= a xor b;
    layer2_outputs(5243) <= b;
    layer2_outputs(5244) <= a xor b;
    layer2_outputs(5245) <= a;
    layer2_outputs(5246) <= a;
    layer2_outputs(5247) <= not (a xor b);
    layer2_outputs(5248) <= b;
    layer2_outputs(5249) <= not (a xor b);
    layer2_outputs(5250) <= a xor b;
    layer2_outputs(5251) <= a xor b;
    layer2_outputs(5252) <= not a;
    layer2_outputs(5253) <= not a;
    layer2_outputs(5254) <= a or b;
    layer2_outputs(5255) <= not b;
    layer2_outputs(5256) <= not b;
    layer2_outputs(5257) <= a or b;
    layer2_outputs(5258) <= b;
    layer2_outputs(5259) <= not a or b;
    layer2_outputs(5260) <= a xor b;
    layer2_outputs(5261) <= a xor b;
    layer2_outputs(5262) <= not b or a;
    layer2_outputs(5263) <= a and not b;
    layer2_outputs(5264) <= not b or a;
    layer2_outputs(5265) <= not a;
    layer2_outputs(5266) <= b and not a;
    layer2_outputs(5267) <= not (a and b);
    layer2_outputs(5268) <= b;
    layer2_outputs(5269) <= b and not a;
    layer2_outputs(5270) <= a and b;
    layer2_outputs(5271) <= a;
    layer2_outputs(5272) <= not b or a;
    layer2_outputs(5273) <= a and b;
    layer2_outputs(5274) <= b;
    layer2_outputs(5275) <= a;
    layer2_outputs(5276) <= a and b;
    layer2_outputs(5277) <= b;
    layer2_outputs(5278) <= b and not a;
    layer2_outputs(5279) <= a xor b;
    layer2_outputs(5280) <= not a;
    layer2_outputs(5281) <= a;
    layer2_outputs(5282) <= not a;
    layer2_outputs(5283) <= not (a or b);
    layer2_outputs(5284) <= not a;
    layer2_outputs(5285) <= not b;
    layer2_outputs(5286) <= a xor b;
    layer2_outputs(5287) <= not b or a;
    layer2_outputs(5288) <= not (a or b);
    layer2_outputs(5289) <= b;
    layer2_outputs(5290) <= not (a xor b);
    layer2_outputs(5291) <= not a;
    layer2_outputs(5292) <= a and b;
    layer2_outputs(5293) <= b;
    layer2_outputs(5294) <= a;
    layer2_outputs(5295) <= a xor b;
    layer2_outputs(5296) <= b;
    layer2_outputs(5297) <= b;
    layer2_outputs(5298) <= a xor b;
    layer2_outputs(5299) <= a and b;
    layer2_outputs(5300) <= not (a and b);
    layer2_outputs(5301) <= b;
    layer2_outputs(5302) <= not b;
    layer2_outputs(5303) <= a;
    layer2_outputs(5304) <= a;
    layer2_outputs(5305) <= not b;
    layer2_outputs(5306) <= a and not b;
    layer2_outputs(5307) <= not (a xor b);
    layer2_outputs(5308) <= a and not b;
    layer2_outputs(5309) <= not b;
    layer2_outputs(5310) <= not a;
    layer2_outputs(5311) <= a and b;
    layer2_outputs(5312) <= a;
    layer2_outputs(5313) <= not (a and b);
    layer2_outputs(5314) <= a and not b;
    layer2_outputs(5315) <= not b or a;
    layer2_outputs(5316) <= a;
    layer2_outputs(5317) <= not b;
    layer2_outputs(5318) <= a xor b;
    layer2_outputs(5319) <= a xor b;
    layer2_outputs(5320) <= b;
    layer2_outputs(5321) <= not b;
    layer2_outputs(5322) <= not a;
    layer2_outputs(5323) <= a xor b;
    layer2_outputs(5324) <= not a or b;
    layer2_outputs(5325) <= not a or b;
    layer2_outputs(5326) <= a;
    layer2_outputs(5327) <= b;
    layer2_outputs(5328) <= b and not a;
    layer2_outputs(5329) <= not (a and b);
    layer2_outputs(5330) <= b;
    layer2_outputs(5331) <= a or b;
    layer2_outputs(5332) <= a;
    layer2_outputs(5333) <= a;
    layer2_outputs(5334) <= b;
    layer2_outputs(5335) <= a xor b;
    layer2_outputs(5336) <= not a;
    layer2_outputs(5337) <= not b;
    layer2_outputs(5338) <= not a;
    layer2_outputs(5339) <= a;
    layer2_outputs(5340) <= not b or a;
    layer2_outputs(5341) <= a xor b;
    layer2_outputs(5342) <= a and b;
    layer2_outputs(5343) <= not b or a;
    layer2_outputs(5344) <= not b or a;
    layer2_outputs(5345) <= a and not b;
    layer2_outputs(5346) <= a and b;
    layer2_outputs(5347) <= a;
    layer2_outputs(5348) <= a or b;
    layer2_outputs(5349) <= a;
    layer2_outputs(5350) <= not b;
    layer2_outputs(5351) <= b;
    layer2_outputs(5352) <= a xor b;
    layer2_outputs(5353) <= b and not a;
    layer2_outputs(5354) <= b;
    layer2_outputs(5355) <= not b;
    layer2_outputs(5356) <= a or b;
    layer2_outputs(5357) <= not (a xor b);
    layer2_outputs(5358) <= a xor b;
    layer2_outputs(5359) <= not b;
    layer2_outputs(5360) <= a;
    layer2_outputs(5361) <= a or b;
    layer2_outputs(5362) <= not a;
    layer2_outputs(5363) <= a xor b;
    layer2_outputs(5364) <= a xor b;
    layer2_outputs(5365) <= not (a xor b);
    layer2_outputs(5366) <= a and not b;
    layer2_outputs(5367) <= not a or b;
    layer2_outputs(5368) <= a and b;
    layer2_outputs(5369) <= a;
    layer2_outputs(5370) <= not b;
    layer2_outputs(5371) <= not b;
    layer2_outputs(5372) <= not (a and b);
    layer2_outputs(5373) <= a xor b;
    layer2_outputs(5374) <= not (a and b);
    layer2_outputs(5375) <= b;
    layer2_outputs(5376) <= b and not a;
    layer2_outputs(5377) <= b;
    layer2_outputs(5378) <= not a;
    layer2_outputs(5379) <= not (a and b);
    layer2_outputs(5380) <= b;
    layer2_outputs(5381) <= a xor b;
    layer2_outputs(5382) <= not (a xor b);
    layer2_outputs(5383) <= not (a xor b);
    layer2_outputs(5384) <= not b;
    layer2_outputs(5385) <= not (a or b);
    layer2_outputs(5386) <= a or b;
    layer2_outputs(5387) <= a;
    layer2_outputs(5388) <= not (a and b);
    layer2_outputs(5389) <= not b;
    layer2_outputs(5390) <= not a;
    layer2_outputs(5391) <= b;
    layer2_outputs(5392) <= not a or b;
    layer2_outputs(5393) <= a;
    layer2_outputs(5394) <= b;
    layer2_outputs(5395) <= a;
    layer2_outputs(5396) <= a;
    layer2_outputs(5397) <= not (a xor b);
    layer2_outputs(5398) <= a and not b;
    layer2_outputs(5399) <= not (a xor b);
    layer2_outputs(5400) <= a;
    layer2_outputs(5401) <= not (a or b);
    layer2_outputs(5402) <= a;
    layer2_outputs(5403) <= b;
    layer2_outputs(5404) <= not b or a;
    layer2_outputs(5405) <= not b;
    layer2_outputs(5406) <= a and b;
    layer2_outputs(5407) <= not b;
    layer2_outputs(5408) <= not b or a;
    layer2_outputs(5409) <= not b;
    layer2_outputs(5410) <= b and not a;
    layer2_outputs(5411) <= not b or a;
    layer2_outputs(5412) <= not (a xor b);
    layer2_outputs(5413) <= not b or a;
    layer2_outputs(5414) <= not a;
    layer2_outputs(5415) <= a and not b;
    layer2_outputs(5416) <= 1'b0;
    layer2_outputs(5417) <= a;
    layer2_outputs(5418) <= a;
    layer2_outputs(5419) <= a and b;
    layer2_outputs(5420) <= not (a xor b);
    layer2_outputs(5421) <= a xor b;
    layer2_outputs(5422) <= a and b;
    layer2_outputs(5423) <= a xor b;
    layer2_outputs(5424) <= a and not b;
    layer2_outputs(5425) <= not (a xor b);
    layer2_outputs(5426) <= a or b;
    layer2_outputs(5427) <= a or b;
    layer2_outputs(5428) <= a xor b;
    layer2_outputs(5429) <= not (a xor b);
    layer2_outputs(5430) <= b;
    layer2_outputs(5431) <= a and b;
    layer2_outputs(5432) <= a or b;
    layer2_outputs(5433) <= not (a xor b);
    layer2_outputs(5434) <= a xor b;
    layer2_outputs(5435) <= not (a xor b);
    layer2_outputs(5436) <= a xor b;
    layer2_outputs(5437) <= not b;
    layer2_outputs(5438) <= a xor b;
    layer2_outputs(5439) <= a xor b;
    layer2_outputs(5440) <= not (a and b);
    layer2_outputs(5441) <= a;
    layer2_outputs(5442) <= a xor b;
    layer2_outputs(5443) <= b;
    layer2_outputs(5444) <= a or b;
    layer2_outputs(5445) <= not a;
    layer2_outputs(5446) <= a xor b;
    layer2_outputs(5447) <= not b or a;
    layer2_outputs(5448) <= a;
    layer2_outputs(5449) <= a and not b;
    layer2_outputs(5450) <= not b;
    layer2_outputs(5451) <= not b or a;
    layer2_outputs(5452) <= b;
    layer2_outputs(5453) <= not (a xor b);
    layer2_outputs(5454) <= not a;
    layer2_outputs(5455) <= b;
    layer2_outputs(5456) <= not (a or b);
    layer2_outputs(5457) <= not a;
    layer2_outputs(5458) <= b and not a;
    layer2_outputs(5459) <= b;
    layer2_outputs(5460) <= not (a xor b);
    layer2_outputs(5461) <= not b or a;
    layer2_outputs(5462) <= not a;
    layer2_outputs(5463) <= not a or b;
    layer2_outputs(5464) <= not a;
    layer2_outputs(5465) <= not b or a;
    layer2_outputs(5466) <= not b;
    layer2_outputs(5467) <= not b or a;
    layer2_outputs(5468) <= not (a xor b);
    layer2_outputs(5469) <= not b or a;
    layer2_outputs(5470) <= not (a and b);
    layer2_outputs(5471) <= a;
    layer2_outputs(5472) <= 1'b1;
    layer2_outputs(5473) <= b;
    layer2_outputs(5474) <= a and not b;
    layer2_outputs(5475) <= not b;
    layer2_outputs(5476) <= b;
    layer2_outputs(5477) <= a xor b;
    layer2_outputs(5478) <= a;
    layer2_outputs(5479) <= a and b;
    layer2_outputs(5480) <= b and not a;
    layer2_outputs(5481) <= not a;
    layer2_outputs(5482) <= b;
    layer2_outputs(5483) <= a;
    layer2_outputs(5484) <= a and b;
    layer2_outputs(5485) <= not (a and b);
    layer2_outputs(5486) <= b and not a;
    layer2_outputs(5487) <= 1'b0;
    layer2_outputs(5488) <= not (a xor b);
    layer2_outputs(5489) <= not (a xor b);
    layer2_outputs(5490) <= a;
    layer2_outputs(5491) <= not (a and b);
    layer2_outputs(5492) <= a;
    layer2_outputs(5493) <= a xor b;
    layer2_outputs(5494) <= a;
    layer2_outputs(5495) <= not b;
    layer2_outputs(5496) <= not (a and b);
    layer2_outputs(5497) <= a xor b;
    layer2_outputs(5498) <= a and not b;
    layer2_outputs(5499) <= not (a xor b);
    layer2_outputs(5500) <= not (a and b);
    layer2_outputs(5501) <= not b or a;
    layer2_outputs(5502) <= a or b;
    layer2_outputs(5503) <= a;
    layer2_outputs(5504) <= a xor b;
    layer2_outputs(5505) <= a;
    layer2_outputs(5506) <= b;
    layer2_outputs(5507) <= not b;
    layer2_outputs(5508) <= not a;
    layer2_outputs(5509) <= not b;
    layer2_outputs(5510) <= 1'b0;
    layer2_outputs(5511) <= a xor b;
    layer2_outputs(5512) <= a and b;
    layer2_outputs(5513) <= b and not a;
    layer2_outputs(5514) <= b;
    layer2_outputs(5515) <= a and not b;
    layer2_outputs(5516) <= a;
    layer2_outputs(5517) <= b;
    layer2_outputs(5518) <= a and b;
    layer2_outputs(5519) <= a;
    layer2_outputs(5520) <= not (a and b);
    layer2_outputs(5521) <= 1'b1;
    layer2_outputs(5522) <= a;
    layer2_outputs(5523) <= a and b;
    layer2_outputs(5524) <= b;
    layer2_outputs(5525) <= not b;
    layer2_outputs(5526) <= a and b;
    layer2_outputs(5527) <= a and b;
    layer2_outputs(5528) <= a xor b;
    layer2_outputs(5529) <= b;
    layer2_outputs(5530) <= not (a and b);
    layer2_outputs(5531) <= not (a xor b);
    layer2_outputs(5532) <= b;
    layer2_outputs(5533) <= a;
    layer2_outputs(5534) <= b;
    layer2_outputs(5535) <= a xor b;
    layer2_outputs(5536) <= not a;
    layer2_outputs(5537) <= not a;
    layer2_outputs(5538) <= a xor b;
    layer2_outputs(5539) <= not (a xor b);
    layer2_outputs(5540) <= a;
    layer2_outputs(5541) <= a;
    layer2_outputs(5542) <= not (a or b);
    layer2_outputs(5543) <= a or b;
    layer2_outputs(5544) <= b;
    layer2_outputs(5545) <= not a;
    layer2_outputs(5546) <= not b or a;
    layer2_outputs(5547) <= not a;
    layer2_outputs(5548) <= a or b;
    layer2_outputs(5549) <= not (a xor b);
    layer2_outputs(5550) <= a xor b;
    layer2_outputs(5551) <= not b or a;
    layer2_outputs(5552) <= b and not a;
    layer2_outputs(5553) <= not b;
    layer2_outputs(5554) <= not b or a;
    layer2_outputs(5555) <= not (a xor b);
    layer2_outputs(5556) <= a and not b;
    layer2_outputs(5557) <= not b;
    layer2_outputs(5558) <= a and b;
    layer2_outputs(5559) <= b;
    layer2_outputs(5560) <= a;
    layer2_outputs(5561) <= not (a or b);
    layer2_outputs(5562) <= not (a or b);
    layer2_outputs(5563) <= a;
    layer2_outputs(5564) <= not (a and b);
    layer2_outputs(5565) <= a;
    layer2_outputs(5566) <= a and b;
    layer2_outputs(5567) <= b;
    layer2_outputs(5568) <= not (a and b);
    layer2_outputs(5569) <= not a or b;
    layer2_outputs(5570) <= a xor b;
    layer2_outputs(5571) <= a xor b;
    layer2_outputs(5572) <= not b;
    layer2_outputs(5573) <= not (a or b);
    layer2_outputs(5574) <= a xor b;
    layer2_outputs(5575) <= not a or b;
    layer2_outputs(5576) <= not a;
    layer2_outputs(5577) <= a xor b;
    layer2_outputs(5578) <= a;
    layer2_outputs(5579) <= a and not b;
    layer2_outputs(5580) <= b and not a;
    layer2_outputs(5581) <= a xor b;
    layer2_outputs(5582) <= not b;
    layer2_outputs(5583) <= a;
    layer2_outputs(5584) <= b and not a;
    layer2_outputs(5585) <= a xor b;
    layer2_outputs(5586) <= a and not b;
    layer2_outputs(5587) <= not (a and b);
    layer2_outputs(5588) <= not b or a;
    layer2_outputs(5589) <= a;
    layer2_outputs(5590) <= not b or a;
    layer2_outputs(5591) <= a and not b;
    layer2_outputs(5592) <= not a;
    layer2_outputs(5593) <= a or b;
    layer2_outputs(5594) <= not (a or b);
    layer2_outputs(5595) <= a or b;
    layer2_outputs(5596) <= a xor b;
    layer2_outputs(5597) <= not (a and b);
    layer2_outputs(5598) <= a xor b;
    layer2_outputs(5599) <= not a or b;
    layer2_outputs(5600) <= not a or b;
    layer2_outputs(5601) <= not a or b;
    layer2_outputs(5602) <= b and not a;
    layer2_outputs(5603) <= b;
    layer2_outputs(5604) <= not (a xor b);
    layer2_outputs(5605) <= b;
    layer2_outputs(5606) <= b;
    layer2_outputs(5607) <= not b;
    layer2_outputs(5608) <= b;
    layer2_outputs(5609) <= not b;
    layer2_outputs(5610) <= not b;
    layer2_outputs(5611) <= not b;
    layer2_outputs(5612) <= b;
    layer2_outputs(5613) <= b and not a;
    layer2_outputs(5614) <= a and not b;
    layer2_outputs(5615) <= not b;
    layer2_outputs(5616) <= b;
    layer2_outputs(5617) <= not a;
    layer2_outputs(5618) <= not a;
    layer2_outputs(5619) <= not (a and b);
    layer2_outputs(5620) <= not b;
    layer2_outputs(5621) <= a;
    layer2_outputs(5622) <= not a;
    layer2_outputs(5623) <= not a or b;
    layer2_outputs(5624) <= b and not a;
    layer2_outputs(5625) <= a xor b;
    layer2_outputs(5626) <= a;
    layer2_outputs(5627) <= not b;
    layer2_outputs(5628) <= not a;
    layer2_outputs(5629) <= not (a and b);
    layer2_outputs(5630) <= not b;
    layer2_outputs(5631) <= a xor b;
    layer2_outputs(5632) <= not b;
    layer2_outputs(5633) <= not b;
    layer2_outputs(5634) <= b and not a;
    layer2_outputs(5635) <= not a;
    layer2_outputs(5636) <= not (a or b);
    layer2_outputs(5637) <= not b or a;
    layer2_outputs(5638) <= a and not b;
    layer2_outputs(5639) <= a and not b;
    layer2_outputs(5640) <= a;
    layer2_outputs(5641) <= not b or a;
    layer2_outputs(5642) <= a;
    layer2_outputs(5643) <= not a;
    layer2_outputs(5644) <= a xor b;
    layer2_outputs(5645) <= b;
    layer2_outputs(5646) <= a;
    layer2_outputs(5647) <= b;
    layer2_outputs(5648) <= not (a xor b);
    layer2_outputs(5649) <= not a;
    layer2_outputs(5650) <= not a or b;
    layer2_outputs(5651) <= b;
    layer2_outputs(5652) <= b;
    layer2_outputs(5653) <= b;
    layer2_outputs(5654) <= a xor b;
    layer2_outputs(5655) <= not b or a;
    layer2_outputs(5656) <= a;
    layer2_outputs(5657) <= a and not b;
    layer2_outputs(5658) <= b;
    layer2_outputs(5659) <= not b or a;
    layer2_outputs(5660) <= not b or a;
    layer2_outputs(5661) <= not a;
    layer2_outputs(5662) <= a;
    layer2_outputs(5663) <= not (a and b);
    layer2_outputs(5664) <= not (a and b);
    layer2_outputs(5665) <= not b or a;
    layer2_outputs(5666) <= b;
    layer2_outputs(5667) <= not (a xor b);
    layer2_outputs(5668) <= 1'b0;
    layer2_outputs(5669) <= a xor b;
    layer2_outputs(5670) <= not b;
    layer2_outputs(5671) <= a;
    layer2_outputs(5672) <= 1'b0;
    layer2_outputs(5673) <= a;
    layer2_outputs(5674) <= b and not a;
    layer2_outputs(5675) <= a;
    layer2_outputs(5676) <= 1'b0;
    layer2_outputs(5677) <= b;
    layer2_outputs(5678) <= not (a xor b);
    layer2_outputs(5679) <= a and b;
    layer2_outputs(5680) <= not (a xor b);
    layer2_outputs(5681) <= b;
    layer2_outputs(5682) <= not b;
    layer2_outputs(5683) <= not b or a;
    layer2_outputs(5684) <= a xor b;
    layer2_outputs(5685) <= a;
    layer2_outputs(5686) <= a;
    layer2_outputs(5687) <= a;
    layer2_outputs(5688) <= not (a xor b);
    layer2_outputs(5689) <= a and b;
    layer2_outputs(5690) <= not (a or b);
    layer2_outputs(5691) <= a;
    layer2_outputs(5692) <= a xor b;
    layer2_outputs(5693) <= a and b;
    layer2_outputs(5694) <= not a;
    layer2_outputs(5695) <= not (a xor b);
    layer2_outputs(5696) <= not a;
    layer2_outputs(5697) <= not b;
    layer2_outputs(5698) <= not b or a;
    layer2_outputs(5699) <= not b or a;
    layer2_outputs(5700) <= b and not a;
    layer2_outputs(5701) <= a and not b;
    layer2_outputs(5702) <= not b;
    layer2_outputs(5703) <= a xor b;
    layer2_outputs(5704) <= b;
    layer2_outputs(5705) <= not (a or b);
    layer2_outputs(5706) <= a and not b;
    layer2_outputs(5707) <= not b;
    layer2_outputs(5708) <= a;
    layer2_outputs(5709) <= a or b;
    layer2_outputs(5710) <= b;
    layer2_outputs(5711) <= not b or a;
    layer2_outputs(5712) <= b;
    layer2_outputs(5713) <= not b or a;
    layer2_outputs(5714) <= b and not a;
    layer2_outputs(5715) <= b;
    layer2_outputs(5716) <= a and not b;
    layer2_outputs(5717) <= a or b;
    layer2_outputs(5718) <= not (a xor b);
    layer2_outputs(5719) <= not (a xor b);
    layer2_outputs(5720) <= a and b;
    layer2_outputs(5721) <= a and not b;
    layer2_outputs(5722) <= a xor b;
    layer2_outputs(5723) <= b and not a;
    layer2_outputs(5724) <= not b or a;
    layer2_outputs(5725) <= not b;
    layer2_outputs(5726) <= not b;
    layer2_outputs(5727) <= not (a or b);
    layer2_outputs(5728) <= not b;
    layer2_outputs(5729) <= a xor b;
    layer2_outputs(5730) <= b;
    layer2_outputs(5731) <= a xor b;
    layer2_outputs(5732) <= a or b;
    layer2_outputs(5733) <= b and not a;
    layer2_outputs(5734) <= not a;
    layer2_outputs(5735) <= not a;
    layer2_outputs(5736) <= a;
    layer2_outputs(5737) <= a xor b;
    layer2_outputs(5738) <= a xor b;
    layer2_outputs(5739) <= a;
    layer2_outputs(5740) <= not a;
    layer2_outputs(5741) <= a xor b;
    layer2_outputs(5742) <= not (a xor b);
    layer2_outputs(5743) <= not a;
    layer2_outputs(5744) <= not b;
    layer2_outputs(5745) <= not (a or b);
    layer2_outputs(5746) <= not b;
    layer2_outputs(5747) <= not (a xor b);
    layer2_outputs(5748) <= a or b;
    layer2_outputs(5749) <= not b;
    layer2_outputs(5750) <= a and b;
    layer2_outputs(5751) <= a and b;
    layer2_outputs(5752) <= b;
    layer2_outputs(5753) <= a and b;
    layer2_outputs(5754) <= b;
    layer2_outputs(5755) <= not (a xor b);
    layer2_outputs(5756) <= not a;
    layer2_outputs(5757) <= a;
    layer2_outputs(5758) <= b;
    layer2_outputs(5759) <= a and not b;
    layer2_outputs(5760) <= not (a or b);
    layer2_outputs(5761) <= not a or b;
    layer2_outputs(5762) <= not a;
    layer2_outputs(5763) <= not b;
    layer2_outputs(5764) <= a;
    layer2_outputs(5765) <= not b;
    layer2_outputs(5766) <= a or b;
    layer2_outputs(5767) <= a;
    layer2_outputs(5768) <= a;
    layer2_outputs(5769) <= not b or a;
    layer2_outputs(5770) <= a or b;
    layer2_outputs(5771) <= a xor b;
    layer2_outputs(5772) <= a xor b;
    layer2_outputs(5773) <= not a or b;
    layer2_outputs(5774) <= not (a xor b);
    layer2_outputs(5775) <= not b or a;
    layer2_outputs(5776) <= a and not b;
    layer2_outputs(5777) <= not (a and b);
    layer2_outputs(5778) <= b;
    layer2_outputs(5779) <= a xor b;
    layer2_outputs(5780) <= not b;
    layer2_outputs(5781) <= not b or a;
    layer2_outputs(5782) <= not (a xor b);
    layer2_outputs(5783) <= b;
    layer2_outputs(5784) <= not b or a;
    layer2_outputs(5785) <= not (a xor b);
    layer2_outputs(5786) <= 1'b1;
    layer2_outputs(5787) <= not (a xor b);
    layer2_outputs(5788) <= a xor b;
    layer2_outputs(5789) <= not b;
    layer2_outputs(5790) <= not b;
    layer2_outputs(5791) <= a and b;
    layer2_outputs(5792) <= not b;
    layer2_outputs(5793) <= a or b;
    layer2_outputs(5794) <= not b or a;
    layer2_outputs(5795) <= not (a or b);
    layer2_outputs(5796) <= not b or a;
    layer2_outputs(5797) <= b;
    layer2_outputs(5798) <= not (a and b);
    layer2_outputs(5799) <= a;
    layer2_outputs(5800) <= not (a and b);
    layer2_outputs(5801) <= a xor b;
    layer2_outputs(5802) <= b;
    layer2_outputs(5803) <= a xor b;
    layer2_outputs(5804) <= not (a xor b);
    layer2_outputs(5805) <= b;
    layer2_outputs(5806) <= not b;
    layer2_outputs(5807) <= not b;
    layer2_outputs(5808) <= b;
    layer2_outputs(5809) <= not b or a;
    layer2_outputs(5810) <= not (a xor b);
    layer2_outputs(5811) <= b and not a;
    layer2_outputs(5812) <= a;
    layer2_outputs(5813) <= not b;
    layer2_outputs(5814) <= a and not b;
    layer2_outputs(5815) <= a xor b;
    layer2_outputs(5816) <= not a;
    layer2_outputs(5817) <= a and not b;
    layer2_outputs(5818) <= not b or a;
    layer2_outputs(5819) <= 1'b0;
    layer2_outputs(5820) <= not (a and b);
    layer2_outputs(5821) <= a;
    layer2_outputs(5822) <= not (a and b);
    layer2_outputs(5823) <= a and b;
    layer2_outputs(5824) <= b and not a;
    layer2_outputs(5825) <= not (a and b);
    layer2_outputs(5826) <= not a;
    layer2_outputs(5827) <= not (a or b);
    layer2_outputs(5828) <= a and not b;
    layer2_outputs(5829) <= a xor b;
    layer2_outputs(5830) <= b;
    layer2_outputs(5831) <= a;
    layer2_outputs(5832) <= not b;
    layer2_outputs(5833) <= a or b;
    layer2_outputs(5834) <= not b or a;
    layer2_outputs(5835) <= not b;
    layer2_outputs(5836) <= not (a and b);
    layer2_outputs(5837) <= not (a xor b);
    layer2_outputs(5838) <= a;
    layer2_outputs(5839) <= a or b;
    layer2_outputs(5840) <= not b;
    layer2_outputs(5841) <= not b;
    layer2_outputs(5842) <= not (a and b);
    layer2_outputs(5843) <= a or b;
    layer2_outputs(5844) <= not (a or b);
    layer2_outputs(5845) <= a;
    layer2_outputs(5846) <= not (a xor b);
    layer2_outputs(5847) <= not (a xor b);
    layer2_outputs(5848) <= a;
    layer2_outputs(5849) <= a and not b;
    layer2_outputs(5850) <= a;
    layer2_outputs(5851) <= not b;
    layer2_outputs(5852) <= a xor b;
    layer2_outputs(5853) <= not b or a;
    layer2_outputs(5854) <= not a;
    layer2_outputs(5855) <= not a or b;
    layer2_outputs(5856) <= not (a or b);
    layer2_outputs(5857) <= b and not a;
    layer2_outputs(5858) <= a;
    layer2_outputs(5859) <= not b;
    layer2_outputs(5860) <= a and not b;
    layer2_outputs(5861) <= b;
    layer2_outputs(5862) <= a or b;
    layer2_outputs(5863) <= not (a and b);
    layer2_outputs(5864) <= not (a and b);
    layer2_outputs(5865) <= not b;
    layer2_outputs(5866) <= not a;
    layer2_outputs(5867) <= a xor b;
    layer2_outputs(5868) <= not (a xor b);
    layer2_outputs(5869) <= b and not a;
    layer2_outputs(5870) <= b;
    layer2_outputs(5871) <= not a;
    layer2_outputs(5872) <= not a or b;
    layer2_outputs(5873) <= not (a and b);
    layer2_outputs(5874) <= not (a and b);
    layer2_outputs(5875) <= not (a xor b);
    layer2_outputs(5876) <= not (a xor b);
    layer2_outputs(5877) <= a xor b;
    layer2_outputs(5878) <= a or b;
    layer2_outputs(5879) <= not b or a;
    layer2_outputs(5880) <= not a or b;
    layer2_outputs(5881) <= not b;
    layer2_outputs(5882) <= a and b;
    layer2_outputs(5883) <= not (a xor b);
    layer2_outputs(5884) <= a or b;
    layer2_outputs(5885) <= b;
    layer2_outputs(5886) <= a xor b;
    layer2_outputs(5887) <= a;
    layer2_outputs(5888) <= b;
    layer2_outputs(5889) <= not (a xor b);
    layer2_outputs(5890) <= b;
    layer2_outputs(5891) <= not a;
    layer2_outputs(5892) <= a and b;
    layer2_outputs(5893) <= not b;
    layer2_outputs(5894) <= b;
    layer2_outputs(5895) <= a;
    layer2_outputs(5896) <= not a or b;
    layer2_outputs(5897) <= a;
    layer2_outputs(5898) <= 1'b0;
    layer2_outputs(5899) <= not a;
    layer2_outputs(5900) <= b;
    layer2_outputs(5901) <= a and b;
    layer2_outputs(5902) <= not b;
    layer2_outputs(5903) <= not (a xor b);
    layer2_outputs(5904) <= not a or b;
    layer2_outputs(5905) <= not b or a;
    layer2_outputs(5906) <= b;
    layer2_outputs(5907) <= not a;
    layer2_outputs(5908) <= not (a xor b);
    layer2_outputs(5909) <= not a or b;
    layer2_outputs(5910) <= a xor b;
    layer2_outputs(5911) <= not (a or b);
    layer2_outputs(5912) <= a or b;
    layer2_outputs(5913) <= a and b;
    layer2_outputs(5914) <= b;
    layer2_outputs(5915) <= a xor b;
    layer2_outputs(5916) <= not b;
    layer2_outputs(5917) <= not a;
    layer2_outputs(5918) <= not b;
    layer2_outputs(5919) <= not b;
    layer2_outputs(5920) <= not a;
    layer2_outputs(5921) <= a and b;
    layer2_outputs(5922) <= b;
    layer2_outputs(5923) <= not a or b;
    layer2_outputs(5924) <= a;
    layer2_outputs(5925) <= a;
    layer2_outputs(5926) <= a;
    layer2_outputs(5927) <= not (a xor b);
    layer2_outputs(5928) <= a;
    layer2_outputs(5929) <= a xor b;
    layer2_outputs(5930) <= not b or a;
    layer2_outputs(5931) <= a xor b;
    layer2_outputs(5932) <= not a;
    layer2_outputs(5933) <= not (a and b);
    layer2_outputs(5934) <= not a;
    layer2_outputs(5935) <= a;
    layer2_outputs(5936) <= not b or a;
    layer2_outputs(5937) <= not b;
    layer2_outputs(5938) <= a and b;
    layer2_outputs(5939) <= a xor b;
    layer2_outputs(5940) <= not b;
    layer2_outputs(5941) <= a or b;
    layer2_outputs(5942) <= a;
    layer2_outputs(5943) <= not a;
    layer2_outputs(5944) <= a and b;
    layer2_outputs(5945) <= not a;
    layer2_outputs(5946) <= not (a and b);
    layer2_outputs(5947) <= not a;
    layer2_outputs(5948) <= a;
    layer2_outputs(5949) <= not a;
    layer2_outputs(5950) <= not (a and b);
    layer2_outputs(5951) <= not (a xor b);
    layer2_outputs(5952) <= not a;
    layer2_outputs(5953) <= not b or a;
    layer2_outputs(5954) <= not b;
    layer2_outputs(5955) <= not (a and b);
    layer2_outputs(5956) <= not (a xor b);
    layer2_outputs(5957) <= not (a xor b);
    layer2_outputs(5958) <= b;
    layer2_outputs(5959) <= a or b;
    layer2_outputs(5960) <= not a or b;
    layer2_outputs(5961) <= not b;
    layer2_outputs(5962) <= a and b;
    layer2_outputs(5963) <= not (a and b);
    layer2_outputs(5964) <= not a;
    layer2_outputs(5965) <= not a;
    layer2_outputs(5966) <= not (a and b);
    layer2_outputs(5967) <= not a or b;
    layer2_outputs(5968) <= not (a and b);
    layer2_outputs(5969) <= not (a and b);
    layer2_outputs(5970) <= b and not a;
    layer2_outputs(5971) <= a;
    layer2_outputs(5972) <= not (a xor b);
    layer2_outputs(5973) <= not b or a;
    layer2_outputs(5974) <= not a;
    layer2_outputs(5975) <= not (a xor b);
    layer2_outputs(5976) <= not (a xor b);
    layer2_outputs(5977) <= not (a xor b);
    layer2_outputs(5978) <= not a;
    layer2_outputs(5979) <= b;
    layer2_outputs(5980) <= b and not a;
    layer2_outputs(5981) <= not (a and b);
    layer2_outputs(5982) <= not (a and b);
    layer2_outputs(5983) <= b;
    layer2_outputs(5984) <= b;
    layer2_outputs(5985) <= not a;
    layer2_outputs(5986) <= not a or b;
    layer2_outputs(5987) <= a;
    layer2_outputs(5988) <= not b or a;
    layer2_outputs(5989) <= not a;
    layer2_outputs(5990) <= not (a xor b);
    layer2_outputs(5991) <= a or b;
    layer2_outputs(5992) <= b and not a;
    layer2_outputs(5993) <= not b;
    layer2_outputs(5994) <= a;
    layer2_outputs(5995) <= b;
    layer2_outputs(5996) <= a xor b;
    layer2_outputs(5997) <= not a;
    layer2_outputs(5998) <= not (a xor b);
    layer2_outputs(5999) <= b;
    layer2_outputs(6000) <= b;
    layer2_outputs(6001) <= a or b;
    layer2_outputs(6002) <= a and b;
    layer2_outputs(6003) <= b;
    layer2_outputs(6004) <= a;
    layer2_outputs(6005) <= a and b;
    layer2_outputs(6006) <= b and not a;
    layer2_outputs(6007) <= not a;
    layer2_outputs(6008) <= not a or b;
    layer2_outputs(6009) <= not b;
    layer2_outputs(6010) <= not (a xor b);
    layer2_outputs(6011) <= not b or a;
    layer2_outputs(6012) <= a;
    layer2_outputs(6013) <= not (a or b);
    layer2_outputs(6014) <= not a;
    layer2_outputs(6015) <= not (a or b);
    layer2_outputs(6016) <= not b or a;
    layer2_outputs(6017) <= a xor b;
    layer2_outputs(6018) <= not a or b;
    layer2_outputs(6019) <= a xor b;
    layer2_outputs(6020) <= not a;
    layer2_outputs(6021) <= not (a xor b);
    layer2_outputs(6022) <= b and not a;
    layer2_outputs(6023) <= a or b;
    layer2_outputs(6024) <= a and b;
    layer2_outputs(6025) <= not b;
    layer2_outputs(6026) <= not (a xor b);
    layer2_outputs(6027) <= a and not b;
    layer2_outputs(6028) <= a;
    layer2_outputs(6029) <= not (a xor b);
    layer2_outputs(6030) <= not b or a;
    layer2_outputs(6031) <= not a;
    layer2_outputs(6032) <= not b;
    layer2_outputs(6033) <= a and not b;
    layer2_outputs(6034) <= b;
    layer2_outputs(6035) <= a xor b;
    layer2_outputs(6036) <= not (a xor b);
    layer2_outputs(6037) <= not b;
    layer2_outputs(6038) <= a and b;
    layer2_outputs(6039) <= not a;
    layer2_outputs(6040) <= b;
    layer2_outputs(6041) <= not a or b;
    layer2_outputs(6042) <= not a;
    layer2_outputs(6043) <= not (a xor b);
    layer2_outputs(6044) <= not a;
    layer2_outputs(6045) <= b and not a;
    layer2_outputs(6046) <= a;
    layer2_outputs(6047) <= a and b;
    layer2_outputs(6048) <= not (a xor b);
    layer2_outputs(6049) <= a;
    layer2_outputs(6050) <= a and b;
    layer2_outputs(6051) <= a or b;
    layer2_outputs(6052) <= b;
    layer2_outputs(6053) <= a;
    layer2_outputs(6054) <= b;
    layer2_outputs(6055) <= b;
    layer2_outputs(6056) <= not (a or b);
    layer2_outputs(6057) <= not (a xor b);
    layer2_outputs(6058) <= not a;
    layer2_outputs(6059) <= not a;
    layer2_outputs(6060) <= b;
    layer2_outputs(6061) <= a or b;
    layer2_outputs(6062) <= not (a xor b);
    layer2_outputs(6063) <= a or b;
    layer2_outputs(6064) <= a xor b;
    layer2_outputs(6065) <= b;
    layer2_outputs(6066) <= not (a and b);
    layer2_outputs(6067) <= a;
    layer2_outputs(6068) <= not (a or b);
    layer2_outputs(6069) <= a xor b;
    layer2_outputs(6070) <= not (a xor b);
    layer2_outputs(6071) <= a;
    layer2_outputs(6072) <= not (a xor b);
    layer2_outputs(6073) <= a and not b;
    layer2_outputs(6074) <= a and not b;
    layer2_outputs(6075) <= not a;
    layer2_outputs(6076) <= a;
    layer2_outputs(6077) <= not (a xor b);
    layer2_outputs(6078) <= not (a xor b);
    layer2_outputs(6079) <= a;
    layer2_outputs(6080) <= not (a or b);
    layer2_outputs(6081) <= not (a and b);
    layer2_outputs(6082) <= b and not a;
    layer2_outputs(6083) <= a;
    layer2_outputs(6084) <= a xor b;
    layer2_outputs(6085) <= a or b;
    layer2_outputs(6086) <= b;
    layer2_outputs(6087) <= not (a and b);
    layer2_outputs(6088) <= a;
    layer2_outputs(6089) <= 1'b1;
    layer2_outputs(6090) <= not (a xor b);
    layer2_outputs(6091) <= not b or a;
    layer2_outputs(6092) <= b and not a;
    layer2_outputs(6093) <= b;
    layer2_outputs(6094) <= not b;
    layer2_outputs(6095) <= a;
    layer2_outputs(6096) <= a xor b;
    layer2_outputs(6097) <= b;
    layer2_outputs(6098) <= not b;
    layer2_outputs(6099) <= not b or a;
    layer2_outputs(6100) <= not (a and b);
    layer2_outputs(6101) <= a;
    layer2_outputs(6102) <= not a;
    layer2_outputs(6103) <= a and not b;
    layer2_outputs(6104) <= b and not a;
    layer2_outputs(6105) <= a xor b;
    layer2_outputs(6106) <= not b;
    layer2_outputs(6107) <= not a;
    layer2_outputs(6108) <= b;
    layer2_outputs(6109) <= b;
    layer2_outputs(6110) <= not a or b;
    layer2_outputs(6111) <= a and not b;
    layer2_outputs(6112) <= not (a xor b);
    layer2_outputs(6113) <= a xor b;
    layer2_outputs(6114) <= a or b;
    layer2_outputs(6115) <= not a or b;
    layer2_outputs(6116) <= a;
    layer2_outputs(6117) <= not b or a;
    layer2_outputs(6118) <= a;
    layer2_outputs(6119) <= not (a or b);
    layer2_outputs(6120) <= not (a xor b);
    layer2_outputs(6121) <= a and b;
    layer2_outputs(6122) <= not a;
    layer2_outputs(6123) <= a;
    layer2_outputs(6124) <= not (a xor b);
    layer2_outputs(6125) <= not b;
    layer2_outputs(6126) <= 1'b0;
    layer2_outputs(6127) <= not a;
    layer2_outputs(6128) <= a or b;
    layer2_outputs(6129) <= b and not a;
    layer2_outputs(6130) <= a xor b;
    layer2_outputs(6131) <= not a or b;
    layer2_outputs(6132) <= not (a xor b);
    layer2_outputs(6133) <= not (a or b);
    layer2_outputs(6134) <= b;
    layer2_outputs(6135) <= not b or a;
    layer2_outputs(6136) <= a;
    layer2_outputs(6137) <= b and not a;
    layer2_outputs(6138) <= a;
    layer2_outputs(6139) <= a xor b;
    layer2_outputs(6140) <= not (a and b);
    layer2_outputs(6141) <= not b;
    layer2_outputs(6142) <= not a;
    layer2_outputs(6143) <= a;
    layer2_outputs(6144) <= b;
    layer2_outputs(6145) <= a or b;
    layer2_outputs(6146) <= a xor b;
    layer2_outputs(6147) <= b;
    layer2_outputs(6148) <= a xor b;
    layer2_outputs(6149) <= not (a and b);
    layer2_outputs(6150) <= not (a xor b);
    layer2_outputs(6151) <= not (a xor b);
    layer2_outputs(6152) <= a or b;
    layer2_outputs(6153) <= a xor b;
    layer2_outputs(6154) <= not (a and b);
    layer2_outputs(6155) <= a and b;
    layer2_outputs(6156) <= a;
    layer2_outputs(6157) <= a;
    layer2_outputs(6158) <= not b;
    layer2_outputs(6159) <= not b or a;
    layer2_outputs(6160) <= not (a or b);
    layer2_outputs(6161) <= not a;
    layer2_outputs(6162) <= a and not b;
    layer2_outputs(6163) <= a and not b;
    layer2_outputs(6164) <= a;
    layer2_outputs(6165) <= a and b;
    layer2_outputs(6166) <= b;
    layer2_outputs(6167) <= not b or a;
    layer2_outputs(6168) <= not a;
    layer2_outputs(6169) <= a and not b;
    layer2_outputs(6170) <= not (a xor b);
    layer2_outputs(6171) <= a;
    layer2_outputs(6172) <= a;
    layer2_outputs(6173) <= not (a xor b);
    layer2_outputs(6174) <= a;
    layer2_outputs(6175) <= a;
    layer2_outputs(6176) <= not a or b;
    layer2_outputs(6177) <= a xor b;
    layer2_outputs(6178) <= not (a and b);
    layer2_outputs(6179) <= a or b;
    layer2_outputs(6180) <= a xor b;
    layer2_outputs(6181) <= a and b;
    layer2_outputs(6182) <= a;
    layer2_outputs(6183) <= not b;
    layer2_outputs(6184) <= not b;
    layer2_outputs(6185) <= b and not a;
    layer2_outputs(6186) <= a and not b;
    layer2_outputs(6187) <= a xor b;
    layer2_outputs(6188) <= not (a and b);
    layer2_outputs(6189) <= not a;
    layer2_outputs(6190) <= a and not b;
    layer2_outputs(6191) <= not (a xor b);
    layer2_outputs(6192) <= a;
    layer2_outputs(6193) <= not (a or b);
    layer2_outputs(6194) <= not a or b;
    layer2_outputs(6195) <= b;
    layer2_outputs(6196) <= not (a or b);
    layer2_outputs(6197) <= a and b;
    layer2_outputs(6198) <= not b;
    layer2_outputs(6199) <= a or b;
    layer2_outputs(6200) <= a;
    layer2_outputs(6201) <= not a or b;
    layer2_outputs(6202) <= b;
    layer2_outputs(6203) <= b;
    layer2_outputs(6204) <= not (a xor b);
    layer2_outputs(6205) <= not (a xor b);
    layer2_outputs(6206) <= not (a and b);
    layer2_outputs(6207) <= b;
    layer2_outputs(6208) <= not (a xor b);
    layer2_outputs(6209) <= a or b;
    layer2_outputs(6210) <= b;
    layer2_outputs(6211) <= not a;
    layer2_outputs(6212) <= a;
    layer2_outputs(6213) <= not b;
    layer2_outputs(6214) <= not (a xor b);
    layer2_outputs(6215) <= a and b;
    layer2_outputs(6216) <= not b;
    layer2_outputs(6217) <= a xor b;
    layer2_outputs(6218) <= not (a or b);
    layer2_outputs(6219) <= not (a xor b);
    layer2_outputs(6220) <= b;
    layer2_outputs(6221) <= not b;
    layer2_outputs(6222) <= b;
    layer2_outputs(6223) <= not b or a;
    layer2_outputs(6224) <= a or b;
    layer2_outputs(6225) <= not a;
    layer2_outputs(6226) <= not b;
    layer2_outputs(6227) <= not (a and b);
    layer2_outputs(6228) <= a;
    layer2_outputs(6229) <= a and not b;
    layer2_outputs(6230) <= a xor b;
    layer2_outputs(6231) <= a or b;
    layer2_outputs(6232) <= a and not b;
    layer2_outputs(6233) <= a and not b;
    layer2_outputs(6234) <= not b or a;
    layer2_outputs(6235) <= not (a and b);
    layer2_outputs(6236) <= a;
    layer2_outputs(6237) <= b and not a;
    layer2_outputs(6238) <= not a;
    layer2_outputs(6239) <= b;
    layer2_outputs(6240) <= not a or b;
    layer2_outputs(6241) <= not b;
    layer2_outputs(6242) <= a xor b;
    layer2_outputs(6243) <= not b;
    layer2_outputs(6244) <= not a or b;
    layer2_outputs(6245) <= not b;
    layer2_outputs(6246) <= not a;
    layer2_outputs(6247) <= not (a xor b);
    layer2_outputs(6248) <= not a;
    layer2_outputs(6249) <= not b or a;
    layer2_outputs(6250) <= not a or b;
    layer2_outputs(6251) <= not b;
    layer2_outputs(6252) <= not b;
    layer2_outputs(6253) <= a or b;
    layer2_outputs(6254) <= not (a xor b);
    layer2_outputs(6255) <= not a or b;
    layer2_outputs(6256) <= not (a or b);
    layer2_outputs(6257) <= not (a xor b);
    layer2_outputs(6258) <= not b;
    layer2_outputs(6259) <= not b;
    layer2_outputs(6260) <= not (a xor b);
    layer2_outputs(6261) <= a and b;
    layer2_outputs(6262) <= not b;
    layer2_outputs(6263) <= not a or b;
    layer2_outputs(6264) <= b;
    layer2_outputs(6265) <= a or b;
    layer2_outputs(6266) <= a xor b;
    layer2_outputs(6267) <= not b;
    layer2_outputs(6268) <= not (a xor b);
    layer2_outputs(6269) <= not b;
    layer2_outputs(6270) <= b;
    layer2_outputs(6271) <= not a;
    layer2_outputs(6272) <= a;
    layer2_outputs(6273) <= not b;
    layer2_outputs(6274) <= a;
    layer2_outputs(6275) <= not a;
    layer2_outputs(6276) <= not (a xor b);
    layer2_outputs(6277) <= a and b;
    layer2_outputs(6278) <= a and not b;
    layer2_outputs(6279) <= a and b;
    layer2_outputs(6280) <= not b or a;
    layer2_outputs(6281) <= a;
    layer2_outputs(6282) <= a;
    layer2_outputs(6283) <= b;
    layer2_outputs(6284) <= not (a xor b);
    layer2_outputs(6285) <= not (a xor b);
    layer2_outputs(6286) <= b;
    layer2_outputs(6287) <= a and b;
    layer2_outputs(6288) <= a xor b;
    layer2_outputs(6289) <= not (a xor b);
    layer2_outputs(6290) <= not (a and b);
    layer2_outputs(6291) <= a and b;
    layer2_outputs(6292) <= not a;
    layer2_outputs(6293) <= not b;
    layer2_outputs(6294) <= not b;
    layer2_outputs(6295) <= a xor b;
    layer2_outputs(6296) <= a or b;
    layer2_outputs(6297) <= a xor b;
    layer2_outputs(6298) <= not a;
    layer2_outputs(6299) <= not b or a;
    layer2_outputs(6300) <= not a;
    layer2_outputs(6301) <= not b;
    layer2_outputs(6302) <= not (a xor b);
    layer2_outputs(6303) <= not b;
    layer2_outputs(6304) <= b;
    layer2_outputs(6305) <= b and not a;
    layer2_outputs(6306) <= not a;
    layer2_outputs(6307) <= a or b;
    layer2_outputs(6308) <= not a;
    layer2_outputs(6309) <= not (a and b);
    layer2_outputs(6310) <= a and b;
    layer2_outputs(6311) <= a or b;
    layer2_outputs(6312) <= a or b;
    layer2_outputs(6313) <= a xor b;
    layer2_outputs(6314) <= not b;
    layer2_outputs(6315) <= not (a or b);
    layer2_outputs(6316) <= not b;
    layer2_outputs(6317) <= not b;
    layer2_outputs(6318) <= a and b;
    layer2_outputs(6319) <= b;
    layer2_outputs(6320) <= b;
    layer2_outputs(6321) <= a or b;
    layer2_outputs(6322) <= b;
    layer2_outputs(6323) <= not a;
    layer2_outputs(6324) <= not (a xor b);
    layer2_outputs(6325) <= a;
    layer2_outputs(6326) <= not b;
    layer2_outputs(6327) <= not (a xor b);
    layer2_outputs(6328) <= a and not b;
    layer2_outputs(6329) <= not (a xor b);
    layer2_outputs(6330) <= not (a or b);
    layer2_outputs(6331) <= a;
    layer2_outputs(6332) <= not b;
    layer2_outputs(6333) <= b;
    layer2_outputs(6334) <= not b;
    layer2_outputs(6335) <= not a;
    layer2_outputs(6336) <= not (a and b);
    layer2_outputs(6337) <= b;
    layer2_outputs(6338) <= not a;
    layer2_outputs(6339) <= not b;
    layer2_outputs(6340) <= b;
    layer2_outputs(6341) <= not (a and b);
    layer2_outputs(6342) <= a or b;
    layer2_outputs(6343) <= b;
    layer2_outputs(6344) <= a or b;
    layer2_outputs(6345) <= b and not a;
    layer2_outputs(6346) <= not (a and b);
    layer2_outputs(6347) <= not a or b;
    layer2_outputs(6348) <= not a;
    layer2_outputs(6349) <= a;
    layer2_outputs(6350) <= a;
    layer2_outputs(6351) <= a and b;
    layer2_outputs(6352) <= not b;
    layer2_outputs(6353) <= a xor b;
    layer2_outputs(6354) <= b;
    layer2_outputs(6355) <= not b;
    layer2_outputs(6356) <= not a or b;
    layer2_outputs(6357) <= not a;
    layer2_outputs(6358) <= a or b;
    layer2_outputs(6359) <= not (a or b);
    layer2_outputs(6360) <= b;
    layer2_outputs(6361) <= a and b;
    layer2_outputs(6362) <= b and not a;
    layer2_outputs(6363) <= not b or a;
    layer2_outputs(6364) <= not b or a;
    layer2_outputs(6365) <= not a;
    layer2_outputs(6366) <= not b;
    layer2_outputs(6367) <= a xor b;
    layer2_outputs(6368) <= not (a or b);
    layer2_outputs(6369) <= a;
    layer2_outputs(6370) <= not (a or b);
    layer2_outputs(6371) <= not b;
    layer2_outputs(6372) <= b;
    layer2_outputs(6373) <= not (a xor b);
    layer2_outputs(6374) <= not (a or b);
    layer2_outputs(6375) <= a xor b;
    layer2_outputs(6376) <= b and not a;
    layer2_outputs(6377) <= not (a or b);
    layer2_outputs(6378) <= not b;
    layer2_outputs(6379) <= a xor b;
    layer2_outputs(6380) <= not (a xor b);
    layer2_outputs(6381) <= not (a and b);
    layer2_outputs(6382) <= not b;
    layer2_outputs(6383) <= b and not a;
    layer2_outputs(6384) <= not b;
    layer2_outputs(6385) <= not a;
    layer2_outputs(6386) <= not (a and b);
    layer2_outputs(6387) <= not (a xor b);
    layer2_outputs(6388) <= not (a xor b);
    layer2_outputs(6389) <= not b;
    layer2_outputs(6390) <= a;
    layer2_outputs(6391) <= not (a or b);
    layer2_outputs(6392) <= a and not b;
    layer2_outputs(6393) <= not (a xor b);
    layer2_outputs(6394) <= a and b;
    layer2_outputs(6395) <= not (a or b);
    layer2_outputs(6396) <= b;
    layer2_outputs(6397) <= a and b;
    layer2_outputs(6398) <= a;
    layer2_outputs(6399) <= not a;
    layer2_outputs(6400) <= a;
    layer2_outputs(6401) <= not b;
    layer2_outputs(6402) <= a;
    layer2_outputs(6403) <= a or b;
    layer2_outputs(6404) <= not (a and b);
    layer2_outputs(6405) <= not b or a;
    layer2_outputs(6406) <= b;
    layer2_outputs(6407) <= not (a xor b);
    layer2_outputs(6408) <= b and not a;
    layer2_outputs(6409) <= not (a xor b);
    layer2_outputs(6410) <= not (a or b);
    layer2_outputs(6411) <= not (a xor b);
    layer2_outputs(6412) <= a and not b;
    layer2_outputs(6413) <= a or b;
    layer2_outputs(6414) <= a xor b;
    layer2_outputs(6415) <= a;
    layer2_outputs(6416) <= a xor b;
    layer2_outputs(6417) <= not b;
    layer2_outputs(6418) <= a and not b;
    layer2_outputs(6419) <= not b;
    layer2_outputs(6420) <= a;
    layer2_outputs(6421) <= not b;
    layer2_outputs(6422) <= b;
    layer2_outputs(6423) <= not a;
    layer2_outputs(6424) <= not (a and b);
    layer2_outputs(6425) <= a and b;
    layer2_outputs(6426) <= not (a xor b);
    layer2_outputs(6427) <= not a;
    layer2_outputs(6428) <= not (a xor b);
    layer2_outputs(6429) <= not a or b;
    layer2_outputs(6430) <= a;
    layer2_outputs(6431) <= not b;
    layer2_outputs(6432) <= a or b;
    layer2_outputs(6433) <= b and not a;
    layer2_outputs(6434) <= a or b;
    layer2_outputs(6435) <= not (a xor b);
    layer2_outputs(6436) <= not (a xor b);
    layer2_outputs(6437) <= not (a xor b);
    layer2_outputs(6438) <= a;
    layer2_outputs(6439) <= not a;
    layer2_outputs(6440) <= a and not b;
    layer2_outputs(6441) <= not a;
    layer2_outputs(6442) <= not a;
    layer2_outputs(6443) <= a or b;
    layer2_outputs(6444) <= b;
    layer2_outputs(6445) <= a;
    layer2_outputs(6446) <= not (a and b);
    layer2_outputs(6447) <= b;
    layer2_outputs(6448) <= a and not b;
    layer2_outputs(6449) <= not (a or b);
    layer2_outputs(6450) <= b;
    layer2_outputs(6451) <= not b;
    layer2_outputs(6452) <= not (a xor b);
    layer2_outputs(6453) <= not b or a;
    layer2_outputs(6454) <= not (a xor b);
    layer2_outputs(6455) <= a;
    layer2_outputs(6456) <= b;
    layer2_outputs(6457) <= not b or a;
    layer2_outputs(6458) <= a xor b;
    layer2_outputs(6459) <= a;
    layer2_outputs(6460) <= not (a xor b);
    layer2_outputs(6461) <= not (a or b);
    layer2_outputs(6462) <= not (a and b);
    layer2_outputs(6463) <= a and not b;
    layer2_outputs(6464) <= not b;
    layer2_outputs(6465) <= b;
    layer2_outputs(6466) <= not (a or b);
    layer2_outputs(6467) <= a;
    layer2_outputs(6468) <= b and not a;
    layer2_outputs(6469) <= not (a xor b);
    layer2_outputs(6470) <= a;
    layer2_outputs(6471) <= not (a xor b);
    layer2_outputs(6472) <= not (a or b);
    layer2_outputs(6473) <= a and not b;
    layer2_outputs(6474) <= not (a or b);
    layer2_outputs(6475) <= not a;
    layer2_outputs(6476) <= not b or a;
    layer2_outputs(6477) <= not (a xor b);
    layer2_outputs(6478) <= not a;
    layer2_outputs(6479) <= not (a and b);
    layer2_outputs(6480) <= b;
    layer2_outputs(6481) <= not (a xor b);
    layer2_outputs(6482) <= a and not b;
    layer2_outputs(6483) <= not b;
    layer2_outputs(6484) <= b and not a;
    layer2_outputs(6485) <= a and not b;
    layer2_outputs(6486) <= a;
    layer2_outputs(6487) <= 1'b1;
    layer2_outputs(6488) <= not (a and b);
    layer2_outputs(6489) <= not b;
    layer2_outputs(6490) <= a;
    layer2_outputs(6491) <= not (a or b);
    layer2_outputs(6492) <= 1'b1;
    layer2_outputs(6493) <= not a;
    layer2_outputs(6494) <= a xor b;
    layer2_outputs(6495) <= a and not b;
    layer2_outputs(6496) <= a xor b;
    layer2_outputs(6497) <= a;
    layer2_outputs(6498) <= a or b;
    layer2_outputs(6499) <= 1'b0;
    layer2_outputs(6500) <= not (a xor b);
    layer2_outputs(6501) <= not b or a;
    layer2_outputs(6502) <= not (a or b);
    layer2_outputs(6503) <= a or b;
    layer2_outputs(6504) <= not (a and b);
    layer2_outputs(6505) <= not (a xor b);
    layer2_outputs(6506) <= not (a or b);
    layer2_outputs(6507) <= b;
    layer2_outputs(6508) <= a xor b;
    layer2_outputs(6509) <= b;
    layer2_outputs(6510) <= a and not b;
    layer2_outputs(6511) <= a xor b;
    layer2_outputs(6512) <= a and not b;
    layer2_outputs(6513) <= not (a and b);
    layer2_outputs(6514) <= not (a xor b);
    layer2_outputs(6515) <= not b;
    layer2_outputs(6516) <= a and b;
    layer2_outputs(6517) <= a;
    layer2_outputs(6518) <= not a or b;
    layer2_outputs(6519) <= b and not a;
    layer2_outputs(6520) <= b and not a;
    layer2_outputs(6521) <= not a;
    layer2_outputs(6522) <= a;
    layer2_outputs(6523) <= b and not a;
    layer2_outputs(6524) <= not (a and b);
    layer2_outputs(6525) <= not (a and b);
    layer2_outputs(6526) <= not b;
    layer2_outputs(6527) <= a xor b;
    layer2_outputs(6528) <= a;
    layer2_outputs(6529) <= not a;
    layer2_outputs(6530) <= not (a or b);
    layer2_outputs(6531) <= not (a xor b);
    layer2_outputs(6532) <= not (a and b);
    layer2_outputs(6533) <= not (a or b);
    layer2_outputs(6534) <= a or b;
    layer2_outputs(6535) <= not b;
    layer2_outputs(6536) <= a xor b;
    layer2_outputs(6537) <= not a;
    layer2_outputs(6538) <= not a;
    layer2_outputs(6539) <= b and not a;
    layer2_outputs(6540) <= a and b;
    layer2_outputs(6541) <= a and not b;
    layer2_outputs(6542) <= b and not a;
    layer2_outputs(6543) <= not b or a;
    layer2_outputs(6544) <= not (a and b);
    layer2_outputs(6545) <= a or b;
    layer2_outputs(6546) <= b and not a;
    layer2_outputs(6547) <= a and not b;
    layer2_outputs(6548) <= not b;
    layer2_outputs(6549) <= a xor b;
    layer2_outputs(6550) <= b and not a;
    layer2_outputs(6551) <= not b or a;
    layer2_outputs(6552) <= not b;
    layer2_outputs(6553) <= not (a xor b);
    layer2_outputs(6554) <= not (a or b);
    layer2_outputs(6555) <= not b;
    layer2_outputs(6556) <= not (a and b);
    layer2_outputs(6557) <= b;
    layer2_outputs(6558) <= a;
    layer2_outputs(6559) <= not (a xor b);
    layer2_outputs(6560) <= b and not a;
    layer2_outputs(6561) <= not a or b;
    layer2_outputs(6562) <= not a;
    layer2_outputs(6563) <= a and b;
    layer2_outputs(6564) <= a xor b;
    layer2_outputs(6565) <= not (a or b);
    layer2_outputs(6566) <= a;
    layer2_outputs(6567) <= not b;
    layer2_outputs(6568) <= a or b;
    layer2_outputs(6569) <= not a;
    layer2_outputs(6570) <= a;
    layer2_outputs(6571) <= not a or b;
    layer2_outputs(6572) <= not b;
    layer2_outputs(6573) <= not (a and b);
    layer2_outputs(6574) <= a and b;
    layer2_outputs(6575) <= not (a xor b);
    layer2_outputs(6576) <= b and not a;
    layer2_outputs(6577) <= a xor b;
    layer2_outputs(6578) <= not a;
    layer2_outputs(6579) <= a xor b;
    layer2_outputs(6580) <= a;
    layer2_outputs(6581) <= a and b;
    layer2_outputs(6582) <= not (a or b);
    layer2_outputs(6583) <= a;
    layer2_outputs(6584) <= a;
    layer2_outputs(6585) <= a;
    layer2_outputs(6586) <= a and b;
    layer2_outputs(6587) <= not a;
    layer2_outputs(6588) <= b;
    layer2_outputs(6589) <= not a or b;
    layer2_outputs(6590) <= not (a or b);
    layer2_outputs(6591) <= a and not b;
    layer2_outputs(6592) <= not (a or b);
    layer2_outputs(6593) <= not a;
    layer2_outputs(6594) <= not b or a;
    layer2_outputs(6595) <= not b or a;
    layer2_outputs(6596) <= not b;
    layer2_outputs(6597) <= not (a xor b);
    layer2_outputs(6598) <= not a;
    layer2_outputs(6599) <= not b;
    layer2_outputs(6600) <= a and not b;
    layer2_outputs(6601) <= not b or a;
    layer2_outputs(6602) <= a xor b;
    layer2_outputs(6603) <= not (a and b);
    layer2_outputs(6604) <= a;
    layer2_outputs(6605) <= not b;
    layer2_outputs(6606) <= b;
    layer2_outputs(6607) <= a xor b;
    layer2_outputs(6608) <= not a;
    layer2_outputs(6609) <= not b;
    layer2_outputs(6610) <= not b or a;
    layer2_outputs(6611) <= a;
    layer2_outputs(6612) <= not a or b;
    layer2_outputs(6613) <= not a or b;
    layer2_outputs(6614) <= not a;
    layer2_outputs(6615) <= a or b;
    layer2_outputs(6616) <= a xor b;
    layer2_outputs(6617) <= not b;
    layer2_outputs(6618) <= not a or b;
    layer2_outputs(6619) <= not (a xor b);
    layer2_outputs(6620) <= not b or a;
    layer2_outputs(6621) <= not a;
    layer2_outputs(6622) <= a and not b;
    layer2_outputs(6623) <= not b;
    layer2_outputs(6624) <= not (a or b);
    layer2_outputs(6625) <= not b;
    layer2_outputs(6626) <= 1'b0;
    layer2_outputs(6627) <= a;
    layer2_outputs(6628) <= a or b;
    layer2_outputs(6629) <= not (a xor b);
    layer2_outputs(6630) <= not a;
    layer2_outputs(6631) <= not b or a;
    layer2_outputs(6632) <= a;
    layer2_outputs(6633) <= not b;
    layer2_outputs(6634) <= a or b;
    layer2_outputs(6635) <= b and not a;
    layer2_outputs(6636) <= not (a and b);
    layer2_outputs(6637) <= not b;
    layer2_outputs(6638) <= b;
    layer2_outputs(6639) <= a;
    layer2_outputs(6640) <= b;
    layer2_outputs(6641) <= not a;
    layer2_outputs(6642) <= b;
    layer2_outputs(6643) <= a and not b;
    layer2_outputs(6644) <= b;
    layer2_outputs(6645) <= b;
    layer2_outputs(6646) <= a;
    layer2_outputs(6647) <= not b;
    layer2_outputs(6648) <= not (a or b);
    layer2_outputs(6649) <= a;
    layer2_outputs(6650) <= b;
    layer2_outputs(6651) <= not a;
    layer2_outputs(6652) <= a or b;
    layer2_outputs(6653) <= not (a and b);
    layer2_outputs(6654) <= a and b;
    layer2_outputs(6655) <= not b;
    layer2_outputs(6656) <= not (a xor b);
    layer2_outputs(6657) <= not a;
    layer2_outputs(6658) <= 1'b0;
    layer2_outputs(6659) <= not b;
    layer2_outputs(6660) <= not a or b;
    layer2_outputs(6661) <= not b;
    layer2_outputs(6662) <= not (a or b);
    layer2_outputs(6663) <= a and not b;
    layer2_outputs(6664) <= a or b;
    layer2_outputs(6665) <= a and not b;
    layer2_outputs(6666) <= a and b;
    layer2_outputs(6667) <= a and b;
    layer2_outputs(6668) <= not (a or b);
    layer2_outputs(6669) <= a xor b;
    layer2_outputs(6670) <= b;
    layer2_outputs(6671) <= not b;
    layer2_outputs(6672) <= not (a and b);
    layer2_outputs(6673) <= not (a xor b);
    layer2_outputs(6674) <= a;
    layer2_outputs(6675) <= a xor b;
    layer2_outputs(6676) <= not a or b;
    layer2_outputs(6677) <= a;
    layer2_outputs(6678) <= a xor b;
    layer2_outputs(6679) <= not a;
    layer2_outputs(6680) <= not (a and b);
    layer2_outputs(6681) <= b;
    layer2_outputs(6682) <= not b;
    layer2_outputs(6683) <= a;
    layer2_outputs(6684) <= not (a xor b);
    layer2_outputs(6685) <= not a or b;
    layer2_outputs(6686) <= not a;
    layer2_outputs(6687) <= not b or a;
    layer2_outputs(6688) <= not a;
    layer2_outputs(6689) <= not (a and b);
    layer2_outputs(6690) <= not b or a;
    layer2_outputs(6691) <= not a;
    layer2_outputs(6692) <= b;
    layer2_outputs(6693) <= a xor b;
    layer2_outputs(6694) <= b;
    layer2_outputs(6695) <= not a;
    layer2_outputs(6696) <= not b;
    layer2_outputs(6697) <= a and not b;
    layer2_outputs(6698) <= a xor b;
    layer2_outputs(6699) <= not a;
    layer2_outputs(6700) <= a;
    layer2_outputs(6701) <= b and not a;
    layer2_outputs(6702) <= not (a and b);
    layer2_outputs(6703) <= not a or b;
    layer2_outputs(6704) <= b and not a;
    layer2_outputs(6705) <= not a;
    layer2_outputs(6706) <= not (a xor b);
    layer2_outputs(6707) <= a and b;
    layer2_outputs(6708) <= a xor b;
    layer2_outputs(6709) <= not a or b;
    layer2_outputs(6710) <= a xor b;
    layer2_outputs(6711) <= not (a xor b);
    layer2_outputs(6712) <= a and b;
    layer2_outputs(6713) <= not (a or b);
    layer2_outputs(6714) <= not (a or b);
    layer2_outputs(6715) <= a and not b;
    layer2_outputs(6716) <= not a;
    layer2_outputs(6717) <= not b or a;
    layer2_outputs(6718) <= not a or b;
    layer2_outputs(6719) <= b;
    layer2_outputs(6720) <= b;
    layer2_outputs(6721) <= b;
    layer2_outputs(6722) <= a xor b;
    layer2_outputs(6723) <= a xor b;
    layer2_outputs(6724) <= a xor b;
    layer2_outputs(6725) <= a xor b;
    layer2_outputs(6726) <= a;
    layer2_outputs(6727) <= a xor b;
    layer2_outputs(6728) <= not (a and b);
    layer2_outputs(6729) <= a or b;
    layer2_outputs(6730) <= a or b;
    layer2_outputs(6731) <= not (a or b);
    layer2_outputs(6732) <= not a;
    layer2_outputs(6733) <= a xor b;
    layer2_outputs(6734) <= not a;
    layer2_outputs(6735) <= not (a xor b);
    layer2_outputs(6736) <= b;
    layer2_outputs(6737) <= a;
    layer2_outputs(6738) <= b;
    layer2_outputs(6739) <= b and not a;
    layer2_outputs(6740) <= a;
    layer2_outputs(6741) <= not a;
    layer2_outputs(6742) <= not b or a;
    layer2_outputs(6743) <= b;
    layer2_outputs(6744) <= not a or b;
    layer2_outputs(6745) <= not (a and b);
    layer2_outputs(6746) <= a;
    layer2_outputs(6747) <= a xor b;
    layer2_outputs(6748) <= not (a xor b);
    layer2_outputs(6749) <= a xor b;
    layer2_outputs(6750) <= a and not b;
    layer2_outputs(6751) <= b;
    layer2_outputs(6752) <= a;
    layer2_outputs(6753) <= not a or b;
    layer2_outputs(6754) <= a and not b;
    layer2_outputs(6755) <= not a;
    layer2_outputs(6756) <= not (a xor b);
    layer2_outputs(6757) <= a xor b;
    layer2_outputs(6758) <= not (a xor b);
    layer2_outputs(6759) <= not b;
    layer2_outputs(6760) <= not (a xor b);
    layer2_outputs(6761) <= b;
    layer2_outputs(6762) <= a xor b;
    layer2_outputs(6763) <= not a;
    layer2_outputs(6764) <= a and b;
    layer2_outputs(6765) <= not a;
    layer2_outputs(6766) <= not b or a;
    layer2_outputs(6767) <= b;
    layer2_outputs(6768) <= a xor b;
    layer2_outputs(6769) <= not b;
    layer2_outputs(6770) <= not a;
    layer2_outputs(6771) <= b;
    layer2_outputs(6772) <= a or b;
    layer2_outputs(6773) <= a;
    layer2_outputs(6774) <= not a;
    layer2_outputs(6775) <= b;
    layer2_outputs(6776) <= a and not b;
    layer2_outputs(6777) <= a xor b;
    layer2_outputs(6778) <= not (a or b);
    layer2_outputs(6779) <= b and not a;
    layer2_outputs(6780) <= a;
    layer2_outputs(6781) <= a;
    layer2_outputs(6782) <= not (a xor b);
    layer2_outputs(6783) <= not (a xor b);
    layer2_outputs(6784) <= a or b;
    layer2_outputs(6785) <= not (a xor b);
    layer2_outputs(6786) <= not b;
    layer2_outputs(6787) <= not (a and b);
    layer2_outputs(6788) <= not (a and b);
    layer2_outputs(6789) <= not a or b;
    layer2_outputs(6790) <= a xor b;
    layer2_outputs(6791) <= not a;
    layer2_outputs(6792) <= not b;
    layer2_outputs(6793) <= a and not b;
    layer2_outputs(6794) <= a xor b;
    layer2_outputs(6795) <= b;
    layer2_outputs(6796) <= not b;
    layer2_outputs(6797) <= a;
    layer2_outputs(6798) <= not a or b;
    layer2_outputs(6799) <= not b or a;
    layer2_outputs(6800) <= b;
    layer2_outputs(6801) <= not (a xor b);
    layer2_outputs(6802) <= not (a xor b);
    layer2_outputs(6803) <= a xor b;
    layer2_outputs(6804) <= a and not b;
    layer2_outputs(6805) <= b;
    layer2_outputs(6806) <= b and not a;
    layer2_outputs(6807) <= not b or a;
    layer2_outputs(6808) <= not (a and b);
    layer2_outputs(6809) <= not b;
    layer2_outputs(6810) <= not b;
    layer2_outputs(6811) <= a xor b;
    layer2_outputs(6812) <= a xor b;
    layer2_outputs(6813) <= not b or a;
    layer2_outputs(6814) <= not b;
    layer2_outputs(6815) <= a xor b;
    layer2_outputs(6816) <= not a;
    layer2_outputs(6817) <= not (a or b);
    layer2_outputs(6818) <= not (a and b);
    layer2_outputs(6819) <= b and not a;
    layer2_outputs(6820) <= a xor b;
    layer2_outputs(6821) <= b;
    layer2_outputs(6822) <= b;
    layer2_outputs(6823) <= not (a xor b);
    layer2_outputs(6824) <= a;
    layer2_outputs(6825) <= not b;
    layer2_outputs(6826) <= a;
    layer2_outputs(6827) <= not b or a;
    layer2_outputs(6828) <= a;
    layer2_outputs(6829) <= not b;
    layer2_outputs(6830) <= a;
    layer2_outputs(6831) <= b;
    layer2_outputs(6832) <= not a;
    layer2_outputs(6833) <= not b;
    layer2_outputs(6834) <= a and not b;
    layer2_outputs(6835) <= b;
    layer2_outputs(6836) <= b;
    layer2_outputs(6837) <= not b;
    layer2_outputs(6838) <= a xor b;
    layer2_outputs(6839) <= not a;
    layer2_outputs(6840) <= not (a xor b);
    layer2_outputs(6841) <= a xor b;
    layer2_outputs(6842) <= b;
    layer2_outputs(6843) <= a or b;
    layer2_outputs(6844) <= not (a xor b);
    layer2_outputs(6845) <= a or b;
    layer2_outputs(6846) <= not a;
    layer2_outputs(6847) <= not a;
    layer2_outputs(6848) <= not (a and b);
    layer2_outputs(6849) <= not b or a;
    layer2_outputs(6850) <= not b;
    layer2_outputs(6851) <= a and b;
    layer2_outputs(6852) <= b;
    layer2_outputs(6853) <= not a;
    layer2_outputs(6854) <= not b;
    layer2_outputs(6855) <= not b;
    layer2_outputs(6856) <= a or b;
    layer2_outputs(6857) <= a xor b;
    layer2_outputs(6858) <= a or b;
    layer2_outputs(6859) <= b;
    layer2_outputs(6860) <= 1'b0;
    layer2_outputs(6861) <= not b;
    layer2_outputs(6862) <= not b or a;
    layer2_outputs(6863) <= not (a and b);
    layer2_outputs(6864) <= a and b;
    layer2_outputs(6865) <= not (a and b);
    layer2_outputs(6866) <= not a;
    layer2_outputs(6867) <= not b;
    layer2_outputs(6868) <= b;
    layer2_outputs(6869) <= a and not b;
    layer2_outputs(6870) <= not b;
    layer2_outputs(6871) <= b and not a;
    layer2_outputs(6872) <= b;
    layer2_outputs(6873) <= not (a xor b);
    layer2_outputs(6874) <= not a or b;
    layer2_outputs(6875) <= not a;
    layer2_outputs(6876) <= not a or b;
    layer2_outputs(6877) <= b and not a;
    layer2_outputs(6878) <= not a;
    layer2_outputs(6879) <= not (a or b);
    layer2_outputs(6880) <= a xor b;
    layer2_outputs(6881) <= not b or a;
    layer2_outputs(6882) <= not (a xor b);
    layer2_outputs(6883) <= a xor b;
    layer2_outputs(6884) <= not (a or b);
    layer2_outputs(6885) <= not (a and b);
    layer2_outputs(6886) <= not (a and b);
    layer2_outputs(6887) <= a;
    layer2_outputs(6888) <= a and not b;
    layer2_outputs(6889) <= not a;
    layer2_outputs(6890) <= not a or b;
    layer2_outputs(6891) <= not b;
    layer2_outputs(6892) <= a or b;
    layer2_outputs(6893) <= a and b;
    layer2_outputs(6894) <= not (a or b);
    layer2_outputs(6895) <= a;
    layer2_outputs(6896) <= b;
    layer2_outputs(6897) <= a and not b;
    layer2_outputs(6898) <= a and not b;
    layer2_outputs(6899) <= not a;
    layer2_outputs(6900) <= a and not b;
    layer2_outputs(6901) <= not a;
    layer2_outputs(6902) <= not b;
    layer2_outputs(6903) <= b and not a;
    layer2_outputs(6904) <= a xor b;
    layer2_outputs(6905) <= a and not b;
    layer2_outputs(6906) <= not b or a;
    layer2_outputs(6907) <= not a;
    layer2_outputs(6908) <= a;
    layer2_outputs(6909) <= a and b;
    layer2_outputs(6910) <= not b;
    layer2_outputs(6911) <= not b;
    layer2_outputs(6912) <= a and b;
    layer2_outputs(6913) <= not b;
    layer2_outputs(6914) <= a xor b;
    layer2_outputs(6915) <= not (a and b);
    layer2_outputs(6916) <= not b;
    layer2_outputs(6917) <= a and b;
    layer2_outputs(6918) <= a;
    layer2_outputs(6919) <= not b;
    layer2_outputs(6920) <= not a or b;
    layer2_outputs(6921) <= b;
    layer2_outputs(6922) <= b and not a;
    layer2_outputs(6923) <= not (a or b);
    layer2_outputs(6924) <= a;
    layer2_outputs(6925) <= not b;
    layer2_outputs(6926) <= not (a xor b);
    layer2_outputs(6927) <= b;
    layer2_outputs(6928) <= not b;
    layer2_outputs(6929) <= a xor b;
    layer2_outputs(6930) <= b;
    layer2_outputs(6931) <= a or b;
    layer2_outputs(6932) <= a xor b;
    layer2_outputs(6933) <= a and b;
    layer2_outputs(6934) <= a xor b;
    layer2_outputs(6935) <= a xor b;
    layer2_outputs(6936) <= a xor b;
    layer2_outputs(6937) <= a xor b;
    layer2_outputs(6938) <= a or b;
    layer2_outputs(6939) <= not a;
    layer2_outputs(6940) <= not b;
    layer2_outputs(6941) <= b;
    layer2_outputs(6942) <= a and b;
    layer2_outputs(6943) <= a xor b;
    layer2_outputs(6944) <= not (a xor b);
    layer2_outputs(6945) <= a xor b;
    layer2_outputs(6946) <= not b;
    layer2_outputs(6947) <= a and b;
    layer2_outputs(6948) <= not b;
    layer2_outputs(6949) <= not a;
    layer2_outputs(6950) <= not b;
    layer2_outputs(6951) <= b;
    layer2_outputs(6952) <= not a;
    layer2_outputs(6953) <= not a;
    layer2_outputs(6954) <= not (a or b);
    layer2_outputs(6955) <= a xor b;
    layer2_outputs(6956) <= b;
    layer2_outputs(6957) <= b;
    layer2_outputs(6958) <= not b or a;
    layer2_outputs(6959) <= a;
    layer2_outputs(6960) <= not b;
    layer2_outputs(6961) <= not a;
    layer2_outputs(6962) <= a and b;
    layer2_outputs(6963) <= a;
    layer2_outputs(6964) <= not (a xor b);
    layer2_outputs(6965) <= not a;
    layer2_outputs(6966) <= a;
    layer2_outputs(6967) <= a;
    layer2_outputs(6968) <= not (a or b);
    layer2_outputs(6969) <= not b;
    layer2_outputs(6970) <= a xor b;
    layer2_outputs(6971) <= not a;
    layer2_outputs(6972) <= not b;
    layer2_outputs(6973) <= not a;
    layer2_outputs(6974) <= a or b;
    layer2_outputs(6975) <= a xor b;
    layer2_outputs(6976) <= a or b;
    layer2_outputs(6977) <= a xor b;
    layer2_outputs(6978) <= a xor b;
    layer2_outputs(6979) <= not (a xor b);
    layer2_outputs(6980) <= a;
    layer2_outputs(6981) <= not b;
    layer2_outputs(6982) <= b;
    layer2_outputs(6983) <= not b or a;
    layer2_outputs(6984) <= not (a xor b);
    layer2_outputs(6985) <= not (a and b);
    layer2_outputs(6986) <= a or b;
    layer2_outputs(6987) <= a;
    layer2_outputs(6988) <= a or b;
    layer2_outputs(6989) <= not b;
    layer2_outputs(6990) <= not (a or b);
    layer2_outputs(6991) <= not b;
    layer2_outputs(6992) <= not b;
    layer2_outputs(6993) <= not a;
    layer2_outputs(6994) <= not b;
    layer2_outputs(6995) <= not b;
    layer2_outputs(6996) <= a xor b;
    layer2_outputs(6997) <= a and not b;
    layer2_outputs(6998) <= b and not a;
    layer2_outputs(6999) <= not b;
    layer2_outputs(7000) <= not b or a;
    layer2_outputs(7001) <= not (a and b);
    layer2_outputs(7002) <= not a;
    layer2_outputs(7003) <= not a;
    layer2_outputs(7004) <= not (a xor b);
    layer2_outputs(7005) <= not a;
    layer2_outputs(7006) <= not a or b;
    layer2_outputs(7007) <= b and not a;
    layer2_outputs(7008) <= not b;
    layer2_outputs(7009) <= not a;
    layer2_outputs(7010) <= not (a or b);
    layer2_outputs(7011) <= not a;
    layer2_outputs(7012) <= not a;
    layer2_outputs(7013) <= a;
    layer2_outputs(7014) <= b;
    layer2_outputs(7015) <= not b;
    layer2_outputs(7016) <= not a;
    layer2_outputs(7017) <= b;
    layer2_outputs(7018) <= not b or a;
    layer2_outputs(7019) <= a;
    layer2_outputs(7020) <= not b;
    layer2_outputs(7021) <= a and not b;
    layer2_outputs(7022) <= not (a xor b);
    layer2_outputs(7023) <= a and not b;
    layer2_outputs(7024) <= a;
    layer2_outputs(7025) <= not b or a;
    layer2_outputs(7026) <= not a;
    layer2_outputs(7027) <= not b;
    layer2_outputs(7028) <= a xor b;
    layer2_outputs(7029) <= not (a or b);
    layer2_outputs(7030) <= not (a and b);
    layer2_outputs(7031) <= b;
    layer2_outputs(7032) <= b and not a;
    layer2_outputs(7033) <= a xor b;
    layer2_outputs(7034) <= not a;
    layer2_outputs(7035) <= a or b;
    layer2_outputs(7036) <= not b;
    layer2_outputs(7037) <= not a;
    layer2_outputs(7038) <= not a;
    layer2_outputs(7039) <= not (a or b);
    layer2_outputs(7040) <= not b;
    layer2_outputs(7041) <= b;
    layer2_outputs(7042) <= not b;
    layer2_outputs(7043) <= not a;
    layer2_outputs(7044) <= b;
    layer2_outputs(7045) <= a xor b;
    layer2_outputs(7046) <= a;
    layer2_outputs(7047) <= not (a xor b);
    layer2_outputs(7048) <= b;
    layer2_outputs(7049) <= b;
    layer2_outputs(7050) <= not a;
    layer2_outputs(7051) <= a or b;
    layer2_outputs(7052) <= not b;
    layer2_outputs(7053) <= b and not a;
    layer2_outputs(7054) <= a and b;
    layer2_outputs(7055) <= not b or a;
    layer2_outputs(7056) <= a;
    layer2_outputs(7057) <= not (a xor b);
    layer2_outputs(7058) <= not a;
    layer2_outputs(7059) <= a or b;
    layer2_outputs(7060) <= a xor b;
    layer2_outputs(7061) <= not (a and b);
    layer2_outputs(7062) <= a and not b;
    layer2_outputs(7063) <= not (a and b);
    layer2_outputs(7064) <= not a;
    layer2_outputs(7065) <= not a;
    layer2_outputs(7066) <= not b;
    layer2_outputs(7067) <= not (a xor b);
    layer2_outputs(7068) <= not a;
    layer2_outputs(7069) <= not b;
    layer2_outputs(7070) <= not b;
    layer2_outputs(7071) <= not (a and b);
    layer2_outputs(7072) <= not a;
    layer2_outputs(7073) <= not (a or b);
    layer2_outputs(7074) <= not (a xor b);
    layer2_outputs(7075) <= not a;
    layer2_outputs(7076) <= a or b;
    layer2_outputs(7077) <= not (a xor b);
    layer2_outputs(7078) <= not a or b;
    layer2_outputs(7079) <= not b or a;
    layer2_outputs(7080) <= a xor b;
    layer2_outputs(7081) <= a and b;
    layer2_outputs(7082) <= not a or b;
    layer2_outputs(7083) <= a and not b;
    layer2_outputs(7084) <= not b;
    layer2_outputs(7085) <= a;
    layer2_outputs(7086) <= not a;
    layer2_outputs(7087) <= not b;
    layer2_outputs(7088) <= b;
    layer2_outputs(7089) <= a;
    layer2_outputs(7090) <= not b;
    layer2_outputs(7091) <= a;
    layer2_outputs(7092) <= not (a xor b);
    layer2_outputs(7093) <= b and not a;
    layer2_outputs(7094) <= not a;
    layer2_outputs(7095) <= a xor b;
    layer2_outputs(7096) <= a;
    layer2_outputs(7097) <= a xor b;
    layer2_outputs(7098) <= not (a xor b);
    layer2_outputs(7099) <= not (a xor b);
    layer2_outputs(7100) <= a;
    layer2_outputs(7101) <= not b or a;
    layer2_outputs(7102) <= a and not b;
    layer2_outputs(7103) <= not b;
    layer2_outputs(7104) <= a or b;
    layer2_outputs(7105) <= a and not b;
    layer2_outputs(7106) <= not b;
    layer2_outputs(7107) <= a or b;
    layer2_outputs(7108) <= not a;
    layer2_outputs(7109) <= b and not a;
    layer2_outputs(7110) <= not (a and b);
    layer2_outputs(7111) <= not (a and b);
    layer2_outputs(7112) <= not (a and b);
    layer2_outputs(7113) <= not b;
    layer2_outputs(7114) <= not a;
    layer2_outputs(7115) <= not (a and b);
    layer2_outputs(7116) <= not a or b;
    layer2_outputs(7117) <= not a;
    layer2_outputs(7118) <= a;
    layer2_outputs(7119) <= not a;
    layer2_outputs(7120) <= not b;
    layer2_outputs(7121) <= b and not a;
    layer2_outputs(7122) <= a;
    layer2_outputs(7123) <= not b;
    layer2_outputs(7124) <= not a or b;
    layer2_outputs(7125) <= a xor b;
    layer2_outputs(7126) <= a xor b;
    layer2_outputs(7127) <= b;
    layer2_outputs(7128) <= b and not a;
    layer2_outputs(7129) <= b;
    layer2_outputs(7130) <= a xor b;
    layer2_outputs(7131) <= a or b;
    layer2_outputs(7132) <= not (a xor b);
    layer2_outputs(7133) <= not a;
    layer2_outputs(7134) <= not (a and b);
    layer2_outputs(7135) <= not b;
    layer2_outputs(7136) <= b;
    layer2_outputs(7137) <= b;
    layer2_outputs(7138) <= not b;
    layer2_outputs(7139) <= a xor b;
    layer2_outputs(7140) <= not (a and b);
    layer2_outputs(7141) <= not b or a;
    layer2_outputs(7142) <= b;
    layer2_outputs(7143) <= not a or b;
    layer2_outputs(7144) <= a xor b;
    layer2_outputs(7145) <= not a;
    layer2_outputs(7146) <= b;
    layer2_outputs(7147) <= not a or b;
    layer2_outputs(7148) <= not b or a;
    layer2_outputs(7149) <= a xor b;
    layer2_outputs(7150) <= not (a and b);
    layer2_outputs(7151) <= not (a xor b);
    layer2_outputs(7152) <= not (a and b);
    layer2_outputs(7153) <= a and b;
    layer2_outputs(7154) <= a;
    layer2_outputs(7155) <= b and not a;
    layer2_outputs(7156) <= not (a and b);
    layer2_outputs(7157) <= a and not b;
    layer2_outputs(7158) <= not a;
    layer2_outputs(7159) <= a and not b;
    layer2_outputs(7160) <= not (a or b);
    layer2_outputs(7161) <= not a;
    layer2_outputs(7162) <= not b or a;
    layer2_outputs(7163) <= a and not b;
    layer2_outputs(7164) <= a xor b;
    layer2_outputs(7165) <= not (a xor b);
    layer2_outputs(7166) <= not b or a;
    layer2_outputs(7167) <= b;
    layer2_outputs(7168) <= a;
    layer2_outputs(7169) <= not (a xor b);
    layer2_outputs(7170) <= not (a and b);
    layer2_outputs(7171) <= a and b;
    layer2_outputs(7172) <= not a or b;
    layer2_outputs(7173) <= b;
    layer2_outputs(7174) <= a and b;
    layer2_outputs(7175) <= not a;
    layer2_outputs(7176) <= not a or b;
    layer2_outputs(7177) <= b;
    layer2_outputs(7178) <= not (a xor b);
    layer2_outputs(7179) <= not (a and b);
    layer2_outputs(7180) <= not a;
    layer2_outputs(7181) <= not b;
    layer2_outputs(7182) <= b;
    layer2_outputs(7183) <= not b;
    layer2_outputs(7184) <= not b;
    layer2_outputs(7185) <= not b;
    layer2_outputs(7186) <= b and not a;
    layer2_outputs(7187) <= a;
    layer2_outputs(7188) <= a;
    layer2_outputs(7189) <= b;
    layer2_outputs(7190) <= a or b;
    layer2_outputs(7191) <= a or b;
    layer2_outputs(7192) <= b;
    layer2_outputs(7193) <= not (a xor b);
    layer2_outputs(7194) <= b;
    layer2_outputs(7195) <= not a or b;
    layer2_outputs(7196) <= a;
    layer2_outputs(7197) <= not (a and b);
    layer2_outputs(7198) <= not a;
    layer2_outputs(7199) <= a;
    layer2_outputs(7200) <= a or b;
    layer2_outputs(7201) <= not (a or b);
    layer2_outputs(7202) <= not b;
    layer2_outputs(7203) <= a or b;
    layer2_outputs(7204) <= b and not a;
    layer2_outputs(7205) <= b;
    layer2_outputs(7206) <= a;
    layer2_outputs(7207) <= not (a and b);
    layer2_outputs(7208) <= a;
    layer2_outputs(7209) <= not (a xor b);
    layer2_outputs(7210) <= not b;
    layer2_outputs(7211) <= b and not a;
    layer2_outputs(7212) <= not b or a;
    layer2_outputs(7213) <= not (a or b);
    layer2_outputs(7214) <= not (a xor b);
    layer2_outputs(7215) <= a or b;
    layer2_outputs(7216) <= a xor b;
    layer2_outputs(7217) <= b and not a;
    layer2_outputs(7218) <= not (a and b);
    layer2_outputs(7219) <= a;
    layer2_outputs(7220) <= not b;
    layer2_outputs(7221) <= a xor b;
    layer2_outputs(7222) <= b;
    layer2_outputs(7223) <= not a;
    layer2_outputs(7224) <= b;
    layer2_outputs(7225) <= not b;
    layer2_outputs(7226) <= a;
    layer2_outputs(7227) <= not a;
    layer2_outputs(7228) <= not b;
    layer2_outputs(7229) <= a and not b;
    layer2_outputs(7230) <= not (a or b);
    layer2_outputs(7231) <= b and not a;
    layer2_outputs(7232) <= not b;
    layer2_outputs(7233) <= not (a xor b);
    layer2_outputs(7234) <= not a;
    layer2_outputs(7235) <= b and not a;
    layer2_outputs(7236) <= not (a xor b);
    layer2_outputs(7237) <= not (a xor b);
    layer2_outputs(7238) <= a and b;
    layer2_outputs(7239) <= not a or b;
    layer2_outputs(7240) <= not (a xor b);
    layer2_outputs(7241) <= not (a xor b);
    layer2_outputs(7242) <= not b;
    layer2_outputs(7243) <= not (a xor b);
    layer2_outputs(7244) <= not a;
    layer2_outputs(7245) <= b and not a;
    layer2_outputs(7246) <= a xor b;
    layer2_outputs(7247) <= b;
    layer2_outputs(7248) <= a xor b;
    layer2_outputs(7249) <= b;
    layer2_outputs(7250) <= a;
    layer2_outputs(7251) <= not b or a;
    layer2_outputs(7252) <= not (a and b);
    layer2_outputs(7253) <= a and not b;
    layer2_outputs(7254) <= a and b;
    layer2_outputs(7255) <= a;
    layer2_outputs(7256) <= a xor b;
    layer2_outputs(7257) <= 1'b1;
    layer2_outputs(7258) <= b;
    layer2_outputs(7259) <= a xor b;
    layer2_outputs(7260) <= not b;
    layer2_outputs(7261) <= not (a and b);
    layer2_outputs(7262) <= not b;
    layer2_outputs(7263) <= not (a or b);
    layer2_outputs(7264) <= not a or b;
    layer2_outputs(7265) <= a;
    layer2_outputs(7266) <= not b or a;
    layer2_outputs(7267) <= not a;
    layer2_outputs(7268) <= b;
    layer2_outputs(7269) <= not b or a;
    layer2_outputs(7270) <= a or b;
    layer2_outputs(7271) <= a;
    layer2_outputs(7272) <= not a;
    layer2_outputs(7273) <= not a;
    layer2_outputs(7274) <= not (a and b);
    layer2_outputs(7275) <= not a;
    layer2_outputs(7276) <= b;
    layer2_outputs(7277) <= not a or b;
    layer2_outputs(7278) <= not a or b;
    layer2_outputs(7279) <= not b;
    layer2_outputs(7280) <= not b;
    layer2_outputs(7281) <= not a;
    layer2_outputs(7282) <= not a;
    layer2_outputs(7283) <= not (a or b);
    layer2_outputs(7284) <= not (a and b);
    layer2_outputs(7285) <= not b;
    layer2_outputs(7286) <= a;
    layer2_outputs(7287) <= a xor b;
    layer2_outputs(7288) <= b and not a;
    layer2_outputs(7289) <= a xor b;
    layer2_outputs(7290) <= a;
    layer2_outputs(7291) <= a xor b;
    layer2_outputs(7292) <= 1'b1;
    layer2_outputs(7293) <= b;
    layer2_outputs(7294) <= a;
    layer2_outputs(7295) <= not (a or b);
    layer2_outputs(7296) <= b and not a;
    layer2_outputs(7297) <= not (a or b);
    layer2_outputs(7298) <= not a;
    layer2_outputs(7299) <= not b;
    layer2_outputs(7300) <= not (a xor b);
    layer2_outputs(7301) <= a and not b;
    layer2_outputs(7302) <= not a;
    layer2_outputs(7303) <= not a;
    layer2_outputs(7304) <= not (a or b);
    layer2_outputs(7305) <= a and not b;
    layer2_outputs(7306) <= not (a xor b);
    layer2_outputs(7307) <= b and not a;
    layer2_outputs(7308) <= not (a xor b);
    layer2_outputs(7309) <= a or b;
    layer2_outputs(7310) <= b;
    layer2_outputs(7311) <= not a or b;
    layer2_outputs(7312) <= a and b;
    layer2_outputs(7313) <= not b;
    layer2_outputs(7314) <= b;
    layer2_outputs(7315) <= not a;
    layer2_outputs(7316) <= not (a or b);
    layer2_outputs(7317) <= a or b;
    layer2_outputs(7318) <= a xor b;
    layer2_outputs(7319) <= not a;
    layer2_outputs(7320) <= a and b;
    layer2_outputs(7321) <= not b;
    layer2_outputs(7322) <= not b;
    layer2_outputs(7323) <= a;
    layer2_outputs(7324) <= not (a xor b);
    layer2_outputs(7325) <= not a;
    layer2_outputs(7326) <= a;
    layer2_outputs(7327) <= not a;
    layer2_outputs(7328) <= a and b;
    layer2_outputs(7329) <= a;
    layer2_outputs(7330) <= not b;
    layer2_outputs(7331) <= not (a xor b);
    layer2_outputs(7332) <= not a or b;
    layer2_outputs(7333) <= a and not b;
    layer2_outputs(7334) <= a and not b;
    layer2_outputs(7335) <= not a or b;
    layer2_outputs(7336) <= b;
    layer2_outputs(7337) <= not (a and b);
    layer2_outputs(7338) <= not b or a;
    layer2_outputs(7339) <= not (a and b);
    layer2_outputs(7340) <= not (a xor b);
    layer2_outputs(7341) <= a and not b;
    layer2_outputs(7342) <= not a;
    layer2_outputs(7343) <= b;
    layer2_outputs(7344) <= not (a or b);
    layer2_outputs(7345) <= not (a or b);
    layer2_outputs(7346) <= a;
    layer2_outputs(7347) <= not (a or b);
    layer2_outputs(7348) <= not b;
    layer2_outputs(7349) <= b and not a;
    layer2_outputs(7350) <= not a;
    layer2_outputs(7351) <= not (a or b);
    layer2_outputs(7352) <= a and not b;
    layer2_outputs(7353) <= not (a xor b);
    layer2_outputs(7354) <= not a;
    layer2_outputs(7355) <= a and not b;
    layer2_outputs(7356) <= b and not a;
    layer2_outputs(7357) <= not a;
    layer2_outputs(7358) <= not (a and b);
    layer2_outputs(7359) <= a xor b;
    layer2_outputs(7360) <= not b;
    layer2_outputs(7361) <= a xor b;
    layer2_outputs(7362) <= a and not b;
    layer2_outputs(7363) <= not (a xor b);
    layer2_outputs(7364) <= not b;
    layer2_outputs(7365) <= a or b;
    layer2_outputs(7366) <= a and not b;
    layer2_outputs(7367) <= not a;
    layer2_outputs(7368) <= not a;
    layer2_outputs(7369) <= a xor b;
    layer2_outputs(7370) <= b and not a;
    layer2_outputs(7371) <= b;
    layer2_outputs(7372) <= 1'b1;
    layer2_outputs(7373) <= not (a or b);
    layer2_outputs(7374) <= not b;
    layer2_outputs(7375) <= b;
    layer2_outputs(7376) <= not (a or b);
    layer2_outputs(7377) <= a xor b;
    layer2_outputs(7378) <= not (a xor b);
    layer2_outputs(7379) <= a;
    layer2_outputs(7380) <= not (a xor b);
    layer2_outputs(7381) <= b and not a;
    layer2_outputs(7382) <= a and b;
    layer2_outputs(7383) <= not a;
    layer2_outputs(7384) <= not a;
    layer2_outputs(7385) <= a and b;
    layer2_outputs(7386) <= a and not b;
    layer2_outputs(7387) <= b;
    layer2_outputs(7388) <= not (a xor b);
    layer2_outputs(7389) <= a;
    layer2_outputs(7390) <= a xor b;
    layer2_outputs(7391) <= a and b;
    layer2_outputs(7392) <= not a;
    layer2_outputs(7393) <= b and not a;
    layer2_outputs(7394) <= not b or a;
    layer2_outputs(7395) <= a and not b;
    layer2_outputs(7396) <= a xor b;
    layer2_outputs(7397) <= not (a xor b);
    layer2_outputs(7398) <= not (a or b);
    layer2_outputs(7399) <= not a;
    layer2_outputs(7400) <= not a or b;
    layer2_outputs(7401) <= a xor b;
    layer2_outputs(7402) <= not b;
    layer2_outputs(7403) <= a or b;
    layer2_outputs(7404) <= a;
    layer2_outputs(7405) <= b;
    layer2_outputs(7406) <= not a;
    layer2_outputs(7407) <= a and not b;
    layer2_outputs(7408) <= not a;
    layer2_outputs(7409) <= b;
    layer2_outputs(7410) <= not (a and b);
    layer2_outputs(7411) <= a;
    layer2_outputs(7412) <= not (a xor b);
    layer2_outputs(7413) <= not a or b;
    layer2_outputs(7414) <= not (a xor b);
    layer2_outputs(7415) <= not a or b;
    layer2_outputs(7416) <= not a or b;
    layer2_outputs(7417) <= not b or a;
    layer2_outputs(7418) <= a xor b;
    layer2_outputs(7419) <= not b;
    layer2_outputs(7420) <= b;
    layer2_outputs(7421) <= not a;
    layer2_outputs(7422) <= a or b;
    layer2_outputs(7423) <= a and b;
    layer2_outputs(7424) <= not a;
    layer2_outputs(7425) <= a or b;
    layer2_outputs(7426) <= not b;
    layer2_outputs(7427) <= a and b;
    layer2_outputs(7428) <= a xor b;
    layer2_outputs(7429) <= b;
    layer2_outputs(7430) <= not (a or b);
    layer2_outputs(7431) <= b;
    layer2_outputs(7432) <= a and not b;
    layer2_outputs(7433) <= not (a or b);
    layer2_outputs(7434) <= not b;
    layer2_outputs(7435) <= a;
    layer2_outputs(7436) <= not a;
    layer2_outputs(7437) <= not (a and b);
    layer2_outputs(7438) <= a xor b;
    layer2_outputs(7439) <= a or b;
    layer2_outputs(7440) <= not (a xor b);
    layer2_outputs(7441) <= a;
    layer2_outputs(7442) <= not b;
    layer2_outputs(7443) <= not a;
    layer2_outputs(7444) <= b and not a;
    layer2_outputs(7445) <= b and not a;
    layer2_outputs(7446) <= not (a or b);
    layer2_outputs(7447) <= a;
    layer2_outputs(7448) <= not a or b;
    layer2_outputs(7449) <= not (a or b);
    layer2_outputs(7450) <= b;
    layer2_outputs(7451) <= not b;
    layer2_outputs(7452) <= a or b;
    layer2_outputs(7453) <= not a;
    layer2_outputs(7454) <= not b;
    layer2_outputs(7455) <= a xor b;
    layer2_outputs(7456) <= a;
    layer2_outputs(7457) <= not a;
    layer2_outputs(7458) <= a and not b;
    layer2_outputs(7459) <= a xor b;
    layer2_outputs(7460) <= a xor b;
    layer2_outputs(7461) <= b and not a;
    layer2_outputs(7462) <= b and not a;
    layer2_outputs(7463) <= b;
    layer2_outputs(7464) <= a and b;
    layer2_outputs(7465) <= not a;
    layer2_outputs(7466) <= a and b;
    layer2_outputs(7467) <= not (a and b);
    layer2_outputs(7468) <= a and b;
    layer2_outputs(7469) <= 1'b0;
    layer2_outputs(7470) <= not (a xor b);
    layer2_outputs(7471) <= not (a or b);
    layer2_outputs(7472) <= a and b;
    layer2_outputs(7473) <= 1'b0;
    layer2_outputs(7474) <= not (a and b);
    layer2_outputs(7475) <= a;
    layer2_outputs(7476) <= not (a or b);
    layer2_outputs(7477) <= a or b;
    layer2_outputs(7478) <= a and not b;
    layer2_outputs(7479) <= b;
    layer2_outputs(7480) <= a and b;
    layer2_outputs(7481) <= a or b;
    layer2_outputs(7482) <= not (a or b);
    layer2_outputs(7483) <= not (a xor b);
    layer2_outputs(7484) <= not a;
    layer2_outputs(7485) <= a;
    layer2_outputs(7486) <= not (a xor b);
    layer2_outputs(7487) <= b;
    layer2_outputs(7488) <= 1'b1;
    layer2_outputs(7489) <= not (a and b);
    layer2_outputs(7490) <= a;
    layer2_outputs(7491) <= b;
    layer2_outputs(7492) <= not b;
    layer2_outputs(7493) <= not (a or b);
    layer2_outputs(7494) <= b;
    layer2_outputs(7495) <= a and b;
    layer2_outputs(7496) <= not (a or b);
    layer2_outputs(7497) <= a xor b;
    layer2_outputs(7498) <= not a;
    layer2_outputs(7499) <= not b;
    layer2_outputs(7500) <= b;
    layer2_outputs(7501) <= a and not b;
    layer2_outputs(7502) <= a;
    layer2_outputs(7503) <= not b or a;
    layer2_outputs(7504) <= b;
    layer2_outputs(7505) <= not a;
    layer2_outputs(7506) <= a;
    layer2_outputs(7507) <= a xor b;
    layer2_outputs(7508) <= a;
    layer2_outputs(7509) <= not a;
    layer2_outputs(7510) <= b;
    layer2_outputs(7511) <= a;
    layer2_outputs(7512) <= a and not b;
    layer2_outputs(7513) <= not a or b;
    layer2_outputs(7514) <= a and not b;
    layer2_outputs(7515) <= a and b;
    layer2_outputs(7516) <= a xor b;
    layer2_outputs(7517) <= not (a xor b);
    layer2_outputs(7518) <= not a;
    layer2_outputs(7519) <= a and b;
    layer2_outputs(7520) <= b;
    layer2_outputs(7521) <= a and not b;
    layer2_outputs(7522) <= a or b;
    layer2_outputs(7523) <= a and not b;
    layer2_outputs(7524) <= not a;
    layer2_outputs(7525) <= not b;
    layer2_outputs(7526) <= not b or a;
    layer2_outputs(7527) <= not b or a;
    layer2_outputs(7528) <= not a;
    layer2_outputs(7529) <= a or b;
    layer2_outputs(7530) <= b and not a;
    layer2_outputs(7531) <= not a;
    layer2_outputs(7532) <= not b;
    layer2_outputs(7533) <= a and b;
    layer2_outputs(7534) <= a and not b;
    layer2_outputs(7535) <= a;
    layer2_outputs(7536) <= not (a xor b);
    layer2_outputs(7537) <= not (a xor b);
    layer2_outputs(7538) <= not b;
    layer2_outputs(7539) <= b and not a;
    layer2_outputs(7540) <= a or b;
    layer2_outputs(7541) <= a or b;
    layer2_outputs(7542) <= a;
    layer2_outputs(7543) <= a and not b;
    layer2_outputs(7544) <= not (a or b);
    layer2_outputs(7545) <= not (a or b);
    layer2_outputs(7546) <= not b;
    layer2_outputs(7547) <= a or b;
    layer2_outputs(7548) <= b;
    layer2_outputs(7549) <= not b or a;
    layer2_outputs(7550) <= b and not a;
    layer2_outputs(7551) <= 1'b0;
    layer2_outputs(7552) <= a and not b;
    layer2_outputs(7553) <= a;
    layer2_outputs(7554) <= a xor b;
    layer2_outputs(7555) <= b;
    layer2_outputs(7556) <= not (a xor b);
    layer2_outputs(7557) <= a;
    layer2_outputs(7558) <= not (a and b);
    layer2_outputs(7559) <= a or b;
    layer2_outputs(7560) <= a and b;
    layer2_outputs(7561) <= not a or b;
    layer2_outputs(7562) <= a or b;
    layer2_outputs(7563) <= a and not b;
    layer2_outputs(7564) <= a and b;
    layer2_outputs(7565) <= a;
    layer2_outputs(7566) <= not a or b;
    layer2_outputs(7567) <= a and not b;
    layer2_outputs(7568) <= a;
    layer2_outputs(7569) <= b;
    layer2_outputs(7570) <= b;
    layer2_outputs(7571) <= not a or b;
    layer2_outputs(7572) <= not (a and b);
    layer2_outputs(7573) <= not a or b;
    layer2_outputs(7574) <= not (a and b);
    layer2_outputs(7575) <= not (a xor b);
    layer2_outputs(7576) <= not b;
    layer2_outputs(7577) <= a xor b;
    layer2_outputs(7578) <= not (a xor b);
    layer2_outputs(7579) <= not (a or b);
    layer2_outputs(7580) <= a;
    layer2_outputs(7581) <= a;
    layer2_outputs(7582) <= not b;
    layer2_outputs(7583) <= not (a or b);
    layer2_outputs(7584) <= not b;
    layer2_outputs(7585) <= b and not a;
    layer2_outputs(7586) <= not a or b;
    layer2_outputs(7587) <= b and not a;
    layer2_outputs(7588) <= b and not a;
    layer2_outputs(7589) <= a and not b;
    layer2_outputs(7590) <= not (a xor b);
    layer2_outputs(7591) <= not (a xor b);
    layer2_outputs(7592) <= not (a and b);
    layer2_outputs(7593) <= not b or a;
    layer2_outputs(7594) <= not a;
    layer2_outputs(7595) <= a and not b;
    layer2_outputs(7596) <= not a;
    layer2_outputs(7597) <= not a;
    layer2_outputs(7598) <= b and not a;
    layer2_outputs(7599) <= a;
    layer2_outputs(7600) <= not (a xor b);
    layer2_outputs(7601) <= a;
    layer2_outputs(7602) <= a or b;
    layer2_outputs(7603) <= b;
    layer2_outputs(7604) <= not (a and b);
    layer2_outputs(7605) <= b and not a;
    layer2_outputs(7606) <= b;
    layer2_outputs(7607) <= not a;
    layer2_outputs(7608) <= a;
    layer2_outputs(7609) <= not a;
    layer2_outputs(7610) <= a or b;
    layer2_outputs(7611) <= a and not b;
    layer2_outputs(7612) <= not b;
    layer2_outputs(7613) <= a or b;
    layer2_outputs(7614) <= not (a and b);
    layer2_outputs(7615) <= not a;
    layer2_outputs(7616) <= a xor b;
    layer2_outputs(7617) <= 1'b1;
    layer2_outputs(7618) <= a;
    layer2_outputs(7619) <= not (a and b);
    layer2_outputs(7620) <= a xor b;
    layer2_outputs(7621) <= not b;
    layer2_outputs(7622) <= a;
    layer2_outputs(7623) <= a;
    layer2_outputs(7624) <= a xor b;
    layer2_outputs(7625) <= not b or a;
    layer2_outputs(7626) <= a;
    layer2_outputs(7627) <= not a or b;
    layer2_outputs(7628) <= a;
    layer2_outputs(7629) <= a or b;
    layer2_outputs(7630) <= a and b;
    layer2_outputs(7631) <= b and not a;
    layer2_outputs(7632) <= not a;
    layer2_outputs(7633) <= a;
    layer2_outputs(7634) <= a;
    layer2_outputs(7635) <= not (a and b);
    layer2_outputs(7636) <= a;
    layer2_outputs(7637) <= not a;
    layer2_outputs(7638) <= not (a or b);
    layer2_outputs(7639) <= a or b;
    layer2_outputs(7640) <= a and not b;
    layer2_outputs(7641) <= not a;
    layer2_outputs(7642) <= not a;
    layer2_outputs(7643) <= b and not a;
    layer2_outputs(7644) <= not (a xor b);
    layer2_outputs(7645) <= not a;
    layer2_outputs(7646) <= not b;
    layer2_outputs(7647) <= not (a or b);
    layer2_outputs(7648) <= a xor b;
    layer2_outputs(7649) <= not b;
    layer2_outputs(7650) <= not b;
    layer2_outputs(7651) <= not (a and b);
    layer2_outputs(7652) <= a xor b;
    layer2_outputs(7653) <= not a or b;
    layer2_outputs(7654) <= not (a xor b);
    layer2_outputs(7655) <= not (a xor b);
    layer2_outputs(7656) <= b;
    layer2_outputs(7657) <= not a;
    layer2_outputs(7658) <= not b;
    layer2_outputs(7659) <= not (a and b);
    layer2_outputs(7660) <= b and not a;
    layer2_outputs(7661) <= not b;
    layer2_outputs(7662) <= not (a xor b);
    layer2_outputs(7663) <= not (a xor b);
    layer2_outputs(7664) <= not b;
    layer2_outputs(7665) <= a and b;
    layer2_outputs(7666) <= b;
    layer2_outputs(7667) <= not (a or b);
    layer2_outputs(7668) <= not b;
    layer2_outputs(7669) <= not b or a;
    layer2_outputs(7670) <= not a;
    layer2_outputs(7671) <= not (a or b);
    layer2_outputs(7672) <= not a;
    layer2_outputs(7673) <= not (a and b);
    layer2_outputs(7674) <= a xor b;
    layer2_outputs(7675) <= b;
    layer2_outputs(7676) <= not (a or b);
    layer2_outputs(7677) <= b;
    layer2_outputs(7678) <= not a;
    layer2_outputs(7679) <= not (a xor b);
    layer2_outputs(7680) <= a or b;
    layer2_outputs(7681) <= not a;
    layer2_outputs(7682) <= a and b;
    layer2_outputs(7683) <= b;
    layer2_outputs(7684) <= not (a and b);
    layer2_outputs(7685) <= b;
    layer2_outputs(7686) <= not a;
    layer2_outputs(7687) <= not b;
    layer2_outputs(7688) <= a;
    layer2_outputs(7689) <= a and not b;
    layer2_outputs(7690) <= a or b;
    layer2_outputs(7691) <= a xor b;
    layer2_outputs(7692) <= a or b;
    layer2_outputs(7693) <= not a;
    layer2_outputs(7694) <= not (a xor b);
    layer2_outputs(7695) <= a or b;
    layer2_outputs(7696) <= not (a xor b);
    layer2_outputs(7697) <= a;
    layer2_outputs(7698) <= not b;
    layer2_outputs(7699) <= not (a xor b);
    layer2_outputs(7700) <= not a;
    layer2_outputs(7701) <= not a or b;
    layer2_outputs(7702) <= not (a xor b);
    layer2_outputs(7703) <= a xor b;
    layer2_outputs(7704) <= not a or b;
    layer2_outputs(7705) <= a;
    layer2_outputs(7706) <= a xor b;
    layer2_outputs(7707) <= a and not b;
    layer2_outputs(7708) <= b;
    layer2_outputs(7709) <= not (a xor b);
    layer2_outputs(7710) <= not a or b;
    layer2_outputs(7711) <= not a or b;
    layer2_outputs(7712) <= a xor b;
    layer2_outputs(7713) <= not a;
    layer2_outputs(7714) <= a or b;
    layer2_outputs(7715) <= a and not b;
    layer2_outputs(7716) <= not (a xor b);
    layer2_outputs(7717) <= not (a or b);
    layer2_outputs(7718) <= not a or b;
    layer2_outputs(7719) <= a;
    layer2_outputs(7720) <= not (a xor b);
    layer2_outputs(7721) <= 1'b0;
    layer2_outputs(7722) <= b;
    layer2_outputs(7723) <= a and b;
    layer2_outputs(7724) <= not b;
    layer2_outputs(7725) <= not b;
    layer2_outputs(7726) <= a and not b;
    layer2_outputs(7727) <= a xor b;
    layer2_outputs(7728) <= not b;
    layer2_outputs(7729) <= a;
    layer2_outputs(7730) <= not a;
    layer2_outputs(7731) <= b;
    layer2_outputs(7732) <= not (a or b);
    layer2_outputs(7733) <= not (a xor b);
    layer2_outputs(7734) <= not (a or b);
    layer2_outputs(7735) <= a;
    layer2_outputs(7736) <= a or b;
    layer2_outputs(7737) <= a xor b;
    layer2_outputs(7738) <= not b or a;
    layer2_outputs(7739) <= not (a and b);
    layer2_outputs(7740) <= not (a or b);
    layer2_outputs(7741) <= b and not a;
    layer2_outputs(7742) <= not b;
    layer2_outputs(7743) <= not (a and b);
    layer2_outputs(7744) <= a and not b;
    layer2_outputs(7745) <= not a or b;
    layer2_outputs(7746) <= not (a and b);
    layer2_outputs(7747) <= b;
    layer2_outputs(7748) <= a;
    layer2_outputs(7749) <= not b;
    layer2_outputs(7750) <= a xor b;
    layer2_outputs(7751) <= a;
    layer2_outputs(7752) <= not a or b;
    layer2_outputs(7753) <= a;
    layer2_outputs(7754) <= not a;
    layer2_outputs(7755) <= not (a xor b);
    layer2_outputs(7756) <= not b;
    layer2_outputs(7757) <= b;
    layer2_outputs(7758) <= not (a or b);
    layer2_outputs(7759) <= a or b;
    layer2_outputs(7760) <= a or b;
    layer2_outputs(7761) <= a;
    layer2_outputs(7762) <= not b or a;
    layer2_outputs(7763) <= a xor b;
    layer2_outputs(7764) <= a and not b;
    layer2_outputs(7765) <= a;
    layer2_outputs(7766) <= 1'b1;
    layer2_outputs(7767) <= b;
    layer2_outputs(7768) <= a;
    layer2_outputs(7769) <= not b or a;
    layer2_outputs(7770) <= not b or a;
    layer2_outputs(7771) <= not b;
    layer2_outputs(7772) <= not b;
    layer2_outputs(7773) <= a and b;
    layer2_outputs(7774) <= not b;
    layer2_outputs(7775) <= b;
    layer2_outputs(7776) <= not a;
    layer2_outputs(7777) <= b;
    layer2_outputs(7778) <= not (a xor b);
    layer2_outputs(7779) <= not (a xor b);
    layer2_outputs(7780) <= not (a or b);
    layer2_outputs(7781) <= not b;
    layer2_outputs(7782) <= not a;
    layer2_outputs(7783) <= not a;
    layer2_outputs(7784) <= not a or b;
    layer2_outputs(7785) <= b and not a;
    layer2_outputs(7786) <= not a;
    layer2_outputs(7787) <= a;
    layer2_outputs(7788) <= not (a and b);
    layer2_outputs(7789) <= not (a or b);
    layer2_outputs(7790) <= a or b;
    layer2_outputs(7791) <= not b;
    layer2_outputs(7792) <= a xor b;
    layer2_outputs(7793) <= not a or b;
    layer2_outputs(7794) <= not a or b;
    layer2_outputs(7795) <= not (a xor b);
    layer2_outputs(7796) <= not a;
    layer2_outputs(7797) <= a and not b;
    layer2_outputs(7798) <= not (a or b);
    layer2_outputs(7799) <= b and not a;
    layer2_outputs(7800) <= not (a or b);
    layer2_outputs(7801) <= b and not a;
    layer2_outputs(7802) <= a;
    layer2_outputs(7803) <= a;
    layer2_outputs(7804) <= a and not b;
    layer2_outputs(7805) <= a and b;
    layer2_outputs(7806) <= a and not b;
    layer2_outputs(7807) <= a;
    layer2_outputs(7808) <= a xor b;
    layer2_outputs(7809) <= not a or b;
    layer2_outputs(7810) <= a or b;
    layer2_outputs(7811) <= not (a or b);
    layer2_outputs(7812) <= not (a or b);
    layer2_outputs(7813) <= not a or b;
    layer2_outputs(7814) <= not b;
    layer2_outputs(7815) <= a and not b;
    layer2_outputs(7816) <= not b or a;
    layer2_outputs(7817) <= not (a and b);
    layer2_outputs(7818) <= b and not a;
    layer2_outputs(7819) <= not a;
    layer2_outputs(7820) <= a;
    layer2_outputs(7821) <= b and not a;
    layer2_outputs(7822) <= not b;
    layer2_outputs(7823) <= not (a xor b);
    layer2_outputs(7824) <= not (a or b);
    layer2_outputs(7825) <= not (a or b);
    layer2_outputs(7826) <= not b;
    layer2_outputs(7827) <= b and not a;
    layer2_outputs(7828) <= not b;
    layer2_outputs(7829) <= b;
    layer2_outputs(7830) <= not a;
    layer2_outputs(7831) <= not (a and b);
    layer2_outputs(7832) <= not a;
    layer2_outputs(7833) <= b and not a;
    layer2_outputs(7834) <= a xor b;
    layer2_outputs(7835) <= not b or a;
    layer2_outputs(7836) <= not b;
    layer2_outputs(7837) <= a or b;
    layer2_outputs(7838) <= b and not a;
    layer2_outputs(7839) <= not (a xor b);
    layer2_outputs(7840) <= not b;
    layer2_outputs(7841) <= a xor b;
    layer2_outputs(7842) <= a;
    layer2_outputs(7843) <= not b;
    layer2_outputs(7844) <= not (a xor b);
    layer2_outputs(7845) <= not (a and b);
    layer2_outputs(7846) <= a xor b;
    layer2_outputs(7847) <= not b;
    layer2_outputs(7848) <= not a;
    layer2_outputs(7849) <= a or b;
    layer2_outputs(7850) <= b;
    layer2_outputs(7851) <= not a;
    layer2_outputs(7852) <= not (a xor b);
    layer2_outputs(7853) <= not b or a;
    layer2_outputs(7854) <= not a;
    layer2_outputs(7855) <= a and b;
    layer2_outputs(7856) <= b;
    layer2_outputs(7857) <= not b or a;
    layer2_outputs(7858) <= not b or a;
    layer2_outputs(7859) <= not a;
    layer2_outputs(7860) <= not a or b;
    layer2_outputs(7861) <= not a;
    layer2_outputs(7862) <= not (a and b);
    layer2_outputs(7863) <= not (a xor b);
    layer2_outputs(7864) <= b and not a;
    layer2_outputs(7865) <= b;
    layer2_outputs(7866) <= b;
    layer2_outputs(7867) <= a xor b;
    layer2_outputs(7868) <= a and not b;
    layer2_outputs(7869) <= not (a xor b);
    layer2_outputs(7870) <= a xor b;
    layer2_outputs(7871) <= not a;
    layer2_outputs(7872) <= a or b;
    layer2_outputs(7873) <= a and not b;
    layer2_outputs(7874) <= a;
    layer2_outputs(7875) <= not b;
    layer2_outputs(7876) <= a;
    layer2_outputs(7877) <= not b or a;
    layer2_outputs(7878) <= not (a and b);
    layer2_outputs(7879) <= not a;
    layer2_outputs(7880) <= a xor b;
    layer2_outputs(7881) <= not b;
    layer2_outputs(7882) <= not (a xor b);
    layer2_outputs(7883) <= a;
    layer2_outputs(7884) <= not (a xor b);
    layer2_outputs(7885) <= a;
    layer2_outputs(7886) <= not b or a;
    layer2_outputs(7887) <= not (a xor b);
    layer2_outputs(7888) <= a or b;
    layer2_outputs(7889) <= not (a xor b);
    layer2_outputs(7890) <= not b or a;
    layer2_outputs(7891) <= a and b;
    layer2_outputs(7892) <= not a;
    layer2_outputs(7893) <= a;
    layer2_outputs(7894) <= a;
    layer2_outputs(7895) <= not (a and b);
    layer2_outputs(7896) <= a or b;
    layer2_outputs(7897) <= b and not a;
    layer2_outputs(7898) <= not b;
    layer2_outputs(7899) <= not a or b;
    layer2_outputs(7900) <= not b;
    layer2_outputs(7901) <= b;
    layer2_outputs(7902) <= not b;
    layer2_outputs(7903) <= not a;
    layer2_outputs(7904) <= a or b;
    layer2_outputs(7905) <= b;
    layer2_outputs(7906) <= not (a xor b);
    layer2_outputs(7907) <= not (a xor b);
    layer2_outputs(7908) <= not a;
    layer2_outputs(7909) <= not (a xor b);
    layer2_outputs(7910) <= b;
    layer2_outputs(7911) <= a xor b;
    layer2_outputs(7912) <= a and b;
    layer2_outputs(7913) <= a xor b;
    layer2_outputs(7914) <= a and b;
    layer2_outputs(7915) <= not a or b;
    layer2_outputs(7916) <= not a or b;
    layer2_outputs(7917) <= not a;
    layer2_outputs(7918) <= a xor b;
    layer2_outputs(7919) <= b and not a;
    layer2_outputs(7920) <= b;
    layer2_outputs(7921) <= not (a or b);
    layer2_outputs(7922) <= a or b;
    layer2_outputs(7923) <= a;
    layer2_outputs(7924) <= not (a or b);
    layer2_outputs(7925) <= not (a and b);
    layer2_outputs(7926) <= b;
    layer2_outputs(7927) <= a or b;
    layer2_outputs(7928) <= not (a and b);
    layer2_outputs(7929) <= not a;
    layer2_outputs(7930) <= a and b;
    layer2_outputs(7931) <= a xor b;
    layer2_outputs(7932) <= not a or b;
    layer2_outputs(7933) <= not a;
    layer2_outputs(7934) <= not (a xor b);
    layer2_outputs(7935) <= not (a xor b);
    layer2_outputs(7936) <= not (a xor b);
    layer2_outputs(7937) <= b;
    layer2_outputs(7938) <= b;
    layer2_outputs(7939) <= a and not b;
    layer2_outputs(7940) <= not b or a;
    layer2_outputs(7941) <= a or b;
    layer2_outputs(7942) <= not (a and b);
    layer2_outputs(7943) <= not a;
    layer2_outputs(7944) <= not (a xor b);
    layer2_outputs(7945) <= not a or b;
    layer2_outputs(7946) <= not a;
    layer2_outputs(7947) <= not (a xor b);
    layer2_outputs(7948) <= a xor b;
    layer2_outputs(7949) <= not (a and b);
    layer2_outputs(7950) <= not (a and b);
    layer2_outputs(7951) <= a xor b;
    layer2_outputs(7952) <= not b or a;
    layer2_outputs(7953) <= a xor b;
    layer2_outputs(7954) <= not b or a;
    layer2_outputs(7955) <= not a or b;
    layer2_outputs(7956) <= not (a or b);
    layer2_outputs(7957) <= a and not b;
    layer2_outputs(7958) <= b;
    layer2_outputs(7959) <= not b;
    layer2_outputs(7960) <= a or b;
    layer2_outputs(7961) <= not a;
    layer2_outputs(7962) <= not b or a;
    layer2_outputs(7963) <= b;
    layer2_outputs(7964) <= a xor b;
    layer2_outputs(7965) <= b and not a;
    layer2_outputs(7966) <= not b or a;
    layer2_outputs(7967) <= not (a or b);
    layer2_outputs(7968) <= a and b;
    layer2_outputs(7969) <= not (a or b);
    layer2_outputs(7970) <= a and b;
    layer2_outputs(7971) <= not (a or b);
    layer2_outputs(7972) <= not (a or b);
    layer2_outputs(7973) <= b and not a;
    layer2_outputs(7974) <= a and b;
    layer2_outputs(7975) <= a or b;
    layer2_outputs(7976) <= not b or a;
    layer2_outputs(7977) <= a and not b;
    layer2_outputs(7978) <= not b;
    layer2_outputs(7979) <= a;
    layer2_outputs(7980) <= a xor b;
    layer2_outputs(7981) <= not b;
    layer2_outputs(7982) <= not b or a;
    layer2_outputs(7983) <= b and not a;
    layer2_outputs(7984) <= a and not b;
    layer2_outputs(7985) <= a and b;
    layer2_outputs(7986) <= a and b;
    layer2_outputs(7987) <= not b;
    layer2_outputs(7988) <= not b;
    layer2_outputs(7989) <= not (a and b);
    layer2_outputs(7990) <= not b;
    layer2_outputs(7991) <= a;
    layer2_outputs(7992) <= not (a xor b);
    layer2_outputs(7993) <= a and not b;
    layer2_outputs(7994) <= a or b;
    layer2_outputs(7995) <= b;
    layer2_outputs(7996) <= a and b;
    layer2_outputs(7997) <= a xor b;
    layer2_outputs(7998) <= not (a or b);
    layer2_outputs(7999) <= not a;
    layer2_outputs(8000) <= not (a xor b);
    layer2_outputs(8001) <= b and not a;
    layer2_outputs(8002) <= a and b;
    layer2_outputs(8003) <= a;
    layer2_outputs(8004) <= not (a xor b);
    layer2_outputs(8005) <= a and not b;
    layer2_outputs(8006) <= a xor b;
    layer2_outputs(8007) <= a xor b;
    layer2_outputs(8008) <= b;
    layer2_outputs(8009) <= a or b;
    layer2_outputs(8010) <= b and not a;
    layer2_outputs(8011) <= not (a xor b);
    layer2_outputs(8012) <= a and not b;
    layer2_outputs(8013) <= b and not a;
    layer2_outputs(8014) <= not a;
    layer2_outputs(8015) <= b;
    layer2_outputs(8016) <= b;
    layer2_outputs(8017) <= not a;
    layer2_outputs(8018) <= b and not a;
    layer2_outputs(8019) <= not a or b;
    layer2_outputs(8020) <= b and not a;
    layer2_outputs(8021) <= not a;
    layer2_outputs(8022) <= not (a xor b);
    layer2_outputs(8023) <= b;
    layer2_outputs(8024) <= b;
    layer2_outputs(8025) <= not a;
    layer2_outputs(8026) <= a;
    layer2_outputs(8027) <= a or b;
    layer2_outputs(8028) <= a and not b;
    layer2_outputs(8029) <= b;
    layer2_outputs(8030) <= b;
    layer2_outputs(8031) <= a;
    layer2_outputs(8032) <= not (a xor b);
    layer2_outputs(8033) <= 1'b0;
    layer2_outputs(8034) <= a and not b;
    layer2_outputs(8035) <= a;
    layer2_outputs(8036) <= a and not b;
    layer2_outputs(8037) <= a;
    layer2_outputs(8038) <= not b;
    layer2_outputs(8039) <= b and not a;
    layer2_outputs(8040) <= a;
    layer2_outputs(8041) <= a xor b;
    layer2_outputs(8042) <= a xor b;
    layer2_outputs(8043) <= a and not b;
    layer2_outputs(8044) <= not b;
    layer2_outputs(8045) <= not (a xor b);
    layer2_outputs(8046) <= a xor b;
    layer2_outputs(8047) <= not a or b;
    layer2_outputs(8048) <= not (a or b);
    layer2_outputs(8049) <= a and b;
    layer2_outputs(8050) <= not b;
    layer2_outputs(8051) <= b;
    layer2_outputs(8052) <= a and b;
    layer2_outputs(8053) <= not a;
    layer2_outputs(8054) <= not a;
    layer2_outputs(8055) <= a;
    layer2_outputs(8056) <= not b or a;
    layer2_outputs(8057) <= b;
    layer2_outputs(8058) <= not (a xor b);
    layer2_outputs(8059) <= not a;
    layer2_outputs(8060) <= not b;
    layer2_outputs(8061) <= not a;
    layer2_outputs(8062) <= not (a xor b);
    layer2_outputs(8063) <= a and not b;
    layer2_outputs(8064) <= not b or a;
    layer2_outputs(8065) <= b and not a;
    layer2_outputs(8066) <= a xor b;
    layer2_outputs(8067) <= not (a or b);
    layer2_outputs(8068) <= not b or a;
    layer2_outputs(8069) <= b;
    layer2_outputs(8070) <= b;
    layer2_outputs(8071) <= a;
    layer2_outputs(8072) <= not b;
    layer2_outputs(8073) <= not a or b;
    layer2_outputs(8074) <= b;
    layer2_outputs(8075) <= not a;
    layer2_outputs(8076) <= not (a xor b);
    layer2_outputs(8077) <= a or b;
    layer2_outputs(8078) <= not b;
    layer2_outputs(8079) <= b and not a;
    layer2_outputs(8080) <= a xor b;
    layer2_outputs(8081) <= not (a and b);
    layer2_outputs(8082) <= not (a and b);
    layer2_outputs(8083) <= not a or b;
    layer2_outputs(8084) <= not a;
    layer2_outputs(8085) <= not a;
    layer2_outputs(8086) <= not (a xor b);
    layer2_outputs(8087) <= not a;
    layer2_outputs(8088) <= not b or a;
    layer2_outputs(8089) <= a or b;
    layer2_outputs(8090) <= b;
    layer2_outputs(8091) <= a and not b;
    layer2_outputs(8092) <= a;
    layer2_outputs(8093) <= b;
    layer2_outputs(8094) <= not (a or b);
    layer2_outputs(8095) <= not (a xor b);
    layer2_outputs(8096) <= a and not b;
    layer2_outputs(8097) <= a and b;
    layer2_outputs(8098) <= not (a xor b);
    layer2_outputs(8099) <= not (a or b);
    layer2_outputs(8100) <= not a;
    layer2_outputs(8101) <= not a;
    layer2_outputs(8102) <= a and not b;
    layer2_outputs(8103) <= not (a or b);
    layer2_outputs(8104) <= b;
    layer2_outputs(8105) <= not b;
    layer2_outputs(8106) <= a xor b;
    layer2_outputs(8107) <= not a;
    layer2_outputs(8108) <= b and not a;
    layer2_outputs(8109) <= 1'b0;
    layer2_outputs(8110) <= not b;
    layer2_outputs(8111) <= b and not a;
    layer2_outputs(8112) <= a xor b;
    layer2_outputs(8113) <= not b or a;
    layer2_outputs(8114) <= b;
    layer2_outputs(8115) <= not (a and b);
    layer2_outputs(8116) <= a and b;
    layer2_outputs(8117) <= not a or b;
    layer2_outputs(8118) <= not (a xor b);
    layer2_outputs(8119) <= a;
    layer2_outputs(8120) <= b;
    layer2_outputs(8121) <= not a;
    layer2_outputs(8122) <= b;
    layer2_outputs(8123) <= not (a or b);
    layer2_outputs(8124) <= a xor b;
    layer2_outputs(8125) <= not b;
    layer2_outputs(8126) <= a;
    layer2_outputs(8127) <= not a;
    layer2_outputs(8128) <= not b or a;
    layer2_outputs(8129) <= not (a and b);
    layer2_outputs(8130) <= not (a or b);
    layer2_outputs(8131) <= a xor b;
    layer2_outputs(8132) <= not (a xor b);
    layer2_outputs(8133) <= not a;
    layer2_outputs(8134) <= not (a and b);
    layer2_outputs(8135) <= b;
    layer2_outputs(8136) <= a and not b;
    layer2_outputs(8137) <= not a or b;
    layer2_outputs(8138) <= not (a or b);
    layer2_outputs(8139) <= a xor b;
    layer2_outputs(8140) <= not a;
    layer2_outputs(8141) <= a or b;
    layer2_outputs(8142) <= not b;
    layer2_outputs(8143) <= a and b;
    layer2_outputs(8144) <= a xor b;
    layer2_outputs(8145) <= a and not b;
    layer2_outputs(8146) <= not (a or b);
    layer2_outputs(8147) <= a and not b;
    layer2_outputs(8148) <= a and not b;
    layer2_outputs(8149) <= b;
    layer2_outputs(8150) <= a or b;
    layer2_outputs(8151) <= a xor b;
    layer2_outputs(8152) <= not b or a;
    layer2_outputs(8153) <= a xor b;
    layer2_outputs(8154) <= not (a xor b);
    layer2_outputs(8155) <= b;
    layer2_outputs(8156) <= not b;
    layer2_outputs(8157) <= not b or a;
    layer2_outputs(8158) <= b;
    layer2_outputs(8159) <= a;
    layer2_outputs(8160) <= a xor b;
    layer2_outputs(8161) <= a or b;
    layer2_outputs(8162) <= not b;
    layer2_outputs(8163) <= not a or b;
    layer2_outputs(8164) <= not b;
    layer2_outputs(8165) <= not a;
    layer2_outputs(8166) <= not a;
    layer2_outputs(8167) <= b and not a;
    layer2_outputs(8168) <= not (a or b);
    layer2_outputs(8169) <= not b or a;
    layer2_outputs(8170) <= a and b;
    layer2_outputs(8171) <= not b or a;
    layer2_outputs(8172) <= 1'b0;
    layer2_outputs(8173) <= not a;
    layer2_outputs(8174) <= a and not b;
    layer2_outputs(8175) <= not a;
    layer2_outputs(8176) <= a;
    layer2_outputs(8177) <= a xor b;
    layer2_outputs(8178) <= a;
    layer2_outputs(8179) <= a and not b;
    layer2_outputs(8180) <= not a or b;
    layer2_outputs(8181) <= not a;
    layer2_outputs(8182) <= not a;
    layer2_outputs(8183) <= not b;
    layer2_outputs(8184) <= a xor b;
    layer2_outputs(8185) <= not a;
    layer2_outputs(8186) <= not (a xor b);
    layer2_outputs(8187) <= a and not b;
    layer2_outputs(8188) <= not a;
    layer2_outputs(8189) <= a;
    layer2_outputs(8190) <= b;
    layer2_outputs(8191) <= b;
    layer2_outputs(8192) <= not (a and b);
    layer2_outputs(8193) <= a;
    layer2_outputs(8194) <= not b;
    layer2_outputs(8195) <= not a or b;
    layer2_outputs(8196) <= not b;
    layer2_outputs(8197) <= not (a xor b);
    layer2_outputs(8198) <= not a;
    layer2_outputs(8199) <= a xor b;
    layer2_outputs(8200) <= b;
    layer2_outputs(8201) <= a or b;
    layer2_outputs(8202) <= not a or b;
    layer2_outputs(8203) <= not b;
    layer2_outputs(8204) <= a xor b;
    layer2_outputs(8205) <= not b or a;
    layer2_outputs(8206) <= not b or a;
    layer2_outputs(8207) <= a;
    layer2_outputs(8208) <= not a;
    layer2_outputs(8209) <= a and b;
    layer2_outputs(8210) <= a xor b;
    layer2_outputs(8211) <= not b or a;
    layer2_outputs(8212) <= a xor b;
    layer2_outputs(8213) <= a xor b;
    layer2_outputs(8214) <= b;
    layer2_outputs(8215) <= not (a xor b);
    layer2_outputs(8216) <= a;
    layer2_outputs(8217) <= a;
    layer2_outputs(8218) <= 1'b0;
    layer2_outputs(8219) <= not (a xor b);
    layer2_outputs(8220) <= b;
    layer2_outputs(8221) <= a xor b;
    layer2_outputs(8222) <= b and not a;
    layer2_outputs(8223) <= not a;
    layer2_outputs(8224) <= not (a xor b);
    layer2_outputs(8225) <= not (a and b);
    layer2_outputs(8226) <= a;
    layer2_outputs(8227) <= not a or b;
    layer2_outputs(8228) <= not b or a;
    layer2_outputs(8229) <= not b or a;
    layer2_outputs(8230) <= b;
    layer2_outputs(8231) <= a and b;
    layer2_outputs(8232) <= not (a xor b);
    layer2_outputs(8233) <= a;
    layer2_outputs(8234) <= not b;
    layer2_outputs(8235) <= b;
    layer2_outputs(8236) <= b;
    layer2_outputs(8237) <= not (a xor b);
    layer2_outputs(8238) <= a and b;
    layer2_outputs(8239) <= not b or a;
    layer2_outputs(8240) <= 1'b1;
    layer2_outputs(8241) <= not (a xor b);
    layer2_outputs(8242) <= not (a xor b);
    layer2_outputs(8243) <= a xor b;
    layer2_outputs(8244) <= 1'b1;
    layer2_outputs(8245) <= not a;
    layer2_outputs(8246) <= not (a or b);
    layer2_outputs(8247) <= a xor b;
    layer2_outputs(8248) <= a;
    layer2_outputs(8249) <= not a;
    layer2_outputs(8250) <= a and b;
    layer2_outputs(8251) <= not a;
    layer2_outputs(8252) <= b;
    layer2_outputs(8253) <= a;
    layer2_outputs(8254) <= a;
    layer2_outputs(8255) <= a;
    layer2_outputs(8256) <= b and not a;
    layer2_outputs(8257) <= a xor b;
    layer2_outputs(8258) <= not b or a;
    layer2_outputs(8259) <= not b or a;
    layer2_outputs(8260) <= a and b;
    layer2_outputs(8261) <= not (a xor b);
    layer2_outputs(8262) <= not b or a;
    layer2_outputs(8263) <= b;
    layer2_outputs(8264) <= not (a or b);
    layer2_outputs(8265) <= not a;
    layer2_outputs(8266) <= not a;
    layer2_outputs(8267) <= a;
    layer2_outputs(8268) <= not (a or b);
    layer2_outputs(8269) <= b and not a;
    layer2_outputs(8270) <= not a;
    layer2_outputs(8271) <= not b or a;
    layer2_outputs(8272) <= not b or a;
    layer2_outputs(8273) <= a;
    layer2_outputs(8274) <= not a;
    layer2_outputs(8275) <= b and not a;
    layer2_outputs(8276) <= a and b;
    layer2_outputs(8277) <= a;
    layer2_outputs(8278) <= not (a xor b);
    layer2_outputs(8279) <= not (a and b);
    layer2_outputs(8280) <= not a or b;
    layer2_outputs(8281) <= not b;
    layer2_outputs(8282) <= a and b;
    layer2_outputs(8283) <= not b;
    layer2_outputs(8284) <= a and not b;
    layer2_outputs(8285) <= not b;
    layer2_outputs(8286) <= not b;
    layer2_outputs(8287) <= not a;
    layer2_outputs(8288) <= a xor b;
    layer2_outputs(8289) <= not (a and b);
    layer2_outputs(8290) <= a xor b;
    layer2_outputs(8291) <= not a or b;
    layer2_outputs(8292) <= not (a xor b);
    layer2_outputs(8293) <= not (a xor b);
    layer2_outputs(8294) <= not b or a;
    layer2_outputs(8295) <= b;
    layer2_outputs(8296) <= b;
    layer2_outputs(8297) <= not a or b;
    layer2_outputs(8298) <= not b or a;
    layer2_outputs(8299) <= b;
    layer2_outputs(8300) <= not (a and b);
    layer2_outputs(8301) <= not (a or b);
    layer2_outputs(8302) <= not a;
    layer2_outputs(8303) <= not (a xor b);
    layer2_outputs(8304) <= a xor b;
    layer2_outputs(8305) <= a or b;
    layer2_outputs(8306) <= a;
    layer2_outputs(8307) <= not b or a;
    layer2_outputs(8308) <= a;
    layer2_outputs(8309) <= b and not a;
    layer2_outputs(8310) <= a;
    layer2_outputs(8311) <= not (a xor b);
    layer2_outputs(8312) <= not (a xor b);
    layer2_outputs(8313) <= a xor b;
    layer2_outputs(8314) <= not (a or b);
    layer2_outputs(8315) <= a xor b;
    layer2_outputs(8316) <= not b;
    layer2_outputs(8317) <= a;
    layer2_outputs(8318) <= not (a and b);
    layer2_outputs(8319) <= not a;
    layer2_outputs(8320) <= a and not b;
    layer2_outputs(8321) <= b;
    layer2_outputs(8322) <= a;
    layer2_outputs(8323) <= a;
    layer2_outputs(8324) <= a and not b;
    layer2_outputs(8325) <= not a or b;
    layer2_outputs(8326) <= not (a xor b);
    layer2_outputs(8327) <= not b;
    layer2_outputs(8328) <= not a;
    layer2_outputs(8329) <= not b or a;
    layer2_outputs(8330) <= not (a xor b);
    layer2_outputs(8331) <= a xor b;
    layer2_outputs(8332) <= b;
    layer2_outputs(8333) <= not b or a;
    layer2_outputs(8334) <= not b or a;
    layer2_outputs(8335) <= b;
    layer2_outputs(8336) <= not (a xor b);
    layer2_outputs(8337) <= not (a and b);
    layer2_outputs(8338) <= not b or a;
    layer2_outputs(8339) <= not (a and b);
    layer2_outputs(8340) <= a or b;
    layer2_outputs(8341) <= not (a xor b);
    layer2_outputs(8342) <= b;
    layer2_outputs(8343) <= a and b;
    layer2_outputs(8344) <= not (a xor b);
    layer2_outputs(8345) <= a;
    layer2_outputs(8346) <= not a;
    layer2_outputs(8347) <= not a;
    layer2_outputs(8348) <= not b or a;
    layer2_outputs(8349) <= a and not b;
    layer2_outputs(8350) <= a xor b;
    layer2_outputs(8351) <= b and not a;
    layer2_outputs(8352) <= not b;
    layer2_outputs(8353) <= b and not a;
    layer2_outputs(8354) <= not a;
    layer2_outputs(8355) <= not (a xor b);
    layer2_outputs(8356) <= not b;
    layer2_outputs(8357) <= not b;
    layer2_outputs(8358) <= a xor b;
    layer2_outputs(8359) <= a;
    layer2_outputs(8360) <= not a;
    layer2_outputs(8361) <= 1'b1;
    layer2_outputs(8362) <= a xor b;
    layer2_outputs(8363) <= not b;
    layer2_outputs(8364) <= a and b;
    layer2_outputs(8365) <= a and b;
    layer2_outputs(8366) <= not b;
    layer2_outputs(8367) <= not b;
    layer2_outputs(8368) <= a and b;
    layer2_outputs(8369) <= b and not a;
    layer2_outputs(8370) <= not (a or b);
    layer2_outputs(8371) <= a;
    layer2_outputs(8372) <= a;
    layer2_outputs(8373) <= a or b;
    layer2_outputs(8374) <= a;
    layer2_outputs(8375) <= a or b;
    layer2_outputs(8376) <= not b;
    layer2_outputs(8377) <= not b or a;
    layer2_outputs(8378) <= not (a or b);
    layer2_outputs(8379) <= not (a or b);
    layer2_outputs(8380) <= a xor b;
    layer2_outputs(8381) <= b;
    layer2_outputs(8382) <= a;
    layer2_outputs(8383) <= not b;
    layer2_outputs(8384) <= a and not b;
    layer2_outputs(8385) <= a xor b;
    layer2_outputs(8386) <= not a;
    layer2_outputs(8387) <= a or b;
    layer2_outputs(8388) <= not (a and b);
    layer2_outputs(8389) <= not a;
    layer2_outputs(8390) <= not a;
    layer2_outputs(8391) <= a xor b;
    layer2_outputs(8392) <= not b;
    layer2_outputs(8393) <= not (a xor b);
    layer2_outputs(8394) <= not (a and b);
    layer2_outputs(8395) <= not (a and b);
    layer2_outputs(8396) <= not (a and b);
    layer2_outputs(8397) <= a xor b;
    layer2_outputs(8398) <= not (a and b);
    layer2_outputs(8399) <= b and not a;
    layer2_outputs(8400) <= a xor b;
    layer2_outputs(8401) <= not b;
    layer2_outputs(8402) <= a and b;
    layer2_outputs(8403) <= not a;
    layer2_outputs(8404) <= not a;
    layer2_outputs(8405) <= b;
    layer2_outputs(8406) <= not a;
    layer2_outputs(8407) <= not b or a;
    layer2_outputs(8408) <= a;
    layer2_outputs(8409) <= not b;
    layer2_outputs(8410) <= a and b;
    layer2_outputs(8411) <= not (a xor b);
    layer2_outputs(8412) <= a xor b;
    layer2_outputs(8413) <= a;
    layer2_outputs(8414) <= a or b;
    layer2_outputs(8415) <= a or b;
    layer2_outputs(8416) <= not b;
    layer2_outputs(8417) <= a or b;
    layer2_outputs(8418) <= not (a or b);
    layer2_outputs(8419) <= a and not b;
    layer2_outputs(8420) <= not b;
    layer2_outputs(8421) <= a and not b;
    layer2_outputs(8422) <= not (a xor b);
    layer2_outputs(8423) <= 1'b1;
    layer2_outputs(8424) <= not (a xor b);
    layer2_outputs(8425) <= b;
    layer2_outputs(8426) <= b;
    layer2_outputs(8427) <= a xor b;
    layer2_outputs(8428) <= not b;
    layer2_outputs(8429) <= a xor b;
    layer2_outputs(8430) <= b;
    layer2_outputs(8431) <= not (a and b);
    layer2_outputs(8432) <= not (a or b);
    layer2_outputs(8433) <= a;
    layer2_outputs(8434) <= b and not a;
    layer2_outputs(8435) <= not b;
    layer2_outputs(8436) <= not b or a;
    layer2_outputs(8437) <= a and b;
    layer2_outputs(8438) <= not (a or b);
    layer2_outputs(8439) <= not a or b;
    layer2_outputs(8440) <= a;
    layer2_outputs(8441) <= not a or b;
    layer2_outputs(8442) <= not (a xor b);
    layer2_outputs(8443) <= not (a and b);
    layer2_outputs(8444) <= not b or a;
    layer2_outputs(8445) <= not a;
    layer2_outputs(8446) <= not b;
    layer2_outputs(8447) <= not a;
    layer2_outputs(8448) <= a xor b;
    layer2_outputs(8449) <= a xor b;
    layer2_outputs(8450) <= not a;
    layer2_outputs(8451) <= a and not b;
    layer2_outputs(8452) <= b and not a;
    layer2_outputs(8453) <= not a or b;
    layer2_outputs(8454) <= a xor b;
    layer2_outputs(8455) <= a and b;
    layer2_outputs(8456) <= not a;
    layer2_outputs(8457) <= b;
    layer2_outputs(8458) <= not b;
    layer2_outputs(8459) <= not (a or b);
    layer2_outputs(8460) <= not (a xor b);
    layer2_outputs(8461) <= not b;
    layer2_outputs(8462) <= a and not b;
    layer2_outputs(8463) <= not (a xor b);
    layer2_outputs(8464) <= a xor b;
    layer2_outputs(8465) <= not b;
    layer2_outputs(8466) <= not b;
    layer2_outputs(8467) <= not a or b;
    layer2_outputs(8468) <= b and not a;
    layer2_outputs(8469) <= a or b;
    layer2_outputs(8470) <= not (a and b);
    layer2_outputs(8471) <= not a;
    layer2_outputs(8472) <= a and not b;
    layer2_outputs(8473) <= 1'b0;
    layer2_outputs(8474) <= not (a xor b);
    layer2_outputs(8475) <= a xor b;
    layer2_outputs(8476) <= a;
    layer2_outputs(8477) <= 1'b1;
    layer2_outputs(8478) <= a;
    layer2_outputs(8479) <= a or b;
    layer2_outputs(8480) <= not b;
    layer2_outputs(8481) <= a xor b;
    layer2_outputs(8482) <= a and b;
    layer2_outputs(8483) <= not b or a;
    layer2_outputs(8484) <= not a;
    layer2_outputs(8485) <= b and not a;
    layer2_outputs(8486) <= b;
    layer2_outputs(8487) <= a and b;
    layer2_outputs(8488) <= not b or a;
    layer2_outputs(8489) <= not b;
    layer2_outputs(8490) <= a and not b;
    layer2_outputs(8491) <= b;
    layer2_outputs(8492) <= not a;
    layer2_outputs(8493) <= not b;
    layer2_outputs(8494) <= not (a xor b);
    layer2_outputs(8495) <= not (a xor b);
    layer2_outputs(8496) <= a xor b;
    layer2_outputs(8497) <= a xor b;
    layer2_outputs(8498) <= a;
    layer2_outputs(8499) <= b;
    layer2_outputs(8500) <= a xor b;
    layer2_outputs(8501) <= a and b;
    layer2_outputs(8502) <= not (a and b);
    layer2_outputs(8503) <= b;
    layer2_outputs(8504) <= not (a or b);
    layer2_outputs(8505) <= a and b;
    layer2_outputs(8506) <= not (a or b);
    layer2_outputs(8507) <= a and not b;
    layer2_outputs(8508) <= a;
    layer2_outputs(8509) <= b;
    layer2_outputs(8510) <= not a;
    layer2_outputs(8511) <= b;
    layer2_outputs(8512) <= not (a xor b);
    layer2_outputs(8513) <= b and not a;
    layer2_outputs(8514) <= not a or b;
    layer2_outputs(8515) <= not (a xor b);
    layer2_outputs(8516) <= a;
    layer2_outputs(8517) <= not b;
    layer2_outputs(8518) <= not a;
    layer2_outputs(8519) <= a and not b;
    layer2_outputs(8520) <= not a;
    layer2_outputs(8521) <= a and not b;
    layer2_outputs(8522) <= not (a xor b);
    layer2_outputs(8523) <= not (a xor b);
    layer2_outputs(8524) <= a xor b;
    layer2_outputs(8525) <= a;
    layer2_outputs(8526) <= a or b;
    layer2_outputs(8527) <= not (a or b);
    layer2_outputs(8528) <= not b;
    layer2_outputs(8529) <= not (a and b);
    layer2_outputs(8530) <= not b or a;
    layer2_outputs(8531) <= a;
    layer2_outputs(8532) <= not (a or b);
    layer2_outputs(8533) <= not (a xor b);
    layer2_outputs(8534) <= not (a xor b);
    layer2_outputs(8535) <= a and not b;
    layer2_outputs(8536) <= b;
    layer2_outputs(8537) <= a or b;
    layer2_outputs(8538) <= not b or a;
    layer2_outputs(8539) <= b and not a;
    layer2_outputs(8540) <= a;
    layer2_outputs(8541) <= not a or b;
    layer2_outputs(8542) <= not (a xor b);
    layer2_outputs(8543) <= not a;
    layer2_outputs(8544) <= not b;
    layer2_outputs(8545) <= b;
    layer2_outputs(8546) <= not (a and b);
    layer2_outputs(8547) <= b and not a;
    layer2_outputs(8548) <= a or b;
    layer2_outputs(8549) <= not (a xor b);
    layer2_outputs(8550) <= not b;
    layer2_outputs(8551) <= not b or a;
    layer2_outputs(8552) <= b;
    layer2_outputs(8553) <= b;
    layer2_outputs(8554) <= b;
    layer2_outputs(8555) <= b;
    layer2_outputs(8556) <= b;
    layer2_outputs(8557) <= not a or b;
    layer2_outputs(8558) <= not a;
    layer2_outputs(8559) <= not b;
    layer2_outputs(8560) <= not b;
    layer2_outputs(8561) <= a or b;
    layer2_outputs(8562) <= a;
    layer2_outputs(8563) <= not b;
    layer2_outputs(8564) <= a xor b;
    layer2_outputs(8565) <= not (a xor b);
    layer2_outputs(8566) <= not a;
    layer2_outputs(8567) <= b;
    layer2_outputs(8568) <= not (a or b);
    layer2_outputs(8569) <= a and b;
    layer2_outputs(8570) <= a xor b;
    layer2_outputs(8571) <= not a;
    layer2_outputs(8572) <= a xor b;
    layer2_outputs(8573) <= b and not a;
    layer2_outputs(8574) <= b;
    layer2_outputs(8575) <= a;
    layer2_outputs(8576) <= not (a xor b);
    layer2_outputs(8577) <= not b;
    layer2_outputs(8578) <= a xor b;
    layer2_outputs(8579) <= b and not a;
    layer2_outputs(8580) <= a or b;
    layer2_outputs(8581) <= a and not b;
    layer2_outputs(8582) <= a and not b;
    layer2_outputs(8583) <= not b;
    layer2_outputs(8584) <= not b or a;
    layer2_outputs(8585) <= not b or a;
    layer2_outputs(8586) <= a and not b;
    layer2_outputs(8587) <= b and not a;
    layer2_outputs(8588) <= not (a xor b);
    layer2_outputs(8589) <= not (a xor b);
    layer2_outputs(8590) <= a and not b;
    layer2_outputs(8591) <= not b;
    layer2_outputs(8592) <= a xor b;
    layer2_outputs(8593) <= b;
    layer2_outputs(8594) <= not (a and b);
    layer2_outputs(8595) <= a and not b;
    layer2_outputs(8596) <= a and b;
    layer2_outputs(8597) <= not b;
    layer2_outputs(8598) <= a;
    layer2_outputs(8599) <= not (a and b);
    layer2_outputs(8600) <= a and not b;
    layer2_outputs(8601) <= not (a xor b);
    layer2_outputs(8602) <= not (a xor b);
    layer2_outputs(8603) <= not b or a;
    layer2_outputs(8604) <= not b;
    layer2_outputs(8605) <= b and not a;
    layer2_outputs(8606) <= a or b;
    layer2_outputs(8607) <= a xor b;
    layer2_outputs(8608) <= a;
    layer2_outputs(8609) <= not (a or b);
    layer2_outputs(8610) <= a;
    layer2_outputs(8611) <= b;
    layer2_outputs(8612) <= b and not a;
    layer2_outputs(8613) <= not b or a;
    layer2_outputs(8614) <= a xor b;
    layer2_outputs(8615) <= b and not a;
    layer2_outputs(8616) <= not a;
    layer2_outputs(8617) <= b;
    layer2_outputs(8618) <= not (a xor b);
    layer2_outputs(8619) <= a xor b;
    layer2_outputs(8620) <= b and not a;
    layer2_outputs(8621) <= a xor b;
    layer2_outputs(8622) <= a or b;
    layer2_outputs(8623) <= not b or a;
    layer2_outputs(8624) <= not (a and b);
    layer2_outputs(8625) <= a or b;
    layer2_outputs(8626) <= not (a xor b);
    layer2_outputs(8627) <= a or b;
    layer2_outputs(8628) <= not (a or b);
    layer2_outputs(8629) <= not (a xor b);
    layer2_outputs(8630) <= not b or a;
    layer2_outputs(8631) <= a;
    layer2_outputs(8632) <= not (a and b);
    layer2_outputs(8633) <= a xor b;
    layer2_outputs(8634) <= not b;
    layer2_outputs(8635) <= not a or b;
    layer2_outputs(8636) <= not (a xor b);
    layer2_outputs(8637) <= b;
    layer2_outputs(8638) <= not (a xor b);
    layer2_outputs(8639) <= a or b;
    layer2_outputs(8640) <= a and not b;
    layer2_outputs(8641) <= a xor b;
    layer2_outputs(8642) <= a and b;
    layer2_outputs(8643) <= not (a xor b);
    layer2_outputs(8644) <= a and b;
    layer2_outputs(8645) <= not b;
    layer2_outputs(8646) <= not (a xor b);
    layer2_outputs(8647) <= a xor b;
    layer2_outputs(8648) <= not (a xor b);
    layer2_outputs(8649) <= b and not a;
    layer2_outputs(8650) <= not a;
    layer2_outputs(8651) <= not a;
    layer2_outputs(8652) <= a;
    layer2_outputs(8653) <= not b;
    layer2_outputs(8654) <= a and not b;
    layer2_outputs(8655) <= not (a xor b);
    layer2_outputs(8656) <= not (a xor b);
    layer2_outputs(8657) <= not (a xor b);
    layer2_outputs(8658) <= a and not b;
    layer2_outputs(8659) <= b and not a;
    layer2_outputs(8660) <= b;
    layer2_outputs(8661) <= b and not a;
    layer2_outputs(8662) <= not a;
    layer2_outputs(8663) <= not (a xor b);
    layer2_outputs(8664) <= a xor b;
    layer2_outputs(8665) <= not b;
    layer2_outputs(8666) <= a xor b;
    layer2_outputs(8667) <= b;
    layer2_outputs(8668) <= not b;
    layer2_outputs(8669) <= not b;
    layer2_outputs(8670) <= not b;
    layer2_outputs(8671) <= b and not a;
    layer2_outputs(8672) <= not (a or b);
    layer2_outputs(8673) <= a;
    layer2_outputs(8674) <= b;
    layer2_outputs(8675) <= not (a or b);
    layer2_outputs(8676) <= a;
    layer2_outputs(8677) <= not b;
    layer2_outputs(8678) <= a or b;
    layer2_outputs(8679) <= a and not b;
    layer2_outputs(8680) <= b and not a;
    layer2_outputs(8681) <= b;
    layer2_outputs(8682) <= a or b;
    layer2_outputs(8683) <= a and not b;
    layer2_outputs(8684) <= b;
    layer2_outputs(8685) <= not b;
    layer2_outputs(8686) <= not b;
    layer2_outputs(8687) <= not (a xor b);
    layer2_outputs(8688) <= not a;
    layer2_outputs(8689) <= a;
    layer2_outputs(8690) <= b;
    layer2_outputs(8691) <= b;
    layer2_outputs(8692) <= a;
    layer2_outputs(8693) <= a xor b;
    layer2_outputs(8694) <= not b;
    layer2_outputs(8695) <= not (a and b);
    layer2_outputs(8696) <= a and not b;
    layer2_outputs(8697) <= b;
    layer2_outputs(8698) <= not (a or b);
    layer2_outputs(8699) <= not a;
    layer2_outputs(8700) <= not a or b;
    layer2_outputs(8701) <= a and not b;
    layer2_outputs(8702) <= not (a and b);
    layer2_outputs(8703) <= b;
    layer2_outputs(8704) <= a xor b;
    layer2_outputs(8705) <= not b;
    layer2_outputs(8706) <= a xor b;
    layer2_outputs(8707) <= not b;
    layer2_outputs(8708) <= b;
    layer2_outputs(8709) <= a and b;
    layer2_outputs(8710) <= b and not a;
    layer2_outputs(8711) <= not b;
    layer2_outputs(8712) <= b and not a;
    layer2_outputs(8713) <= not a;
    layer2_outputs(8714) <= a and b;
    layer2_outputs(8715) <= a or b;
    layer2_outputs(8716) <= not (a and b);
    layer2_outputs(8717) <= not a;
    layer2_outputs(8718) <= not (a or b);
    layer2_outputs(8719) <= not b or a;
    layer2_outputs(8720) <= a and b;
    layer2_outputs(8721) <= not b;
    layer2_outputs(8722) <= not (a xor b);
    layer2_outputs(8723) <= a or b;
    layer2_outputs(8724) <= not (a xor b);
    layer2_outputs(8725) <= not a or b;
    layer2_outputs(8726) <= a;
    layer2_outputs(8727) <= not b;
    layer2_outputs(8728) <= b;
    layer2_outputs(8729) <= a or b;
    layer2_outputs(8730) <= a or b;
    layer2_outputs(8731) <= not b;
    layer2_outputs(8732) <= a;
    layer2_outputs(8733) <= not b;
    layer2_outputs(8734) <= not a or b;
    layer2_outputs(8735) <= not b or a;
    layer2_outputs(8736) <= b;
    layer2_outputs(8737) <= not b or a;
    layer2_outputs(8738) <= a or b;
    layer2_outputs(8739) <= not b or a;
    layer2_outputs(8740) <= a and not b;
    layer2_outputs(8741) <= b;
    layer2_outputs(8742) <= a or b;
    layer2_outputs(8743) <= a;
    layer2_outputs(8744) <= a xor b;
    layer2_outputs(8745) <= a;
    layer2_outputs(8746) <= not a;
    layer2_outputs(8747) <= not (a or b);
    layer2_outputs(8748) <= b;
    layer2_outputs(8749) <= b;
    layer2_outputs(8750) <= not a;
    layer2_outputs(8751) <= not (a or b);
    layer2_outputs(8752) <= a;
    layer2_outputs(8753) <= not b;
    layer2_outputs(8754) <= b;
    layer2_outputs(8755) <= not a;
    layer2_outputs(8756) <= b;
    layer2_outputs(8757) <= a xor b;
    layer2_outputs(8758) <= a xor b;
    layer2_outputs(8759) <= not a;
    layer2_outputs(8760) <= not a;
    layer2_outputs(8761) <= not a;
    layer2_outputs(8762) <= not b or a;
    layer2_outputs(8763) <= a or b;
    layer2_outputs(8764) <= not b or a;
    layer2_outputs(8765) <= b;
    layer2_outputs(8766) <= a or b;
    layer2_outputs(8767) <= b;
    layer2_outputs(8768) <= a xor b;
    layer2_outputs(8769) <= not (a and b);
    layer2_outputs(8770) <= not a;
    layer2_outputs(8771) <= not (a and b);
    layer2_outputs(8772) <= a;
    layer2_outputs(8773) <= not (a xor b);
    layer2_outputs(8774) <= b and not a;
    layer2_outputs(8775) <= not (a xor b);
    layer2_outputs(8776) <= a;
    layer2_outputs(8777) <= a;
    layer2_outputs(8778) <= not b;
    layer2_outputs(8779) <= not b or a;
    layer2_outputs(8780) <= a;
    layer2_outputs(8781) <= a;
    layer2_outputs(8782) <= not a or b;
    layer2_outputs(8783) <= not b;
    layer2_outputs(8784) <= a or b;
    layer2_outputs(8785) <= a and not b;
    layer2_outputs(8786) <= not (a or b);
    layer2_outputs(8787) <= b and not a;
    layer2_outputs(8788) <= a and b;
    layer2_outputs(8789) <= a;
    layer2_outputs(8790) <= not b or a;
    layer2_outputs(8791) <= not a;
    layer2_outputs(8792) <= not b;
    layer2_outputs(8793) <= b;
    layer2_outputs(8794) <= not (a or b);
    layer2_outputs(8795) <= b and not a;
    layer2_outputs(8796) <= not b;
    layer2_outputs(8797) <= a;
    layer2_outputs(8798) <= b;
    layer2_outputs(8799) <= b;
    layer2_outputs(8800) <= not b;
    layer2_outputs(8801) <= not b or a;
    layer2_outputs(8802) <= a and not b;
    layer2_outputs(8803) <= not a;
    layer2_outputs(8804) <= not (a or b);
    layer2_outputs(8805) <= a xor b;
    layer2_outputs(8806) <= not a or b;
    layer2_outputs(8807) <= a or b;
    layer2_outputs(8808) <= not (a xor b);
    layer2_outputs(8809) <= not (a and b);
    layer2_outputs(8810) <= b;
    layer2_outputs(8811) <= not (a or b);
    layer2_outputs(8812) <= b;
    layer2_outputs(8813) <= not a or b;
    layer2_outputs(8814) <= a and not b;
    layer2_outputs(8815) <= not b;
    layer2_outputs(8816) <= a and not b;
    layer2_outputs(8817) <= not (a or b);
    layer2_outputs(8818) <= a and b;
    layer2_outputs(8819) <= not a;
    layer2_outputs(8820) <= not (a xor b);
    layer2_outputs(8821) <= not b or a;
    layer2_outputs(8822) <= b;
    layer2_outputs(8823) <= a or b;
    layer2_outputs(8824) <= not a or b;
    layer2_outputs(8825) <= not a;
    layer2_outputs(8826) <= a xor b;
    layer2_outputs(8827) <= not b or a;
    layer2_outputs(8828) <= not (a and b);
    layer2_outputs(8829) <= not b or a;
    layer2_outputs(8830) <= a;
    layer2_outputs(8831) <= a and b;
    layer2_outputs(8832) <= a and b;
    layer2_outputs(8833) <= 1'b0;
    layer2_outputs(8834) <= not b or a;
    layer2_outputs(8835) <= b;
    layer2_outputs(8836) <= a or b;
    layer2_outputs(8837) <= b;
    layer2_outputs(8838) <= not (a and b);
    layer2_outputs(8839) <= a;
    layer2_outputs(8840) <= not a;
    layer2_outputs(8841) <= a xor b;
    layer2_outputs(8842) <= not (a and b);
    layer2_outputs(8843) <= not a or b;
    layer2_outputs(8844) <= not (a and b);
    layer2_outputs(8845) <= not (a or b);
    layer2_outputs(8846) <= a xor b;
    layer2_outputs(8847) <= b and not a;
    layer2_outputs(8848) <= not (a xor b);
    layer2_outputs(8849) <= not a;
    layer2_outputs(8850) <= a xor b;
    layer2_outputs(8851) <= b and not a;
    layer2_outputs(8852) <= not (a and b);
    layer2_outputs(8853) <= a and not b;
    layer2_outputs(8854) <= b and not a;
    layer2_outputs(8855) <= 1'b1;
    layer2_outputs(8856) <= a and b;
    layer2_outputs(8857) <= not b;
    layer2_outputs(8858) <= not a;
    layer2_outputs(8859) <= not a;
    layer2_outputs(8860) <= not (a and b);
    layer2_outputs(8861) <= b;
    layer2_outputs(8862) <= not a or b;
    layer2_outputs(8863) <= not b;
    layer2_outputs(8864) <= a xor b;
    layer2_outputs(8865) <= not (a xor b);
    layer2_outputs(8866) <= not b;
    layer2_outputs(8867) <= not a;
    layer2_outputs(8868) <= not (a xor b);
    layer2_outputs(8869) <= not (a xor b);
    layer2_outputs(8870) <= a and b;
    layer2_outputs(8871) <= b;
    layer2_outputs(8872) <= a;
    layer2_outputs(8873) <= not a or b;
    layer2_outputs(8874) <= not (a xor b);
    layer2_outputs(8875) <= b;
    layer2_outputs(8876) <= not b;
    layer2_outputs(8877) <= not b;
    layer2_outputs(8878) <= b;
    layer2_outputs(8879) <= not a or b;
    layer2_outputs(8880) <= not (a and b);
    layer2_outputs(8881) <= not (a and b);
    layer2_outputs(8882) <= not (a or b);
    layer2_outputs(8883) <= b;
    layer2_outputs(8884) <= not (a xor b);
    layer2_outputs(8885) <= not a or b;
    layer2_outputs(8886) <= a xor b;
    layer2_outputs(8887) <= a xor b;
    layer2_outputs(8888) <= b and not a;
    layer2_outputs(8889) <= not (a and b);
    layer2_outputs(8890) <= a;
    layer2_outputs(8891) <= not (a or b);
    layer2_outputs(8892) <= a;
    layer2_outputs(8893) <= b;
    layer2_outputs(8894) <= a xor b;
    layer2_outputs(8895) <= not (a and b);
    layer2_outputs(8896) <= not b;
    layer2_outputs(8897) <= not a;
    layer2_outputs(8898) <= not b;
    layer2_outputs(8899) <= b;
    layer2_outputs(8900) <= a;
    layer2_outputs(8901) <= a and not b;
    layer2_outputs(8902) <= a;
    layer2_outputs(8903) <= b;
    layer2_outputs(8904) <= a or b;
    layer2_outputs(8905) <= a;
    layer2_outputs(8906) <= not (a or b);
    layer2_outputs(8907) <= not (a xor b);
    layer2_outputs(8908) <= not (a or b);
    layer2_outputs(8909) <= 1'b1;
    layer2_outputs(8910) <= a xor b;
    layer2_outputs(8911) <= a;
    layer2_outputs(8912) <= b;
    layer2_outputs(8913) <= a;
    layer2_outputs(8914) <= b;
    layer2_outputs(8915) <= not (a xor b);
    layer2_outputs(8916) <= a and b;
    layer2_outputs(8917) <= b and not a;
    layer2_outputs(8918) <= not b;
    layer2_outputs(8919) <= a;
    layer2_outputs(8920) <= a;
    layer2_outputs(8921) <= not a or b;
    layer2_outputs(8922) <= not (a or b);
    layer2_outputs(8923) <= a and not b;
    layer2_outputs(8924) <= not b;
    layer2_outputs(8925) <= a xor b;
    layer2_outputs(8926) <= not (a and b);
    layer2_outputs(8927) <= not a or b;
    layer2_outputs(8928) <= not (a or b);
    layer2_outputs(8929) <= a xor b;
    layer2_outputs(8930) <= not a;
    layer2_outputs(8931) <= not b;
    layer2_outputs(8932) <= b and not a;
    layer2_outputs(8933) <= not b;
    layer2_outputs(8934) <= a or b;
    layer2_outputs(8935) <= not a;
    layer2_outputs(8936) <= not (a xor b);
    layer2_outputs(8937) <= a and not b;
    layer2_outputs(8938) <= not (a xor b);
    layer2_outputs(8939) <= not b;
    layer2_outputs(8940) <= a;
    layer2_outputs(8941) <= not b;
    layer2_outputs(8942) <= a;
    layer2_outputs(8943) <= not b or a;
    layer2_outputs(8944) <= not (a or b);
    layer2_outputs(8945) <= not a or b;
    layer2_outputs(8946) <= not b or a;
    layer2_outputs(8947) <= not (a and b);
    layer2_outputs(8948) <= a or b;
    layer2_outputs(8949) <= b and not a;
    layer2_outputs(8950) <= not (a and b);
    layer2_outputs(8951) <= not a or b;
    layer2_outputs(8952) <= not (a xor b);
    layer2_outputs(8953) <= b;
    layer2_outputs(8954) <= a xor b;
    layer2_outputs(8955) <= not b or a;
    layer2_outputs(8956) <= a and b;
    layer2_outputs(8957) <= not a;
    layer2_outputs(8958) <= a;
    layer2_outputs(8959) <= not (a and b);
    layer2_outputs(8960) <= not b or a;
    layer2_outputs(8961) <= not (a xor b);
    layer2_outputs(8962) <= not (a or b);
    layer2_outputs(8963) <= not a;
    layer2_outputs(8964) <= not b;
    layer2_outputs(8965) <= not (a xor b);
    layer2_outputs(8966) <= b;
    layer2_outputs(8967) <= not (a xor b);
    layer2_outputs(8968) <= not (a xor b);
    layer2_outputs(8969) <= not a;
    layer2_outputs(8970) <= not (a xor b);
    layer2_outputs(8971) <= b;
    layer2_outputs(8972) <= not b;
    layer2_outputs(8973) <= b;
    layer2_outputs(8974) <= not (a and b);
    layer2_outputs(8975) <= not a;
    layer2_outputs(8976) <= a;
    layer2_outputs(8977) <= not (a xor b);
    layer2_outputs(8978) <= not (a or b);
    layer2_outputs(8979) <= not a;
    layer2_outputs(8980) <= a and b;
    layer2_outputs(8981) <= not a or b;
    layer2_outputs(8982) <= not a;
    layer2_outputs(8983) <= b;
    layer2_outputs(8984) <= not b or a;
    layer2_outputs(8985) <= not (a and b);
    layer2_outputs(8986) <= b;
    layer2_outputs(8987) <= a;
    layer2_outputs(8988) <= not a;
    layer2_outputs(8989) <= not b or a;
    layer2_outputs(8990) <= a xor b;
    layer2_outputs(8991) <= b;
    layer2_outputs(8992) <= not (a and b);
    layer2_outputs(8993) <= a and not b;
    layer2_outputs(8994) <= a xor b;
    layer2_outputs(8995) <= a;
    layer2_outputs(8996) <= a or b;
    layer2_outputs(8997) <= a or b;
    layer2_outputs(8998) <= not a;
    layer2_outputs(8999) <= not b or a;
    layer2_outputs(9000) <= not (a xor b);
    layer2_outputs(9001) <= a xor b;
    layer2_outputs(9002) <= a and not b;
    layer2_outputs(9003) <= not (a xor b);
    layer2_outputs(9004) <= b and not a;
    layer2_outputs(9005) <= b;
    layer2_outputs(9006) <= a;
    layer2_outputs(9007) <= a xor b;
    layer2_outputs(9008) <= b;
    layer2_outputs(9009) <= not b;
    layer2_outputs(9010) <= a and b;
    layer2_outputs(9011) <= a;
    layer2_outputs(9012) <= not (a or b);
    layer2_outputs(9013) <= b;
    layer2_outputs(9014) <= a;
    layer2_outputs(9015) <= a;
    layer2_outputs(9016) <= a;
    layer2_outputs(9017) <= not (a xor b);
    layer2_outputs(9018) <= a or b;
    layer2_outputs(9019) <= not (a xor b);
    layer2_outputs(9020) <= not a or b;
    layer2_outputs(9021) <= a xor b;
    layer2_outputs(9022) <= not b;
    layer2_outputs(9023) <= b and not a;
    layer2_outputs(9024) <= b;
    layer2_outputs(9025) <= b;
    layer2_outputs(9026) <= not a;
    layer2_outputs(9027) <= a xor b;
    layer2_outputs(9028) <= a;
    layer2_outputs(9029) <= not (a xor b);
    layer2_outputs(9030) <= a;
    layer2_outputs(9031) <= not (a xor b);
    layer2_outputs(9032) <= not a;
    layer2_outputs(9033) <= b;
    layer2_outputs(9034) <= a xor b;
    layer2_outputs(9035) <= a xor b;
    layer2_outputs(9036) <= b and not a;
    layer2_outputs(9037) <= not (a xor b);
    layer2_outputs(9038) <= a;
    layer2_outputs(9039) <= a or b;
    layer2_outputs(9040) <= a xor b;
    layer2_outputs(9041) <= b;
    layer2_outputs(9042) <= not a or b;
    layer2_outputs(9043) <= not b or a;
    layer2_outputs(9044) <= b;
    layer2_outputs(9045) <= not (a xor b);
    layer2_outputs(9046) <= a and not b;
    layer2_outputs(9047) <= a and not b;
    layer2_outputs(9048) <= b;
    layer2_outputs(9049) <= not (a or b);
    layer2_outputs(9050) <= not b;
    layer2_outputs(9051) <= a xor b;
    layer2_outputs(9052) <= not a or b;
    layer2_outputs(9053) <= not (a and b);
    layer2_outputs(9054) <= not (a xor b);
    layer2_outputs(9055) <= a;
    layer2_outputs(9056) <= a and not b;
    layer2_outputs(9057) <= a and not b;
    layer2_outputs(9058) <= a or b;
    layer2_outputs(9059) <= a xor b;
    layer2_outputs(9060) <= not (a or b);
    layer2_outputs(9061) <= a and b;
    layer2_outputs(9062) <= not a or b;
    layer2_outputs(9063) <= not (a or b);
    layer2_outputs(9064) <= not (a xor b);
    layer2_outputs(9065) <= not (a xor b);
    layer2_outputs(9066) <= a;
    layer2_outputs(9067) <= a;
    layer2_outputs(9068) <= not b;
    layer2_outputs(9069) <= a and not b;
    layer2_outputs(9070) <= not (a and b);
    layer2_outputs(9071) <= b;
    layer2_outputs(9072) <= a;
    layer2_outputs(9073) <= not (a or b);
    layer2_outputs(9074) <= b;
    layer2_outputs(9075) <= not (a xor b);
    layer2_outputs(9076) <= not b;
    layer2_outputs(9077) <= not (a or b);
    layer2_outputs(9078) <= not (a xor b);
    layer2_outputs(9079) <= a;
    layer2_outputs(9080) <= b and not a;
    layer2_outputs(9081) <= a;
    layer2_outputs(9082) <= b and not a;
    layer2_outputs(9083) <= b;
    layer2_outputs(9084) <= a and b;
    layer2_outputs(9085) <= not (a and b);
    layer2_outputs(9086) <= not a or b;
    layer2_outputs(9087) <= a xor b;
    layer2_outputs(9088) <= a or b;
    layer2_outputs(9089) <= not b or a;
    layer2_outputs(9090) <= a and not b;
    layer2_outputs(9091) <= a and b;
    layer2_outputs(9092) <= not a or b;
    layer2_outputs(9093) <= a and b;
    layer2_outputs(9094) <= a xor b;
    layer2_outputs(9095) <= not b;
    layer2_outputs(9096) <= not (a xor b);
    layer2_outputs(9097) <= not (a xor b);
    layer2_outputs(9098) <= not a or b;
    layer2_outputs(9099) <= a and b;
    layer2_outputs(9100) <= not (a xor b);
    layer2_outputs(9101) <= not b;
    layer2_outputs(9102) <= not a or b;
    layer2_outputs(9103) <= a;
    layer2_outputs(9104) <= a;
    layer2_outputs(9105) <= not b;
    layer2_outputs(9106) <= not a;
    layer2_outputs(9107) <= b;
    layer2_outputs(9108) <= a;
    layer2_outputs(9109) <= a xor b;
    layer2_outputs(9110) <= not a or b;
    layer2_outputs(9111) <= not (a xor b);
    layer2_outputs(9112) <= not a or b;
    layer2_outputs(9113) <= not (a xor b);
    layer2_outputs(9114) <= b;
    layer2_outputs(9115) <= a xor b;
    layer2_outputs(9116) <= b and not a;
    layer2_outputs(9117) <= not (a xor b);
    layer2_outputs(9118) <= not (a xor b);
    layer2_outputs(9119) <= not a;
    layer2_outputs(9120) <= a;
    layer2_outputs(9121) <= a xor b;
    layer2_outputs(9122) <= not b;
    layer2_outputs(9123) <= b and not a;
    layer2_outputs(9124) <= not a;
    layer2_outputs(9125) <= not a;
    layer2_outputs(9126) <= b;
    layer2_outputs(9127) <= not (a or b);
    layer2_outputs(9128) <= b;
    layer2_outputs(9129) <= not (a xor b);
    layer2_outputs(9130) <= a and b;
    layer2_outputs(9131) <= not b or a;
    layer2_outputs(9132) <= not b or a;
    layer2_outputs(9133) <= not (a and b);
    layer2_outputs(9134) <= not a or b;
    layer2_outputs(9135) <= b;
    layer2_outputs(9136) <= not a;
    layer2_outputs(9137) <= not b;
    layer2_outputs(9138) <= not a;
    layer2_outputs(9139) <= a and b;
    layer2_outputs(9140) <= not b;
    layer2_outputs(9141) <= not b;
    layer2_outputs(9142) <= a;
    layer2_outputs(9143) <= not (a or b);
    layer2_outputs(9144) <= b and not a;
    layer2_outputs(9145) <= a;
    layer2_outputs(9146) <= not (a xor b);
    layer2_outputs(9147) <= b;
    layer2_outputs(9148) <= b and not a;
    layer2_outputs(9149) <= not a;
    layer2_outputs(9150) <= b and not a;
    layer2_outputs(9151) <= not b or a;
    layer2_outputs(9152) <= not b;
    layer2_outputs(9153) <= b;
    layer2_outputs(9154) <= not (a or b);
    layer2_outputs(9155) <= not b;
    layer2_outputs(9156) <= not a;
    layer2_outputs(9157) <= b and not a;
    layer2_outputs(9158) <= not (a and b);
    layer2_outputs(9159) <= not (a and b);
    layer2_outputs(9160) <= a;
    layer2_outputs(9161) <= not (a or b);
    layer2_outputs(9162) <= not (a and b);
    layer2_outputs(9163) <= b;
    layer2_outputs(9164) <= a;
    layer2_outputs(9165) <= not (a xor b);
    layer2_outputs(9166) <= not a;
    layer2_outputs(9167) <= a;
    layer2_outputs(9168) <= not (a xor b);
    layer2_outputs(9169) <= not (a and b);
    layer2_outputs(9170) <= a xor b;
    layer2_outputs(9171) <= a and not b;
    layer2_outputs(9172) <= not a or b;
    layer2_outputs(9173) <= b and not a;
    layer2_outputs(9174) <= b;
    layer2_outputs(9175) <= not a or b;
    layer2_outputs(9176) <= a xor b;
    layer2_outputs(9177) <= not b;
    layer2_outputs(9178) <= a or b;
    layer2_outputs(9179) <= not a;
    layer2_outputs(9180) <= not b;
    layer2_outputs(9181) <= a xor b;
    layer2_outputs(9182) <= not (a or b);
    layer2_outputs(9183) <= not b or a;
    layer2_outputs(9184) <= a and b;
    layer2_outputs(9185) <= b;
    layer2_outputs(9186) <= a xor b;
    layer2_outputs(9187) <= a;
    layer2_outputs(9188) <= a or b;
    layer2_outputs(9189) <= a;
    layer2_outputs(9190) <= not (a xor b);
    layer2_outputs(9191) <= not (a xor b);
    layer2_outputs(9192) <= not b;
    layer2_outputs(9193) <= a and not b;
    layer2_outputs(9194) <= b and not a;
    layer2_outputs(9195) <= a xor b;
    layer2_outputs(9196) <= not (a xor b);
    layer2_outputs(9197) <= b;
    layer2_outputs(9198) <= a xor b;
    layer2_outputs(9199) <= a and b;
    layer2_outputs(9200) <= a xor b;
    layer2_outputs(9201) <= a xor b;
    layer2_outputs(9202) <= b and not a;
    layer2_outputs(9203) <= not b;
    layer2_outputs(9204) <= b and not a;
    layer2_outputs(9205) <= a or b;
    layer2_outputs(9206) <= not a or b;
    layer2_outputs(9207) <= not (a xor b);
    layer2_outputs(9208) <= a;
    layer2_outputs(9209) <= a xor b;
    layer2_outputs(9210) <= not a or b;
    layer2_outputs(9211) <= b and not a;
    layer2_outputs(9212) <= not a;
    layer2_outputs(9213) <= a or b;
    layer2_outputs(9214) <= b;
    layer2_outputs(9215) <= not (a or b);
    layer2_outputs(9216) <= a xor b;
    layer2_outputs(9217) <= a xor b;
    layer2_outputs(9218) <= a xor b;
    layer2_outputs(9219) <= not b;
    layer2_outputs(9220) <= not a;
    layer2_outputs(9221) <= a;
    layer2_outputs(9222) <= not a;
    layer2_outputs(9223) <= not a or b;
    layer2_outputs(9224) <= not a;
    layer2_outputs(9225) <= b and not a;
    layer2_outputs(9226) <= a;
    layer2_outputs(9227) <= not a;
    layer2_outputs(9228) <= not b or a;
    layer2_outputs(9229) <= a;
    layer2_outputs(9230) <= not b;
    layer2_outputs(9231) <= a and b;
    layer2_outputs(9232) <= not b;
    layer2_outputs(9233) <= b;
    layer2_outputs(9234) <= not b or a;
    layer2_outputs(9235) <= a;
    layer2_outputs(9236) <= not a;
    layer2_outputs(9237) <= not b;
    layer2_outputs(9238) <= not a;
    layer2_outputs(9239) <= not a;
    layer2_outputs(9240) <= a or b;
    layer2_outputs(9241) <= a xor b;
    layer2_outputs(9242) <= a or b;
    layer2_outputs(9243) <= not b;
    layer2_outputs(9244) <= not a;
    layer2_outputs(9245) <= not (a xor b);
    layer2_outputs(9246) <= not b or a;
    layer2_outputs(9247) <= a;
    layer2_outputs(9248) <= b;
    layer2_outputs(9249) <= b;
    layer2_outputs(9250) <= a;
    layer2_outputs(9251) <= not (a and b);
    layer2_outputs(9252) <= not b;
    layer2_outputs(9253) <= b;
    layer2_outputs(9254) <= not b;
    layer2_outputs(9255) <= a and not b;
    layer2_outputs(9256) <= a;
    layer2_outputs(9257) <= not b;
    layer2_outputs(9258) <= a;
    layer2_outputs(9259) <= a and not b;
    layer2_outputs(9260) <= a or b;
    layer2_outputs(9261) <= not a;
    layer2_outputs(9262) <= not b;
    layer2_outputs(9263) <= not a;
    layer2_outputs(9264) <= b and not a;
    layer2_outputs(9265) <= b;
    layer2_outputs(9266) <= a and b;
    layer2_outputs(9267) <= a and b;
    layer2_outputs(9268) <= not a or b;
    layer2_outputs(9269) <= not b;
    layer2_outputs(9270) <= not b;
    layer2_outputs(9271) <= a xor b;
    layer2_outputs(9272) <= not b;
    layer2_outputs(9273) <= b;
    layer2_outputs(9274) <= not b;
    layer2_outputs(9275) <= b;
    layer2_outputs(9276) <= not a;
    layer2_outputs(9277) <= a and b;
    layer2_outputs(9278) <= not a;
    layer2_outputs(9279) <= not b;
    layer2_outputs(9280) <= a xor b;
    layer2_outputs(9281) <= not (a and b);
    layer2_outputs(9282) <= a and not b;
    layer2_outputs(9283) <= not (a or b);
    layer2_outputs(9284) <= not a;
    layer2_outputs(9285) <= not a;
    layer2_outputs(9286) <= not (a xor b);
    layer2_outputs(9287) <= not (a or b);
    layer2_outputs(9288) <= a;
    layer2_outputs(9289) <= not b;
    layer2_outputs(9290) <= not (a xor b);
    layer2_outputs(9291) <= b;
    layer2_outputs(9292) <= a and b;
    layer2_outputs(9293) <= a;
    layer2_outputs(9294) <= not a;
    layer2_outputs(9295) <= not (a or b);
    layer2_outputs(9296) <= a and not b;
    layer2_outputs(9297) <= a;
    layer2_outputs(9298) <= not b or a;
    layer2_outputs(9299) <= b;
    layer2_outputs(9300) <= not a;
    layer2_outputs(9301) <= not (a or b);
    layer2_outputs(9302) <= b;
    layer2_outputs(9303) <= a and b;
    layer2_outputs(9304) <= a;
    layer2_outputs(9305) <= a and not b;
    layer2_outputs(9306) <= a;
    layer2_outputs(9307) <= a xor b;
    layer2_outputs(9308) <= not (a and b);
    layer2_outputs(9309) <= a and b;
    layer2_outputs(9310) <= a xor b;
    layer2_outputs(9311) <= b and not a;
    layer2_outputs(9312) <= a and not b;
    layer2_outputs(9313) <= a xor b;
    layer2_outputs(9314) <= b;
    layer2_outputs(9315) <= a or b;
    layer2_outputs(9316) <= b;
    layer2_outputs(9317) <= a and not b;
    layer2_outputs(9318) <= not a or b;
    layer2_outputs(9319) <= a and not b;
    layer2_outputs(9320) <= a or b;
    layer2_outputs(9321) <= a;
    layer2_outputs(9322) <= a or b;
    layer2_outputs(9323) <= not (a and b);
    layer2_outputs(9324) <= a and b;
    layer2_outputs(9325) <= not a;
    layer2_outputs(9326) <= a and b;
    layer2_outputs(9327) <= not (a xor b);
    layer2_outputs(9328) <= not b;
    layer2_outputs(9329) <= b;
    layer2_outputs(9330) <= not (a xor b);
    layer2_outputs(9331) <= not (a xor b);
    layer2_outputs(9332) <= not (a xor b);
    layer2_outputs(9333) <= a or b;
    layer2_outputs(9334) <= b;
    layer2_outputs(9335) <= a and b;
    layer2_outputs(9336) <= b and not a;
    layer2_outputs(9337) <= not a;
    layer2_outputs(9338) <= a and b;
    layer2_outputs(9339) <= b;
    layer2_outputs(9340) <= a;
    layer2_outputs(9341) <= 1'b1;
    layer2_outputs(9342) <= not (a or b);
    layer2_outputs(9343) <= b;
    layer2_outputs(9344) <= a and b;
    layer2_outputs(9345) <= b;
    layer2_outputs(9346) <= not (a xor b);
    layer2_outputs(9347) <= not a or b;
    layer2_outputs(9348) <= a and not b;
    layer2_outputs(9349) <= a xor b;
    layer2_outputs(9350) <= not a;
    layer2_outputs(9351) <= not b;
    layer2_outputs(9352) <= b;
    layer2_outputs(9353) <= not a;
    layer2_outputs(9354) <= b and not a;
    layer2_outputs(9355) <= a;
    layer2_outputs(9356) <= not a;
    layer2_outputs(9357) <= a;
    layer2_outputs(9358) <= a or b;
    layer2_outputs(9359) <= a xor b;
    layer2_outputs(9360) <= not a;
    layer2_outputs(9361) <= not (a xor b);
    layer2_outputs(9362) <= a;
    layer2_outputs(9363) <= b;
    layer2_outputs(9364) <= a and not b;
    layer2_outputs(9365) <= b and not a;
    layer2_outputs(9366) <= a and b;
    layer2_outputs(9367) <= not (a or b);
    layer2_outputs(9368) <= a;
    layer2_outputs(9369) <= not (a xor b);
    layer2_outputs(9370) <= not a or b;
    layer2_outputs(9371) <= not b;
    layer2_outputs(9372) <= not (a xor b);
    layer2_outputs(9373) <= not (a xor b);
    layer2_outputs(9374) <= not (a and b);
    layer2_outputs(9375) <= not a;
    layer2_outputs(9376) <= not b;
    layer2_outputs(9377) <= not b;
    layer2_outputs(9378) <= not (a xor b);
    layer2_outputs(9379) <= not a;
    layer2_outputs(9380) <= a xor b;
    layer2_outputs(9381) <= not (a and b);
    layer2_outputs(9382) <= not a;
    layer2_outputs(9383) <= not (a and b);
    layer2_outputs(9384) <= not b;
    layer2_outputs(9385) <= not (a xor b);
    layer2_outputs(9386) <= not a;
    layer2_outputs(9387) <= not b;
    layer2_outputs(9388) <= a;
    layer2_outputs(9389) <= a and b;
    layer2_outputs(9390) <= not b;
    layer2_outputs(9391) <= a;
    layer2_outputs(9392) <= not (a xor b);
    layer2_outputs(9393) <= a or b;
    layer2_outputs(9394) <= not b;
    layer2_outputs(9395) <= a or b;
    layer2_outputs(9396) <= not b;
    layer2_outputs(9397) <= a xor b;
    layer2_outputs(9398) <= a and not b;
    layer2_outputs(9399) <= not a;
    layer2_outputs(9400) <= b;
    layer2_outputs(9401) <= a;
    layer2_outputs(9402) <= a xor b;
    layer2_outputs(9403) <= not b or a;
    layer2_outputs(9404) <= not (a xor b);
    layer2_outputs(9405) <= a;
    layer2_outputs(9406) <= b;
    layer2_outputs(9407) <= not b or a;
    layer2_outputs(9408) <= b;
    layer2_outputs(9409) <= a;
    layer2_outputs(9410) <= a xor b;
    layer2_outputs(9411) <= b and not a;
    layer2_outputs(9412) <= a or b;
    layer2_outputs(9413) <= not (a xor b);
    layer2_outputs(9414) <= a and not b;
    layer2_outputs(9415) <= a;
    layer2_outputs(9416) <= a;
    layer2_outputs(9417) <= not a or b;
    layer2_outputs(9418) <= not b or a;
    layer2_outputs(9419) <= a xor b;
    layer2_outputs(9420) <= not (a xor b);
    layer2_outputs(9421) <= a and not b;
    layer2_outputs(9422) <= not (a xor b);
    layer2_outputs(9423) <= not (a xor b);
    layer2_outputs(9424) <= a and b;
    layer2_outputs(9425) <= a xor b;
    layer2_outputs(9426) <= not b;
    layer2_outputs(9427) <= b;
    layer2_outputs(9428) <= not (a xor b);
    layer2_outputs(9429) <= not b;
    layer2_outputs(9430) <= a xor b;
    layer2_outputs(9431) <= not b;
    layer2_outputs(9432) <= a and b;
    layer2_outputs(9433) <= a xor b;
    layer2_outputs(9434) <= a and not b;
    layer2_outputs(9435) <= not b;
    layer2_outputs(9436) <= not (a or b);
    layer2_outputs(9437) <= not (a xor b);
    layer2_outputs(9438) <= a;
    layer2_outputs(9439) <= not b;
    layer2_outputs(9440) <= b;
    layer2_outputs(9441) <= not b;
    layer2_outputs(9442) <= a;
    layer2_outputs(9443) <= not (a or b);
    layer2_outputs(9444) <= a and b;
    layer2_outputs(9445) <= b;
    layer2_outputs(9446) <= not a or b;
    layer2_outputs(9447) <= not b;
    layer2_outputs(9448) <= a xor b;
    layer2_outputs(9449) <= not (a or b);
    layer2_outputs(9450) <= a and b;
    layer2_outputs(9451) <= a xor b;
    layer2_outputs(9452) <= not a;
    layer2_outputs(9453) <= not b;
    layer2_outputs(9454) <= not a or b;
    layer2_outputs(9455) <= not (a xor b);
    layer2_outputs(9456) <= a xor b;
    layer2_outputs(9457) <= not (a or b);
    layer2_outputs(9458) <= a xor b;
    layer2_outputs(9459) <= a;
    layer2_outputs(9460) <= not b;
    layer2_outputs(9461) <= not (a and b);
    layer2_outputs(9462) <= b and not a;
    layer2_outputs(9463) <= a and not b;
    layer2_outputs(9464) <= not (a xor b);
    layer2_outputs(9465) <= a or b;
    layer2_outputs(9466) <= not b;
    layer2_outputs(9467) <= not a;
    layer2_outputs(9468) <= a;
    layer2_outputs(9469) <= not (a or b);
    layer2_outputs(9470) <= b and not a;
    layer2_outputs(9471) <= a and b;
    layer2_outputs(9472) <= a xor b;
    layer2_outputs(9473) <= a xor b;
    layer2_outputs(9474) <= not (a xor b);
    layer2_outputs(9475) <= a xor b;
    layer2_outputs(9476) <= a or b;
    layer2_outputs(9477) <= b and not a;
    layer2_outputs(9478) <= a and b;
    layer2_outputs(9479) <= a and b;
    layer2_outputs(9480) <= b;
    layer2_outputs(9481) <= a;
    layer2_outputs(9482) <= not b;
    layer2_outputs(9483) <= a xor b;
    layer2_outputs(9484) <= a xor b;
    layer2_outputs(9485) <= not b or a;
    layer2_outputs(9486) <= not b or a;
    layer2_outputs(9487) <= b;
    layer2_outputs(9488) <= a;
    layer2_outputs(9489) <= a or b;
    layer2_outputs(9490) <= a;
    layer2_outputs(9491) <= a xor b;
    layer2_outputs(9492) <= not b or a;
    layer2_outputs(9493) <= not b;
    layer2_outputs(9494) <= a xor b;
    layer2_outputs(9495) <= a and not b;
    layer2_outputs(9496) <= not (a or b);
    layer2_outputs(9497) <= a or b;
    layer2_outputs(9498) <= a xor b;
    layer2_outputs(9499) <= b and not a;
    layer2_outputs(9500) <= not (a or b);
    layer2_outputs(9501) <= not b;
    layer2_outputs(9502) <= a xor b;
    layer2_outputs(9503) <= a;
    layer2_outputs(9504) <= not (a and b);
    layer2_outputs(9505) <= a xor b;
    layer2_outputs(9506) <= b and not a;
    layer2_outputs(9507) <= a;
    layer2_outputs(9508) <= not a;
    layer2_outputs(9509) <= not b;
    layer2_outputs(9510) <= a xor b;
    layer2_outputs(9511) <= b;
    layer2_outputs(9512) <= not b;
    layer2_outputs(9513) <= a and b;
    layer2_outputs(9514) <= not a;
    layer2_outputs(9515) <= not a;
    layer2_outputs(9516) <= not a;
    layer2_outputs(9517) <= not b or a;
    layer2_outputs(9518) <= 1'b1;
    layer2_outputs(9519) <= not b;
    layer2_outputs(9520) <= a;
    layer2_outputs(9521) <= a xor b;
    layer2_outputs(9522) <= b;
    layer2_outputs(9523) <= not (a and b);
    layer2_outputs(9524) <= not a;
    layer2_outputs(9525) <= not b or a;
    layer2_outputs(9526) <= not (a and b);
    layer2_outputs(9527) <= not b;
    layer2_outputs(9528) <= not a;
    layer2_outputs(9529) <= 1'b1;
    layer2_outputs(9530) <= a and b;
    layer2_outputs(9531) <= not a;
    layer2_outputs(9532) <= not (a xor b);
    layer2_outputs(9533) <= b and not a;
    layer2_outputs(9534) <= a xor b;
    layer2_outputs(9535) <= not a or b;
    layer2_outputs(9536) <= a;
    layer2_outputs(9537) <= a xor b;
    layer2_outputs(9538) <= not (a xor b);
    layer2_outputs(9539) <= not (a or b);
    layer2_outputs(9540) <= not (a or b);
    layer2_outputs(9541) <= 1'b0;
    layer2_outputs(9542) <= not b;
    layer2_outputs(9543) <= a xor b;
    layer2_outputs(9544) <= b;
    layer2_outputs(9545) <= a xor b;
    layer2_outputs(9546) <= not a;
    layer2_outputs(9547) <= not (a and b);
    layer2_outputs(9548) <= not a;
    layer2_outputs(9549) <= not a;
    layer2_outputs(9550) <= not (a or b);
    layer2_outputs(9551) <= b;
    layer2_outputs(9552) <= not b;
    layer2_outputs(9553) <= a;
    layer2_outputs(9554) <= not b or a;
    layer2_outputs(9555) <= a and not b;
    layer2_outputs(9556) <= not a;
    layer2_outputs(9557) <= not b;
    layer2_outputs(9558) <= b and not a;
    layer2_outputs(9559) <= b;
    layer2_outputs(9560) <= not b or a;
    layer2_outputs(9561) <= b;
    layer2_outputs(9562) <= b;
    layer2_outputs(9563) <= a xor b;
    layer2_outputs(9564) <= a and b;
    layer2_outputs(9565) <= not a;
    layer2_outputs(9566) <= b;
    layer2_outputs(9567) <= not (a xor b);
    layer2_outputs(9568) <= not a or b;
    layer2_outputs(9569) <= not a;
    layer2_outputs(9570) <= not (a xor b);
    layer2_outputs(9571) <= b and not a;
    layer2_outputs(9572) <= a and not b;
    layer2_outputs(9573) <= not b;
    layer2_outputs(9574) <= a and not b;
    layer2_outputs(9575) <= not (a and b);
    layer2_outputs(9576) <= a and not b;
    layer2_outputs(9577) <= a xor b;
    layer2_outputs(9578) <= b;
    layer2_outputs(9579) <= a;
    layer2_outputs(9580) <= not b or a;
    layer2_outputs(9581) <= not (a xor b);
    layer2_outputs(9582) <= a xor b;
    layer2_outputs(9583) <= not a;
    layer2_outputs(9584) <= a or b;
    layer2_outputs(9585) <= a and not b;
    layer2_outputs(9586) <= a or b;
    layer2_outputs(9587) <= b;
    layer2_outputs(9588) <= b;
    layer2_outputs(9589) <= not (a xor b);
    layer2_outputs(9590) <= not a;
    layer2_outputs(9591) <= a xor b;
    layer2_outputs(9592) <= a and not b;
    layer2_outputs(9593) <= 1'b1;
    layer2_outputs(9594) <= a xor b;
    layer2_outputs(9595) <= a xor b;
    layer2_outputs(9596) <= b and not a;
    layer2_outputs(9597) <= not b;
    layer2_outputs(9598) <= not (a xor b);
    layer2_outputs(9599) <= not (a xor b);
    layer2_outputs(9600) <= not a;
    layer2_outputs(9601) <= not a;
    layer2_outputs(9602) <= a;
    layer2_outputs(9603) <= not (a xor b);
    layer2_outputs(9604) <= not b;
    layer2_outputs(9605) <= a and b;
    layer2_outputs(9606) <= a and not b;
    layer2_outputs(9607) <= not a;
    layer2_outputs(9608) <= not b;
    layer2_outputs(9609) <= a xor b;
    layer2_outputs(9610) <= not (a xor b);
    layer2_outputs(9611) <= not (a xor b);
    layer2_outputs(9612) <= not b or a;
    layer2_outputs(9613) <= not a;
    layer2_outputs(9614) <= a;
    layer2_outputs(9615) <= not b or a;
    layer2_outputs(9616) <= not (a xor b);
    layer2_outputs(9617) <= not b;
    layer2_outputs(9618) <= not b;
    layer2_outputs(9619) <= a xor b;
    layer2_outputs(9620) <= a and b;
    layer2_outputs(9621) <= not a;
    layer2_outputs(9622) <= not a;
    layer2_outputs(9623) <= not (a and b);
    layer2_outputs(9624) <= not (a and b);
    layer2_outputs(9625) <= b and not a;
    layer2_outputs(9626) <= a;
    layer2_outputs(9627) <= a xor b;
    layer2_outputs(9628) <= not b;
    layer2_outputs(9629) <= not a or b;
    layer2_outputs(9630) <= b;
    layer2_outputs(9631) <= a or b;
    layer2_outputs(9632) <= a and not b;
    layer2_outputs(9633) <= a xor b;
    layer2_outputs(9634) <= not a or b;
    layer2_outputs(9635) <= not b;
    layer2_outputs(9636) <= not a;
    layer2_outputs(9637) <= not a or b;
    layer2_outputs(9638) <= not (a xor b);
    layer2_outputs(9639) <= not a;
    layer2_outputs(9640) <= a or b;
    layer2_outputs(9641) <= not a;
    layer2_outputs(9642) <= a and b;
    layer2_outputs(9643) <= a or b;
    layer2_outputs(9644) <= a and b;
    layer2_outputs(9645) <= 1'b1;
    layer2_outputs(9646) <= not b;
    layer2_outputs(9647) <= b;
    layer2_outputs(9648) <= not (a xor b);
    layer2_outputs(9649) <= b;
    layer2_outputs(9650) <= a and b;
    layer2_outputs(9651) <= a;
    layer2_outputs(9652) <= not b;
    layer2_outputs(9653) <= not b;
    layer2_outputs(9654) <= a;
    layer2_outputs(9655) <= a;
    layer2_outputs(9656) <= not (a xor b);
    layer2_outputs(9657) <= not (a or b);
    layer2_outputs(9658) <= not (a xor b);
    layer2_outputs(9659) <= not a or b;
    layer2_outputs(9660) <= a and not b;
    layer2_outputs(9661) <= a and not b;
    layer2_outputs(9662) <= b;
    layer2_outputs(9663) <= a and not b;
    layer2_outputs(9664) <= a xor b;
    layer2_outputs(9665) <= not (a xor b);
    layer2_outputs(9666) <= not b or a;
    layer2_outputs(9667) <= a;
    layer2_outputs(9668) <= not a or b;
    layer2_outputs(9669) <= a xor b;
    layer2_outputs(9670) <= a and b;
    layer2_outputs(9671) <= b;
    layer2_outputs(9672) <= b;
    layer2_outputs(9673) <= a;
    layer2_outputs(9674) <= a;
    layer2_outputs(9675) <= not (a or b);
    layer2_outputs(9676) <= not (a or b);
    layer2_outputs(9677) <= not a;
    layer2_outputs(9678) <= b;
    layer2_outputs(9679) <= a;
    layer2_outputs(9680) <= a or b;
    layer2_outputs(9681) <= a xor b;
    layer2_outputs(9682) <= a xor b;
    layer2_outputs(9683) <= b;
    layer2_outputs(9684) <= a xor b;
    layer2_outputs(9685) <= b;
    layer2_outputs(9686) <= b;
    layer2_outputs(9687) <= not b or a;
    layer2_outputs(9688) <= not (a xor b);
    layer2_outputs(9689) <= not (a xor b);
    layer2_outputs(9690) <= b;
    layer2_outputs(9691) <= a;
    layer2_outputs(9692) <= a xor b;
    layer2_outputs(9693) <= a;
    layer2_outputs(9694) <= a;
    layer2_outputs(9695) <= a;
    layer2_outputs(9696) <= not a;
    layer2_outputs(9697) <= a and not b;
    layer2_outputs(9698) <= a or b;
    layer2_outputs(9699) <= not a;
    layer2_outputs(9700) <= not a or b;
    layer2_outputs(9701) <= a and b;
    layer2_outputs(9702) <= b;
    layer2_outputs(9703) <= a xor b;
    layer2_outputs(9704) <= b;
    layer2_outputs(9705) <= not b or a;
    layer2_outputs(9706) <= a xor b;
    layer2_outputs(9707) <= not (a xor b);
    layer2_outputs(9708) <= b and not a;
    layer2_outputs(9709) <= a and b;
    layer2_outputs(9710) <= a xor b;
    layer2_outputs(9711) <= not b;
    layer2_outputs(9712) <= a xor b;
    layer2_outputs(9713) <= b;
    layer2_outputs(9714) <= not b;
    layer2_outputs(9715) <= a xor b;
    layer2_outputs(9716) <= not a or b;
    layer2_outputs(9717) <= not (a and b);
    layer2_outputs(9718) <= b;
    layer2_outputs(9719) <= b;
    layer2_outputs(9720) <= not b;
    layer2_outputs(9721) <= not a;
    layer2_outputs(9722) <= not a;
    layer2_outputs(9723) <= a;
    layer2_outputs(9724) <= not (a xor b);
    layer2_outputs(9725) <= b;
    layer2_outputs(9726) <= not a or b;
    layer2_outputs(9727) <= a xor b;
    layer2_outputs(9728) <= not (a xor b);
    layer2_outputs(9729) <= b;
    layer2_outputs(9730) <= a and not b;
    layer2_outputs(9731) <= a or b;
    layer2_outputs(9732) <= not (a xor b);
    layer2_outputs(9733) <= a and not b;
    layer2_outputs(9734) <= not a;
    layer2_outputs(9735) <= not a;
    layer2_outputs(9736) <= a or b;
    layer2_outputs(9737) <= not (a xor b);
    layer2_outputs(9738) <= not b;
    layer2_outputs(9739) <= a and not b;
    layer2_outputs(9740) <= not (a or b);
    layer2_outputs(9741) <= not (a xor b);
    layer2_outputs(9742) <= b;
    layer2_outputs(9743) <= not a;
    layer2_outputs(9744) <= a;
    layer2_outputs(9745) <= not (a or b);
    layer2_outputs(9746) <= b;
    layer2_outputs(9747) <= a;
    layer2_outputs(9748) <= a;
    layer2_outputs(9749) <= not a or b;
    layer2_outputs(9750) <= b and not a;
    layer2_outputs(9751) <= b;
    layer2_outputs(9752) <= not b or a;
    layer2_outputs(9753) <= b and not a;
    layer2_outputs(9754) <= b;
    layer2_outputs(9755) <= a and not b;
    layer2_outputs(9756) <= a xor b;
    layer2_outputs(9757) <= not (a xor b);
    layer2_outputs(9758) <= not b;
    layer2_outputs(9759) <= not a;
    layer2_outputs(9760) <= not b;
    layer2_outputs(9761) <= not a or b;
    layer2_outputs(9762) <= a or b;
    layer2_outputs(9763) <= b and not a;
    layer2_outputs(9764) <= b;
    layer2_outputs(9765) <= not (a and b);
    layer2_outputs(9766) <= a and b;
    layer2_outputs(9767) <= not a;
    layer2_outputs(9768) <= b;
    layer2_outputs(9769) <= a xor b;
    layer2_outputs(9770) <= not b;
    layer2_outputs(9771) <= a or b;
    layer2_outputs(9772) <= not (a xor b);
    layer2_outputs(9773) <= not a;
    layer2_outputs(9774) <= a or b;
    layer2_outputs(9775) <= a;
    layer2_outputs(9776) <= not (a or b);
    layer2_outputs(9777) <= a;
    layer2_outputs(9778) <= a;
    layer2_outputs(9779) <= not (a and b);
    layer2_outputs(9780) <= not b or a;
    layer2_outputs(9781) <= not (a and b);
    layer2_outputs(9782) <= not (a xor b);
    layer2_outputs(9783) <= not (a xor b);
    layer2_outputs(9784) <= not a;
    layer2_outputs(9785) <= not b;
    layer2_outputs(9786) <= not a or b;
    layer2_outputs(9787) <= a xor b;
    layer2_outputs(9788) <= a;
    layer2_outputs(9789) <= a and b;
    layer2_outputs(9790) <= not a or b;
    layer2_outputs(9791) <= not (a xor b);
    layer2_outputs(9792) <= not a;
    layer2_outputs(9793) <= a and b;
    layer2_outputs(9794) <= not b;
    layer2_outputs(9795) <= not (a xor b);
    layer2_outputs(9796) <= not a or b;
    layer2_outputs(9797) <= a;
    layer2_outputs(9798) <= not a;
    layer2_outputs(9799) <= not a;
    layer2_outputs(9800) <= not (a or b);
    layer2_outputs(9801) <= a;
    layer2_outputs(9802) <= not a;
    layer2_outputs(9803) <= a xor b;
    layer2_outputs(9804) <= not a or b;
    layer2_outputs(9805) <= b;
    layer2_outputs(9806) <= not (a xor b);
    layer2_outputs(9807) <= not (a xor b);
    layer2_outputs(9808) <= not (a xor b);
    layer2_outputs(9809) <= not a;
    layer2_outputs(9810) <= not (a and b);
    layer2_outputs(9811) <= b;
    layer2_outputs(9812) <= not b;
    layer2_outputs(9813) <= not a;
    layer2_outputs(9814) <= not (a or b);
    layer2_outputs(9815) <= b;
    layer2_outputs(9816) <= a;
    layer2_outputs(9817) <= not (a and b);
    layer2_outputs(9818) <= a xor b;
    layer2_outputs(9819) <= b and not a;
    layer2_outputs(9820) <= not b;
    layer2_outputs(9821) <= not (a xor b);
    layer2_outputs(9822) <= a or b;
    layer2_outputs(9823) <= not b;
    layer2_outputs(9824) <= not (a xor b);
    layer2_outputs(9825) <= not a;
    layer2_outputs(9826) <= a and not b;
    layer2_outputs(9827) <= b;
    layer2_outputs(9828) <= 1'b0;
    layer2_outputs(9829) <= b and not a;
    layer2_outputs(9830) <= a xor b;
    layer2_outputs(9831) <= a xor b;
    layer2_outputs(9832) <= not (a xor b);
    layer2_outputs(9833) <= not a;
    layer2_outputs(9834) <= a and b;
    layer2_outputs(9835) <= not (a and b);
    layer2_outputs(9836) <= a xor b;
    layer2_outputs(9837) <= a and not b;
    layer2_outputs(9838) <= a and not b;
    layer2_outputs(9839) <= not (a or b);
    layer2_outputs(9840) <= not (a xor b);
    layer2_outputs(9841) <= not b;
    layer2_outputs(9842) <= not a or b;
    layer2_outputs(9843) <= b;
    layer2_outputs(9844) <= not a;
    layer2_outputs(9845) <= not b;
    layer2_outputs(9846) <= b;
    layer2_outputs(9847) <= not a or b;
    layer2_outputs(9848) <= a and not b;
    layer2_outputs(9849) <= a;
    layer2_outputs(9850) <= not a;
    layer2_outputs(9851) <= a xor b;
    layer2_outputs(9852) <= b;
    layer2_outputs(9853) <= a and not b;
    layer2_outputs(9854) <= a;
    layer2_outputs(9855) <= a or b;
    layer2_outputs(9856) <= a xor b;
    layer2_outputs(9857) <= not a;
    layer2_outputs(9858) <= 1'b1;
    layer2_outputs(9859) <= not a;
    layer2_outputs(9860) <= not (a or b);
    layer2_outputs(9861) <= a and b;
    layer2_outputs(9862) <= b and not a;
    layer2_outputs(9863) <= a and b;
    layer2_outputs(9864) <= a and b;
    layer2_outputs(9865) <= not b or a;
    layer2_outputs(9866) <= not (a xor b);
    layer2_outputs(9867) <= not a;
    layer2_outputs(9868) <= not a;
    layer2_outputs(9869) <= not (a xor b);
    layer2_outputs(9870) <= not a;
    layer2_outputs(9871) <= not (a and b);
    layer2_outputs(9872) <= b and not a;
    layer2_outputs(9873) <= a;
    layer2_outputs(9874) <= b;
    layer2_outputs(9875) <= a and b;
    layer2_outputs(9876) <= not b;
    layer2_outputs(9877) <= a;
    layer2_outputs(9878) <= not a or b;
    layer2_outputs(9879) <= not (a xor b);
    layer2_outputs(9880) <= b;
    layer2_outputs(9881) <= a xor b;
    layer2_outputs(9882) <= b and not a;
    layer2_outputs(9883) <= not (a xor b);
    layer2_outputs(9884) <= a xor b;
    layer2_outputs(9885) <= a and b;
    layer2_outputs(9886) <= not a;
    layer2_outputs(9887) <= not b or a;
    layer2_outputs(9888) <= not a;
    layer2_outputs(9889) <= not a;
    layer2_outputs(9890) <= not (a xor b);
    layer2_outputs(9891) <= 1'b0;
    layer2_outputs(9892) <= not (a or b);
    layer2_outputs(9893) <= not a;
    layer2_outputs(9894) <= not a or b;
    layer2_outputs(9895) <= a;
    layer2_outputs(9896) <= a and not b;
    layer2_outputs(9897) <= b;
    layer2_outputs(9898) <= a;
    layer2_outputs(9899) <= a and b;
    layer2_outputs(9900) <= b;
    layer2_outputs(9901) <= not a or b;
    layer2_outputs(9902) <= a;
    layer2_outputs(9903) <= b and not a;
    layer2_outputs(9904) <= not a;
    layer2_outputs(9905) <= a and b;
    layer2_outputs(9906) <= a and not b;
    layer2_outputs(9907) <= not (a xor b);
    layer2_outputs(9908) <= not a;
    layer2_outputs(9909) <= a and not b;
    layer2_outputs(9910) <= not b;
    layer2_outputs(9911) <= a;
    layer2_outputs(9912) <= not a or b;
    layer2_outputs(9913) <= a;
    layer2_outputs(9914) <= a;
    layer2_outputs(9915) <= a xor b;
    layer2_outputs(9916) <= not b;
    layer2_outputs(9917) <= not a;
    layer2_outputs(9918) <= 1'b0;
    layer2_outputs(9919) <= not (a and b);
    layer2_outputs(9920) <= a;
    layer2_outputs(9921) <= not b or a;
    layer2_outputs(9922) <= a;
    layer2_outputs(9923) <= not (a or b);
    layer2_outputs(9924) <= not (a xor b);
    layer2_outputs(9925) <= not b;
    layer2_outputs(9926) <= b;
    layer2_outputs(9927) <= not (a and b);
    layer2_outputs(9928) <= a and b;
    layer2_outputs(9929) <= a;
    layer2_outputs(9930) <= b;
    layer2_outputs(9931) <= a or b;
    layer2_outputs(9932) <= not a;
    layer2_outputs(9933) <= not (a or b);
    layer2_outputs(9934) <= not b;
    layer2_outputs(9935) <= a and b;
    layer2_outputs(9936) <= not (a xor b);
    layer2_outputs(9937) <= a and not b;
    layer2_outputs(9938) <= not a or b;
    layer2_outputs(9939) <= b;
    layer2_outputs(9940) <= a or b;
    layer2_outputs(9941) <= not (a xor b);
    layer2_outputs(9942) <= b;
    layer2_outputs(9943) <= not (a xor b);
    layer2_outputs(9944) <= not a or b;
    layer2_outputs(9945) <= a;
    layer2_outputs(9946) <= b and not a;
    layer2_outputs(9947) <= not b;
    layer2_outputs(9948) <= a and not b;
    layer2_outputs(9949) <= not (a xor b);
    layer2_outputs(9950) <= b;
    layer2_outputs(9951) <= a or b;
    layer2_outputs(9952) <= not b;
    layer2_outputs(9953) <= not b or a;
    layer2_outputs(9954) <= a xor b;
    layer2_outputs(9955) <= b;
    layer2_outputs(9956) <= not (a xor b);
    layer2_outputs(9957) <= not a or b;
    layer2_outputs(9958) <= not b;
    layer2_outputs(9959) <= not (a and b);
    layer2_outputs(9960) <= a and b;
    layer2_outputs(9961) <= b;
    layer2_outputs(9962) <= not a;
    layer2_outputs(9963) <= not b;
    layer2_outputs(9964) <= not (a xor b);
    layer2_outputs(9965) <= not b;
    layer2_outputs(9966) <= a;
    layer2_outputs(9967) <= a and not b;
    layer2_outputs(9968) <= a;
    layer2_outputs(9969) <= a and not b;
    layer2_outputs(9970) <= b;
    layer2_outputs(9971) <= a xor b;
    layer2_outputs(9972) <= not b;
    layer2_outputs(9973) <= a and not b;
    layer2_outputs(9974) <= not b;
    layer2_outputs(9975) <= a;
    layer2_outputs(9976) <= not a;
    layer2_outputs(9977) <= not b;
    layer2_outputs(9978) <= b;
    layer2_outputs(9979) <= not (a and b);
    layer2_outputs(9980) <= b and not a;
    layer2_outputs(9981) <= not a;
    layer2_outputs(9982) <= not b or a;
    layer2_outputs(9983) <= not b;
    layer2_outputs(9984) <= not b or a;
    layer2_outputs(9985) <= a;
    layer2_outputs(9986) <= b;
    layer2_outputs(9987) <= not a or b;
    layer2_outputs(9988) <= a;
    layer2_outputs(9989) <= a xor b;
    layer2_outputs(9990) <= a and not b;
    layer2_outputs(9991) <= a;
    layer2_outputs(9992) <= not (a and b);
    layer2_outputs(9993) <= not (a or b);
    layer2_outputs(9994) <= not a or b;
    layer2_outputs(9995) <= a and b;
    layer2_outputs(9996) <= not (a xor b);
    layer2_outputs(9997) <= a;
    layer2_outputs(9998) <= not (a xor b);
    layer2_outputs(9999) <= not (a xor b);
    layer2_outputs(10000) <= not (a xor b);
    layer2_outputs(10001) <= not a;
    layer2_outputs(10002) <= not (a xor b);
    layer2_outputs(10003) <= a;
    layer2_outputs(10004) <= not a or b;
    layer2_outputs(10005) <= not b;
    layer2_outputs(10006) <= b and not a;
    layer2_outputs(10007) <= a or b;
    layer2_outputs(10008) <= b;
    layer2_outputs(10009) <= a or b;
    layer2_outputs(10010) <= a xor b;
    layer2_outputs(10011) <= not a;
    layer2_outputs(10012) <= not a;
    layer2_outputs(10013) <= not (a and b);
    layer2_outputs(10014) <= not (a or b);
    layer2_outputs(10015) <= a;
    layer2_outputs(10016) <= not b;
    layer2_outputs(10017) <= not b;
    layer2_outputs(10018) <= b and not a;
    layer2_outputs(10019) <= b and not a;
    layer2_outputs(10020) <= a;
    layer2_outputs(10021) <= not a;
    layer2_outputs(10022) <= not b;
    layer2_outputs(10023) <= not a;
    layer2_outputs(10024) <= not b or a;
    layer2_outputs(10025) <= b;
    layer2_outputs(10026) <= not (a and b);
    layer2_outputs(10027) <= a xor b;
    layer2_outputs(10028) <= a or b;
    layer2_outputs(10029) <= not (a xor b);
    layer2_outputs(10030) <= not (a xor b);
    layer2_outputs(10031) <= a or b;
    layer2_outputs(10032) <= not (a xor b);
    layer2_outputs(10033) <= b;
    layer2_outputs(10034) <= not (a xor b);
    layer2_outputs(10035) <= b and not a;
    layer2_outputs(10036) <= a or b;
    layer2_outputs(10037) <= not a;
    layer2_outputs(10038) <= not b or a;
    layer2_outputs(10039) <= a;
    layer2_outputs(10040) <= not a;
    layer2_outputs(10041) <= b;
    layer2_outputs(10042) <= a and not b;
    layer2_outputs(10043) <= a xor b;
    layer2_outputs(10044) <= not b or a;
    layer2_outputs(10045) <= a xor b;
    layer2_outputs(10046) <= b;
    layer2_outputs(10047) <= not a;
    layer2_outputs(10048) <= a xor b;
    layer2_outputs(10049) <= not a or b;
    layer2_outputs(10050) <= b;
    layer2_outputs(10051) <= a and b;
    layer2_outputs(10052) <= not (a and b);
    layer2_outputs(10053) <= not (a or b);
    layer2_outputs(10054) <= a xor b;
    layer2_outputs(10055) <= not (a and b);
    layer2_outputs(10056) <= a xor b;
    layer2_outputs(10057) <= a;
    layer2_outputs(10058) <= not (a xor b);
    layer2_outputs(10059) <= b;
    layer2_outputs(10060) <= not b or a;
    layer2_outputs(10061) <= not (a xor b);
    layer2_outputs(10062) <= a or b;
    layer2_outputs(10063) <= not b or a;
    layer2_outputs(10064) <= not a;
    layer2_outputs(10065) <= not a;
    layer2_outputs(10066) <= not (a and b);
    layer2_outputs(10067) <= a xor b;
    layer2_outputs(10068) <= a;
    layer2_outputs(10069) <= a;
    layer2_outputs(10070) <= a;
    layer2_outputs(10071) <= not (a xor b);
    layer2_outputs(10072) <= not b;
    layer2_outputs(10073) <= b;
    layer2_outputs(10074) <= a;
    layer2_outputs(10075) <= not b or a;
    layer2_outputs(10076) <= not b or a;
    layer2_outputs(10077) <= not a or b;
    layer2_outputs(10078) <= not b or a;
    layer2_outputs(10079) <= a xor b;
    layer2_outputs(10080) <= b;
    layer2_outputs(10081) <= b;
    layer2_outputs(10082) <= not a;
    layer2_outputs(10083) <= a xor b;
    layer2_outputs(10084) <= b;
    layer2_outputs(10085) <= a;
    layer2_outputs(10086) <= not a;
    layer2_outputs(10087) <= b;
    layer2_outputs(10088) <= a;
    layer2_outputs(10089) <= not b;
    layer2_outputs(10090) <= b;
    layer2_outputs(10091) <= not (a xor b);
    layer2_outputs(10092) <= a xor b;
    layer2_outputs(10093) <= a xor b;
    layer2_outputs(10094) <= not a or b;
    layer2_outputs(10095) <= a xor b;
    layer2_outputs(10096) <= a xor b;
    layer2_outputs(10097) <= a or b;
    layer2_outputs(10098) <= not (a xor b);
    layer2_outputs(10099) <= not (a or b);
    layer2_outputs(10100) <= not (a xor b);
    layer2_outputs(10101) <= a xor b;
    layer2_outputs(10102) <= a;
    layer2_outputs(10103) <= not b;
    layer2_outputs(10104) <= b;
    layer2_outputs(10105) <= b;
    layer2_outputs(10106) <= not b;
    layer2_outputs(10107) <= not a;
    layer2_outputs(10108) <= a;
    layer2_outputs(10109) <= a xor b;
    layer2_outputs(10110) <= a or b;
    layer2_outputs(10111) <= a and b;
    layer2_outputs(10112) <= not b or a;
    layer2_outputs(10113) <= b and not a;
    layer2_outputs(10114) <= not (a or b);
    layer2_outputs(10115) <= a;
    layer2_outputs(10116) <= not a;
    layer2_outputs(10117) <= b;
    layer2_outputs(10118) <= a;
    layer2_outputs(10119) <= b;
    layer2_outputs(10120) <= a xor b;
    layer2_outputs(10121) <= a and b;
    layer2_outputs(10122) <= not (a and b);
    layer2_outputs(10123) <= b;
    layer2_outputs(10124) <= not a or b;
    layer2_outputs(10125) <= b and not a;
    layer2_outputs(10126) <= not (a xor b);
    layer2_outputs(10127) <= not b;
    layer2_outputs(10128) <= not a;
    layer2_outputs(10129) <= not (a and b);
    layer2_outputs(10130) <= a and not b;
    layer2_outputs(10131) <= a;
    layer2_outputs(10132) <= not a;
    layer2_outputs(10133) <= not (a or b);
    layer2_outputs(10134) <= not a or b;
    layer2_outputs(10135) <= a or b;
    layer2_outputs(10136) <= not a or b;
    layer2_outputs(10137) <= a xor b;
    layer2_outputs(10138) <= not (a xor b);
    layer2_outputs(10139) <= not b or a;
    layer2_outputs(10140) <= a and b;
    layer2_outputs(10141) <= b;
    layer2_outputs(10142) <= not b or a;
    layer2_outputs(10143) <= b and not a;
    layer2_outputs(10144) <= a xor b;
    layer2_outputs(10145) <= b;
    layer2_outputs(10146) <= b;
    layer2_outputs(10147) <= a;
    layer2_outputs(10148) <= not a;
    layer2_outputs(10149) <= a or b;
    layer2_outputs(10150) <= not a;
    layer2_outputs(10151) <= not a;
    layer2_outputs(10152) <= not b;
    layer2_outputs(10153) <= a;
    layer2_outputs(10154) <= not (a xor b);
    layer2_outputs(10155) <= a or b;
    layer2_outputs(10156) <= not (a xor b);
    layer2_outputs(10157) <= b;
    layer2_outputs(10158) <= b;
    layer2_outputs(10159) <= a and not b;
    layer2_outputs(10160) <= not b;
    layer2_outputs(10161) <= a;
    layer2_outputs(10162) <= b;
    layer2_outputs(10163) <= not b or a;
    layer2_outputs(10164) <= not a;
    layer2_outputs(10165) <= a;
    layer2_outputs(10166) <= not a;
    layer2_outputs(10167) <= a and not b;
    layer2_outputs(10168) <= not a;
    layer2_outputs(10169) <= a xor b;
    layer2_outputs(10170) <= a and not b;
    layer2_outputs(10171) <= b;
    layer2_outputs(10172) <= a xor b;
    layer2_outputs(10173) <= not (a or b);
    layer2_outputs(10174) <= a or b;
    layer2_outputs(10175) <= not (a xor b);
    layer2_outputs(10176) <= b and not a;
    layer2_outputs(10177) <= not (a and b);
    layer2_outputs(10178) <= not (a xor b);
    layer2_outputs(10179) <= a;
    layer2_outputs(10180) <= b;
    layer2_outputs(10181) <= not a;
    layer2_outputs(10182) <= not a;
    layer2_outputs(10183) <= not (a and b);
    layer2_outputs(10184) <= a;
    layer2_outputs(10185) <= a xor b;
    layer2_outputs(10186) <= not a;
    layer2_outputs(10187) <= a and not b;
    layer2_outputs(10188) <= not a or b;
    layer2_outputs(10189) <= not (a and b);
    layer2_outputs(10190) <= not b;
    layer2_outputs(10191) <= not a;
    layer2_outputs(10192) <= a;
    layer2_outputs(10193) <= not a;
    layer2_outputs(10194) <= a or b;
    layer2_outputs(10195) <= b;
    layer2_outputs(10196) <= not a or b;
    layer2_outputs(10197) <= a xor b;
    layer2_outputs(10198) <= not (a and b);
    layer2_outputs(10199) <= a xor b;
    layer2_outputs(10200) <= a;
    layer2_outputs(10201) <= not (a and b);
    layer2_outputs(10202) <= not (a and b);
    layer2_outputs(10203) <= b and not a;
    layer2_outputs(10204) <= a;
    layer2_outputs(10205) <= a xor b;
    layer2_outputs(10206) <= a;
    layer2_outputs(10207) <= a xor b;
    layer2_outputs(10208) <= a xor b;
    layer2_outputs(10209) <= a xor b;
    layer2_outputs(10210) <= a;
    layer2_outputs(10211) <= not a or b;
    layer2_outputs(10212) <= not b;
    layer2_outputs(10213) <= not b;
    layer2_outputs(10214) <= b;
    layer2_outputs(10215) <= not (a xor b);
    layer2_outputs(10216) <= a xor b;
    layer2_outputs(10217) <= b and not a;
    layer2_outputs(10218) <= not a;
    layer2_outputs(10219) <= a and not b;
    layer2_outputs(10220) <= a or b;
    layer2_outputs(10221) <= b;
    layer2_outputs(10222) <= b;
    layer2_outputs(10223) <= not a;
    layer2_outputs(10224) <= a;
    layer2_outputs(10225) <= b;
    layer2_outputs(10226) <= not (a xor b);
    layer2_outputs(10227) <= not a;
    layer2_outputs(10228) <= b;
    layer2_outputs(10229) <= b;
    layer2_outputs(10230) <= not b or a;
    layer2_outputs(10231) <= not b;
    layer2_outputs(10232) <= a and b;
    layer2_outputs(10233) <= not b;
    layer2_outputs(10234) <= not a;
    layer2_outputs(10235) <= b and not a;
    layer2_outputs(10236) <= a and not b;
    layer2_outputs(10237) <= a and b;
    layer2_outputs(10238) <= b;
    layer2_outputs(10239) <= a and not b;
    layer2_outputs(10240) <= not (a xor b);
    layer2_outputs(10241) <= not a or b;
    layer2_outputs(10242) <= not (a xor b);
    layer2_outputs(10243) <= not (a and b);
    layer2_outputs(10244) <= a and b;
    layer2_outputs(10245) <= not a or b;
    layer2_outputs(10246) <= not (a xor b);
    layer2_outputs(10247) <= not a;
    layer2_outputs(10248) <= not (a xor b);
    layer2_outputs(10249) <= not a;
    layer2_outputs(10250) <= a xor b;
    layer2_outputs(10251) <= not a or b;
    layer2_outputs(10252) <= not (a and b);
    layer2_outputs(10253) <= a;
    layer2_outputs(10254) <= a xor b;
    layer2_outputs(10255) <= a and not b;
    layer2_outputs(10256) <= a and not b;
    layer2_outputs(10257) <= not a;
    layer2_outputs(10258) <= not (a and b);
    layer2_outputs(10259) <= not (a and b);
    layer2_outputs(10260) <= a;
    layer2_outputs(10261) <= not (a xor b);
    layer2_outputs(10262) <= a and not b;
    layer2_outputs(10263) <= b and not a;
    layer2_outputs(10264) <= b;
    layer2_outputs(10265) <= not a;
    layer2_outputs(10266) <= b;
    layer2_outputs(10267) <= b;
    layer2_outputs(10268) <= not (a or b);
    layer2_outputs(10269) <= not b or a;
    layer2_outputs(10270) <= not b or a;
    layer2_outputs(10271) <= a and not b;
    layer2_outputs(10272) <= not a or b;
    layer2_outputs(10273) <= not (a or b);
    layer2_outputs(10274) <= a or b;
    layer2_outputs(10275) <= not b;
    layer2_outputs(10276) <= a and b;
    layer2_outputs(10277) <= not (a and b);
    layer2_outputs(10278) <= a;
    layer2_outputs(10279) <= not a;
    layer2_outputs(10280) <= not a;
    layer2_outputs(10281) <= not (a or b);
    layer2_outputs(10282) <= not (a xor b);
    layer2_outputs(10283) <= a and not b;
    layer2_outputs(10284) <= not (a and b);
    layer2_outputs(10285) <= b and not a;
    layer2_outputs(10286) <= not (a xor b);
    layer2_outputs(10287) <= not (a xor b);
    layer2_outputs(10288) <= not (a and b);
    layer2_outputs(10289) <= b;
    layer2_outputs(10290) <= not b;
    layer2_outputs(10291) <= a xor b;
    layer2_outputs(10292) <= not (a xor b);
    layer2_outputs(10293) <= not b;
    layer2_outputs(10294) <= a;
    layer2_outputs(10295) <= b and not a;
    layer2_outputs(10296) <= a xor b;
    layer2_outputs(10297) <= a xor b;
    layer2_outputs(10298) <= not a or b;
    layer2_outputs(10299) <= b;
    layer2_outputs(10300) <= a;
    layer2_outputs(10301) <= b;
    layer2_outputs(10302) <= b;
    layer2_outputs(10303) <= not (a xor b);
    layer2_outputs(10304) <= a and not b;
    layer2_outputs(10305) <= not b;
    layer2_outputs(10306) <= a;
    layer2_outputs(10307) <= not b;
    layer2_outputs(10308) <= b;
    layer2_outputs(10309) <= not b or a;
    layer2_outputs(10310) <= b and not a;
    layer2_outputs(10311) <= a;
    layer2_outputs(10312) <= a and not b;
    layer2_outputs(10313) <= not (a xor b);
    layer2_outputs(10314) <= not b or a;
    layer2_outputs(10315) <= b;
    layer2_outputs(10316) <= a;
    layer2_outputs(10317) <= not a or b;
    layer2_outputs(10318) <= a;
    layer2_outputs(10319) <= not b;
    layer2_outputs(10320) <= a xor b;
    layer2_outputs(10321) <= not (a xor b);
    layer2_outputs(10322) <= a xor b;
    layer2_outputs(10323) <= not a;
    layer2_outputs(10324) <= not (a xor b);
    layer2_outputs(10325) <= not a;
    layer2_outputs(10326) <= b and not a;
    layer2_outputs(10327) <= a and b;
    layer2_outputs(10328) <= b;
    layer2_outputs(10329) <= not a;
    layer2_outputs(10330) <= a xor b;
    layer2_outputs(10331) <= b;
    layer2_outputs(10332) <= not b;
    layer2_outputs(10333) <= b and not a;
    layer2_outputs(10334) <= a and b;
    layer2_outputs(10335) <= b;
    layer2_outputs(10336) <= a xor b;
    layer2_outputs(10337) <= not (a xor b);
    layer2_outputs(10338) <= b;
    layer2_outputs(10339) <= not (a and b);
    layer2_outputs(10340) <= a and not b;
    layer2_outputs(10341) <= b;
    layer2_outputs(10342) <= b;
    layer2_outputs(10343) <= not b;
    layer2_outputs(10344) <= not b;
    layer2_outputs(10345) <= not a or b;
    layer2_outputs(10346) <= not b;
    layer2_outputs(10347) <= a;
    layer2_outputs(10348) <= not a;
    layer2_outputs(10349) <= a xor b;
    layer2_outputs(10350) <= not (a xor b);
    layer2_outputs(10351) <= not (a xor b);
    layer2_outputs(10352) <= a xor b;
    layer2_outputs(10353) <= not b or a;
    layer2_outputs(10354) <= a;
    layer2_outputs(10355) <= not b;
    layer2_outputs(10356) <= not a;
    layer2_outputs(10357) <= a xor b;
    layer2_outputs(10358) <= not b;
    layer2_outputs(10359) <= b;
    layer2_outputs(10360) <= a xor b;
    layer2_outputs(10361) <= not b or a;
    layer2_outputs(10362) <= not (a or b);
    layer2_outputs(10363) <= b;
    layer2_outputs(10364) <= not a or b;
    layer2_outputs(10365) <= not (a xor b);
    layer2_outputs(10366) <= a;
    layer2_outputs(10367) <= not b;
    layer2_outputs(10368) <= b;
    layer2_outputs(10369) <= not (a xor b);
    layer2_outputs(10370) <= not b;
    layer2_outputs(10371) <= b;
    layer2_outputs(10372) <= b;
    layer2_outputs(10373) <= not b;
    layer2_outputs(10374) <= not a;
    layer2_outputs(10375) <= not (a or b);
    layer2_outputs(10376) <= not b;
    layer2_outputs(10377) <= not a;
    layer2_outputs(10378) <= not b;
    layer2_outputs(10379) <= not (a and b);
    layer2_outputs(10380) <= a xor b;
    layer2_outputs(10381) <= a or b;
    layer2_outputs(10382) <= a;
    layer2_outputs(10383) <= not (a xor b);
    layer2_outputs(10384) <= b;
    layer2_outputs(10385) <= a xor b;
    layer2_outputs(10386) <= not (a or b);
    layer2_outputs(10387) <= not (a and b);
    layer2_outputs(10388) <= not (a xor b);
    layer2_outputs(10389) <= a xor b;
    layer2_outputs(10390) <= not (a and b);
    layer2_outputs(10391) <= b;
    layer2_outputs(10392) <= a xor b;
    layer2_outputs(10393) <= a xor b;
    layer2_outputs(10394) <= not b;
    layer2_outputs(10395) <= not a;
    layer2_outputs(10396) <= a xor b;
    layer2_outputs(10397) <= not (a xor b);
    layer2_outputs(10398) <= not a;
    layer2_outputs(10399) <= not a or b;
    layer2_outputs(10400) <= a;
    layer2_outputs(10401) <= not a or b;
    layer2_outputs(10402) <= not a;
    layer2_outputs(10403) <= 1'b0;
    layer2_outputs(10404) <= a or b;
    layer2_outputs(10405) <= not a or b;
    layer2_outputs(10406) <= a xor b;
    layer2_outputs(10407) <= not b or a;
    layer2_outputs(10408) <= b;
    layer2_outputs(10409) <= a and not b;
    layer2_outputs(10410) <= a and not b;
    layer2_outputs(10411) <= not (a xor b);
    layer2_outputs(10412) <= not (a xor b);
    layer2_outputs(10413) <= not (a and b);
    layer2_outputs(10414) <= a and b;
    layer2_outputs(10415) <= a xor b;
    layer2_outputs(10416) <= not (a and b);
    layer2_outputs(10417) <= not (a and b);
    layer2_outputs(10418) <= not a or b;
    layer2_outputs(10419) <= not (a or b);
    layer2_outputs(10420) <= not b or a;
    layer2_outputs(10421) <= not b or a;
    layer2_outputs(10422) <= a and b;
    layer2_outputs(10423) <= not b;
    layer2_outputs(10424) <= not b;
    layer2_outputs(10425) <= not a or b;
    layer2_outputs(10426) <= a xor b;
    layer2_outputs(10427) <= a or b;
    layer2_outputs(10428) <= not (a xor b);
    layer2_outputs(10429) <= not b;
    layer2_outputs(10430) <= not b;
    layer2_outputs(10431) <= a xor b;
    layer2_outputs(10432) <= not b or a;
    layer2_outputs(10433) <= a xor b;
    layer2_outputs(10434) <= not b;
    layer2_outputs(10435) <= b;
    layer2_outputs(10436) <= a;
    layer2_outputs(10437) <= b;
    layer2_outputs(10438) <= not a;
    layer2_outputs(10439) <= b and not a;
    layer2_outputs(10440) <= a xor b;
    layer2_outputs(10441) <= not b;
    layer2_outputs(10442) <= a and b;
    layer2_outputs(10443) <= a;
    layer2_outputs(10444) <= not b or a;
    layer2_outputs(10445) <= a and b;
    layer2_outputs(10446) <= b and not a;
    layer2_outputs(10447) <= not a or b;
    layer2_outputs(10448) <= a;
    layer2_outputs(10449) <= a;
    layer2_outputs(10450) <= not (a xor b);
    layer2_outputs(10451) <= a;
    layer2_outputs(10452) <= not (a xor b);
    layer2_outputs(10453) <= a;
    layer2_outputs(10454) <= a or b;
    layer2_outputs(10455) <= a and not b;
    layer2_outputs(10456) <= not a or b;
    layer2_outputs(10457) <= not (a xor b);
    layer2_outputs(10458) <= a and not b;
    layer2_outputs(10459) <= not (a xor b);
    layer2_outputs(10460) <= b and not a;
    layer2_outputs(10461) <= not (a xor b);
    layer2_outputs(10462) <= a and not b;
    layer2_outputs(10463) <= a and b;
    layer2_outputs(10464) <= 1'b1;
    layer2_outputs(10465) <= b and not a;
    layer2_outputs(10466) <= not (a and b);
    layer2_outputs(10467) <= a or b;
    layer2_outputs(10468) <= not a;
    layer2_outputs(10469) <= not (a and b);
    layer2_outputs(10470) <= not (a xor b);
    layer2_outputs(10471) <= a or b;
    layer2_outputs(10472) <= a;
    layer2_outputs(10473) <= not (a or b);
    layer2_outputs(10474) <= b;
    layer2_outputs(10475) <= not (a xor b);
    layer2_outputs(10476) <= a or b;
    layer2_outputs(10477) <= b;
    layer2_outputs(10478) <= not a;
    layer2_outputs(10479) <= not a or b;
    layer2_outputs(10480) <= b;
    layer2_outputs(10481) <= not b;
    layer2_outputs(10482) <= not b or a;
    layer2_outputs(10483) <= b;
    layer2_outputs(10484) <= a;
    layer2_outputs(10485) <= a xor b;
    layer2_outputs(10486) <= a;
    layer2_outputs(10487) <= not a;
    layer2_outputs(10488) <= not b;
    layer2_outputs(10489) <= a and b;
    layer2_outputs(10490) <= a xor b;
    layer2_outputs(10491) <= not (a xor b);
    layer2_outputs(10492) <= a xor b;
    layer2_outputs(10493) <= b and not a;
    layer2_outputs(10494) <= a;
    layer2_outputs(10495) <= not (a xor b);
    layer2_outputs(10496) <= a and b;
    layer2_outputs(10497) <= not a;
    layer2_outputs(10498) <= not (a xor b);
    layer2_outputs(10499) <= not (a and b);
    layer2_outputs(10500) <= a;
    layer2_outputs(10501) <= a;
    layer2_outputs(10502) <= a xor b;
    layer2_outputs(10503) <= not a or b;
    layer2_outputs(10504) <= a and b;
    layer2_outputs(10505) <= a;
    layer2_outputs(10506) <= a or b;
    layer2_outputs(10507) <= a and b;
    layer2_outputs(10508) <= a and not b;
    layer2_outputs(10509) <= a xor b;
    layer2_outputs(10510) <= not b;
    layer2_outputs(10511) <= not b;
    layer2_outputs(10512) <= a;
    layer2_outputs(10513) <= a;
    layer2_outputs(10514) <= not b;
    layer2_outputs(10515) <= a;
    layer2_outputs(10516) <= not b or a;
    layer2_outputs(10517) <= not (a and b);
    layer2_outputs(10518) <= a and not b;
    layer2_outputs(10519) <= a and b;
    layer2_outputs(10520) <= not b or a;
    layer2_outputs(10521) <= not (a and b);
    layer2_outputs(10522) <= not b or a;
    layer2_outputs(10523) <= not (a xor b);
    layer2_outputs(10524) <= not a or b;
    layer2_outputs(10525) <= a and not b;
    layer2_outputs(10526) <= a xor b;
    layer2_outputs(10527) <= a or b;
    layer2_outputs(10528) <= not (a or b);
    layer2_outputs(10529) <= not (a and b);
    layer2_outputs(10530) <= a or b;
    layer2_outputs(10531) <= a and not b;
    layer2_outputs(10532) <= a;
    layer2_outputs(10533) <= not b or a;
    layer2_outputs(10534) <= not a or b;
    layer2_outputs(10535) <= a;
    layer2_outputs(10536) <= a;
    layer2_outputs(10537) <= b;
    layer2_outputs(10538) <= not (a and b);
    layer2_outputs(10539) <= not b;
    layer2_outputs(10540) <= a;
    layer2_outputs(10541) <= a;
    layer2_outputs(10542) <= not b or a;
    layer2_outputs(10543) <= not a or b;
    layer2_outputs(10544) <= not (a and b);
    layer2_outputs(10545) <= b;
    layer2_outputs(10546) <= not b;
    layer2_outputs(10547) <= b;
    layer2_outputs(10548) <= a;
    layer2_outputs(10549) <= b;
    layer2_outputs(10550) <= b;
    layer2_outputs(10551) <= a;
    layer2_outputs(10552) <= not (a and b);
    layer2_outputs(10553) <= not b;
    layer2_outputs(10554) <= a and b;
    layer2_outputs(10555) <= a xor b;
    layer2_outputs(10556) <= a or b;
    layer2_outputs(10557) <= 1'b1;
    layer2_outputs(10558) <= b;
    layer2_outputs(10559) <= not b;
    layer2_outputs(10560) <= b and not a;
    layer2_outputs(10561) <= not (a xor b);
    layer2_outputs(10562) <= a or b;
    layer2_outputs(10563) <= a;
    layer2_outputs(10564) <= not a;
    layer2_outputs(10565) <= not b;
    layer2_outputs(10566) <= a xor b;
    layer2_outputs(10567) <= not (a xor b);
    layer2_outputs(10568) <= a and not b;
    layer2_outputs(10569) <= a;
    layer2_outputs(10570) <= not b;
    layer2_outputs(10571) <= not (a or b);
    layer2_outputs(10572) <= b;
    layer2_outputs(10573) <= b and not a;
    layer2_outputs(10574) <= not a or b;
    layer2_outputs(10575) <= b;
    layer2_outputs(10576) <= a and b;
    layer2_outputs(10577) <= b;
    layer2_outputs(10578) <= not (a xor b);
    layer2_outputs(10579) <= a;
    layer2_outputs(10580) <= a;
    layer2_outputs(10581) <= not (a or b);
    layer2_outputs(10582) <= not a or b;
    layer2_outputs(10583) <= a or b;
    layer2_outputs(10584) <= b and not a;
    layer2_outputs(10585) <= b;
    layer2_outputs(10586) <= not a;
    layer2_outputs(10587) <= not (a xor b);
    layer2_outputs(10588) <= b;
    layer2_outputs(10589) <= not b;
    layer2_outputs(10590) <= a and not b;
    layer2_outputs(10591) <= a;
    layer2_outputs(10592) <= not (a xor b);
    layer2_outputs(10593) <= b;
    layer2_outputs(10594) <= not (a or b);
    layer2_outputs(10595) <= not b;
    layer2_outputs(10596) <= not (a xor b);
    layer2_outputs(10597) <= not a;
    layer2_outputs(10598) <= a;
    layer2_outputs(10599) <= not b;
    layer2_outputs(10600) <= a;
    layer2_outputs(10601) <= a;
    layer2_outputs(10602) <= a;
    layer2_outputs(10603) <= not (a or b);
    layer2_outputs(10604) <= not a;
    layer2_outputs(10605) <= a xor b;
    layer2_outputs(10606) <= not a;
    layer2_outputs(10607) <= a and b;
    layer2_outputs(10608) <= not a or b;
    layer2_outputs(10609) <= b;
    layer2_outputs(10610) <= not a or b;
    layer2_outputs(10611) <= not b or a;
    layer2_outputs(10612) <= b;
    layer2_outputs(10613) <= not b or a;
    layer2_outputs(10614) <= not (a xor b);
    layer2_outputs(10615) <= a xor b;
    layer2_outputs(10616) <= not (a xor b);
    layer2_outputs(10617) <= not a or b;
    layer2_outputs(10618) <= not b;
    layer2_outputs(10619) <= not (a or b);
    layer2_outputs(10620) <= a xor b;
    layer2_outputs(10621) <= not b;
    layer2_outputs(10622) <= a xor b;
    layer2_outputs(10623) <= not b or a;
    layer2_outputs(10624) <= a or b;
    layer2_outputs(10625) <= a;
    layer2_outputs(10626) <= 1'b0;
    layer2_outputs(10627) <= not a;
    layer2_outputs(10628) <= not b;
    layer2_outputs(10629) <= b and not a;
    layer2_outputs(10630) <= not (a xor b);
    layer2_outputs(10631) <= b;
    layer2_outputs(10632) <= a xor b;
    layer2_outputs(10633) <= not b;
    layer2_outputs(10634) <= not (a and b);
    layer2_outputs(10635) <= not (a and b);
    layer2_outputs(10636) <= not b;
    layer2_outputs(10637) <= not a;
    layer2_outputs(10638) <= a;
    layer2_outputs(10639) <= b and not a;
    layer2_outputs(10640) <= a xor b;
    layer2_outputs(10641) <= not (a and b);
    layer2_outputs(10642) <= a;
    layer2_outputs(10643) <= a and not b;
    layer2_outputs(10644) <= not (a or b);
    layer2_outputs(10645) <= a xor b;
    layer2_outputs(10646) <= not b;
    layer2_outputs(10647) <= b and not a;
    layer2_outputs(10648) <= a;
    layer2_outputs(10649) <= a;
    layer2_outputs(10650) <= a xor b;
    layer2_outputs(10651) <= not (a xor b);
    layer2_outputs(10652) <= not a;
    layer2_outputs(10653) <= not a or b;
    layer2_outputs(10654) <= a xor b;
    layer2_outputs(10655) <= a or b;
    layer2_outputs(10656) <= a and not b;
    layer2_outputs(10657) <= not (a and b);
    layer2_outputs(10658) <= not (a xor b);
    layer2_outputs(10659) <= a and b;
    layer2_outputs(10660) <= not (a xor b);
    layer2_outputs(10661) <= not a or b;
    layer2_outputs(10662) <= not b;
    layer2_outputs(10663) <= not b or a;
    layer2_outputs(10664) <= not a or b;
    layer2_outputs(10665) <= a;
    layer2_outputs(10666) <= a or b;
    layer2_outputs(10667) <= a and b;
    layer2_outputs(10668) <= a;
    layer2_outputs(10669) <= not (a xor b);
    layer2_outputs(10670) <= not a;
    layer2_outputs(10671) <= 1'b0;
    layer2_outputs(10672) <= a and b;
    layer2_outputs(10673) <= b and not a;
    layer2_outputs(10674) <= a and b;
    layer2_outputs(10675) <= a and b;
    layer2_outputs(10676) <= not (a and b);
    layer2_outputs(10677) <= not b or a;
    layer2_outputs(10678) <= not a;
    layer2_outputs(10679) <= a or b;
    layer2_outputs(10680) <= not b or a;
    layer2_outputs(10681) <= b;
    layer2_outputs(10682) <= not a;
    layer2_outputs(10683) <= a and not b;
    layer2_outputs(10684) <= not b;
    layer2_outputs(10685) <= not a;
    layer2_outputs(10686) <= not a or b;
    layer2_outputs(10687) <= not b;
    layer2_outputs(10688) <= b and not a;
    layer2_outputs(10689) <= not b or a;
    layer2_outputs(10690) <= not (a and b);
    layer2_outputs(10691) <= not b;
    layer2_outputs(10692) <= a;
    layer2_outputs(10693) <= not (a and b);
    layer2_outputs(10694) <= not (a xor b);
    layer2_outputs(10695) <= not a;
    layer2_outputs(10696) <= not (a xor b);
    layer2_outputs(10697) <= b;
    layer2_outputs(10698) <= not (a or b);
    layer2_outputs(10699) <= b;
    layer2_outputs(10700) <= 1'b0;
    layer2_outputs(10701) <= not a or b;
    layer2_outputs(10702) <= b;
    layer2_outputs(10703) <= not a or b;
    layer2_outputs(10704) <= a and b;
    layer2_outputs(10705) <= a or b;
    layer2_outputs(10706) <= a;
    layer2_outputs(10707) <= not a or b;
    layer2_outputs(10708) <= b;
    layer2_outputs(10709) <= b;
    layer2_outputs(10710) <= a and b;
    layer2_outputs(10711) <= not b;
    layer2_outputs(10712) <= b;
    layer2_outputs(10713) <= a and b;
    layer2_outputs(10714) <= not b or a;
    layer2_outputs(10715) <= not b;
    layer2_outputs(10716) <= a xor b;
    layer2_outputs(10717) <= not (a or b);
    layer2_outputs(10718) <= not (a xor b);
    layer2_outputs(10719) <= not a;
    layer2_outputs(10720) <= a or b;
    layer2_outputs(10721) <= a and not b;
    layer2_outputs(10722) <= not (a xor b);
    layer2_outputs(10723) <= a and not b;
    layer2_outputs(10724) <= b;
    layer2_outputs(10725) <= not a;
    layer2_outputs(10726) <= not a;
    layer2_outputs(10727) <= b and not a;
    layer2_outputs(10728) <= not a or b;
    layer2_outputs(10729) <= not b;
    layer2_outputs(10730) <= 1'b0;
    layer2_outputs(10731) <= not (a or b);
    layer2_outputs(10732) <= a and b;
    layer2_outputs(10733) <= not (a and b);
    layer2_outputs(10734) <= not b;
    layer2_outputs(10735) <= not (a and b);
    layer2_outputs(10736) <= not (a xor b);
    layer2_outputs(10737) <= not b or a;
    layer2_outputs(10738) <= not b;
    layer2_outputs(10739) <= not a;
    layer2_outputs(10740) <= b;
    layer2_outputs(10741) <= a;
    layer2_outputs(10742) <= not (a xor b);
    layer2_outputs(10743) <= a xor b;
    layer2_outputs(10744) <= a;
    layer2_outputs(10745) <= b;
    layer2_outputs(10746) <= not (a and b);
    layer2_outputs(10747) <= a or b;
    layer2_outputs(10748) <= a;
    layer2_outputs(10749) <= not b;
    layer2_outputs(10750) <= a and not b;
    layer2_outputs(10751) <= not (a or b);
    layer2_outputs(10752) <= not a;
    layer2_outputs(10753) <= not (a xor b);
    layer2_outputs(10754) <= not a or b;
    layer2_outputs(10755) <= not b or a;
    layer2_outputs(10756) <= not (a xor b);
    layer2_outputs(10757) <= not b;
    layer2_outputs(10758) <= not (a or b);
    layer2_outputs(10759) <= a or b;
    layer2_outputs(10760) <= b;
    layer2_outputs(10761) <= not b or a;
    layer2_outputs(10762) <= a xor b;
    layer2_outputs(10763) <= a and b;
    layer2_outputs(10764) <= b;
    layer2_outputs(10765) <= b;
    layer2_outputs(10766) <= a xor b;
    layer2_outputs(10767) <= not b;
    layer2_outputs(10768) <= a;
    layer2_outputs(10769) <= not b or a;
    layer2_outputs(10770) <= a;
    layer2_outputs(10771) <= b;
    layer2_outputs(10772) <= a;
    layer2_outputs(10773) <= not (a xor b);
    layer2_outputs(10774) <= a;
    layer2_outputs(10775) <= not (a or b);
    layer2_outputs(10776) <= a and b;
    layer2_outputs(10777) <= a;
    layer2_outputs(10778) <= not a;
    layer2_outputs(10779) <= not a;
    layer2_outputs(10780) <= b and not a;
    layer2_outputs(10781) <= not a;
    layer2_outputs(10782) <= not (a or b);
    layer2_outputs(10783) <= not (a xor b);
    layer2_outputs(10784) <= not b;
    layer2_outputs(10785) <= not (a or b);
    layer2_outputs(10786) <= not a;
    layer2_outputs(10787) <= a;
    layer2_outputs(10788) <= not b;
    layer2_outputs(10789) <= not (a xor b);
    layer2_outputs(10790) <= not (a xor b);
    layer2_outputs(10791) <= not b or a;
    layer2_outputs(10792) <= not a;
    layer2_outputs(10793) <= not b;
    layer2_outputs(10794) <= not (a or b);
    layer2_outputs(10795) <= not (a and b);
    layer2_outputs(10796) <= not b or a;
    layer2_outputs(10797) <= not a;
    layer2_outputs(10798) <= not b or a;
    layer2_outputs(10799) <= a;
    layer2_outputs(10800) <= b;
    layer2_outputs(10801) <= a;
    layer2_outputs(10802) <= b;
    layer2_outputs(10803) <= not (a or b);
    layer2_outputs(10804) <= not b;
    layer2_outputs(10805) <= not a or b;
    layer2_outputs(10806) <= b;
    layer2_outputs(10807) <= b and not a;
    layer2_outputs(10808) <= b;
    layer2_outputs(10809) <= not b;
    layer2_outputs(10810) <= b;
    layer2_outputs(10811) <= not (a and b);
    layer2_outputs(10812) <= not (a or b);
    layer2_outputs(10813) <= not a;
    layer2_outputs(10814) <= not b or a;
    layer2_outputs(10815) <= a xor b;
    layer2_outputs(10816) <= a;
    layer2_outputs(10817) <= a;
    layer2_outputs(10818) <= b;
    layer2_outputs(10819) <= not (a and b);
    layer2_outputs(10820) <= not (a xor b);
    layer2_outputs(10821) <= a;
    layer2_outputs(10822) <= not a;
    layer2_outputs(10823) <= b and not a;
    layer2_outputs(10824) <= a xor b;
    layer2_outputs(10825) <= b and not a;
    layer2_outputs(10826) <= not a;
    layer2_outputs(10827) <= not (a xor b);
    layer2_outputs(10828) <= not b;
    layer2_outputs(10829) <= a xor b;
    layer2_outputs(10830) <= a xor b;
    layer2_outputs(10831) <= not a;
    layer2_outputs(10832) <= not (a xor b);
    layer2_outputs(10833) <= not (a xor b);
    layer2_outputs(10834) <= b;
    layer2_outputs(10835) <= not b;
    layer2_outputs(10836) <= a and not b;
    layer2_outputs(10837) <= b and not a;
    layer2_outputs(10838) <= not b;
    layer2_outputs(10839) <= a xor b;
    layer2_outputs(10840) <= not (a and b);
    layer2_outputs(10841) <= not (a and b);
    layer2_outputs(10842) <= a xor b;
    layer2_outputs(10843) <= b;
    layer2_outputs(10844) <= not a or b;
    layer2_outputs(10845) <= b;
    layer2_outputs(10846) <= a and b;
    layer2_outputs(10847) <= a;
    layer2_outputs(10848) <= not (a or b);
    layer2_outputs(10849) <= not a or b;
    layer2_outputs(10850) <= a or b;
    layer2_outputs(10851) <= a xor b;
    layer2_outputs(10852) <= not b;
    layer2_outputs(10853) <= not a;
    layer2_outputs(10854) <= not b;
    layer2_outputs(10855) <= not b or a;
    layer2_outputs(10856) <= a;
    layer2_outputs(10857) <= b;
    layer2_outputs(10858) <= a;
    layer2_outputs(10859) <= b;
    layer2_outputs(10860) <= not b;
    layer2_outputs(10861) <= not (a xor b);
    layer2_outputs(10862) <= not (a xor b);
    layer2_outputs(10863) <= a xor b;
    layer2_outputs(10864) <= not a;
    layer2_outputs(10865) <= not a;
    layer2_outputs(10866) <= not a or b;
    layer2_outputs(10867) <= a;
    layer2_outputs(10868) <= not b;
    layer2_outputs(10869) <= a;
    layer2_outputs(10870) <= not b or a;
    layer2_outputs(10871) <= a and not b;
    layer2_outputs(10872) <= not (a and b);
    layer2_outputs(10873) <= a;
    layer2_outputs(10874) <= a and not b;
    layer2_outputs(10875) <= not (a xor b);
    layer2_outputs(10876) <= not a or b;
    layer2_outputs(10877) <= a xor b;
    layer2_outputs(10878) <= not (a xor b);
    layer2_outputs(10879) <= a;
    layer2_outputs(10880) <= a and b;
    layer2_outputs(10881) <= not (a or b);
    layer2_outputs(10882) <= not (a xor b);
    layer2_outputs(10883) <= not b;
    layer2_outputs(10884) <= not (a xor b);
    layer2_outputs(10885) <= not a;
    layer2_outputs(10886) <= not b;
    layer2_outputs(10887) <= not a;
    layer2_outputs(10888) <= b;
    layer2_outputs(10889) <= not b;
    layer2_outputs(10890) <= a and not b;
    layer2_outputs(10891) <= not a;
    layer2_outputs(10892) <= b;
    layer2_outputs(10893) <= a or b;
    layer2_outputs(10894) <= not a;
    layer2_outputs(10895) <= not a or b;
    layer2_outputs(10896) <= not (a xor b);
    layer2_outputs(10897) <= not (a xor b);
    layer2_outputs(10898) <= not a;
    layer2_outputs(10899) <= b and not a;
    layer2_outputs(10900) <= a or b;
    layer2_outputs(10901) <= not b or a;
    layer2_outputs(10902) <= a and b;
    layer2_outputs(10903) <= a;
    layer2_outputs(10904) <= a and b;
    layer2_outputs(10905) <= a xor b;
    layer2_outputs(10906) <= not (a and b);
    layer2_outputs(10907) <= not b;
    layer2_outputs(10908) <= not (a and b);
    layer2_outputs(10909) <= a and b;
    layer2_outputs(10910) <= not (a or b);
    layer2_outputs(10911) <= not b;
    layer2_outputs(10912) <= not (a or b);
    layer2_outputs(10913) <= not b;
    layer2_outputs(10914) <= a;
    layer2_outputs(10915) <= not (a and b);
    layer2_outputs(10916) <= a and b;
    layer2_outputs(10917) <= not b;
    layer2_outputs(10918) <= not b;
    layer2_outputs(10919) <= not (a and b);
    layer2_outputs(10920) <= not a;
    layer2_outputs(10921) <= b;
    layer2_outputs(10922) <= not a;
    layer2_outputs(10923) <= a xor b;
    layer2_outputs(10924) <= a and not b;
    layer2_outputs(10925) <= not b or a;
    layer2_outputs(10926) <= b and not a;
    layer2_outputs(10927) <= a xor b;
    layer2_outputs(10928) <= a or b;
    layer2_outputs(10929) <= not (a or b);
    layer2_outputs(10930) <= a;
    layer2_outputs(10931) <= b and not a;
    layer2_outputs(10932) <= not a;
    layer2_outputs(10933) <= not (a xor b);
    layer2_outputs(10934) <= 1'b0;
    layer2_outputs(10935) <= not (a and b);
    layer2_outputs(10936) <= not (a or b);
    layer2_outputs(10937) <= a xor b;
    layer2_outputs(10938) <= not (a or b);
    layer2_outputs(10939) <= a;
    layer2_outputs(10940) <= a xor b;
    layer2_outputs(10941) <= not a or b;
    layer2_outputs(10942) <= 1'b1;
    layer2_outputs(10943) <= not (a or b);
    layer2_outputs(10944) <= not a or b;
    layer2_outputs(10945) <= not a;
    layer2_outputs(10946) <= not (a xor b);
    layer2_outputs(10947) <= a xor b;
    layer2_outputs(10948) <= b;
    layer2_outputs(10949) <= a;
    layer2_outputs(10950) <= not (a and b);
    layer2_outputs(10951) <= a xor b;
    layer2_outputs(10952) <= not b;
    layer2_outputs(10953) <= not (a or b);
    layer2_outputs(10954) <= a xor b;
    layer2_outputs(10955) <= not a;
    layer2_outputs(10956) <= a;
    layer2_outputs(10957) <= a and not b;
    layer2_outputs(10958) <= not b;
    layer2_outputs(10959) <= a;
    layer2_outputs(10960) <= b;
    layer2_outputs(10961) <= a xor b;
    layer2_outputs(10962) <= a and b;
    layer2_outputs(10963) <= a xor b;
    layer2_outputs(10964) <= not b;
    layer2_outputs(10965) <= b;
    layer2_outputs(10966) <= a;
    layer2_outputs(10967) <= a;
    layer2_outputs(10968) <= not a;
    layer2_outputs(10969) <= not b;
    layer2_outputs(10970) <= not a;
    layer2_outputs(10971) <= a;
    layer2_outputs(10972) <= a xor b;
    layer2_outputs(10973) <= not b;
    layer2_outputs(10974) <= not (a xor b);
    layer2_outputs(10975) <= a and b;
    layer2_outputs(10976) <= a or b;
    layer2_outputs(10977) <= not (a xor b);
    layer2_outputs(10978) <= not (a xor b);
    layer2_outputs(10979) <= not (a and b);
    layer2_outputs(10980) <= a;
    layer2_outputs(10981) <= not (a xor b);
    layer2_outputs(10982) <= not (a and b);
    layer2_outputs(10983) <= not a;
    layer2_outputs(10984) <= a and not b;
    layer2_outputs(10985) <= not (a xor b);
    layer2_outputs(10986) <= not (a and b);
    layer2_outputs(10987) <= not b or a;
    layer2_outputs(10988) <= a xor b;
    layer2_outputs(10989) <= a xor b;
    layer2_outputs(10990) <= a;
    layer2_outputs(10991) <= not b;
    layer2_outputs(10992) <= not (a or b);
    layer2_outputs(10993) <= not b or a;
    layer2_outputs(10994) <= not (a or b);
    layer2_outputs(10995) <= b and not a;
    layer2_outputs(10996) <= b;
    layer2_outputs(10997) <= not (a xor b);
    layer2_outputs(10998) <= a;
    layer2_outputs(10999) <= b;
    layer2_outputs(11000) <= not (a xor b);
    layer2_outputs(11001) <= not a;
    layer2_outputs(11002) <= not (a xor b);
    layer2_outputs(11003) <= not (a and b);
    layer2_outputs(11004) <= not b;
    layer2_outputs(11005) <= b and not a;
    layer2_outputs(11006) <= b;
    layer2_outputs(11007) <= not (a or b);
    layer2_outputs(11008) <= a xor b;
    layer2_outputs(11009) <= not (a or b);
    layer2_outputs(11010) <= a or b;
    layer2_outputs(11011) <= not (a xor b);
    layer2_outputs(11012) <= a;
    layer2_outputs(11013) <= not (a or b);
    layer2_outputs(11014) <= a and b;
    layer2_outputs(11015) <= b;
    layer2_outputs(11016) <= not a;
    layer2_outputs(11017) <= a and not b;
    layer2_outputs(11018) <= b;
    layer2_outputs(11019) <= not b or a;
    layer2_outputs(11020) <= a;
    layer2_outputs(11021) <= a and b;
    layer2_outputs(11022) <= b;
    layer2_outputs(11023) <= a;
    layer2_outputs(11024) <= not b;
    layer2_outputs(11025) <= not a;
    layer2_outputs(11026) <= a and not b;
    layer2_outputs(11027) <= a and not b;
    layer2_outputs(11028) <= not a or b;
    layer2_outputs(11029) <= b and not a;
    layer2_outputs(11030) <= b and not a;
    layer2_outputs(11031) <= a xor b;
    layer2_outputs(11032) <= a xor b;
    layer2_outputs(11033) <= not a;
    layer2_outputs(11034) <= a;
    layer2_outputs(11035) <= not a or b;
    layer2_outputs(11036) <= b;
    layer2_outputs(11037) <= a;
    layer2_outputs(11038) <= b;
    layer2_outputs(11039) <= b and not a;
    layer2_outputs(11040) <= not a or b;
    layer2_outputs(11041) <= not (a and b);
    layer2_outputs(11042) <= not a;
    layer2_outputs(11043) <= b;
    layer2_outputs(11044) <= a or b;
    layer2_outputs(11045) <= not (a or b);
    layer2_outputs(11046) <= not b or a;
    layer2_outputs(11047) <= a or b;
    layer2_outputs(11048) <= b;
    layer2_outputs(11049) <= b and not a;
    layer2_outputs(11050) <= not a;
    layer2_outputs(11051) <= not (a or b);
    layer2_outputs(11052) <= not b;
    layer2_outputs(11053) <= a or b;
    layer2_outputs(11054) <= not a or b;
    layer2_outputs(11055) <= not b;
    layer2_outputs(11056) <= not a;
    layer2_outputs(11057) <= not (a and b);
    layer2_outputs(11058) <= not (a and b);
    layer2_outputs(11059) <= not (a and b);
    layer2_outputs(11060) <= not b or a;
    layer2_outputs(11061) <= b;
    layer2_outputs(11062) <= not b;
    layer2_outputs(11063) <= a;
    layer2_outputs(11064) <= not b;
    layer2_outputs(11065) <= a xor b;
    layer2_outputs(11066) <= not b or a;
    layer2_outputs(11067) <= a or b;
    layer2_outputs(11068) <= not a or b;
    layer2_outputs(11069) <= a;
    layer2_outputs(11070) <= a or b;
    layer2_outputs(11071) <= not (a xor b);
    layer2_outputs(11072) <= a and b;
    layer2_outputs(11073) <= not (a or b);
    layer2_outputs(11074) <= b;
    layer2_outputs(11075) <= 1'b0;
    layer2_outputs(11076) <= not b;
    layer2_outputs(11077) <= not b;
    layer2_outputs(11078) <= not b;
    layer2_outputs(11079) <= 1'b1;
    layer2_outputs(11080) <= b and not a;
    layer2_outputs(11081) <= a or b;
    layer2_outputs(11082) <= a xor b;
    layer2_outputs(11083) <= not b or a;
    layer2_outputs(11084) <= a or b;
    layer2_outputs(11085) <= not b;
    layer2_outputs(11086) <= b and not a;
    layer2_outputs(11087) <= not a;
    layer2_outputs(11088) <= a and not b;
    layer2_outputs(11089) <= not a;
    layer2_outputs(11090) <= not a or b;
    layer2_outputs(11091) <= not (a xor b);
    layer2_outputs(11092) <= b;
    layer2_outputs(11093) <= a xor b;
    layer2_outputs(11094) <= a;
    layer2_outputs(11095) <= not (a and b);
    layer2_outputs(11096) <= a xor b;
    layer2_outputs(11097) <= a;
    layer2_outputs(11098) <= not a;
    layer2_outputs(11099) <= not (a and b);
    layer2_outputs(11100) <= a and not b;
    layer2_outputs(11101) <= not a;
    layer2_outputs(11102) <= a;
    layer2_outputs(11103) <= a or b;
    layer2_outputs(11104) <= not a;
    layer2_outputs(11105) <= a or b;
    layer2_outputs(11106) <= a;
    layer2_outputs(11107) <= b;
    layer2_outputs(11108) <= a;
    layer2_outputs(11109) <= not (a xor b);
    layer2_outputs(11110) <= a and b;
    layer2_outputs(11111) <= b;
    layer2_outputs(11112) <= b and not a;
    layer2_outputs(11113) <= not a;
    layer2_outputs(11114) <= b;
    layer2_outputs(11115) <= a and not b;
    layer2_outputs(11116) <= not b;
    layer2_outputs(11117) <= not (a or b);
    layer2_outputs(11118) <= not (a and b);
    layer2_outputs(11119) <= b;
    layer2_outputs(11120) <= not b;
    layer2_outputs(11121) <= not a;
    layer2_outputs(11122) <= not (a or b);
    layer2_outputs(11123) <= a;
    layer2_outputs(11124) <= not (a or b);
    layer2_outputs(11125) <= not (a xor b);
    layer2_outputs(11126) <= b;
    layer2_outputs(11127) <= a or b;
    layer2_outputs(11128) <= not (a xor b);
    layer2_outputs(11129) <= not a or b;
    layer2_outputs(11130) <= not b;
    layer2_outputs(11131) <= not a;
    layer2_outputs(11132) <= a;
    layer2_outputs(11133) <= a and not b;
    layer2_outputs(11134) <= b;
    layer2_outputs(11135) <= not b or a;
    layer2_outputs(11136) <= b;
    layer2_outputs(11137) <= not a;
    layer2_outputs(11138) <= not (a xor b);
    layer2_outputs(11139) <= a xor b;
    layer2_outputs(11140) <= not b;
    layer2_outputs(11141) <= b;
    layer2_outputs(11142) <= not b;
    layer2_outputs(11143) <= not (a or b);
    layer2_outputs(11144) <= a;
    layer2_outputs(11145) <= a xor b;
    layer2_outputs(11146) <= not a or b;
    layer2_outputs(11147) <= a and not b;
    layer2_outputs(11148) <= not a;
    layer2_outputs(11149) <= a;
    layer2_outputs(11150) <= not a;
    layer2_outputs(11151) <= not a;
    layer2_outputs(11152) <= a xor b;
    layer2_outputs(11153) <= b;
    layer2_outputs(11154) <= not b;
    layer2_outputs(11155) <= b;
    layer2_outputs(11156) <= not (a xor b);
    layer2_outputs(11157) <= a xor b;
    layer2_outputs(11158) <= not (a xor b);
    layer2_outputs(11159) <= a;
    layer2_outputs(11160) <= not (a xor b);
    layer2_outputs(11161) <= a xor b;
    layer2_outputs(11162) <= b;
    layer2_outputs(11163) <= b and not a;
    layer2_outputs(11164) <= not (a or b);
    layer2_outputs(11165) <= b;
    layer2_outputs(11166) <= a and b;
    layer2_outputs(11167) <= a and b;
    layer2_outputs(11168) <= not (a xor b);
    layer2_outputs(11169) <= a xor b;
    layer2_outputs(11170) <= a xor b;
    layer2_outputs(11171) <= a;
    layer2_outputs(11172) <= not (a xor b);
    layer2_outputs(11173) <= a or b;
    layer2_outputs(11174) <= not a;
    layer2_outputs(11175) <= not a;
    layer2_outputs(11176) <= not b;
    layer2_outputs(11177) <= not a;
    layer2_outputs(11178) <= not b;
    layer2_outputs(11179) <= not b;
    layer2_outputs(11180) <= not a or b;
    layer2_outputs(11181) <= a or b;
    layer2_outputs(11182) <= not b;
    layer2_outputs(11183) <= b;
    layer2_outputs(11184) <= a and not b;
    layer2_outputs(11185) <= a and not b;
    layer2_outputs(11186) <= a;
    layer2_outputs(11187) <= b;
    layer2_outputs(11188) <= not a or b;
    layer2_outputs(11189) <= a or b;
    layer2_outputs(11190) <= not (a xor b);
    layer2_outputs(11191) <= a and b;
    layer2_outputs(11192) <= not (a and b);
    layer2_outputs(11193) <= a;
    layer2_outputs(11194) <= a xor b;
    layer2_outputs(11195) <= not b;
    layer2_outputs(11196) <= a xor b;
    layer2_outputs(11197) <= b;
    layer2_outputs(11198) <= not (a xor b);
    layer2_outputs(11199) <= not (a or b);
    layer2_outputs(11200) <= a or b;
    layer2_outputs(11201) <= not (a and b);
    layer2_outputs(11202) <= a and b;
    layer2_outputs(11203) <= not (a xor b);
    layer2_outputs(11204) <= not b or a;
    layer2_outputs(11205) <= not (a or b);
    layer2_outputs(11206) <= not (a xor b);
    layer2_outputs(11207) <= not (a and b);
    layer2_outputs(11208) <= b and not a;
    layer2_outputs(11209) <= b and not a;
    layer2_outputs(11210) <= not a;
    layer2_outputs(11211) <= a or b;
    layer2_outputs(11212) <= a xor b;
    layer2_outputs(11213) <= a xor b;
    layer2_outputs(11214) <= not b;
    layer2_outputs(11215) <= b;
    layer2_outputs(11216) <= a or b;
    layer2_outputs(11217) <= a xor b;
    layer2_outputs(11218) <= a xor b;
    layer2_outputs(11219) <= not (a xor b);
    layer2_outputs(11220) <= not a or b;
    layer2_outputs(11221) <= not a;
    layer2_outputs(11222) <= a or b;
    layer2_outputs(11223) <= not (a and b);
    layer2_outputs(11224) <= a xor b;
    layer2_outputs(11225) <= a;
    layer2_outputs(11226) <= not a;
    layer2_outputs(11227) <= a and b;
    layer2_outputs(11228) <= b;
    layer2_outputs(11229) <= b;
    layer2_outputs(11230) <= a and not b;
    layer2_outputs(11231) <= not a;
    layer2_outputs(11232) <= not b;
    layer2_outputs(11233) <= not b;
    layer2_outputs(11234) <= a and b;
    layer2_outputs(11235) <= a xor b;
    layer2_outputs(11236) <= a xor b;
    layer2_outputs(11237) <= a;
    layer2_outputs(11238) <= not (a xor b);
    layer2_outputs(11239) <= a;
    layer2_outputs(11240) <= b;
    layer2_outputs(11241) <= a xor b;
    layer2_outputs(11242) <= b;
    layer2_outputs(11243) <= a xor b;
    layer2_outputs(11244) <= not (a and b);
    layer2_outputs(11245) <= not b;
    layer2_outputs(11246) <= a;
    layer2_outputs(11247) <= a or b;
    layer2_outputs(11248) <= a;
    layer2_outputs(11249) <= not b;
    layer2_outputs(11250) <= b;
    layer2_outputs(11251) <= not a or b;
    layer2_outputs(11252) <= not (a xor b);
    layer2_outputs(11253) <= b and not a;
    layer2_outputs(11254) <= a or b;
    layer2_outputs(11255) <= a xor b;
    layer2_outputs(11256) <= b;
    layer2_outputs(11257) <= not a or b;
    layer2_outputs(11258) <= a;
    layer2_outputs(11259) <= a xor b;
    layer2_outputs(11260) <= not (a xor b);
    layer2_outputs(11261) <= a;
    layer2_outputs(11262) <= b;
    layer2_outputs(11263) <= not b or a;
    layer2_outputs(11264) <= not b or a;
    layer2_outputs(11265) <= a and b;
    layer2_outputs(11266) <= not (a or b);
    layer2_outputs(11267) <= a and not b;
    layer2_outputs(11268) <= b;
    layer2_outputs(11269) <= a;
    layer2_outputs(11270) <= not (a xor b);
    layer2_outputs(11271) <= not b;
    layer2_outputs(11272) <= not (a or b);
    layer2_outputs(11273) <= b;
    layer2_outputs(11274) <= a xor b;
    layer2_outputs(11275) <= not a;
    layer2_outputs(11276) <= a xor b;
    layer2_outputs(11277) <= a or b;
    layer2_outputs(11278) <= b;
    layer2_outputs(11279) <= b;
    layer2_outputs(11280) <= a and not b;
    layer2_outputs(11281) <= b;
    layer2_outputs(11282) <= not (a or b);
    layer2_outputs(11283) <= a;
    layer2_outputs(11284) <= not (a and b);
    layer2_outputs(11285) <= not a;
    layer2_outputs(11286) <= a;
    layer2_outputs(11287) <= a xor b;
    layer2_outputs(11288) <= not b;
    layer2_outputs(11289) <= a and not b;
    layer2_outputs(11290) <= b;
    layer2_outputs(11291) <= not a or b;
    layer2_outputs(11292) <= a;
    layer2_outputs(11293) <= a xor b;
    layer2_outputs(11294) <= not (a and b);
    layer2_outputs(11295) <= a or b;
    layer2_outputs(11296) <= not a;
    layer2_outputs(11297) <= b;
    layer2_outputs(11298) <= a or b;
    layer2_outputs(11299) <= a and b;
    layer2_outputs(11300) <= not a;
    layer2_outputs(11301) <= not a or b;
    layer2_outputs(11302) <= not b or a;
    layer2_outputs(11303) <= a xor b;
    layer2_outputs(11304) <= a;
    layer2_outputs(11305) <= not a;
    layer2_outputs(11306) <= b and not a;
    layer2_outputs(11307) <= a and not b;
    layer2_outputs(11308) <= not b or a;
    layer2_outputs(11309) <= not b;
    layer2_outputs(11310) <= a;
    layer2_outputs(11311) <= a and b;
    layer2_outputs(11312) <= not b;
    layer2_outputs(11313) <= not (a xor b);
    layer2_outputs(11314) <= a or b;
    layer2_outputs(11315) <= b;
    layer2_outputs(11316) <= a and b;
    layer2_outputs(11317) <= not (a and b);
    layer2_outputs(11318) <= a xor b;
    layer2_outputs(11319) <= not a;
    layer2_outputs(11320) <= not (a and b);
    layer2_outputs(11321) <= not (a and b);
    layer2_outputs(11322) <= a;
    layer2_outputs(11323) <= not (a xor b);
    layer2_outputs(11324) <= not a or b;
    layer2_outputs(11325) <= not b;
    layer2_outputs(11326) <= a or b;
    layer2_outputs(11327) <= a and not b;
    layer2_outputs(11328) <= not a;
    layer2_outputs(11329) <= a;
    layer2_outputs(11330) <= not a;
    layer2_outputs(11331) <= a or b;
    layer2_outputs(11332) <= not (a and b);
    layer2_outputs(11333) <= b;
    layer2_outputs(11334) <= not a or b;
    layer2_outputs(11335) <= b;
    layer2_outputs(11336) <= b and not a;
    layer2_outputs(11337) <= a and not b;
    layer2_outputs(11338) <= a and b;
    layer2_outputs(11339) <= not (a xor b);
    layer2_outputs(11340) <= a xor b;
    layer2_outputs(11341) <= a;
    layer2_outputs(11342) <= a and b;
    layer2_outputs(11343) <= not b;
    layer2_outputs(11344) <= a and not b;
    layer2_outputs(11345) <= not (a xor b);
    layer2_outputs(11346) <= a xor b;
    layer2_outputs(11347) <= not a or b;
    layer2_outputs(11348) <= a and not b;
    layer2_outputs(11349) <= not b;
    layer2_outputs(11350) <= a;
    layer2_outputs(11351) <= a and b;
    layer2_outputs(11352) <= not (a xor b);
    layer2_outputs(11353) <= not a or b;
    layer2_outputs(11354) <= b and not a;
    layer2_outputs(11355) <= not b;
    layer2_outputs(11356) <= b and not a;
    layer2_outputs(11357) <= a;
    layer2_outputs(11358) <= b;
    layer2_outputs(11359) <= a xor b;
    layer2_outputs(11360) <= b;
    layer2_outputs(11361) <= a and not b;
    layer2_outputs(11362) <= b;
    layer2_outputs(11363) <= a and b;
    layer2_outputs(11364) <= a or b;
    layer2_outputs(11365) <= not (a and b);
    layer2_outputs(11366) <= a and not b;
    layer2_outputs(11367) <= a xor b;
    layer2_outputs(11368) <= not a;
    layer2_outputs(11369) <= a;
    layer2_outputs(11370) <= a;
    layer2_outputs(11371) <= not (a xor b);
    layer2_outputs(11372) <= a;
    layer2_outputs(11373) <= not b;
    layer2_outputs(11374) <= not b or a;
    layer2_outputs(11375) <= a or b;
    layer2_outputs(11376) <= not a or b;
    layer2_outputs(11377) <= not a or b;
    layer2_outputs(11378) <= not (a xor b);
    layer2_outputs(11379) <= not (a xor b);
    layer2_outputs(11380) <= not b;
    layer2_outputs(11381) <= a;
    layer2_outputs(11382) <= not (a or b);
    layer2_outputs(11383) <= a;
    layer2_outputs(11384) <= a;
    layer2_outputs(11385) <= a or b;
    layer2_outputs(11386) <= a xor b;
    layer2_outputs(11387) <= a and not b;
    layer2_outputs(11388) <= not (a and b);
    layer2_outputs(11389) <= b;
    layer2_outputs(11390) <= not b;
    layer2_outputs(11391) <= b;
    layer2_outputs(11392) <= not a;
    layer2_outputs(11393) <= not a or b;
    layer2_outputs(11394) <= b and not a;
    layer2_outputs(11395) <= b and not a;
    layer2_outputs(11396) <= not (a or b);
    layer2_outputs(11397) <= b and not a;
    layer2_outputs(11398) <= a;
    layer2_outputs(11399) <= a;
    layer2_outputs(11400) <= not (a and b);
    layer2_outputs(11401) <= not (a xor b);
    layer2_outputs(11402) <= not (a xor b);
    layer2_outputs(11403) <= not a or b;
    layer2_outputs(11404) <= not (a xor b);
    layer2_outputs(11405) <= a and not b;
    layer2_outputs(11406) <= not b;
    layer2_outputs(11407) <= not a;
    layer2_outputs(11408) <= b and not a;
    layer2_outputs(11409) <= b;
    layer2_outputs(11410) <= not (a and b);
    layer2_outputs(11411) <= not a;
    layer2_outputs(11412) <= a;
    layer2_outputs(11413) <= not (a or b);
    layer2_outputs(11414) <= not b;
    layer2_outputs(11415) <= not b;
    layer2_outputs(11416) <= not b;
    layer2_outputs(11417) <= not (a or b);
    layer2_outputs(11418) <= a and not b;
    layer2_outputs(11419) <= 1'b0;
    layer2_outputs(11420) <= not a;
    layer2_outputs(11421) <= not (a and b);
    layer2_outputs(11422) <= a;
    layer2_outputs(11423) <= not b or a;
    layer2_outputs(11424) <= not a;
    layer2_outputs(11425) <= not a or b;
    layer2_outputs(11426) <= b and not a;
    layer2_outputs(11427) <= b;
    layer2_outputs(11428) <= a and not b;
    layer2_outputs(11429) <= a;
    layer2_outputs(11430) <= not a;
    layer2_outputs(11431) <= not b or a;
    layer2_outputs(11432) <= b;
    layer2_outputs(11433) <= not a;
    layer2_outputs(11434) <= not (a or b);
    layer2_outputs(11435) <= b;
    layer2_outputs(11436) <= a xor b;
    layer2_outputs(11437) <= a and b;
    layer2_outputs(11438) <= b;
    layer2_outputs(11439) <= not b;
    layer2_outputs(11440) <= not b;
    layer2_outputs(11441) <= not b;
    layer2_outputs(11442) <= not (a and b);
    layer2_outputs(11443) <= not b;
    layer2_outputs(11444) <= not a;
    layer2_outputs(11445) <= not (a xor b);
    layer2_outputs(11446) <= b and not a;
    layer2_outputs(11447) <= a and not b;
    layer2_outputs(11448) <= a and b;
    layer2_outputs(11449) <= not a;
    layer2_outputs(11450) <= a xor b;
    layer2_outputs(11451) <= a;
    layer2_outputs(11452) <= not (a xor b);
    layer2_outputs(11453) <= a xor b;
    layer2_outputs(11454) <= a xor b;
    layer2_outputs(11455) <= b;
    layer2_outputs(11456) <= not a or b;
    layer2_outputs(11457) <= not b;
    layer2_outputs(11458) <= a or b;
    layer2_outputs(11459) <= not (a and b);
    layer2_outputs(11460) <= b;
    layer2_outputs(11461) <= a xor b;
    layer2_outputs(11462) <= b;
    layer2_outputs(11463) <= a;
    layer2_outputs(11464) <= b and not a;
    layer2_outputs(11465) <= a and not b;
    layer2_outputs(11466) <= not b;
    layer2_outputs(11467) <= not b;
    layer2_outputs(11468) <= not b;
    layer2_outputs(11469) <= not (a xor b);
    layer2_outputs(11470) <= a and b;
    layer2_outputs(11471) <= a;
    layer2_outputs(11472) <= not (a xor b);
    layer2_outputs(11473) <= a and b;
    layer2_outputs(11474) <= not b;
    layer2_outputs(11475) <= a or b;
    layer2_outputs(11476) <= not b or a;
    layer2_outputs(11477) <= not (a or b);
    layer2_outputs(11478) <= not b;
    layer2_outputs(11479) <= a or b;
    layer2_outputs(11480) <= not a or b;
    layer2_outputs(11481) <= a;
    layer2_outputs(11482) <= a;
    layer2_outputs(11483) <= not b or a;
    layer2_outputs(11484) <= a;
    layer2_outputs(11485) <= not (a or b);
    layer2_outputs(11486) <= not b;
    layer2_outputs(11487) <= a and b;
    layer2_outputs(11488) <= not b or a;
    layer2_outputs(11489) <= a and not b;
    layer2_outputs(11490) <= a;
    layer2_outputs(11491) <= not b or a;
    layer2_outputs(11492) <= a xor b;
    layer2_outputs(11493) <= not (a and b);
    layer2_outputs(11494) <= not a;
    layer2_outputs(11495) <= a xor b;
    layer2_outputs(11496) <= not b;
    layer2_outputs(11497) <= not (a or b);
    layer2_outputs(11498) <= a or b;
    layer2_outputs(11499) <= a;
    layer2_outputs(11500) <= not (a xor b);
    layer2_outputs(11501) <= not b or a;
    layer2_outputs(11502) <= not b;
    layer2_outputs(11503) <= a xor b;
    layer2_outputs(11504) <= b;
    layer2_outputs(11505) <= a;
    layer2_outputs(11506) <= not (a or b);
    layer2_outputs(11507) <= a and b;
    layer2_outputs(11508) <= a xor b;
    layer2_outputs(11509) <= 1'b1;
    layer2_outputs(11510) <= not b;
    layer2_outputs(11511) <= not a or b;
    layer2_outputs(11512) <= a xor b;
    layer2_outputs(11513) <= not (a xor b);
    layer2_outputs(11514) <= not b or a;
    layer2_outputs(11515) <= b;
    layer2_outputs(11516) <= b;
    layer2_outputs(11517) <= not b;
    layer2_outputs(11518) <= not a;
    layer2_outputs(11519) <= 1'b1;
    layer2_outputs(11520) <= not b;
    layer2_outputs(11521) <= b;
    layer2_outputs(11522) <= not a;
    layer2_outputs(11523) <= a and not b;
    layer2_outputs(11524) <= not b;
    layer2_outputs(11525) <= not (a or b);
    layer2_outputs(11526) <= a;
    layer2_outputs(11527) <= not a;
    layer2_outputs(11528) <= a and b;
    layer2_outputs(11529) <= not b;
    layer2_outputs(11530) <= not b or a;
    layer2_outputs(11531) <= not (a xor b);
    layer2_outputs(11532) <= b;
    layer2_outputs(11533) <= not a;
    layer2_outputs(11534) <= not (a and b);
    layer2_outputs(11535) <= not a;
    layer2_outputs(11536) <= not (a xor b);
    layer2_outputs(11537) <= b;
    layer2_outputs(11538) <= a and not b;
    layer2_outputs(11539) <= a;
    layer2_outputs(11540) <= not b or a;
    layer2_outputs(11541) <= b and not a;
    layer2_outputs(11542) <= b;
    layer2_outputs(11543) <= not (a and b);
    layer2_outputs(11544) <= not (a and b);
    layer2_outputs(11545) <= a and not b;
    layer2_outputs(11546) <= b;
    layer2_outputs(11547) <= not b;
    layer2_outputs(11548) <= not b;
    layer2_outputs(11549) <= 1'b0;
    layer2_outputs(11550) <= not b or a;
    layer2_outputs(11551) <= b;
    layer2_outputs(11552) <= a xor b;
    layer2_outputs(11553) <= a xor b;
    layer2_outputs(11554) <= a xor b;
    layer2_outputs(11555) <= a or b;
    layer2_outputs(11556) <= not b;
    layer2_outputs(11557) <= a xor b;
    layer2_outputs(11558) <= b and not a;
    layer2_outputs(11559) <= not (a xor b);
    layer2_outputs(11560) <= a xor b;
    layer2_outputs(11561) <= not a;
    layer2_outputs(11562) <= a xor b;
    layer2_outputs(11563) <= not (a and b);
    layer2_outputs(11564) <= a and b;
    layer2_outputs(11565) <= a;
    layer2_outputs(11566) <= b and not a;
    layer2_outputs(11567) <= not (a xor b);
    layer2_outputs(11568) <= not b;
    layer2_outputs(11569) <= not b;
    layer2_outputs(11570) <= a;
    layer2_outputs(11571) <= not (a xor b);
    layer2_outputs(11572) <= a xor b;
    layer2_outputs(11573) <= not b;
    layer2_outputs(11574) <= b;
    layer2_outputs(11575) <= not b;
    layer2_outputs(11576) <= not b;
    layer2_outputs(11577) <= a xor b;
    layer2_outputs(11578) <= not a;
    layer2_outputs(11579) <= a or b;
    layer2_outputs(11580) <= a;
    layer2_outputs(11581) <= a;
    layer2_outputs(11582) <= not b;
    layer2_outputs(11583) <= a or b;
    layer2_outputs(11584) <= a;
    layer2_outputs(11585) <= not b;
    layer2_outputs(11586) <= not b;
    layer2_outputs(11587) <= not a;
    layer2_outputs(11588) <= a and not b;
    layer2_outputs(11589) <= a xor b;
    layer2_outputs(11590) <= 1'b0;
    layer2_outputs(11591) <= not b or a;
    layer2_outputs(11592) <= a xor b;
    layer2_outputs(11593) <= not a;
    layer2_outputs(11594) <= not (a and b);
    layer2_outputs(11595) <= not (a and b);
    layer2_outputs(11596) <= not b;
    layer2_outputs(11597) <= not (a and b);
    layer2_outputs(11598) <= not (a xor b);
    layer2_outputs(11599) <= a xor b;
    layer2_outputs(11600) <= a;
    layer2_outputs(11601) <= not b;
    layer2_outputs(11602) <= b;
    layer2_outputs(11603) <= not b;
    layer2_outputs(11604) <= not (a and b);
    layer2_outputs(11605) <= not (a and b);
    layer2_outputs(11606) <= not b;
    layer2_outputs(11607) <= a xor b;
    layer2_outputs(11608) <= not a or b;
    layer2_outputs(11609) <= a and b;
    layer2_outputs(11610) <= a xor b;
    layer2_outputs(11611) <= not (a xor b);
    layer2_outputs(11612) <= not (a or b);
    layer2_outputs(11613) <= a and b;
    layer2_outputs(11614) <= a and b;
    layer2_outputs(11615) <= not (a and b);
    layer2_outputs(11616) <= a;
    layer2_outputs(11617) <= a and not b;
    layer2_outputs(11618) <= not (a xor b);
    layer2_outputs(11619) <= a and b;
    layer2_outputs(11620) <= not (a xor b);
    layer2_outputs(11621) <= not (a or b);
    layer2_outputs(11622) <= not a;
    layer2_outputs(11623) <= a xor b;
    layer2_outputs(11624) <= not (a or b);
    layer2_outputs(11625) <= not b;
    layer2_outputs(11626) <= a xor b;
    layer2_outputs(11627) <= not (a xor b);
    layer2_outputs(11628) <= not (a xor b);
    layer2_outputs(11629) <= not a;
    layer2_outputs(11630) <= not (a xor b);
    layer2_outputs(11631) <= a xor b;
    layer2_outputs(11632) <= b;
    layer2_outputs(11633) <= not b;
    layer2_outputs(11634) <= not (a xor b);
    layer2_outputs(11635) <= not (a xor b);
    layer2_outputs(11636) <= a xor b;
    layer2_outputs(11637) <= not b;
    layer2_outputs(11638) <= b and not a;
    layer2_outputs(11639) <= not a;
    layer2_outputs(11640) <= a;
    layer2_outputs(11641) <= a;
    layer2_outputs(11642) <= b and not a;
    layer2_outputs(11643) <= not (a or b);
    layer2_outputs(11644) <= a;
    layer2_outputs(11645) <= b and not a;
    layer2_outputs(11646) <= a;
    layer2_outputs(11647) <= a and b;
    layer2_outputs(11648) <= b and not a;
    layer2_outputs(11649) <= b;
    layer2_outputs(11650) <= a;
    layer2_outputs(11651) <= a;
    layer2_outputs(11652) <= not b;
    layer2_outputs(11653) <= not (a or b);
    layer2_outputs(11654) <= not (a or b);
    layer2_outputs(11655) <= b;
    layer2_outputs(11656) <= not b;
    layer2_outputs(11657) <= a xor b;
    layer2_outputs(11658) <= not (a xor b);
    layer2_outputs(11659) <= b;
    layer2_outputs(11660) <= not a or b;
    layer2_outputs(11661) <= not a;
    layer2_outputs(11662) <= a or b;
    layer2_outputs(11663) <= not (a xor b);
    layer2_outputs(11664) <= not b or a;
    layer2_outputs(11665) <= b;
    layer2_outputs(11666) <= not (a xor b);
    layer2_outputs(11667) <= a;
    layer2_outputs(11668) <= not b;
    layer2_outputs(11669) <= not b;
    layer2_outputs(11670) <= a xor b;
    layer2_outputs(11671) <= b;
    layer2_outputs(11672) <= a;
    layer2_outputs(11673) <= a and b;
    layer2_outputs(11674) <= a and b;
    layer2_outputs(11675) <= a or b;
    layer2_outputs(11676) <= not (a xor b);
    layer2_outputs(11677) <= not b or a;
    layer2_outputs(11678) <= a;
    layer2_outputs(11679) <= b;
    layer2_outputs(11680) <= a or b;
    layer2_outputs(11681) <= not b;
    layer2_outputs(11682) <= a;
    layer2_outputs(11683) <= a;
    layer2_outputs(11684) <= not b;
    layer2_outputs(11685) <= a xor b;
    layer2_outputs(11686) <= not (a or b);
    layer2_outputs(11687) <= b;
    layer2_outputs(11688) <= a;
    layer2_outputs(11689) <= a and not b;
    layer2_outputs(11690) <= a;
    layer2_outputs(11691) <= not b;
    layer2_outputs(11692) <= a and b;
    layer2_outputs(11693) <= a;
    layer2_outputs(11694) <= not (a xor b);
    layer2_outputs(11695) <= a or b;
    layer2_outputs(11696) <= not a;
    layer2_outputs(11697) <= b;
    layer2_outputs(11698) <= not b or a;
    layer2_outputs(11699) <= b;
    layer2_outputs(11700) <= not b;
    layer2_outputs(11701) <= a;
    layer2_outputs(11702) <= not a or b;
    layer2_outputs(11703) <= not b or a;
    layer2_outputs(11704) <= b;
    layer2_outputs(11705) <= not a or b;
    layer2_outputs(11706) <= b;
    layer2_outputs(11707) <= a xor b;
    layer2_outputs(11708) <= not b or a;
    layer2_outputs(11709) <= a xor b;
    layer2_outputs(11710) <= not a;
    layer2_outputs(11711) <= a xor b;
    layer2_outputs(11712) <= a xor b;
    layer2_outputs(11713) <= a and not b;
    layer2_outputs(11714) <= b;
    layer2_outputs(11715) <= not a;
    layer2_outputs(11716) <= not a;
    layer2_outputs(11717) <= b and not a;
    layer2_outputs(11718) <= b;
    layer2_outputs(11719) <= a xor b;
    layer2_outputs(11720) <= not (a and b);
    layer2_outputs(11721) <= not a;
    layer2_outputs(11722) <= not b;
    layer2_outputs(11723) <= a and b;
    layer2_outputs(11724) <= not a;
    layer2_outputs(11725) <= not (a or b);
    layer2_outputs(11726) <= not (a xor b);
    layer2_outputs(11727) <= a;
    layer2_outputs(11728) <= a and not b;
    layer2_outputs(11729) <= a xor b;
    layer2_outputs(11730) <= not (a xor b);
    layer2_outputs(11731) <= not b;
    layer2_outputs(11732) <= not b;
    layer2_outputs(11733) <= a;
    layer2_outputs(11734) <= a or b;
    layer2_outputs(11735) <= not (a or b);
    layer2_outputs(11736) <= a;
    layer2_outputs(11737) <= b;
    layer2_outputs(11738) <= not (a and b);
    layer2_outputs(11739) <= not (a and b);
    layer2_outputs(11740) <= not b;
    layer2_outputs(11741) <= not a;
    layer2_outputs(11742) <= a xor b;
    layer2_outputs(11743) <= not a;
    layer2_outputs(11744) <= a and not b;
    layer2_outputs(11745) <= not b or a;
    layer2_outputs(11746) <= not b;
    layer2_outputs(11747) <= not (a xor b);
    layer2_outputs(11748) <= b;
    layer2_outputs(11749) <= not (a xor b);
    layer2_outputs(11750) <= not b or a;
    layer2_outputs(11751) <= not b;
    layer2_outputs(11752) <= b;
    layer2_outputs(11753) <= a;
    layer2_outputs(11754) <= a and not b;
    layer2_outputs(11755) <= not (a xor b);
    layer2_outputs(11756) <= not a;
    layer2_outputs(11757) <= not (a and b);
    layer2_outputs(11758) <= a xor b;
    layer2_outputs(11759) <= not (a or b);
    layer2_outputs(11760) <= not b;
    layer2_outputs(11761) <= b and not a;
    layer2_outputs(11762) <= a xor b;
    layer2_outputs(11763) <= not b;
    layer2_outputs(11764) <= not b;
    layer2_outputs(11765) <= b;
    layer2_outputs(11766) <= not (a xor b);
    layer2_outputs(11767) <= a and b;
    layer2_outputs(11768) <= not (a or b);
    layer2_outputs(11769) <= not (a or b);
    layer2_outputs(11770) <= a or b;
    layer2_outputs(11771) <= 1'b0;
    layer2_outputs(11772) <= a or b;
    layer2_outputs(11773) <= a and b;
    layer2_outputs(11774) <= b;
    layer2_outputs(11775) <= a xor b;
    layer2_outputs(11776) <= not a or b;
    layer2_outputs(11777) <= not (a xor b);
    layer2_outputs(11778) <= not (a xor b);
    layer2_outputs(11779) <= not b or a;
    layer2_outputs(11780) <= a xor b;
    layer2_outputs(11781) <= b;
    layer2_outputs(11782) <= a or b;
    layer2_outputs(11783) <= not a;
    layer2_outputs(11784) <= a and b;
    layer2_outputs(11785) <= not (a xor b);
    layer2_outputs(11786) <= not (a xor b);
    layer2_outputs(11787) <= a xor b;
    layer2_outputs(11788) <= a and b;
    layer2_outputs(11789) <= not (a and b);
    layer2_outputs(11790) <= not a or b;
    layer2_outputs(11791) <= a;
    layer2_outputs(11792) <= a;
    layer2_outputs(11793) <= a;
    layer2_outputs(11794) <= b and not a;
    layer2_outputs(11795) <= b;
    layer2_outputs(11796) <= not a;
    layer2_outputs(11797) <= b;
    layer2_outputs(11798) <= b;
    layer2_outputs(11799) <= a or b;
    layer2_outputs(11800) <= not (a xor b);
    layer2_outputs(11801) <= not (a xor b);
    layer2_outputs(11802) <= not (a and b);
    layer2_outputs(11803) <= not a or b;
    layer2_outputs(11804) <= not (a xor b);
    layer2_outputs(11805) <= not (a or b);
    layer2_outputs(11806) <= not (a and b);
    layer2_outputs(11807) <= a and b;
    layer2_outputs(11808) <= not a;
    layer2_outputs(11809) <= b and not a;
    layer2_outputs(11810) <= a xor b;
    layer2_outputs(11811) <= not (a or b);
    layer2_outputs(11812) <= a;
    layer2_outputs(11813) <= a xor b;
    layer2_outputs(11814) <= b;
    layer2_outputs(11815) <= not b or a;
    layer2_outputs(11816) <= not (a xor b);
    layer2_outputs(11817) <= not (a and b);
    layer2_outputs(11818) <= a xor b;
    layer2_outputs(11819) <= not a;
    layer2_outputs(11820) <= not (a xor b);
    layer2_outputs(11821) <= not a;
    layer2_outputs(11822) <= a;
    layer2_outputs(11823) <= not b or a;
    layer2_outputs(11824) <= not a;
    layer2_outputs(11825) <= not b;
    layer2_outputs(11826) <= not b;
    layer2_outputs(11827) <= a;
    layer2_outputs(11828) <= not (a or b);
    layer2_outputs(11829) <= a and b;
    layer2_outputs(11830) <= a;
    layer2_outputs(11831) <= a or b;
    layer2_outputs(11832) <= not a;
    layer2_outputs(11833) <= a and not b;
    layer2_outputs(11834) <= a and b;
    layer2_outputs(11835) <= b;
    layer2_outputs(11836) <= a and b;
    layer2_outputs(11837) <= a xor b;
    layer2_outputs(11838) <= not (a and b);
    layer2_outputs(11839) <= a or b;
    layer2_outputs(11840) <= not (a xor b);
    layer2_outputs(11841) <= not (a xor b);
    layer2_outputs(11842) <= not (a and b);
    layer2_outputs(11843) <= a xor b;
    layer2_outputs(11844) <= b;
    layer2_outputs(11845) <= a and not b;
    layer2_outputs(11846) <= not b;
    layer2_outputs(11847) <= a xor b;
    layer2_outputs(11848) <= a;
    layer2_outputs(11849) <= not (a and b);
    layer2_outputs(11850) <= not b or a;
    layer2_outputs(11851) <= b;
    layer2_outputs(11852) <= not (a xor b);
    layer2_outputs(11853) <= a;
    layer2_outputs(11854) <= a and not b;
    layer2_outputs(11855) <= not b;
    layer2_outputs(11856) <= a xor b;
    layer2_outputs(11857) <= b and not a;
    layer2_outputs(11858) <= a xor b;
    layer2_outputs(11859) <= a and b;
    layer2_outputs(11860) <= not b or a;
    layer2_outputs(11861) <= not a;
    layer2_outputs(11862) <= a and b;
    layer2_outputs(11863) <= not a;
    layer2_outputs(11864) <= not (a and b);
    layer2_outputs(11865) <= a;
    layer2_outputs(11866) <= a and b;
    layer2_outputs(11867) <= 1'b1;
    layer2_outputs(11868) <= not a;
    layer2_outputs(11869) <= a xor b;
    layer2_outputs(11870) <= not b or a;
    layer2_outputs(11871) <= not (a and b);
    layer2_outputs(11872) <= not (a xor b);
    layer2_outputs(11873) <= b and not a;
    layer2_outputs(11874) <= 1'b1;
    layer2_outputs(11875) <= not (a xor b);
    layer2_outputs(11876) <= b and not a;
    layer2_outputs(11877) <= not (a xor b);
    layer2_outputs(11878) <= a or b;
    layer2_outputs(11879) <= a xor b;
    layer2_outputs(11880) <= b;
    layer2_outputs(11881) <= a and b;
    layer2_outputs(11882) <= not b or a;
    layer2_outputs(11883) <= not a or b;
    layer2_outputs(11884) <= b and not a;
    layer2_outputs(11885) <= not a;
    layer2_outputs(11886) <= a or b;
    layer2_outputs(11887) <= a or b;
    layer2_outputs(11888) <= not a;
    layer2_outputs(11889) <= b and not a;
    layer2_outputs(11890) <= not b or a;
    layer2_outputs(11891) <= a;
    layer2_outputs(11892) <= a and not b;
    layer2_outputs(11893) <= a xor b;
    layer2_outputs(11894) <= a;
    layer2_outputs(11895) <= b;
    layer2_outputs(11896) <= not (a xor b);
    layer2_outputs(11897) <= not a;
    layer2_outputs(11898) <= a xor b;
    layer2_outputs(11899) <= a or b;
    layer2_outputs(11900) <= not a;
    layer2_outputs(11901) <= not a;
    layer2_outputs(11902) <= not (a xor b);
    layer2_outputs(11903) <= not a or b;
    layer2_outputs(11904) <= a and not b;
    layer2_outputs(11905) <= not a or b;
    layer2_outputs(11906) <= not a or b;
    layer2_outputs(11907) <= b;
    layer2_outputs(11908) <= not a or b;
    layer2_outputs(11909) <= a;
    layer2_outputs(11910) <= b and not a;
    layer2_outputs(11911) <= b;
    layer2_outputs(11912) <= a xor b;
    layer2_outputs(11913) <= a or b;
    layer2_outputs(11914) <= not (a and b);
    layer2_outputs(11915) <= a xor b;
    layer2_outputs(11916) <= not a;
    layer2_outputs(11917) <= not (a and b);
    layer2_outputs(11918) <= a;
    layer2_outputs(11919) <= not b;
    layer2_outputs(11920) <= not (a xor b);
    layer2_outputs(11921) <= b;
    layer2_outputs(11922) <= a;
    layer2_outputs(11923) <= not (a xor b);
    layer2_outputs(11924) <= a and b;
    layer2_outputs(11925) <= not (a xor b);
    layer2_outputs(11926) <= a and not b;
    layer2_outputs(11927) <= a or b;
    layer2_outputs(11928) <= not a;
    layer2_outputs(11929) <= not b or a;
    layer2_outputs(11930) <= a or b;
    layer2_outputs(11931) <= not (a xor b);
    layer2_outputs(11932) <= not b;
    layer2_outputs(11933) <= a or b;
    layer2_outputs(11934) <= not (a xor b);
    layer2_outputs(11935) <= a xor b;
    layer2_outputs(11936) <= a and not b;
    layer2_outputs(11937) <= not b or a;
    layer2_outputs(11938) <= b;
    layer2_outputs(11939) <= not (a xor b);
    layer2_outputs(11940) <= a and not b;
    layer2_outputs(11941) <= a xor b;
    layer2_outputs(11942) <= not (a and b);
    layer2_outputs(11943) <= b and not a;
    layer2_outputs(11944) <= a xor b;
    layer2_outputs(11945) <= b and not a;
    layer2_outputs(11946) <= b and not a;
    layer2_outputs(11947) <= b;
    layer2_outputs(11948) <= b;
    layer2_outputs(11949) <= not a;
    layer2_outputs(11950) <= not (a xor b);
    layer2_outputs(11951) <= b;
    layer2_outputs(11952) <= not b;
    layer2_outputs(11953) <= not (a or b);
    layer2_outputs(11954) <= not b;
    layer2_outputs(11955) <= a and b;
    layer2_outputs(11956) <= a xor b;
    layer2_outputs(11957) <= not (a xor b);
    layer2_outputs(11958) <= b and not a;
    layer2_outputs(11959) <= not a or b;
    layer2_outputs(11960) <= b;
    layer2_outputs(11961) <= b and not a;
    layer2_outputs(11962) <= not (a xor b);
    layer2_outputs(11963) <= b;
    layer2_outputs(11964) <= a or b;
    layer2_outputs(11965) <= b and not a;
    layer2_outputs(11966) <= not b;
    layer2_outputs(11967) <= not a;
    layer2_outputs(11968) <= a xor b;
    layer2_outputs(11969) <= a;
    layer2_outputs(11970) <= a xor b;
    layer2_outputs(11971) <= not (a and b);
    layer2_outputs(11972) <= not (a xor b);
    layer2_outputs(11973) <= not (a or b);
    layer2_outputs(11974) <= not b;
    layer2_outputs(11975) <= not a;
    layer2_outputs(11976) <= not a;
    layer2_outputs(11977) <= b;
    layer2_outputs(11978) <= not a;
    layer2_outputs(11979) <= not a;
    layer2_outputs(11980) <= b and not a;
    layer2_outputs(11981) <= a or b;
    layer2_outputs(11982) <= b;
    layer2_outputs(11983) <= b;
    layer2_outputs(11984) <= a;
    layer2_outputs(11985) <= not (a or b);
    layer2_outputs(11986) <= a and b;
    layer2_outputs(11987) <= a xor b;
    layer2_outputs(11988) <= a;
    layer2_outputs(11989) <= a xor b;
    layer2_outputs(11990) <= not b;
    layer2_outputs(11991) <= a xor b;
    layer2_outputs(11992) <= not b;
    layer2_outputs(11993) <= a;
    layer2_outputs(11994) <= not b;
    layer2_outputs(11995) <= not (a or b);
    layer2_outputs(11996) <= not b;
    layer2_outputs(11997) <= a;
    layer2_outputs(11998) <= a;
    layer2_outputs(11999) <= not (a xor b);
    layer2_outputs(12000) <= a;
    layer2_outputs(12001) <= not (a or b);
    layer2_outputs(12002) <= a;
    layer2_outputs(12003) <= a;
    layer2_outputs(12004) <= b and not a;
    layer2_outputs(12005) <= b;
    layer2_outputs(12006) <= 1'b0;
    layer2_outputs(12007) <= a and b;
    layer2_outputs(12008) <= a xor b;
    layer2_outputs(12009) <= a;
    layer2_outputs(12010) <= a or b;
    layer2_outputs(12011) <= not a;
    layer2_outputs(12012) <= a;
    layer2_outputs(12013) <= not b;
    layer2_outputs(12014) <= a xor b;
    layer2_outputs(12015) <= a xor b;
    layer2_outputs(12016) <= a xor b;
    layer2_outputs(12017) <= b;
    layer2_outputs(12018) <= not (a and b);
    layer2_outputs(12019) <= not a;
    layer2_outputs(12020) <= a and b;
    layer2_outputs(12021) <= a;
    layer2_outputs(12022) <= not (a or b);
    layer2_outputs(12023) <= not a;
    layer2_outputs(12024) <= not b;
    layer2_outputs(12025) <= not (a xor b);
    layer2_outputs(12026) <= b;
    layer2_outputs(12027) <= not a or b;
    layer2_outputs(12028) <= not b;
    layer2_outputs(12029) <= not a or b;
    layer2_outputs(12030) <= a;
    layer2_outputs(12031) <= not a or b;
    layer2_outputs(12032) <= a;
    layer2_outputs(12033) <= not (a or b);
    layer2_outputs(12034) <= not b;
    layer2_outputs(12035) <= not a;
    layer2_outputs(12036) <= not a;
    layer2_outputs(12037) <= not a;
    layer2_outputs(12038) <= a xor b;
    layer2_outputs(12039) <= not a or b;
    layer2_outputs(12040) <= not (a xor b);
    layer2_outputs(12041) <= a;
    layer2_outputs(12042) <= not b;
    layer2_outputs(12043) <= b;
    layer2_outputs(12044) <= a;
    layer2_outputs(12045) <= not b or a;
    layer2_outputs(12046) <= a;
    layer2_outputs(12047) <= a or b;
    layer2_outputs(12048) <= not a;
    layer2_outputs(12049) <= not b;
    layer2_outputs(12050) <= a;
    layer2_outputs(12051) <= not (a or b);
    layer2_outputs(12052) <= not a;
    layer2_outputs(12053) <= a xor b;
    layer2_outputs(12054) <= b and not a;
    layer2_outputs(12055) <= not b;
    layer2_outputs(12056) <= a and b;
    layer2_outputs(12057) <= a xor b;
    layer2_outputs(12058) <= a xor b;
    layer2_outputs(12059) <= not b;
    layer2_outputs(12060) <= a xor b;
    layer2_outputs(12061) <= not a or b;
    layer2_outputs(12062) <= a or b;
    layer2_outputs(12063) <= not (a xor b);
    layer2_outputs(12064) <= not b or a;
    layer2_outputs(12065) <= a;
    layer2_outputs(12066) <= not a;
    layer2_outputs(12067) <= a;
    layer2_outputs(12068) <= not (a xor b);
    layer2_outputs(12069) <= not (a xor b);
    layer2_outputs(12070) <= not (a xor b);
    layer2_outputs(12071) <= not a;
    layer2_outputs(12072) <= a;
    layer2_outputs(12073) <= not (a xor b);
    layer2_outputs(12074) <= not b or a;
    layer2_outputs(12075) <= not (a xor b);
    layer2_outputs(12076) <= not b or a;
    layer2_outputs(12077) <= a xor b;
    layer2_outputs(12078) <= not a;
    layer2_outputs(12079) <= a;
    layer2_outputs(12080) <= not (a xor b);
    layer2_outputs(12081) <= not b;
    layer2_outputs(12082) <= b and not a;
    layer2_outputs(12083) <= not b or a;
    layer2_outputs(12084) <= a and b;
    layer2_outputs(12085) <= b;
    layer2_outputs(12086) <= a;
    layer2_outputs(12087) <= not a;
    layer2_outputs(12088) <= not a or b;
    layer2_outputs(12089) <= not a;
    layer2_outputs(12090) <= a;
    layer2_outputs(12091) <= a;
    layer2_outputs(12092) <= b and not a;
    layer2_outputs(12093) <= a;
    layer2_outputs(12094) <= a;
    layer2_outputs(12095) <= a and b;
    layer2_outputs(12096) <= not a;
    layer2_outputs(12097) <= not (a xor b);
    layer2_outputs(12098) <= not b or a;
    layer2_outputs(12099) <= b;
    layer2_outputs(12100) <= not a;
    layer2_outputs(12101) <= not a;
    layer2_outputs(12102) <= a;
    layer2_outputs(12103) <= not b;
    layer2_outputs(12104) <= not (a xor b);
    layer2_outputs(12105) <= not a or b;
    layer2_outputs(12106) <= a;
    layer2_outputs(12107) <= a;
    layer2_outputs(12108) <= b;
    layer2_outputs(12109) <= not (a or b);
    layer2_outputs(12110) <= not (a xor b);
    layer2_outputs(12111) <= a;
    layer2_outputs(12112) <= a or b;
    layer2_outputs(12113) <= not a;
    layer2_outputs(12114) <= a and b;
    layer2_outputs(12115) <= not b or a;
    layer2_outputs(12116) <= a and not b;
    layer2_outputs(12117) <= not b or a;
    layer2_outputs(12118) <= not (a or b);
    layer2_outputs(12119) <= not a;
    layer2_outputs(12120) <= a or b;
    layer2_outputs(12121) <= a or b;
    layer2_outputs(12122) <= a and not b;
    layer2_outputs(12123) <= not (a or b);
    layer2_outputs(12124) <= a or b;
    layer2_outputs(12125) <= not b or a;
    layer2_outputs(12126) <= not b;
    layer2_outputs(12127) <= a and not b;
    layer2_outputs(12128) <= not (a xor b);
    layer2_outputs(12129) <= b and not a;
    layer2_outputs(12130) <= not b or a;
    layer2_outputs(12131) <= not a;
    layer2_outputs(12132) <= b and not a;
    layer2_outputs(12133) <= not a or b;
    layer2_outputs(12134) <= not (a xor b);
    layer2_outputs(12135) <= not b;
    layer2_outputs(12136) <= not b;
    layer2_outputs(12137) <= b;
    layer2_outputs(12138) <= a or b;
    layer2_outputs(12139) <= not a;
    layer2_outputs(12140) <= not a or b;
    layer2_outputs(12141) <= not (a xor b);
    layer2_outputs(12142) <= a xor b;
    layer2_outputs(12143) <= not b;
    layer2_outputs(12144) <= not (a and b);
    layer2_outputs(12145) <= not a or b;
    layer2_outputs(12146) <= not a;
    layer2_outputs(12147) <= not b or a;
    layer2_outputs(12148) <= b;
    layer2_outputs(12149) <= b and not a;
    layer2_outputs(12150) <= a;
    layer2_outputs(12151) <= not b or a;
    layer2_outputs(12152) <= b;
    layer2_outputs(12153) <= not a or b;
    layer2_outputs(12154) <= not (a or b);
    layer2_outputs(12155) <= b;
    layer2_outputs(12156) <= not a or b;
    layer2_outputs(12157) <= b;
    layer2_outputs(12158) <= b and not a;
    layer2_outputs(12159) <= a and not b;
    layer2_outputs(12160) <= b;
    layer2_outputs(12161) <= b;
    layer2_outputs(12162) <= not (a or b);
    layer2_outputs(12163) <= not b;
    layer2_outputs(12164) <= not (a xor b);
    layer2_outputs(12165) <= b;
    layer2_outputs(12166) <= b;
    layer2_outputs(12167) <= a or b;
    layer2_outputs(12168) <= a and b;
    layer2_outputs(12169) <= a and not b;
    layer2_outputs(12170) <= not (a and b);
    layer2_outputs(12171) <= not (a or b);
    layer2_outputs(12172) <= not a;
    layer2_outputs(12173) <= not a;
    layer2_outputs(12174) <= not a or b;
    layer2_outputs(12175) <= not a;
    layer2_outputs(12176) <= a xor b;
    layer2_outputs(12177) <= not (a xor b);
    layer2_outputs(12178) <= b;
    layer2_outputs(12179) <= a and b;
    layer2_outputs(12180) <= b;
    layer2_outputs(12181) <= a xor b;
    layer2_outputs(12182) <= not b or a;
    layer2_outputs(12183) <= a xor b;
    layer2_outputs(12184) <= not b;
    layer2_outputs(12185) <= not a;
    layer2_outputs(12186) <= not a;
    layer2_outputs(12187) <= b and not a;
    layer2_outputs(12188) <= b and not a;
    layer2_outputs(12189) <= not (a xor b);
    layer2_outputs(12190) <= a xor b;
    layer2_outputs(12191) <= not a;
    layer2_outputs(12192) <= a xor b;
    layer2_outputs(12193) <= not b;
    layer2_outputs(12194) <= not (a and b);
    layer2_outputs(12195) <= a or b;
    layer2_outputs(12196) <= not a or b;
    layer2_outputs(12197) <= not a or b;
    layer2_outputs(12198) <= not (a xor b);
    layer2_outputs(12199) <= a and b;
    layer2_outputs(12200) <= not a;
    layer2_outputs(12201) <= a xor b;
    layer2_outputs(12202) <= not a;
    layer2_outputs(12203) <= not a;
    layer2_outputs(12204) <= not (a and b);
    layer2_outputs(12205) <= not (a and b);
    layer2_outputs(12206) <= a and b;
    layer2_outputs(12207) <= a;
    layer2_outputs(12208) <= b;
    layer2_outputs(12209) <= 1'b1;
    layer2_outputs(12210) <= not a;
    layer2_outputs(12211) <= a or b;
    layer2_outputs(12212) <= not a or b;
    layer2_outputs(12213) <= not (a and b);
    layer2_outputs(12214) <= a;
    layer2_outputs(12215) <= not a;
    layer2_outputs(12216) <= b and not a;
    layer2_outputs(12217) <= a and b;
    layer2_outputs(12218) <= b;
    layer2_outputs(12219) <= a xor b;
    layer2_outputs(12220) <= a;
    layer2_outputs(12221) <= not b;
    layer2_outputs(12222) <= a xor b;
    layer2_outputs(12223) <= not a or b;
    layer2_outputs(12224) <= b;
    layer2_outputs(12225) <= a;
    layer2_outputs(12226) <= not (a and b);
    layer2_outputs(12227) <= not (a or b);
    layer2_outputs(12228) <= not (a and b);
    layer2_outputs(12229) <= a and b;
    layer2_outputs(12230) <= b;
    layer2_outputs(12231) <= a;
    layer2_outputs(12232) <= b;
    layer2_outputs(12233) <= not a or b;
    layer2_outputs(12234) <= b and not a;
    layer2_outputs(12235) <= not a;
    layer2_outputs(12236) <= a xor b;
    layer2_outputs(12237) <= not b;
    layer2_outputs(12238) <= not b;
    layer2_outputs(12239) <= not a;
    layer2_outputs(12240) <= a;
    layer2_outputs(12241) <= b;
    layer2_outputs(12242) <= not b;
    layer2_outputs(12243) <= not b or a;
    layer2_outputs(12244) <= a xor b;
    layer2_outputs(12245) <= a xor b;
    layer2_outputs(12246) <= not (a or b);
    layer2_outputs(12247) <= a xor b;
    layer2_outputs(12248) <= a and b;
    layer2_outputs(12249) <= a xor b;
    layer2_outputs(12250) <= not b;
    layer2_outputs(12251) <= a and not b;
    layer2_outputs(12252) <= not b;
    layer2_outputs(12253) <= a or b;
    layer2_outputs(12254) <= b and not a;
    layer2_outputs(12255) <= not (a xor b);
    layer2_outputs(12256) <= not (a or b);
    layer2_outputs(12257) <= a and not b;
    layer2_outputs(12258) <= a xor b;
    layer2_outputs(12259) <= b;
    layer2_outputs(12260) <= not (a and b);
    layer2_outputs(12261) <= not b or a;
    layer2_outputs(12262) <= b;
    layer2_outputs(12263) <= a xor b;
    layer2_outputs(12264) <= not b;
    layer2_outputs(12265) <= a and not b;
    layer2_outputs(12266) <= not b;
    layer2_outputs(12267) <= not a or b;
    layer2_outputs(12268) <= not (a or b);
    layer2_outputs(12269) <= b;
    layer2_outputs(12270) <= not a or b;
    layer2_outputs(12271) <= a xor b;
    layer2_outputs(12272) <= b;
    layer2_outputs(12273) <= a and b;
    layer2_outputs(12274) <= not (a or b);
    layer2_outputs(12275) <= not a;
    layer2_outputs(12276) <= b;
    layer2_outputs(12277) <= not a;
    layer2_outputs(12278) <= a xor b;
    layer2_outputs(12279) <= b;
    layer2_outputs(12280) <= not b;
    layer2_outputs(12281) <= b;
    layer2_outputs(12282) <= b;
    layer2_outputs(12283) <= not a;
    layer2_outputs(12284) <= not a;
    layer2_outputs(12285) <= b;
    layer2_outputs(12286) <= a xor b;
    layer2_outputs(12287) <= not a or b;
    layer2_outputs(12288) <= not (a xor b);
    layer2_outputs(12289) <= b and not a;
    layer2_outputs(12290) <= a and not b;
    layer2_outputs(12291) <= not b;
    layer2_outputs(12292) <= a xor b;
    layer2_outputs(12293) <= not b;
    layer2_outputs(12294) <= not (a xor b);
    layer2_outputs(12295) <= not (a xor b);
    layer2_outputs(12296) <= a and not b;
    layer2_outputs(12297) <= a and not b;
    layer2_outputs(12298) <= not (a and b);
    layer2_outputs(12299) <= b;
    layer2_outputs(12300) <= a and not b;
    layer2_outputs(12301) <= not a;
    layer2_outputs(12302) <= not (a xor b);
    layer2_outputs(12303) <= a and not b;
    layer2_outputs(12304) <= not (a xor b);
    layer2_outputs(12305) <= not b;
    layer2_outputs(12306) <= a and b;
    layer2_outputs(12307) <= not b;
    layer2_outputs(12308) <= not a;
    layer2_outputs(12309) <= a;
    layer2_outputs(12310) <= not (a or b);
    layer2_outputs(12311) <= not (a and b);
    layer2_outputs(12312) <= a and not b;
    layer2_outputs(12313) <= not a;
    layer2_outputs(12314) <= a and not b;
    layer2_outputs(12315) <= a and b;
    layer2_outputs(12316) <= not a;
    layer2_outputs(12317) <= a xor b;
    layer2_outputs(12318) <= not a;
    layer2_outputs(12319) <= a;
    layer2_outputs(12320) <= not b;
    layer2_outputs(12321) <= not a;
    layer2_outputs(12322) <= b;
    layer2_outputs(12323) <= b;
    layer2_outputs(12324) <= not a;
    layer2_outputs(12325) <= a xor b;
    layer2_outputs(12326) <= a;
    layer2_outputs(12327) <= b and not a;
    layer2_outputs(12328) <= not (a or b);
    layer2_outputs(12329) <= a xor b;
    layer2_outputs(12330) <= not (a xor b);
    layer2_outputs(12331) <= not b or a;
    layer2_outputs(12332) <= not (a and b);
    layer2_outputs(12333) <= not a or b;
    layer2_outputs(12334) <= b and not a;
    layer2_outputs(12335) <= b and not a;
    layer2_outputs(12336) <= a or b;
    layer2_outputs(12337) <= a and b;
    layer2_outputs(12338) <= not b;
    layer2_outputs(12339) <= not b or a;
    layer2_outputs(12340) <= b and not a;
    layer2_outputs(12341) <= not a or b;
    layer2_outputs(12342) <= not (a or b);
    layer2_outputs(12343) <= b;
    layer2_outputs(12344) <= b;
    layer2_outputs(12345) <= b;
    layer2_outputs(12346) <= b and not a;
    layer2_outputs(12347) <= not a;
    layer2_outputs(12348) <= a xor b;
    layer2_outputs(12349) <= a and b;
    layer2_outputs(12350) <= a;
    layer2_outputs(12351) <= not b;
    layer2_outputs(12352) <= a xor b;
    layer2_outputs(12353) <= not a;
    layer2_outputs(12354) <= not (a xor b);
    layer2_outputs(12355) <= not a or b;
    layer2_outputs(12356) <= not (a and b);
    layer2_outputs(12357) <= not (a or b);
    layer2_outputs(12358) <= not (a and b);
    layer2_outputs(12359) <= not b;
    layer2_outputs(12360) <= not a;
    layer2_outputs(12361) <= not a;
    layer2_outputs(12362) <= not b or a;
    layer2_outputs(12363) <= a;
    layer2_outputs(12364) <= a or b;
    layer2_outputs(12365) <= b;
    layer2_outputs(12366) <= not a;
    layer2_outputs(12367) <= not b;
    layer2_outputs(12368) <= not b;
    layer2_outputs(12369) <= a;
    layer2_outputs(12370) <= b;
    layer2_outputs(12371) <= not b;
    layer2_outputs(12372) <= b;
    layer2_outputs(12373) <= a;
    layer2_outputs(12374) <= b and not a;
    layer2_outputs(12375) <= not b or a;
    layer2_outputs(12376) <= a;
    layer2_outputs(12377) <= b;
    layer2_outputs(12378) <= not b;
    layer2_outputs(12379) <= not (a xor b);
    layer2_outputs(12380) <= a;
    layer2_outputs(12381) <= not (a or b);
    layer2_outputs(12382) <= not a;
    layer2_outputs(12383) <= not (a xor b);
    layer2_outputs(12384) <= b and not a;
    layer2_outputs(12385) <= a xor b;
    layer2_outputs(12386) <= not (a and b);
    layer2_outputs(12387) <= a xor b;
    layer2_outputs(12388) <= a and not b;
    layer2_outputs(12389) <= a or b;
    layer2_outputs(12390) <= b;
    layer2_outputs(12391) <= not b;
    layer2_outputs(12392) <= b;
    layer2_outputs(12393) <= not b;
    layer2_outputs(12394) <= a xor b;
    layer2_outputs(12395) <= not (a xor b);
    layer2_outputs(12396) <= a xor b;
    layer2_outputs(12397) <= a;
    layer2_outputs(12398) <= not (a xor b);
    layer2_outputs(12399) <= not a;
    layer2_outputs(12400) <= not (a or b);
    layer2_outputs(12401) <= not a;
    layer2_outputs(12402) <= b;
    layer2_outputs(12403) <= not a or b;
    layer2_outputs(12404) <= b and not a;
    layer2_outputs(12405) <= not b or a;
    layer2_outputs(12406) <= not (a and b);
    layer2_outputs(12407) <= not b;
    layer2_outputs(12408) <= a;
    layer2_outputs(12409) <= a;
    layer2_outputs(12410) <= b;
    layer2_outputs(12411) <= not b;
    layer2_outputs(12412) <= a;
    layer2_outputs(12413) <= not b or a;
    layer2_outputs(12414) <= not b;
    layer2_outputs(12415) <= not (a xor b);
    layer2_outputs(12416) <= not a;
    layer2_outputs(12417) <= not (a and b);
    layer2_outputs(12418) <= a and not b;
    layer2_outputs(12419) <= b;
    layer2_outputs(12420) <= a;
    layer2_outputs(12421) <= not (a or b);
    layer2_outputs(12422) <= a;
    layer2_outputs(12423) <= not a;
    layer2_outputs(12424) <= b and not a;
    layer2_outputs(12425) <= b and not a;
    layer2_outputs(12426) <= not b or a;
    layer2_outputs(12427) <= a xor b;
    layer2_outputs(12428) <= a xor b;
    layer2_outputs(12429) <= b;
    layer2_outputs(12430) <= not b;
    layer2_outputs(12431) <= b;
    layer2_outputs(12432) <= a and not b;
    layer2_outputs(12433) <= b;
    layer2_outputs(12434) <= not b;
    layer2_outputs(12435) <= not b;
    layer2_outputs(12436) <= a and b;
    layer2_outputs(12437) <= not (a xor b);
    layer2_outputs(12438) <= not (a xor b);
    layer2_outputs(12439) <= b;
    layer2_outputs(12440) <= a;
    layer2_outputs(12441) <= b;
    layer2_outputs(12442) <= not b or a;
    layer2_outputs(12443) <= not b;
    layer2_outputs(12444) <= not a;
    layer2_outputs(12445) <= not a or b;
    layer2_outputs(12446) <= a xor b;
    layer2_outputs(12447) <= not (a xor b);
    layer2_outputs(12448) <= not a or b;
    layer2_outputs(12449) <= a and not b;
    layer2_outputs(12450) <= not (a or b);
    layer2_outputs(12451) <= not (a or b);
    layer2_outputs(12452) <= not a;
    layer2_outputs(12453) <= not b;
    layer2_outputs(12454) <= b;
    layer2_outputs(12455) <= a and not b;
    layer2_outputs(12456) <= a and b;
    layer2_outputs(12457) <= a;
    layer2_outputs(12458) <= not a;
    layer2_outputs(12459) <= a or b;
    layer2_outputs(12460) <= b and not a;
    layer2_outputs(12461) <= not b;
    layer2_outputs(12462) <= not (a xor b);
    layer2_outputs(12463) <= not (a xor b);
    layer2_outputs(12464) <= not b;
    layer2_outputs(12465) <= a;
    layer2_outputs(12466) <= not b or a;
    layer2_outputs(12467) <= not (a and b);
    layer2_outputs(12468) <= b and not a;
    layer2_outputs(12469) <= not (a and b);
    layer2_outputs(12470) <= not a;
    layer2_outputs(12471) <= a and not b;
    layer2_outputs(12472) <= not a or b;
    layer2_outputs(12473) <= not a or b;
    layer2_outputs(12474) <= a or b;
    layer2_outputs(12475) <= a or b;
    layer2_outputs(12476) <= a and not b;
    layer2_outputs(12477) <= not (a xor b);
    layer2_outputs(12478) <= not (a xor b);
    layer2_outputs(12479) <= not (a xor b);
    layer2_outputs(12480) <= not a;
    layer2_outputs(12481) <= not (a and b);
    layer2_outputs(12482) <= not (a xor b);
    layer2_outputs(12483) <= not (a xor b);
    layer2_outputs(12484) <= not (a xor b);
    layer2_outputs(12485) <= a and not b;
    layer2_outputs(12486) <= not b or a;
    layer2_outputs(12487) <= 1'b0;
    layer2_outputs(12488) <= not a;
    layer2_outputs(12489) <= a;
    layer2_outputs(12490) <= a;
    layer2_outputs(12491) <= not (a xor b);
    layer2_outputs(12492) <= b and not a;
    layer2_outputs(12493) <= not (a xor b);
    layer2_outputs(12494) <= not b;
    layer2_outputs(12495) <= not a;
    layer2_outputs(12496) <= b and not a;
    layer2_outputs(12497) <= a xor b;
    layer2_outputs(12498) <= a xor b;
    layer2_outputs(12499) <= b and not a;
    layer2_outputs(12500) <= a;
    layer2_outputs(12501) <= not a;
    layer2_outputs(12502) <= not b;
    layer2_outputs(12503) <= not a or b;
    layer2_outputs(12504) <= b;
    layer2_outputs(12505) <= a and b;
    layer2_outputs(12506) <= not (a xor b);
    layer2_outputs(12507) <= not b or a;
    layer2_outputs(12508) <= not (a xor b);
    layer2_outputs(12509) <= not b;
    layer2_outputs(12510) <= a and b;
    layer2_outputs(12511) <= b;
    layer2_outputs(12512) <= not a;
    layer2_outputs(12513) <= not a or b;
    layer2_outputs(12514) <= not (a xor b);
    layer2_outputs(12515) <= a or b;
    layer2_outputs(12516) <= not (a or b);
    layer2_outputs(12517) <= a and b;
    layer2_outputs(12518) <= a and not b;
    layer2_outputs(12519) <= a and b;
    layer2_outputs(12520) <= b and not a;
    layer2_outputs(12521) <= not (a and b);
    layer2_outputs(12522) <= not (a and b);
    layer2_outputs(12523) <= not b;
    layer2_outputs(12524) <= not (a xor b);
    layer2_outputs(12525) <= b and not a;
    layer2_outputs(12526) <= a and b;
    layer2_outputs(12527) <= b;
    layer2_outputs(12528) <= b;
    layer2_outputs(12529) <= 1'b0;
    layer2_outputs(12530) <= a xor b;
    layer2_outputs(12531) <= a xor b;
    layer2_outputs(12532) <= a;
    layer2_outputs(12533) <= a xor b;
    layer2_outputs(12534) <= a and b;
    layer2_outputs(12535) <= not a;
    layer2_outputs(12536) <= b;
    layer2_outputs(12537) <= not (a xor b);
    layer2_outputs(12538) <= b;
    layer2_outputs(12539) <= not (a xor b);
    layer2_outputs(12540) <= b;
    layer2_outputs(12541) <= b and not a;
    layer2_outputs(12542) <= not b;
    layer2_outputs(12543) <= not b;
    layer2_outputs(12544) <= a and not b;
    layer2_outputs(12545) <= not (a xor b);
    layer2_outputs(12546) <= a and b;
    layer2_outputs(12547) <= a and not b;
    layer2_outputs(12548) <= a xor b;
    layer2_outputs(12549) <= not b;
    layer2_outputs(12550) <= a;
    layer2_outputs(12551) <= a xor b;
    layer2_outputs(12552) <= not a;
    layer2_outputs(12553) <= not b;
    layer2_outputs(12554) <= a and not b;
    layer2_outputs(12555) <= a and not b;
    layer2_outputs(12556) <= a and b;
    layer2_outputs(12557) <= a and not b;
    layer2_outputs(12558) <= a xor b;
    layer2_outputs(12559) <= not (a and b);
    layer2_outputs(12560) <= a xor b;
    layer2_outputs(12561) <= a;
    layer2_outputs(12562) <= not a or b;
    layer2_outputs(12563) <= b;
    layer2_outputs(12564) <= b;
    layer2_outputs(12565) <= not a;
    layer2_outputs(12566) <= a;
    layer2_outputs(12567) <= a xor b;
    layer2_outputs(12568) <= a or b;
    layer2_outputs(12569) <= not (a xor b);
    layer2_outputs(12570) <= not b;
    layer2_outputs(12571) <= not (a or b);
    layer2_outputs(12572) <= a;
    layer2_outputs(12573) <= not b;
    layer2_outputs(12574) <= not a;
    layer2_outputs(12575) <= not b;
    layer2_outputs(12576) <= b;
    layer2_outputs(12577) <= b and not a;
    layer2_outputs(12578) <= a or b;
    layer2_outputs(12579) <= not (a xor b);
    layer2_outputs(12580) <= a xor b;
    layer2_outputs(12581) <= b;
    layer2_outputs(12582) <= not (a and b);
    layer2_outputs(12583) <= a or b;
    layer2_outputs(12584) <= not b or a;
    layer2_outputs(12585) <= a or b;
    layer2_outputs(12586) <= b and not a;
    layer2_outputs(12587) <= not (a xor b);
    layer2_outputs(12588) <= not a;
    layer2_outputs(12589) <= not (a and b);
    layer2_outputs(12590) <= a and not b;
    layer2_outputs(12591) <= a xor b;
    layer2_outputs(12592) <= b;
    layer2_outputs(12593) <= a or b;
    layer2_outputs(12594) <= not a;
    layer2_outputs(12595) <= b;
    layer2_outputs(12596) <= not (a or b);
    layer2_outputs(12597) <= a and b;
    layer2_outputs(12598) <= a or b;
    layer2_outputs(12599) <= not b or a;
    layer2_outputs(12600) <= b;
    layer2_outputs(12601) <= not a;
    layer2_outputs(12602) <= a xor b;
    layer2_outputs(12603) <= b and not a;
    layer2_outputs(12604) <= a;
    layer2_outputs(12605) <= not (a and b);
    layer2_outputs(12606) <= a xor b;
    layer2_outputs(12607) <= b;
    layer2_outputs(12608) <= not (a and b);
    layer2_outputs(12609) <= a or b;
    layer2_outputs(12610) <= a;
    layer2_outputs(12611) <= a and b;
    layer2_outputs(12612) <= not b;
    layer2_outputs(12613) <= not (a xor b);
    layer2_outputs(12614) <= b and not a;
    layer2_outputs(12615) <= not b;
    layer2_outputs(12616) <= not a;
    layer2_outputs(12617) <= not a or b;
    layer2_outputs(12618) <= a and not b;
    layer2_outputs(12619) <= not a;
    layer2_outputs(12620) <= not b;
    layer2_outputs(12621) <= a and b;
    layer2_outputs(12622) <= not (a and b);
    layer2_outputs(12623) <= not b or a;
    layer2_outputs(12624) <= b;
    layer2_outputs(12625) <= a or b;
    layer2_outputs(12626) <= not a;
    layer2_outputs(12627) <= a and not b;
    layer2_outputs(12628) <= not (a xor b);
    layer2_outputs(12629) <= not (a or b);
    layer2_outputs(12630) <= a and b;
    layer2_outputs(12631) <= a xor b;
    layer2_outputs(12632) <= b;
    layer2_outputs(12633) <= a;
    layer2_outputs(12634) <= not (a and b);
    layer2_outputs(12635) <= not (a and b);
    layer2_outputs(12636) <= not (a xor b);
    layer2_outputs(12637) <= not b;
    layer2_outputs(12638) <= a xor b;
    layer2_outputs(12639) <= a and b;
    layer2_outputs(12640) <= not b;
    layer2_outputs(12641) <= b;
    layer2_outputs(12642) <= a;
    layer2_outputs(12643) <= a and not b;
    layer2_outputs(12644) <= not b or a;
    layer2_outputs(12645) <= not a;
    layer2_outputs(12646) <= a and b;
    layer2_outputs(12647) <= a;
    layer2_outputs(12648) <= b;
    layer2_outputs(12649) <= not b;
    layer2_outputs(12650) <= b;
    layer2_outputs(12651) <= not (a or b);
    layer2_outputs(12652) <= not (a xor b);
    layer2_outputs(12653) <= a and b;
    layer2_outputs(12654) <= not b;
    layer2_outputs(12655) <= a and not b;
    layer2_outputs(12656) <= b and not a;
    layer2_outputs(12657) <= not a;
    layer2_outputs(12658) <= a xor b;
    layer2_outputs(12659) <= not b or a;
    layer2_outputs(12660) <= a and b;
    layer2_outputs(12661) <= a or b;
    layer2_outputs(12662) <= a;
    layer2_outputs(12663) <= not a or b;
    layer2_outputs(12664) <= not b;
    layer2_outputs(12665) <= a and b;
    layer2_outputs(12666) <= a;
    layer2_outputs(12667) <= a xor b;
    layer2_outputs(12668) <= a or b;
    layer2_outputs(12669) <= b;
    layer2_outputs(12670) <= a xor b;
    layer2_outputs(12671) <= not (a xor b);
    layer2_outputs(12672) <= not b or a;
    layer2_outputs(12673) <= not (a xor b);
    layer2_outputs(12674) <= a xor b;
    layer2_outputs(12675) <= a;
    layer2_outputs(12676) <= a and b;
    layer2_outputs(12677) <= not a;
    layer2_outputs(12678) <= b and not a;
    layer2_outputs(12679) <= not b;
    layer2_outputs(12680) <= a;
    layer2_outputs(12681) <= not a;
    layer2_outputs(12682) <= not b;
    layer2_outputs(12683) <= not b;
    layer2_outputs(12684) <= a xor b;
    layer2_outputs(12685) <= not b;
    layer2_outputs(12686) <= not b;
    layer2_outputs(12687) <= a and b;
    layer2_outputs(12688) <= not (a xor b);
    layer2_outputs(12689) <= not b;
    layer2_outputs(12690) <= not b;
    layer2_outputs(12691) <= a and not b;
    layer2_outputs(12692) <= a or b;
    layer2_outputs(12693) <= not (a xor b);
    layer2_outputs(12694) <= a and not b;
    layer2_outputs(12695) <= not b or a;
    layer2_outputs(12696) <= a and not b;
    layer2_outputs(12697) <= b;
    layer2_outputs(12698) <= not (a xor b);
    layer2_outputs(12699) <= not a or b;
    layer2_outputs(12700) <= not (a or b);
    layer2_outputs(12701) <= not (a or b);
    layer2_outputs(12702) <= a;
    layer2_outputs(12703) <= not a;
    layer2_outputs(12704) <= not b;
    layer2_outputs(12705) <= not (a and b);
    layer2_outputs(12706) <= b;
    layer2_outputs(12707) <= not (a or b);
    layer2_outputs(12708) <= not (a or b);
    layer2_outputs(12709) <= not b;
    layer2_outputs(12710) <= not b or a;
    layer2_outputs(12711) <= a and not b;
    layer2_outputs(12712) <= a and not b;
    layer2_outputs(12713) <= a;
    layer2_outputs(12714) <= not b;
    layer2_outputs(12715) <= a and not b;
    layer2_outputs(12716) <= a and not b;
    layer2_outputs(12717) <= not (a xor b);
    layer2_outputs(12718) <= not (a or b);
    layer2_outputs(12719) <= not b;
    layer2_outputs(12720) <= b and not a;
    layer2_outputs(12721) <= a or b;
    layer2_outputs(12722) <= not b;
    layer2_outputs(12723) <= not (a xor b);
    layer2_outputs(12724) <= b;
    layer2_outputs(12725) <= not a;
    layer2_outputs(12726) <= a xor b;
    layer2_outputs(12727) <= a xor b;
    layer2_outputs(12728) <= a xor b;
    layer2_outputs(12729) <= not b;
    layer2_outputs(12730) <= not a;
    layer2_outputs(12731) <= not b or a;
    layer2_outputs(12732) <= not (a xor b);
    layer2_outputs(12733) <= a;
    layer2_outputs(12734) <= a xor b;
    layer2_outputs(12735) <= not a;
    layer2_outputs(12736) <= not (a xor b);
    layer2_outputs(12737) <= not a;
    layer2_outputs(12738) <= a and not b;
    layer2_outputs(12739) <= not (a and b);
    layer2_outputs(12740) <= not a;
    layer2_outputs(12741) <= not a;
    layer2_outputs(12742) <= not a;
    layer2_outputs(12743) <= b;
    layer2_outputs(12744) <= not b or a;
    layer2_outputs(12745) <= not a;
    layer2_outputs(12746) <= not (a and b);
    layer2_outputs(12747) <= b;
    layer2_outputs(12748) <= a;
    layer2_outputs(12749) <= not b or a;
    layer2_outputs(12750) <= not a;
    layer2_outputs(12751) <= not b or a;
    layer2_outputs(12752) <= not a or b;
    layer2_outputs(12753) <= b;
    layer2_outputs(12754) <= a and not b;
    layer2_outputs(12755) <= a or b;
    layer2_outputs(12756) <= not a or b;
    layer2_outputs(12757) <= not (a or b);
    layer2_outputs(12758) <= a xor b;
    layer2_outputs(12759) <= not (a xor b);
    layer2_outputs(12760) <= a and not b;
    layer2_outputs(12761) <= not a;
    layer2_outputs(12762) <= a xor b;
    layer2_outputs(12763) <= not b;
    layer2_outputs(12764) <= a;
    layer2_outputs(12765) <= a or b;
    layer2_outputs(12766) <= a or b;
    layer2_outputs(12767) <= a and not b;
    layer2_outputs(12768) <= a or b;
    layer2_outputs(12769) <= not (a or b);
    layer2_outputs(12770) <= a and not b;
    layer2_outputs(12771) <= not b;
    layer2_outputs(12772) <= b;
    layer2_outputs(12773) <= not a;
    layer2_outputs(12774) <= a or b;
    layer2_outputs(12775) <= a and not b;
    layer2_outputs(12776) <= a xor b;
    layer2_outputs(12777) <= not a;
    layer2_outputs(12778) <= a;
    layer2_outputs(12779) <= not a or b;
    layer2_outputs(12780) <= not (a xor b);
    layer2_outputs(12781) <= a;
    layer2_outputs(12782) <= not (a xor b);
    layer2_outputs(12783) <= not a;
    layer2_outputs(12784) <= not a;
    layer2_outputs(12785) <= not b;
    layer2_outputs(12786) <= a or b;
    layer2_outputs(12787) <= a and b;
    layer2_outputs(12788) <= b;
    layer2_outputs(12789) <= not b;
    layer2_outputs(12790) <= not b or a;
    layer2_outputs(12791) <= a xor b;
    layer2_outputs(12792) <= not a or b;
    layer2_outputs(12793) <= not a;
    layer2_outputs(12794) <= not (a and b);
    layer2_outputs(12795) <= b;
    layer2_outputs(12796) <= not (a and b);
    layer2_outputs(12797) <= a and not b;
    layer2_outputs(12798) <= not a;
    layer2_outputs(12799) <= not a;
    outputs(0) <= not b;
    outputs(1) <= not b;
    outputs(2) <= a xor b;
    outputs(3) <= a and not b;
    outputs(4) <= not (a xor b);
    outputs(5) <= a xor b;
    outputs(6) <= b;
    outputs(7) <= not (a xor b);
    outputs(8) <= not a;
    outputs(9) <= not a;
    outputs(10) <= not (a xor b);
    outputs(11) <= b;
    outputs(12) <= not b;
    outputs(13) <= b;
    outputs(14) <= a;
    outputs(15) <= not a;
    outputs(16) <= not b;
    outputs(17) <= a xor b;
    outputs(18) <= not a;
    outputs(19) <= a xor b;
    outputs(20) <= a and b;
    outputs(21) <= b;
    outputs(22) <= a xor b;
    outputs(23) <= a xor b;
    outputs(24) <= a xor b;
    outputs(25) <= a xor b;
    outputs(26) <= a xor b;
    outputs(27) <= a;
    outputs(28) <= not (a xor b);
    outputs(29) <= not (a xor b);
    outputs(30) <= not a;
    outputs(31) <= b;
    outputs(32) <= not a;
    outputs(33) <= not (a or b);
    outputs(34) <= b;
    outputs(35) <= not (a xor b);
    outputs(36) <= not b;
    outputs(37) <= not (a xor b);
    outputs(38) <= a xor b;
    outputs(39) <= not (a xor b);
    outputs(40) <= not a;
    outputs(41) <= b;
    outputs(42) <= not a;
    outputs(43) <= b and not a;
    outputs(44) <= not b;
    outputs(45) <= a;
    outputs(46) <= not (a xor b);
    outputs(47) <= not (a xor b);
    outputs(48) <= not (a xor b);
    outputs(49) <= a;
    outputs(50) <= a and b;
    outputs(51) <= a and b;
    outputs(52) <= not b or a;
    outputs(53) <= not (a xor b);
    outputs(54) <= a xor b;
    outputs(55) <= a xor b;
    outputs(56) <= a;
    outputs(57) <= a and b;
    outputs(58) <= a xor b;
    outputs(59) <= b;
    outputs(60) <= not a;
    outputs(61) <= b;
    outputs(62) <= a;
    outputs(63) <= b;
    outputs(64) <= not (a xor b);
    outputs(65) <= not (a xor b);
    outputs(66) <= not a;
    outputs(67) <= not (a xor b);
    outputs(68) <= b;
    outputs(69) <= a xor b;
    outputs(70) <= a xor b;
    outputs(71) <= not a or b;
    outputs(72) <= not (a or b);
    outputs(73) <= a or b;
    outputs(74) <= a xor b;
    outputs(75) <= b and not a;
    outputs(76) <= a;
    outputs(77) <= not a;
    outputs(78) <= not (a xor b);
    outputs(79) <= a;
    outputs(80) <= a or b;
    outputs(81) <= a;
    outputs(82) <= a and not b;
    outputs(83) <= a and not b;
    outputs(84) <= not a;
    outputs(85) <= not b;
    outputs(86) <= not (a xor b);
    outputs(87) <= not (a xor b);
    outputs(88) <= a;
    outputs(89) <= b;
    outputs(90) <= b;
    outputs(91) <= not (a xor b);
    outputs(92) <= not (a or b);
    outputs(93) <= not (a and b);
    outputs(94) <= not a;
    outputs(95) <= not (a and b);
    outputs(96) <= not b or a;
    outputs(97) <= b and not a;
    outputs(98) <= a and b;
    outputs(99) <= not b or a;
    outputs(100) <= a xor b;
    outputs(101) <= not a;
    outputs(102) <= not (a xor b);
    outputs(103) <= a;
    outputs(104) <= a xor b;
    outputs(105) <= not b or a;
    outputs(106) <= b;
    outputs(107) <= not (a and b);
    outputs(108) <= a;
    outputs(109) <= b and not a;
    outputs(110) <= not b;
    outputs(111) <= a xor b;
    outputs(112) <= not a;
    outputs(113) <= not b or a;
    outputs(114) <= a;
    outputs(115) <= a and b;
    outputs(116) <= not a;
    outputs(117) <= a xor b;
    outputs(118) <= not (a and b);
    outputs(119) <= not a;
    outputs(120) <= not (a xor b);
    outputs(121) <= not a;
    outputs(122) <= not a;
    outputs(123) <= a or b;
    outputs(124) <= a or b;
    outputs(125) <= a and b;
    outputs(126) <= not a or b;
    outputs(127) <= a and b;
    outputs(128) <= not (a xor b);
    outputs(129) <= b and not a;
    outputs(130) <= a xor b;
    outputs(131) <= not b;
    outputs(132) <= not b;
    outputs(133) <= not b;
    outputs(134) <= a;
    outputs(135) <= not b;
    outputs(136) <= b;
    outputs(137) <= a xor b;
    outputs(138) <= a;
    outputs(139) <= a;
    outputs(140) <= a or b;
    outputs(141) <= not (a xor b);
    outputs(142) <= a xor b;
    outputs(143) <= not (a xor b);
    outputs(144) <= b;
    outputs(145) <= b and not a;
    outputs(146) <= not a;
    outputs(147) <= not b;
    outputs(148) <= not (a xor b);
    outputs(149) <= a;
    outputs(150) <= not b;
    outputs(151) <= a xor b;
    outputs(152) <= a;
    outputs(153) <= not (a xor b);
    outputs(154) <= a and not b;
    outputs(155) <= a;
    outputs(156) <= not b;
    outputs(157) <= not b or a;
    outputs(158) <= b;
    outputs(159) <= a and not b;
    outputs(160) <= not (a xor b);
    outputs(161) <= not (a xor b);
    outputs(162) <= not (a xor b);
    outputs(163) <= b;
    outputs(164) <= a and not b;
    outputs(165) <= a and not b;
    outputs(166) <= not a;
    outputs(167) <= not b;
    outputs(168) <= not a;
    outputs(169) <= b;
    outputs(170) <= not (a xor b);
    outputs(171) <= a xor b;
    outputs(172) <= a and b;
    outputs(173) <= a and not b;
    outputs(174) <= not (a xor b);
    outputs(175) <= not (a xor b);
    outputs(176) <= b;
    outputs(177) <= not (a xor b);
    outputs(178) <= a xor b;
    outputs(179) <= not a or b;
    outputs(180) <= a and not b;
    outputs(181) <= a xor b;
    outputs(182) <= b;
    outputs(183) <= not (a xor b);
    outputs(184) <= not (a xor b);
    outputs(185) <= not b;
    outputs(186) <= not (a or b);
    outputs(187) <= a xor b;
    outputs(188) <= not b;
    outputs(189) <= not (a xor b);
    outputs(190) <= not a;
    outputs(191) <= a xor b;
    outputs(192) <= not a;
    outputs(193) <= not (a xor b);
    outputs(194) <= not b;
    outputs(195) <= not b;
    outputs(196) <= a and not b;
    outputs(197) <= not b;
    outputs(198) <= a xor b;
    outputs(199) <= not b or a;
    outputs(200) <= b;
    outputs(201) <= not a;
    outputs(202) <= b;
    outputs(203) <= b;
    outputs(204) <= not (a and b);
    outputs(205) <= not b;
    outputs(206) <= b;
    outputs(207) <= not b;
    outputs(208) <= not a;
    outputs(209) <= not a;
    outputs(210) <= not b or a;
    outputs(211) <= not (a xor b);
    outputs(212) <= a or b;
    outputs(213) <= b;
    outputs(214) <= not b;
    outputs(215) <= not b;
    outputs(216) <= a and not b;
    outputs(217) <= not (a xor b);
    outputs(218) <= b;
    outputs(219) <= a xor b;
    outputs(220) <= a and b;
    outputs(221) <= a xor b;
    outputs(222) <= not b;
    outputs(223) <= b;
    outputs(224) <= b;
    outputs(225) <= not b;
    outputs(226) <= not (a xor b);
    outputs(227) <= not a or b;
    outputs(228) <= not b;
    outputs(229) <= a xor b;
    outputs(230) <= a xor b;
    outputs(231) <= not b;
    outputs(232) <= a;
    outputs(233) <= not b;
    outputs(234) <= a xor b;
    outputs(235) <= not a;
    outputs(236) <= not b;
    outputs(237) <= a or b;
    outputs(238) <= not a;
    outputs(239) <= not b;
    outputs(240) <= a and not b;
    outputs(241) <= a and b;
    outputs(242) <= not a;
    outputs(243) <= a;
    outputs(244) <= not b;
    outputs(245) <= b;
    outputs(246) <= a and not b;
    outputs(247) <= not b;
    outputs(248) <= not b or a;
    outputs(249) <= a xor b;
    outputs(250) <= a xor b;
    outputs(251) <= a;
    outputs(252) <= not b;
    outputs(253) <= not b;
    outputs(254) <= a xor b;
    outputs(255) <= b;
    outputs(256) <= not a;
    outputs(257) <= a xor b;
    outputs(258) <= a and not b;
    outputs(259) <= b and not a;
    outputs(260) <= not (a and b);
    outputs(261) <= not b or a;
    outputs(262) <= a xor b;
    outputs(263) <= a xor b;
    outputs(264) <= not a;
    outputs(265) <= not b or a;
    outputs(266) <= b;
    outputs(267) <= a;
    outputs(268) <= not a;
    outputs(269) <= not b;
    outputs(270) <= a;
    outputs(271) <= a and b;
    outputs(272) <= b;
    outputs(273) <= a and not b;
    outputs(274) <= b;
    outputs(275) <= not (a xor b);
    outputs(276) <= not (a xor b);
    outputs(277) <= b;
    outputs(278) <= not b;
    outputs(279) <= b;
    outputs(280) <= a and b;
    outputs(281) <= not a;
    outputs(282) <= a and not b;
    outputs(283) <= a xor b;
    outputs(284) <= a xor b;
    outputs(285) <= a xor b;
    outputs(286) <= not a;
    outputs(287) <= b;
    outputs(288) <= b;
    outputs(289) <= b;
    outputs(290) <= a and b;
    outputs(291) <= b;
    outputs(292) <= a;
    outputs(293) <= not (a xor b);
    outputs(294) <= not b;
    outputs(295) <= not (a or b);
    outputs(296) <= not (a or b);
    outputs(297) <= a;
    outputs(298) <= a xor b;
    outputs(299) <= b;
    outputs(300) <= a;
    outputs(301) <= a xor b;
    outputs(302) <= not a;
    outputs(303) <= not a;
    outputs(304) <= not a;
    outputs(305) <= b and not a;
    outputs(306) <= a;
    outputs(307) <= not (a and b);
    outputs(308) <= a;
    outputs(309) <= a;
    outputs(310) <= not a;
    outputs(311) <= not (a or b);
    outputs(312) <= not (a xor b);
    outputs(313) <= a and b;
    outputs(314) <= not b;
    outputs(315) <= not a or b;
    outputs(316) <= not a or b;
    outputs(317) <= a;
    outputs(318) <= not a;
    outputs(319) <= a and b;
    outputs(320) <= a;
    outputs(321) <= not (a xor b);
    outputs(322) <= not (a xor b);
    outputs(323) <= b;
    outputs(324) <= a;
    outputs(325) <= b;
    outputs(326) <= not a;
    outputs(327) <= not (a and b);
    outputs(328) <= a and not b;
    outputs(329) <= not b;
    outputs(330) <= a and not b;
    outputs(331) <= a xor b;
    outputs(332) <= not b;
    outputs(333) <= b and not a;
    outputs(334) <= not a;
    outputs(335) <= not (a xor b);
    outputs(336) <= not b or a;
    outputs(337) <= not b;
    outputs(338) <= a xor b;
    outputs(339) <= not a;
    outputs(340) <= not a;
    outputs(341) <= not b or a;
    outputs(342) <= a;
    outputs(343) <= a;
    outputs(344) <= a xor b;
    outputs(345) <= not (a xor b);
    outputs(346) <= a xor b;
    outputs(347) <= not (a or b);
    outputs(348) <= b;
    outputs(349) <= a xor b;
    outputs(350) <= a;
    outputs(351) <= a;
    outputs(352) <= not a;
    outputs(353) <= b;
    outputs(354) <= b and not a;
    outputs(355) <= not b;
    outputs(356) <= not b;
    outputs(357) <= b;
    outputs(358) <= not b;
    outputs(359) <= a xor b;
    outputs(360) <= not (a xor b);
    outputs(361) <= not (a xor b);
    outputs(362) <= a and not b;
    outputs(363) <= not b;
    outputs(364) <= not a;
    outputs(365) <= not (a xor b);
    outputs(366) <= not a;
    outputs(367) <= a and b;
    outputs(368) <= a xor b;
    outputs(369) <= a;
    outputs(370) <= not (a xor b);
    outputs(371) <= not a;
    outputs(372) <= not (a or b);
    outputs(373) <= not (a or b);
    outputs(374) <= a;
    outputs(375) <= a xor b;
    outputs(376) <= not a;
    outputs(377) <= b;
    outputs(378) <= b and not a;
    outputs(379) <= not a;
    outputs(380) <= a;
    outputs(381) <= b;
    outputs(382) <= not b;
    outputs(383) <= not a;
    outputs(384) <= a and b;
    outputs(385) <= a xor b;
    outputs(386) <= a;
    outputs(387) <= b;
    outputs(388) <= a xor b;
    outputs(389) <= not (a xor b);
    outputs(390) <= not b or a;
    outputs(391) <= a xor b;
    outputs(392) <= a;
    outputs(393) <= a xor b;
    outputs(394) <= a;
    outputs(395) <= a;
    outputs(396) <= not (a xor b);
    outputs(397) <= not a;
    outputs(398) <= not a or b;
    outputs(399) <= a and not b;
    outputs(400) <= not b;
    outputs(401) <= not a;
    outputs(402) <= not (a xor b);
    outputs(403) <= a and not b;
    outputs(404) <= not b or a;
    outputs(405) <= not a;
    outputs(406) <= not b;
    outputs(407) <= not a;
    outputs(408) <= not a;
    outputs(409) <= b;
    outputs(410) <= not b or a;
    outputs(411) <= a xor b;
    outputs(412) <= not (a xor b);
    outputs(413) <= not b;
    outputs(414) <= b;
    outputs(415) <= a;
    outputs(416) <= not a;
    outputs(417) <= not (a xor b);
    outputs(418) <= b;
    outputs(419) <= b and not a;
    outputs(420) <= b;
    outputs(421) <= not b;
    outputs(422) <= not a or b;
    outputs(423) <= not (a or b);
    outputs(424) <= not b;
    outputs(425) <= not (a or b);
    outputs(426) <= not (a xor b);
    outputs(427) <= a;
    outputs(428) <= a xor b;
    outputs(429) <= a xor b;
    outputs(430) <= a;
    outputs(431) <= a xor b;
    outputs(432) <= not b;
    outputs(433) <= not (a xor b);
    outputs(434) <= a or b;
    outputs(435) <= a xor b;
    outputs(436) <= a;
    outputs(437) <= not (a xor b);
    outputs(438) <= b;
    outputs(439) <= b;
    outputs(440) <= a;
    outputs(441) <= a;
    outputs(442) <= b;
    outputs(443) <= a xor b;
    outputs(444) <= not a;
    outputs(445) <= not a or b;
    outputs(446) <= not b;
    outputs(447) <= b and not a;
    outputs(448) <= b;
    outputs(449) <= b and not a;
    outputs(450) <= not (a xor b);
    outputs(451) <= not (a xor b);
    outputs(452) <= not b or a;
    outputs(453) <= not (a xor b);
    outputs(454) <= not a;
    outputs(455) <= not a;
    outputs(456) <= not b;
    outputs(457) <= not a;
    outputs(458) <= a and b;
    outputs(459) <= a;
    outputs(460) <= not b or a;
    outputs(461) <= not a;
    outputs(462) <= a or b;
    outputs(463) <= a;
    outputs(464) <= a and not b;
    outputs(465) <= not (a xor b);
    outputs(466) <= a and b;
    outputs(467) <= not (a and b);
    outputs(468) <= not (a xor b);
    outputs(469) <= not a;
    outputs(470) <= a;
    outputs(471) <= b;
    outputs(472) <= b and not a;
    outputs(473) <= a xor b;
    outputs(474) <= a;
    outputs(475) <= b;
    outputs(476) <= a;
    outputs(477) <= a;
    outputs(478) <= not (a or b);
    outputs(479) <= not (a xor b);
    outputs(480) <= not a;
    outputs(481) <= a xor b;
    outputs(482) <= a xor b;
    outputs(483) <= a and not b;
    outputs(484) <= not (a xor b);
    outputs(485) <= not a;
    outputs(486) <= a and b;
    outputs(487) <= not (a xor b);
    outputs(488) <= a xor b;
    outputs(489) <= a xor b;
    outputs(490) <= not (a xor b);
    outputs(491) <= a and not b;
    outputs(492) <= a or b;
    outputs(493) <= not a;
    outputs(494) <= not (a xor b);
    outputs(495) <= b;
    outputs(496) <= a xor b;
    outputs(497) <= b and not a;
    outputs(498) <= b;
    outputs(499) <= not (a xor b);
    outputs(500) <= not a;
    outputs(501) <= not a;
    outputs(502) <= not (a xor b);
    outputs(503) <= a xor b;
    outputs(504) <= b;
    outputs(505) <= a or b;
    outputs(506) <= a;
    outputs(507) <= a;
    outputs(508) <= a or b;
    outputs(509) <= not a;
    outputs(510) <= a;
    outputs(511) <= not a;
    outputs(512) <= a;
    outputs(513) <= not b;
    outputs(514) <= not a;
    outputs(515) <= not (a xor b);
    outputs(516) <= b;
    outputs(517) <= a;
    outputs(518) <= not (a or b);
    outputs(519) <= b and not a;
    outputs(520) <= a and not b;
    outputs(521) <= not b;
    outputs(522) <= a;
    outputs(523) <= a and b;
    outputs(524) <= not (a xor b);
    outputs(525) <= a;
    outputs(526) <= b;
    outputs(527) <= a and b;
    outputs(528) <= a xor b;
    outputs(529) <= a and b;
    outputs(530) <= a and b;
    outputs(531) <= a xor b;
    outputs(532) <= not (a xor b);
    outputs(533) <= a;
    outputs(534) <= not (a xor b);
    outputs(535) <= a xor b;
    outputs(536) <= a;
    outputs(537) <= a;
    outputs(538) <= a xor b;
    outputs(539) <= not (a xor b);
    outputs(540) <= a xor b;
    outputs(541) <= b;
    outputs(542) <= a;
    outputs(543) <= a or b;
    outputs(544) <= not b or a;
    outputs(545) <= a and not b;
    outputs(546) <= a xor b;
    outputs(547) <= a or b;
    outputs(548) <= a;
    outputs(549) <= not b or a;
    outputs(550) <= b;
    outputs(551) <= not a or b;
    outputs(552) <= a and not b;
    outputs(553) <= not (a xor b);
    outputs(554) <= not a;
    outputs(555) <= b;
    outputs(556) <= a xor b;
    outputs(557) <= not b;
    outputs(558) <= a;
    outputs(559) <= a xor b;
    outputs(560) <= a xor b;
    outputs(561) <= a xor b;
    outputs(562) <= a;
    outputs(563) <= a;
    outputs(564) <= not a;
    outputs(565) <= a xor b;
    outputs(566) <= not a;
    outputs(567) <= not (a xor b);
    outputs(568) <= not b or a;
    outputs(569) <= a and not b;
    outputs(570) <= not b or a;
    outputs(571) <= not a;
    outputs(572) <= not a;
    outputs(573) <= not a;
    outputs(574) <= not b;
    outputs(575) <= not (a xor b);
    outputs(576) <= b;
    outputs(577) <= not (a xor b);
    outputs(578) <= not b;
    outputs(579) <= not a;
    outputs(580) <= a;
    outputs(581) <= not a;
    outputs(582) <= not (a xor b);
    outputs(583) <= a xor b;
    outputs(584) <= not (a or b);
    outputs(585) <= not a;
    outputs(586) <= b;
    outputs(587) <= not a;
    outputs(588) <= a;
    outputs(589) <= b;
    outputs(590) <= not (a xor b);
    outputs(591) <= not b;
    outputs(592) <= a;
    outputs(593) <= a xor b;
    outputs(594) <= not (a xor b);
    outputs(595) <= a and b;
    outputs(596) <= a xor b;
    outputs(597) <= not (a and b);
    outputs(598) <= not b or a;
    outputs(599) <= not a;
    outputs(600) <= a xor b;
    outputs(601) <= not a;
    outputs(602) <= b;
    outputs(603) <= not a;
    outputs(604) <= not b;
    outputs(605) <= not b;
    outputs(606) <= not (a and b);
    outputs(607) <= a xor b;
    outputs(608) <= not (a xor b);
    outputs(609) <= a xor b;
    outputs(610) <= not a;
    outputs(611) <= not (a xor b);
    outputs(612) <= a and b;
    outputs(613) <= not a;
    outputs(614) <= b;
    outputs(615) <= a and not b;
    outputs(616) <= a xor b;
    outputs(617) <= b and not a;
    outputs(618) <= a;
    outputs(619) <= a or b;
    outputs(620) <= b;
    outputs(621) <= not b;
    outputs(622) <= not a;
    outputs(623) <= a and not b;
    outputs(624) <= not (a or b);
    outputs(625) <= not (a xor b);
    outputs(626) <= not (a xor b);
    outputs(627) <= a xor b;
    outputs(628) <= not b;
    outputs(629) <= not (a xor b);
    outputs(630) <= not (a or b);
    outputs(631) <= not a;
    outputs(632) <= not b;
    outputs(633) <= a xor b;
    outputs(634) <= a and b;
    outputs(635) <= not a;
    outputs(636) <= a and not b;
    outputs(637) <= b;
    outputs(638) <= not (a xor b);
    outputs(639) <= a xor b;
    outputs(640) <= not (a or b);
    outputs(641) <= not a;
    outputs(642) <= not b;
    outputs(643) <= a xor b;
    outputs(644) <= not a;
    outputs(645) <= b;
    outputs(646) <= a xor b;
    outputs(647) <= a xor b;
    outputs(648) <= not a;
    outputs(649) <= a xor b;
    outputs(650) <= not b;
    outputs(651) <= not (a and b);
    outputs(652) <= a;
    outputs(653) <= not (a xor b);
    outputs(654) <= not (a or b);
    outputs(655) <= not b;
    outputs(656) <= a and b;
    outputs(657) <= not (a xor b);
    outputs(658) <= not a;
    outputs(659) <= not (a and b);
    outputs(660) <= b;
    outputs(661) <= not b or a;
    outputs(662) <= not (a xor b);
    outputs(663) <= not (a and b);
    outputs(664) <= b;
    outputs(665) <= not a;
    outputs(666) <= b;
    outputs(667) <= not a;
    outputs(668) <= b and not a;
    outputs(669) <= not a;
    outputs(670) <= not (a xor b);
    outputs(671) <= b;
    outputs(672) <= a and not b;
    outputs(673) <= a xor b;
    outputs(674) <= not b;
    outputs(675) <= not a;
    outputs(676) <= a and not b;
    outputs(677) <= not (a and b);
    outputs(678) <= a xor b;
    outputs(679) <= not a or b;
    outputs(680) <= a and not b;
    outputs(681) <= not a;
    outputs(682) <= a;
    outputs(683) <= a and not b;
    outputs(684) <= a xor b;
    outputs(685) <= not a;
    outputs(686) <= not b;
    outputs(687) <= a xor b;
    outputs(688) <= a xor b;
    outputs(689) <= a or b;
    outputs(690) <= not a;
    outputs(691) <= b;
    outputs(692) <= a and b;
    outputs(693) <= not b;
    outputs(694) <= not b;
    outputs(695) <= b and not a;
    outputs(696) <= b;
    outputs(697) <= not b;
    outputs(698) <= a;
    outputs(699) <= a;
    outputs(700) <= not a;
    outputs(701) <= not b;
    outputs(702) <= a and b;
    outputs(703) <= a xor b;
    outputs(704) <= a;
    outputs(705) <= not b;
    outputs(706) <= not b;
    outputs(707) <= a xor b;
    outputs(708) <= a;
    outputs(709) <= b and not a;
    outputs(710) <= not a or b;
    outputs(711) <= not (a and b);
    outputs(712) <= not a or b;
    outputs(713) <= not b or a;
    outputs(714) <= not a or b;
    outputs(715) <= not b;
    outputs(716) <= not b or a;
    outputs(717) <= not (a or b);
    outputs(718) <= not (a or b);
    outputs(719) <= a or b;
    outputs(720) <= not (a xor b);
    outputs(721) <= a;
    outputs(722) <= not (a or b);
    outputs(723) <= not b;
    outputs(724) <= a and not b;
    outputs(725) <= a or b;
    outputs(726) <= not b;
    outputs(727) <= b and not a;
    outputs(728) <= b;
    outputs(729) <= not a;
    outputs(730) <= not (a xor b);
    outputs(731) <= not b or a;
    outputs(732) <= not a;
    outputs(733) <= not (a xor b);
    outputs(734) <= b;
    outputs(735) <= not a or b;
    outputs(736) <= b;
    outputs(737) <= not b;
    outputs(738) <= a xor b;
    outputs(739) <= a;
    outputs(740) <= a or b;
    outputs(741) <= not a;
    outputs(742) <= a and b;
    outputs(743) <= not (a and b);
    outputs(744) <= not b;
    outputs(745) <= a or b;
    outputs(746) <= a and b;
    outputs(747) <= not b;
    outputs(748) <= a xor b;
    outputs(749) <= not (a xor b);
    outputs(750) <= a xor b;
    outputs(751) <= not a;
    outputs(752) <= b;
    outputs(753) <= a xor b;
    outputs(754) <= not b;
    outputs(755) <= not a;
    outputs(756) <= b;
    outputs(757) <= b;
    outputs(758) <= not (a xor b);
    outputs(759) <= a xor b;
    outputs(760) <= a or b;
    outputs(761) <= a xor b;
    outputs(762) <= not b or a;
    outputs(763) <= a xor b;
    outputs(764) <= not (a xor b);
    outputs(765) <= a xor b;
    outputs(766) <= not a;
    outputs(767) <= not (a or b);
    outputs(768) <= not a;
    outputs(769) <= a xor b;
    outputs(770) <= a and b;
    outputs(771) <= b;
    outputs(772) <= b;
    outputs(773) <= a and b;
    outputs(774) <= not (a or b);
    outputs(775) <= a xor b;
    outputs(776) <= a and b;
    outputs(777) <= not b or a;
    outputs(778) <= not (a xor b);
    outputs(779) <= a and not b;
    outputs(780) <= not a;
    outputs(781) <= b;
    outputs(782) <= a xor b;
    outputs(783) <= a xor b;
    outputs(784) <= not b or a;
    outputs(785) <= b and not a;
    outputs(786) <= b and not a;
    outputs(787) <= not a;
    outputs(788) <= a;
    outputs(789) <= a;
    outputs(790) <= a;
    outputs(791) <= a;
    outputs(792) <= a xor b;
    outputs(793) <= a;
    outputs(794) <= a and not b;
    outputs(795) <= not b;
    outputs(796) <= not b or a;
    outputs(797) <= a and b;
    outputs(798) <= a xor b;
    outputs(799) <= a;
    outputs(800) <= not (a xor b);
    outputs(801) <= a;
    outputs(802) <= not b or a;
    outputs(803) <= a;
    outputs(804) <= not (a xor b);
    outputs(805) <= not a;
    outputs(806) <= a and b;
    outputs(807) <= not (a xor b);
    outputs(808) <= a xor b;
    outputs(809) <= not b or a;
    outputs(810) <= not a;
    outputs(811) <= a xor b;
    outputs(812) <= not b;
    outputs(813) <= not b;
    outputs(814) <= a xor b;
    outputs(815) <= b;
    outputs(816) <= not (a or b);
    outputs(817) <= not a;
    outputs(818) <= a xor b;
    outputs(819) <= not a;
    outputs(820) <= a;
    outputs(821) <= not (a xor b);
    outputs(822) <= not a or b;
    outputs(823) <= a xor b;
    outputs(824) <= a;
    outputs(825) <= not (a and b);
    outputs(826) <= a;
    outputs(827) <= a;
    outputs(828) <= not b;
    outputs(829) <= a;
    outputs(830) <= b;
    outputs(831) <= not b;
    outputs(832) <= b;
    outputs(833) <= b and not a;
    outputs(834) <= b;
    outputs(835) <= b;
    outputs(836) <= not (a xor b);
    outputs(837) <= b;
    outputs(838) <= b;
    outputs(839) <= not (a or b);
    outputs(840) <= not a;
    outputs(841) <= a xor b;
    outputs(842) <= not (a xor b);
    outputs(843) <= b and not a;
    outputs(844) <= a or b;
    outputs(845) <= not a;
    outputs(846) <= not (a xor b);
    outputs(847) <= not a;
    outputs(848) <= not a or b;
    outputs(849) <= b;
    outputs(850) <= a xor b;
    outputs(851) <= a;
    outputs(852) <= not a;
    outputs(853) <= a xor b;
    outputs(854) <= a;
    outputs(855) <= a;
    outputs(856) <= a;
    outputs(857) <= b;
    outputs(858) <= not (a xor b);
    outputs(859) <= not b;
    outputs(860) <= not b;
    outputs(861) <= not (a xor b);
    outputs(862) <= not (a xor b);
    outputs(863) <= a and b;
    outputs(864) <= not (a or b);
    outputs(865) <= not a;
    outputs(866) <= a xor b;
    outputs(867) <= a xor b;
    outputs(868) <= a xor b;
    outputs(869) <= a xor b;
    outputs(870) <= a;
    outputs(871) <= a;
    outputs(872) <= not a;
    outputs(873) <= not b;
    outputs(874) <= a;
    outputs(875) <= not (a xor b);
    outputs(876) <= not a;
    outputs(877) <= a xor b;
    outputs(878) <= a xor b;
    outputs(879) <= b;
    outputs(880) <= b;
    outputs(881) <= not a or b;
    outputs(882) <= not (a xor b);
    outputs(883) <= a xor b;
    outputs(884) <= b;
    outputs(885) <= b;
    outputs(886) <= not b;
    outputs(887) <= not b;
    outputs(888) <= not (a xor b);
    outputs(889) <= a xor b;
    outputs(890) <= a;
    outputs(891) <= a and not b;
    outputs(892) <= a and not b;
    outputs(893) <= not a or b;
    outputs(894) <= a and not b;
    outputs(895) <= not a or b;
    outputs(896) <= not b;
    outputs(897) <= b;
    outputs(898) <= a xor b;
    outputs(899) <= not (a and b);
    outputs(900) <= not (a xor b);
    outputs(901) <= not a;
    outputs(902) <= a or b;
    outputs(903) <= b;
    outputs(904) <= a xor b;
    outputs(905) <= not (a xor b);
    outputs(906) <= b;
    outputs(907) <= a;
    outputs(908) <= a and not b;
    outputs(909) <= not a;
    outputs(910) <= a;
    outputs(911) <= a xor b;
    outputs(912) <= not (a or b);
    outputs(913) <= not b;
    outputs(914) <= not (a xor b);
    outputs(915) <= not (a or b);
    outputs(916) <= not a;
    outputs(917) <= a xor b;
    outputs(918) <= not (a xor b);
    outputs(919) <= a and b;
    outputs(920) <= not b;
    outputs(921) <= b and not a;
    outputs(922) <= not b or a;
    outputs(923) <= a;
    outputs(924) <= not (a xor b);
    outputs(925) <= not (a and b);
    outputs(926) <= not (a xor b);
    outputs(927) <= a and b;
    outputs(928) <= a xor b;
    outputs(929) <= b;
    outputs(930) <= not b;
    outputs(931) <= not a;
    outputs(932) <= not b;
    outputs(933) <= a;
    outputs(934) <= not (a xor b);
    outputs(935) <= a;
    outputs(936) <= not (a xor b);
    outputs(937) <= a;
    outputs(938) <= b;
    outputs(939) <= a xor b;
    outputs(940) <= a or b;
    outputs(941) <= a;
    outputs(942) <= a;
    outputs(943) <= not (a xor b);
    outputs(944) <= not b;
    outputs(945) <= a and not b;
    outputs(946) <= not (a or b);
    outputs(947) <= not b;
    outputs(948) <= b;
    outputs(949) <= not (a xor b);
    outputs(950) <= b and not a;
    outputs(951) <= not (a xor b);
    outputs(952) <= a and not b;
    outputs(953) <= a and b;
    outputs(954) <= not (a xor b);
    outputs(955) <= a;
    outputs(956) <= not b;
    outputs(957) <= a or b;
    outputs(958) <= b;
    outputs(959) <= a and not b;
    outputs(960) <= a;
    outputs(961) <= not a;
    outputs(962) <= a xor b;
    outputs(963) <= not a;
    outputs(964) <= not b or a;
    outputs(965) <= not b;
    outputs(966) <= not (a xor b);
    outputs(967) <= a xor b;
    outputs(968) <= not b;
    outputs(969) <= not b;
    outputs(970) <= not a;
    outputs(971) <= not (a xor b);
    outputs(972) <= a xor b;
    outputs(973) <= not b;
    outputs(974) <= not b;
    outputs(975) <= a;
    outputs(976) <= not (a xor b);
    outputs(977) <= a xor b;
    outputs(978) <= b;
    outputs(979) <= not b;
    outputs(980) <= b;
    outputs(981) <= not b or a;
    outputs(982) <= a xor b;
    outputs(983) <= not b;
    outputs(984) <= not b;
    outputs(985) <= a xor b;
    outputs(986) <= not b;
    outputs(987) <= not (a or b);
    outputs(988) <= b;
    outputs(989) <= not a;
    outputs(990) <= b;
    outputs(991) <= not b;
    outputs(992) <= b and not a;
    outputs(993) <= a and b;
    outputs(994) <= a xor b;
    outputs(995) <= not a or b;
    outputs(996) <= b;
    outputs(997) <= not (a and b);
    outputs(998) <= not (a or b);
    outputs(999) <= not b;
    outputs(1000) <= a xor b;
    outputs(1001) <= a and not b;
    outputs(1002) <= not (a and b);
    outputs(1003) <= a;
    outputs(1004) <= not b;
    outputs(1005) <= not a;
    outputs(1006) <= not b;
    outputs(1007) <= b and not a;
    outputs(1008) <= b;
    outputs(1009) <= not (a xor b);
    outputs(1010) <= a;
    outputs(1011) <= b;
    outputs(1012) <= a xor b;
    outputs(1013) <= a or b;
    outputs(1014) <= a xor b;
    outputs(1015) <= b;
    outputs(1016) <= not (a xor b);
    outputs(1017) <= b;
    outputs(1018) <= b;
    outputs(1019) <= a xor b;
    outputs(1020) <= a;
    outputs(1021) <= a or b;
    outputs(1022) <= not a;
    outputs(1023) <= not b;
    outputs(1024) <= not b or a;
    outputs(1025) <= not b;
    outputs(1026) <= not b;
    outputs(1027) <= not a;
    outputs(1028) <= not a or b;
    outputs(1029) <= not a;
    outputs(1030) <= a;
    outputs(1031) <= b;
    outputs(1032) <= not b;
    outputs(1033) <= a and b;
    outputs(1034) <= a xor b;
    outputs(1035) <= not (a xor b);
    outputs(1036) <= not a;
    outputs(1037) <= a and not b;
    outputs(1038) <= not (a and b);
    outputs(1039) <= b;
    outputs(1040) <= not (a xor b);
    outputs(1041) <= b;
    outputs(1042) <= b;
    outputs(1043) <= not (a and b);
    outputs(1044) <= a xor b;
    outputs(1045) <= not b;
    outputs(1046) <= a;
    outputs(1047) <= not (a or b);
    outputs(1048) <= b;
    outputs(1049) <= not (a and b);
    outputs(1050) <= not b;
    outputs(1051) <= not a;
    outputs(1052) <= not b;
    outputs(1053) <= not a;
    outputs(1054) <= not (a xor b);
    outputs(1055) <= not (a xor b);
    outputs(1056) <= not (a xor b);
    outputs(1057) <= not a;
    outputs(1058) <= not b;
    outputs(1059) <= a and b;
    outputs(1060) <= b;
    outputs(1061) <= not (a xor b);
    outputs(1062) <= not (a and b);
    outputs(1063) <= not (a xor b);
    outputs(1064) <= not (a xor b);
    outputs(1065) <= not a;
    outputs(1066) <= not (a xor b);
    outputs(1067) <= a xor b;
    outputs(1068) <= a xor b;
    outputs(1069) <= not a;
    outputs(1070) <= a;
    outputs(1071) <= not (a xor b);
    outputs(1072) <= a xor b;
    outputs(1073) <= not a;
    outputs(1074) <= not a;
    outputs(1075) <= a xor b;
    outputs(1076) <= not b;
    outputs(1077) <= a and not b;
    outputs(1078) <= not (a xor b);
    outputs(1079) <= not a;
    outputs(1080) <= not (a or b);
    outputs(1081) <= a xor b;
    outputs(1082) <= b;
    outputs(1083) <= not a or b;
    outputs(1084) <= a;
    outputs(1085) <= not b;
    outputs(1086) <= a or b;
    outputs(1087) <= not b;
    outputs(1088) <= b and not a;
    outputs(1089) <= a;
    outputs(1090) <= not a;
    outputs(1091) <= b and not a;
    outputs(1092) <= a or b;
    outputs(1093) <= a;
    outputs(1094) <= not a;
    outputs(1095) <= a;
    outputs(1096) <= b;
    outputs(1097) <= not a;
    outputs(1098) <= a xor b;
    outputs(1099) <= not b;
    outputs(1100) <= a;
    outputs(1101) <= not b;
    outputs(1102) <= not b or a;
    outputs(1103) <= b;
    outputs(1104) <= not (a xor b);
    outputs(1105) <= a;
    outputs(1106) <= not b;
    outputs(1107) <= not (a xor b);
    outputs(1108) <= b;
    outputs(1109) <= a;
    outputs(1110) <= not b;
    outputs(1111) <= a and b;
    outputs(1112) <= a xor b;
    outputs(1113) <= not (a xor b);
    outputs(1114) <= not a;
    outputs(1115) <= b and not a;
    outputs(1116) <= not (a or b);
    outputs(1117) <= not (a xor b);
    outputs(1118) <= a xor b;
    outputs(1119) <= not (a xor b);
    outputs(1120) <= not a or b;
    outputs(1121) <= not (a xor b);
    outputs(1122) <= a and b;
    outputs(1123) <= not (a or b);
    outputs(1124) <= a xor b;
    outputs(1125) <= a xor b;
    outputs(1126) <= not a;
    outputs(1127) <= not (a and b);
    outputs(1128) <= not a;
    outputs(1129) <= b and not a;
    outputs(1130) <= not b;
    outputs(1131) <= not (a and b);
    outputs(1132) <= not (a xor b);
    outputs(1133) <= not a;
    outputs(1134) <= a;
    outputs(1135) <= not b or a;
    outputs(1136) <= not b;
    outputs(1137) <= a or b;
    outputs(1138) <= a xor b;
    outputs(1139) <= a xor b;
    outputs(1140) <= b;
    outputs(1141) <= not b;
    outputs(1142) <= not (a xor b);
    outputs(1143) <= not (a and b);
    outputs(1144) <= not b;
    outputs(1145) <= a;
    outputs(1146) <= not b;
    outputs(1147) <= a;
    outputs(1148) <= not (a xor b);
    outputs(1149) <= a;
    outputs(1150) <= not (a xor b);
    outputs(1151) <= not b;
    outputs(1152) <= not b;
    outputs(1153) <= b;
    outputs(1154) <= a;
    outputs(1155) <= not b or a;
    outputs(1156) <= a and b;
    outputs(1157) <= a;
    outputs(1158) <= not b;
    outputs(1159) <= not (a and b);
    outputs(1160) <= not (a xor b);
    outputs(1161) <= not b;
    outputs(1162) <= not b;
    outputs(1163) <= b;
    outputs(1164) <= not a;
    outputs(1165) <= a;
    outputs(1166) <= a;
    outputs(1167) <= a;
    outputs(1168) <= not a;
    outputs(1169) <= not b;
    outputs(1170) <= not (a xor b);
    outputs(1171) <= a xor b;
    outputs(1172) <= not a or b;
    outputs(1173) <= a xor b;
    outputs(1174) <= not b;
    outputs(1175) <= b;
    outputs(1176) <= not b;
    outputs(1177) <= b;
    outputs(1178) <= b;
    outputs(1179) <= not b;
    outputs(1180) <= not (a xor b);
    outputs(1181) <= not a;
    outputs(1182) <= not b;
    outputs(1183) <= a and b;
    outputs(1184) <= a or b;
    outputs(1185) <= not b;
    outputs(1186) <= a and not b;
    outputs(1187) <= not a;
    outputs(1188) <= a;
    outputs(1189) <= not a;
    outputs(1190) <= a;
    outputs(1191) <= a;
    outputs(1192) <= a xor b;
    outputs(1193) <= a and b;
    outputs(1194) <= a;
    outputs(1195) <= a and b;
    outputs(1196) <= a and b;
    outputs(1197) <= a xor b;
    outputs(1198) <= a xor b;
    outputs(1199) <= b and not a;
    outputs(1200) <= b;
    outputs(1201) <= not (a or b);
    outputs(1202) <= not (a and b);
    outputs(1203) <= a or b;
    outputs(1204) <= b and not a;
    outputs(1205) <= a and not b;
    outputs(1206) <= not a;
    outputs(1207) <= not (a or b);
    outputs(1208) <= not b;
    outputs(1209) <= a;
    outputs(1210) <= a xor b;
    outputs(1211) <= not (a xor b);
    outputs(1212) <= a and b;
    outputs(1213) <= a and b;
    outputs(1214) <= a or b;
    outputs(1215) <= a xor b;
    outputs(1216) <= not (a xor b);
    outputs(1217) <= a and b;
    outputs(1218) <= not (a xor b);
    outputs(1219) <= not b or a;
    outputs(1220) <= not b;
    outputs(1221) <= not b;
    outputs(1222) <= not a;
    outputs(1223) <= not b or a;
    outputs(1224) <= not b;
    outputs(1225) <= not (a and b);
    outputs(1226) <= not b or a;
    outputs(1227) <= not a;
    outputs(1228) <= not (a xor b);
    outputs(1229) <= not (a xor b);
    outputs(1230) <= b and not a;
    outputs(1231) <= a;
    outputs(1232) <= not (a xor b);
    outputs(1233) <= not (a xor b);
    outputs(1234) <= not b;
    outputs(1235) <= a;
    outputs(1236) <= a;
    outputs(1237) <= not b or a;
    outputs(1238) <= a and not b;
    outputs(1239) <= not a or b;
    outputs(1240) <= b;
    outputs(1241) <= b;
    outputs(1242) <= a and not b;
    outputs(1243) <= not b;
    outputs(1244) <= not (a and b);
    outputs(1245) <= not (a xor b);
    outputs(1246) <= a or b;
    outputs(1247) <= a or b;
    outputs(1248) <= a;
    outputs(1249) <= a xor b;
    outputs(1250) <= a;
    outputs(1251) <= not a;
    outputs(1252) <= not (a or b);
    outputs(1253) <= a;
    outputs(1254) <= a xor b;
    outputs(1255) <= not (a xor b);
    outputs(1256) <= a or b;
    outputs(1257) <= not (a or b);
    outputs(1258) <= b;
    outputs(1259) <= a;
    outputs(1260) <= not (a xor b);
    outputs(1261) <= not (a xor b);
    outputs(1262) <= not (a xor b);
    outputs(1263) <= not (a and b);
    outputs(1264) <= a;
    outputs(1265) <= not (a xor b);
    outputs(1266) <= a and not b;
    outputs(1267) <= not (a xor b);
    outputs(1268) <= b;
    outputs(1269) <= b and not a;
    outputs(1270) <= a;
    outputs(1271) <= a xor b;
    outputs(1272) <= a xor b;
    outputs(1273) <= b;
    outputs(1274) <= a;
    outputs(1275) <= a xor b;
    outputs(1276) <= not b;
    outputs(1277) <= a and b;
    outputs(1278) <= a and not b;
    outputs(1279) <= b;
    outputs(1280) <= not (a xor b);
    outputs(1281) <= b and not a;
    outputs(1282) <= not (a or b);
    outputs(1283) <= a xor b;
    outputs(1284) <= a xor b;
    outputs(1285) <= a xor b;
    outputs(1286) <= a and not b;
    outputs(1287) <= 1'b0;
    outputs(1288) <= not (a or b);
    outputs(1289) <= a xor b;
    outputs(1290) <= not a or b;
    outputs(1291) <= not b;
    outputs(1292) <= a xor b;
    outputs(1293) <= not (a or b);
    outputs(1294) <= a xor b;
    outputs(1295) <= not (a or b);
    outputs(1296) <= a and not b;
    outputs(1297) <= not b;
    outputs(1298) <= not (a or b);
    outputs(1299) <= not b;
    outputs(1300) <= a;
    outputs(1301) <= a xor b;
    outputs(1302) <= not a;
    outputs(1303) <= a and b;
    outputs(1304) <= not (a or b);
    outputs(1305) <= not a;
    outputs(1306) <= not b;
    outputs(1307) <= not b;
    outputs(1308) <= not (a or b);
    outputs(1309) <= not a;
    outputs(1310) <= a;
    outputs(1311) <= not (a or b);
    outputs(1312) <= a;
    outputs(1313) <= a or b;
    outputs(1314) <= a;
    outputs(1315) <= a xor b;
    outputs(1316) <= not (a or b);
    outputs(1317) <= not (a or b);
    outputs(1318) <= not (a or b);
    outputs(1319) <= not (a or b);
    outputs(1320) <= not a;
    outputs(1321) <= a;
    outputs(1322) <= b and not a;
    outputs(1323) <= not b;
    outputs(1324) <= a xor b;
    outputs(1325) <= a xor b;
    outputs(1326) <= a and not b;
    outputs(1327) <= a xor b;
    outputs(1328) <= a and not b;
    outputs(1329) <= a;
    outputs(1330) <= b;
    outputs(1331) <= a xor b;
    outputs(1332) <= a and not b;
    outputs(1333) <= a and b;
    outputs(1334) <= not (a xor b);
    outputs(1335) <= not b;
    outputs(1336) <= not (a xor b);
    outputs(1337) <= a;
    outputs(1338) <= a and b;
    outputs(1339) <= not b or a;
    outputs(1340) <= a and not b;
    outputs(1341) <= b and not a;
    outputs(1342) <= a xor b;
    outputs(1343) <= not (a xor b);
    outputs(1344) <= not (a xor b);
    outputs(1345) <= a xor b;
    outputs(1346) <= a or b;
    outputs(1347) <= not (a xor b);
    outputs(1348) <= not a;
    outputs(1349) <= not (a xor b);
    outputs(1350) <= b and not a;
    outputs(1351) <= not (a xor b);
    outputs(1352) <= a xor b;
    outputs(1353) <= not a;
    outputs(1354) <= a and not b;
    outputs(1355) <= a xor b;
    outputs(1356) <= not a;
    outputs(1357) <= not b;
    outputs(1358) <= 1'b0;
    outputs(1359) <= not (a or b);
    outputs(1360) <= a xor b;
    outputs(1361) <= b and not a;
    outputs(1362) <= not (a or b);
    outputs(1363) <= a and b;
    outputs(1364) <= not a;
    outputs(1365) <= b and not a;
    outputs(1366) <= a;
    outputs(1367) <= not b;
    outputs(1368) <= a;
    outputs(1369) <= not b;
    outputs(1370) <= a xor b;
    outputs(1371) <= a and not b;
    outputs(1372) <= a xor b;
    outputs(1373) <= b;
    outputs(1374) <= a and not b;
    outputs(1375) <= not a;
    outputs(1376) <= a;
    outputs(1377) <= a xor b;
    outputs(1378) <= b and not a;
    outputs(1379) <= not (a or b);
    outputs(1380) <= a and not b;
    outputs(1381) <= a or b;
    outputs(1382) <= b and not a;
    outputs(1383) <= a xor b;
    outputs(1384) <= a xor b;
    outputs(1385) <= b;
    outputs(1386) <= a and not b;
    outputs(1387) <= a and not b;
    outputs(1388) <= a;
    outputs(1389) <= not a;
    outputs(1390) <= a;
    outputs(1391) <= a and not b;
    outputs(1392) <= not b;
    outputs(1393) <= b;
    outputs(1394) <= a and not b;
    outputs(1395) <= b;
    outputs(1396) <= a xor b;
    outputs(1397) <= a xor b;
    outputs(1398) <= not (a or b);
    outputs(1399) <= not b;
    outputs(1400) <= b and not a;
    outputs(1401) <= a xor b;
    outputs(1402) <= a xor b;
    outputs(1403) <= b and not a;
    outputs(1404) <= not b;
    outputs(1405) <= not b;
    outputs(1406) <= a xor b;
    outputs(1407) <= not b;
    outputs(1408) <= a xor b;
    outputs(1409) <= b;
    outputs(1410) <= not (a xor b);
    outputs(1411) <= a xor b;
    outputs(1412) <= a;
    outputs(1413) <= not b;
    outputs(1414) <= not b;
    outputs(1415) <= a xor b;
    outputs(1416) <= a and not b;
    outputs(1417) <= a;
    outputs(1418) <= not (a or b);
    outputs(1419) <= a and not b;
    outputs(1420) <= a xor b;
    outputs(1421) <= a and b;
    outputs(1422) <= not b;
    outputs(1423) <= a;
    outputs(1424) <= b;
    outputs(1425) <= a xor b;
    outputs(1426) <= not b;
    outputs(1427) <= not (a xor b);
    outputs(1428) <= b and not a;
    outputs(1429) <= b and not a;
    outputs(1430) <= a xor b;
    outputs(1431) <= not (a and b);
    outputs(1432) <= a xor b;
    outputs(1433) <= b and not a;
    outputs(1434) <= not (a xor b);
    outputs(1435) <= not b;
    outputs(1436) <= a and not b;
    outputs(1437) <= not (a xor b);
    outputs(1438) <= not (a or b);
    outputs(1439) <= b;
    outputs(1440) <= a xor b;
    outputs(1441) <= a and not b;
    outputs(1442) <= not (a or b);
    outputs(1443) <= a;
    outputs(1444) <= b and not a;
    outputs(1445) <= a and b;
    outputs(1446) <= not b;
    outputs(1447) <= a xor b;
    outputs(1448) <= a;
    outputs(1449) <= a xor b;
    outputs(1450) <= b and not a;
    outputs(1451) <= not (a xor b);
    outputs(1452) <= a xor b;
    outputs(1453) <= a and b;
    outputs(1454) <= a xor b;
    outputs(1455) <= not (a xor b);
    outputs(1456) <= not (a xor b);
    outputs(1457) <= b and not a;
    outputs(1458) <= a xor b;
    outputs(1459) <= a xor b;
    outputs(1460) <= b and not a;
    outputs(1461) <= a xor b;
    outputs(1462) <= not b;
    outputs(1463) <= b and not a;
    outputs(1464) <= a and b;
    outputs(1465) <= not (a or b);
    outputs(1466) <= not (a xor b);
    outputs(1467) <= a and not b;
    outputs(1468) <= a xor b;
    outputs(1469) <= a;
    outputs(1470) <= a;
    outputs(1471) <= b;
    outputs(1472) <= a and b;
    outputs(1473) <= b and not a;
    outputs(1474) <= a;
    outputs(1475) <= 1'b0;
    outputs(1476) <= b and not a;
    outputs(1477) <= not a;
    outputs(1478) <= a and b;
    outputs(1479) <= not (a xor b);
    outputs(1480) <= not (a xor b);
    outputs(1481) <= a and not b;
    outputs(1482) <= a and not b;
    outputs(1483) <= b;
    outputs(1484) <= a and b;
    outputs(1485) <= not (a or b);
    outputs(1486) <= a xor b;
    outputs(1487) <= b and not a;
    outputs(1488) <= not (a xor b);
    outputs(1489) <= not (a or b);
    outputs(1490) <= a xor b;
    outputs(1491) <= b;
    outputs(1492) <= not (a or b);
    outputs(1493) <= not (a or b);
    outputs(1494) <= a and b;
    outputs(1495) <= b and not a;
    outputs(1496) <= not b;
    outputs(1497) <= not (a xor b);
    outputs(1498) <= a and b;
    outputs(1499) <= a xor b;
    outputs(1500) <= not b;
    outputs(1501) <= not b;
    outputs(1502) <= a xor b;
    outputs(1503) <= a or b;
    outputs(1504) <= a and not b;
    outputs(1505) <= not b;
    outputs(1506) <= a xor b;
    outputs(1507) <= not (a xor b);
    outputs(1508) <= a xor b;
    outputs(1509) <= b and not a;
    outputs(1510) <= a and b;
    outputs(1511) <= a xor b;
    outputs(1512) <= not b;
    outputs(1513) <= a and not b;
    outputs(1514) <= not (a xor b);
    outputs(1515) <= a xor b;
    outputs(1516) <= not b;
    outputs(1517) <= a;
    outputs(1518) <= b and not a;
    outputs(1519) <= not (a xor b);
    outputs(1520) <= a and b;
    outputs(1521) <= not a or b;
    outputs(1522) <= a and b;
    outputs(1523) <= a and not b;
    outputs(1524) <= b;
    outputs(1525) <= not (a or b);
    outputs(1526) <= not (a xor b);
    outputs(1527) <= a xor b;
    outputs(1528) <= not b or a;
    outputs(1529) <= not (a xor b);
    outputs(1530) <= a and not b;
    outputs(1531) <= not (a xor b);
    outputs(1532) <= not b;
    outputs(1533) <= b;
    outputs(1534) <= a xor b;
    outputs(1535) <= not (a xor b);
    outputs(1536) <= a and b;
    outputs(1537) <= a and b;
    outputs(1538) <= a xor b;
    outputs(1539) <= not (a xor b);
    outputs(1540) <= not (a or b);
    outputs(1541) <= not (a xor b);
    outputs(1542) <= a and b;
    outputs(1543) <= a;
    outputs(1544) <= b and not a;
    outputs(1545) <= 1'b0;
    outputs(1546) <= a xor b;
    outputs(1547) <= b;
    outputs(1548) <= a;
    outputs(1549) <= a and not b;
    outputs(1550) <= not b;
    outputs(1551) <= a or b;
    outputs(1552) <= a xor b;
    outputs(1553) <= a xor b;
    outputs(1554) <= not a;
    outputs(1555) <= not (a xor b);
    outputs(1556) <= a and not b;
    outputs(1557) <= b and not a;
    outputs(1558) <= b;
    outputs(1559) <= b;
    outputs(1560) <= a and b;
    outputs(1561) <= b;
    outputs(1562) <= a;
    outputs(1563) <= not b or a;
    outputs(1564) <= not (a xor b);
    outputs(1565) <= a xor b;
    outputs(1566) <= a xor b;
    outputs(1567) <= b and not a;
    outputs(1568) <= not (a xor b);
    outputs(1569) <= b and not a;
    outputs(1570) <= not (a xor b);
    outputs(1571) <= b;
    outputs(1572) <= not a;
    outputs(1573) <= a and b;
    outputs(1574) <= a xor b;
    outputs(1575) <= not (a or b);
    outputs(1576) <= a or b;
    outputs(1577) <= not b;
    outputs(1578) <= not (a xor b);
    outputs(1579) <= b and not a;
    outputs(1580) <= a and b;
    outputs(1581) <= a xor b;
    outputs(1582) <= not b;
    outputs(1583) <= b;
    outputs(1584) <= not (a xor b);
    outputs(1585) <= b;
    outputs(1586) <= not a;
    outputs(1587) <= b and not a;
    outputs(1588) <= not b;
    outputs(1589) <= b;
    outputs(1590) <= not a;
    outputs(1591) <= b;
    outputs(1592) <= a xor b;
    outputs(1593) <= a and b;
    outputs(1594) <= b;
    outputs(1595) <= not b;
    outputs(1596) <= not (a xor b);
    outputs(1597) <= not (a xor b);
    outputs(1598) <= a and not b;
    outputs(1599) <= b;
    outputs(1600) <= not (a xor b);
    outputs(1601) <= not b or a;
    outputs(1602) <= not (a or b);
    outputs(1603) <= not (a or b);
    outputs(1604) <= a and b;
    outputs(1605) <= a;
    outputs(1606) <= not (a or b);
    outputs(1607) <= a and b;
    outputs(1608) <= not a;
    outputs(1609) <= not b;
    outputs(1610) <= not (a xor b);
    outputs(1611) <= a xor b;
    outputs(1612) <= not (a xor b);
    outputs(1613) <= not a or b;
    outputs(1614) <= not (a xor b);
    outputs(1615) <= not (a or b);
    outputs(1616) <= not (a or b);
    outputs(1617) <= a;
    outputs(1618) <= a and b;
    outputs(1619) <= a xor b;
    outputs(1620) <= not (a xor b);
    outputs(1621) <= b;
    outputs(1622) <= a xor b;
    outputs(1623) <= a and b;
    outputs(1624) <= not (a xor b);
    outputs(1625) <= a;
    outputs(1626) <= not (a or b);
    outputs(1627) <= a;
    outputs(1628) <= a;
    outputs(1629) <= a;
    outputs(1630) <= a;
    outputs(1631) <= a and b;
    outputs(1632) <= not b;
    outputs(1633) <= not b;
    outputs(1634) <= a;
    outputs(1635) <= a xor b;
    outputs(1636) <= not (a or b);
    outputs(1637) <= not (a xor b);
    outputs(1638) <= not (a xor b);
    outputs(1639) <= not a or b;
    outputs(1640) <= not b;
    outputs(1641) <= a xor b;
    outputs(1642) <= a and b;
    outputs(1643) <= not (a xor b);
    outputs(1644) <= a xor b;
    outputs(1645) <= 1'b0;
    outputs(1646) <= not (a and b);
    outputs(1647) <= not b;
    outputs(1648) <= a and not b;
    outputs(1649) <= not (a xor b);
    outputs(1650) <= not (a xor b);
    outputs(1651) <= a;
    outputs(1652) <= a xor b;
    outputs(1653) <= b and not a;
    outputs(1654) <= not a;
    outputs(1655) <= not a;
    outputs(1656) <= b and not a;
    outputs(1657) <= a and b;
    outputs(1658) <= not a;
    outputs(1659) <= not b;
    outputs(1660) <= a and not b;
    outputs(1661) <= a and not b;
    outputs(1662) <= b;
    outputs(1663) <= not (a xor b);
    outputs(1664) <= not (a xor b);
    outputs(1665) <= a and not b;
    outputs(1666) <= not (a xor b);
    outputs(1667) <= a xor b;
    outputs(1668) <= not b;
    outputs(1669) <= b and not a;
    outputs(1670) <= not b;
    outputs(1671) <= not (a or b);
    outputs(1672) <= a and not b;
    outputs(1673) <= not (a xor b);
    outputs(1674) <= a xor b;
    outputs(1675) <= a or b;
    outputs(1676) <= a or b;
    outputs(1677) <= b;
    outputs(1678) <= not a;
    outputs(1679) <= a and b;
    outputs(1680) <= not a or b;
    outputs(1681) <= a xor b;
    outputs(1682) <= not (a xor b);
    outputs(1683) <= a;
    outputs(1684) <= a;
    outputs(1685) <= a xor b;
    outputs(1686) <= b and not a;
    outputs(1687) <= a;
    outputs(1688) <= a and b;
    outputs(1689) <= not b;
    outputs(1690) <= b and not a;
    outputs(1691) <= not (a xor b);
    outputs(1692) <= a xor b;
    outputs(1693) <= b;
    outputs(1694) <= not b;
    outputs(1695) <= a and not b;
    outputs(1696) <= a xor b;
    outputs(1697) <= not b;
    outputs(1698) <= b;
    outputs(1699) <= a xor b;
    outputs(1700) <= not (a xor b);
    outputs(1701) <= a xor b;
    outputs(1702) <= b and not a;
    outputs(1703) <= b;
    outputs(1704) <= 1'b0;
    outputs(1705) <= a xor b;
    outputs(1706) <= b;
    outputs(1707) <= not b;
    outputs(1708) <= not (a or b);
    outputs(1709) <= not b;
    outputs(1710) <= b and not a;
    outputs(1711) <= not (a xor b);
    outputs(1712) <= not a;
    outputs(1713) <= not a;
    outputs(1714) <= a and b;
    outputs(1715) <= not (a xor b);
    outputs(1716) <= a and b;
    outputs(1717) <= b and not a;
    outputs(1718) <= a and not b;
    outputs(1719) <= not (a and b);
    outputs(1720) <= a or b;
    outputs(1721) <= not (a or b);
    outputs(1722) <= not (a xor b);
    outputs(1723) <= a and not b;
    outputs(1724) <= a and b;
    outputs(1725) <= a xor b;
    outputs(1726) <= a xor b;
    outputs(1727) <= b and not a;
    outputs(1728) <= a xor b;
    outputs(1729) <= a and not b;
    outputs(1730) <= a and not b;
    outputs(1731) <= not (a xor b);
    outputs(1732) <= a xor b;
    outputs(1733) <= not (a xor b);
    outputs(1734) <= b and not a;
    outputs(1735) <= not b;
    outputs(1736) <= a and not b;
    outputs(1737) <= not b;
    outputs(1738) <= not (a or b);
    outputs(1739) <= 1'b0;
    outputs(1740) <= a xor b;
    outputs(1741) <= b;
    outputs(1742) <= not (a or b);
    outputs(1743) <= a and not b;
    outputs(1744) <= a;
    outputs(1745) <= b;
    outputs(1746) <= b and not a;
    outputs(1747) <= not a;
    outputs(1748) <= a and not b;
    outputs(1749) <= a and not b;
    outputs(1750) <= not b;
    outputs(1751) <= a xor b;
    outputs(1752) <= b and not a;
    outputs(1753) <= a or b;
    outputs(1754) <= a;
    outputs(1755) <= a xor b;
    outputs(1756) <= a xor b;
    outputs(1757) <= not b;
    outputs(1758) <= b;
    outputs(1759) <= a xor b;
    outputs(1760) <= not a;
    outputs(1761) <= a;
    outputs(1762) <= not (a xor b);
    outputs(1763) <= a;
    outputs(1764) <= not (a or b);
    outputs(1765) <= not (a or b);
    outputs(1766) <= a and b;
    outputs(1767) <= not a;
    outputs(1768) <= not (a and b);
    outputs(1769) <= not (a xor b);
    outputs(1770) <= a xor b;
    outputs(1771) <= not (a or b);
    outputs(1772) <= a xor b;
    outputs(1773) <= not (a or b);
    outputs(1774) <= not a;
    outputs(1775) <= b;
    outputs(1776) <= not b;
    outputs(1777) <= a xor b;
    outputs(1778) <= not (a xor b);
    outputs(1779) <= not (a xor b);
    outputs(1780) <= b and not a;
    outputs(1781) <= b and not a;
    outputs(1782) <= not (a xor b);
    outputs(1783) <= not b;
    outputs(1784) <= a and b;
    outputs(1785) <= not (a xor b);
    outputs(1786) <= b;
    outputs(1787) <= a and b;
    outputs(1788) <= a and not b;
    outputs(1789) <= a xor b;
    outputs(1790) <= b and not a;
    outputs(1791) <= a and not b;
    outputs(1792) <= b;
    outputs(1793) <= a xor b;
    outputs(1794) <= a xor b;
    outputs(1795) <= a and b;
    outputs(1796) <= not (a or b);
    outputs(1797) <= a;
    outputs(1798) <= a;
    outputs(1799) <= not b;
    outputs(1800) <= a;
    outputs(1801) <= a xor b;
    outputs(1802) <= a xor b;
    outputs(1803) <= b and not a;
    outputs(1804) <= b and not a;
    outputs(1805) <= not (a or b);
    outputs(1806) <= not a;
    outputs(1807) <= not (a or b);
    outputs(1808) <= not b;
    outputs(1809) <= a xor b;
    outputs(1810) <= a xor b;
    outputs(1811) <= not a;
    outputs(1812) <= a xor b;
    outputs(1813) <= a and not b;
    outputs(1814) <= not a;
    outputs(1815) <= b and not a;
    outputs(1816) <= b;
    outputs(1817) <= a xor b;
    outputs(1818) <= a and b;
    outputs(1819) <= not b;
    outputs(1820) <= not (a or b);
    outputs(1821) <= a and not b;
    outputs(1822) <= not a;
    outputs(1823) <= a xor b;
    outputs(1824) <= a and not b;
    outputs(1825) <= not b;
    outputs(1826) <= b;
    outputs(1827) <= not b;
    outputs(1828) <= a and not b;
    outputs(1829) <= a;
    outputs(1830) <= a;
    outputs(1831) <= not a;
    outputs(1832) <= not (a xor b);
    outputs(1833) <= not a;
    outputs(1834) <= not a;
    outputs(1835) <= a;
    outputs(1836) <= not (a xor b);
    outputs(1837) <= a and b;
    outputs(1838) <= a xor b;
    outputs(1839) <= not (a xor b);
    outputs(1840) <= not (a xor b);
    outputs(1841) <= not (a xor b);
    outputs(1842) <= a xor b;
    outputs(1843) <= not a;
    outputs(1844) <= not a or b;
    outputs(1845) <= b;
    outputs(1846) <= not (a xor b);
    outputs(1847) <= b and not a;
    outputs(1848) <= not (a or b);
    outputs(1849) <= not (a or b);
    outputs(1850) <= a xor b;
    outputs(1851) <= 1'b0;
    outputs(1852) <= a and not b;
    outputs(1853) <= not (a xor b);
    outputs(1854) <= a xor b;
    outputs(1855) <= b;
    outputs(1856) <= not (a or b);
    outputs(1857) <= not (a or b);
    outputs(1858) <= b and not a;
    outputs(1859) <= a and not b;
    outputs(1860) <= not b;
    outputs(1861) <= a;
    outputs(1862) <= not (a xor b);
    outputs(1863) <= a and not b;
    outputs(1864) <= a and not b;
    outputs(1865) <= not b or a;
    outputs(1866) <= not a;
    outputs(1867) <= a xor b;
    outputs(1868) <= not (a or b);
    outputs(1869) <= not a;
    outputs(1870) <= a xor b;
    outputs(1871) <= not (a xor b);
    outputs(1872) <= a;
    outputs(1873) <= not a;
    outputs(1874) <= b;
    outputs(1875) <= 1'b0;
    outputs(1876) <= a and not b;
    outputs(1877) <= not b;
    outputs(1878) <= a and not b;
    outputs(1879) <= not (a xor b);
    outputs(1880) <= not b;
    outputs(1881) <= not b;
    outputs(1882) <= a;
    outputs(1883) <= not a;
    outputs(1884) <= a and not b;
    outputs(1885) <= not (a xor b);
    outputs(1886) <= a;
    outputs(1887) <= b;
    outputs(1888) <= b and not a;
    outputs(1889) <= not (a xor b);
    outputs(1890) <= b;
    outputs(1891) <= a xor b;
    outputs(1892) <= not a;
    outputs(1893) <= not b;
    outputs(1894) <= a and not b;
    outputs(1895) <= b and not a;
    outputs(1896) <= a and b;
    outputs(1897) <= a and b;
    outputs(1898) <= a xor b;
    outputs(1899) <= b;
    outputs(1900) <= not (a xor b);
    outputs(1901) <= a and b;
    outputs(1902) <= b;
    outputs(1903) <= not a;
    outputs(1904) <= b and not a;
    outputs(1905) <= a xor b;
    outputs(1906) <= a and not b;
    outputs(1907) <= not b or a;
    outputs(1908) <= b;
    outputs(1909) <= not (a or b);
    outputs(1910) <= not (a or b);
    outputs(1911) <= a and not b;
    outputs(1912) <= a;
    outputs(1913) <= a and b;
    outputs(1914) <= not (a xor b);
    outputs(1915) <= not (a xor b);
    outputs(1916) <= not (a xor b);
    outputs(1917) <= not (a or b);
    outputs(1918) <= a xor b;
    outputs(1919) <= b and not a;
    outputs(1920) <= not b;
    outputs(1921) <= not b or a;
    outputs(1922) <= a and b;
    outputs(1923) <= not a;
    outputs(1924) <= b;
    outputs(1925) <= not (a xor b);
    outputs(1926) <= b and not a;
    outputs(1927) <= not b;
    outputs(1928) <= a xor b;
    outputs(1929) <= not a;
    outputs(1930) <= a and not b;
    outputs(1931) <= not (a xor b);
    outputs(1932) <= a and b;
    outputs(1933) <= not b;
    outputs(1934) <= not (a or b);
    outputs(1935) <= b;
    outputs(1936) <= not b;
    outputs(1937) <= a and not b;
    outputs(1938) <= not (a xor b);
    outputs(1939) <= a and not b;
    outputs(1940) <= b;
    outputs(1941) <= a and b;
    outputs(1942) <= not a;
    outputs(1943) <= not (a xor b);
    outputs(1944) <= not a;
    outputs(1945) <= not (a xor b);
    outputs(1946) <= a xor b;
    outputs(1947) <= not b or a;
    outputs(1948) <= not (a xor b);
    outputs(1949) <= b and not a;
    outputs(1950) <= a;
    outputs(1951) <= a and not b;
    outputs(1952) <= not (a or b);
    outputs(1953) <= not (a xor b);
    outputs(1954) <= a xor b;
    outputs(1955) <= a;
    outputs(1956) <= not b;
    outputs(1957) <= a and not b;
    outputs(1958) <= b;
    outputs(1959) <= not b;
    outputs(1960) <= a xor b;
    outputs(1961) <= a xor b;
    outputs(1962) <= b and not a;
    outputs(1963) <= a or b;
    outputs(1964) <= a xor b;
    outputs(1965) <= a;
    outputs(1966) <= a and not b;
    outputs(1967) <= a;
    outputs(1968) <= b;
    outputs(1969) <= not a;
    outputs(1970) <= not (a xor b);
    outputs(1971) <= not (a or b);
    outputs(1972) <= a or b;
    outputs(1973) <= not (a xor b);
    outputs(1974) <= not a;
    outputs(1975) <= a xor b;
    outputs(1976) <= a xor b;
    outputs(1977) <= b;
    outputs(1978) <= not b;
    outputs(1979) <= a and b;
    outputs(1980) <= not (a or b);
    outputs(1981) <= a;
    outputs(1982) <= not (a or b);
    outputs(1983) <= a or b;
    outputs(1984) <= not (a or b);
    outputs(1985) <= not (a xor b);
    outputs(1986) <= a xor b;
    outputs(1987) <= not (a xor b);
    outputs(1988) <= not (a xor b);
    outputs(1989) <= a xor b;
    outputs(1990) <= not a;
    outputs(1991) <= not a;
    outputs(1992) <= b;
    outputs(1993) <= not b;
    outputs(1994) <= b;
    outputs(1995) <= not a;
    outputs(1996) <= not b;
    outputs(1997) <= not (a or b);
    outputs(1998) <= not b;
    outputs(1999) <= not b;
    outputs(2000) <= a and not b;
    outputs(2001) <= not b;
    outputs(2002) <= a and b;
    outputs(2003) <= not (a xor b);
    outputs(2004) <= a xor b;
    outputs(2005) <= not a;
    outputs(2006) <= not (a or b);
    outputs(2007) <= not (a or b);
    outputs(2008) <= b and not a;
    outputs(2009) <= b and not a;
    outputs(2010) <= not a;
    outputs(2011) <= b and not a;
    outputs(2012) <= b and not a;
    outputs(2013) <= not b;
    outputs(2014) <= not (a or b);
    outputs(2015) <= a;
    outputs(2016) <= b;
    outputs(2017) <= b and not a;
    outputs(2018) <= not (a xor b);
    outputs(2019) <= a and not b;
    outputs(2020) <= b;
    outputs(2021) <= not (a or b);
    outputs(2022) <= not (a or b);
    outputs(2023) <= not (a xor b);
    outputs(2024) <= a xor b;
    outputs(2025) <= a and b;
    outputs(2026) <= a and b;
    outputs(2027) <= not (a xor b);
    outputs(2028) <= b and not a;
    outputs(2029) <= a xor b;
    outputs(2030) <= not (a xor b);
    outputs(2031) <= b;
    outputs(2032) <= not a;
    outputs(2033) <= b and not a;
    outputs(2034) <= not a;
    outputs(2035) <= a;
    outputs(2036) <= a xor b;
    outputs(2037) <= not (a xor b);
    outputs(2038) <= a and b;
    outputs(2039) <= not (a xor b);
    outputs(2040) <= b;
    outputs(2041) <= a;
    outputs(2042) <= b and not a;
    outputs(2043) <= b and not a;
    outputs(2044) <= not a;
    outputs(2045) <= a;
    outputs(2046) <= a;
    outputs(2047) <= a xor b;
    outputs(2048) <= a and b;
    outputs(2049) <= a xor b;
    outputs(2050) <= not (a or b);
    outputs(2051) <= not (a xor b);
    outputs(2052) <= a and not b;
    outputs(2053) <= not a;
    outputs(2054) <= b;
    outputs(2055) <= not a;
    outputs(2056) <= a and not b;
    outputs(2057) <= not (a xor b);
    outputs(2058) <= a xor b;
    outputs(2059) <= a xor b;
    outputs(2060) <= a and not b;
    outputs(2061) <= b and not a;
    outputs(2062) <= a;
    outputs(2063) <= b and not a;
    outputs(2064) <= not a;
    outputs(2065) <= b and not a;
    outputs(2066) <= not (a xor b);
    outputs(2067) <= not b;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= a and not b;
    outputs(2070) <= not (a or b);
    outputs(2071) <= a and not b;
    outputs(2072) <= a and b;
    outputs(2073) <= a and not b;
    outputs(2074) <= not (a xor b);
    outputs(2075) <= a and not b;
    outputs(2076) <= a and not b;
    outputs(2077) <= not b;
    outputs(2078) <= a and b;
    outputs(2079) <= b;
    outputs(2080) <= not a;
    outputs(2081) <= a and not b;
    outputs(2082) <= not (a xor b);
    outputs(2083) <= not (a or b);
    outputs(2084) <= a xor b;
    outputs(2085) <= a xor b;
    outputs(2086) <= b and not a;
    outputs(2087) <= a and b;
    outputs(2088) <= b and not a;
    outputs(2089) <= a and not b;
    outputs(2090) <= a xor b;
    outputs(2091) <= a xor b;
    outputs(2092) <= a and b;
    outputs(2093) <= a and b;
    outputs(2094) <= not (a xor b);
    outputs(2095) <= not b;
    outputs(2096) <= not (a xor b);
    outputs(2097) <= not b;
    outputs(2098) <= a and b;
    outputs(2099) <= not a;
    outputs(2100) <= a;
    outputs(2101) <= not (a or b);
    outputs(2102) <= a xor b;
    outputs(2103) <= not (a xor b);
    outputs(2104) <= a xor b;
    outputs(2105) <= a and b;
    outputs(2106) <= not (a xor b);
    outputs(2107) <= not a;
    outputs(2108) <= not b;
    outputs(2109) <= a and not b;
    outputs(2110) <= a;
    outputs(2111) <= not a;
    outputs(2112) <= a xor b;
    outputs(2113) <= a;
    outputs(2114) <= a and not b;
    outputs(2115) <= b;
    outputs(2116) <= b and not a;
    outputs(2117) <= not (a xor b);
    outputs(2118) <= not a;
    outputs(2119) <= not (a xor b);
    outputs(2120) <= a xor b;
    outputs(2121) <= a xor b;
    outputs(2122) <= a and b;
    outputs(2123) <= a xor b;
    outputs(2124) <= a xor b;
    outputs(2125) <= not b;
    outputs(2126) <= b;
    outputs(2127) <= not (a or b);
    outputs(2128) <= a;
    outputs(2129) <= not (a xor b);
    outputs(2130) <= not (a xor b);
    outputs(2131) <= not b;
    outputs(2132) <= a and b;
    outputs(2133) <= not b;
    outputs(2134) <= a xor b;
    outputs(2135) <= b;
    outputs(2136) <= a and b;
    outputs(2137) <= not (a xor b);
    outputs(2138) <= not (a xor b);
    outputs(2139) <= not a;
    outputs(2140) <= b and not a;
    outputs(2141) <= a xor b;
    outputs(2142) <= not b;
    outputs(2143) <= a and b;
    outputs(2144) <= a xor b;
    outputs(2145) <= a and not b;
    outputs(2146) <= not (a xor b);
    outputs(2147) <= b;
    outputs(2148) <= not b;
    outputs(2149) <= not (a xor b);
    outputs(2150) <= b;
    outputs(2151) <= not a;
    outputs(2152) <= not a;
    outputs(2153) <= a xor b;
    outputs(2154) <= a xor b;
    outputs(2155) <= not (a or b);
    outputs(2156) <= a xor b;
    outputs(2157) <= a and b;
    outputs(2158) <= a;
    outputs(2159) <= not (a or b);
    outputs(2160) <= b and not a;
    outputs(2161) <= a xor b;
    outputs(2162) <= not (a or b);
    outputs(2163) <= b;
    outputs(2164) <= a;
    outputs(2165) <= a xor b;
    outputs(2166) <= not b;
    outputs(2167) <= a xor b;
    outputs(2168) <= a;
    outputs(2169) <= a xor b;
    outputs(2170) <= not b or a;
    outputs(2171) <= a;
    outputs(2172) <= not a;
    outputs(2173) <= b and not a;
    outputs(2174) <= not b;
    outputs(2175) <= not a;
    outputs(2176) <= not b;
    outputs(2177) <= a xor b;
    outputs(2178) <= not (a xor b);
    outputs(2179) <= a xor b;
    outputs(2180) <= a and b;
    outputs(2181) <= not a or b;
    outputs(2182) <= not b;
    outputs(2183) <= a and not b;
    outputs(2184) <= a and not b;
    outputs(2185) <= b and not a;
    outputs(2186) <= not b;
    outputs(2187) <= a and not b;
    outputs(2188) <= b and not a;
    outputs(2189) <= a and b;
    outputs(2190) <= a xor b;
    outputs(2191) <= a;
    outputs(2192) <= not (a xor b);
    outputs(2193) <= not (a xor b);
    outputs(2194) <= not a;
    outputs(2195) <= a xor b;
    outputs(2196) <= a and not b;
    outputs(2197) <= a xor b;
    outputs(2198) <= not (a xor b);
    outputs(2199) <= a;
    outputs(2200) <= a xor b;
    outputs(2201) <= not (a xor b);
    outputs(2202) <= not (a xor b);
    outputs(2203) <= not a;
    outputs(2204) <= not (a or b);
    outputs(2205) <= a xor b;
    outputs(2206) <= b and not a;
    outputs(2207) <= not (a xor b);
    outputs(2208) <= a xor b;
    outputs(2209) <= a and b;
    outputs(2210) <= a xor b;
    outputs(2211) <= b;
    outputs(2212) <= b;
    outputs(2213) <= not b;
    outputs(2214) <= a and b;
    outputs(2215) <= not a;
    outputs(2216) <= not (a or b);
    outputs(2217) <= not (a xor b);
    outputs(2218) <= b;
    outputs(2219) <= not (a xor b);
    outputs(2220) <= b;
    outputs(2221) <= a;
    outputs(2222) <= not (a or b);
    outputs(2223) <= not (a xor b);
    outputs(2224) <= b;
    outputs(2225) <= not (a xor b);
    outputs(2226) <= a and b;
    outputs(2227) <= a xor b;
    outputs(2228) <= 1'b0;
    outputs(2229) <= not (a xor b);
    outputs(2230) <= a xor b;
    outputs(2231) <= a and not b;
    outputs(2232) <= not (a xor b);
    outputs(2233) <= not a;
    outputs(2234) <= a and not b;
    outputs(2235) <= not a;
    outputs(2236) <= b;
    outputs(2237) <= not (a xor b);
    outputs(2238) <= a xor b;
    outputs(2239) <= a xor b;
    outputs(2240) <= not b or a;
    outputs(2241) <= b;
    outputs(2242) <= not b;
    outputs(2243) <= not (a or b);
    outputs(2244) <= a and not b;
    outputs(2245) <= a and b;
    outputs(2246) <= not (a xor b);
    outputs(2247) <= b and not a;
    outputs(2248) <= not (a xor b);
    outputs(2249) <= not (a or b);
    outputs(2250) <= a;
    outputs(2251) <= not (a xor b);
    outputs(2252) <= a xor b;
    outputs(2253) <= not (a xor b);
    outputs(2254) <= b and not a;
    outputs(2255) <= not (a xor b);
    outputs(2256) <= not (a and b);
    outputs(2257) <= a;
    outputs(2258) <= b and not a;
    outputs(2259) <= b;
    outputs(2260) <= not a;
    outputs(2261) <= b and not a;
    outputs(2262) <= a and b;
    outputs(2263) <= not a;
    outputs(2264) <= not (a xor b);
    outputs(2265) <= not (a xor b);
    outputs(2266) <= not (a or b);
    outputs(2267) <= not (a xor b);
    outputs(2268) <= a xor b;
    outputs(2269) <= b and not a;
    outputs(2270) <= a xor b;
    outputs(2271) <= a;
    outputs(2272) <= a xor b;
    outputs(2273) <= a;
    outputs(2274) <= b and not a;
    outputs(2275) <= a xor b;
    outputs(2276) <= a and not b;
    outputs(2277) <= a and not b;
    outputs(2278) <= a xor b;
    outputs(2279) <= not (a xor b);
    outputs(2280) <= not a;
    outputs(2281) <= not b;
    outputs(2282) <= not (a xor b);
    outputs(2283) <= b;
    outputs(2284) <= 1'b0;
    outputs(2285) <= a and b;
    outputs(2286) <= not (a or b);
    outputs(2287) <= a xor b;
    outputs(2288) <= not (a xor b);
    outputs(2289) <= not b;
    outputs(2290) <= not a;
    outputs(2291) <= a and b;
    outputs(2292) <= not (a xor b);
    outputs(2293) <= not (a or b);
    outputs(2294) <= a xor b;
    outputs(2295) <= not (a xor b);
    outputs(2296) <= a xor b;
    outputs(2297) <= b and not a;
    outputs(2298) <= a and not b;
    outputs(2299) <= not b;
    outputs(2300) <= not b;
    outputs(2301) <= a and not b;
    outputs(2302) <= a and b;
    outputs(2303) <= not (a xor b);
    outputs(2304) <= a xor b;
    outputs(2305) <= not b;
    outputs(2306) <= a;
    outputs(2307) <= a and b;
    outputs(2308) <= not a;
    outputs(2309) <= b;
    outputs(2310) <= not a;
    outputs(2311) <= b;
    outputs(2312) <= b;
    outputs(2313) <= a and not b;
    outputs(2314) <= 1'b0;
    outputs(2315) <= b and not a;
    outputs(2316) <= 1'b0;
    outputs(2317) <= not (a xor b);
    outputs(2318) <= not b;
    outputs(2319) <= a and not b;
    outputs(2320) <= not (a or b);
    outputs(2321) <= not (a xor b);
    outputs(2322) <= not b;
    outputs(2323) <= b;
    outputs(2324) <= not (a or b);
    outputs(2325) <= a;
    outputs(2326) <= a and not b;
    outputs(2327) <= b;
    outputs(2328) <= a xor b;
    outputs(2329) <= a;
    outputs(2330) <= not a;
    outputs(2331) <= not (a or b);
    outputs(2332) <= b;
    outputs(2333) <= b;
    outputs(2334) <= a xor b;
    outputs(2335) <= a;
    outputs(2336) <= a and b;
    outputs(2337) <= a xor b;
    outputs(2338) <= b and not a;
    outputs(2339) <= a xor b;
    outputs(2340) <= a;
    outputs(2341) <= not b or a;
    outputs(2342) <= b and not a;
    outputs(2343) <= not (a or b);
    outputs(2344) <= not b;
    outputs(2345) <= not (a xor b);
    outputs(2346) <= b and not a;
    outputs(2347) <= not (a or b);
    outputs(2348) <= not a;
    outputs(2349) <= a xor b;
    outputs(2350) <= a and b;
    outputs(2351) <= b and not a;
    outputs(2352) <= not (a xor b);
    outputs(2353) <= b and not a;
    outputs(2354) <= a and not b;
    outputs(2355) <= not (a xor b);
    outputs(2356) <= not (a xor b);
    outputs(2357) <= not (a or b);
    outputs(2358) <= not b;
    outputs(2359) <= not (a xor b);
    outputs(2360) <= a xor b;
    outputs(2361) <= b;
    outputs(2362) <= not a or b;
    outputs(2363) <= a;
    outputs(2364) <= not (a xor b);
    outputs(2365) <= not (a or b);
    outputs(2366) <= a;
    outputs(2367) <= not b;
    outputs(2368) <= b;
    outputs(2369) <= b;
    outputs(2370) <= not b or a;
    outputs(2371) <= not (a xor b);
    outputs(2372) <= b;
    outputs(2373) <= b and not a;
    outputs(2374) <= a;
    outputs(2375) <= not a;
    outputs(2376) <= not (a or b);
    outputs(2377) <= not (a or b);
    outputs(2378) <= b and not a;
    outputs(2379) <= 1'b0;
    outputs(2380) <= a and b;
    outputs(2381) <= a and b;
    outputs(2382) <= not a;
    outputs(2383) <= b;
    outputs(2384) <= a and not b;
    outputs(2385) <= a;
    outputs(2386) <= b and not a;
    outputs(2387) <= not (a xor b);
    outputs(2388) <= a;
    outputs(2389) <= not (a or b);
    outputs(2390) <= a xor b;
    outputs(2391) <= not (a or b);
    outputs(2392) <= b and not a;
    outputs(2393) <= not (a or b);
    outputs(2394) <= a xor b;
    outputs(2395) <= 1'b0;
    outputs(2396) <= a and b;
    outputs(2397) <= not b;
    outputs(2398) <= a;
    outputs(2399) <= a and b;
    outputs(2400) <= a xor b;
    outputs(2401) <= a and b;
    outputs(2402) <= b and not a;
    outputs(2403) <= a xor b;
    outputs(2404) <= not (a or b);
    outputs(2405) <= not (a xor b);
    outputs(2406) <= a and b;
    outputs(2407) <= b and not a;
    outputs(2408) <= a and not b;
    outputs(2409) <= a xor b;
    outputs(2410) <= b;
    outputs(2411) <= not (a xor b);
    outputs(2412) <= a and b;
    outputs(2413) <= a;
    outputs(2414) <= b;
    outputs(2415) <= b;
    outputs(2416) <= b and not a;
    outputs(2417) <= not b;
    outputs(2418) <= not a;
    outputs(2419) <= a;
    outputs(2420) <= a xor b;
    outputs(2421) <= a;
    outputs(2422) <= b;
    outputs(2423) <= not (a and b);
    outputs(2424) <= b;
    outputs(2425) <= not (a xor b);
    outputs(2426) <= a;
    outputs(2427) <= a;
    outputs(2428) <= b;
    outputs(2429) <= a and not b;
    outputs(2430) <= not (a xor b);
    outputs(2431) <= a xor b;
    outputs(2432) <= a xor b;
    outputs(2433) <= not b;
    outputs(2434) <= a and not b;
    outputs(2435) <= a and b;
    outputs(2436) <= a and not b;
    outputs(2437) <= a and b;
    outputs(2438) <= a xor b;
    outputs(2439) <= a and b;
    outputs(2440) <= not a;
    outputs(2441) <= a xor b;
    outputs(2442) <= a xor b;
    outputs(2443) <= b;
    outputs(2444) <= a and not b;
    outputs(2445) <= not (a xor b);
    outputs(2446) <= not b;
    outputs(2447) <= not a;
    outputs(2448) <= a and b;
    outputs(2449) <= not (a xor b);
    outputs(2450) <= not (a xor b);
    outputs(2451) <= a xor b;
    outputs(2452) <= not (a xor b);
    outputs(2453) <= not (a or b);
    outputs(2454) <= 1'b0;
    outputs(2455) <= a and not b;
    outputs(2456) <= not (a or b);
    outputs(2457) <= b and not a;
    outputs(2458) <= a xor b;
    outputs(2459) <= a xor b;
    outputs(2460) <= not (a xor b);
    outputs(2461) <= a xor b;
    outputs(2462) <= a and not b;
    outputs(2463) <= a and not b;
    outputs(2464) <= not b;
    outputs(2465) <= not (a xor b);
    outputs(2466) <= not (a or b);
    outputs(2467) <= a xor b;
    outputs(2468) <= not a;
    outputs(2469) <= b;
    outputs(2470) <= b;
    outputs(2471) <= a or b;
    outputs(2472) <= a and not b;
    outputs(2473) <= a xor b;
    outputs(2474) <= not b or a;
    outputs(2475) <= b and not a;
    outputs(2476) <= a xor b;
    outputs(2477) <= b and not a;
    outputs(2478) <= a and not b;
    outputs(2479) <= a and not b;
    outputs(2480) <= a xor b;
    outputs(2481) <= not (a xor b);
    outputs(2482) <= b;
    outputs(2483) <= a xor b;
    outputs(2484) <= not (a xor b);
    outputs(2485) <= a and not b;
    outputs(2486) <= not (a xor b);
    outputs(2487) <= not a;
    outputs(2488) <= a and not b;
    outputs(2489) <= not b;
    outputs(2490) <= a;
    outputs(2491) <= a xor b;
    outputs(2492) <= a xor b;
    outputs(2493) <= a and not b;
    outputs(2494) <= a and b;
    outputs(2495) <= a and not b;
    outputs(2496) <= a;
    outputs(2497) <= not (a xor b);
    outputs(2498) <= a xor b;
    outputs(2499) <= b;
    outputs(2500) <= not a;
    outputs(2501) <= not a;
    outputs(2502) <= not a;
    outputs(2503) <= not (a or b);
    outputs(2504) <= b and not a;
    outputs(2505) <= 1'b0;
    outputs(2506) <= not (a xor b);
    outputs(2507) <= a and not b;
    outputs(2508) <= a and b;
    outputs(2509) <= a xor b;
    outputs(2510) <= a xor b;
    outputs(2511) <= not b;
    outputs(2512) <= not b;
    outputs(2513) <= a and b;
    outputs(2514) <= a xor b;
    outputs(2515) <= a;
    outputs(2516) <= a;
    outputs(2517) <= not (a or b);
    outputs(2518) <= a and b;
    outputs(2519) <= a;
    outputs(2520) <= not a;
    outputs(2521) <= b;
    outputs(2522) <= not (a or b);
    outputs(2523) <= not b;
    outputs(2524) <= a;
    outputs(2525) <= a xor b;
    outputs(2526) <= not b;
    outputs(2527) <= b and not a;
    outputs(2528) <= not (a xor b);
    outputs(2529) <= not a;
    outputs(2530) <= a or b;
    outputs(2531) <= a xor b;
    outputs(2532) <= a and b;
    outputs(2533) <= a and b;
    outputs(2534) <= not b;
    outputs(2535) <= a and not b;
    outputs(2536) <= a and b;
    outputs(2537) <= a or b;
    outputs(2538) <= b;
    outputs(2539) <= not (a or b);
    outputs(2540) <= not (a or b);
    outputs(2541) <= a and b;
    outputs(2542) <= not (a xor b);
    outputs(2543) <= not b;
    outputs(2544) <= not (a or b);
    outputs(2545) <= not b or a;
    outputs(2546) <= 1'b0;
    outputs(2547) <= not b;
    outputs(2548) <= a and not b;
    outputs(2549) <= not b;
    outputs(2550) <= a xor b;
    outputs(2551) <= not a;
    outputs(2552) <= a and not b;
    outputs(2553) <= b and not a;
    outputs(2554) <= b and not a;
    outputs(2555) <= not b;
    outputs(2556) <= b and not a;
    outputs(2557) <= not b;
    outputs(2558) <= a xor b;
    outputs(2559) <= not (a xor b);
    outputs(2560) <= not (a xor b);
    outputs(2561) <= b and not a;
    outputs(2562) <= not a or b;
    outputs(2563) <= not b;
    outputs(2564) <= not b or a;
    outputs(2565) <= not b or a;
    outputs(2566) <= a and not b;
    outputs(2567) <= a xor b;
    outputs(2568) <= a xor b;
    outputs(2569) <= a xor b;
    outputs(2570) <= not b;
    outputs(2571) <= a;
    outputs(2572) <= a;
    outputs(2573) <= a xor b;
    outputs(2574) <= b;
    outputs(2575) <= a xor b;
    outputs(2576) <= a;
    outputs(2577) <= b;
    outputs(2578) <= b and not a;
    outputs(2579) <= not a;
    outputs(2580) <= not b;
    outputs(2581) <= not (a or b);
    outputs(2582) <= a;
    outputs(2583) <= not b or a;
    outputs(2584) <= not (a xor b);
    outputs(2585) <= b and not a;
    outputs(2586) <= a;
    outputs(2587) <= not (a xor b);
    outputs(2588) <= not (a xor b);
    outputs(2589) <= not (a xor b);
    outputs(2590) <= not (a xor b);
    outputs(2591) <= not a;
    outputs(2592) <= not (a xor b);
    outputs(2593) <= b;
    outputs(2594) <= a xor b;
    outputs(2595) <= not b;
    outputs(2596) <= not b or a;
    outputs(2597) <= a and b;
    outputs(2598) <= not a;
    outputs(2599) <= not a;
    outputs(2600) <= a;
    outputs(2601) <= not a;
    outputs(2602) <= a;
    outputs(2603) <= not (a xor b);
    outputs(2604) <= not b;
    outputs(2605) <= b;
    outputs(2606) <= b;
    outputs(2607) <= not (a xor b);
    outputs(2608) <= a and not b;
    outputs(2609) <= a xor b;
    outputs(2610) <= b and not a;
    outputs(2611) <= not a;
    outputs(2612) <= not (a or b);
    outputs(2613) <= a or b;
    outputs(2614) <= not (a or b);
    outputs(2615) <= b and not a;
    outputs(2616) <= a;
    outputs(2617) <= not (a or b);
    outputs(2618) <= b;
    outputs(2619) <= not a;
    outputs(2620) <= b;
    outputs(2621) <= b;
    outputs(2622) <= not a;
    outputs(2623) <= a;
    outputs(2624) <= not b or a;
    outputs(2625) <= a and not b;
    outputs(2626) <= not b;
    outputs(2627) <= b and not a;
    outputs(2628) <= not a;
    outputs(2629) <= b;
    outputs(2630) <= a;
    outputs(2631) <= a or b;
    outputs(2632) <= a xor b;
    outputs(2633) <= not (a xor b);
    outputs(2634) <= not a;
    outputs(2635) <= not (a xor b);
    outputs(2636) <= not a;
    outputs(2637) <= not (a xor b);
    outputs(2638) <= not (a xor b);
    outputs(2639) <= not a;
    outputs(2640) <= not (a xor b);
    outputs(2641) <= a and b;
    outputs(2642) <= b;
    outputs(2643) <= b;
    outputs(2644) <= not a or b;
    outputs(2645) <= a and b;
    outputs(2646) <= a and not b;
    outputs(2647) <= a xor b;
    outputs(2648) <= not (a xor b);
    outputs(2649) <= not (a xor b);
    outputs(2650) <= not b or a;
    outputs(2651) <= a xor b;
    outputs(2652) <= not (a xor b);
    outputs(2653) <= a;
    outputs(2654) <= a xor b;
    outputs(2655) <= not a;
    outputs(2656) <= not b;
    outputs(2657) <= not (a xor b);
    outputs(2658) <= not a;
    outputs(2659) <= not a;
    outputs(2660) <= b;
    outputs(2661) <= b;
    outputs(2662) <= a xor b;
    outputs(2663) <= a and b;
    outputs(2664) <= not (a xor b);
    outputs(2665) <= not (a xor b);
    outputs(2666) <= a or b;
    outputs(2667) <= not b;
    outputs(2668) <= not (a or b);
    outputs(2669) <= not (a and b);
    outputs(2670) <= not (a xor b);
    outputs(2671) <= not (a xor b);
    outputs(2672) <= a;
    outputs(2673) <= a xor b;
    outputs(2674) <= a xor b;
    outputs(2675) <= a;
    outputs(2676) <= not b;
    outputs(2677) <= a xor b;
    outputs(2678) <= not (a xor b);
    outputs(2679) <= a and not b;
    outputs(2680) <= not b;
    outputs(2681) <= not (a or b);
    outputs(2682) <= a and not b;
    outputs(2683) <= a;
    outputs(2684) <= not (a xor b);
    outputs(2685) <= not (a xor b);
    outputs(2686) <= a;
    outputs(2687) <= not b;
    outputs(2688) <= not a;
    outputs(2689) <= not b;
    outputs(2690) <= not (a xor b);
    outputs(2691) <= a and not b;
    outputs(2692) <= a and b;
    outputs(2693) <= a;
    outputs(2694) <= not b;
    outputs(2695) <= not (a xor b);
    outputs(2696) <= b and not a;
    outputs(2697) <= not (a xor b);
    outputs(2698) <= not b;
    outputs(2699) <= b and not a;
    outputs(2700) <= not (a xor b);
    outputs(2701) <= not a;
    outputs(2702) <= b;
    outputs(2703) <= not b;
    outputs(2704) <= b and not a;
    outputs(2705) <= a;
    outputs(2706) <= not a or b;
    outputs(2707) <= a and b;
    outputs(2708) <= not a;
    outputs(2709) <= b and not a;
    outputs(2710) <= not (a xor b);
    outputs(2711) <= b;
    outputs(2712) <= not a;
    outputs(2713) <= not (a xor b);
    outputs(2714) <= not (a xor b);
    outputs(2715) <= a or b;
    outputs(2716) <= a;
    outputs(2717) <= a xor b;
    outputs(2718) <= not (a xor b);
    outputs(2719) <= a xor b;
    outputs(2720) <= not a;
    outputs(2721) <= not (a and b);
    outputs(2722) <= a and b;
    outputs(2723) <= not b or a;
    outputs(2724) <= not (a xor b);
    outputs(2725) <= not (a xor b);
    outputs(2726) <= a;
    outputs(2727) <= a xor b;
    outputs(2728) <= not a or b;
    outputs(2729) <= not (a and b);
    outputs(2730) <= a xor b;
    outputs(2731) <= not b;
    outputs(2732) <= a and not b;
    outputs(2733) <= not b;
    outputs(2734) <= a or b;
    outputs(2735) <= a xor b;
    outputs(2736) <= not b;
    outputs(2737) <= b;
    outputs(2738) <= b;
    outputs(2739) <= not b or a;
    outputs(2740) <= b;
    outputs(2741) <= a and b;
    outputs(2742) <= not b;
    outputs(2743) <= not (a xor b);
    outputs(2744) <= a;
    outputs(2745) <= b;
    outputs(2746) <= b;
    outputs(2747) <= not b;
    outputs(2748) <= not (a xor b);
    outputs(2749) <= a or b;
    outputs(2750) <= not (a xor b);
    outputs(2751) <= not a;
    outputs(2752) <= a xor b;
    outputs(2753) <= not b or a;
    outputs(2754) <= not a;
    outputs(2755) <= a xor b;
    outputs(2756) <= a or b;
    outputs(2757) <= a;
    outputs(2758) <= a xor b;
    outputs(2759) <= a xor b;
    outputs(2760) <= a and not b;
    outputs(2761) <= b;
    outputs(2762) <= a;
    outputs(2763) <= not a;
    outputs(2764) <= a xor b;
    outputs(2765) <= not (a xor b);
    outputs(2766) <= not b;
    outputs(2767) <= not (a or b);
    outputs(2768) <= not (a xor b);
    outputs(2769) <= not b;
    outputs(2770) <= not b;
    outputs(2771) <= a;
    outputs(2772) <= a xor b;
    outputs(2773) <= not a or b;
    outputs(2774) <= a;
    outputs(2775) <= not (a xor b);
    outputs(2776) <= not b;
    outputs(2777) <= a xor b;
    outputs(2778) <= a xor b;
    outputs(2779) <= a;
    outputs(2780) <= b;
    outputs(2781) <= not a;
    outputs(2782) <= b;
    outputs(2783) <= a xor b;
    outputs(2784) <= a xor b;
    outputs(2785) <= not b or a;
    outputs(2786) <= a and not b;
    outputs(2787) <= not b or a;
    outputs(2788) <= not a or b;
    outputs(2789) <= not b or a;
    outputs(2790) <= a xor b;
    outputs(2791) <= b;
    outputs(2792) <= not (a or b);
    outputs(2793) <= a;
    outputs(2794) <= not a or b;
    outputs(2795) <= not b;
    outputs(2796) <= a or b;
    outputs(2797) <= a;
    outputs(2798) <= not (a xor b);
    outputs(2799) <= a xor b;
    outputs(2800) <= b;
    outputs(2801) <= a or b;
    outputs(2802) <= a xor b;
    outputs(2803) <= not (a xor b);
    outputs(2804) <= not b or a;
    outputs(2805) <= b;
    outputs(2806) <= not a or b;
    outputs(2807) <= not (a xor b);
    outputs(2808) <= a xor b;
    outputs(2809) <= not (a xor b);
    outputs(2810) <= not (a xor b);
    outputs(2811) <= not b;
    outputs(2812) <= not b;
    outputs(2813) <= b;
    outputs(2814) <= not (a and b);
    outputs(2815) <= not a or b;
    outputs(2816) <= not a or b;
    outputs(2817) <= a and b;
    outputs(2818) <= not b or a;
    outputs(2819) <= not (a xor b);
    outputs(2820) <= not b;
    outputs(2821) <= not (a xor b);
    outputs(2822) <= not b or a;
    outputs(2823) <= not (a xor b);
    outputs(2824) <= a;
    outputs(2825) <= a;
    outputs(2826) <= b;
    outputs(2827) <= a and b;
    outputs(2828) <= not (a xor b);
    outputs(2829) <= a;
    outputs(2830) <= not (a xor b);
    outputs(2831) <= not b;
    outputs(2832) <= a xor b;
    outputs(2833) <= a and not b;
    outputs(2834) <= b;
    outputs(2835) <= not b;
    outputs(2836) <= not a;
    outputs(2837) <= a xor b;
    outputs(2838) <= not a;
    outputs(2839) <= a or b;
    outputs(2840) <= b;
    outputs(2841) <= b and not a;
    outputs(2842) <= a;
    outputs(2843) <= b and not a;
    outputs(2844) <= not (a xor b);
    outputs(2845) <= a and b;
    outputs(2846) <= a xor b;
    outputs(2847) <= 1'b1;
    outputs(2848) <= not b or a;
    outputs(2849) <= b and not a;
    outputs(2850) <= a xor b;
    outputs(2851) <= not (a and b);
    outputs(2852) <= not b;
    outputs(2853) <= not a;
    outputs(2854) <= not (a or b);
    outputs(2855) <= a and not b;
    outputs(2856) <= not (a and b);
    outputs(2857) <= a xor b;
    outputs(2858) <= a;
    outputs(2859) <= a;
    outputs(2860) <= not (a xor b);
    outputs(2861) <= a xor b;
    outputs(2862) <= not (a xor b);
    outputs(2863) <= not a;
    outputs(2864) <= b;
    outputs(2865) <= not a;
    outputs(2866) <= b;
    outputs(2867) <= b and not a;
    outputs(2868) <= not (a xor b);
    outputs(2869) <= a xor b;
    outputs(2870) <= not (a xor b);
    outputs(2871) <= not (a xor b);
    outputs(2872) <= not a;
    outputs(2873) <= a xor b;
    outputs(2874) <= b;
    outputs(2875) <= b;
    outputs(2876) <= a and b;
    outputs(2877) <= a xor b;
    outputs(2878) <= not a;
    outputs(2879) <= a;
    outputs(2880) <= not b or a;
    outputs(2881) <= not a or b;
    outputs(2882) <= not (a and b);
    outputs(2883) <= not b or a;
    outputs(2884) <= a xor b;
    outputs(2885) <= a and not b;
    outputs(2886) <= not a;
    outputs(2887) <= b;
    outputs(2888) <= not a;
    outputs(2889) <= not b;
    outputs(2890) <= b;
    outputs(2891) <= not a;
    outputs(2892) <= a;
    outputs(2893) <= not a;
    outputs(2894) <= b;
    outputs(2895) <= not b;
    outputs(2896) <= a xor b;
    outputs(2897) <= not b;
    outputs(2898) <= a and b;
    outputs(2899) <= a xor b;
    outputs(2900) <= a or b;
    outputs(2901) <= not (a xor b);
    outputs(2902) <= not a or b;
    outputs(2903) <= not (a xor b);
    outputs(2904) <= not (a or b);
    outputs(2905) <= not a or b;
    outputs(2906) <= a and not b;
    outputs(2907) <= a xor b;
    outputs(2908) <= a xor b;
    outputs(2909) <= not a;
    outputs(2910) <= b;
    outputs(2911) <= not (a xor b);
    outputs(2912) <= b;
    outputs(2913) <= b;
    outputs(2914) <= not (a and b);
    outputs(2915) <= a and not b;
    outputs(2916) <= not a or b;
    outputs(2917) <= b;
    outputs(2918) <= not (a or b);
    outputs(2919) <= b;
    outputs(2920) <= not a;
    outputs(2921) <= not a;
    outputs(2922) <= a or b;
    outputs(2923) <= a;
    outputs(2924) <= b;
    outputs(2925) <= not a;
    outputs(2926) <= a xor b;
    outputs(2927) <= b;
    outputs(2928) <= not a;
    outputs(2929) <= not b or a;
    outputs(2930) <= a or b;
    outputs(2931) <= b and not a;
    outputs(2932) <= a;
    outputs(2933) <= not a;
    outputs(2934) <= not a or b;
    outputs(2935) <= a xor b;
    outputs(2936) <= not b or a;
    outputs(2937) <= not b;
    outputs(2938) <= a;
    outputs(2939) <= not a or b;
    outputs(2940) <= b;
    outputs(2941) <= not (a xor b);
    outputs(2942) <= not b;
    outputs(2943) <= not a;
    outputs(2944) <= not (a and b);
    outputs(2945) <= not (a xor b);
    outputs(2946) <= b and not a;
    outputs(2947) <= not (a xor b);
    outputs(2948) <= a xor b;
    outputs(2949) <= a and not b;
    outputs(2950) <= not b or a;
    outputs(2951) <= not b;
    outputs(2952) <= a and not b;
    outputs(2953) <= b;
    outputs(2954) <= not (a xor b);
    outputs(2955) <= b;
    outputs(2956) <= not (a xor b);
    outputs(2957) <= a xor b;
    outputs(2958) <= b and not a;
    outputs(2959) <= b;
    outputs(2960) <= not b;
    outputs(2961) <= a xor b;
    outputs(2962) <= b;
    outputs(2963) <= a and b;
    outputs(2964) <= b and not a;
    outputs(2965) <= a;
    outputs(2966) <= a xor b;
    outputs(2967) <= not a;
    outputs(2968) <= a;
    outputs(2969) <= not (a xor b);
    outputs(2970) <= not a or b;
    outputs(2971) <= not a or b;
    outputs(2972) <= not (a xor b);
    outputs(2973) <= a;
    outputs(2974) <= not (a xor b);
    outputs(2975) <= a;
    outputs(2976) <= not b or a;
    outputs(2977) <= not (a xor b);
    outputs(2978) <= a or b;
    outputs(2979) <= not (a xor b);
    outputs(2980) <= not a;
    outputs(2981) <= b;
    outputs(2982) <= not a or b;
    outputs(2983) <= b;
    outputs(2984) <= not b;
    outputs(2985) <= not (a and b);
    outputs(2986) <= a and b;
    outputs(2987) <= not (a xor b);
    outputs(2988) <= not a or b;
    outputs(2989) <= not (a or b);
    outputs(2990) <= not b;
    outputs(2991) <= a;
    outputs(2992) <= not a;
    outputs(2993) <= not (a xor b);
    outputs(2994) <= not (a or b);
    outputs(2995) <= not b;
    outputs(2996) <= not (a xor b);
    outputs(2997) <= not a;
    outputs(2998) <= a xor b;
    outputs(2999) <= not (a xor b);
    outputs(3000) <= not (a xor b);
    outputs(3001) <= a and not b;
    outputs(3002) <= not a;
    outputs(3003) <= a;
    outputs(3004) <= a and b;
    outputs(3005) <= a;
    outputs(3006) <= b and not a;
    outputs(3007) <= a and b;
    outputs(3008) <= not (a xor b);
    outputs(3009) <= not a;
    outputs(3010) <= not b or a;
    outputs(3011) <= a and b;
    outputs(3012) <= b;
    outputs(3013) <= not a;
    outputs(3014) <= not (a xor b);
    outputs(3015) <= not a;
    outputs(3016) <= a xor b;
    outputs(3017) <= not b or a;
    outputs(3018) <= a;
    outputs(3019) <= a xor b;
    outputs(3020) <= not a;
    outputs(3021) <= a;
    outputs(3022) <= not (a xor b);
    outputs(3023) <= a xor b;
    outputs(3024) <= b;
    outputs(3025) <= b;
    outputs(3026) <= a xor b;
    outputs(3027) <= not a or b;
    outputs(3028) <= not a;
    outputs(3029) <= b;
    outputs(3030) <= not a;
    outputs(3031) <= not (a xor b);
    outputs(3032) <= not (a xor b);
    outputs(3033) <= a xor b;
    outputs(3034) <= not (a xor b);
    outputs(3035) <= b;
    outputs(3036) <= a;
    outputs(3037) <= not (a xor b);
    outputs(3038) <= not (a xor b);
    outputs(3039) <= not (a xor b);
    outputs(3040) <= not (a xor b);
    outputs(3041) <= not (a and b);
    outputs(3042) <= not (a xor b);
    outputs(3043) <= not (a and b);
    outputs(3044) <= not (a or b);
    outputs(3045) <= not (a xor b);
    outputs(3046) <= not b;
    outputs(3047) <= not a or b;
    outputs(3048) <= not b;
    outputs(3049) <= a xor b;
    outputs(3050) <= b and not a;
    outputs(3051) <= a xor b;
    outputs(3052) <= not (a xor b);
    outputs(3053) <= b;
    outputs(3054) <= b;
    outputs(3055) <= a and not b;
    outputs(3056) <= a;
    outputs(3057) <= not a or b;
    outputs(3058) <= not b;
    outputs(3059) <= not (a xor b);
    outputs(3060) <= not (a or b);
    outputs(3061) <= b;
    outputs(3062) <= not (a xor b);
    outputs(3063) <= not (a xor b);
    outputs(3064) <= a xor b;
    outputs(3065) <= a;
    outputs(3066) <= a;
    outputs(3067) <= a xor b;
    outputs(3068) <= not (a xor b);
    outputs(3069) <= not (a xor b);
    outputs(3070) <= a and b;
    outputs(3071) <= not a;
    outputs(3072) <= a xor b;
    outputs(3073) <= a xor b;
    outputs(3074) <= a xor b;
    outputs(3075) <= not (a xor b);
    outputs(3076) <= not b or a;
    outputs(3077) <= not a;
    outputs(3078) <= not (a xor b);
    outputs(3079) <= a xor b;
    outputs(3080) <= not b;
    outputs(3081) <= not a or b;
    outputs(3082) <= a;
    outputs(3083) <= not (a xor b);
    outputs(3084) <= not a;
    outputs(3085) <= b;
    outputs(3086) <= a xor b;
    outputs(3087) <= a and not b;
    outputs(3088) <= not a or b;
    outputs(3089) <= not (a xor b);
    outputs(3090) <= a;
    outputs(3091) <= not (a xor b);
    outputs(3092) <= a and b;
    outputs(3093) <= not a or b;
    outputs(3094) <= not b;
    outputs(3095) <= b;
    outputs(3096) <= not a or b;
    outputs(3097) <= not a;
    outputs(3098) <= not (a and b);
    outputs(3099) <= not b or a;
    outputs(3100) <= a and not b;
    outputs(3101) <= not (a and b);
    outputs(3102) <= not a;
    outputs(3103) <= a xor b;
    outputs(3104) <= not (a xor b);
    outputs(3105) <= not (a xor b);
    outputs(3106) <= b;
    outputs(3107) <= a;
    outputs(3108) <= not b;
    outputs(3109) <= a;
    outputs(3110) <= a xor b;
    outputs(3111) <= not a;
    outputs(3112) <= not b;
    outputs(3113) <= not (a xor b);
    outputs(3114) <= not b;
    outputs(3115) <= not a;
    outputs(3116) <= a or b;
    outputs(3117) <= a and b;
    outputs(3118) <= a xor b;
    outputs(3119) <= a or b;
    outputs(3120) <= a xor b;
    outputs(3121) <= a and b;
    outputs(3122) <= a xor b;
    outputs(3123) <= not b;
    outputs(3124) <= a or b;
    outputs(3125) <= b;
    outputs(3126) <= a;
    outputs(3127) <= a xor b;
    outputs(3128) <= a;
    outputs(3129) <= not (a xor b);
    outputs(3130) <= not (a xor b);
    outputs(3131) <= not (a xor b);
    outputs(3132) <= a xor b;
    outputs(3133) <= not a;
    outputs(3134) <= a xor b;
    outputs(3135) <= a and not b;
    outputs(3136) <= b;
    outputs(3137) <= not (a xor b);
    outputs(3138) <= not a;
    outputs(3139) <= a or b;
    outputs(3140) <= not b;
    outputs(3141) <= a xor b;
    outputs(3142) <= a xor b;
    outputs(3143) <= not a;
    outputs(3144) <= b;
    outputs(3145) <= a and not b;
    outputs(3146) <= a;
    outputs(3147) <= a xor b;
    outputs(3148) <= not a or b;
    outputs(3149) <= a and not b;
    outputs(3150) <= not (a xor b);
    outputs(3151) <= a xor b;
    outputs(3152) <= a;
    outputs(3153) <= a xor b;
    outputs(3154) <= not a;
    outputs(3155) <= a xor b;
    outputs(3156) <= a xor b;
    outputs(3157) <= not a;
    outputs(3158) <= not (a xor b);
    outputs(3159) <= not b;
    outputs(3160) <= not a;
    outputs(3161) <= not a;
    outputs(3162) <= a xor b;
    outputs(3163) <= a xor b;
    outputs(3164) <= not a or b;
    outputs(3165) <= not (a xor b);
    outputs(3166) <= not a;
    outputs(3167) <= not a;
    outputs(3168) <= not a or b;
    outputs(3169) <= a xor b;
    outputs(3170) <= a xor b;
    outputs(3171) <= a;
    outputs(3172) <= b;
    outputs(3173) <= a;
    outputs(3174) <= not (a and b);
    outputs(3175) <= not (a and b);
    outputs(3176) <= not a;
    outputs(3177) <= not (a or b);
    outputs(3178) <= not b;
    outputs(3179) <= not b;
    outputs(3180) <= a;
    outputs(3181) <= not (a xor b);
    outputs(3182) <= a xor b;
    outputs(3183) <= a;
    outputs(3184) <= not b;
    outputs(3185) <= a and b;
    outputs(3186) <= b;
    outputs(3187) <= b;
    outputs(3188) <= not a;
    outputs(3189) <= b;
    outputs(3190) <= a xor b;
    outputs(3191) <= a xor b;
    outputs(3192) <= not (a and b);
    outputs(3193) <= a xor b;
    outputs(3194) <= not b;
    outputs(3195) <= not (a xor b);
    outputs(3196) <= a;
    outputs(3197) <= not (a xor b);
    outputs(3198) <= not (a xor b);
    outputs(3199) <= not b;
    outputs(3200) <= not a;
    outputs(3201) <= not b;
    outputs(3202) <= not a;
    outputs(3203) <= a;
    outputs(3204) <= a and not b;
    outputs(3205) <= not (a xor b);
    outputs(3206) <= not (a xor b);
    outputs(3207) <= b;
    outputs(3208) <= not (a or b);
    outputs(3209) <= not (a xor b);
    outputs(3210) <= b;
    outputs(3211) <= a or b;
    outputs(3212) <= not b;
    outputs(3213) <= a xor b;
    outputs(3214) <= b;
    outputs(3215) <= not b or a;
    outputs(3216) <= not b or a;
    outputs(3217) <= a xor b;
    outputs(3218) <= a;
    outputs(3219) <= not (a or b);
    outputs(3220) <= not (a xor b);
    outputs(3221) <= not (a and b);
    outputs(3222) <= not (a xor b);
    outputs(3223) <= a xor b;
    outputs(3224) <= not (a xor b);
    outputs(3225) <= not (a xor b);
    outputs(3226) <= not (a and b);
    outputs(3227) <= a xor b;
    outputs(3228) <= b;
    outputs(3229) <= a and not b;
    outputs(3230) <= a and not b;
    outputs(3231) <= not b;
    outputs(3232) <= a xor b;
    outputs(3233) <= b;
    outputs(3234) <= a or b;
    outputs(3235) <= a xor b;
    outputs(3236) <= a;
    outputs(3237) <= not b;
    outputs(3238) <= b and not a;
    outputs(3239) <= not (a xor b);
    outputs(3240) <= b and not a;
    outputs(3241) <= b;
    outputs(3242) <= a xor b;
    outputs(3243) <= not (a xor b);
    outputs(3244) <= a and b;
    outputs(3245) <= b;
    outputs(3246) <= not b;
    outputs(3247) <= b;
    outputs(3248) <= b and not a;
    outputs(3249) <= a or b;
    outputs(3250) <= not (a xor b);
    outputs(3251) <= not (a or b);
    outputs(3252) <= a xor b;
    outputs(3253) <= a xor b;
    outputs(3254) <= a xor b;
    outputs(3255) <= not b or a;
    outputs(3256) <= a xor b;
    outputs(3257) <= a;
    outputs(3258) <= not b;
    outputs(3259) <= not (a xor b);
    outputs(3260) <= a;
    outputs(3261) <= a xor b;
    outputs(3262) <= not b;
    outputs(3263) <= not (a xor b);
    outputs(3264) <= not a;
    outputs(3265) <= not a;
    outputs(3266) <= a and not b;
    outputs(3267) <= not (a or b);
    outputs(3268) <= not a;
    outputs(3269) <= a and b;
    outputs(3270) <= not a or b;
    outputs(3271) <= a and b;
    outputs(3272) <= a or b;
    outputs(3273) <= not (a xor b);
    outputs(3274) <= a and not b;
    outputs(3275) <= a xor b;
    outputs(3276) <= not b;
    outputs(3277) <= not a;
    outputs(3278) <= a;
    outputs(3279) <= a and b;
    outputs(3280) <= b;
    outputs(3281) <= a;
    outputs(3282) <= a xor b;
    outputs(3283) <= not a or b;
    outputs(3284) <= not a or b;
    outputs(3285) <= a xor b;
    outputs(3286) <= not (a and b);
    outputs(3287) <= not (a xor b);
    outputs(3288) <= a and b;
    outputs(3289) <= not (a or b);
    outputs(3290) <= not a;
    outputs(3291) <= b;
    outputs(3292) <= not (a xor b);
    outputs(3293) <= not (a xor b);
    outputs(3294) <= b;
    outputs(3295) <= a or b;
    outputs(3296) <= not b or a;
    outputs(3297) <= b;
    outputs(3298) <= b and not a;
    outputs(3299) <= not a;
    outputs(3300) <= a;
    outputs(3301) <= a xor b;
    outputs(3302) <= not b;
    outputs(3303) <= not (a xor b);
    outputs(3304) <= not b;
    outputs(3305) <= not (a and b);
    outputs(3306) <= a xor b;
    outputs(3307) <= a;
    outputs(3308) <= not (a or b);
    outputs(3309) <= a xor b;
    outputs(3310) <= not (a and b);
    outputs(3311) <= not b;
    outputs(3312) <= not a;
    outputs(3313) <= not (a xor b);
    outputs(3314) <= a xor b;
    outputs(3315) <= a xor b;
    outputs(3316) <= b;
    outputs(3317) <= not a;
    outputs(3318) <= not (a xor b);
    outputs(3319) <= a;
    outputs(3320) <= not b;
    outputs(3321) <= a xor b;
    outputs(3322) <= not a;
    outputs(3323) <= not (a and b);
    outputs(3324) <= a xor b;
    outputs(3325) <= not (a or b);
    outputs(3326) <= not b;
    outputs(3327) <= not b or a;
    outputs(3328) <= b and not a;
    outputs(3329) <= not (a xor b);
    outputs(3330) <= not b;
    outputs(3331) <= a xor b;
    outputs(3332) <= a or b;
    outputs(3333) <= not (a xor b);
    outputs(3334) <= not a;
    outputs(3335) <= a xor b;
    outputs(3336) <= b and not a;
    outputs(3337) <= not b;
    outputs(3338) <= b;
    outputs(3339) <= not (a xor b);
    outputs(3340) <= not (a xor b);
    outputs(3341) <= not b;
    outputs(3342) <= b;
    outputs(3343) <= a and not b;
    outputs(3344) <= a and b;
    outputs(3345) <= b;
    outputs(3346) <= not (a xor b);
    outputs(3347) <= b;
    outputs(3348) <= not a;
    outputs(3349) <= not (a xor b);
    outputs(3350) <= not b;
    outputs(3351) <= a;
    outputs(3352) <= not (a xor b);
    outputs(3353) <= not a;
    outputs(3354) <= not a or b;
    outputs(3355) <= not b;
    outputs(3356) <= a and not b;
    outputs(3357) <= not a or b;
    outputs(3358) <= b;
    outputs(3359) <= not a;
    outputs(3360) <= not a;
    outputs(3361) <= a xor b;
    outputs(3362) <= not (a and b);
    outputs(3363) <= a xor b;
    outputs(3364) <= a or b;
    outputs(3365) <= not (a xor b);
    outputs(3366) <= b;
    outputs(3367) <= a xor b;
    outputs(3368) <= a and b;
    outputs(3369) <= not a;
    outputs(3370) <= a xor b;
    outputs(3371) <= not a;
    outputs(3372) <= a;
    outputs(3373) <= not (a xor b);
    outputs(3374) <= not a or b;
    outputs(3375) <= not (a xor b);
    outputs(3376) <= not (a or b);
    outputs(3377) <= not a or b;
    outputs(3378) <= a and b;
    outputs(3379) <= not a;
    outputs(3380) <= a;
    outputs(3381) <= not (a xor b);
    outputs(3382) <= not b;
    outputs(3383) <= a or b;
    outputs(3384) <= not b;
    outputs(3385) <= not b;
    outputs(3386) <= not b;
    outputs(3387) <= a xor b;
    outputs(3388) <= a or b;
    outputs(3389) <= b;
    outputs(3390) <= not a;
    outputs(3391) <= a xor b;
    outputs(3392) <= not b;
    outputs(3393) <= not (a xor b);
    outputs(3394) <= not a;
    outputs(3395) <= b and not a;
    outputs(3396) <= b;
    outputs(3397) <= not (a xor b);
    outputs(3398) <= a and not b;
    outputs(3399) <= a and b;
    outputs(3400) <= b and not a;
    outputs(3401) <= not a;
    outputs(3402) <= b;
    outputs(3403) <= not (a and b);
    outputs(3404) <= not (a and b);
    outputs(3405) <= a xor b;
    outputs(3406) <= a xor b;
    outputs(3407) <= not b;
    outputs(3408) <= not (a xor b);
    outputs(3409) <= a;
    outputs(3410) <= not a;
    outputs(3411) <= not a or b;
    outputs(3412) <= a xor b;
    outputs(3413) <= not (a and b);
    outputs(3414) <= b;
    outputs(3415) <= a and b;
    outputs(3416) <= a xor b;
    outputs(3417) <= not (a xor b);
    outputs(3418) <= b;
    outputs(3419) <= not (a xor b);
    outputs(3420) <= not (a or b);
    outputs(3421) <= not b;
    outputs(3422) <= not b;
    outputs(3423) <= a;
    outputs(3424) <= a;
    outputs(3425) <= b and not a;
    outputs(3426) <= not a or b;
    outputs(3427) <= not a;
    outputs(3428) <= a and b;
    outputs(3429) <= not (a xor b);
    outputs(3430) <= a xor b;
    outputs(3431) <= not a;
    outputs(3432) <= not (a or b);
    outputs(3433) <= a xor b;
    outputs(3434) <= b and not a;
    outputs(3435) <= not a or b;
    outputs(3436) <= not (a and b);
    outputs(3437) <= not (a xor b);
    outputs(3438) <= b and not a;
    outputs(3439) <= a and b;
    outputs(3440) <= not b;
    outputs(3441) <= not a;
    outputs(3442) <= a xor b;
    outputs(3443) <= not (a xor b);
    outputs(3444) <= a or b;
    outputs(3445) <= not b;
    outputs(3446) <= a;
    outputs(3447) <= a;
    outputs(3448) <= not a or b;
    outputs(3449) <= b;
    outputs(3450) <= not b;
    outputs(3451) <= not b or a;
    outputs(3452) <= a and b;
    outputs(3453) <= a or b;
    outputs(3454) <= a xor b;
    outputs(3455) <= a xor b;
    outputs(3456) <= b;
    outputs(3457) <= a or b;
    outputs(3458) <= not b or a;
    outputs(3459) <= not (a or b);
    outputs(3460) <= a xor b;
    outputs(3461) <= not b or a;
    outputs(3462) <= a xor b;
    outputs(3463) <= a and not b;
    outputs(3464) <= not b;
    outputs(3465) <= not b or a;
    outputs(3466) <= b;
    outputs(3467) <= a;
    outputs(3468) <= not b;
    outputs(3469) <= not b;
    outputs(3470) <= not (a xor b);
    outputs(3471) <= not b;
    outputs(3472) <= not a;
    outputs(3473) <= not a;
    outputs(3474) <= a xor b;
    outputs(3475) <= a xor b;
    outputs(3476) <= not a;
    outputs(3477) <= not a;
    outputs(3478) <= b and not a;
    outputs(3479) <= a;
    outputs(3480) <= not a;
    outputs(3481) <= not a;
    outputs(3482) <= not (a xor b);
    outputs(3483) <= a;
    outputs(3484) <= not b;
    outputs(3485) <= a or b;
    outputs(3486) <= not (a xor b);
    outputs(3487) <= not (a xor b);
    outputs(3488) <= not b;
    outputs(3489) <= a;
    outputs(3490) <= b;
    outputs(3491) <= not a;
    outputs(3492) <= not b or a;
    outputs(3493) <= a or b;
    outputs(3494) <= a and b;
    outputs(3495) <= not b;
    outputs(3496) <= a xor b;
    outputs(3497) <= not (a xor b);
    outputs(3498) <= not a or b;
    outputs(3499) <= b;
    outputs(3500) <= not a or b;
    outputs(3501) <= not (a xor b);
    outputs(3502) <= not b;
    outputs(3503) <= a and not b;
    outputs(3504) <= not b;
    outputs(3505) <= b;
    outputs(3506) <= not (a and b);
    outputs(3507) <= not a;
    outputs(3508) <= not a;
    outputs(3509) <= not b;
    outputs(3510) <= a xor b;
    outputs(3511) <= not (a xor b);
    outputs(3512) <= b;
    outputs(3513) <= a;
    outputs(3514) <= a xor b;
    outputs(3515) <= not (a and b);
    outputs(3516) <= not b;
    outputs(3517) <= not a or b;
    outputs(3518) <= a xor b;
    outputs(3519) <= b;
    outputs(3520) <= not a or b;
    outputs(3521) <= a;
    outputs(3522) <= a xor b;
    outputs(3523) <= a;
    outputs(3524) <= b;
    outputs(3525) <= a or b;
    outputs(3526) <= a xor b;
    outputs(3527) <= not a;
    outputs(3528) <= b;
    outputs(3529) <= not a;
    outputs(3530) <= not a;
    outputs(3531) <= a or b;
    outputs(3532) <= not b;
    outputs(3533) <= not a;
    outputs(3534) <= not a;
    outputs(3535) <= not a;
    outputs(3536) <= not b or a;
    outputs(3537) <= not a;
    outputs(3538) <= not a;
    outputs(3539) <= a;
    outputs(3540) <= not (a xor b);
    outputs(3541) <= b;
    outputs(3542) <= a xor b;
    outputs(3543) <= a;
    outputs(3544) <= not b;
    outputs(3545) <= not a;
    outputs(3546) <= not (a xor b);
    outputs(3547) <= not (a and b);
    outputs(3548) <= a;
    outputs(3549) <= not a or b;
    outputs(3550) <= a and b;
    outputs(3551) <= a or b;
    outputs(3552) <= a;
    outputs(3553) <= not (a and b);
    outputs(3554) <= a or b;
    outputs(3555) <= not b or a;
    outputs(3556) <= not a;
    outputs(3557) <= not (a xor b);
    outputs(3558) <= not (a xor b);
    outputs(3559) <= not b;
    outputs(3560) <= not (a xor b);
    outputs(3561) <= a and not b;
    outputs(3562) <= not a;
    outputs(3563) <= b;
    outputs(3564) <= not (a xor b);
    outputs(3565) <= not b;
    outputs(3566) <= a and not b;
    outputs(3567) <= a xor b;
    outputs(3568) <= not a;
    outputs(3569) <= b;
    outputs(3570) <= b;
    outputs(3571) <= not b;
    outputs(3572) <= not a;
    outputs(3573) <= not (a xor b);
    outputs(3574) <= a or b;
    outputs(3575) <= not (a xor b);
    outputs(3576) <= not (a and b);
    outputs(3577) <= a xor b;
    outputs(3578) <= a;
    outputs(3579) <= a xor b;
    outputs(3580) <= not a or b;
    outputs(3581) <= a xor b;
    outputs(3582) <= a xor b;
    outputs(3583) <= not a or b;
    outputs(3584) <= b;
    outputs(3585) <= a xor b;
    outputs(3586) <= not (a and b);
    outputs(3587) <= not a or b;
    outputs(3588) <= not (a xor b);
    outputs(3589) <= not b or a;
    outputs(3590) <= b and not a;
    outputs(3591) <= b;
    outputs(3592) <= b;
    outputs(3593) <= a or b;
    outputs(3594) <= not (a xor b);
    outputs(3595) <= b and not a;
    outputs(3596) <= not b;
    outputs(3597) <= not (a xor b);
    outputs(3598) <= a or b;
    outputs(3599) <= a and not b;
    outputs(3600) <= a and not b;
    outputs(3601) <= a;
    outputs(3602) <= not (a xor b);
    outputs(3603) <= b;
    outputs(3604) <= not (a xor b);
    outputs(3605) <= a or b;
    outputs(3606) <= not b;
    outputs(3607) <= a xor b;
    outputs(3608) <= a xor b;
    outputs(3609) <= a and b;
    outputs(3610) <= a or b;
    outputs(3611) <= not (a and b);
    outputs(3612) <= not a;
    outputs(3613) <= not (a or b);
    outputs(3614) <= a and b;
    outputs(3615) <= a or b;
    outputs(3616) <= a xor b;
    outputs(3617) <= not b;
    outputs(3618) <= a and not b;
    outputs(3619) <= not a;
    outputs(3620) <= a xor b;
    outputs(3621) <= not (a or b);
    outputs(3622) <= b and not a;
    outputs(3623) <= a and b;
    outputs(3624) <= a xor b;
    outputs(3625) <= a xor b;
    outputs(3626) <= b;
    outputs(3627) <= a xor b;
    outputs(3628) <= a or b;
    outputs(3629) <= a or b;
    outputs(3630) <= not a;
    outputs(3631) <= not (a xor b);
    outputs(3632) <= not b;
    outputs(3633) <= not (a xor b);
    outputs(3634) <= a;
    outputs(3635) <= a xor b;
    outputs(3636) <= a or b;
    outputs(3637) <= not (a xor b);
    outputs(3638) <= not (a xor b);
    outputs(3639) <= not (a xor b);
    outputs(3640) <= not (a or b);
    outputs(3641) <= not (a xor b);
    outputs(3642) <= not (a xor b);
    outputs(3643) <= not (a or b);
    outputs(3644) <= a;
    outputs(3645) <= not a;
    outputs(3646) <= a and b;
    outputs(3647) <= not (a xor b);
    outputs(3648) <= a xor b;
    outputs(3649) <= not b;
    outputs(3650) <= a or b;
    outputs(3651) <= a and b;
    outputs(3652) <= a xor b;
    outputs(3653) <= not (a xor b);
    outputs(3654) <= a;
    outputs(3655) <= a;
    outputs(3656) <= not b;
    outputs(3657) <= a xor b;
    outputs(3658) <= not b;
    outputs(3659) <= a xor b;
    outputs(3660) <= a and b;
    outputs(3661) <= not (a xor b);
    outputs(3662) <= a xor b;
    outputs(3663) <= not b;
    outputs(3664) <= not a;
    outputs(3665) <= a and not b;
    outputs(3666) <= a and b;
    outputs(3667) <= a xor b;
    outputs(3668) <= not a or b;
    outputs(3669) <= not b or a;
    outputs(3670) <= not b;
    outputs(3671) <= not a;
    outputs(3672) <= not (a or b);
    outputs(3673) <= a;
    outputs(3674) <= not b;
    outputs(3675) <= a and b;
    outputs(3676) <= not (a and b);
    outputs(3677) <= a xor b;
    outputs(3678) <= not (a xor b);
    outputs(3679) <= a and not b;
    outputs(3680) <= a;
    outputs(3681) <= a or b;
    outputs(3682) <= a xor b;
    outputs(3683) <= a;
    outputs(3684) <= a or b;
    outputs(3685) <= a xor b;
    outputs(3686) <= b;
    outputs(3687) <= not (a xor b);
    outputs(3688) <= not (a xor b);
    outputs(3689) <= b;
    outputs(3690) <= not (a xor b);
    outputs(3691) <= not b;
    outputs(3692) <= not a or b;
    outputs(3693) <= not (a and b);
    outputs(3694) <= b;
    outputs(3695) <= b;
    outputs(3696) <= not (a xor b);
    outputs(3697) <= a xor b;
    outputs(3698) <= b;
    outputs(3699) <= a xor b;
    outputs(3700) <= a or b;
    outputs(3701) <= not (a xor b);
    outputs(3702) <= not a or b;
    outputs(3703) <= a;
    outputs(3704) <= b;
    outputs(3705) <= not (a xor b);
    outputs(3706) <= a;
    outputs(3707) <= not (a xor b);
    outputs(3708) <= not b or a;
    outputs(3709) <= not (a xor b);
    outputs(3710) <= b and not a;
    outputs(3711) <= not a or b;
    outputs(3712) <= not (a xor b);
    outputs(3713) <= a or b;
    outputs(3714) <= a or b;
    outputs(3715) <= not b or a;
    outputs(3716) <= not b;
    outputs(3717) <= not b;
    outputs(3718) <= b;
    outputs(3719) <= not b;
    outputs(3720) <= a;
    outputs(3721) <= b;
    outputs(3722) <= not b;
    outputs(3723) <= not a;
    outputs(3724) <= a;
    outputs(3725) <= a;
    outputs(3726) <= b;
    outputs(3727) <= b;
    outputs(3728) <= not a;
    outputs(3729) <= not (a xor b);
    outputs(3730) <= a xor b;
    outputs(3731) <= not a or b;
    outputs(3732) <= not (a xor b);
    outputs(3733) <= a xor b;
    outputs(3734) <= a or b;
    outputs(3735) <= not (a or b);
    outputs(3736) <= not (a xor b);
    outputs(3737) <= not (a xor b);
    outputs(3738) <= a xor b;
    outputs(3739) <= not a or b;
    outputs(3740) <= not a or b;
    outputs(3741) <= not b;
    outputs(3742) <= a xor b;
    outputs(3743) <= not b;
    outputs(3744) <= a xor b;
    outputs(3745) <= not a or b;
    outputs(3746) <= a and not b;
    outputs(3747) <= a xor b;
    outputs(3748) <= not a;
    outputs(3749) <= not b or a;
    outputs(3750) <= a;
    outputs(3751) <= not (a xor b);
    outputs(3752) <= a;
    outputs(3753) <= b and not a;
    outputs(3754) <= not b;
    outputs(3755) <= not b;
    outputs(3756) <= a xor b;
    outputs(3757) <= b;
    outputs(3758) <= not a;
    outputs(3759) <= not (a xor b);
    outputs(3760) <= a;
    outputs(3761) <= not (a xor b);
    outputs(3762) <= a;
    outputs(3763) <= not b or a;
    outputs(3764) <= not a;
    outputs(3765) <= b;
    outputs(3766) <= a xor b;
    outputs(3767) <= b;
    outputs(3768) <= a xor b;
    outputs(3769) <= not (a xor b);
    outputs(3770) <= a xor b;
    outputs(3771) <= b and not a;
    outputs(3772) <= not a;
    outputs(3773) <= not (a or b);
    outputs(3774) <= not (a xor b);
    outputs(3775) <= a;
    outputs(3776) <= a xor b;
    outputs(3777) <= b and not a;
    outputs(3778) <= not a or b;
    outputs(3779) <= not a;
    outputs(3780) <= a or b;
    outputs(3781) <= a or b;
    outputs(3782) <= a;
    outputs(3783) <= not a or b;
    outputs(3784) <= a xor b;
    outputs(3785) <= not (a xor b);
    outputs(3786) <= not a or b;
    outputs(3787) <= a xor b;
    outputs(3788) <= a or b;
    outputs(3789) <= a;
    outputs(3790) <= a;
    outputs(3791) <= b;
    outputs(3792) <= not (a and b);
    outputs(3793) <= not a;
    outputs(3794) <= a xor b;
    outputs(3795) <= not b;
    outputs(3796) <= not (a xor b);
    outputs(3797) <= a and not b;
    outputs(3798) <= not b or a;
    outputs(3799) <= b;
    outputs(3800) <= not (a xor b);
    outputs(3801) <= a;
    outputs(3802) <= a;
    outputs(3803) <= a and b;
    outputs(3804) <= a and b;
    outputs(3805) <= not a;
    outputs(3806) <= not a;
    outputs(3807) <= a;
    outputs(3808) <= a xor b;
    outputs(3809) <= a;
    outputs(3810) <= not b;
    outputs(3811) <= b;
    outputs(3812) <= a xor b;
    outputs(3813) <= not (a xor b);
    outputs(3814) <= not b;
    outputs(3815) <= not (a and b);
    outputs(3816) <= not a;
    outputs(3817) <= b;
    outputs(3818) <= not a;
    outputs(3819) <= not b;
    outputs(3820) <= not b;
    outputs(3821) <= not a;
    outputs(3822) <= not (a and b);
    outputs(3823) <= a and not b;
    outputs(3824) <= b;
    outputs(3825) <= not a;
    outputs(3826) <= a xor b;
    outputs(3827) <= a;
    outputs(3828) <= not b;
    outputs(3829) <= not b;
    outputs(3830) <= a xor b;
    outputs(3831) <= a and b;
    outputs(3832) <= not b;
    outputs(3833) <= not (a xor b);
    outputs(3834) <= not a;
    outputs(3835) <= not (a xor b);
    outputs(3836) <= a;
    outputs(3837) <= b;
    outputs(3838) <= a xor b;
    outputs(3839) <= a and b;
    outputs(3840) <= not (a xor b);
    outputs(3841) <= not a;
    outputs(3842) <= a;
    outputs(3843) <= a;
    outputs(3844) <= a xor b;
    outputs(3845) <= not a or b;
    outputs(3846) <= b and not a;
    outputs(3847) <= a;
    outputs(3848) <= not b;
    outputs(3849) <= not (a or b);
    outputs(3850) <= not (a and b);
    outputs(3851) <= not (a xor b);
    outputs(3852) <= not (a xor b);
    outputs(3853) <= not b;
    outputs(3854) <= not (a xor b);
    outputs(3855) <= not a;
    outputs(3856) <= a xor b;
    outputs(3857) <= not b;
    outputs(3858) <= not (a and b);
    outputs(3859) <= a;
    outputs(3860) <= b and not a;
    outputs(3861) <= not (a xor b);
    outputs(3862) <= not a or b;
    outputs(3863) <= a;
    outputs(3864) <= a and b;
    outputs(3865) <= a and not b;
    outputs(3866) <= not b;
    outputs(3867) <= a or b;
    outputs(3868) <= not b;
    outputs(3869) <= not (a xor b);
    outputs(3870) <= b and not a;
    outputs(3871) <= a xor b;
    outputs(3872) <= not a;
    outputs(3873) <= b;
    outputs(3874) <= a xor b;
    outputs(3875) <= not b or a;
    outputs(3876) <= not (a xor b);
    outputs(3877) <= b and not a;
    outputs(3878) <= not b or a;
    outputs(3879) <= not a;
    outputs(3880) <= not (a xor b);
    outputs(3881) <= not (a xor b);
    outputs(3882) <= not (a xor b);
    outputs(3883) <= not (a or b);
    outputs(3884) <= not (a xor b);
    outputs(3885) <= b;
    outputs(3886) <= not (a xor b);
    outputs(3887) <= not b;
    outputs(3888) <= not (a and b);
    outputs(3889) <= a xor b;
    outputs(3890) <= a;
    outputs(3891) <= not (a xor b);
    outputs(3892) <= a and b;
    outputs(3893) <= not (a xor b);
    outputs(3894) <= a xor b;
    outputs(3895) <= a;
    outputs(3896) <= b;
    outputs(3897) <= a and not b;
    outputs(3898) <= a xor b;
    outputs(3899) <= not (a and b);
    outputs(3900) <= a or b;
    outputs(3901) <= not a;
    outputs(3902) <= b and not a;
    outputs(3903) <= not (a xor b);
    outputs(3904) <= a xor b;
    outputs(3905) <= not (a xor b);
    outputs(3906) <= not (a xor b);
    outputs(3907) <= not (a xor b);
    outputs(3908) <= b;
    outputs(3909) <= not b;
    outputs(3910) <= a;
    outputs(3911) <= b;
    outputs(3912) <= not (a and b);
    outputs(3913) <= a xor b;
    outputs(3914) <= b;
    outputs(3915) <= a xor b;
    outputs(3916) <= not (a xor b);
    outputs(3917) <= a xor b;
    outputs(3918) <= a xor b;
    outputs(3919) <= a xor b;
    outputs(3920) <= a;
    outputs(3921) <= not (a xor b);
    outputs(3922) <= not (a xor b);
    outputs(3923) <= not (a xor b);
    outputs(3924) <= a;
    outputs(3925) <= not (a or b);
    outputs(3926) <= a xor b;
    outputs(3927) <= not (a or b);
    outputs(3928) <= not a or b;
    outputs(3929) <= a xor b;
    outputs(3930) <= not (a or b);
    outputs(3931) <= not (a xor b);
    outputs(3932) <= not (a xor b);
    outputs(3933) <= not b;
    outputs(3934) <= b;
    outputs(3935) <= a xor b;
    outputs(3936) <= a;
    outputs(3937) <= a and not b;
    outputs(3938) <= not a;
    outputs(3939) <= not b or a;
    outputs(3940) <= a;
    outputs(3941) <= not b;
    outputs(3942) <= not (a xor b);
    outputs(3943) <= not (a xor b);
    outputs(3944) <= b;
    outputs(3945) <= not a or b;
    outputs(3946) <= not b;
    outputs(3947) <= not b;
    outputs(3948) <= not a;
    outputs(3949) <= not (a and b);
    outputs(3950) <= a and b;
    outputs(3951) <= a;
    outputs(3952) <= not b;
    outputs(3953) <= not b;
    outputs(3954) <= b;
    outputs(3955) <= a;
    outputs(3956) <= a xor b;
    outputs(3957) <= not b;
    outputs(3958) <= not a;
    outputs(3959) <= a and not b;
    outputs(3960) <= a xor b;
    outputs(3961) <= not (a and b);
    outputs(3962) <= a xor b;
    outputs(3963) <= b and not a;
    outputs(3964) <= not a;
    outputs(3965) <= not (a xor b);
    outputs(3966) <= not b;
    outputs(3967) <= not b;
    outputs(3968) <= not b;
    outputs(3969) <= not b;
    outputs(3970) <= not (a xor b);
    outputs(3971) <= a and b;
    outputs(3972) <= a xor b;
    outputs(3973) <= not (a xor b);
    outputs(3974) <= not (a or b);
    outputs(3975) <= not b;
    outputs(3976) <= b and not a;
    outputs(3977) <= a and not b;
    outputs(3978) <= not (a xor b);
    outputs(3979) <= a;
    outputs(3980) <= a;
    outputs(3981) <= not a;
    outputs(3982) <= not a;
    outputs(3983) <= not a;
    outputs(3984) <= a;
    outputs(3985) <= a and not b;
    outputs(3986) <= a xor b;
    outputs(3987) <= a xor b;
    outputs(3988) <= a xor b;
    outputs(3989) <= a;
    outputs(3990) <= a and b;
    outputs(3991) <= not (a and b);
    outputs(3992) <= not (a xor b);
    outputs(3993) <= not a;
    outputs(3994) <= not (a and b);
    outputs(3995) <= not a;
    outputs(3996) <= not a;
    outputs(3997) <= b and not a;
    outputs(3998) <= b and not a;
    outputs(3999) <= b;
    outputs(4000) <= not (a xor b);
    outputs(4001) <= not a or b;
    outputs(4002) <= a xor b;
    outputs(4003) <= not b;
    outputs(4004) <= not (a xor b);
    outputs(4005) <= not (a or b);
    outputs(4006) <= not a or b;
    outputs(4007) <= not b;
    outputs(4008) <= not (a xor b);
    outputs(4009) <= not b;
    outputs(4010) <= a xor b;
    outputs(4011) <= a;
    outputs(4012) <= not a or b;
    outputs(4013) <= a xor b;
    outputs(4014) <= a;
    outputs(4015) <= a;
    outputs(4016) <= a xor b;
    outputs(4017) <= a and not b;
    outputs(4018) <= b;
    outputs(4019) <= a;
    outputs(4020) <= b;
    outputs(4021) <= a xor b;
    outputs(4022) <= a and b;
    outputs(4023) <= not b;
    outputs(4024) <= not a;
    outputs(4025) <= a;
    outputs(4026) <= not (a xor b);
    outputs(4027) <= not (a and b);
    outputs(4028) <= a;
    outputs(4029) <= not (a xor b);
    outputs(4030) <= a xor b;
    outputs(4031) <= a;
    outputs(4032) <= not b;
    outputs(4033) <= a xor b;
    outputs(4034) <= not a;
    outputs(4035) <= a xor b;
    outputs(4036) <= not a or b;
    outputs(4037) <= a xor b;
    outputs(4038) <= a xor b;
    outputs(4039) <= not a;
    outputs(4040) <= not (a and b);
    outputs(4041) <= b and not a;
    outputs(4042) <= a and not b;
    outputs(4043) <= not b or a;
    outputs(4044) <= a or b;
    outputs(4045) <= a;
    outputs(4046) <= not b;
    outputs(4047) <= not (a xor b);
    outputs(4048) <= b;
    outputs(4049) <= not (a and b);
    outputs(4050) <= not (a and b);
    outputs(4051) <= a xor b;
    outputs(4052) <= a and b;
    outputs(4053) <= a xor b;
    outputs(4054) <= a xor b;
    outputs(4055) <= a;
    outputs(4056) <= not (a xor b);
    outputs(4057) <= not b;
    outputs(4058) <= not (a xor b);
    outputs(4059) <= not b;
    outputs(4060) <= not a;
    outputs(4061) <= not a;
    outputs(4062) <= a or b;
    outputs(4063) <= b;
    outputs(4064) <= not b;
    outputs(4065) <= not (a or b);
    outputs(4066) <= a;
    outputs(4067) <= not a;
    outputs(4068) <= a;
    outputs(4069) <= not (a and b);
    outputs(4070) <= a xor b;
    outputs(4071) <= not (a xor b);
    outputs(4072) <= b;
    outputs(4073) <= not a;
    outputs(4074) <= not (a xor b);
    outputs(4075) <= b;
    outputs(4076) <= not b;
    outputs(4077) <= not (a xor b);
    outputs(4078) <= b and not a;
    outputs(4079) <= b;
    outputs(4080) <= a and not b;
    outputs(4081) <= not (a xor b);
    outputs(4082) <= not (a xor b);
    outputs(4083) <= a;
    outputs(4084) <= a and b;
    outputs(4085) <= b;
    outputs(4086) <= not a;
    outputs(4087) <= a and not b;
    outputs(4088) <= b;
    outputs(4089) <= not b or a;
    outputs(4090) <= a xor b;
    outputs(4091) <= not b;
    outputs(4092) <= not a;
    outputs(4093) <= not b;
    outputs(4094) <= a;
    outputs(4095) <= a xor b;
    outputs(4096) <= b;
    outputs(4097) <= not b or a;
    outputs(4098) <= b;
    outputs(4099) <= not b;
    outputs(4100) <= not b or a;
    outputs(4101) <= not (a xor b);
    outputs(4102) <= not a;
    outputs(4103) <= a;
    outputs(4104) <= a and not b;
    outputs(4105) <= a;
    outputs(4106) <= not b;
    outputs(4107) <= b;
    outputs(4108) <= a;
    outputs(4109) <= b;
    outputs(4110) <= not a or b;
    outputs(4111) <= not (a and b);
    outputs(4112) <= a or b;
    outputs(4113) <= not a or b;
    outputs(4114) <= a xor b;
    outputs(4115) <= not a or b;
    outputs(4116) <= a;
    outputs(4117) <= not (a xor b);
    outputs(4118) <= not (a xor b);
    outputs(4119) <= a;
    outputs(4120) <= a xor b;
    outputs(4121) <= not b;
    outputs(4122) <= a xor b;
    outputs(4123) <= b;
    outputs(4124) <= not b;
    outputs(4125) <= not (a or b);
    outputs(4126) <= a xor b;
    outputs(4127) <= not (a or b);
    outputs(4128) <= b;
    outputs(4129) <= not (a xor b);
    outputs(4130) <= not b;
    outputs(4131) <= not (a xor b);
    outputs(4132) <= not b;
    outputs(4133) <= not b;
    outputs(4134) <= not a;
    outputs(4135) <= a or b;
    outputs(4136) <= a xor b;
    outputs(4137) <= not b;
    outputs(4138) <= b;
    outputs(4139) <= not (a xor b);
    outputs(4140) <= a and b;
    outputs(4141) <= a xor b;
    outputs(4142) <= a xor b;
    outputs(4143) <= not b;
    outputs(4144) <= not a;
    outputs(4145) <= b;
    outputs(4146) <= a;
    outputs(4147) <= a xor b;
    outputs(4148) <= a and b;
    outputs(4149) <= not (a xor b);
    outputs(4150) <= not (a and b);
    outputs(4151) <= not (a xor b);
    outputs(4152) <= not (a and b);
    outputs(4153) <= not b;
    outputs(4154) <= b;
    outputs(4155) <= not a;
    outputs(4156) <= not (a xor b);
    outputs(4157) <= not (a xor b);
    outputs(4158) <= not (a xor b);
    outputs(4159) <= not b;
    outputs(4160) <= b;
    outputs(4161) <= not a or b;
    outputs(4162) <= not a;
    outputs(4163) <= b;
    outputs(4164) <= a xor b;
    outputs(4165) <= a xor b;
    outputs(4166) <= a xor b;
    outputs(4167) <= a xor b;
    outputs(4168) <= a xor b;
    outputs(4169) <= not a;
    outputs(4170) <= not (a xor b);
    outputs(4171) <= a xor b;
    outputs(4172) <= b and not a;
    outputs(4173) <= a;
    outputs(4174) <= a xor b;
    outputs(4175) <= not (a or b);
    outputs(4176) <= not a;
    outputs(4177) <= not b;
    outputs(4178) <= not (a or b);
    outputs(4179) <= a xor b;
    outputs(4180) <= a;
    outputs(4181) <= a;
    outputs(4182) <= a and not b;
    outputs(4183) <= a or b;
    outputs(4184) <= a xor b;
    outputs(4185) <= b and not a;
    outputs(4186) <= a;
    outputs(4187) <= a xor b;
    outputs(4188) <= not (a xor b);
    outputs(4189) <= not (a xor b);
    outputs(4190) <= a;
    outputs(4191) <= not (a xor b);
    outputs(4192) <= b;
    outputs(4193) <= a and b;
    outputs(4194) <= a xor b;
    outputs(4195) <= not b;
    outputs(4196) <= not a;
    outputs(4197) <= a xor b;
    outputs(4198) <= not (a or b);
    outputs(4199) <= a;
    outputs(4200) <= not (a xor b);
    outputs(4201) <= a xor b;
    outputs(4202) <= not a;
    outputs(4203) <= a xor b;
    outputs(4204) <= b;
    outputs(4205) <= a xor b;
    outputs(4206) <= not a;
    outputs(4207) <= not (a xor b);
    outputs(4208) <= not (a xor b);
    outputs(4209) <= a xor b;
    outputs(4210) <= b;
    outputs(4211) <= a and not b;
    outputs(4212) <= not a;
    outputs(4213) <= a xor b;
    outputs(4214) <= not b;
    outputs(4215) <= not (a xor b);
    outputs(4216) <= not (a xor b);
    outputs(4217) <= a xor b;
    outputs(4218) <= not (a xor b);
    outputs(4219) <= not (a xor b);
    outputs(4220) <= not b or a;
    outputs(4221) <= not a or b;
    outputs(4222) <= not a;
    outputs(4223) <= not a;
    outputs(4224) <= not (a xor b);
    outputs(4225) <= b;
    outputs(4226) <= not (a xor b);
    outputs(4227) <= b and not a;
    outputs(4228) <= a and not b;
    outputs(4229) <= not a;
    outputs(4230) <= not a or b;
    outputs(4231) <= a and not b;
    outputs(4232) <= not b or a;
    outputs(4233) <= not a;
    outputs(4234) <= a;
    outputs(4235) <= not a;
    outputs(4236) <= not a;
    outputs(4237) <= not a;
    outputs(4238) <= a or b;
    outputs(4239) <= a xor b;
    outputs(4240) <= a;
    outputs(4241) <= not a or b;
    outputs(4242) <= not (a xor b);
    outputs(4243) <= a or b;
    outputs(4244) <= a;
    outputs(4245) <= not (a xor b);
    outputs(4246) <= not (a xor b);
    outputs(4247) <= a xor b;
    outputs(4248) <= not (a xor b);
    outputs(4249) <= a;
    outputs(4250) <= not a;
    outputs(4251) <= a xor b;
    outputs(4252) <= b and not a;
    outputs(4253) <= a xor b;
    outputs(4254) <= not b or a;
    outputs(4255) <= not a;
    outputs(4256) <= not a or b;
    outputs(4257) <= not b;
    outputs(4258) <= not (a xor b);
    outputs(4259) <= not b;
    outputs(4260) <= not (a and b);
    outputs(4261) <= not b;
    outputs(4262) <= not (a xor b);
    outputs(4263) <= b;
    outputs(4264) <= not (a and b);
    outputs(4265) <= not (a xor b);
    outputs(4266) <= a xor b;
    outputs(4267) <= not (a xor b);
    outputs(4268) <= a;
    outputs(4269) <= not a or b;
    outputs(4270) <= a xor b;
    outputs(4271) <= not b or a;
    outputs(4272) <= b;
    outputs(4273) <= not a;
    outputs(4274) <= a xor b;
    outputs(4275) <= not b;
    outputs(4276) <= b;
    outputs(4277) <= not a or b;
    outputs(4278) <= a xor b;
    outputs(4279) <= a xor b;
    outputs(4280) <= b;
    outputs(4281) <= not b;
    outputs(4282) <= not (a and b);
    outputs(4283) <= a and not b;
    outputs(4284) <= b;
    outputs(4285) <= not (a xor b);
    outputs(4286) <= not b;
    outputs(4287) <= b;
    outputs(4288) <= b;
    outputs(4289) <= not (a xor b);
    outputs(4290) <= a xor b;
    outputs(4291) <= not (a xor b);
    outputs(4292) <= not (a xor b);
    outputs(4293) <= not b;
    outputs(4294) <= not (a xor b);
    outputs(4295) <= not (a xor b);
    outputs(4296) <= not (a or b);
    outputs(4297) <= a xor b;
    outputs(4298) <= a and not b;
    outputs(4299) <= not (a xor b);
    outputs(4300) <= not a;
    outputs(4301) <= a xor b;
    outputs(4302) <= b;
    outputs(4303) <= a;
    outputs(4304) <= not (a xor b);
    outputs(4305) <= a;
    outputs(4306) <= a xor b;
    outputs(4307) <= not (a xor b);
    outputs(4308) <= not b;
    outputs(4309) <= a and b;
    outputs(4310) <= a xor b;
    outputs(4311) <= a;
    outputs(4312) <= not b;
    outputs(4313) <= not b or a;
    outputs(4314) <= b;
    outputs(4315) <= not b;
    outputs(4316) <= a xor b;
    outputs(4317) <= a xor b;
    outputs(4318) <= not a or b;
    outputs(4319) <= not (a xor b);
    outputs(4320) <= not (a xor b);
    outputs(4321) <= a and b;
    outputs(4322) <= a xor b;
    outputs(4323) <= not (a and b);
    outputs(4324) <= not (a or b);
    outputs(4325) <= not b;
    outputs(4326) <= not (a or b);
    outputs(4327) <= a;
    outputs(4328) <= not (a and b);
    outputs(4329) <= a and b;
    outputs(4330) <= not b;
    outputs(4331) <= b;
    outputs(4332) <= b;
    outputs(4333) <= not b or a;
    outputs(4334) <= a;
    outputs(4335) <= b and not a;
    outputs(4336) <= b;
    outputs(4337) <= a xor b;
    outputs(4338) <= a xor b;
    outputs(4339) <= a xor b;
    outputs(4340) <= a xor b;
    outputs(4341) <= not (a or b);
    outputs(4342) <= not a or b;
    outputs(4343) <= a xor b;
    outputs(4344) <= not (a xor b);
    outputs(4345) <= a and b;
    outputs(4346) <= not b;
    outputs(4347) <= a and not b;
    outputs(4348) <= a and not b;
    outputs(4349) <= not (a and b);
    outputs(4350) <= b;
    outputs(4351) <= a xor b;
    outputs(4352) <= not a;
    outputs(4353) <= b;
    outputs(4354) <= a xor b;
    outputs(4355) <= not (a xor b);
    outputs(4356) <= not a or b;
    outputs(4357) <= not (a and b);
    outputs(4358) <= b;
    outputs(4359) <= a xor b;
    outputs(4360) <= not (a or b);
    outputs(4361) <= not a;
    outputs(4362) <= not b;
    outputs(4363) <= not (a and b);
    outputs(4364) <= a xor b;
    outputs(4365) <= not (a xor b);
    outputs(4366) <= a;
    outputs(4367) <= a xor b;
    outputs(4368) <= not (a xor b);
    outputs(4369) <= a xor b;
    outputs(4370) <= a xor b;
    outputs(4371) <= not (a xor b);
    outputs(4372) <= a xor b;
    outputs(4373) <= b and not a;
    outputs(4374) <= a;
    outputs(4375) <= b;
    outputs(4376) <= not a;
    outputs(4377) <= not b or a;
    outputs(4378) <= a;
    outputs(4379) <= a xor b;
    outputs(4380) <= b and not a;
    outputs(4381) <= not (a xor b);
    outputs(4382) <= a;
    outputs(4383) <= not a;
    outputs(4384) <= a and b;
    outputs(4385) <= a;
    outputs(4386) <= a xor b;
    outputs(4387) <= not (a xor b);
    outputs(4388) <= not (a and b);
    outputs(4389) <= a;
    outputs(4390) <= not b;
    outputs(4391) <= not (a xor b);
    outputs(4392) <= not (a xor b);
    outputs(4393) <= a xor b;
    outputs(4394) <= not (a xor b);
    outputs(4395) <= not b;
    outputs(4396) <= not a or b;
    outputs(4397) <= a and b;
    outputs(4398) <= not b;
    outputs(4399) <= b;
    outputs(4400) <= not a or b;
    outputs(4401) <= not (a and b);
    outputs(4402) <= not a;
    outputs(4403) <= b and not a;
    outputs(4404) <= a xor b;
    outputs(4405) <= a xor b;
    outputs(4406) <= a;
    outputs(4407) <= b and not a;
    outputs(4408) <= a and b;
    outputs(4409) <= not (a and b);
    outputs(4410) <= a;
    outputs(4411) <= not a;
    outputs(4412) <= not a;
    outputs(4413) <= b;
    outputs(4414) <= not a;
    outputs(4415) <= b and not a;
    outputs(4416) <= not (a xor b);
    outputs(4417) <= a or b;
    outputs(4418) <= b;
    outputs(4419) <= not a;
    outputs(4420) <= b and not a;
    outputs(4421) <= not (a or b);
    outputs(4422) <= not (a and b);
    outputs(4423) <= not (a xor b);
    outputs(4424) <= not a;
    outputs(4425) <= not (a xor b);
    outputs(4426) <= not (a xor b);
    outputs(4427) <= a and not b;
    outputs(4428) <= not a;
    outputs(4429) <= b and not a;
    outputs(4430) <= a xor b;
    outputs(4431) <= a xor b;
    outputs(4432) <= not (a and b);
    outputs(4433) <= not (a xor b);
    outputs(4434) <= not (a or b);
    outputs(4435) <= not a;
    outputs(4436) <= b and not a;
    outputs(4437) <= not a;
    outputs(4438) <= b;
    outputs(4439) <= not (a xor b);
    outputs(4440) <= not a;
    outputs(4441) <= not (a xor b);
    outputs(4442) <= not b or a;
    outputs(4443) <= a;
    outputs(4444) <= a and not b;
    outputs(4445) <= a xor b;
    outputs(4446) <= not b or a;
    outputs(4447) <= not (a or b);
    outputs(4448) <= not (a xor b);
    outputs(4449) <= not b;
    outputs(4450) <= not (a xor b);
    outputs(4451) <= a or b;
    outputs(4452) <= a xor b;
    outputs(4453) <= a or b;
    outputs(4454) <= not b;
    outputs(4455) <= a;
    outputs(4456) <= not (a xor b);
    outputs(4457) <= not a;
    outputs(4458) <= not (a or b);
    outputs(4459) <= not b;
    outputs(4460) <= a xor b;
    outputs(4461) <= a xor b;
    outputs(4462) <= a xor b;
    outputs(4463) <= not b;
    outputs(4464) <= not b or a;
    outputs(4465) <= b;
    outputs(4466) <= a;
    outputs(4467) <= a xor b;
    outputs(4468) <= not a or b;
    outputs(4469) <= a;
    outputs(4470) <= not b;
    outputs(4471) <= not (a and b);
    outputs(4472) <= not (a xor b);
    outputs(4473) <= a xor b;
    outputs(4474) <= not (a xor b);
    outputs(4475) <= not a;
    outputs(4476) <= a xor b;
    outputs(4477) <= not (a xor b);
    outputs(4478) <= not b;
    outputs(4479) <= not b;
    outputs(4480) <= not a or b;
    outputs(4481) <= not a;
    outputs(4482) <= not (a xor b);
    outputs(4483) <= b;
    outputs(4484) <= a and not b;
    outputs(4485) <= not b or a;
    outputs(4486) <= not b;
    outputs(4487) <= b;
    outputs(4488) <= a or b;
    outputs(4489) <= b;
    outputs(4490) <= not (a xor b);
    outputs(4491) <= b and not a;
    outputs(4492) <= not b;
    outputs(4493) <= not b;
    outputs(4494) <= not a;
    outputs(4495) <= a xor b;
    outputs(4496) <= not a;
    outputs(4497) <= b and not a;
    outputs(4498) <= not b;
    outputs(4499) <= a;
    outputs(4500) <= b;
    outputs(4501) <= a xor b;
    outputs(4502) <= a;
    outputs(4503) <= not b or a;
    outputs(4504) <= a xor b;
    outputs(4505) <= not b;
    outputs(4506) <= not a;
    outputs(4507) <= not a;
    outputs(4508) <= not (a xor b);
    outputs(4509) <= not (a and b);
    outputs(4510) <= not (a xor b);
    outputs(4511) <= a;
    outputs(4512) <= a xor b;
    outputs(4513) <= a and not b;
    outputs(4514) <= a and not b;
    outputs(4515) <= not a;
    outputs(4516) <= b;
    outputs(4517) <= a xor b;
    outputs(4518) <= not (a xor b);
    outputs(4519) <= b;
    outputs(4520) <= a;
    outputs(4521) <= not (a xor b);
    outputs(4522) <= not a;
    outputs(4523) <= not b;
    outputs(4524) <= a;
    outputs(4525) <= not (a or b);
    outputs(4526) <= not a;
    outputs(4527) <= not (a or b);
    outputs(4528) <= a xor b;
    outputs(4529) <= a;
    outputs(4530) <= not (a xor b);
    outputs(4531) <= not a;
    outputs(4532) <= not (a xor b);
    outputs(4533) <= a and not b;
    outputs(4534) <= a;
    outputs(4535) <= a xor b;
    outputs(4536) <= not (a or b);
    outputs(4537) <= a xor b;
    outputs(4538) <= b and not a;
    outputs(4539) <= not a or b;
    outputs(4540) <= b;
    outputs(4541) <= b and not a;
    outputs(4542) <= a xor b;
    outputs(4543) <= not a or b;
    outputs(4544) <= b;
    outputs(4545) <= not a or b;
    outputs(4546) <= not b;
    outputs(4547) <= b;
    outputs(4548) <= a or b;
    outputs(4549) <= not (a xor b);
    outputs(4550) <= a xor b;
    outputs(4551) <= a xor b;
    outputs(4552) <= b;
    outputs(4553) <= b and not a;
    outputs(4554) <= not a;
    outputs(4555) <= not b;
    outputs(4556) <= a;
    outputs(4557) <= a xor b;
    outputs(4558) <= a xor b;
    outputs(4559) <= b and not a;
    outputs(4560) <= a xor b;
    outputs(4561) <= not (a xor b);
    outputs(4562) <= not (a xor b);
    outputs(4563) <= a or b;
    outputs(4564) <= not (a xor b);
    outputs(4565) <= a or b;
    outputs(4566) <= b and not a;
    outputs(4567) <= a;
    outputs(4568) <= a and b;
    outputs(4569) <= not (a and b);
    outputs(4570) <= not (a xor b);
    outputs(4571) <= a;
    outputs(4572) <= not (a xor b);
    outputs(4573) <= not b or a;
    outputs(4574) <= not b;
    outputs(4575) <= a and not b;
    outputs(4576) <= not a;
    outputs(4577) <= a;
    outputs(4578) <= not (a xor b);
    outputs(4579) <= b;
    outputs(4580) <= not (a and b);
    outputs(4581) <= not b;
    outputs(4582) <= not (a and b);
    outputs(4583) <= a and not b;
    outputs(4584) <= a xor b;
    outputs(4585) <= b;
    outputs(4586) <= a xor b;
    outputs(4587) <= not (a or b);
    outputs(4588) <= not a;
    outputs(4589) <= a xor b;
    outputs(4590) <= a and b;
    outputs(4591) <= b;
    outputs(4592) <= a xor b;
    outputs(4593) <= not (a xor b);
    outputs(4594) <= not (a xor b);
    outputs(4595) <= not (a xor b);
    outputs(4596) <= b;
    outputs(4597) <= not (a xor b);
    outputs(4598) <= a and b;
    outputs(4599) <= not b;
    outputs(4600) <= not b or a;
    outputs(4601) <= a or b;
    outputs(4602) <= not (a xor b);
    outputs(4603) <= not (a xor b);
    outputs(4604) <= a;
    outputs(4605) <= b;
    outputs(4606) <= not (a xor b);
    outputs(4607) <= a;
    outputs(4608) <= a xor b;
    outputs(4609) <= not b;
    outputs(4610) <= a and b;
    outputs(4611) <= a;
    outputs(4612) <= a xor b;
    outputs(4613) <= not a;
    outputs(4614) <= a;
    outputs(4615) <= not b;
    outputs(4616) <= not a;
    outputs(4617) <= b;
    outputs(4618) <= not (a xor b);
    outputs(4619) <= a;
    outputs(4620) <= not a;
    outputs(4621) <= a xor b;
    outputs(4622) <= a;
    outputs(4623) <= b;
    outputs(4624) <= not b;
    outputs(4625) <= not a or b;
    outputs(4626) <= not (a or b);
    outputs(4627) <= b;
    outputs(4628) <= not (a or b);
    outputs(4629) <= not b;
    outputs(4630) <= a and b;
    outputs(4631) <= not a or b;
    outputs(4632) <= not (a xor b);
    outputs(4633) <= b;
    outputs(4634) <= not (a xor b);
    outputs(4635) <= not a;
    outputs(4636) <= not b;
    outputs(4637) <= a and b;
    outputs(4638) <= not a;
    outputs(4639) <= not (a or b);
    outputs(4640) <= not b or a;
    outputs(4641) <= a xor b;
    outputs(4642) <= not (a xor b);
    outputs(4643) <= not b or a;
    outputs(4644) <= a;
    outputs(4645) <= not (a or b);
    outputs(4646) <= not (a or b);
    outputs(4647) <= b;
    outputs(4648) <= a xor b;
    outputs(4649) <= not a;
    outputs(4650) <= a and b;
    outputs(4651) <= b;
    outputs(4652) <= not a;
    outputs(4653) <= not a or b;
    outputs(4654) <= not a;
    outputs(4655) <= a xor b;
    outputs(4656) <= a xor b;
    outputs(4657) <= not (a or b);
    outputs(4658) <= not (a xor b);
    outputs(4659) <= a xor b;
    outputs(4660) <= not b;
    outputs(4661) <= a xor b;
    outputs(4662) <= a;
    outputs(4663) <= a xor b;
    outputs(4664) <= a xor b;
    outputs(4665) <= a xor b;
    outputs(4666) <= not a;
    outputs(4667) <= a;
    outputs(4668) <= not (a xor b);
    outputs(4669) <= not (a xor b);
    outputs(4670) <= a;
    outputs(4671) <= not (a xor b);
    outputs(4672) <= not (a or b);
    outputs(4673) <= a xor b;
    outputs(4674) <= b and not a;
    outputs(4675) <= a xor b;
    outputs(4676) <= not (a xor b);
    outputs(4677) <= not b;
    outputs(4678) <= not (a and b);
    outputs(4679) <= a xor b;
    outputs(4680) <= a;
    outputs(4681) <= a xor b;
    outputs(4682) <= not b or a;
    outputs(4683) <= not a or b;
    outputs(4684) <= a xor b;
    outputs(4685) <= not (a xor b);
    outputs(4686) <= not (a and b);
    outputs(4687) <= a xor b;
    outputs(4688) <= a;
    outputs(4689) <= not (a and b);
    outputs(4690) <= a and b;
    outputs(4691) <= a xor b;
    outputs(4692) <= a;
    outputs(4693) <= not b or a;
    outputs(4694) <= not (a and b);
    outputs(4695) <= a;
    outputs(4696) <= not b;
    outputs(4697) <= b and not a;
    outputs(4698) <= a and b;
    outputs(4699) <= not (a xor b);
    outputs(4700) <= a and b;
    outputs(4701) <= not b;
    outputs(4702) <= b;
    outputs(4703) <= not (a or b);
    outputs(4704) <= a xor b;
    outputs(4705) <= a;
    outputs(4706) <= a xor b;
    outputs(4707) <= a xor b;
    outputs(4708) <= not b;
    outputs(4709) <= a xor b;
    outputs(4710) <= not b;
    outputs(4711) <= a or b;
    outputs(4712) <= not a;
    outputs(4713) <= a or b;
    outputs(4714) <= b and not a;
    outputs(4715) <= a;
    outputs(4716) <= b and not a;
    outputs(4717) <= b;
    outputs(4718) <= not (a xor b);
    outputs(4719) <= not a;
    outputs(4720) <= not b or a;
    outputs(4721) <= not b;
    outputs(4722) <= not (a or b);
    outputs(4723) <= not (a xor b);
    outputs(4724) <= not (a xor b);
    outputs(4725) <= a;
    outputs(4726) <= a;
    outputs(4727) <= not (a or b);
    outputs(4728) <= not b;
    outputs(4729) <= a xor b;
    outputs(4730) <= not a or b;
    outputs(4731) <= a xor b;
    outputs(4732) <= not a;
    outputs(4733) <= not (a xor b);
    outputs(4734) <= a xor b;
    outputs(4735) <= not b;
    outputs(4736) <= a;
    outputs(4737) <= not b;
    outputs(4738) <= not (a xor b);
    outputs(4739) <= a;
    outputs(4740) <= not b;
    outputs(4741) <= not b or a;
    outputs(4742) <= b and not a;
    outputs(4743) <= not b;
    outputs(4744) <= not b;
    outputs(4745) <= a;
    outputs(4746) <= a xor b;
    outputs(4747) <= b;
    outputs(4748) <= not (a xor b);
    outputs(4749) <= not a;
    outputs(4750) <= a xor b;
    outputs(4751) <= a;
    outputs(4752) <= b;
    outputs(4753) <= not b or a;
    outputs(4754) <= not (a xor b);
    outputs(4755) <= not (a xor b);
    outputs(4756) <= b and not a;
    outputs(4757) <= not a or b;
    outputs(4758) <= a;
    outputs(4759) <= not b;
    outputs(4760) <= not (a xor b);
    outputs(4761) <= a;
    outputs(4762) <= not b;
    outputs(4763) <= a;
    outputs(4764) <= a xor b;
    outputs(4765) <= not (a xor b);
    outputs(4766) <= a;
    outputs(4767) <= not (a xor b);
    outputs(4768) <= not (a xor b);
    outputs(4769) <= b;
    outputs(4770) <= not (a xor b);
    outputs(4771) <= a xor b;
    outputs(4772) <= a and not b;
    outputs(4773) <= not (a xor b);
    outputs(4774) <= a xor b;
    outputs(4775) <= a xor b;
    outputs(4776) <= not (a xor b);
    outputs(4777) <= a xor b;
    outputs(4778) <= a;
    outputs(4779) <= b;
    outputs(4780) <= not b;
    outputs(4781) <= b;
    outputs(4782) <= a xor b;
    outputs(4783) <= not (a xor b);
    outputs(4784) <= not (a xor b);
    outputs(4785) <= a;
    outputs(4786) <= not (a or b);
    outputs(4787) <= a xor b;
    outputs(4788) <= not (a xor b);
    outputs(4789) <= a or b;
    outputs(4790) <= not (a or b);
    outputs(4791) <= not (a xor b);
    outputs(4792) <= b;
    outputs(4793) <= a xor b;
    outputs(4794) <= not b or a;
    outputs(4795) <= not b or a;
    outputs(4796) <= not (a xor b);
    outputs(4797) <= not (a xor b);
    outputs(4798) <= a or b;
    outputs(4799) <= not b or a;
    outputs(4800) <= b;
    outputs(4801) <= not a;
    outputs(4802) <= a xor b;
    outputs(4803) <= not (a and b);
    outputs(4804) <= b and not a;
    outputs(4805) <= not b;
    outputs(4806) <= b;
    outputs(4807) <= not b or a;
    outputs(4808) <= not a;
    outputs(4809) <= not (a or b);
    outputs(4810) <= a xor b;
    outputs(4811) <= not a;
    outputs(4812) <= a xor b;
    outputs(4813) <= a and b;
    outputs(4814) <= a xor b;
    outputs(4815) <= not a or b;
    outputs(4816) <= not (a or b);
    outputs(4817) <= a and not b;
    outputs(4818) <= not b;
    outputs(4819) <= b;
    outputs(4820) <= a xor b;
    outputs(4821) <= not (a xor b);
    outputs(4822) <= not a;
    outputs(4823) <= not a;
    outputs(4824) <= a xor b;
    outputs(4825) <= a and b;
    outputs(4826) <= b and not a;
    outputs(4827) <= b and not a;
    outputs(4828) <= not (a and b);
    outputs(4829) <= a or b;
    outputs(4830) <= a xor b;
    outputs(4831) <= not (a and b);
    outputs(4832) <= a xor b;
    outputs(4833) <= b;
    outputs(4834) <= not b;
    outputs(4835) <= b and not a;
    outputs(4836) <= a xor b;
    outputs(4837) <= not (a or b);
    outputs(4838) <= not b;
    outputs(4839) <= not b;
    outputs(4840) <= not (a xor b);
    outputs(4841) <= not a or b;
    outputs(4842) <= a xor b;
    outputs(4843) <= not a or b;
    outputs(4844) <= a xor b;
    outputs(4845) <= not (a xor b);
    outputs(4846) <= not b;
    outputs(4847) <= not (a or b);
    outputs(4848) <= a and b;
    outputs(4849) <= not (a and b);
    outputs(4850) <= a xor b;
    outputs(4851) <= not b or a;
    outputs(4852) <= a and not b;
    outputs(4853) <= b and not a;
    outputs(4854) <= not (a xor b);
    outputs(4855) <= a or b;
    outputs(4856) <= not b;
    outputs(4857) <= not b or a;
    outputs(4858) <= b;
    outputs(4859) <= not a;
    outputs(4860) <= not a;
    outputs(4861) <= not a;
    outputs(4862) <= not (a xor b);
    outputs(4863) <= b;
    outputs(4864) <= not (a xor b);
    outputs(4865) <= a xor b;
    outputs(4866) <= b;
    outputs(4867) <= not (a xor b);
    outputs(4868) <= not b or a;
    outputs(4869) <= not a;
    outputs(4870) <= b;
    outputs(4871) <= a xor b;
    outputs(4872) <= a;
    outputs(4873) <= not a;
    outputs(4874) <= not a;
    outputs(4875) <= b;
    outputs(4876) <= a;
    outputs(4877) <= not (a xor b);
    outputs(4878) <= not b;
    outputs(4879) <= a xor b;
    outputs(4880) <= not b;
    outputs(4881) <= not (a xor b);
    outputs(4882) <= not b or a;
    outputs(4883) <= a xor b;
    outputs(4884) <= not (a or b);
    outputs(4885) <= not b;
    outputs(4886) <= b;
    outputs(4887) <= not b;
    outputs(4888) <= a or b;
    outputs(4889) <= not (a xor b);
    outputs(4890) <= a or b;
    outputs(4891) <= b;
    outputs(4892) <= a;
    outputs(4893) <= not (a xor b);
    outputs(4894) <= a;
    outputs(4895) <= a;
    outputs(4896) <= not (a xor b);
    outputs(4897) <= b;
    outputs(4898) <= not b or a;
    outputs(4899) <= a xor b;
    outputs(4900) <= a xor b;
    outputs(4901) <= a xor b;
    outputs(4902) <= not (a xor b);
    outputs(4903) <= a and not b;
    outputs(4904) <= not b;
    outputs(4905) <= a xor b;
    outputs(4906) <= a xor b;
    outputs(4907) <= a;
    outputs(4908) <= b;
    outputs(4909) <= a xor b;
    outputs(4910) <= a and b;
    outputs(4911) <= a and not b;
    outputs(4912) <= a xor b;
    outputs(4913) <= not b;
    outputs(4914) <= not a;
    outputs(4915) <= a and not b;
    outputs(4916) <= not (a xor b);
    outputs(4917) <= not (a xor b);
    outputs(4918) <= not a;
    outputs(4919) <= a xor b;
    outputs(4920) <= not (a xor b);
    outputs(4921) <= not b;
    outputs(4922) <= a or b;
    outputs(4923) <= a xor b;
    outputs(4924) <= a xor b;
    outputs(4925) <= not a;
    outputs(4926) <= a xor b;
    outputs(4927) <= a;
    outputs(4928) <= not (a xor b);
    outputs(4929) <= a xor b;
    outputs(4930) <= not (a and b);
    outputs(4931) <= not b or a;
    outputs(4932) <= a or b;
    outputs(4933) <= a or b;
    outputs(4934) <= not a;
    outputs(4935) <= a or b;
    outputs(4936) <= not (a or b);
    outputs(4937) <= a;
    outputs(4938) <= not (a xor b);
    outputs(4939) <= not b;
    outputs(4940) <= not (a xor b);
    outputs(4941) <= not b or a;
    outputs(4942) <= not (a and b);
    outputs(4943) <= not b;
    outputs(4944) <= not b;
    outputs(4945) <= not b;
    outputs(4946) <= a;
    outputs(4947) <= not a or b;
    outputs(4948) <= not (a xor b);
    outputs(4949) <= b and not a;
    outputs(4950) <= not b;
    outputs(4951) <= a;
    outputs(4952) <= a;
    outputs(4953) <= a and b;
    outputs(4954) <= not (a xor b);
    outputs(4955) <= not a;
    outputs(4956) <= not (a or b);
    outputs(4957) <= a and b;
    outputs(4958) <= not (a xor b);
    outputs(4959) <= not b or a;
    outputs(4960) <= not a;
    outputs(4961) <= a;
    outputs(4962) <= a xor b;
    outputs(4963) <= a or b;
    outputs(4964) <= not b or a;
    outputs(4965) <= a or b;
    outputs(4966) <= a;
    outputs(4967) <= a;
    outputs(4968) <= a;
    outputs(4969) <= not (a xor b);
    outputs(4970) <= not (a or b);
    outputs(4971) <= a;
    outputs(4972) <= not b or a;
    outputs(4973) <= not (a xor b);
    outputs(4974) <= b and not a;
    outputs(4975) <= not a or b;
    outputs(4976) <= b;
    outputs(4977) <= a xor b;
    outputs(4978) <= not (a xor b);
    outputs(4979) <= not (a xor b);
    outputs(4980) <= not b;
    outputs(4981) <= a and not b;
    outputs(4982) <= not (a xor b);
    outputs(4983) <= b;
    outputs(4984) <= not (a and b);
    outputs(4985) <= a or b;
    outputs(4986) <= not a;
    outputs(4987) <= b;
    outputs(4988) <= not a;
    outputs(4989) <= b;
    outputs(4990) <= b;
    outputs(4991) <= b;
    outputs(4992) <= not (a xor b);
    outputs(4993) <= b;
    outputs(4994) <= not (a xor b);
    outputs(4995) <= not a;
    outputs(4996) <= not a;
    outputs(4997) <= not (a and b);
    outputs(4998) <= not b or a;
    outputs(4999) <= b;
    outputs(5000) <= a;
    outputs(5001) <= a xor b;
    outputs(5002) <= not (a xor b);
    outputs(5003) <= a xor b;
    outputs(5004) <= a xor b;
    outputs(5005) <= not (a xor b);
    outputs(5006) <= not b;
    outputs(5007) <= a xor b;
    outputs(5008) <= not (a xor b);
    outputs(5009) <= not a;
    outputs(5010) <= a;
    outputs(5011) <= a;
    outputs(5012) <= not (a xor b);
    outputs(5013) <= a xor b;
    outputs(5014) <= not a;
    outputs(5015) <= a and b;
    outputs(5016) <= not a;
    outputs(5017) <= not b or a;
    outputs(5018) <= not a or b;
    outputs(5019) <= b;
    outputs(5020) <= not (a xor b);
    outputs(5021) <= a;
    outputs(5022) <= not b;
    outputs(5023) <= not b;
    outputs(5024) <= a xor b;
    outputs(5025) <= not (a or b);
    outputs(5026) <= not b;
    outputs(5027) <= a and not b;
    outputs(5028) <= not b;
    outputs(5029) <= not a;
    outputs(5030) <= a xor b;
    outputs(5031) <= not a;
    outputs(5032) <= not a;
    outputs(5033) <= a xor b;
    outputs(5034) <= a xor b;
    outputs(5035) <= not (a and b);
    outputs(5036) <= a;
    outputs(5037) <= not a or b;
    outputs(5038) <= a xor b;
    outputs(5039) <= not a;
    outputs(5040) <= not (a xor b);
    outputs(5041) <= not b or a;
    outputs(5042) <= a xor b;
    outputs(5043) <= a;
    outputs(5044) <= not a;
    outputs(5045) <= not (a xor b);
    outputs(5046) <= a;
    outputs(5047) <= a xor b;
    outputs(5048) <= not a;
    outputs(5049) <= not b;
    outputs(5050) <= a;
    outputs(5051) <= not b;
    outputs(5052) <= not b or a;
    outputs(5053) <= b;
    outputs(5054) <= a xor b;
    outputs(5055) <= b;
    outputs(5056) <= not (a xor b);
    outputs(5057) <= a xor b;
    outputs(5058) <= not (a or b);
    outputs(5059) <= a;
    outputs(5060) <= a;
    outputs(5061) <= not (a xor b);
    outputs(5062) <= not b or a;
    outputs(5063) <= not a or b;
    outputs(5064) <= not (a xor b);
    outputs(5065) <= b;
    outputs(5066) <= not (a and b);
    outputs(5067) <= not a;
    outputs(5068) <= b;
    outputs(5069) <= a xor b;
    outputs(5070) <= a xor b;
    outputs(5071) <= not b;
    outputs(5072) <= a xor b;
    outputs(5073) <= a xor b;
    outputs(5074) <= not a or b;
    outputs(5075) <= not (a xor b);
    outputs(5076) <= not a;
    outputs(5077) <= not (a xor b);
    outputs(5078) <= b;
    outputs(5079) <= not (a xor b);
    outputs(5080) <= not a or b;
    outputs(5081) <= a;
    outputs(5082) <= not (a or b);
    outputs(5083) <= a xor b;
    outputs(5084) <= a and b;
    outputs(5085) <= not b or a;
    outputs(5086) <= not b or a;
    outputs(5087) <= a xor b;
    outputs(5088) <= not (a and b);
    outputs(5089) <= b;
    outputs(5090) <= not (a or b);
    outputs(5091) <= b;
    outputs(5092) <= not a or b;
    outputs(5093) <= b and not a;
    outputs(5094) <= a;
    outputs(5095) <= a;
    outputs(5096) <= not (a xor b);
    outputs(5097) <= a xor b;
    outputs(5098) <= not (a xor b);
    outputs(5099) <= not (a xor b);
    outputs(5100) <= a;
    outputs(5101) <= not (a or b);
    outputs(5102) <= not (a and b);
    outputs(5103) <= a or b;
    outputs(5104) <= a xor b;
    outputs(5105) <= a xor b;
    outputs(5106) <= a;
    outputs(5107) <= not (a or b);
    outputs(5108) <= not a;
    outputs(5109) <= a;
    outputs(5110) <= a and b;
    outputs(5111) <= a xor b;
    outputs(5112) <= not (a or b);
    outputs(5113) <= a and b;
    outputs(5114) <= not (a xor b);
    outputs(5115) <= not (a xor b);
    outputs(5116) <= not b;
    outputs(5117) <= not (a or b);
    outputs(5118) <= not (a xor b);
    outputs(5119) <= b and not a;
    outputs(5120) <= a xor b;
    outputs(5121) <= b;
    outputs(5122) <= b;
    outputs(5123) <= b;
    outputs(5124) <= not a;
    outputs(5125) <= not a;
    outputs(5126) <= not a;
    outputs(5127) <= not (a or b);
    outputs(5128) <= not (a or b);
    outputs(5129) <= not (a and b);
    outputs(5130) <= a xor b;
    outputs(5131) <= not b or a;
    outputs(5132) <= not a or b;
    outputs(5133) <= a xor b;
    outputs(5134) <= not (a xor b);
    outputs(5135) <= a and b;
    outputs(5136) <= not (a xor b);
    outputs(5137) <= a xor b;
    outputs(5138) <= not a or b;
    outputs(5139) <= not a;
    outputs(5140) <= b;
    outputs(5141) <= a and b;
    outputs(5142) <= a;
    outputs(5143) <= not b;
    outputs(5144) <= not a or b;
    outputs(5145) <= not (a xor b);
    outputs(5146) <= a and not b;
    outputs(5147) <= not b;
    outputs(5148) <= a and b;
    outputs(5149) <= not b;
    outputs(5150) <= a xor b;
    outputs(5151) <= not (a xor b);
    outputs(5152) <= not b;
    outputs(5153) <= not (a xor b);
    outputs(5154) <= not (a and b);
    outputs(5155) <= a xor b;
    outputs(5156) <= not (a xor b);
    outputs(5157) <= a;
    outputs(5158) <= b;
    outputs(5159) <= not b or a;
    outputs(5160) <= a;
    outputs(5161) <= a xor b;
    outputs(5162) <= a or b;
    outputs(5163) <= not a;
    outputs(5164) <= not (a xor b);
    outputs(5165) <= b;
    outputs(5166) <= not (a xor b);
    outputs(5167) <= a and b;
    outputs(5168) <= not a or b;
    outputs(5169) <= not (a xor b);
    outputs(5170) <= not (a xor b);
    outputs(5171) <= b and not a;
    outputs(5172) <= a xor b;
    outputs(5173) <= a xor b;
    outputs(5174) <= a;
    outputs(5175) <= b;
    outputs(5176) <= a xor b;
    outputs(5177) <= not (a xor b);
    outputs(5178) <= a xor b;
    outputs(5179) <= not (a xor b);
    outputs(5180) <= b;
    outputs(5181) <= a xor b;
    outputs(5182) <= a and not b;
    outputs(5183) <= a and not b;
    outputs(5184) <= b;
    outputs(5185) <= not b;
    outputs(5186) <= not b;
    outputs(5187) <= b;
    outputs(5188) <= a xor b;
    outputs(5189) <= not b;
    outputs(5190) <= not b;
    outputs(5191) <= a;
    outputs(5192) <= a;
    outputs(5193) <= b;
    outputs(5194) <= a xor b;
    outputs(5195) <= not (a or b);
    outputs(5196) <= not b;
    outputs(5197) <= a;
    outputs(5198) <= not b;
    outputs(5199) <= a and not b;
    outputs(5200) <= not (a xor b);
    outputs(5201) <= a xor b;
    outputs(5202) <= not (a xor b);
    outputs(5203) <= not (a xor b);
    outputs(5204) <= a;
    outputs(5205) <= a xor b;
    outputs(5206) <= a;
    outputs(5207) <= a xor b;
    outputs(5208) <= not b;
    outputs(5209) <= not (a or b);
    outputs(5210) <= not (a xor b);
    outputs(5211) <= a;
    outputs(5212) <= not (a xor b);
    outputs(5213) <= not a;
    outputs(5214) <= not a;
    outputs(5215) <= b;
    outputs(5216) <= a;
    outputs(5217) <= not b;
    outputs(5218) <= a;
    outputs(5219) <= a and not b;
    outputs(5220) <= not b;
    outputs(5221) <= a xor b;
    outputs(5222) <= not b;
    outputs(5223) <= b;
    outputs(5224) <= a xor b;
    outputs(5225) <= b and not a;
    outputs(5226) <= b and not a;
    outputs(5227) <= a;
    outputs(5228) <= a xor b;
    outputs(5229) <= not a;
    outputs(5230) <= b;
    outputs(5231) <= a and not b;
    outputs(5232) <= not (a xor b);
    outputs(5233) <= not b;
    outputs(5234) <= not (a or b);
    outputs(5235) <= b;
    outputs(5236) <= a xor b;
    outputs(5237) <= b;
    outputs(5238) <= a or b;
    outputs(5239) <= not (a xor b);
    outputs(5240) <= a xor b;
    outputs(5241) <= b;
    outputs(5242) <= not b;
    outputs(5243) <= b;
    outputs(5244) <= b;
    outputs(5245) <= not (a xor b);
    outputs(5246) <= not (a or b);
    outputs(5247) <= a xor b;
    outputs(5248) <= b;
    outputs(5249) <= not (a or b);
    outputs(5250) <= not (a xor b);
    outputs(5251) <= b and not a;
    outputs(5252) <= not (a or b);
    outputs(5253) <= b and not a;
    outputs(5254) <= a xor b;
    outputs(5255) <= a;
    outputs(5256) <= b;
    outputs(5257) <= not (a or b);
    outputs(5258) <= not (a xor b);
    outputs(5259) <= not a;
    outputs(5260) <= not (a xor b);
    outputs(5261) <= not a;
    outputs(5262) <= not (a xor b);
    outputs(5263) <= not a;
    outputs(5264) <= not a;
    outputs(5265) <= not (a xor b);
    outputs(5266) <= not (a xor b);
    outputs(5267) <= a xor b;
    outputs(5268) <= a and b;
    outputs(5269) <= a;
    outputs(5270) <= a;
    outputs(5271) <= a xor b;
    outputs(5272) <= not (a xor b);
    outputs(5273) <= not (a xor b);
    outputs(5274) <= not (a xor b);
    outputs(5275) <= b;
    outputs(5276) <= b;
    outputs(5277) <= a;
    outputs(5278) <= a;
    outputs(5279) <= not (a xor b);
    outputs(5280) <= a xor b;
    outputs(5281) <= not (a or b);
    outputs(5282) <= not b;
    outputs(5283) <= not a or b;
    outputs(5284) <= not b;
    outputs(5285) <= a xor b;
    outputs(5286) <= b and not a;
    outputs(5287) <= not (a or b);
    outputs(5288) <= not (a or b);
    outputs(5289) <= a;
    outputs(5290) <= not (a xor b);
    outputs(5291) <= not b;
    outputs(5292) <= not b;
    outputs(5293) <= not a;
    outputs(5294) <= a xor b;
    outputs(5295) <= a xor b;
    outputs(5296) <= a or b;
    outputs(5297) <= b;
    outputs(5298) <= a;
    outputs(5299) <= not a or b;
    outputs(5300) <= not (a xor b);
    outputs(5301) <= not (a xor b);
    outputs(5302) <= a;
    outputs(5303) <= b;
    outputs(5304) <= a xor b;
    outputs(5305) <= not b or a;
    outputs(5306) <= not (a xor b);
    outputs(5307) <= not b;
    outputs(5308) <= not b;
    outputs(5309) <= not (a or b);
    outputs(5310) <= not a;
    outputs(5311) <= b;
    outputs(5312) <= a xor b;
    outputs(5313) <= a;
    outputs(5314) <= not a;
    outputs(5315) <= a;
    outputs(5316) <= not (a xor b);
    outputs(5317) <= b;
    outputs(5318) <= not b or a;
    outputs(5319) <= not (a xor b);
    outputs(5320) <= not a;
    outputs(5321) <= not a;
    outputs(5322) <= not b;
    outputs(5323) <= a xor b;
    outputs(5324) <= not (a or b);
    outputs(5325) <= not a;
    outputs(5326) <= not a;
    outputs(5327) <= not (a xor b);
    outputs(5328) <= not b;
    outputs(5329) <= b;
    outputs(5330) <= not (a xor b);
    outputs(5331) <= a and b;
    outputs(5332) <= not (a xor b);
    outputs(5333) <= not (a xor b);
    outputs(5334) <= not b or a;
    outputs(5335) <= a xor b;
    outputs(5336) <= a xor b;
    outputs(5337) <= a or b;
    outputs(5338) <= b and not a;
    outputs(5339) <= not (a or b);
    outputs(5340) <= not a;
    outputs(5341) <= not (a xor b);
    outputs(5342) <= not b;
    outputs(5343) <= b;
    outputs(5344) <= not (a xor b);
    outputs(5345) <= a and b;
    outputs(5346) <= not (a or b);
    outputs(5347) <= a;
    outputs(5348) <= not b;
    outputs(5349) <= a and not b;
    outputs(5350) <= b and not a;
    outputs(5351) <= b;
    outputs(5352) <= b;
    outputs(5353) <= not a;
    outputs(5354) <= a xor b;
    outputs(5355) <= a xor b;
    outputs(5356) <= a xor b;
    outputs(5357) <= a;
    outputs(5358) <= not (a xor b);
    outputs(5359) <= a or b;
    outputs(5360) <= not (a or b);
    outputs(5361) <= a;
    outputs(5362) <= not a;
    outputs(5363) <= not a or b;
    outputs(5364) <= b;
    outputs(5365) <= not a;
    outputs(5366) <= b;
    outputs(5367) <= b and not a;
    outputs(5368) <= b;
    outputs(5369) <= a and not b;
    outputs(5370) <= a and not b;
    outputs(5371) <= b and not a;
    outputs(5372) <= not b;
    outputs(5373) <= not a or b;
    outputs(5374) <= b;
    outputs(5375) <= a and b;
    outputs(5376) <= a or b;
    outputs(5377) <= b;
    outputs(5378) <= not b;
    outputs(5379) <= not b or a;
    outputs(5380) <= a xor b;
    outputs(5381) <= not a;
    outputs(5382) <= not (a xor b);
    outputs(5383) <= b and not a;
    outputs(5384) <= b;
    outputs(5385) <= a and not b;
    outputs(5386) <= a and b;
    outputs(5387) <= not (a or b);
    outputs(5388) <= not (a xor b);
    outputs(5389) <= not (a xor b);
    outputs(5390) <= not b;
    outputs(5391) <= not b;
    outputs(5392) <= not a;
    outputs(5393) <= not b;
    outputs(5394) <= a and b;
    outputs(5395) <= not (a xor b);
    outputs(5396) <= a xor b;
    outputs(5397) <= a;
    outputs(5398) <= b and not a;
    outputs(5399) <= b and not a;
    outputs(5400) <= b and not a;
    outputs(5401) <= not b or a;
    outputs(5402) <= not (a xor b);
    outputs(5403) <= not (a xor b);
    outputs(5404) <= not (a or b);
    outputs(5405) <= a;
    outputs(5406) <= a xor b;
    outputs(5407) <= a xor b;
    outputs(5408) <= not b;
    outputs(5409) <= b;
    outputs(5410) <= b;
    outputs(5411) <= a xor b;
    outputs(5412) <= not a;
    outputs(5413) <= a xor b;
    outputs(5414) <= not (a xor b);
    outputs(5415) <= not (a or b);
    outputs(5416) <= a;
    outputs(5417) <= a xor b;
    outputs(5418) <= not b;
    outputs(5419) <= not (a or b);
    outputs(5420) <= not a;
    outputs(5421) <= b;
    outputs(5422) <= b;
    outputs(5423) <= not (a xor b);
    outputs(5424) <= a xor b;
    outputs(5425) <= a xor b;
    outputs(5426) <= a xor b;
    outputs(5427) <= b;
    outputs(5428) <= a;
    outputs(5429) <= a xor b;
    outputs(5430) <= a or b;
    outputs(5431) <= a;
    outputs(5432) <= a xor b;
    outputs(5433) <= b and not a;
    outputs(5434) <= b;
    outputs(5435) <= not a;
    outputs(5436) <= a and b;
    outputs(5437) <= a and b;
    outputs(5438) <= b;
    outputs(5439) <= not (a or b);
    outputs(5440) <= a;
    outputs(5441) <= a and not b;
    outputs(5442) <= not b;
    outputs(5443) <= a;
    outputs(5444) <= a xor b;
    outputs(5445) <= not (a xor b);
    outputs(5446) <= not (a or b);
    outputs(5447) <= a xor b;
    outputs(5448) <= not b;
    outputs(5449) <= b;
    outputs(5450) <= not a;
    outputs(5451) <= not a;
    outputs(5452) <= a xor b;
    outputs(5453) <= a xor b;
    outputs(5454) <= not a;
    outputs(5455) <= b and not a;
    outputs(5456) <= a and b;
    outputs(5457) <= not b;
    outputs(5458) <= not (a and b);
    outputs(5459) <= a;
    outputs(5460) <= not b;
    outputs(5461) <= not (a xor b);
    outputs(5462) <= not (a xor b);
    outputs(5463) <= b and not a;
    outputs(5464) <= not (a xor b);
    outputs(5465) <= not b;
    outputs(5466) <= not (a xor b);
    outputs(5467) <= b;
    outputs(5468) <= not (a xor b);
    outputs(5469) <= a xor b;
    outputs(5470) <= a and b;
    outputs(5471) <= b;
    outputs(5472) <= not b;
    outputs(5473) <= b;
    outputs(5474) <= b;
    outputs(5475) <= not (a xor b);
    outputs(5476) <= not (a or b);
    outputs(5477) <= not (a or b);
    outputs(5478) <= not b;
    outputs(5479) <= a xor b;
    outputs(5480) <= a xor b;
    outputs(5481) <= not (a xor b);
    outputs(5482) <= a and b;
    outputs(5483) <= a and not b;
    outputs(5484) <= a or b;
    outputs(5485) <= a and b;
    outputs(5486) <= a xor b;
    outputs(5487) <= not b;
    outputs(5488) <= b;
    outputs(5489) <= a and not b;
    outputs(5490) <= b;
    outputs(5491) <= b;
    outputs(5492) <= b;
    outputs(5493) <= not (a xor b);
    outputs(5494) <= a;
    outputs(5495) <= not (a xor b);
    outputs(5496) <= not (a xor b);
    outputs(5497) <= not a;
    outputs(5498) <= a xor b;
    outputs(5499) <= not a;
    outputs(5500) <= a xor b;
    outputs(5501) <= a and b;
    outputs(5502) <= not b;
    outputs(5503) <= not b;
    outputs(5504) <= a;
    outputs(5505) <= a;
    outputs(5506) <= not (a xor b);
    outputs(5507) <= a xor b;
    outputs(5508) <= not a;
    outputs(5509) <= a and b;
    outputs(5510) <= not a;
    outputs(5511) <= not (a xor b);
    outputs(5512) <= b;
    outputs(5513) <= a and b;
    outputs(5514) <= a and not b;
    outputs(5515) <= not b;
    outputs(5516) <= not b;
    outputs(5517) <= a and not b;
    outputs(5518) <= not (a xor b);
    outputs(5519) <= a xor b;
    outputs(5520) <= a xor b;
    outputs(5521) <= a xor b;
    outputs(5522) <= a;
    outputs(5523) <= not b;
    outputs(5524) <= not b;
    outputs(5525) <= not a;
    outputs(5526) <= a xor b;
    outputs(5527) <= not b;
    outputs(5528) <= b;
    outputs(5529) <= b and not a;
    outputs(5530) <= a and not b;
    outputs(5531) <= a xor b;
    outputs(5532) <= b;
    outputs(5533) <= not (a xor b);
    outputs(5534) <= a xor b;
    outputs(5535) <= a xor b;
    outputs(5536) <= not (a xor b);
    outputs(5537) <= not (a xor b);
    outputs(5538) <= a;
    outputs(5539) <= b;
    outputs(5540) <= a and b;
    outputs(5541) <= not (a xor b);
    outputs(5542) <= not a;
    outputs(5543) <= a and not b;
    outputs(5544) <= a;
    outputs(5545) <= not b;
    outputs(5546) <= a;
    outputs(5547) <= not a;
    outputs(5548) <= not b or a;
    outputs(5549) <= not a;
    outputs(5550) <= a;
    outputs(5551) <= not (a xor b);
    outputs(5552) <= a xor b;
    outputs(5553) <= a;
    outputs(5554) <= a and b;
    outputs(5555) <= b;
    outputs(5556) <= a xor b;
    outputs(5557) <= not a;
    outputs(5558) <= not (a xor b);
    outputs(5559) <= b;
    outputs(5560) <= a xor b;
    outputs(5561) <= a xor b;
    outputs(5562) <= not (a xor b);
    outputs(5563) <= a xor b;
    outputs(5564) <= b;
    outputs(5565) <= a or b;
    outputs(5566) <= not (a xor b);
    outputs(5567) <= b;
    outputs(5568) <= a;
    outputs(5569) <= not (a or b);
    outputs(5570) <= not a;
    outputs(5571) <= not b or a;
    outputs(5572) <= a xor b;
    outputs(5573) <= not (a xor b);
    outputs(5574) <= not a;
    outputs(5575) <= a xor b;
    outputs(5576) <= a and not b;
    outputs(5577) <= not a;
    outputs(5578) <= a xor b;
    outputs(5579) <= not (a xor b);
    outputs(5580) <= not b or a;
    outputs(5581) <= not (a xor b);
    outputs(5582) <= not b;
    outputs(5583) <= not (a and b);
    outputs(5584) <= a and not b;
    outputs(5585) <= a;
    outputs(5586) <= a xor b;
    outputs(5587) <= b and not a;
    outputs(5588) <= not b;
    outputs(5589) <= a xor b;
    outputs(5590) <= not b;
    outputs(5591) <= not (a or b);
    outputs(5592) <= b;
    outputs(5593) <= b;
    outputs(5594) <= not (a xor b);
    outputs(5595) <= a xor b;
    outputs(5596) <= a and b;
    outputs(5597) <= b;
    outputs(5598) <= a xor b;
    outputs(5599) <= a and b;
    outputs(5600) <= not (a or b);
    outputs(5601) <= not (a and b);
    outputs(5602) <= a or b;
    outputs(5603) <= a;
    outputs(5604) <= a and b;
    outputs(5605) <= b;
    outputs(5606) <= b and not a;
    outputs(5607) <= b and not a;
    outputs(5608) <= a and b;
    outputs(5609) <= not b;
    outputs(5610) <= not b or a;
    outputs(5611) <= a xor b;
    outputs(5612) <= not b;
    outputs(5613) <= not b;
    outputs(5614) <= b;
    outputs(5615) <= not (a xor b);
    outputs(5616) <= b;
    outputs(5617) <= not (a xor b);
    outputs(5618) <= not b;
    outputs(5619) <= not b;
    outputs(5620) <= a and not b;
    outputs(5621) <= not (a xor b);
    outputs(5622) <= not a;
    outputs(5623) <= a xor b;
    outputs(5624) <= not b or a;
    outputs(5625) <= b;
    outputs(5626) <= not b;
    outputs(5627) <= a and not b;
    outputs(5628) <= not (a xor b);
    outputs(5629) <= a and b;
    outputs(5630) <= a or b;
    outputs(5631) <= not a;
    outputs(5632) <= not (a xor b);
    outputs(5633) <= not b;
    outputs(5634) <= a;
    outputs(5635) <= not a;
    outputs(5636) <= not b;
    outputs(5637) <= not b;
    outputs(5638) <= not (a xor b);
    outputs(5639) <= not (a or b);
    outputs(5640) <= not a;
    outputs(5641) <= not (a or b);
    outputs(5642) <= b;
    outputs(5643) <= not a;
    outputs(5644) <= not a;
    outputs(5645) <= not b;
    outputs(5646) <= b;
    outputs(5647) <= not (a xor b);
    outputs(5648) <= b;
    outputs(5649) <= a and b;
    outputs(5650) <= not a;
    outputs(5651) <= a or b;
    outputs(5652) <= a and b;
    outputs(5653) <= not (a and b);
    outputs(5654) <= not a;
    outputs(5655) <= not a;
    outputs(5656) <= not (a or b);
    outputs(5657) <= not (a xor b);
    outputs(5658) <= not (a xor b);
    outputs(5659) <= b;
    outputs(5660) <= a xor b;
    outputs(5661) <= b;
    outputs(5662) <= not (a xor b);
    outputs(5663) <= not a or b;
    outputs(5664) <= not (a xor b);
    outputs(5665) <= not (a xor b);
    outputs(5666) <= a;
    outputs(5667) <= not a;
    outputs(5668) <= a or b;
    outputs(5669) <= a and b;
    outputs(5670) <= a xor b;
    outputs(5671) <= not (a xor b);
    outputs(5672) <= a;
    outputs(5673) <= a;
    outputs(5674) <= not b or a;
    outputs(5675) <= a xor b;
    outputs(5676) <= not b;
    outputs(5677) <= a xor b;
    outputs(5678) <= not (a xor b);
    outputs(5679) <= a and not b;
    outputs(5680) <= not a;
    outputs(5681) <= a xor b;
    outputs(5682) <= a and not b;
    outputs(5683) <= not a or b;
    outputs(5684) <= a;
    outputs(5685) <= not a;
    outputs(5686) <= not (a xor b);
    outputs(5687) <= not a or b;
    outputs(5688) <= a;
    outputs(5689) <= not (a or b);
    outputs(5690) <= not (a xor b);
    outputs(5691) <= not b;
    outputs(5692) <= a;
    outputs(5693) <= not b;
    outputs(5694) <= b;
    outputs(5695) <= not b;
    outputs(5696) <= not b;
    outputs(5697) <= a xor b;
    outputs(5698) <= not (a xor b);
    outputs(5699) <= a xor b;
    outputs(5700) <= a;
    outputs(5701) <= not a;
    outputs(5702) <= a;
    outputs(5703) <= a;
    outputs(5704) <= not (a xor b);
    outputs(5705) <= not b;
    outputs(5706) <= a xor b;
    outputs(5707) <= b and not a;
    outputs(5708) <= not (a xor b);
    outputs(5709) <= not a;
    outputs(5710) <= not a;
    outputs(5711) <= not (a xor b);
    outputs(5712) <= b;
    outputs(5713) <= not (a or b);
    outputs(5714) <= a;
    outputs(5715) <= not b;
    outputs(5716) <= not a;
    outputs(5717) <= not (a or b);
    outputs(5718) <= not a;
    outputs(5719) <= not a;
    outputs(5720) <= not b;
    outputs(5721) <= a xor b;
    outputs(5722) <= not b;
    outputs(5723) <= not a;
    outputs(5724) <= not b;
    outputs(5725) <= not a;
    outputs(5726) <= not (a xor b);
    outputs(5727) <= b and not a;
    outputs(5728) <= not b;
    outputs(5729) <= not (a and b);
    outputs(5730) <= b and not a;
    outputs(5731) <= not (a or b);
    outputs(5732) <= b;
    outputs(5733) <= not (a xor b);
    outputs(5734) <= a xor b;
    outputs(5735) <= a and b;
    outputs(5736) <= a;
    outputs(5737) <= b and not a;
    outputs(5738) <= not b;
    outputs(5739) <= b and not a;
    outputs(5740) <= a xor b;
    outputs(5741) <= not b;
    outputs(5742) <= a xor b;
    outputs(5743) <= a;
    outputs(5744) <= b;
    outputs(5745) <= not (a xor b);
    outputs(5746) <= not b;
    outputs(5747) <= a or b;
    outputs(5748) <= a and not b;
    outputs(5749) <= not a;
    outputs(5750) <= b;
    outputs(5751) <= b;
    outputs(5752) <= a and not b;
    outputs(5753) <= not b or a;
    outputs(5754) <= not (a xor b);
    outputs(5755) <= a xor b;
    outputs(5756) <= b;
    outputs(5757) <= not a;
    outputs(5758) <= b;
    outputs(5759) <= not b;
    outputs(5760) <= a;
    outputs(5761) <= a xor b;
    outputs(5762) <= b;
    outputs(5763) <= not (a xor b);
    outputs(5764) <= a;
    outputs(5765) <= b;
    outputs(5766) <= not b;
    outputs(5767) <= not b or a;
    outputs(5768) <= a and b;
    outputs(5769) <= a xor b;
    outputs(5770) <= b and not a;
    outputs(5771) <= a or b;
    outputs(5772) <= a;
    outputs(5773) <= not (a xor b);
    outputs(5774) <= a xor b;
    outputs(5775) <= not (a xor b);
    outputs(5776) <= not b;
    outputs(5777) <= b;
    outputs(5778) <= b;
    outputs(5779) <= a and b;
    outputs(5780) <= b;
    outputs(5781) <= not (a xor b);
    outputs(5782) <= not a or b;
    outputs(5783) <= not b;
    outputs(5784) <= not b;
    outputs(5785) <= b;
    outputs(5786) <= not a;
    outputs(5787) <= not (a xor b);
    outputs(5788) <= not b;
    outputs(5789) <= not (a or b);
    outputs(5790) <= a;
    outputs(5791) <= a xor b;
    outputs(5792) <= not (a xor b);
    outputs(5793) <= not a;
    outputs(5794) <= not b;
    outputs(5795) <= not b;
    outputs(5796) <= not (a or b);
    outputs(5797) <= not a or b;
    outputs(5798) <= a xor b;
    outputs(5799) <= a and not b;
    outputs(5800) <= a;
    outputs(5801) <= a xor b;
    outputs(5802) <= not (a or b);
    outputs(5803) <= not a;
    outputs(5804) <= not b;
    outputs(5805) <= a xor b;
    outputs(5806) <= a xor b;
    outputs(5807) <= a and not b;
    outputs(5808) <= a;
    outputs(5809) <= not (a xor b);
    outputs(5810) <= not a;
    outputs(5811) <= b;
    outputs(5812) <= b;
    outputs(5813) <= not (a xor b);
    outputs(5814) <= not (a xor b);
    outputs(5815) <= a or b;
    outputs(5816) <= not a;
    outputs(5817) <= not (a xor b);
    outputs(5818) <= a xor b;
    outputs(5819) <= a or b;
    outputs(5820) <= not b;
    outputs(5821) <= a;
    outputs(5822) <= a and not b;
    outputs(5823) <= not b;
    outputs(5824) <= a xor b;
    outputs(5825) <= a;
    outputs(5826) <= b and not a;
    outputs(5827) <= a and b;
    outputs(5828) <= a and not b;
    outputs(5829) <= b;
    outputs(5830) <= a or b;
    outputs(5831) <= not a;
    outputs(5832) <= b;
    outputs(5833) <= b and not a;
    outputs(5834) <= not (a xor b);
    outputs(5835) <= b;
    outputs(5836) <= not (a or b);
    outputs(5837) <= b;
    outputs(5838) <= not a;
    outputs(5839) <= a;
    outputs(5840) <= not a;
    outputs(5841) <= not (a xor b);
    outputs(5842) <= a xor b;
    outputs(5843) <= not b;
    outputs(5844) <= a xor b;
    outputs(5845) <= a and b;
    outputs(5846) <= not (a or b);
    outputs(5847) <= a and not b;
    outputs(5848) <= a xor b;
    outputs(5849) <= b;
    outputs(5850) <= a;
    outputs(5851) <= a and not b;
    outputs(5852) <= a;
    outputs(5853) <= a;
    outputs(5854) <= not b;
    outputs(5855) <= a xor b;
    outputs(5856) <= not a;
    outputs(5857) <= not (a xor b);
    outputs(5858) <= a;
    outputs(5859) <= a and not b;
    outputs(5860) <= a xor b;
    outputs(5861) <= b;
    outputs(5862) <= not a;
    outputs(5863) <= not (a and b);
    outputs(5864) <= a;
    outputs(5865) <= not (a or b);
    outputs(5866) <= a and not b;
    outputs(5867) <= not a;
    outputs(5868) <= a xor b;
    outputs(5869) <= a xor b;
    outputs(5870) <= not b;
    outputs(5871) <= 1'b0;
    outputs(5872) <= b;
    outputs(5873) <= not (a xor b);
    outputs(5874) <= not (a xor b);
    outputs(5875) <= a and not b;
    outputs(5876) <= a xor b;
    outputs(5877) <= not b or a;
    outputs(5878) <= a and not b;
    outputs(5879) <= not b;
    outputs(5880) <= b;
    outputs(5881) <= not (a or b);
    outputs(5882) <= not (a xor b);
    outputs(5883) <= a xor b;
    outputs(5884) <= not a;
    outputs(5885) <= a and not b;
    outputs(5886) <= a;
    outputs(5887) <= a xor b;
    outputs(5888) <= not a;
    outputs(5889) <= a;
    outputs(5890) <= not (a or b);
    outputs(5891) <= not b;
    outputs(5892) <= not a;
    outputs(5893) <= a xor b;
    outputs(5894) <= not a;
    outputs(5895) <= a xor b;
    outputs(5896) <= not (a xor b);
    outputs(5897) <= a;
    outputs(5898) <= a;
    outputs(5899) <= a and b;
    outputs(5900) <= not b;
    outputs(5901) <= not (a xor b);
    outputs(5902) <= not (a xor b);
    outputs(5903) <= not a;
    outputs(5904) <= a;
    outputs(5905) <= not (a or b);
    outputs(5906) <= not (a xor b);
    outputs(5907) <= a;
    outputs(5908) <= b;
    outputs(5909) <= a xor b;
    outputs(5910) <= not b;
    outputs(5911) <= a xor b;
    outputs(5912) <= a xor b;
    outputs(5913) <= not (a or b);
    outputs(5914) <= not (a xor b);
    outputs(5915) <= not (a or b);
    outputs(5916) <= b;
    outputs(5917) <= b and not a;
    outputs(5918) <= a xor b;
    outputs(5919) <= not (a and b);
    outputs(5920) <= b;
    outputs(5921) <= b;
    outputs(5922) <= a and b;
    outputs(5923) <= not a;
    outputs(5924) <= a and not b;
    outputs(5925) <= a xor b;
    outputs(5926) <= b;
    outputs(5927) <= not a or b;
    outputs(5928) <= not (a xor b);
    outputs(5929) <= a;
    outputs(5930) <= not a;
    outputs(5931) <= not (a xor b);
    outputs(5932) <= not (a or b);
    outputs(5933) <= not a;
    outputs(5934) <= not a;
    outputs(5935) <= a xor b;
    outputs(5936) <= b;
    outputs(5937) <= not a;
    outputs(5938) <= b and not a;
    outputs(5939) <= a and b;
    outputs(5940) <= not (a xor b);
    outputs(5941) <= a and b;
    outputs(5942) <= b;
    outputs(5943) <= not a;
    outputs(5944) <= a and b;
    outputs(5945) <= a xor b;
    outputs(5946) <= not (a or b);
    outputs(5947) <= not a;
    outputs(5948) <= not a;
    outputs(5949) <= not b;
    outputs(5950) <= a;
    outputs(5951) <= b and not a;
    outputs(5952) <= not a;
    outputs(5953) <= a and b;
    outputs(5954) <= not (a xor b);
    outputs(5955) <= a and not b;
    outputs(5956) <= not (a or b);
    outputs(5957) <= not b;
    outputs(5958) <= not (a xor b);
    outputs(5959) <= not (a xor b);
    outputs(5960) <= not (a xor b);
    outputs(5961) <= not a;
    outputs(5962) <= not a;
    outputs(5963) <= a;
    outputs(5964) <= b;
    outputs(5965) <= a xor b;
    outputs(5966) <= a xor b;
    outputs(5967) <= not b;
    outputs(5968) <= not (a and b);
    outputs(5969) <= not b or a;
    outputs(5970) <= a;
    outputs(5971) <= not b;
    outputs(5972) <= b;
    outputs(5973) <= not b;
    outputs(5974) <= not (a xor b);
    outputs(5975) <= a xor b;
    outputs(5976) <= not a;
    outputs(5977) <= not a;
    outputs(5978) <= not b;
    outputs(5979) <= not b or a;
    outputs(5980) <= not a;
    outputs(5981) <= a xor b;
    outputs(5982) <= a;
    outputs(5983) <= a and not b;
    outputs(5984) <= a;
    outputs(5985) <= a or b;
    outputs(5986) <= not b;
    outputs(5987) <= a xor b;
    outputs(5988) <= a and b;
    outputs(5989) <= not (a xor b);
    outputs(5990) <= not b;
    outputs(5991) <= a xor b;
    outputs(5992) <= a and not b;
    outputs(5993) <= a xor b;
    outputs(5994) <= not b;
    outputs(5995) <= not b;
    outputs(5996) <= a and not b;
    outputs(5997) <= a xor b;
    outputs(5998) <= a;
    outputs(5999) <= not a;
    outputs(6000) <= not (a xor b);
    outputs(6001) <= b;
    outputs(6002) <= a;
    outputs(6003) <= b;
    outputs(6004) <= a and b;
    outputs(6005) <= a xor b;
    outputs(6006) <= b;
    outputs(6007) <= b and not a;
    outputs(6008) <= b;
    outputs(6009) <= not (a xor b);
    outputs(6010) <= not b;
    outputs(6011) <= a;
    outputs(6012) <= a xor b;
    outputs(6013) <= a xor b;
    outputs(6014) <= not b;
    outputs(6015) <= not (a xor b);
    outputs(6016) <= a and b;
    outputs(6017) <= not a;
    outputs(6018) <= not (a xor b);
    outputs(6019) <= b and not a;
    outputs(6020) <= a xor b;
    outputs(6021) <= not b;
    outputs(6022) <= a;
    outputs(6023) <= a and b;
    outputs(6024) <= a;
    outputs(6025) <= a;
    outputs(6026) <= not b;
    outputs(6027) <= not b or a;
    outputs(6028) <= not a or b;
    outputs(6029) <= not a;
    outputs(6030) <= not a;
    outputs(6031) <= a or b;
    outputs(6032) <= not b;
    outputs(6033) <= not b or a;
    outputs(6034) <= not a;
    outputs(6035) <= not (a or b);
    outputs(6036) <= not b or a;
    outputs(6037) <= not b;
    outputs(6038) <= a xor b;
    outputs(6039) <= a xor b;
    outputs(6040) <= a;
    outputs(6041) <= a and b;
    outputs(6042) <= not b;
    outputs(6043) <= not (a xor b);
    outputs(6044) <= not (a xor b);
    outputs(6045) <= not b;
    outputs(6046) <= not (a xor b);
    outputs(6047) <= a and b;
    outputs(6048) <= not b;
    outputs(6049) <= b;
    outputs(6050) <= a xor b;
    outputs(6051) <= a xor b;
    outputs(6052) <= not a;
    outputs(6053) <= b;
    outputs(6054) <= not b;
    outputs(6055) <= a or b;
    outputs(6056) <= not (a xor b);
    outputs(6057) <= b and not a;
    outputs(6058) <= a and not b;
    outputs(6059) <= b;
    outputs(6060) <= not b;
    outputs(6061) <= a;
    outputs(6062) <= not (a xor b);
    outputs(6063) <= b and not a;
    outputs(6064) <= b;
    outputs(6065) <= a xor b;
    outputs(6066) <= a and b;
    outputs(6067) <= not a;
    outputs(6068) <= not (a xor b);
    outputs(6069) <= a and not b;
    outputs(6070) <= a xor b;
    outputs(6071) <= not a;
    outputs(6072) <= not (a xor b);
    outputs(6073) <= a;
    outputs(6074) <= not (a xor b);
    outputs(6075) <= not b or a;
    outputs(6076) <= not b;
    outputs(6077) <= b;
    outputs(6078) <= a and b;
    outputs(6079) <= a and not b;
    outputs(6080) <= a xor b;
    outputs(6081) <= a;
    outputs(6082) <= not (a xor b);
    outputs(6083) <= a and b;
    outputs(6084) <= a;
    outputs(6085) <= a xor b;
    outputs(6086) <= not a;
    outputs(6087) <= not b;
    outputs(6088) <= b and not a;
    outputs(6089) <= a xor b;
    outputs(6090) <= not (a or b);
    outputs(6091) <= not a or b;
    outputs(6092) <= not (a xor b);
    outputs(6093) <= b;
    outputs(6094) <= b;
    outputs(6095) <= a and b;
    outputs(6096) <= not a or b;
    outputs(6097) <= not (a or b);
    outputs(6098) <= a or b;
    outputs(6099) <= not (a xor b);
    outputs(6100) <= a xor b;
    outputs(6101) <= a;
    outputs(6102) <= a xor b;
    outputs(6103) <= not (a xor b);
    outputs(6104) <= not b or a;
    outputs(6105) <= b;
    outputs(6106) <= not (a xor b);
    outputs(6107) <= not (a xor b);
    outputs(6108) <= b;
    outputs(6109) <= a;
    outputs(6110) <= not (a xor b);
    outputs(6111) <= a xor b;
    outputs(6112) <= not a or b;
    outputs(6113) <= b;
    outputs(6114) <= a xor b;
    outputs(6115) <= b;
    outputs(6116) <= b and not a;
    outputs(6117) <= a and not b;
    outputs(6118) <= not (a xor b);
    outputs(6119) <= b and not a;
    outputs(6120) <= not b;
    outputs(6121) <= a xor b;
    outputs(6122) <= a xor b;
    outputs(6123) <= not a or b;
    outputs(6124) <= a xor b;
    outputs(6125) <= a xor b;
    outputs(6126) <= not (a xor b);
    outputs(6127) <= not a or b;
    outputs(6128) <= not (a xor b);
    outputs(6129) <= a xor b;
    outputs(6130) <= not b;
    outputs(6131) <= not (a or b);
    outputs(6132) <= a and b;
    outputs(6133) <= b;
    outputs(6134) <= not (a xor b);
    outputs(6135) <= not a;
    outputs(6136) <= b;
    outputs(6137) <= not (a or b);
    outputs(6138) <= a and not b;
    outputs(6139) <= b;
    outputs(6140) <= a xor b;
    outputs(6141) <= a;
    outputs(6142) <= not (a xor b);
    outputs(6143) <= not a;
    outputs(6144) <= b;
    outputs(6145) <= b;
    outputs(6146) <= a xor b;
    outputs(6147) <= not a;
    outputs(6148) <= not (a or b);
    outputs(6149) <= a;
    outputs(6150) <= a;
    outputs(6151) <= a xor b;
    outputs(6152) <= b;
    outputs(6153) <= a and b;
    outputs(6154) <= a and b;
    outputs(6155) <= not (a or b);
    outputs(6156) <= a xor b;
    outputs(6157) <= b and not a;
    outputs(6158) <= not (a and b);
    outputs(6159) <= a xor b;
    outputs(6160) <= not a;
    outputs(6161) <= b;
    outputs(6162) <= not a;
    outputs(6163) <= not (a xor b);
    outputs(6164) <= not (a or b);
    outputs(6165) <= a;
    outputs(6166) <= a xor b;
    outputs(6167) <= not (a or b);
    outputs(6168) <= a xor b;
    outputs(6169) <= not (a and b);
    outputs(6170) <= b;
    outputs(6171) <= a xor b;
    outputs(6172) <= not a;
    outputs(6173) <= a and b;
    outputs(6174) <= a xor b;
    outputs(6175) <= b and not a;
    outputs(6176) <= a and not b;
    outputs(6177) <= a and b;
    outputs(6178) <= not a;
    outputs(6179) <= not b;
    outputs(6180) <= not a;
    outputs(6181) <= not a;
    outputs(6182) <= b and not a;
    outputs(6183) <= a;
    outputs(6184) <= not (a xor b);
    outputs(6185) <= a xor b;
    outputs(6186) <= a xor b;
    outputs(6187) <= a xor b;
    outputs(6188) <= a;
    outputs(6189) <= b and not a;
    outputs(6190) <= a and not b;
    outputs(6191) <= not b;
    outputs(6192) <= not b;
    outputs(6193) <= a;
    outputs(6194) <= a xor b;
    outputs(6195) <= not b;
    outputs(6196) <= b;
    outputs(6197) <= a xor b;
    outputs(6198) <= not (a or b);
    outputs(6199) <= b;
    outputs(6200) <= not (a xor b);
    outputs(6201) <= not b;
    outputs(6202) <= not (a xor b);
    outputs(6203) <= b and not a;
    outputs(6204) <= a;
    outputs(6205) <= b;
    outputs(6206) <= a xor b;
    outputs(6207) <= b;
    outputs(6208) <= not a;
    outputs(6209) <= a xor b;
    outputs(6210) <= not (a xor b);
    outputs(6211) <= a and not b;
    outputs(6212) <= b and not a;
    outputs(6213) <= not (a and b);
    outputs(6214) <= a xor b;
    outputs(6215) <= not (a or b);
    outputs(6216) <= a xor b;
    outputs(6217) <= b;
    outputs(6218) <= a and b;
    outputs(6219) <= a;
    outputs(6220) <= not b;
    outputs(6221) <= a xor b;
    outputs(6222) <= a;
    outputs(6223) <= not b;
    outputs(6224) <= a and b;
    outputs(6225) <= not b or a;
    outputs(6226) <= a and b;
    outputs(6227) <= b;
    outputs(6228) <= a and not b;
    outputs(6229) <= a or b;
    outputs(6230) <= not a;
    outputs(6231) <= not (a and b);
    outputs(6232) <= not a;
    outputs(6233) <= a and b;
    outputs(6234) <= a;
    outputs(6235) <= not (a xor b);
    outputs(6236) <= not a;
    outputs(6237) <= a xor b;
    outputs(6238) <= a;
    outputs(6239) <= a and not b;
    outputs(6240) <= a;
    outputs(6241) <= a xor b;
    outputs(6242) <= not (a xor b);
    outputs(6243) <= not (a xor b);
    outputs(6244) <= not (a and b);
    outputs(6245) <= not b or a;
    outputs(6246) <= a xor b;
    outputs(6247) <= not (a xor b);
    outputs(6248) <= not a;
    outputs(6249) <= not (a xor b);
    outputs(6250) <= a and not b;
    outputs(6251) <= not (a xor b);
    outputs(6252) <= a xor b;
    outputs(6253) <= not a;
    outputs(6254) <= b;
    outputs(6255) <= not b;
    outputs(6256) <= not a;
    outputs(6257) <= a and not b;
    outputs(6258) <= not (a xor b);
    outputs(6259) <= not (a xor b);
    outputs(6260) <= b;
    outputs(6261) <= not b;
    outputs(6262) <= not (a xor b);
    outputs(6263) <= a or b;
    outputs(6264) <= not (a xor b);
    outputs(6265) <= a xor b;
    outputs(6266) <= not a;
    outputs(6267) <= a or b;
    outputs(6268) <= not (a xor b);
    outputs(6269) <= a;
    outputs(6270) <= not (a xor b);
    outputs(6271) <= not (a xor b);
    outputs(6272) <= b;
    outputs(6273) <= not (a xor b);
    outputs(6274) <= a;
    outputs(6275) <= b;
    outputs(6276) <= a xor b;
    outputs(6277) <= b;
    outputs(6278) <= b and not a;
    outputs(6279) <= not a;
    outputs(6280) <= a xor b;
    outputs(6281) <= a xor b;
    outputs(6282) <= not (a xor b);
    outputs(6283) <= not a;
    outputs(6284) <= a xor b;
    outputs(6285) <= not (a xor b);
    outputs(6286) <= not (a xor b);
    outputs(6287) <= not a or b;
    outputs(6288) <= b and not a;
    outputs(6289) <= a and not b;
    outputs(6290) <= not (a and b);
    outputs(6291) <= a xor b;
    outputs(6292) <= not (a or b);
    outputs(6293) <= not a or b;
    outputs(6294) <= not b;
    outputs(6295) <= a xor b;
    outputs(6296) <= not a;
    outputs(6297) <= b;
    outputs(6298) <= not b;
    outputs(6299) <= not (a xor b);
    outputs(6300) <= not a;
    outputs(6301) <= not (a xor b);
    outputs(6302) <= not (a xor b);
    outputs(6303) <= a and not b;
    outputs(6304) <= b and not a;
    outputs(6305) <= not (a xor b);
    outputs(6306) <= not b;
    outputs(6307) <= not (a xor b);
    outputs(6308) <= a;
    outputs(6309) <= a xor b;
    outputs(6310) <= a xor b;
    outputs(6311) <= a xor b;
    outputs(6312) <= not (a xor b);
    outputs(6313) <= not (a xor b);
    outputs(6314) <= a xor b;
    outputs(6315) <= a and not b;
    outputs(6316) <= a and b;
    outputs(6317) <= a;
    outputs(6318) <= not a;
    outputs(6319) <= not (a xor b);
    outputs(6320) <= not b;
    outputs(6321) <= not (a xor b);
    outputs(6322) <= not b;
    outputs(6323) <= not b;
    outputs(6324) <= not (a or b);
    outputs(6325) <= not (a xor b);
    outputs(6326) <= b;
    outputs(6327) <= not b;
    outputs(6328) <= not a;
    outputs(6329) <= not b;
    outputs(6330) <= b;
    outputs(6331) <= a xor b;
    outputs(6332) <= not a or b;
    outputs(6333) <= not (a xor b);
    outputs(6334) <= not (a xor b);
    outputs(6335) <= a xor b;
    outputs(6336) <= not b;
    outputs(6337) <= not (a xor b);
    outputs(6338) <= b;
    outputs(6339) <= not (a xor b);
    outputs(6340) <= not (a xor b);
    outputs(6341) <= not b;
    outputs(6342) <= not (a and b);
    outputs(6343) <= not a;
    outputs(6344) <= not (a xor b);
    outputs(6345) <= a xor b;
    outputs(6346) <= b and not a;
    outputs(6347) <= not (a or b);
    outputs(6348) <= a and not b;
    outputs(6349) <= b and not a;
    outputs(6350) <= not (a xor b);
    outputs(6351) <= not a;
    outputs(6352) <= a;
    outputs(6353) <= not (a or b);
    outputs(6354) <= not a;
    outputs(6355) <= a;
    outputs(6356) <= a and b;
    outputs(6357) <= not (a and b);
    outputs(6358) <= b and not a;
    outputs(6359) <= b and not a;
    outputs(6360) <= a and not b;
    outputs(6361) <= not a;
    outputs(6362) <= not (a or b);
    outputs(6363) <= not (a xor b);
    outputs(6364) <= not b;
    outputs(6365) <= a xor b;
    outputs(6366) <= a;
    outputs(6367) <= not b;
    outputs(6368) <= a xor b;
    outputs(6369) <= b;
    outputs(6370) <= not (a xor b);
    outputs(6371) <= not (a xor b);
    outputs(6372) <= b;
    outputs(6373) <= a and b;
    outputs(6374) <= a xor b;
    outputs(6375) <= not b;
    outputs(6376) <= not (a xor b);
    outputs(6377) <= not b;
    outputs(6378) <= b;
    outputs(6379) <= not a;
    outputs(6380) <= not (a xor b);
    outputs(6381) <= a;
    outputs(6382) <= not a or b;
    outputs(6383) <= a or b;
    outputs(6384) <= not a;
    outputs(6385) <= not a;
    outputs(6386) <= not (a xor b);
    outputs(6387) <= a xor b;
    outputs(6388) <= a xor b;
    outputs(6389) <= a xor b;
    outputs(6390) <= a xor b;
    outputs(6391) <= b and not a;
    outputs(6392) <= not (a or b);
    outputs(6393) <= a and not b;
    outputs(6394) <= not a;
    outputs(6395) <= a and b;
    outputs(6396) <= not (a xor b);
    outputs(6397) <= b and not a;
    outputs(6398) <= not (a xor b);
    outputs(6399) <= not b or a;
    outputs(6400) <= a xor b;
    outputs(6401) <= not (a or b);
    outputs(6402) <= not (a and b);
    outputs(6403) <= a xor b;
    outputs(6404) <= a or b;
    outputs(6405) <= a xor b;
    outputs(6406) <= a xor b;
    outputs(6407) <= b;
    outputs(6408) <= a xor b;
    outputs(6409) <= a xor b;
    outputs(6410) <= a xor b;
    outputs(6411) <= not b;
    outputs(6412) <= not b or a;
    outputs(6413) <= not a;
    outputs(6414) <= not b;
    outputs(6415) <= not b or a;
    outputs(6416) <= not b;
    outputs(6417) <= a or b;
    outputs(6418) <= a;
    outputs(6419) <= a xor b;
    outputs(6420) <= a xor b;
    outputs(6421) <= a;
    outputs(6422) <= a and not b;
    outputs(6423) <= a and not b;
    outputs(6424) <= not (a or b);
    outputs(6425) <= not a;
    outputs(6426) <= b;
    outputs(6427) <= a and b;
    outputs(6428) <= not (a and b);
    outputs(6429) <= a;
    outputs(6430) <= not (a and b);
    outputs(6431) <= not (a xor b);
    outputs(6432) <= a;
    outputs(6433) <= a;
    outputs(6434) <= a;
    outputs(6435) <= not a;
    outputs(6436) <= not (a or b);
    outputs(6437) <= a xor b;
    outputs(6438) <= a;
    outputs(6439) <= a xor b;
    outputs(6440) <= not b;
    outputs(6441) <= b;
    outputs(6442) <= b;
    outputs(6443) <= b and not a;
    outputs(6444) <= a xor b;
    outputs(6445) <= b and not a;
    outputs(6446) <= a;
    outputs(6447) <= a;
    outputs(6448) <= a;
    outputs(6449) <= a xor b;
    outputs(6450) <= not a or b;
    outputs(6451) <= a;
    outputs(6452) <= a xor b;
    outputs(6453) <= not a;
    outputs(6454) <= a xor b;
    outputs(6455) <= b;
    outputs(6456) <= a;
    outputs(6457) <= a;
    outputs(6458) <= not b or a;
    outputs(6459) <= b;
    outputs(6460) <= not (a xor b);
    outputs(6461) <= a;
    outputs(6462) <= a xor b;
    outputs(6463) <= not a;
    outputs(6464) <= not (a xor b);
    outputs(6465) <= not (a xor b);
    outputs(6466) <= b and not a;
    outputs(6467) <= a xor b;
    outputs(6468) <= a or b;
    outputs(6469) <= not b or a;
    outputs(6470) <= not a;
    outputs(6471) <= not (a xor b);
    outputs(6472) <= not b;
    outputs(6473) <= not (a xor b);
    outputs(6474) <= a xor b;
    outputs(6475) <= a;
    outputs(6476) <= a;
    outputs(6477) <= not (a xor b);
    outputs(6478) <= a xor b;
    outputs(6479) <= a xor b;
    outputs(6480) <= not a;
    outputs(6481) <= a and not b;
    outputs(6482) <= a and b;
    outputs(6483) <= not b;
    outputs(6484) <= not (a and b);
    outputs(6485) <= a;
    outputs(6486) <= not (a xor b);
    outputs(6487) <= not (a and b);
    outputs(6488) <= not (a and b);
    outputs(6489) <= not (a xor b);
    outputs(6490) <= not (a xor b);
    outputs(6491) <= b;
    outputs(6492) <= not b;
    outputs(6493) <= a xor b;
    outputs(6494) <= b and not a;
    outputs(6495) <= not (a xor b);
    outputs(6496) <= not (a xor b);
    outputs(6497) <= a and b;
    outputs(6498) <= a;
    outputs(6499) <= a xor b;
    outputs(6500) <= a xor b;
    outputs(6501) <= not (a or b);
    outputs(6502) <= not (a xor b);
    outputs(6503) <= not b or a;
    outputs(6504) <= b;
    outputs(6505) <= not a;
    outputs(6506) <= a xor b;
    outputs(6507) <= not b;
    outputs(6508) <= a xor b;
    outputs(6509) <= a;
    outputs(6510) <= not (a and b);
    outputs(6511) <= a xor b;
    outputs(6512) <= not b;
    outputs(6513) <= not (a xor b);
    outputs(6514) <= a xor b;
    outputs(6515) <= a xor b;
    outputs(6516) <= not (a and b);
    outputs(6517) <= b;
    outputs(6518) <= a xor b;
    outputs(6519) <= a xor b;
    outputs(6520) <= not (a xor b);
    outputs(6521) <= not (a xor b);
    outputs(6522) <= a xor b;
    outputs(6523) <= a;
    outputs(6524) <= not (a xor b);
    outputs(6525) <= b;
    outputs(6526) <= a;
    outputs(6527) <= b;
    outputs(6528) <= not b;
    outputs(6529) <= a;
    outputs(6530) <= a xor b;
    outputs(6531) <= a xor b;
    outputs(6532) <= not b or a;
    outputs(6533) <= a xor b;
    outputs(6534) <= not (a xor b);
    outputs(6535) <= not b;
    outputs(6536) <= a xor b;
    outputs(6537) <= b;
    outputs(6538) <= b;
    outputs(6539) <= b;
    outputs(6540) <= not (a xor b);
    outputs(6541) <= a;
    outputs(6542) <= b;
    outputs(6543) <= a;
    outputs(6544) <= not a or b;
    outputs(6545) <= not (a xor b);
    outputs(6546) <= not a;
    outputs(6547) <= a and b;
    outputs(6548) <= b;
    outputs(6549) <= not b;
    outputs(6550) <= a xor b;
    outputs(6551) <= a xor b;
    outputs(6552) <= a or b;
    outputs(6553) <= not a or b;
    outputs(6554) <= not (a or b);
    outputs(6555) <= not (a xor b);
    outputs(6556) <= not (a xor b);
    outputs(6557) <= a xor b;
    outputs(6558) <= not a or b;
    outputs(6559) <= a xor b;
    outputs(6560) <= b;
    outputs(6561) <= a xor b;
    outputs(6562) <= not (a or b);
    outputs(6563) <= not a;
    outputs(6564) <= not a;
    outputs(6565) <= not a;
    outputs(6566) <= a;
    outputs(6567) <= not (a xor b);
    outputs(6568) <= a;
    outputs(6569) <= a xor b;
    outputs(6570) <= a and not b;
    outputs(6571) <= not b or a;
    outputs(6572) <= not (a xor b);
    outputs(6573) <= a or b;
    outputs(6574) <= a or b;
    outputs(6575) <= not (a xor b);
    outputs(6576) <= a xor b;
    outputs(6577) <= not (a xor b);
    outputs(6578) <= a xor b;
    outputs(6579) <= not b;
    outputs(6580) <= not a;
    outputs(6581) <= not (a and b);
    outputs(6582) <= not (a or b);
    outputs(6583) <= a xor b;
    outputs(6584) <= not b;
    outputs(6585) <= not a;
    outputs(6586) <= b;
    outputs(6587) <= not a;
    outputs(6588) <= not a;
    outputs(6589) <= not b;
    outputs(6590) <= a;
    outputs(6591) <= not b;
    outputs(6592) <= a xor b;
    outputs(6593) <= a xor b;
    outputs(6594) <= not (a xor b);
    outputs(6595) <= a or b;
    outputs(6596) <= a and not b;
    outputs(6597) <= not a;
    outputs(6598) <= not a or b;
    outputs(6599) <= a xor b;
    outputs(6600) <= not a;
    outputs(6601) <= b;
    outputs(6602) <= not (a and b);
    outputs(6603) <= a;
    outputs(6604) <= not (a or b);
    outputs(6605) <= not b or a;
    outputs(6606) <= not b;
    outputs(6607) <= not a;
    outputs(6608) <= not b;
    outputs(6609) <= a xor b;
    outputs(6610) <= a and b;
    outputs(6611) <= not (a or b);
    outputs(6612) <= a xor b;
    outputs(6613) <= a;
    outputs(6614) <= not a;
    outputs(6615) <= not (a xor b);
    outputs(6616) <= not (a xor b);
    outputs(6617) <= b;
    outputs(6618) <= not (a xor b);
    outputs(6619) <= a xor b;
    outputs(6620) <= not b or a;
    outputs(6621) <= not (a xor b);
    outputs(6622) <= not (a xor b);
    outputs(6623) <= a;
    outputs(6624) <= a;
    outputs(6625) <= not b or a;
    outputs(6626) <= a xor b;
    outputs(6627) <= a;
    outputs(6628) <= a xor b;
    outputs(6629) <= not a;
    outputs(6630) <= a xor b;
    outputs(6631) <= a xor b;
    outputs(6632) <= b;
    outputs(6633) <= b;
    outputs(6634) <= not (a xor b);
    outputs(6635) <= not (a xor b);
    outputs(6636) <= a xor b;
    outputs(6637) <= not (a xor b);
    outputs(6638) <= not (a or b);
    outputs(6639) <= not (a xor b);
    outputs(6640) <= a and b;
    outputs(6641) <= not b or a;
    outputs(6642) <= not b or a;
    outputs(6643) <= b;
    outputs(6644) <= a xor b;
    outputs(6645) <= a xor b;
    outputs(6646) <= not b;
    outputs(6647) <= a xor b;
    outputs(6648) <= a xor b;
    outputs(6649) <= a xor b;
    outputs(6650) <= not a;
    outputs(6651) <= a xor b;
    outputs(6652) <= not a;
    outputs(6653) <= a xor b;
    outputs(6654) <= b;
    outputs(6655) <= not (a xor b);
    outputs(6656) <= a and not b;
    outputs(6657) <= not (a or b);
    outputs(6658) <= not b;
    outputs(6659) <= not b;
    outputs(6660) <= not a or b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= a and not b;
    outputs(6663) <= a xor b;
    outputs(6664) <= a or b;
    outputs(6665) <= a xor b;
    outputs(6666) <= a or b;
    outputs(6667) <= a and b;
    outputs(6668) <= a xor b;
    outputs(6669) <= a xor b;
    outputs(6670) <= not a or b;
    outputs(6671) <= a or b;
    outputs(6672) <= not b;
    outputs(6673) <= a xor b;
    outputs(6674) <= not a;
    outputs(6675) <= not (a and b);
    outputs(6676) <= b;
    outputs(6677) <= not (a xor b);
    outputs(6678) <= not (a xor b);
    outputs(6679) <= a and not b;
    outputs(6680) <= a xor b;
    outputs(6681) <= a xor b;
    outputs(6682) <= a;
    outputs(6683) <= a and b;
    outputs(6684) <= a or b;
    outputs(6685) <= not a or b;
    outputs(6686) <= a or b;
    outputs(6687) <= not b or a;
    outputs(6688) <= not a;
    outputs(6689) <= a xor b;
    outputs(6690) <= a;
    outputs(6691) <= not b;
    outputs(6692) <= not (a xor b);
    outputs(6693) <= a;
    outputs(6694) <= not b;
    outputs(6695) <= not (a xor b);
    outputs(6696) <= not a or b;
    outputs(6697) <= a and b;
    outputs(6698) <= not a;
    outputs(6699) <= a xor b;
    outputs(6700) <= a and not b;
    outputs(6701) <= not a;
    outputs(6702) <= a;
    outputs(6703) <= not (a xor b);
    outputs(6704) <= a or b;
    outputs(6705) <= a or b;
    outputs(6706) <= not (a xor b);
    outputs(6707) <= a xor b;
    outputs(6708) <= a;
    outputs(6709) <= a;
    outputs(6710) <= not (a xor b);
    outputs(6711) <= b;
    outputs(6712) <= a or b;
    outputs(6713) <= a xor b;
    outputs(6714) <= not a;
    outputs(6715) <= a or b;
    outputs(6716) <= not (a xor b);
    outputs(6717) <= b and not a;
    outputs(6718) <= not b or a;
    outputs(6719) <= not (a or b);
    outputs(6720) <= not b;
    outputs(6721) <= a;
    outputs(6722) <= not a;
    outputs(6723) <= not (a xor b);
    outputs(6724) <= a;
    outputs(6725) <= not (a xor b);
    outputs(6726) <= a or b;
    outputs(6727) <= a;
    outputs(6728) <= a;
    outputs(6729) <= not (a or b);
    outputs(6730) <= b;
    outputs(6731) <= not b;
    outputs(6732) <= a;
    outputs(6733) <= not (a xor b);
    outputs(6734) <= a or b;
    outputs(6735) <= not (a xor b);
    outputs(6736) <= a or b;
    outputs(6737) <= a xor b;
    outputs(6738) <= not b;
    outputs(6739) <= a xor b;
    outputs(6740) <= a xor b;
    outputs(6741) <= a xor b;
    outputs(6742) <= a xor b;
    outputs(6743) <= not (a xor b);
    outputs(6744) <= not a;
    outputs(6745) <= not a;
    outputs(6746) <= a;
    outputs(6747) <= not b;
    outputs(6748) <= not a;
    outputs(6749) <= not (a or b);
    outputs(6750) <= b;
    outputs(6751) <= not b;
    outputs(6752) <= a;
    outputs(6753) <= a xor b;
    outputs(6754) <= a xor b;
    outputs(6755) <= a;
    outputs(6756) <= b;
    outputs(6757) <= a;
    outputs(6758) <= a xor b;
    outputs(6759) <= not a;
    outputs(6760) <= a;
    outputs(6761) <= not (a xor b);
    outputs(6762) <= a or b;
    outputs(6763) <= not (a xor b);
    outputs(6764) <= not (a xor b);
    outputs(6765) <= not a;
    outputs(6766) <= not (a and b);
    outputs(6767) <= not (a or b);
    outputs(6768) <= not (a xor b);
    outputs(6769) <= b;
    outputs(6770) <= not b;
    outputs(6771) <= not a;
    outputs(6772) <= a and not b;
    outputs(6773) <= a and not b;
    outputs(6774) <= not (a xor b);
    outputs(6775) <= not a;
    outputs(6776) <= a or b;
    outputs(6777) <= a and b;
    outputs(6778) <= not (a xor b);
    outputs(6779) <= not b;
    outputs(6780) <= not (a xor b);
    outputs(6781) <= not (a xor b);
    outputs(6782) <= a xor b;
    outputs(6783) <= a;
    outputs(6784) <= not (a xor b);
    outputs(6785) <= a;
    outputs(6786) <= not (a and b);
    outputs(6787) <= not (a or b);
    outputs(6788) <= not (a xor b);
    outputs(6789) <= not a;
    outputs(6790) <= a xor b;
    outputs(6791) <= not (a or b);
    outputs(6792) <= not (a xor b);
    outputs(6793) <= b and not a;
    outputs(6794) <= not a;
    outputs(6795) <= a xor b;
    outputs(6796) <= not (a xor b);
    outputs(6797) <= b;
    outputs(6798) <= not a;
    outputs(6799) <= a;
    outputs(6800) <= not a;
    outputs(6801) <= not b;
    outputs(6802) <= a or b;
    outputs(6803) <= a;
    outputs(6804) <= not a;
    outputs(6805) <= not a or b;
    outputs(6806) <= not (a xor b);
    outputs(6807) <= not (a xor b);
    outputs(6808) <= not b;
    outputs(6809) <= b and not a;
    outputs(6810) <= a and b;
    outputs(6811) <= a or b;
    outputs(6812) <= b;
    outputs(6813) <= not a or b;
    outputs(6814) <= a or b;
    outputs(6815) <= not b;
    outputs(6816) <= b;
    outputs(6817) <= not b;
    outputs(6818) <= b and not a;
    outputs(6819) <= a xor b;
    outputs(6820) <= not (a xor b);
    outputs(6821) <= a xor b;
    outputs(6822) <= a;
    outputs(6823) <= not (a xor b);
    outputs(6824) <= not b or a;
    outputs(6825) <= not (a xor b);
    outputs(6826) <= not (a or b);
    outputs(6827) <= not (a xor b);
    outputs(6828) <= a xor b;
    outputs(6829) <= not a;
    outputs(6830) <= not a;
    outputs(6831) <= not b;
    outputs(6832) <= not a;
    outputs(6833) <= not (a xor b);
    outputs(6834) <= not (a xor b);
    outputs(6835) <= not (a and b);
    outputs(6836) <= not (a xor b);
    outputs(6837) <= a xor b;
    outputs(6838) <= not (a or b);
    outputs(6839) <= not b;
    outputs(6840) <= not a or b;
    outputs(6841) <= a;
    outputs(6842) <= not a;
    outputs(6843) <= not (a xor b);
    outputs(6844) <= b;
    outputs(6845) <= a xor b;
    outputs(6846) <= a;
    outputs(6847) <= not (a xor b);
    outputs(6848) <= a;
    outputs(6849) <= a;
    outputs(6850) <= a and not b;
    outputs(6851) <= not (a xor b);
    outputs(6852) <= not (a xor b);
    outputs(6853) <= not (a or b);
    outputs(6854) <= b and not a;
    outputs(6855) <= a xor b;
    outputs(6856) <= not a or b;
    outputs(6857) <= not a or b;
    outputs(6858) <= not (a or b);
    outputs(6859) <= a xor b;
    outputs(6860) <= a;
    outputs(6861) <= not (a xor b);
    outputs(6862) <= not b;
    outputs(6863) <= b;
    outputs(6864) <= a xor b;
    outputs(6865) <= not a;
    outputs(6866) <= not b;
    outputs(6867) <= not (a or b);
    outputs(6868) <= not b;
    outputs(6869) <= a;
    outputs(6870) <= a xor b;
    outputs(6871) <= a xor b;
    outputs(6872) <= not a;
    outputs(6873) <= not b;
    outputs(6874) <= not b or a;
    outputs(6875) <= not a or b;
    outputs(6876) <= not (a xor b);
    outputs(6877) <= not a or b;
    outputs(6878) <= not (a and b);
    outputs(6879) <= b;
    outputs(6880) <= a and b;
    outputs(6881) <= not (a xor b);
    outputs(6882) <= not b;
    outputs(6883) <= not (a xor b);
    outputs(6884) <= not a;
    outputs(6885) <= a and b;
    outputs(6886) <= b and not a;
    outputs(6887) <= not a;
    outputs(6888) <= not b;
    outputs(6889) <= b and not a;
    outputs(6890) <= a and b;
    outputs(6891) <= a xor b;
    outputs(6892) <= a xor b;
    outputs(6893) <= not (a xor b);
    outputs(6894) <= not b;
    outputs(6895) <= not (a xor b);
    outputs(6896) <= a;
    outputs(6897) <= a xor b;
    outputs(6898) <= a xor b;
    outputs(6899) <= not (a xor b);
    outputs(6900) <= not (a and b);
    outputs(6901) <= a xor b;
    outputs(6902) <= a;
    outputs(6903) <= not (a xor b);
    outputs(6904) <= a and not b;
    outputs(6905) <= a xor b;
    outputs(6906) <= b;
    outputs(6907) <= b;
    outputs(6908) <= not b;
    outputs(6909) <= b;
    outputs(6910) <= b;
    outputs(6911) <= not a;
    outputs(6912) <= not (a or b);
    outputs(6913) <= not (a xor b);
    outputs(6914) <= not a;
    outputs(6915) <= b;
    outputs(6916) <= not (a or b);
    outputs(6917) <= b;
    outputs(6918) <= a and not b;
    outputs(6919) <= a and b;
    outputs(6920) <= not (a xor b);
    outputs(6921) <= not b;
    outputs(6922) <= b;
    outputs(6923) <= b;
    outputs(6924) <= not b;
    outputs(6925) <= a xor b;
    outputs(6926) <= not b;
    outputs(6927) <= a xor b;
    outputs(6928) <= not a;
    outputs(6929) <= not (a or b);
    outputs(6930) <= not (a xor b);
    outputs(6931) <= a xor b;
    outputs(6932) <= not (a xor b);
    outputs(6933) <= not (a or b);
    outputs(6934) <= a xor b;
    outputs(6935) <= a;
    outputs(6936) <= not (a xor b);
    outputs(6937) <= a and not b;
    outputs(6938) <= a;
    outputs(6939) <= not a;
    outputs(6940) <= not b;
    outputs(6941) <= a xor b;
    outputs(6942) <= not (a xor b);
    outputs(6943) <= a;
    outputs(6944) <= a or b;
    outputs(6945) <= not (a xor b);
    outputs(6946) <= b;
    outputs(6947) <= b;
    outputs(6948) <= not a;
    outputs(6949) <= a and not b;
    outputs(6950) <= a;
    outputs(6951) <= a;
    outputs(6952) <= not a;
    outputs(6953) <= b;
    outputs(6954) <= not a;
    outputs(6955) <= not a or b;
    outputs(6956) <= a;
    outputs(6957) <= b;
    outputs(6958) <= b and not a;
    outputs(6959) <= a;
    outputs(6960) <= not a;
    outputs(6961) <= b;
    outputs(6962) <= not a;
    outputs(6963) <= not b;
    outputs(6964) <= a;
    outputs(6965) <= not a;
    outputs(6966) <= b;
    outputs(6967) <= a xor b;
    outputs(6968) <= not (a xor b);
    outputs(6969) <= not b;
    outputs(6970) <= a xor b;
    outputs(6971) <= b;
    outputs(6972) <= b;
    outputs(6973) <= a xor b;
    outputs(6974) <= not (a xor b);
    outputs(6975) <= not (a xor b);
    outputs(6976) <= b;
    outputs(6977) <= not a or b;
    outputs(6978) <= a xor b;
    outputs(6979) <= not b;
    outputs(6980) <= a;
    outputs(6981) <= not b;
    outputs(6982) <= b;
    outputs(6983) <= not (a xor b);
    outputs(6984) <= a;
    outputs(6985) <= a xor b;
    outputs(6986) <= b and not a;
    outputs(6987) <= not b;
    outputs(6988) <= a;
    outputs(6989) <= not a;
    outputs(6990) <= a;
    outputs(6991) <= not b;
    outputs(6992) <= not b;
    outputs(6993) <= a xor b;
    outputs(6994) <= not (a xor b);
    outputs(6995) <= not (a xor b);
    outputs(6996) <= not b;
    outputs(6997) <= not (a xor b);
    outputs(6998) <= not a or b;
    outputs(6999) <= not b;
    outputs(7000) <= not b;
    outputs(7001) <= not b;
    outputs(7002) <= not (a xor b);
    outputs(7003) <= a;
    outputs(7004) <= a and not b;
    outputs(7005) <= not b or a;
    outputs(7006) <= not (a xor b);
    outputs(7007) <= not a;
    outputs(7008) <= not (a xor b);
    outputs(7009) <= b and not a;
    outputs(7010) <= not a or b;
    outputs(7011) <= a xor b;
    outputs(7012) <= not a;
    outputs(7013) <= not b;
    outputs(7014) <= a xor b;
    outputs(7015) <= a;
    outputs(7016) <= a and not b;
    outputs(7017) <= not (a or b);
    outputs(7018) <= a xor b;
    outputs(7019) <= b;
    outputs(7020) <= a;
    outputs(7021) <= not b;
    outputs(7022) <= not (a xor b);
    outputs(7023) <= a;
    outputs(7024) <= b;
    outputs(7025) <= a xor b;
    outputs(7026) <= a xor b;
    outputs(7027) <= a xor b;
    outputs(7028) <= not (a xor b);
    outputs(7029) <= a xor b;
    outputs(7030) <= not a;
    outputs(7031) <= not (a xor b);
    outputs(7032) <= not b;
    outputs(7033) <= b;
    outputs(7034) <= b and not a;
    outputs(7035) <= b;
    outputs(7036) <= not a;
    outputs(7037) <= a and not b;
    outputs(7038) <= not (a xor b);
    outputs(7039) <= not (a xor b);
    outputs(7040) <= a xor b;
    outputs(7041) <= a xor b;
    outputs(7042) <= a and b;
    outputs(7043) <= a xor b;
    outputs(7044) <= not a;
    outputs(7045) <= b;
    outputs(7046) <= not b;
    outputs(7047) <= a xor b;
    outputs(7048) <= a xor b;
    outputs(7049) <= not a;
    outputs(7050) <= not a;
    outputs(7051) <= a xor b;
    outputs(7052) <= a xor b;
    outputs(7053) <= b;
    outputs(7054) <= not (a xor b);
    outputs(7055) <= not b;
    outputs(7056) <= a and not b;
    outputs(7057) <= not b;
    outputs(7058) <= not (a xor b);
    outputs(7059) <= not (a xor b);
    outputs(7060) <= not (a xor b);
    outputs(7061) <= not (a xor b);
    outputs(7062) <= not (a xor b);
    outputs(7063) <= a;
    outputs(7064) <= not (a xor b);
    outputs(7065) <= a xor b;
    outputs(7066) <= a xor b;
    outputs(7067) <= a and not b;
    outputs(7068) <= not b;
    outputs(7069) <= a;
    outputs(7070) <= a;
    outputs(7071) <= a and not b;
    outputs(7072) <= a xor b;
    outputs(7073) <= not b;
    outputs(7074) <= a and not b;
    outputs(7075) <= a and not b;
    outputs(7076) <= not (a xor b);
    outputs(7077) <= not a;
    outputs(7078) <= a xor b;
    outputs(7079) <= a xor b;
    outputs(7080) <= not a or b;
    outputs(7081) <= not (a xor b);
    outputs(7082) <= not (a and b);
    outputs(7083) <= a;
    outputs(7084) <= not b;
    outputs(7085) <= a xor b;
    outputs(7086) <= not a or b;
    outputs(7087) <= a xor b;
    outputs(7088) <= b and not a;
    outputs(7089) <= a and b;
    outputs(7090) <= not (a and b);
    outputs(7091) <= not a or b;
    outputs(7092) <= not (a and b);
    outputs(7093) <= not (a xor b);
    outputs(7094) <= not (a xor b);
    outputs(7095) <= a xor b;
    outputs(7096) <= not b;
    outputs(7097) <= not b;
    outputs(7098) <= a;
    outputs(7099) <= not (a xor b);
    outputs(7100) <= not b;
    outputs(7101) <= not (a xor b);
    outputs(7102) <= not (a xor b);
    outputs(7103) <= a and not b;
    outputs(7104) <= not (a xor b);
    outputs(7105) <= not (a or b);
    outputs(7106) <= not (a xor b);
    outputs(7107) <= a;
    outputs(7108) <= not b;
    outputs(7109) <= b;
    outputs(7110) <= not (a xor b);
    outputs(7111) <= not (a xor b);
    outputs(7112) <= a or b;
    outputs(7113) <= not (a xor b);
    outputs(7114) <= b;
    outputs(7115) <= not (a xor b);
    outputs(7116) <= not a;
    outputs(7117) <= a xor b;
    outputs(7118) <= not a;
    outputs(7119) <= not (a and b);
    outputs(7120) <= b and not a;
    outputs(7121) <= a;
    outputs(7122) <= a;
    outputs(7123) <= not b;
    outputs(7124) <= a xor b;
    outputs(7125) <= a xor b;
    outputs(7126) <= not b;
    outputs(7127) <= a;
    outputs(7128) <= a xor b;
    outputs(7129) <= not (a xor b);
    outputs(7130) <= not (a xor b);
    outputs(7131) <= a xor b;
    outputs(7132) <= not b or a;
    outputs(7133) <= not (a and b);
    outputs(7134) <= not a;
    outputs(7135) <= not a;
    outputs(7136) <= b and not a;
    outputs(7137) <= b;
    outputs(7138) <= not b or a;
    outputs(7139) <= a xor b;
    outputs(7140) <= a;
    outputs(7141) <= not (a or b);
    outputs(7142) <= not a or b;
    outputs(7143) <= not (a xor b);
    outputs(7144) <= a and b;
    outputs(7145) <= not b;
    outputs(7146) <= not (a and b);
    outputs(7147) <= a;
    outputs(7148) <= a;
    outputs(7149) <= not (a xor b);
    outputs(7150) <= not a;
    outputs(7151) <= a;
    outputs(7152) <= not (a xor b);
    outputs(7153) <= not a;
    outputs(7154) <= not b or a;
    outputs(7155) <= not a;
    outputs(7156) <= a xor b;
    outputs(7157) <= not a;
    outputs(7158) <= not b;
    outputs(7159) <= a and b;
    outputs(7160) <= not (a or b);
    outputs(7161) <= a xor b;
    outputs(7162) <= a xor b;
    outputs(7163) <= not (a xor b);
    outputs(7164) <= not (a xor b);
    outputs(7165) <= a xor b;
    outputs(7166) <= b;
    outputs(7167) <= not a;
    outputs(7168) <= b;
    outputs(7169) <= a and b;
    outputs(7170) <= a xor b;
    outputs(7171) <= not (a xor b);
    outputs(7172) <= not (a xor b);
    outputs(7173) <= not a;
    outputs(7174) <= not b or a;
    outputs(7175) <= b;
    outputs(7176) <= a xor b;
    outputs(7177) <= a xor b;
    outputs(7178) <= not (a xor b);
    outputs(7179) <= a xor b;
    outputs(7180) <= not (a and b);
    outputs(7181) <= not (a xor b);
    outputs(7182) <= a or b;
    outputs(7183) <= a;
    outputs(7184) <= not b;
    outputs(7185) <= a and not b;
    outputs(7186) <= b and not a;
    outputs(7187) <= not a;
    outputs(7188) <= a xor b;
    outputs(7189) <= not (a xor b);
    outputs(7190) <= not (a and b);
    outputs(7191) <= not a;
    outputs(7192) <= not b;
    outputs(7193) <= a or b;
    outputs(7194) <= a;
    outputs(7195) <= not b;
    outputs(7196) <= not a;
    outputs(7197) <= not (a xor b);
    outputs(7198) <= a xor b;
    outputs(7199) <= a;
    outputs(7200) <= not (a xor b);
    outputs(7201) <= b;
    outputs(7202) <= a;
    outputs(7203) <= a xor b;
    outputs(7204) <= a xor b;
    outputs(7205) <= not (a and b);
    outputs(7206) <= b;
    outputs(7207) <= not b;
    outputs(7208) <= b;
    outputs(7209) <= a xor b;
    outputs(7210) <= a xor b;
    outputs(7211) <= not a;
    outputs(7212) <= not (a xor b);
    outputs(7213) <= a xor b;
    outputs(7214) <= b;
    outputs(7215) <= a;
    outputs(7216) <= not (a xor b);
    outputs(7217) <= not b;
    outputs(7218) <= a;
    outputs(7219) <= a xor b;
    outputs(7220) <= a and not b;
    outputs(7221) <= a and not b;
    outputs(7222) <= a xor b;
    outputs(7223) <= not a;
    outputs(7224) <= a and not b;
    outputs(7225) <= b;
    outputs(7226) <= a xor b;
    outputs(7227) <= a or b;
    outputs(7228) <= a xor b;
    outputs(7229) <= b;
    outputs(7230) <= a;
    outputs(7231) <= not (a xor b);
    outputs(7232) <= not (a xor b);
    outputs(7233) <= not b;
    outputs(7234) <= a xor b;
    outputs(7235) <= a xor b;
    outputs(7236) <= a;
    outputs(7237) <= b;
    outputs(7238) <= a xor b;
    outputs(7239) <= not (a and b);
    outputs(7240) <= b;
    outputs(7241) <= b and not a;
    outputs(7242) <= b;
    outputs(7243) <= not a;
    outputs(7244) <= not (a xor b);
    outputs(7245) <= not (a or b);
    outputs(7246) <= not a;
    outputs(7247) <= b;
    outputs(7248) <= not b;
    outputs(7249) <= b;
    outputs(7250) <= a xor b;
    outputs(7251) <= a xor b;
    outputs(7252) <= a xor b;
    outputs(7253) <= not (a or b);
    outputs(7254) <= b;
    outputs(7255) <= not (a or b);
    outputs(7256) <= not a;
    outputs(7257) <= b and not a;
    outputs(7258) <= not b;
    outputs(7259) <= not (a xor b);
    outputs(7260) <= a xor b;
    outputs(7261) <= not b;
    outputs(7262) <= not b or a;
    outputs(7263) <= a and not b;
    outputs(7264) <= b;
    outputs(7265) <= not (a xor b);
    outputs(7266) <= a or b;
    outputs(7267) <= a and b;
    outputs(7268) <= a xor b;
    outputs(7269) <= not (a xor b);
    outputs(7270) <= not (a xor b);
    outputs(7271) <= a xor b;
    outputs(7272) <= a;
    outputs(7273) <= not (a xor b);
    outputs(7274) <= not a;
    outputs(7275) <= b;
    outputs(7276) <= not (a xor b);
    outputs(7277) <= not b;
    outputs(7278) <= not (a xor b);
    outputs(7279) <= not b;
    outputs(7280) <= a and not b;
    outputs(7281) <= a;
    outputs(7282) <= b;
    outputs(7283) <= not (a xor b);
    outputs(7284) <= not (a xor b);
    outputs(7285) <= a xor b;
    outputs(7286) <= a xor b;
    outputs(7287) <= not b;
    outputs(7288) <= a;
    outputs(7289) <= a or b;
    outputs(7290) <= not (a xor b);
    outputs(7291) <= not a or b;
    outputs(7292) <= not a or b;
    outputs(7293) <= not (a and b);
    outputs(7294) <= b;
    outputs(7295) <= not b;
    outputs(7296) <= a;
    outputs(7297) <= not a;
    outputs(7298) <= not b;
    outputs(7299) <= not b;
    outputs(7300) <= a or b;
    outputs(7301) <= not (a xor b);
    outputs(7302) <= a xor b;
    outputs(7303) <= not (a xor b);
    outputs(7304) <= not (a xor b);
    outputs(7305) <= a and not b;
    outputs(7306) <= not b;
    outputs(7307) <= not (a xor b);
    outputs(7308) <= a xor b;
    outputs(7309) <= not a;
    outputs(7310) <= a xor b;
    outputs(7311) <= not (a xor b);
    outputs(7312) <= a xor b;
    outputs(7313) <= a;
    outputs(7314) <= b;
    outputs(7315) <= a xor b;
    outputs(7316) <= a or b;
    outputs(7317) <= a and not b;
    outputs(7318) <= not (a or b);
    outputs(7319) <= not (a xor b);
    outputs(7320) <= a;
    outputs(7321) <= a xor b;
    outputs(7322) <= b;
    outputs(7323) <= not a;
    outputs(7324) <= a;
    outputs(7325) <= b;
    outputs(7326) <= not a;
    outputs(7327) <= b;
    outputs(7328) <= not b or a;
    outputs(7329) <= not (a xor b);
    outputs(7330) <= b;
    outputs(7331) <= not (a xor b);
    outputs(7332) <= b and not a;
    outputs(7333) <= not a;
    outputs(7334) <= a and b;
    outputs(7335) <= a xor b;
    outputs(7336) <= not (a xor b);
    outputs(7337) <= not b;
    outputs(7338) <= not a or b;
    outputs(7339) <= not a;
    outputs(7340) <= a or b;
    outputs(7341) <= a xor b;
    outputs(7342) <= b;
    outputs(7343) <= b;
    outputs(7344) <= not (a or b);
    outputs(7345) <= b;
    outputs(7346) <= a xor b;
    outputs(7347) <= not b;
    outputs(7348) <= a;
    outputs(7349) <= a xor b;
    outputs(7350) <= not (a xor b);
    outputs(7351) <= a;
    outputs(7352) <= a xor b;
    outputs(7353) <= a and b;
    outputs(7354) <= not b;
    outputs(7355) <= b and not a;
    outputs(7356) <= a xor b;
    outputs(7357) <= a xor b;
    outputs(7358) <= not (a xor b);
    outputs(7359) <= not a;
    outputs(7360) <= not b;
    outputs(7361) <= a;
    outputs(7362) <= a;
    outputs(7363) <= b;
    outputs(7364) <= not b;
    outputs(7365) <= b;
    outputs(7366) <= not (a xor b);
    outputs(7367) <= not (a or b);
    outputs(7368) <= not (a and b);
    outputs(7369) <= not (a or b);
    outputs(7370) <= not b or a;
    outputs(7371) <= not b or a;
    outputs(7372) <= a or b;
    outputs(7373) <= a;
    outputs(7374) <= not a;
    outputs(7375) <= not a;
    outputs(7376) <= a xor b;
    outputs(7377) <= not b;
    outputs(7378) <= not (a xor b);
    outputs(7379) <= a xor b;
    outputs(7380) <= not b or a;
    outputs(7381) <= not (a xor b);
    outputs(7382) <= not b;
    outputs(7383) <= a;
    outputs(7384) <= a and not b;
    outputs(7385) <= not b;
    outputs(7386) <= a or b;
    outputs(7387) <= not (a xor b);
    outputs(7388) <= not b;
    outputs(7389) <= b;
    outputs(7390) <= not (a xor b);
    outputs(7391) <= not (a xor b);
    outputs(7392) <= not a;
    outputs(7393) <= not (a and b);
    outputs(7394) <= a xor b;
    outputs(7395) <= a xor b;
    outputs(7396) <= not a;
    outputs(7397) <= not a or b;
    outputs(7398) <= not (a xor b);
    outputs(7399) <= not b;
    outputs(7400) <= not b;
    outputs(7401) <= not a;
    outputs(7402) <= not b;
    outputs(7403) <= a xor b;
    outputs(7404) <= not b;
    outputs(7405) <= not b;
    outputs(7406) <= a;
    outputs(7407) <= a xor b;
    outputs(7408) <= not (a xor b);
    outputs(7409) <= not a or b;
    outputs(7410) <= not a;
    outputs(7411) <= a xor b;
    outputs(7412) <= not (a xor b);
    outputs(7413) <= not a;
    outputs(7414) <= a xor b;
    outputs(7415) <= not a or b;
    outputs(7416) <= not b or a;
    outputs(7417) <= a xor b;
    outputs(7418) <= a xor b;
    outputs(7419) <= not (a xor b);
    outputs(7420) <= a or b;
    outputs(7421) <= not b;
    outputs(7422) <= a or b;
    outputs(7423) <= not (a xor b);
    outputs(7424) <= not (a or b);
    outputs(7425) <= b;
    outputs(7426) <= not (a xor b);
    outputs(7427) <= a xor b;
    outputs(7428) <= not a;
    outputs(7429) <= not (a xor b);
    outputs(7430) <= b;
    outputs(7431) <= b;
    outputs(7432) <= b;
    outputs(7433) <= not (a or b);
    outputs(7434) <= not b;
    outputs(7435) <= b;
    outputs(7436) <= b;
    outputs(7437) <= a xor b;
    outputs(7438) <= a;
    outputs(7439) <= not (a xor b);
    outputs(7440) <= not b;
    outputs(7441) <= a xor b;
    outputs(7442) <= not a;
    outputs(7443) <= not b;
    outputs(7444) <= not b or a;
    outputs(7445) <= a;
    outputs(7446) <= a xor b;
    outputs(7447) <= a;
    outputs(7448) <= a or b;
    outputs(7449) <= not (a xor b);
    outputs(7450) <= not b or a;
    outputs(7451) <= a and not b;
    outputs(7452) <= not (a xor b);
    outputs(7453) <= a;
    outputs(7454) <= b;
    outputs(7455) <= b;
    outputs(7456) <= a;
    outputs(7457) <= a xor b;
    outputs(7458) <= not (a xor b);
    outputs(7459) <= not a;
    outputs(7460) <= a xor b;
    outputs(7461) <= b;
    outputs(7462) <= b;
    outputs(7463) <= a;
    outputs(7464) <= not (a and b);
    outputs(7465) <= not b;
    outputs(7466) <= not (a xor b);
    outputs(7467) <= a xor b;
    outputs(7468) <= a xor b;
    outputs(7469) <= a xor b;
    outputs(7470) <= b;
    outputs(7471) <= a xor b;
    outputs(7472) <= not (a xor b);
    outputs(7473) <= a xor b;
    outputs(7474) <= not (a xor b);
    outputs(7475) <= a xor b;
    outputs(7476) <= b;
    outputs(7477) <= not a;
    outputs(7478) <= not (a xor b);
    outputs(7479) <= a;
    outputs(7480) <= a xor b;
    outputs(7481) <= a;
    outputs(7482) <= a xor b;
    outputs(7483) <= not b or a;
    outputs(7484) <= a and b;
    outputs(7485) <= a;
    outputs(7486) <= not (a xor b);
    outputs(7487) <= not (a xor b);
    outputs(7488) <= not (a or b);
    outputs(7489) <= not a or b;
    outputs(7490) <= not b;
    outputs(7491) <= a;
    outputs(7492) <= a xor b;
    outputs(7493) <= not (a xor b);
    outputs(7494) <= not a or b;
    outputs(7495) <= b;
    outputs(7496) <= not a;
    outputs(7497) <= not b;
    outputs(7498) <= a or b;
    outputs(7499) <= not (a xor b);
    outputs(7500) <= not (a and b);
    outputs(7501) <= b;
    outputs(7502) <= b;
    outputs(7503) <= a xor b;
    outputs(7504) <= b;
    outputs(7505) <= a and not b;
    outputs(7506) <= b;
    outputs(7507) <= not b or a;
    outputs(7508) <= a xor b;
    outputs(7509) <= not (a and b);
    outputs(7510) <= a or b;
    outputs(7511) <= a xor b;
    outputs(7512) <= not a;
    outputs(7513) <= not b or a;
    outputs(7514) <= a xor b;
    outputs(7515) <= a;
    outputs(7516) <= b;
    outputs(7517) <= a or b;
    outputs(7518) <= not a;
    outputs(7519) <= not b or a;
    outputs(7520) <= b;
    outputs(7521) <= not b;
    outputs(7522) <= not b;
    outputs(7523) <= a and b;
    outputs(7524) <= a xor b;
    outputs(7525) <= not (a xor b);
    outputs(7526) <= not b or a;
    outputs(7527) <= a xor b;
    outputs(7528) <= not (a or b);
    outputs(7529) <= not b;
    outputs(7530) <= not b;
    outputs(7531) <= b;
    outputs(7532) <= not a;
    outputs(7533) <= a xor b;
    outputs(7534) <= not (a or b);
    outputs(7535) <= a;
    outputs(7536) <= b;
    outputs(7537) <= not a;
    outputs(7538) <= not (a xor b);
    outputs(7539) <= not (a xor b);
    outputs(7540) <= a xor b;
    outputs(7541) <= not (a xor b);
    outputs(7542) <= not (a xor b);
    outputs(7543) <= not (a xor b);
    outputs(7544) <= b;
    outputs(7545) <= not a;
    outputs(7546) <= a;
    outputs(7547) <= b and not a;
    outputs(7548) <= not (a xor b);
    outputs(7549) <= a;
    outputs(7550) <= not a;
    outputs(7551) <= a and not b;
    outputs(7552) <= not (a or b);
    outputs(7553) <= a xor b;
    outputs(7554) <= not (a xor b);
    outputs(7555) <= not b or a;
    outputs(7556) <= not b;
    outputs(7557) <= a xor b;
    outputs(7558) <= not a;
    outputs(7559) <= not b;
    outputs(7560) <= not a;
    outputs(7561) <= b;
    outputs(7562) <= not a;
    outputs(7563) <= a xor b;
    outputs(7564) <= not b;
    outputs(7565) <= b;
    outputs(7566) <= not b or a;
    outputs(7567) <= not (a xor b);
    outputs(7568) <= a xor b;
    outputs(7569) <= a;
    outputs(7570) <= not b;
    outputs(7571) <= not b;
    outputs(7572) <= not b or a;
    outputs(7573) <= not b;
    outputs(7574) <= a;
    outputs(7575) <= not b;
    outputs(7576) <= a xor b;
    outputs(7577) <= b and not a;
    outputs(7578) <= not a;
    outputs(7579) <= not b or a;
    outputs(7580) <= a;
    outputs(7581) <= not b or a;
    outputs(7582) <= not (a xor b);
    outputs(7583) <= b;
    outputs(7584) <= a xor b;
    outputs(7585) <= b;
    outputs(7586) <= a and b;
    outputs(7587) <= b and not a;
    outputs(7588) <= not (a or b);
    outputs(7589) <= not (a xor b);
    outputs(7590) <= not (a xor b);
    outputs(7591) <= a xor b;
    outputs(7592) <= not (a xor b);
    outputs(7593) <= not a;
    outputs(7594) <= not (a xor b);
    outputs(7595) <= not b;
    outputs(7596) <= not (a xor b);
    outputs(7597) <= a;
    outputs(7598) <= b;
    outputs(7599) <= a xor b;
    outputs(7600) <= not (a xor b);
    outputs(7601) <= not (a and b);
    outputs(7602) <= a xor b;
    outputs(7603) <= a or b;
    outputs(7604) <= not (a xor b);
    outputs(7605) <= not (a xor b);
    outputs(7606) <= not (a xor b);
    outputs(7607) <= not (a or b);
    outputs(7608) <= not (a xor b);
    outputs(7609) <= a;
    outputs(7610) <= not b;
    outputs(7611) <= not (a or b);
    outputs(7612) <= not (a and b);
    outputs(7613) <= b;
    outputs(7614) <= a;
    outputs(7615) <= not a;
    outputs(7616) <= not b;
    outputs(7617) <= not (a xor b);
    outputs(7618) <= b;
    outputs(7619) <= a xor b;
    outputs(7620) <= not b;
    outputs(7621) <= a;
    outputs(7622) <= a xor b;
    outputs(7623) <= not (a xor b);
    outputs(7624) <= a xor b;
    outputs(7625) <= a and b;
    outputs(7626) <= a xor b;
    outputs(7627) <= a xor b;
    outputs(7628) <= not b or a;
    outputs(7629) <= a or b;
    outputs(7630) <= not (a xor b);
    outputs(7631) <= not a;
    outputs(7632) <= b and not a;
    outputs(7633) <= a xor b;
    outputs(7634) <= not a;
    outputs(7635) <= not b or a;
    outputs(7636) <= a xor b;
    outputs(7637) <= not (a xor b);
    outputs(7638) <= not (a or b);
    outputs(7639) <= not (a and b);
    outputs(7640) <= a and not b;
    outputs(7641) <= not (a xor b);
    outputs(7642) <= a xor b;
    outputs(7643) <= b and not a;
    outputs(7644) <= a;
    outputs(7645) <= not b;
    outputs(7646) <= not (a and b);
    outputs(7647) <= not b;
    outputs(7648) <= not (a xor b);
    outputs(7649) <= a xor b;
    outputs(7650) <= not (a xor b);
    outputs(7651) <= not (a and b);
    outputs(7652) <= b and not a;
    outputs(7653) <= a;
    outputs(7654) <= not b;
    outputs(7655) <= b;
    outputs(7656) <= not b;
    outputs(7657) <= a and not b;
    outputs(7658) <= not b;
    outputs(7659) <= a xor b;
    outputs(7660) <= not (a xor b);
    outputs(7661) <= a;
    outputs(7662) <= a xor b;
    outputs(7663) <= not a;
    outputs(7664) <= a;
    outputs(7665) <= a;
    outputs(7666) <= a;
    outputs(7667) <= not (a xor b);
    outputs(7668) <= b;
    outputs(7669) <= a;
    outputs(7670) <= not (a xor b);
    outputs(7671) <= not (a xor b);
    outputs(7672) <= not (a xor b);
    outputs(7673) <= a;
    outputs(7674) <= not a;
    outputs(7675) <= b;
    outputs(7676) <= b;
    outputs(7677) <= not (a xor b);
    outputs(7678) <= not b;
    outputs(7679) <= a xor b;
    outputs(7680) <= b;
    outputs(7681) <= not a;
    outputs(7682) <= a;
    outputs(7683) <= not b;
    outputs(7684) <= not a or b;
    outputs(7685) <= not a;
    outputs(7686) <= not b;
    outputs(7687) <= not (a xor b);
    outputs(7688) <= a xor b;
    outputs(7689) <= b;
    outputs(7690) <= a xor b;
    outputs(7691) <= not (a xor b);
    outputs(7692) <= a;
    outputs(7693) <= not (a xor b);
    outputs(7694) <= not (a xor b);
    outputs(7695) <= not (a xor b);
    outputs(7696) <= not b;
    outputs(7697) <= a xor b;
    outputs(7698) <= not b;
    outputs(7699) <= a or b;
    outputs(7700) <= a and not b;
    outputs(7701) <= a and b;
    outputs(7702) <= a or b;
    outputs(7703) <= not a;
    outputs(7704) <= not b or a;
    outputs(7705) <= not b;
    outputs(7706) <= a;
    outputs(7707) <= not (a and b);
    outputs(7708) <= a;
    outputs(7709) <= a xor b;
    outputs(7710) <= not (a xor b);
    outputs(7711) <= not a or b;
    outputs(7712) <= a;
    outputs(7713) <= a xor b;
    outputs(7714) <= not b;
    outputs(7715) <= a and not b;
    outputs(7716) <= b;
    outputs(7717) <= b;
    outputs(7718) <= not (a xor b);
    outputs(7719) <= b;
    outputs(7720) <= a and not b;
    outputs(7721) <= a xor b;
    outputs(7722) <= a xor b;
    outputs(7723) <= a xor b;
    outputs(7724) <= not (a xor b);
    outputs(7725) <= not (a xor b);
    outputs(7726) <= not (a xor b);
    outputs(7727) <= b;
    outputs(7728) <= not a or b;
    outputs(7729) <= a and not b;
    outputs(7730) <= not b;
    outputs(7731) <= not (a xor b);
    outputs(7732) <= not b or a;
    outputs(7733) <= a xor b;
    outputs(7734) <= a xor b;
    outputs(7735) <= b and not a;
    outputs(7736) <= a xor b;
    outputs(7737) <= a or b;
    outputs(7738) <= not (a xor b);
    outputs(7739) <= a and b;
    outputs(7740) <= not b;
    outputs(7741) <= not a or b;
    outputs(7742) <= not b;
    outputs(7743) <= b and not a;
    outputs(7744) <= b;
    outputs(7745) <= a xor b;
    outputs(7746) <= not b;
    outputs(7747) <= a and b;
    outputs(7748) <= not (a and b);
    outputs(7749) <= a and b;
    outputs(7750) <= not a;
    outputs(7751) <= not (a xor b);
    outputs(7752) <= not (a xor b);
    outputs(7753) <= a and b;
    outputs(7754) <= b;
    outputs(7755) <= a xor b;
    outputs(7756) <= not b;
    outputs(7757) <= not (a xor b);
    outputs(7758) <= not b;
    outputs(7759) <= a;
    outputs(7760) <= not (a xor b);
    outputs(7761) <= a;
    outputs(7762) <= b;
    outputs(7763) <= not b;
    outputs(7764) <= a or b;
    outputs(7765) <= not b;
    outputs(7766) <= b;
    outputs(7767) <= a;
    outputs(7768) <= not (a xor b);
    outputs(7769) <= not b;
    outputs(7770) <= not (a xor b);
    outputs(7771) <= b and not a;
    outputs(7772) <= a;
    outputs(7773) <= not (a or b);
    outputs(7774) <= not (a xor b);
    outputs(7775) <= not a;
    outputs(7776) <= b;
    outputs(7777) <= b;
    outputs(7778) <= b and not a;
    outputs(7779) <= not (a xor b);
    outputs(7780) <= not b;
    outputs(7781) <= not a;
    outputs(7782) <= a xor b;
    outputs(7783) <= not b or a;
    outputs(7784) <= a and b;
    outputs(7785) <= not (a xor b);
    outputs(7786) <= not (a xor b);
    outputs(7787) <= not (a xor b);
    outputs(7788) <= a xor b;
    outputs(7789) <= a and b;
    outputs(7790) <= not (a or b);
    outputs(7791) <= b and not a;
    outputs(7792) <= a;
    outputs(7793) <= b and not a;
    outputs(7794) <= a;
    outputs(7795) <= a and not b;
    outputs(7796) <= not b;
    outputs(7797) <= not (a or b);
    outputs(7798) <= not a or b;
    outputs(7799) <= not (a xor b);
    outputs(7800) <= a xor b;
    outputs(7801) <= a;
    outputs(7802) <= a and b;
    outputs(7803) <= not a;
    outputs(7804) <= not (a xor b);
    outputs(7805) <= a;
    outputs(7806) <= not (a xor b);
    outputs(7807) <= a and b;
    outputs(7808) <= a xor b;
    outputs(7809) <= not (a xor b);
    outputs(7810) <= not b;
    outputs(7811) <= not (a or b);
    outputs(7812) <= a and b;
    outputs(7813) <= b;
    outputs(7814) <= not (a xor b);
    outputs(7815) <= not (a xor b);
    outputs(7816) <= a;
    outputs(7817) <= not b or a;
    outputs(7818) <= a;
    outputs(7819) <= not a;
    outputs(7820) <= not b;
    outputs(7821) <= a xor b;
    outputs(7822) <= not (a or b);
    outputs(7823) <= a xor b;
    outputs(7824) <= not (a xor b);
    outputs(7825) <= b;
    outputs(7826) <= not (a xor b);
    outputs(7827) <= not b;
    outputs(7828) <= not (a xor b);
    outputs(7829) <= not b;
    outputs(7830) <= b;
    outputs(7831) <= a xor b;
    outputs(7832) <= a xor b;
    outputs(7833) <= not b;
    outputs(7834) <= b and not a;
    outputs(7835) <= not a;
    outputs(7836) <= b;
    outputs(7837) <= not a;
    outputs(7838) <= a and b;
    outputs(7839) <= not b;
    outputs(7840) <= b;
    outputs(7841) <= not (a xor b);
    outputs(7842) <= a and not b;
    outputs(7843) <= not a;
    outputs(7844) <= a;
    outputs(7845) <= b and not a;
    outputs(7846) <= not (a or b);
    outputs(7847) <= not a;
    outputs(7848) <= a;
    outputs(7849) <= not b;
    outputs(7850) <= not b;
    outputs(7851) <= a and b;
    outputs(7852) <= not (a xor b);
    outputs(7853) <= not (a and b);
    outputs(7854) <= not (a xor b);
    outputs(7855) <= b;
    outputs(7856) <= not (a xor b);
    outputs(7857) <= not b;
    outputs(7858) <= a;
    outputs(7859) <= not a;
    outputs(7860) <= not a;
    outputs(7861) <= not b;
    outputs(7862) <= b and not a;
    outputs(7863) <= not a;
    outputs(7864) <= a;
    outputs(7865) <= not a;
    outputs(7866) <= not b;
    outputs(7867) <= a xor b;
    outputs(7868) <= not (a xor b);
    outputs(7869) <= not b;
    outputs(7870) <= not b or a;
    outputs(7871) <= a xor b;
    outputs(7872) <= a and not b;
    outputs(7873) <= a and b;
    outputs(7874) <= not a or b;
    outputs(7875) <= not (a xor b);
    outputs(7876) <= not a;
    outputs(7877) <= a and b;
    outputs(7878) <= b;
    outputs(7879) <= not (a xor b);
    outputs(7880) <= a and b;
    outputs(7881) <= not (a xor b);
    outputs(7882) <= a xor b;
    outputs(7883) <= a and not b;
    outputs(7884) <= not a;
    outputs(7885) <= a;
    outputs(7886) <= a xor b;
    outputs(7887) <= a;
    outputs(7888) <= a;
    outputs(7889) <= a and b;
    outputs(7890) <= a and not b;
    outputs(7891) <= a xor b;
    outputs(7892) <= b;
    outputs(7893) <= a xor b;
    outputs(7894) <= a and b;
    outputs(7895) <= not a;
    outputs(7896) <= a;
    outputs(7897) <= not b;
    outputs(7898) <= a and not b;
    outputs(7899) <= a;
    outputs(7900) <= not b;
    outputs(7901) <= a xor b;
    outputs(7902) <= not (a xor b);
    outputs(7903) <= a xor b;
    outputs(7904) <= a;
    outputs(7905) <= a xor b;
    outputs(7906) <= not (a xor b);
    outputs(7907) <= b;
    outputs(7908) <= not (a xor b);
    outputs(7909) <= b;
    outputs(7910) <= a;
    outputs(7911) <= a;
    outputs(7912) <= not (a or b);
    outputs(7913) <= a and not b;
    outputs(7914) <= not a;
    outputs(7915) <= b;
    outputs(7916) <= a and b;
    outputs(7917) <= a and not b;
    outputs(7918) <= not (a xor b);
    outputs(7919) <= a and b;
    outputs(7920) <= a and not b;
    outputs(7921) <= not a or b;
    outputs(7922) <= b;
    outputs(7923) <= a xor b;
    outputs(7924) <= a;
    outputs(7925) <= not (a xor b);
    outputs(7926) <= a xor b;
    outputs(7927) <= a and not b;
    outputs(7928) <= not a;
    outputs(7929) <= b;
    outputs(7930) <= a xor b;
    outputs(7931) <= not (a xor b);
    outputs(7932) <= b;
    outputs(7933) <= not b;
    outputs(7934) <= not a;
    outputs(7935) <= not (a xor b);
    outputs(7936) <= a and not b;
    outputs(7937) <= b and not a;
    outputs(7938) <= not b;
    outputs(7939) <= b;
    outputs(7940) <= a xor b;
    outputs(7941) <= not (a xor b);
    outputs(7942) <= not b;
    outputs(7943) <= a;
    outputs(7944) <= a and b;
    outputs(7945) <= not (a or b);
    outputs(7946) <= not (a xor b);
    outputs(7947) <= b;
    outputs(7948) <= b;
    outputs(7949) <= a xor b;
    outputs(7950) <= a xor b;
    outputs(7951) <= a;
    outputs(7952) <= not b or a;
    outputs(7953) <= not b;
    outputs(7954) <= not (a or b);
    outputs(7955) <= a or b;
    outputs(7956) <= b;
    outputs(7957) <= a or b;
    outputs(7958) <= a;
    outputs(7959) <= b and not a;
    outputs(7960) <= not (a or b);
    outputs(7961) <= not (a or b);
    outputs(7962) <= a xor b;
    outputs(7963) <= a and b;
    outputs(7964) <= not (a xor b);
    outputs(7965) <= not (a xor b);
    outputs(7966) <= a;
    outputs(7967) <= not (a xor b);
    outputs(7968) <= a;
    outputs(7969) <= not a;
    outputs(7970) <= a and not b;
    outputs(7971) <= not a;
    outputs(7972) <= a;
    outputs(7973) <= a xor b;
    outputs(7974) <= b;
    outputs(7975) <= not b;
    outputs(7976) <= a and b;
    outputs(7977) <= a xor b;
    outputs(7978) <= b;
    outputs(7979) <= not (a or b);
    outputs(7980) <= a;
    outputs(7981) <= not a;
    outputs(7982) <= a;
    outputs(7983) <= b;
    outputs(7984) <= not (a xor b);
    outputs(7985) <= b and not a;
    outputs(7986) <= a and b;
    outputs(7987) <= a xor b;
    outputs(7988) <= not b;
    outputs(7989) <= a;
    outputs(7990) <= not b;
    outputs(7991) <= a;
    outputs(7992) <= not a or b;
    outputs(7993) <= not a;
    outputs(7994) <= not a;
    outputs(7995) <= a;
    outputs(7996) <= not a;
    outputs(7997) <= not b;
    outputs(7998) <= not b;
    outputs(7999) <= b;
    outputs(8000) <= not (a xor b);
    outputs(8001) <= b and not a;
    outputs(8002) <= a;
    outputs(8003) <= not (a or b);
    outputs(8004) <= b;
    outputs(8005) <= not a;
    outputs(8006) <= a xor b;
    outputs(8007) <= a;
    outputs(8008) <= a;
    outputs(8009) <= not (a xor b);
    outputs(8010) <= not a or b;
    outputs(8011) <= not a;
    outputs(8012) <= a xor b;
    outputs(8013) <= a;
    outputs(8014) <= b;
    outputs(8015) <= not (a or b);
    outputs(8016) <= b;
    outputs(8017) <= not (a xor b);
    outputs(8018) <= a;
    outputs(8019) <= a xor b;
    outputs(8020) <= not (a xor b);
    outputs(8021) <= not (a xor b);
    outputs(8022) <= not (a xor b);
    outputs(8023) <= not a;
    outputs(8024) <= a;
    outputs(8025) <= not (a or b);
    outputs(8026) <= a;
    outputs(8027) <= a;
    outputs(8028) <= a and not b;
    outputs(8029) <= b;
    outputs(8030) <= not a;
    outputs(8031) <= not (a xor b);
    outputs(8032) <= not (a xor b);
    outputs(8033) <= a and b;
    outputs(8034) <= b;
    outputs(8035) <= not b;
    outputs(8036) <= not a;
    outputs(8037) <= b;
    outputs(8038) <= not a;
    outputs(8039) <= a or b;
    outputs(8040) <= not a;
    outputs(8041) <= not b;
    outputs(8042) <= not a;
    outputs(8043) <= not a;
    outputs(8044) <= not a;
    outputs(8045) <= a;
    outputs(8046) <= a xor b;
    outputs(8047) <= a xor b;
    outputs(8048) <= not (a xor b);
    outputs(8049) <= not a;
    outputs(8050) <= a xor b;
    outputs(8051) <= b and not a;
    outputs(8052) <= a xor b;
    outputs(8053) <= b;
    outputs(8054) <= not a or b;
    outputs(8055) <= b and not a;
    outputs(8056) <= a xor b;
    outputs(8057) <= not a;
    outputs(8058) <= a and not b;
    outputs(8059) <= not a;
    outputs(8060) <= a and b;
    outputs(8061) <= not b;
    outputs(8062) <= not (a or b);
    outputs(8063) <= not (a or b);
    outputs(8064) <= not (a and b);
    outputs(8065) <= b;
    outputs(8066) <= not (a xor b);
    outputs(8067) <= b;
    outputs(8068) <= b;
    outputs(8069) <= a xor b;
    outputs(8070) <= a;
    outputs(8071) <= not a;
    outputs(8072) <= not b;
    outputs(8073) <= not (a or b);
    outputs(8074) <= not b;
    outputs(8075) <= not b;
    outputs(8076) <= a xor b;
    outputs(8077) <= not b;
    outputs(8078) <= not a;
    outputs(8079) <= a;
    outputs(8080) <= not (a or b);
    outputs(8081) <= a xor b;
    outputs(8082) <= a xor b;
    outputs(8083) <= not b or a;
    outputs(8084) <= a xor b;
    outputs(8085) <= b;
    outputs(8086) <= a xor b;
    outputs(8087) <= not (a or b);
    outputs(8088) <= not a;
    outputs(8089) <= not (a and b);
    outputs(8090) <= not a;
    outputs(8091) <= a and b;
    outputs(8092) <= a and not b;
    outputs(8093) <= not (a xor b);
    outputs(8094) <= a;
    outputs(8095) <= a;
    outputs(8096) <= not a;
    outputs(8097) <= not (a xor b);
    outputs(8098) <= a and not b;
    outputs(8099) <= a xor b;
    outputs(8100) <= a xor b;
    outputs(8101) <= not b;
    outputs(8102) <= a;
    outputs(8103) <= not a;
    outputs(8104) <= not (a xor b);
    outputs(8105) <= not a or b;
    outputs(8106) <= a;
    outputs(8107) <= a;
    outputs(8108) <= b;
    outputs(8109) <= a xor b;
    outputs(8110) <= not a;
    outputs(8111) <= not (a xor b);
    outputs(8112) <= a;
    outputs(8113) <= a;
    outputs(8114) <= a;
    outputs(8115) <= b;
    outputs(8116) <= not (a or b);
    outputs(8117) <= not (a or b);
    outputs(8118) <= not a;
    outputs(8119) <= b;
    outputs(8120) <= not b or a;
    outputs(8121) <= not b;
    outputs(8122) <= b;
    outputs(8123) <= b and not a;
    outputs(8124) <= not b;
    outputs(8125) <= not a;
    outputs(8126) <= a;
    outputs(8127) <= a;
    outputs(8128) <= not (a xor b);
    outputs(8129) <= a xor b;
    outputs(8130) <= not (a or b);
    outputs(8131) <= a;
    outputs(8132) <= not b;
    outputs(8133) <= a xor b;
    outputs(8134) <= not b;
    outputs(8135) <= a;
    outputs(8136) <= a;
    outputs(8137) <= not a;
    outputs(8138) <= not b;
    outputs(8139) <= not b or a;
    outputs(8140) <= b;
    outputs(8141) <= a;
    outputs(8142) <= a;
    outputs(8143) <= not (a xor b);
    outputs(8144) <= not a or b;
    outputs(8145) <= a;
    outputs(8146) <= not (a xor b);
    outputs(8147) <= b and not a;
    outputs(8148) <= not (a xor b);
    outputs(8149) <= b and not a;
    outputs(8150) <= a xor b;
    outputs(8151) <= a and b;
    outputs(8152) <= a xor b;
    outputs(8153) <= a xor b;
    outputs(8154) <= a;
    outputs(8155) <= a;
    outputs(8156) <= b;
    outputs(8157) <= a xor b;
    outputs(8158) <= b;
    outputs(8159) <= a xor b;
    outputs(8160) <= b;
    outputs(8161) <= a xor b;
    outputs(8162) <= not b;
    outputs(8163) <= a and not b;
    outputs(8164) <= b;
    outputs(8165) <= b;
    outputs(8166) <= not (a xor b);
    outputs(8167) <= a and b;
    outputs(8168) <= not (a or b);
    outputs(8169) <= not (a xor b);
    outputs(8170) <= a;
    outputs(8171) <= a and not b;
    outputs(8172) <= a xor b;
    outputs(8173) <= a and not b;
    outputs(8174) <= not (a or b);
    outputs(8175) <= a xor b;
    outputs(8176) <= b;
    outputs(8177) <= not a or b;
    outputs(8178) <= not b;
    outputs(8179) <= not a;
    outputs(8180) <= a xor b;
    outputs(8181) <= not a;
    outputs(8182) <= not (a xor b);
    outputs(8183) <= not a;
    outputs(8184) <= not a or b;
    outputs(8185) <= a;
    outputs(8186) <= a and b;
    outputs(8187) <= a;
    outputs(8188) <= a;
    outputs(8189) <= a and b;
    outputs(8190) <= not b;
    outputs(8191) <= not a;
    outputs(8192) <= not b;
    outputs(8193) <= not b;
    outputs(8194) <= a xor b;
    outputs(8195) <= a;
    outputs(8196) <= not (a xor b);
    outputs(8197) <= not a;
    outputs(8198) <= not a or b;
    outputs(8199) <= not b or a;
    outputs(8200) <= not (a xor b);
    outputs(8201) <= not (a and b);
    outputs(8202) <= not b;
    outputs(8203) <= a;
    outputs(8204) <= not b;
    outputs(8205) <= a and not b;
    outputs(8206) <= a;
    outputs(8207) <= a xor b;
    outputs(8208) <= b;
    outputs(8209) <= a and b;
    outputs(8210) <= not (a and b);
    outputs(8211) <= b and not a;
    outputs(8212) <= not (a xor b);
    outputs(8213) <= a and b;
    outputs(8214) <= not a;
    outputs(8215) <= not (a xor b);
    outputs(8216) <= a xor b;
    outputs(8217) <= not (a and b);
    outputs(8218) <= not b;
    outputs(8219) <= not (a xor b);
    outputs(8220) <= b;
    outputs(8221) <= a xor b;
    outputs(8222) <= not (a xor b);
    outputs(8223) <= not b;
    outputs(8224) <= not b or a;
    outputs(8225) <= not (a xor b);
    outputs(8226) <= b and not a;
    outputs(8227) <= a and b;
    outputs(8228) <= a;
    outputs(8229) <= not b;
    outputs(8230) <= a and b;
    outputs(8231) <= b and not a;
    outputs(8232) <= not (a and b);
    outputs(8233) <= not a;
    outputs(8234) <= not (a xor b);
    outputs(8235) <= not (a or b);
    outputs(8236) <= not b;
    outputs(8237) <= a xor b;
    outputs(8238) <= b;
    outputs(8239) <= not (a or b);
    outputs(8240) <= not a;
    outputs(8241) <= not a;
    outputs(8242) <= not (a or b);
    outputs(8243) <= a;
    outputs(8244) <= a xor b;
    outputs(8245) <= not (a xor b);
    outputs(8246) <= not b;
    outputs(8247) <= not b;
    outputs(8248) <= not a or b;
    outputs(8249) <= a;
    outputs(8250) <= b;
    outputs(8251) <= a or b;
    outputs(8252) <= b and not a;
    outputs(8253) <= not b;
    outputs(8254) <= b;
    outputs(8255) <= b and not a;
    outputs(8256) <= not (a and b);
    outputs(8257) <= not a;
    outputs(8258) <= not (a or b);
    outputs(8259) <= not a;
    outputs(8260) <= a;
    outputs(8261) <= not (a xor b);
    outputs(8262) <= a and not b;
    outputs(8263) <= not (a xor b);
    outputs(8264) <= not a;
    outputs(8265) <= a;
    outputs(8266) <= not (a xor b);
    outputs(8267) <= b;
    outputs(8268) <= a or b;
    outputs(8269) <= a and not b;
    outputs(8270) <= b;
    outputs(8271) <= a xor b;
    outputs(8272) <= not (a xor b);
    outputs(8273) <= not a;
    outputs(8274) <= not b;
    outputs(8275) <= a;
    outputs(8276) <= not b or a;
    outputs(8277) <= a and b;
    outputs(8278) <= not (a and b);
    outputs(8279) <= a xor b;
    outputs(8280) <= not (a or b);
    outputs(8281) <= not b;
    outputs(8282) <= not b;
    outputs(8283) <= b and not a;
    outputs(8284) <= not (a xor b);
    outputs(8285) <= a;
    outputs(8286) <= not (a or b);
    outputs(8287) <= not (a and b);
    outputs(8288) <= b;
    outputs(8289) <= a xor b;
    outputs(8290) <= not b;
    outputs(8291) <= not (a xor b);
    outputs(8292) <= not b;
    outputs(8293) <= not (a xor b);
    outputs(8294) <= not (a xor b);
    outputs(8295) <= not (a xor b);
    outputs(8296) <= a and not b;
    outputs(8297) <= not b or a;
    outputs(8298) <= a xor b;
    outputs(8299) <= a and b;
    outputs(8300) <= not (a or b);
    outputs(8301) <= b;
    outputs(8302) <= a and not b;
    outputs(8303) <= not b or a;
    outputs(8304) <= a xor b;
    outputs(8305) <= a xor b;
    outputs(8306) <= not a;
    outputs(8307) <= not a or b;
    outputs(8308) <= not b;
    outputs(8309) <= a xor b;
    outputs(8310) <= not (a xor b);
    outputs(8311) <= not a;
    outputs(8312) <= a;
    outputs(8313) <= a;
    outputs(8314) <= a;
    outputs(8315) <= b;
    outputs(8316) <= not (a xor b);
    outputs(8317) <= not (a or b);
    outputs(8318) <= not b;
    outputs(8319) <= a and b;
    outputs(8320) <= not (a xor b);
    outputs(8321) <= b and not a;
    outputs(8322) <= b;
    outputs(8323) <= b;
    outputs(8324) <= a;
    outputs(8325) <= not b;
    outputs(8326) <= a or b;
    outputs(8327) <= not (a xor b);
    outputs(8328) <= not a;
    outputs(8329) <= a and not b;
    outputs(8330) <= a xor b;
    outputs(8331) <= not (a xor b);
    outputs(8332) <= not (a xor b);
    outputs(8333) <= not (a or b);
    outputs(8334) <= not (a or b);
    outputs(8335) <= a xor b;
    outputs(8336) <= not b or a;
    outputs(8337) <= not b;
    outputs(8338) <= not (a xor b);
    outputs(8339) <= not a;
    outputs(8340) <= a xor b;
    outputs(8341) <= a xor b;
    outputs(8342) <= a;
    outputs(8343) <= not (a or b);
    outputs(8344) <= a or b;
    outputs(8345) <= not b;
    outputs(8346) <= not (a and b);
    outputs(8347) <= a or b;
    outputs(8348) <= a and b;
    outputs(8349) <= not a;
    outputs(8350) <= a and not b;
    outputs(8351) <= not b;
    outputs(8352) <= not b or a;
    outputs(8353) <= b;
    outputs(8354) <= not b;
    outputs(8355) <= not (a or b);
    outputs(8356) <= not a;
    outputs(8357) <= not b;
    outputs(8358) <= not (a xor b);
    outputs(8359) <= not (a xor b);
    outputs(8360) <= not (a or b);
    outputs(8361) <= b;
    outputs(8362) <= not (a or b);
    outputs(8363) <= b;
    outputs(8364) <= not b;
    outputs(8365) <= b and not a;
    outputs(8366) <= a xor b;
    outputs(8367) <= 1'b1;
    outputs(8368) <= not (a xor b);
    outputs(8369) <= a and b;
    outputs(8370) <= not b;
    outputs(8371) <= not (a xor b);
    outputs(8372) <= not (a or b);
    outputs(8373) <= a and not b;
    outputs(8374) <= a;
    outputs(8375) <= not b;
    outputs(8376) <= not a;
    outputs(8377) <= b;
    outputs(8378) <= a and not b;
    outputs(8379) <= a;
    outputs(8380) <= a xor b;
    outputs(8381) <= not (a or b);
    outputs(8382) <= not (a or b);
    outputs(8383) <= a and b;
    outputs(8384) <= not b;
    outputs(8385) <= not (a xor b);
    outputs(8386) <= a xor b;
    outputs(8387) <= b;
    outputs(8388) <= not (a xor b);
    outputs(8389) <= a xor b;
    outputs(8390) <= not b;
    outputs(8391) <= not a;
    outputs(8392) <= not a;
    outputs(8393) <= b;
    outputs(8394) <= not (a xor b);
    outputs(8395) <= b;
    outputs(8396) <= a;
    outputs(8397) <= a;
    outputs(8398) <= not a;
    outputs(8399) <= b and not a;
    outputs(8400) <= b;
    outputs(8401) <= a;
    outputs(8402) <= a;
    outputs(8403) <= a xor b;
    outputs(8404) <= not (a and b);
    outputs(8405) <= not b;
    outputs(8406) <= a xor b;
    outputs(8407) <= not b;
    outputs(8408) <= not (a or b);
    outputs(8409) <= not b;
    outputs(8410) <= not a or b;
    outputs(8411) <= a;
    outputs(8412) <= a and not b;
    outputs(8413) <= not a or b;
    outputs(8414) <= not (a and b);
    outputs(8415) <= a xor b;
    outputs(8416) <= a;
    outputs(8417) <= a xor b;
    outputs(8418) <= not b;
    outputs(8419) <= b;
    outputs(8420) <= not (a or b);
    outputs(8421) <= not (a or b);
    outputs(8422) <= b;
    outputs(8423) <= b and not a;
    outputs(8424) <= b;
    outputs(8425) <= not a or b;
    outputs(8426) <= not (a xor b);
    outputs(8427) <= a xor b;
    outputs(8428) <= b;
    outputs(8429) <= a;
    outputs(8430) <= b;
    outputs(8431) <= a xor b;
    outputs(8432) <= b and not a;
    outputs(8433) <= not (a xor b);
    outputs(8434) <= not b;
    outputs(8435) <= a;
    outputs(8436) <= not b or a;
    outputs(8437) <= not b;
    outputs(8438) <= a;
    outputs(8439) <= not b or a;
    outputs(8440) <= a;
    outputs(8441) <= not b;
    outputs(8442) <= not b;
    outputs(8443) <= not b;
    outputs(8444) <= a;
    outputs(8445) <= not a;
    outputs(8446) <= not a;
    outputs(8447) <= not (a xor b);
    outputs(8448) <= a or b;
    outputs(8449) <= a xor b;
    outputs(8450) <= not b;
    outputs(8451) <= not (a xor b);
    outputs(8452) <= not b;
    outputs(8453) <= a xor b;
    outputs(8454) <= not b or a;
    outputs(8455) <= not (a xor b);
    outputs(8456) <= not (a xor b);
    outputs(8457) <= a and b;
    outputs(8458) <= b;
    outputs(8459) <= not (a or b);
    outputs(8460) <= a xor b;
    outputs(8461) <= not (a xor b);
    outputs(8462) <= a xor b;
    outputs(8463) <= not b;
    outputs(8464) <= not (a xor b);
    outputs(8465) <= not b;
    outputs(8466) <= a xor b;
    outputs(8467) <= a or b;
    outputs(8468) <= not (a xor b);
    outputs(8469) <= a and not b;
    outputs(8470) <= a and b;
    outputs(8471) <= a and not b;
    outputs(8472) <= b;
    outputs(8473) <= not a;
    outputs(8474) <= not (a xor b);
    outputs(8475) <= a and b;
    outputs(8476) <= a;
    outputs(8477) <= a and not b;
    outputs(8478) <= not (a or b);
    outputs(8479) <= not b;
    outputs(8480) <= not b or a;
    outputs(8481) <= b and not a;
    outputs(8482) <= not (a or b);
    outputs(8483) <= not a or b;
    outputs(8484) <= a xor b;
    outputs(8485) <= a and b;
    outputs(8486) <= a;
    outputs(8487) <= a;
    outputs(8488) <= a xor b;
    outputs(8489) <= not b;
    outputs(8490) <= not (a xor b);
    outputs(8491) <= not (a xor b);
    outputs(8492) <= not a;
    outputs(8493) <= a xor b;
    outputs(8494) <= not (a xor b);
    outputs(8495) <= a xor b;
    outputs(8496) <= a;
    outputs(8497) <= a and b;
    outputs(8498) <= not (a xor b);
    outputs(8499) <= a xor b;
    outputs(8500) <= b;
    outputs(8501) <= a xor b;
    outputs(8502) <= a;
    outputs(8503) <= not (a xor b);
    outputs(8504) <= not a;
    outputs(8505) <= not b;
    outputs(8506) <= not a or b;
    outputs(8507) <= not b or a;
    outputs(8508) <= a xor b;
    outputs(8509) <= not b;
    outputs(8510) <= not b;
    outputs(8511) <= not b or a;
    outputs(8512) <= a or b;
    outputs(8513) <= a;
    outputs(8514) <= not a;
    outputs(8515) <= a and not b;
    outputs(8516) <= not a or b;
    outputs(8517) <= b;
    outputs(8518) <= b;
    outputs(8519) <= a;
    outputs(8520) <= not a;
    outputs(8521) <= b and not a;
    outputs(8522) <= a;
    outputs(8523) <= b;
    outputs(8524) <= a xor b;
    outputs(8525) <= a;
    outputs(8526) <= not a;
    outputs(8527) <= a or b;
    outputs(8528) <= b;
    outputs(8529) <= not (a xor b);
    outputs(8530) <= b;
    outputs(8531) <= not (a or b);
    outputs(8532) <= not b;
    outputs(8533) <= not a;
    outputs(8534) <= a;
    outputs(8535) <= b and not a;
    outputs(8536) <= not (a xor b);
    outputs(8537) <= not b or a;
    outputs(8538) <= not (a xor b);
    outputs(8539) <= not (a xor b);
    outputs(8540) <= not b;
    outputs(8541) <= not a or b;
    outputs(8542) <= not a;
    outputs(8543) <= not b;
    outputs(8544) <= not a;
    outputs(8545) <= b and not a;
    outputs(8546) <= b and not a;
    outputs(8547) <= a xor b;
    outputs(8548) <= a xor b;
    outputs(8549) <= not (a xor b);
    outputs(8550) <= a and not b;
    outputs(8551) <= a;
    outputs(8552) <= a;
    outputs(8553) <= b;
    outputs(8554) <= not (a xor b);
    outputs(8555) <= not a;
    outputs(8556) <= a and b;
    outputs(8557) <= a xor b;
    outputs(8558) <= not (a xor b);
    outputs(8559) <= a;
    outputs(8560) <= a xor b;
    outputs(8561) <= b;
    outputs(8562) <= not b;
    outputs(8563) <= not b;
    outputs(8564) <= a;
    outputs(8565) <= a or b;
    outputs(8566) <= a xor b;
    outputs(8567) <= not a;
    outputs(8568) <= b;
    outputs(8569) <= not b or a;
    outputs(8570) <= a xor b;
    outputs(8571) <= not b;
    outputs(8572) <= a xor b;
    outputs(8573) <= a;
    outputs(8574) <= a xor b;
    outputs(8575) <= not (a or b);
    outputs(8576) <= not a or b;
    outputs(8577) <= a xor b;
    outputs(8578) <= a or b;
    outputs(8579) <= b;
    outputs(8580) <= not b;
    outputs(8581) <= a xor b;
    outputs(8582) <= b and not a;
    outputs(8583) <= not (a xor b);
    outputs(8584) <= not (a xor b);
    outputs(8585) <= a;
    outputs(8586) <= not (a xor b);
    outputs(8587) <= not (a xor b);
    outputs(8588) <= a;
    outputs(8589) <= a;
    outputs(8590) <= a;
    outputs(8591) <= a xor b;
    outputs(8592) <= a;
    outputs(8593) <= not (a xor b);
    outputs(8594) <= b and not a;
    outputs(8595) <= not a or b;
    outputs(8596) <= a and not b;
    outputs(8597) <= a and b;
    outputs(8598) <= not a;
    outputs(8599) <= a xor b;
    outputs(8600) <= not (a xor b);
    outputs(8601) <= not b;
    outputs(8602) <= not a;
    outputs(8603) <= not (a xor b);
    outputs(8604) <= a xor b;
    outputs(8605) <= a;
    outputs(8606) <= not b;
    outputs(8607) <= b;
    outputs(8608) <= not (a xor b);
    outputs(8609) <= not (a xor b);
    outputs(8610) <= not b;
    outputs(8611) <= b and not a;
    outputs(8612) <= not a;
    outputs(8613) <= a;
    outputs(8614) <= not a;
    outputs(8615) <= not (a or b);
    outputs(8616) <= a xor b;
    outputs(8617) <= a xor b;
    outputs(8618) <= not b;
    outputs(8619) <= not (a or b);
    outputs(8620) <= a xor b;
    outputs(8621) <= a and not b;
    outputs(8622) <= a and b;
    outputs(8623) <= not (a xor b);
    outputs(8624) <= not (a or b);
    outputs(8625) <= not (a xor b);
    outputs(8626) <= a xor b;
    outputs(8627) <= b;
    outputs(8628) <= a xor b;
    outputs(8629) <= b and not a;
    outputs(8630) <= b and not a;
    outputs(8631) <= a xor b;
    outputs(8632) <= not b;
    outputs(8633) <= not b;
    outputs(8634) <= a;
    outputs(8635) <= not (a xor b);
    outputs(8636) <= a xor b;
    outputs(8637) <= not (a and b);
    outputs(8638) <= not b;
    outputs(8639) <= a;
    outputs(8640) <= b;
    outputs(8641) <= b;
    outputs(8642) <= a xor b;
    outputs(8643) <= a;
    outputs(8644) <= a or b;
    outputs(8645) <= a xor b;
    outputs(8646) <= a xor b;
    outputs(8647) <= not b;
    outputs(8648) <= b;
    outputs(8649) <= a and b;
    outputs(8650) <= b and not a;
    outputs(8651) <= not a;
    outputs(8652) <= not a;
    outputs(8653) <= a xor b;
    outputs(8654) <= not (a xor b);
    outputs(8655) <= a and not b;
    outputs(8656) <= not (a xor b);
    outputs(8657) <= b and not a;
    outputs(8658) <= b and not a;
    outputs(8659) <= a or b;
    outputs(8660) <= not (a or b);
    outputs(8661) <= b;
    outputs(8662) <= a and not b;
    outputs(8663) <= not b;
    outputs(8664) <= b and not a;
    outputs(8665) <= not a;
    outputs(8666) <= a xor b;
    outputs(8667) <= b;
    outputs(8668) <= b;
    outputs(8669) <= not a;
    outputs(8670) <= a xor b;
    outputs(8671) <= b;
    outputs(8672) <= a and b;
    outputs(8673) <= a and b;
    outputs(8674) <= not (a xor b);
    outputs(8675) <= a and b;
    outputs(8676) <= b;
    outputs(8677) <= a;
    outputs(8678) <= b;
    outputs(8679) <= not b;
    outputs(8680) <= a xor b;
    outputs(8681) <= not b;
    outputs(8682) <= not (a xor b);
    outputs(8683) <= not a;
    outputs(8684) <= b;
    outputs(8685) <= a and not b;
    outputs(8686) <= not a;
    outputs(8687) <= a and b;
    outputs(8688) <= a;
    outputs(8689) <= b;
    outputs(8690) <= a and not b;
    outputs(8691) <= a xor b;
    outputs(8692) <= not a;
    outputs(8693) <= not a;
    outputs(8694) <= not (a xor b);
    outputs(8695) <= a and b;
    outputs(8696) <= b;
    outputs(8697) <= a and not b;
    outputs(8698) <= b and not a;
    outputs(8699) <= not (a xor b);
    outputs(8700) <= a xor b;
    outputs(8701) <= not a;
    outputs(8702) <= not (a xor b);
    outputs(8703) <= not a;
    outputs(8704) <= a xor b;
    outputs(8705) <= not (a and b);
    outputs(8706) <= a;
    outputs(8707) <= not (a or b);
    outputs(8708) <= a;
    outputs(8709) <= a;
    outputs(8710) <= not (a xor b);
    outputs(8711) <= b;
    outputs(8712) <= not a;
    outputs(8713) <= not b;
    outputs(8714) <= a;
    outputs(8715) <= not (a and b);
    outputs(8716) <= a and not b;
    outputs(8717) <= a and b;
    outputs(8718) <= not (a xor b);
    outputs(8719) <= a;
    outputs(8720) <= b;
    outputs(8721) <= a xor b;
    outputs(8722) <= b;
    outputs(8723) <= not b;
    outputs(8724) <= a;
    outputs(8725) <= b;
    outputs(8726) <= a xor b;
    outputs(8727) <= b;
    outputs(8728) <= a xor b;
    outputs(8729) <= not a;
    outputs(8730) <= a;
    outputs(8731) <= not b;
    outputs(8732) <= a and not b;
    outputs(8733) <= b;
    outputs(8734) <= a and not b;
    outputs(8735) <= a xor b;
    outputs(8736) <= b;
    outputs(8737) <= b;
    outputs(8738) <= a and not b;
    outputs(8739) <= a;
    outputs(8740) <= a and not b;
    outputs(8741) <= a xor b;
    outputs(8742) <= b and not a;
    outputs(8743) <= not (a xor b);
    outputs(8744) <= a xor b;
    outputs(8745) <= not b;
    outputs(8746) <= b and not a;
    outputs(8747) <= not a;
    outputs(8748) <= not (a xor b);
    outputs(8749) <= not a;
    outputs(8750) <= b;
    outputs(8751) <= a xor b;
    outputs(8752) <= a and not b;
    outputs(8753) <= b;
    outputs(8754) <= not a;
    outputs(8755) <= not b;
    outputs(8756) <= a and b;
    outputs(8757) <= not b;
    outputs(8758) <= not (a xor b);
    outputs(8759) <= not (a xor b);
    outputs(8760) <= not (a xor b);
    outputs(8761) <= a and b;
    outputs(8762) <= not (a xor b);
    outputs(8763) <= b and not a;
    outputs(8764) <= a xor b;
    outputs(8765) <= not b;
    outputs(8766) <= not b;
    outputs(8767) <= a;
    outputs(8768) <= a and not b;
    outputs(8769) <= not a;
    outputs(8770) <= not a;
    outputs(8771) <= a;
    outputs(8772) <= not b;
    outputs(8773) <= not b;
    outputs(8774) <= a;
    outputs(8775) <= not (a or b);
    outputs(8776) <= not (a xor b);
    outputs(8777) <= not b;
    outputs(8778) <= a and not b;
    outputs(8779) <= not (a or b);
    outputs(8780) <= not (a xor b);
    outputs(8781) <= a xor b;
    outputs(8782) <= b;
    outputs(8783) <= not (a xor b);
    outputs(8784) <= not a;
    outputs(8785) <= a or b;
    outputs(8786) <= b;
    outputs(8787) <= a xor b;
    outputs(8788) <= a;
    outputs(8789) <= not (a xor b);
    outputs(8790) <= b and not a;
    outputs(8791) <= not b or a;
    outputs(8792) <= b and not a;
    outputs(8793) <= a;
    outputs(8794) <= b and not a;
    outputs(8795) <= a;
    outputs(8796) <= a xor b;
    outputs(8797) <= a xor b;
    outputs(8798) <= a;
    outputs(8799) <= a xor b;
    outputs(8800) <= not (a or b);
    outputs(8801) <= b and not a;
    outputs(8802) <= a and not b;
    outputs(8803) <= b;
    outputs(8804) <= b;
    outputs(8805) <= b and not a;
    outputs(8806) <= a xor b;
    outputs(8807) <= b;
    outputs(8808) <= not a;
    outputs(8809) <= a and not b;
    outputs(8810) <= b and not a;
    outputs(8811) <= a and not b;
    outputs(8812) <= b;
    outputs(8813) <= a;
    outputs(8814) <= not b;
    outputs(8815) <= a;
    outputs(8816) <= a and not b;
    outputs(8817) <= not (a xor b);
    outputs(8818) <= a xor b;
    outputs(8819) <= not (a or b);
    outputs(8820) <= not (a xor b);
    outputs(8821) <= not a;
    outputs(8822) <= not a or b;
    outputs(8823) <= a and not b;
    outputs(8824) <= a;
    outputs(8825) <= a xor b;
    outputs(8826) <= a xor b;
    outputs(8827) <= not (a or b);
    outputs(8828) <= a xor b;
    outputs(8829) <= a and not b;
    outputs(8830) <= a;
    outputs(8831) <= not (a or b);
    outputs(8832) <= not (a xor b);
    outputs(8833) <= b;
    outputs(8834) <= not a;
    outputs(8835) <= a and b;
    outputs(8836) <= a xor b;
    outputs(8837) <= not (a xor b);
    outputs(8838) <= not (a xor b);
    outputs(8839) <= b;
    outputs(8840) <= not (a and b);
    outputs(8841) <= a;
    outputs(8842) <= a xor b;
    outputs(8843) <= a or b;
    outputs(8844) <= not (a xor b);
    outputs(8845) <= not a or b;
    outputs(8846) <= a xor b;
    outputs(8847) <= a xor b;
    outputs(8848) <= b and not a;
    outputs(8849) <= not b;
    outputs(8850) <= not b;
    outputs(8851) <= not (a and b);
    outputs(8852) <= a xor b;
    outputs(8853) <= not (a xor b);
    outputs(8854) <= a and b;
    outputs(8855) <= not (a or b);
    outputs(8856) <= not (a xor b);
    outputs(8857) <= not b or a;
    outputs(8858) <= not (a xor b);
    outputs(8859) <= not a;
    outputs(8860) <= a xor b;
    outputs(8861) <= a xor b;
    outputs(8862) <= not a;
    outputs(8863) <= a xor b;
    outputs(8864) <= not (a xor b);
    outputs(8865) <= a and not b;
    outputs(8866) <= a and b;
    outputs(8867) <= b;
    outputs(8868) <= not (a xor b);
    outputs(8869) <= a and not b;
    outputs(8870) <= not b;
    outputs(8871) <= not (a or b);
    outputs(8872) <= not (a xor b);
    outputs(8873) <= a and b;
    outputs(8874) <= a;
    outputs(8875) <= a and b;
    outputs(8876) <= not (a and b);
    outputs(8877) <= not b;
    outputs(8878) <= a and b;
    outputs(8879) <= not (a xor b);
    outputs(8880) <= not a or b;
    outputs(8881) <= not (a or b);
    outputs(8882) <= not b;
    outputs(8883) <= b;
    outputs(8884) <= a and b;
    outputs(8885) <= not a or b;
    outputs(8886) <= a xor b;
    outputs(8887) <= a and not b;
    outputs(8888) <= not b;
    outputs(8889) <= not a;
    outputs(8890) <= a and not b;
    outputs(8891) <= b and not a;
    outputs(8892) <= not (a or b);
    outputs(8893) <= not a;
    outputs(8894) <= not (a xor b);
    outputs(8895) <= b;
    outputs(8896) <= not a;
    outputs(8897) <= not b;
    outputs(8898) <= b;
    outputs(8899) <= not (a xor b);
    outputs(8900) <= b;
    outputs(8901) <= a xor b;
    outputs(8902) <= a and not b;
    outputs(8903) <= not (a xor b);
    outputs(8904) <= a;
    outputs(8905) <= a and not b;
    outputs(8906) <= a xor b;
    outputs(8907) <= b;
    outputs(8908) <= a;
    outputs(8909) <= a;
    outputs(8910) <= not (a xor b);
    outputs(8911) <= not (a xor b);
    outputs(8912) <= not a;
    outputs(8913) <= not (a xor b);
    outputs(8914) <= a;
    outputs(8915) <= not a or b;
    outputs(8916) <= not (a xor b);
    outputs(8917) <= not a;
    outputs(8918) <= not (a and b);
    outputs(8919) <= not a;
    outputs(8920) <= a and b;
    outputs(8921) <= a xor b;
    outputs(8922) <= not a;
    outputs(8923) <= not b;
    outputs(8924) <= not b;
    outputs(8925) <= not a;
    outputs(8926) <= a;
    outputs(8927) <= b;
    outputs(8928) <= b and not a;
    outputs(8929) <= not a or b;
    outputs(8930) <= not b;
    outputs(8931) <= a or b;
    outputs(8932) <= not (a xor b);
    outputs(8933) <= a xor b;
    outputs(8934) <= not a;
    outputs(8935) <= not b;
    outputs(8936) <= not (a xor b);
    outputs(8937) <= a xor b;
    outputs(8938) <= a and b;
    outputs(8939) <= not b;
    outputs(8940) <= a and b;
    outputs(8941) <= not b;
    outputs(8942) <= not (a and b);
    outputs(8943) <= not a;
    outputs(8944) <= not b;
    outputs(8945) <= a or b;
    outputs(8946) <= a;
    outputs(8947) <= not b;
    outputs(8948) <= b;
    outputs(8949) <= a xor b;
    outputs(8950) <= not (a xor b);
    outputs(8951) <= not (a xor b);
    outputs(8952) <= a and not b;
    outputs(8953) <= a xor b;
    outputs(8954) <= b and not a;
    outputs(8955) <= b;
    outputs(8956) <= not (a and b);
    outputs(8957) <= a;
    outputs(8958) <= a and b;
    outputs(8959) <= not (a xor b);
    outputs(8960) <= a and b;
    outputs(8961) <= not (a xor b);
    outputs(8962) <= not (a xor b);
    outputs(8963) <= a xor b;
    outputs(8964) <= not b;
    outputs(8965) <= not b;
    outputs(8966) <= not a;
    outputs(8967) <= b and not a;
    outputs(8968) <= not a;
    outputs(8969) <= not b;
    outputs(8970) <= b and not a;
    outputs(8971) <= not b;
    outputs(8972) <= b and not a;
    outputs(8973) <= not b;
    outputs(8974) <= a;
    outputs(8975) <= a xor b;
    outputs(8976) <= a xor b;
    outputs(8977) <= not a;
    outputs(8978) <= b;
    outputs(8979) <= a xor b;
    outputs(8980) <= not a;
    outputs(8981) <= a and not b;
    outputs(8982) <= a;
    outputs(8983) <= not (a xor b);
    outputs(8984) <= a and b;
    outputs(8985) <= not (a or b);
    outputs(8986) <= not a;
    outputs(8987) <= not (a or b);
    outputs(8988) <= not (a xor b);
    outputs(8989) <= not (a or b);
    outputs(8990) <= b;
    outputs(8991) <= a xor b;
    outputs(8992) <= not a;
    outputs(8993) <= a or b;
    outputs(8994) <= not b;
    outputs(8995) <= b and not a;
    outputs(8996) <= not a;
    outputs(8997) <= a;
    outputs(8998) <= a xor b;
    outputs(8999) <= a;
    outputs(9000) <= b and not a;
    outputs(9001) <= not b;
    outputs(9002) <= not b;
    outputs(9003) <= not b;
    outputs(9004) <= a xor b;
    outputs(9005) <= a and b;
    outputs(9006) <= a;
    outputs(9007) <= not b;
    outputs(9008) <= not a;
    outputs(9009) <= a or b;
    outputs(9010) <= b and not a;
    outputs(9011) <= a xor b;
    outputs(9012) <= a and not b;
    outputs(9013) <= not a or b;
    outputs(9014) <= not (a xor b);
    outputs(9015) <= a and not b;
    outputs(9016) <= not (a xor b);
    outputs(9017) <= not (a and b);
    outputs(9018) <= a and b;
    outputs(9019) <= a and not b;
    outputs(9020) <= not b or a;
    outputs(9021) <= not (a and b);
    outputs(9022) <= a xor b;
    outputs(9023) <= not (a or b);
    outputs(9024) <= b and not a;
    outputs(9025) <= not b or a;
    outputs(9026) <= not (a xor b);
    outputs(9027) <= a xor b;
    outputs(9028) <= not (a and b);
    outputs(9029) <= b;
    outputs(9030) <= b and not a;
    outputs(9031) <= b;
    outputs(9032) <= b;
    outputs(9033) <= a;
    outputs(9034) <= b;
    outputs(9035) <= a and not b;
    outputs(9036) <= b;
    outputs(9037) <= not b;
    outputs(9038) <= not (a xor b);
    outputs(9039) <= a or b;
    outputs(9040) <= b and not a;
    outputs(9041) <= not (a or b);
    outputs(9042) <= a and b;
    outputs(9043) <= not a;
    outputs(9044) <= a;
    outputs(9045) <= a;
    outputs(9046) <= not a or b;
    outputs(9047) <= not a;
    outputs(9048) <= not (a xor b);
    outputs(9049) <= not (a xor b);
    outputs(9050) <= not b or a;
    outputs(9051) <= not a;
    outputs(9052) <= not a;
    outputs(9053) <= a xor b;
    outputs(9054) <= not (a xor b);
    outputs(9055) <= not (a xor b);
    outputs(9056) <= not (a or b);
    outputs(9057) <= not (a or b);
    outputs(9058) <= b and not a;
    outputs(9059) <= b;
    outputs(9060) <= not a;
    outputs(9061) <= a;
    outputs(9062) <= a xor b;
    outputs(9063) <= b;
    outputs(9064) <= b and not a;
    outputs(9065) <= not a;
    outputs(9066) <= b;
    outputs(9067) <= b and not a;
    outputs(9068) <= not (a or b);
    outputs(9069) <= a;
    outputs(9070) <= a xor b;
    outputs(9071) <= a and b;
    outputs(9072) <= not a;
    outputs(9073) <= a and b;
    outputs(9074) <= b;
    outputs(9075) <= a xor b;
    outputs(9076) <= not (a xor b);
    outputs(9077) <= a xor b;
    outputs(9078) <= b and not a;
    outputs(9079) <= not b;
    outputs(9080) <= a xor b;
    outputs(9081) <= a and not b;
    outputs(9082) <= b;
    outputs(9083) <= not (a xor b);
    outputs(9084) <= a xor b;
    outputs(9085) <= not (a or b);
    outputs(9086) <= b;
    outputs(9087) <= b;
    outputs(9088) <= b and not a;
    outputs(9089) <= a;
    outputs(9090) <= a xor b;
    outputs(9091) <= not (a or b);
    outputs(9092) <= not a;
    outputs(9093) <= a and b;
    outputs(9094) <= a;
    outputs(9095) <= not (a or b);
    outputs(9096) <= a xor b;
    outputs(9097) <= a xor b;
    outputs(9098) <= not a;
    outputs(9099) <= a and not b;
    outputs(9100) <= b;
    outputs(9101) <= a and not b;
    outputs(9102) <= a xor b;
    outputs(9103) <= b;
    outputs(9104) <= a xor b;
    outputs(9105) <= not (a or b);
    outputs(9106) <= not (a xor b);
    outputs(9107) <= a xor b;
    outputs(9108) <= a and b;
    outputs(9109) <= not a;
    outputs(9110) <= not (a xor b);
    outputs(9111) <= a xor b;
    outputs(9112) <= b;
    outputs(9113) <= not (a xor b);
    outputs(9114) <= a;
    outputs(9115) <= not b;
    outputs(9116) <= not b or a;
    outputs(9117) <= a;
    outputs(9118) <= a;
    outputs(9119) <= not b or a;
    outputs(9120) <= not (a xor b);
    outputs(9121) <= not a;
    outputs(9122) <= b;
    outputs(9123) <= a xor b;
    outputs(9124) <= a;
    outputs(9125) <= b;
    outputs(9126) <= a xor b;
    outputs(9127) <= b;
    outputs(9128) <= not (a xor b);
    outputs(9129) <= b and not a;
    outputs(9130) <= not a;
    outputs(9131) <= not (a xor b);
    outputs(9132) <= not (a xor b);
    outputs(9133) <= not b;
    outputs(9134) <= a xor b;
    outputs(9135) <= not b;
    outputs(9136) <= not (a xor b);
    outputs(9137) <= a xor b;
    outputs(9138) <= b;
    outputs(9139) <= not (a xor b);
    outputs(9140) <= not (a xor b);
    outputs(9141) <= not a;
    outputs(9142) <= not a;
    outputs(9143) <= not a;
    outputs(9144) <= a xor b;
    outputs(9145) <= a;
    outputs(9146) <= not a;
    outputs(9147) <= not a;
    outputs(9148) <= not a;
    outputs(9149) <= not a or b;
    outputs(9150) <= not b;
    outputs(9151) <= a;
    outputs(9152) <= not (a or b);
    outputs(9153) <= a xor b;
    outputs(9154) <= a and b;
    outputs(9155) <= a and b;
    outputs(9156) <= a and not b;
    outputs(9157) <= 1'b0;
    outputs(9158) <= not (a xor b);
    outputs(9159) <= not b;
    outputs(9160) <= b;
    outputs(9161) <= b and not a;
    outputs(9162) <= b;
    outputs(9163) <= not a;
    outputs(9164) <= not (a and b);
    outputs(9165) <= not (a xor b);
    outputs(9166) <= not b;
    outputs(9167) <= not (a xor b);
    outputs(9168) <= not b;
    outputs(9169) <= not (a xor b);
    outputs(9170) <= not b;
    outputs(9171) <= a;
    outputs(9172) <= b;
    outputs(9173) <= b;
    outputs(9174) <= not (a xor b);
    outputs(9175) <= not a or b;
    outputs(9176) <= a xor b;
    outputs(9177) <= a xor b;
    outputs(9178) <= b;
    outputs(9179) <= b and not a;
    outputs(9180) <= a xor b;
    outputs(9181) <= a xor b;
    outputs(9182) <= not (a or b);
    outputs(9183) <= not a or b;
    outputs(9184) <= a xor b;
    outputs(9185) <= a and not b;
    outputs(9186) <= not a or b;
    outputs(9187) <= not b;
    outputs(9188) <= not (a xor b);
    outputs(9189) <= not b;
    outputs(9190) <= a xor b;
    outputs(9191) <= a;
    outputs(9192) <= a xor b;
    outputs(9193) <= not (a or b);
    outputs(9194) <= not (a or b);
    outputs(9195) <= not b;
    outputs(9196) <= a and b;
    outputs(9197) <= not (a xor b);
    outputs(9198) <= b and not a;
    outputs(9199) <= a xor b;
    outputs(9200) <= not (a or b);
    outputs(9201) <= a;
    outputs(9202) <= b;
    outputs(9203) <= not (a or b);
    outputs(9204) <= not a;
    outputs(9205) <= a or b;
    outputs(9206) <= not b;
    outputs(9207) <= not a;
    outputs(9208) <= a;
    outputs(9209) <= b;
    outputs(9210) <= not b;
    outputs(9211) <= b and not a;
    outputs(9212) <= not a;
    outputs(9213) <= a xor b;
    outputs(9214) <= a and b;
    outputs(9215) <= not (a xor b);
    outputs(9216) <= not (a or b);
    outputs(9217) <= b and not a;
    outputs(9218) <= not b or a;
    outputs(9219) <= a;
    outputs(9220) <= not (a or b);
    outputs(9221) <= not a;
    outputs(9222) <= not b;
    outputs(9223) <= b and not a;
    outputs(9224) <= a xor b;
    outputs(9225) <= not a;
    outputs(9226) <= not (a and b);
    outputs(9227) <= not (a and b);
    outputs(9228) <= not b;
    outputs(9229) <= b and not a;
    outputs(9230) <= a and b;
    outputs(9231) <= not a or b;
    outputs(9232) <= not (a and b);
    outputs(9233) <= not (a xor b);
    outputs(9234) <= a xor b;
    outputs(9235) <= a and b;
    outputs(9236) <= a and not b;
    outputs(9237) <= b;
    outputs(9238) <= b and not a;
    outputs(9239) <= not (a and b);
    outputs(9240) <= a xor b;
    outputs(9241) <= not a;
    outputs(9242) <= a and not b;
    outputs(9243) <= a and b;
    outputs(9244) <= a and b;
    outputs(9245) <= b;
    outputs(9246) <= not a;
    outputs(9247) <= not (a xor b);
    outputs(9248) <= a;
    outputs(9249) <= a xor b;
    outputs(9250) <= not (a xor b);
    outputs(9251) <= a xor b;
    outputs(9252) <= not a;
    outputs(9253) <= a xor b;
    outputs(9254) <= b and not a;
    outputs(9255) <= a xor b;
    outputs(9256) <= a and not b;
    outputs(9257) <= a xor b;
    outputs(9258) <= b and not a;
    outputs(9259) <= a and b;
    outputs(9260) <= a and b;
    outputs(9261) <= a;
    outputs(9262) <= b;
    outputs(9263) <= not (a xor b);
    outputs(9264) <= not (a xor b);
    outputs(9265) <= a;
    outputs(9266) <= b;
    outputs(9267) <= a and not b;
    outputs(9268) <= a or b;
    outputs(9269) <= a;
    outputs(9270) <= a and b;
    outputs(9271) <= b;
    outputs(9272) <= not a;
    outputs(9273) <= not (a and b);
    outputs(9274) <= a and not b;
    outputs(9275) <= not b;
    outputs(9276) <= not a;
    outputs(9277) <= a;
    outputs(9278) <= b and not a;
    outputs(9279) <= not a;
    outputs(9280) <= not b;
    outputs(9281) <= a and b;
    outputs(9282) <= a or b;
    outputs(9283) <= not a;
    outputs(9284) <= not (a xor b);
    outputs(9285) <= b and not a;
    outputs(9286) <= a xor b;
    outputs(9287) <= a xor b;
    outputs(9288) <= a and not b;
    outputs(9289) <= a or b;
    outputs(9290) <= not b or a;
    outputs(9291) <= not a;
    outputs(9292) <= a xor b;
    outputs(9293) <= a xor b;
    outputs(9294) <= a or b;
    outputs(9295) <= not (a xor b);
    outputs(9296) <= a;
    outputs(9297) <= not a or b;
    outputs(9298) <= not a;
    outputs(9299) <= not b;
    outputs(9300) <= not (a xor b);
    outputs(9301) <= not a;
    outputs(9302) <= a xor b;
    outputs(9303) <= not (a xor b);
    outputs(9304) <= not (a xor b);
    outputs(9305) <= a and b;
    outputs(9306) <= not (a xor b);
    outputs(9307) <= b;
    outputs(9308) <= a xor b;
    outputs(9309) <= a;
    outputs(9310) <= a and b;
    outputs(9311) <= not a;
    outputs(9312) <= not b;
    outputs(9313) <= not b;
    outputs(9314) <= a;
    outputs(9315) <= a;
    outputs(9316) <= not a;
    outputs(9317) <= not (a xor b);
    outputs(9318) <= not a;
    outputs(9319) <= a or b;
    outputs(9320) <= a and b;
    outputs(9321) <= a and b;
    outputs(9322) <= a xor b;
    outputs(9323) <= a or b;
    outputs(9324) <= not b;
    outputs(9325) <= a xor b;
    outputs(9326) <= a and b;
    outputs(9327) <= b;
    outputs(9328) <= not (a or b);
    outputs(9329) <= b;
    outputs(9330) <= a;
    outputs(9331) <= not (a or b);
    outputs(9332) <= not (a xor b);
    outputs(9333) <= not b;
    outputs(9334) <= a and not b;
    outputs(9335) <= a and not b;
    outputs(9336) <= not (a xor b);
    outputs(9337) <= not a;
    outputs(9338) <= a xor b;
    outputs(9339) <= not a;
    outputs(9340) <= a xor b;
    outputs(9341) <= a xor b;
    outputs(9342) <= a xor b;
    outputs(9343) <= not (a xor b);
    outputs(9344) <= a and b;
    outputs(9345) <= a;
    outputs(9346) <= a;
    outputs(9347) <= not b;
    outputs(9348) <= a;
    outputs(9349) <= a xor b;
    outputs(9350) <= not (a and b);
    outputs(9351) <= b;
    outputs(9352) <= not (a xor b);
    outputs(9353) <= not a;
    outputs(9354) <= not b;
    outputs(9355) <= not b;
    outputs(9356) <= a xor b;
    outputs(9357) <= a and b;
    outputs(9358) <= a;
    outputs(9359) <= not (a or b);
    outputs(9360) <= a xor b;
    outputs(9361) <= a and b;
    outputs(9362) <= a and b;
    outputs(9363) <= not (a xor b);
    outputs(9364) <= a xor b;
    outputs(9365) <= a and not b;
    outputs(9366) <= a;
    outputs(9367) <= not (a and b);
    outputs(9368) <= not (a xor b);
    outputs(9369) <= not b;
    outputs(9370) <= a;
    outputs(9371) <= not b;
    outputs(9372) <= not b;
    outputs(9373) <= b and not a;
    outputs(9374) <= not (a and b);
    outputs(9375) <= b;
    outputs(9376) <= not b;
    outputs(9377) <= not (a or b);
    outputs(9378) <= not a or b;
    outputs(9379) <= not b or a;
    outputs(9380) <= b;
    outputs(9381) <= not a;
    outputs(9382) <= a and not b;
    outputs(9383) <= b and not a;
    outputs(9384) <= not a;
    outputs(9385) <= b;
    outputs(9386) <= not (a or b);
    outputs(9387) <= a xor b;
    outputs(9388) <= not a;
    outputs(9389) <= not (a xor b);
    outputs(9390) <= b and not a;
    outputs(9391) <= a xor b;
    outputs(9392) <= a and not b;
    outputs(9393) <= a;
    outputs(9394) <= not a;
    outputs(9395) <= b;
    outputs(9396) <= a or b;
    outputs(9397) <= not (a xor b);
    outputs(9398) <= not (a and b);
    outputs(9399) <= b and not a;
    outputs(9400) <= a and b;
    outputs(9401) <= a xor b;
    outputs(9402) <= b;
    outputs(9403) <= not (a xor b);
    outputs(9404) <= not b or a;
    outputs(9405) <= not (a and b);
    outputs(9406) <= not (a xor b);
    outputs(9407) <= a;
    outputs(9408) <= not (a or b);
    outputs(9409) <= a xor b;
    outputs(9410) <= not (a xor b);
    outputs(9411) <= not b;
    outputs(9412) <= not (a xor b);
    outputs(9413) <= a;
    outputs(9414) <= not (a or b);
    outputs(9415) <= b;
    outputs(9416) <= b and not a;
    outputs(9417) <= not (a or b);
    outputs(9418) <= not b;
    outputs(9419) <= b;
    outputs(9420) <= not (a or b);
    outputs(9421) <= not b;
    outputs(9422) <= not (a xor b);
    outputs(9423) <= not (a or b);
    outputs(9424) <= a;
    outputs(9425) <= a xor b;
    outputs(9426) <= not (a or b);
    outputs(9427) <= not (a xor b);
    outputs(9428) <= not a;
    outputs(9429) <= not (a or b);
    outputs(9430) <= not (a and b);
    outputs(9431) <= a and b;
    outputs(9432) <= a xor b;
    outputs(9433) <= a and b;
    outputs(9434) <= not (a or b);
    outputs(9435) <= a or b;
    outputs(9436) <= b;
    outputs(9437) <= not a;
    outputs(9438) <= not a;
    outputs(9439) <= not b;
    outputs(9440) <= b and not a;
    outputs(9441) <= b;
    outputs(9442) <= a and not b;
    outputs(9443) <= b and not a;
    outputs(9444) <= a xor b;
    outputs(9445) <= not (a xor b);
    outputs(9446) <= not (a xor b);
    outputs(9447) <= not a;
    outputs(9448) <= not b;
    outputs(9449) <= a and not b;
    outputs(9450) <= b and not a;
    outputs(9451) <= b and not a;
    outputs(9452) <= not (a xor b);
    outputs(9453) <= not a;
    outputs(9454) <= a xor b;
    outputs(9455) <= b;
    outputs(9456) <= not a;
    outputs(9457) <= b;
    outputs(9458) <= b;
    outputs(9459) <= not b;
    outputs(9460) <= a;
    outputs(9461) <= not a;
    outputs(9462) <= a and not b;
    outputs(9463) <= a;
    outputs(9464) <= b and not a;
    outputs(9465) <= b;
    outputs(9466) <= a xor b;
    outputs(9467) <= not b;
    outputs(9468) <= b;
    outputs(9469) <= a xor b;
    outputs(9470) <= b;
    outputs(9471) <= not (a xor b);
    outputs(9472) <= not b;
    outputs(9473) <= not (a and b);
    outputs(9474) <= not a or b;
    outputs(9475) <= not (a and b);
    outputs(9476) <= not a;
    outputs(9477) <= not (a and b);
    outputs(9478) <= not (a xor b);
    outputs(9479) <= not (a xor b);
    outputs(9480) <= b;
    outputs(9481) <= not b;
    outputs(9482) <= not a;
    outputs(9483) <= not (a or b);
    outputs(9484) <= b;
    outputs(9485) <= a xor b;
    outputs(9486) <= a;
    outputs(9487) <= not a;
    outputs(9488) <= 1'b0;
    outputs(9489) <= a xor b;
    outputs(9490) <= not (a or b);
    outputs(9491) <= not b;
    outputs(9492) <= a;
    outputs(9493) <= b;
    outputs(9494) <= not (a xor b);
    outputs(9495) <= not a or b;
    outputs(9496) <= a and b;
    outputs(9497) <= b and not a;
    outputs(9498) <= not (a and b);
    outputs(9499) <= a and b;
    outputs(9500) <= a xor b;
    outputs(9501) <= not (a xor b);
    outputs(9502) <= a or b;
    outputs(9503) <= not b or a;
    outputs(9504) <= b and not a;
    outputs(9505) <= a;
    outputs(9506) <= not a;
    outputs(9507) <= a xor b;
    outputs(9508) <= not a;
    outputs(9509) <= a and not b;
    outputs(9510) <= not (a xor b);
    outputs(9511) <= not (a xor b);
    outputs(9512) <= not (a or b);
    outputs(9513) <= a xor b;
    outputs(9514) <= not (a or b);
    outputs(9515) <= a;
    outputs(9516) <= not a or b;
    outputs(9517) <= a xor b;
    outputs(9518) <= a xor b;
    outputs(9519) <= a;
    outputs(9520) <= not b;
    outputs(9521) <= not (a and b);
    outputs(9522) <= not b;
    outputs(9523) <= a;
    outputs(9524) <= a xor b;
    outputs(9525) <= a;
    outputs(9526) <= a and b;
    outputs(9527) <= a xor b;
    outputs(9528) <= not a;
    outputs(9529) <= not (a xor b);
    outputs(9530) <= a and not b;
    outputs(9531) <= not (a xor b);
    outputs(9532) <= not (a xor b);
    outputs(9533) <= not a;
    outputs(9534) <= not a;
    outputs(9535) <= b and not a;
    outputs(9536) <= not (a or b);
    outputs(9537) <= b;
    outputs(9538) <= not (a xor b);
    outputs(9539) <= not b;
    outputs(9540) <= a and not b;
    outputs(9541) <= not a;
    outputs(9542) <= not (a xor b);
    outputs(9543) <= not (a xor b);
    outputs(9544) <= a and not b;
    outputs(9545) <= a xor b;
    outputs(9546) <= a;
    outputs(9547) <= not b;
    outputs(9548) <= a;
    outputs(9549) <= a and b;
    outputs(9550) <= not b or a;
    outputs(9551) <= not a;
    outputs(9552) <= a xor b;
    outputs(9553) <= not (a xor b);
    outputs(9554) <= a and b;
    outputs(9555) <= a and b;
    outputs(9556) <= a;
    outputs(9557) <= a xor b;
    outputs(9558) <= not (a xor b);
    outputs(9559) <= b;
    outputs(9560) <= not (a xor b);
    outputs(9561) <= a and b;
    outputs(9562) <= b;
    outputs(9563) <= a;
    outputs(9564) <= not b;
    outputs(9565) <= a xor b;
    outputs(9566) <= a;
    outputs(9567) <= a or b;
    outputs(9568) <= b;
    outputs(9569) <= not a;
    outputs(9570) <= b and not a;
    outputs(9571) <= a and b;
    outputs(9572) <= not a;
    outputs(9573) <= not b or a;
    outputs(9574) <= a;
    outputs(9575) <= not b or a;
    outputs(9576) <= a and not b;
    outputs(9577) <= b;
    outputs(9578) <= a and not b;
    outputs(9579) <= b;
    outputs(9580) <= b;
    outputs(9581) <= not b;
    outputs(9582) <= a or b;
    outputs(9583) <= not b;
    outputs(9584) <= a;
    outputs(9585) <= a xor b;
    outputs(9586) <= b;
    outputs(9587) <= a xor b;
    outputs(9588) <= a and not b;
    outputs(9589) <= not (a xor b);
    outputs(9590) <= b;
    outputs(9591) <= not a;
    outputs(9592) <= a xor b;
    outputs(9593) <= not b;
    outputs(9594) <= not (a xor b);
    outputs(9595) <= not (a or b);
    outputs(9596) <= not (a xor b);
    outputs(9597) <= not a or b;
    outputs(9598) <= not (a and b);
    outputs(9599) <= not (a and b);
    outputs(9600) <= not a;
    outputs(9601) <= a xor b;
    outputs(9602) <= not (a or b);
    outputs(9603) <= a xor b;
    outputs(9604) <= not (a xor b);
    outputs(9605) <= not b;
    outputs(9606) <= b;
    outputs(9607) <= not a;
    outputs(9608) <= a;
    outputs(9609) <= not b;
    outputs(9610) <= not (a xor b);
    outputs(9611) <= not b;
    outputs(9612) <= not b;
    outputs(9613) <= a;
    outputs(9614) <= not (a or b);
    outputs(9615) <= b and not a;
    outputs(9616) <= not b;
    outputs(9617) <= not (a xor b);
    outputs(9618) <= a xor b;
    outputs(9619) <= a;
    outputs(9620) <= not (a xor b);
    outputs(9621) <= a and b;
    outputs(9622) <= a xor b;
    outputs(9623) <= a xor b;
    outputs(9624) <= b;
    outputs(9625) <= a and not b;
    outputs(9626) <= a or b;
    outputs(9627) <= a xor b;
    outputs(9628) <= a and not b;
    outputs(9629) <= b;
    outputs(9630) <= a xor b;
    outputs(9631) <= not b;
    outputs(9632) <= a xor b;
    outputs(9633) <= not (a or b);
    outputs(9634) <= b;
    outputs(9635) <= a or b;
    outputs(9636) <= not (a xor b);
    outputs(9637) <= not (a or b);
    outputs(9638) <= b;
    outputs(9639) <= b;
    outputs(9640) <= a xor b;
    outputs(9641) <= a xor b;
    outputs(9642) <= not b;
    outputs(9643) <= b;
    outputs(9644) <= not (a xor b);
    outputs(9645) <= a;
    outputs(9646) <= not b;
    outputs(9647) <= not b;
    outputs(9648) <= a xor b;
    outputs(9649) <= b and not a;
    outputs(9650) <= not a;
    outputs(9651) <= b;
    outputs(9652) <= a xor b;
    outputs(9653) <= not (a or b);
    outputs(9654) <= not b;
    outputs(9655) <= b and not a;
    outputs(9656) <= not (a xor b);
    outputs(9657) <= not b;
    outputs(9658) <= a and not b;
    outputs(9659) <= not b;
    outputs(9660) <= not (a or b);
    outputs(9661) <= a or b;
    outputs(9662) <= not (a xor b);
    outputs(9663) <= not a;
    outputs(9664) <= b;
    outputs(9665) <= a;
    outputs(9666) <= not a or b;
    outputs(9667) <= a xor b;
    outputs(9668) <= b;
    outputs(9669) <= a;
    outputs(9670) <= not (a xor b);
    outputs(9671) <= a;
    outputs(9672) <= a and b;
    outputs(9673) <= a xor b;
    outputs(9674) <= b;
    outputs(9675) <= not a;
    outputs(9676) <= not b or a;
    outputs(9677) <= b;
    outputs(9678) <= not b;
    outputs(9679) <= not a;
    outputs(9680) <= not a;
    outputs(9681) <= not (a xor b);
    outputs(9682) <= not (a or b);
    outputs(9683) <= a;
    outputs(9684) <= not (a xor b);
    outputs(9685) <= not b or a;
    outputs(9686) <= not (a xor b);
    outputs(9687) <= a;
    outputs(9688) <= not (a xor b);
    outputs(9689) <= a or b;
    outputs(9690) <= not a;
    outputs(9691) <= not a;
    outputs(9692) <= a and not b;
    outputs(9693) <= not (a xor b);
    outputs(9694) <= not (a or b);
    outputs(9695) <= a;
    outputs(9696) <= a and b;
    outputs(9697) <= 1'b0;
    outputs(9698) <= a xor b;
    outputs(9699) <= b;
    outputs(9700) <= not (a xor b);
    outputs(9701) <= a;
    outputs(9702) <= not a;
    outputs(9703) <= a and b;
    outputs(9704) <= a;
    outputs(9705) <= a;
    outputs(9706) <= b and not a;
    outputs(9707) <= not (a or b);
    outputs(9708) <= not (a or b);
    outputs(9709) <= not a;
    outputs(9710) <= not b;
    outputs(9711) <= a and not b;
    outputs(9712) <= not a;
    outputs(9713) <= not (a and b);
    outputs(9714) <= not b;
    outputs(9715) <= a;
    outputs(9716) <= a and b;
    outputs(9717) <= a xor b;
    outputs(9718) <= a and b;
    outputs(9719) <= not b;
    outputs(9720) <= a and not b;
    outputs(9721) <= not a;
    outputs(9722) <= a;
    outputs(9723) <= not (a xor b);
    outputs(9724) <= b;
    outputs(9725) <= not (a xor b);
    outputs(9726) <= not (a xor b);
    outputs(9727) <= a xor b;
    outputs(9728) <= a and not b;
    outputs(9729) <= a xor b;
    outputs(9730) <= not (a or b);
    outputs(9731) <= not (a and b);
    outputs(9732) <= not (a xor b);
    outputs(9733) <= a xor b;
    outputs(9734) <= not b or a;
    outputs(9735) <= not (a xor b);
    outputs(9736) <= a xor b;
    outputs(9737) <= a xor b;
    outputs(9738) <= not a;
    outputs(9739) <= not b;
    outputs(9740) <= not b;
    outputs(9741) <= a;
    outputs(9742) <= a xor b;
    outputs(9743) <= a xor b;
    outputs(9744) <= a xor b;
    outputs(9745) <= not a;
    outputs(9746) <= a and not b;
    outputs(9747) <= b;
    outputs(9748) <= a and b;
    outputs(9749) <= a xor b;
    outputs(9750) <= a or b;
    outputs(9751) <= b;
    outputs(9752) <= a xor b;
    outputs(9753) <= not b;
    outputs(9754) <= not (a or b);
    outputs(9755) <= a and not b;
    outputs(9756) <= not b;
    outputs(9757) <= a xor b;
    outputs(9758) <= not b;
    outputs(9759) <= not b;
    outputs(9760) <= a and not b;
    outputs(9761) <= not (a or b);
    outputs(9762) <= not b;
    outputs(9763) <= not (a xor b);
    outputs(9764) <= b and not a;
    outputs(9765) <= not (a or b);
    outputs(9766) <= not (a xor b);
    outputs(9767) <= a xor b;
    outputs(9768) <= a and b;
    outputs(9769) <= b;
    outputs(9770) <= a xor b;
    outputs(9771) <= not (a xor b);
    outputs(9772) <= not (a xor b);
    outputs(9773) <= a xor b;
    outputs(9774) <= a xor b;
    outputs(9775) <= a and b;
    outputs(9776) <= not (a xor b);
    outputs(9777) <= not a or b;
    outputs(9778) <= a;
    outputs(9779) <= not (a xor b);
    outputs(9780) <= not b;
    outputs(9781) <= a xor b;
    outputs(9782) <= not (a xor b);
    outputs(9783) <= not (a xor b);
    outputs(9784) <= b;
    outputs(9785) <= not b;
    outputs(9786) <= not (a xor b);
    outputs(9787) <= a xor b;
    outputs(9788) <= not (a xor b);
    outputs(9789) <= b;
    outputs(9790) <= b;
    outputs(9791) <= not a;
    outputs(9792) <= not (a xor b);
    outputs(9793) <= a;
    outputs(9794) <= a or b;
    outputs(9795) <= not b;
    outputs(9796) <= a xor b;
    outputs(9797) <= a xor b;
    outputs(9798) <= not (a xor b);
    outputs(9799) <= not (a xor b);
    outputs(9800) <= a;
    outputs(9801) <= a and not b;
    outputs(9802) <= b and not a;
    outputs(9803) <= not a;
    outputs(9804) <= not a;
    outputs(9805) <= a xor b;
    outputs(9806) <= a and b;
    outputs(9807) <= not (a xor b);
    outputs(9808) <= not a;
    outputs(9809) <= not (a or b);
    outputs(9810) <= a;
    outputs(9811) <= not b;
    outputs(9812) <= a;
    outputs(9813) <= a xor b;
    outputs(9814) <= a and b;
    outputs(9815) <= not a;
    outputs(9816) <= b;
    outputs(9817) <= a and b;
    outputs(9818) <= b;
    outputs(9819) <= not (a xor b);
    outputs(9820) <= not b;
    outputs(9821) <= not (a and b);
    outputs(9822) <= a;
    outputs(9823) <= b and not a;
    outputs(9824) <= not (a xor b);
    outputs(9825) <= b;
    outputs(9826) <= not (a xor b);
    outputs(9827) <= not (a xor b);
    outputs(9828) <= not (a xor b);
    outputs(9829) <= not b;
    outputs(9830) <= a;
    outputs(9831) <= b and not a;
    outputs(9832) <= b;
    outputs(9833) <= b and not a;
    outputs(9834) <= not (a or b);
    outputs(9835) <= b and not a;
    outputs(9836) <= a xor b;
    outputs(9837) <= not (a or b);
    outputs(9838) <= b and not a;
    outputs(9839) <= a and b;
    outputs(9840) <= b;
    outputs(9841) <= b;
    outputs(9842) <= not (a and b);
    outputs(9843) <= not (a or b);
    outputs(9844) <= a xor b;
    outputs(9845) <= b;
    outputs(9846) <= not b;
    outputs(9847) <= a;
    outputs(9848) <= not a or b;
    outputs(9849) <= a and not b;
    outputs(9850) <= not a or b;
    outputs(9851) <= a and not b;
    outputs(9852) <= b;
    outputs(9853) <= a and not b;
    outputs(9854) <= a xor b;
    outputs(9855) <= a and not b;
    outputs(9856) <= not (a or b);
    outputs(9857) <= not b;
    outputs(9858) <= a xor b;
    outputs(9859) <= not (a xor b);
    outputs(9860) <= not b or a;
    outputs(9861) <= b;
    outputs(9862) <= not (a xor b);
    outputs(9863) <= not (a and b);
    outputs(9864) <= not (a or b);
    outputs(9865) <= not (a xor b);
    outputs(9866) <= a xor b;
    outputs(9867) <= not b;
    outputs(9868) <= not b;
    outputs(9869) <= not a;
    outputs(9870) <= not a;
    outputs(9871) <= not a;
    outputs(9872) <= b and not a;
    outputs(9873) <= b;
    outputs(9874) <= a xor b;
    outputs(9875) <= not (a or b);
    outputs(9876) <= a xor b;
    outputs(9877) <= a xor b;
    outputs(9878) <= a or b;
    outputs(9879) <= a and b;
    outputs(9880) <= not (a xor b);
    outputs(9881) <= b and not a;
    outputs(9882) <= a xor b;
    outputs(9883) <= a and b;
    outputs(9884) <= not b;
    outputs(9885) <= b and not a;
    outputs(9886) <= a xor b;
    outputs(9887) <= a and b;
    outputs(9888) <= not a;
    outputs(9889) <= not (a xor b);
    outputs(9890) <= a xor b;
    outputs(9891) <= not a;
    outputs(9892) <= not b or a;
    outputs(9893) <= a xor b;
    outputs(9894) <= not (a xor b);
    outputs(9895) <= not b;
    outputs(9896) <= a xor b;
    outputs(9897) <= not a;
    outputs(9898) <= a or b;
    outputs(9899) <= not (a xor b);
    outputs(9900) <= not b or a;
    outputs(9901) <= a and b;
    outputs(9902) <= a;
    outputs(9903) <= not (a or b);
    outputs(9904) <= a xor b;
    outputs(9905) <= a and not b;
    outputs(9906) <= b;
    outputs(9907) <= not (a or b);
    outputs(9908) <= a xor b;
    outputs(9909) <= a xor b;
    outputs(9910) <= a;
    outputs(9911) <= b;
    outputs(9912) <= a;
    outputs(9913) <= not (a xor b);
    outputs(9914) <= not (a xor b);
    outputs(9915) <= not (a xor b);
    outputs(9916) <= a and b;
    outputs(9917) <= a;
    outputs(9918) <= not b;
    outputs(9919) <= not (a xor b);
    outputs(9920) <= a and b;
    outputs(9921) <= not (a or b);
    outputs(9922) <= not b;
    outputs(9923) <= not a;
    outputs(9924) <= not (a or b);
    outputs(9925) <= b;
    outputs(9926) <= not (a and b);
    outputs(9927) <= a xor b;
    outputs(9928) <= not (a xor b);
    outputs(9929) <= b;
    outputs(9930) <= a and not b;
    outputs(9931) <= a and b;
    outputs(9932) <= not (a xor b);
    outputs(9933) <= not (a xor b);
    outputs(9934) <= not a;
    outputs(9935) <= not (a or b);
    outputs(9936) <= not (a or b);
    outputs(9937) <= a and b;
    outputs(9938) <= a and b;
    outputs(9939) <= not a;
    outputs(9940) <= a and b;
    outputs(9941) <= b and not a;
    outputs(9942) <= a xor b;
    outputs(9943) <= not (a xor b);
    outputs(9944) <= not (a xor b);
    outputs(9945) <= a and not b;
    outputs(9946) <= a;
    outputs(9947) <= not a or b;
    outputs(9948) <= not b;
    outputs(9949) <= a xor b;
    outputs(9950) <= not (a xor b);
    outputs(9951) <= b;
    outputs(9952) <= not (a or b);
    outputs(9953) <= not a;
    outputs(9954) <= b;
    outputs(9955) <= not b;
    outputs(9956) <= a xor b;
    outputs(9957) <= b and not a;
    outputs(9958) <= not b;
    outputs(9959) <= not (a or b);
    outputs(9960) <= a and b;
    outputs(9961) <= not (a or b);
    outputs(9962) <= not (a xor b);
    outputs(9963) <= a;
    outputs(9964) <= b;
    outputs(9965) <= a xor b;
    outputs(9966) <= not a;
    outputs(9967) <= b;
    outputs(9968) <= b;
    outputs(9969) <= not a;
    outputs(9970) <= not (a xor b);
    outputs(9971) <= not a;
    outputs(9972) <= a and not b;
    outputs(9973) <= b;
    outputs(9974) <= a xor b;
    outputs(9975) <= not (a or b);
    outputs(9976) <= not a;
    outputs(9977) <= not (a xor b);
    outputs(9978) <= not (a or b);
    outputs(9979) <= not (a xor b);
    outputs(9980) <= not b or a;
    outputs(9981) <= a and b;
    outputs(9982) <= a;
    outputs(9983) <= a;
    outputs(9984) <= a and not b;
    outputs(9985) <= a and not b;
    outputs(9986) <= not a;
    outputs(9987) <= b;
    outputs(9988) <= not (a xor b);
    outputs(9989) <= a;
    outputs(9990) <= b;
    outputs(9991) <= not a;
    outputs(9992) <= a xor b;
    outputs(9993) <= not (a xor b);
    outputs(9994) <= b and not a;
    outputs(9995) <= b and not a;
    outputs(9996) <= a xor b;
    outputs(9997) <= a xor b;
    outputs(9998) <= 1'b0;
    outputs(9999) <= a xor b;
    outputs(10000) <= b and not a;
    outputs(10001) <= a;
    outputs(10002) <= not a or b;
    outputs(10003) <= a and b;
    outputs(10004) <= not (a xor b);
    outputs(10005) <= not a;
    outputs(10006) <= b;
    outputs(10007) <= a and b;
    outputs(10008) <= not a or b;
    outputs(10009) <= a xor b;
    outputs(10010) <= not (a xor b);
    outputs(10011) <= a;
    outputs(10012) <= not (a or b);
    outputs(10013) <= not (a or b);
    outputs(10014) <= not b or a;
    outputs(10015) <= b and not a;
    outputs(10016) <= a xor b;
    outputs(10017) <= a and b;
    outputs(10018) <= b;
    outputs(10019) <= not (a or b);
    outputs(10020) <= a or b;
    outputs(10021) <= not (a xor b);
    outputs(10022) <= a;
    outputs(10023) <= a xor b;
    outputs(10024) <= not b;
    outputs(10025) <= not b or a;
    outputs(10026) <= not b;
    outputs(10027) <= a and not b;
    outputs(10028) <= a or b;
    outputs(10029) <= a xor b;
    outputs(10030) <= a and b;
    outputs(10031) <= b and not a;
    outputs(10032) <= not a;
    outputs(10033) <= not a;
    outputs(10034) <= a xor b;
    outputs(10035) <= b and not a;
    outputs(10036) <= a;
    outputs(10037) <= not (a xor b);
    outputs(10038) <= not a;
    outputs(10039) <= b and not a;
    outputs(10040) <= not (a xor b);
    outputs(10041) <= a xor b;
    outputs(10042) <= a xor b;
    outputs(10043) <= a and b;
    outputs(10044) <= not a;
    outputs(10045) <= a;
    outputs(10046) <= not b or a;
    outputs(10047) <= a;
    outputs(10048) <= b and not a;
    outputs(10049) <= a xor b;
    outputs(10050) <= a;
    outputs(10051) <= b;
    outputs(10052) <= a xor b;
    outputs(10053) <= not b;
    outputs(10054) <= a and b;
    outputs(10055) <= a;
    outputs(10056) <= a xor b;
    outputs(10057) <= a or b;
    outputs(10058) <= not (a xor b);
    outputs(10059) <= a;
    outputs(10060) <= a xor b;
    outputs(10061) <= a xor b;
    outputs(10062) <= b and not a;
    outputs(10063) <= a;
    outputs(10064) <= a;
    outputs(10065) <= a xor b;
    outputs(10066) <= not a;
    outputs(10067) <= a;
    outputs(10068) <= not b;
    outputs(10069) <= a;
    outputs(10070) <= not b;
    outputs(10071) <= b;
    outputs(10072) <= b;
    outputs(10073) <= a xor b;
    outputs(10074) <= not b or a;
    outputs(10075) <= a and b;
    outputs(10076) <= a xor b;
    outputs(10077) <= a xor b;
    outputs(10078) <= b and not a;
    outputs(10079) <= b;
    outputs(10080) <= not b or a;
    outputs(10081) <= not (a or b);
    outputs(10082) <= not (a or b);
    outputs(10083) <= not (a xor b);
    outputs(10084) <= a xor b;
    outputs(10085) <= a;
    outputs(10086) <= not a;
    outputs(10087) <= b;
    outputs(10088) <= not (a or b);
    outputs(10089) <= b and not a;
    outputs(10090) <= a;
    outputs(10091) <= a and not b;
    outputs(10092) <= b;
    outputs(10093) <= b;
    outputs(10094) <= a and not b;
    outputs(10095) <= a xor b;
    outputs(10096) <= not a;
    outputs(10097) <= a and b;
    outputs(10098) <= a xor b;
    outputs(10099) <= a xor b;
    outputs(10100) <= a xor b;
    outputs(10101) <= not b;
    outputs(10102) <= a xor b;
    outputs(10103) <= not a;
    outputs(10104) <= not a or b;
    outputs(10105) <= not (a or b);
    outputs(10106) <= a or b;
    outputs(10107) <= b and not a;
    outputs(10108) <= a and b;
    outputs(10109) <= a;
    outputs(10110) <= a;
    outputs(10111) <= not b;
    outputs(10112) <= a xor b;
    outputs(10113) <= a xor b;
    outputs(10114) <= b and not a;
    outputs(10115) <= not (a xor b);
    outputs(10116) <= a xor b;
    outputs(10117) <= b;
    outputs(10118) <= a;
    outputs(10119) <= a xor b;
    outputs(10120) <= a xor b;
    outputs(10121) <= b and not a;
    outputs(10122) <= not a;
    outputs(10123) <= not b;
    outputs(10124) <= not a;
    outputs(10125) <= a;
    outputs(10126) <= a and b;
    outputs(10127) <= not a or b;
    outputs(10128) <= not (a and b);
    outputs(10129) <= not (a xor b);
    outputs(10130) <= not (a xor b);
    outputs(10131) <= not (a or b);
    outputs(10132) <= a xor b;
    outputs(10133) <= not a or b;
    outputs(10134) <= a or b;
    outputs(10135) <= b and not a;
    outputs(10136) <= a;
    outputs(10137) <= not (a or b);
    outputs(10138) <= a and b;
    outputs(10139) <= b and not a;
    outputs(10140) <= not (a xor b);
    outputs(10141) <= not a;
    outputs(10142) <= b;
    outputs(10143) <= a;
    outputs(10144) <= not b;
    outputs(10145) <= not (a and b);
    outputs(10146) <= not b;
    outputs(10147) <= b;
    outputs(10148) <= not b;
    outputs(10149) <= a and not b;
    outputs(10150) <= not (a xor b);
    outputs(10151) <= b and not a;
    outputs(10152) <= a and not b;
    outputs(10153) <= a;
    outputs(10154) <= not (a xor b);
    outputs(10155) <= not b;
    outputs(10156) <= not (a or b);
    outputs(10157) <= not a;
    outputs(10158) <= not (a xor b);
    outputs(10159) <= a xor b;
    outputs(10160) <= not a;
    outputs(10161) <= a and b;
    outputs(10162) <= a and not b;
    outputs(10163) <= not a;
    outputs(10164) <= not (a xor b);
    outputs(10165) <= not b;
    outputs(10166) <= a xor b;
    outputs(10167) <= not b;
    outputs(10168) <= b;
    outputs(10169) <= not (a and b);
    outputs(10170) <= a and not b;
    outputs(10171) <= not b or a;
    outputs(10172) <= a xor b;
    outputs(10173) <= a and b;
    outputs(10174) <= a xor b;
    outputs(10175) <= not (a xor b);
    outputs(10176) <= a xor b;
    outputs(10177) <= a xor b;
    outputs(10178) <= not a;
    outputs(10179) <= not b;
    outputs(10180) <= b and not a;
    outputs(10181) <= not b;
    outputs(10182) <= a;
    outputs(10183) <= not b;
    outputs(10184) <= b and not a;
    outputs(10185) <= b;
    outputs(10186) <= b;
    outputs(10187) <= not (a or b);
    outputs(10188) <= not (a xor b);
    outputs(10189) <= b and not a;
    outputs(10190) <= not b;
    outputs(10191) <= b;
    outputs(10192) <= not b;
    outputs(10193) <= a and not b;
    outputs(10194) <= b;
    outputs(10195) <= not (a xor b);
    outputs(10196) <= a or b;
    outputs(10197) <= a;
    outputs(10198) <= not (a and b);
    outputs(10199) <= b and not a;
    outputs(10200) <= not (a xor b);
    outputs(10201) <= not b or a;
    outputs(10202) <= b;
    outputs(10203) <= not (a xor b);
    outputs(10204) <= a;
    outputs(10205) <= a;
    outputs(10206) <= not a or b;
    outputs(10207) <= a xor b;
    outputs(10208) <= a and b;
    outputs(10209) <= not a;
    outputs(10210) <= not b;
    outputs(10211) <= not a;
    outputs(10212) <= b;
    outputs(10213) <= not (a xor b);
    outputs(10214) <= not a;
    outputs(10215) <= b;
    outputs(10216) <= not (a xor b);
    outputs(10217) <= not (a xor b);
    outputs(10218) <= b;
    outputs(10219) <= a and not b;
    outputs(10220) <= not a;
    outputs(10221) <= a xor b;
    outputs(10222) <= b;
    outputs(10223) <= not (a xor b);
    outputs(10224) <= not b or a;
    outputs(10225) <= not (a xor b);
    outputs(10226) <= a xor b;
    outputs(10227) <= not (a xor b);
    outputs(10228) <= a xor b;
    outputs(10229) <= b;
    outputs(10230) <= a xor b;
    outputs(10231) <= a and not b;
    outputs(10232) <= not (a xor b);
    outputs(10233) <= not a;
    outputs(10234) <= b;
    outputs(10235) <= not (a xor b);
    outputs(10236) <= a and not b;
    outputs(10237) <= a and not b;
    outputs(10238) <= not (a xor b);
    outputs(10239) <= not (a xor b);
    outputs(10240) <= not a;
    outputs(10241) <= not b;
    outputs(10242) <= b;
    outputs(10243) <= not (a and b);
    outputs(10244) <= not b or a;
    outputs(10245) <= a xor b;
    outputs(10246) <= b and not a;
    outputs(10247) <= not b;
    outputs(10248) <= not b or a;
    outputs(10249) <= not (a or b);
    outputs(10250) <= a xor b;
    outputs(10251) <= a;
    outputs(10252) <= a and b;
    outputs(10253) <= b;
    outputs(10254) <= not (a xor b);
    outputs(10255) <= not b;
    outputs(10256) <= not (a xor b);
    outputs(10257) <= not b or a;
    outputs(10258) <= not b or a;
    outputs(10259) <= not (a xor b);
    outputs(10260) <= not (a and b);
    outputs(10261) <= a;
    outputs(10262) <= not a;
    outputs(10263) <= a xor b;
    outputs(10264) <= not a or b;
    outputs(10265) <= not (a or b);
    outputs(10266) <= not (a xor b);
    outputs(10267) <= a xor b;
    outputs(10268) <= a or b;
    outputs(10269) <= b and not a;
    outputs(10270) <= a;
    outputs(10271) <= a and not b;
    outputs(10272) <= a or b;
    outputs(10273) <= a;
    outputs(10274) <= not a or b;
    outputs(10275) <= a;
    outputs(10276) <= not b;
    outputs(10277) <= not a;
    outputs(10278) <= not (a xor b);
    outputs(10279) <= not b;
    outputs(10280) <= a or b;
    outputs(10281) <= a;
    outputs(10282) <= a xor b;
    outputs(10283) <= a or b;
    outputs(10284) <= a;
    outputs(10285) <= a;
    outputs(10286) <= not (a xor b);
    outputs(10287) <= a;
    outputs(10288) <= a xor b;
    outputs(10289) <= a xor b;
    outputs(10290) <= b and not a;
    outputs(10291) <= a and b;
    outputs(10292) <= not b;
    outputs(10293) <= not a;
    outputs(10294) <= not a;
    outputs(10295) <= not (a or b);
    outputs(10296) <= not b;
    outputs(10297) <= not b;
    outputs(10298) <= b;
    outputs(10299) <= a;
    outputs(10300) <= a xor b;
    outputs(10301) <= b;
    outputs(10302) <= not (a xor b);
    outputs(10303) <= not (a or b);
    outputs(10304) <= a xor b;
    outputs(10305) <= not (a and b);
    outputs(10306) <= a or b;
    outputs(10307) <= not (a xor b);
    outputs(10308) <= not b;
    outputs(10309) <= b;
    outputs(10310) <= b and not a;
    outputs(10311) <= a xor b;
    outputs(10312) <= not (a and b);
    outputs(10313) <= a xor b;
    outputs(10314) <= a xor b;
    outputs(10315) <= b and not a;
    outputs(10316) <= a;
    outputs(10317) <= a or b;
    outputs(10318) <= a or b;
    outputs(10319) <= a xor b;
    outputs(10320) <= not a;
    outputs(10321) <= not (a and b);
    outputs(10322) <= not a;
    outputs(10323) <= not b;
    outputs(10324) <= not (a xor b);
    outputs(10325) <= not a or b;
    outputs(10326) <= not b or a;
    outputs(10327) <= a xor b;
    outputs(10328) <= not b or a;
    outputs(10329) <= a xor b;
    outputs(10330) <= a xor b;
    outputs(10331) <= a;
    outputs(10332) <= a or b;
    outputs(10333) <= not b;
    outputs(10334) <= a xor b;
    outputs(10335) <= not (a xor b);
    outputs(10336) <= a;
    outputs(10337) <= not b;
    outputs(10338) <= not b or a;
    outputs(10339) <= a;
    outputs(10340) <= not b;
    outputs(10341) <= not (a and b);
    outputs(10342) <= a;
    outputs(10343) <= a;
    outputs(10344) <= a xor b;
    outputs(10345) <= a;
    outputs(10346) <= b;
    outputs(10347) <= a or b;
    outputs(10348) <= a;
    outputs(10349) <= a xor b;
    outputs(10350) <= not b;
    outputs(10351) <= not (a xor b);
    outputs(10352) <= not a or b;
    outputs(10353) <= not (a xor b);
    outputs(10354) <= not (a or b);
    outputs(10355) <= a xor b;
    outputs(10356) <= not (a xor b);
    outputs(10357) <= b and not a;
    outputs(10358) <= not (a and b);
    outputs(10359) <= not b;
    outputs(10360) <= a and not b;
    outputs(10361) <= not a;
    outputs(10362) <= a xor b;
    outputs(10363) <= a xor b;
    outputs(10364) <= a or b;
    outputs(10365) <= a or b;
    outputs(10366) <= not a;
    outputs(10367) <= not (a and b);
    outputs(10368) <= a xor b;
    outputs(10369) <= a xor b;
    outputs(10370) <= not b;
    outputs(10371) <= not b;
    outputs(10372) <= b;
    outputs(10373) <= not (a or b);
    outputs(10374) <= a;
    outputs(10375) <= not a;
    outputs(10376) <= not a;
    outputs(10377) <= not (a xor b);
    outputs(10378) <= a;
    outputs(10379) <= not a;
    outputs(10380) <= not (a xor b);
    outputs(10381) <= a;
    outputs(10382) <= not b or a;
    outputs(10383) <= a or b;
    outputs(10384) <= b;
    outputs(10385) <= not (a xor b);
    outputs(10386) <= not (a xor b);
    outputs(10387) <= b;
    outputs(10388) <= a;
    outputs(10389) <= not a or b;
    outputs(10390) <= a xor b;
    outputs(10391) <= a xor b;
    outputs(10392) <= not b or a;
    outputs(10393) <= not b or a;
    outputs(10394) <= not (a xor b);
    outputs(10395) <= not b;
    outputs(10396) <= a and b;
    outputs(10397) <= not b or a;
    outputs(10398) <= not (a xor b);
    outputs(10399) <= a or b;
    outputs(10400) <= a xor b;
    outputs(10401) <= a or b;
    outputs(10402) <= a;
    outputs(10403) <= a;
    outputs(10404) <= not a;
    outputs(10405) <= not (a xor b);
    outputs(10406) <= b;
    outputs(10407) <= b;
    outputs(10408) <= not b or a;
    outputs(10409) <= not (a xor b);
    outputs(10410) <= not (a xor b);
    outputs(10411) <= a;
    outputs(10412) <= not (a xor b);
    outputs(10413) <= a or b;
    outputs(10414) <= b;
    outputs(10415) <= not (a or b);
    outputs(10416) <= b;
    outputs(10417) <= a xor b;
    outputs(10418) <= a and not b;
    outputs(10419) <= not a or b;
    outputs(10420) <= not b or a;
    outputs(10421) <= a;
    outputs(10422) <= not (a xor b);
    outputs(10423) <= not b or a;
    outputs(10424) <= not (a xor b);
    outputs(10425) <= a;
    outputs(10426) <= a;
    outputs(10427) <= a xor b;
    outputs(10428) <= b;
    outputs(10429) <= not a;
    outputs(10430) <= not a or b;
    outputs(10431) <= not a;
    outputs(10432) <= a xor b;
    outputs(10433) <= not b or a;
    outputs(10434) <= not b;
    outputs(10435) <= not (a xor b);
    outputs(10436) <= not (a and b);
    outputs(10437) <= not (a xor b);
    outputs(10438) <= not b;
    outputs(10439) <= not b;
    outputs(10440) <= not b;
    outputs(10441) <= a;
    outputs(10442) <= a and not b;
    outputs(10443) <= not (a xor b);
    outputs(10444) <= a or b;
    outputs(10445) <= not (a xor b);
    outputs(10446) <= a;
    outputs(10447) <= not (a xor b);
    outputs(10448) <= b;
    outputs(10449) <= a and b;
    outputs(10450) <= a or b;
    outputs(10451) <= b and not a;
    outputs(10452) <= not b;
    outputs(10453) <= not (a xor b);
    outputs(10454) <= a xor b;
    outputs(10455) <= not (a xor b);
    outputs(10456) <= not b or a;
    outputs(10457) <= b;
    outputs(10458) <= not b or a;
    outputs(10459) <= b;
    outputs(10460) <= a xor b;
    outputs(10461) <= a xor b;
    outputs(10462) <= not a;
    outputs(10463) <= b and not a;
    outputs(10464) <= not a;
    outputs(10465) <= b and not a;
    outputs(10466) <= b;
    outputs(10467) <= b;
    outputs(10468) <= not a;
    outputs(10469) <= b;
    outputs(10470) <= b;
    outputs(10471) <= not (a xor b);
    outputs(10472) <= not (a xor b);
    outputs(10473) <= not b;
    outputs(10474) <= b;
    outputs(10475) <= a xor b;
    outputs(10476) <= a xor b;
    outputs(10477) <= b;
    outputs(10478) <= not (a xor b);
    outputs(10479) <= a and b;
    outputs(10480) <= not b or a;
    outputs(10481) <= a;
    outputs(10482) <= not a;
    outputs(10483) <= a and not b;
    outputs(10484) <= a;
    outputs(10485) <= a xor b;
    outputs(10486) <= b;
    outputs(10487) <= a xor b;
    outputs(10488) <= a or b;
    outputs(10489) <= a xor b;
    outputs(10490) <= a and b;
    outputs(10491) <= not (a xor b);
    outputs(10492) <= a xor b;
    outputs(10493) <= not a or b;
    outputs(10494) <= a;
    outputs(10495) <= not (a xor b);
    outputs(10496) <= a xor b;
    outputs(10497) <= not a;
    outputs(10498) <= not (a xor b);
    outputs(10499) <= a;
    outputs(10500) <= a xor b;
    outputs(10501) <= not a;
    outputs(10502) <= b;
    outputs(10503) <= not a or b;
    outputs(10504) <= a;
    outputs(10505) <= not (a xor b);
    outputs(10506) <= a or b;
    outputs(10507) <= not (a xor b);
    outputs(10508) <= not b;
    outputs(10509) <= not b or a;
    outputs(10510) <= not a;
    outputs(10511) <= a or b;
    outputs(10512) <= a xor b;
    outputs(10513) <= b;
    outputs(10514) <= not b or a;
    outputs(10515) <= not (a and b);
    outputs(10516) <= not a or b;
    outputs(10517) <= not (a xor b);
    outputs(10518) <= not b;
    outputs(10519) <= a xor b;
    outputs(10520) <= not a or b;
    outputs(10521) <= not b or a;
    outputs(10522) <= a xor b;
    outputs(10523) <= b and not a;
    outputs(10524) <= a xor b;
    outputs(10525) <= not (a xor b);
    outputs(10526) <= not b;
    outputs(10527) <= a and not b;
    outputs(10528) <= a;
    outputs(10529) <= a;
    outputs(10530) <= not (a and b);
    outputs(10531) <= not b;
    outputs(10532) <= not (a or b);
    outputs(10533) <= a and b;
    outputs(10534) <= not b or a;
    outputs(10535) <= not b or a;
    outputs(10536) <= not (a xor b);
    outputs(10537) <= a;
    outputs(10538) <= not a;
    outputs(10539) <= a xor b;
    outputs(10540) <= not (a and b);
    outputs(10541) <= a xor b;
    outputs(10542) <= not (a xor b);
    outputs(10543) <= not (a and b);
    outputs(10544) <= a and not b;
    outputs(10545) <= not b;
    outputs(10546) <= b;
    outputs(10547) <= not b or a;
    outputs(10548) <= not b or a;
    outputs(10549) <= not (a xor b);
    outputs(10550) <= a;
    outputs(10551) <= a or b;
    outputs(10552) <= a xor b;
    outputs(10553) <= a;
    outputs(10554) <= a;
    outputs(10555) <= b;
    outputs(10556) <= a;
    outputs(10557) <= a;
    outputs(10558) <= b and not a;
    outputs(10559) <= not (a and b);
    outputs(10560) <= a or b;
    outputs(10561) <= not b or a;
    outputs(10562) <= b and not a;
    outputs(10563) <= a and b;
    outputs(10564) <= not (a and b);
    outputs(10565) <= b;
    outputs(10566) <= b and not a;
    outputs(10567) <= not b;
    outputs(10568) <= a and not b;
    outputs(10569) <= not b;
    outputs(10570) <= not (a xor b);
    outputs(10571) <= b and not a;
    outputs(10572) <= a xor b;
    outputs(10573) <= not b;
    outputs(10574) <= not (a xor b);
    outputs(10575) <= not b or a;
    outputs(10576) <= b;
    outputs(10577) <= not a;
    outputs(10578) <= a and not b;
    outputs(10579) <= b and not a;
    outputs(10580) <= not a;
    outputs(10581) <= a xor b;
    outputs(10582) <= a or b;
    outputs(10583) <= not a;
    outputs(10584) <= a xor b;
    outputs(10585) <= not b or a;
    outputs(10586) <= not b;
    outputs(10587) <= a or b;
    outputs(10588) <= a;
    outputs(10589) <= b;
    outputs(10590) <= a xor b;
    outputs(10591) <= not (a and b);
    outputs(10592) <= not (a xor b);
    outputs(10593) <= not (a or b);
    outputs(10594) <= not (a xor b);
    outputs(10595) <= a xor b;
    outputs(10596) <= not (a or b);
    outputs(10597) <= a;
    outputs(10598) <= a xor b;
    outputs(10599) <= not (a xor b);
    outputs(10600) <= a xor b;
    outputs(10601) <= not (a xor b);
    outputs(10602) <= not a;
    outputs(10603) <= not b;
    outputs(10604) <= b;
    outputs(10605) <= a;
    outputs(10606) <= not (a xor b);
    outputs(10607) <= not b or a;
    outputs(10608) <= a or b;
    outputs(10609) <= b;
    outputs(10610) <= not a;
    outputs(10611) <= a xor b;
    outputs(10612) <= a xor b;
    outputs(10613) <= a;
    outputs(10614) <= not (a xor b);
    outputs(10615) <= a;
    outputs(10616) <= a xor b;
    outputs(10617) <= a and not b;
    outputs(10618) <= not a;
    outputs(10619) <= a;
    outputs(10620) <= a xor b;
    outputs(10621) <= not a;
    outputs(10622) <= not (a or b);
    outputs(10623) <= a;
    outputs(10624) <= not a;
    outputs(10625) <= a xor b;
    outputs(10626) <= b and not a;
    outputs(10627) <= not a;
    outputs(10628) <= not (a xor b);
    outputs(10629) <= not b;
    outputs(10630) <= not b;
    outputs(10631) <= not b;
    outputs(10632) <= not b;
    outputs(10633) <= a xor b;
    outputs(10634) <= a xor b;
    outputs(10635) <= a;
    outputs(10636) <= a and not b;
    outputs(10637) <= not (a xor b);
    outputs(10638) <= not a or b;
    outputs(10639) <= b;
    outputs(10640) <= a xor b;
    outputs(10641) <= a xor b;
    outputs(10642) <= b;
    outputs(10643) <= a xor b;
    outputs(10644) <= not (a xor b);
    outputs(10645) <= a xor b;
    outputs(10646) <= a;
    outputs(10647) <= a xor b;
    outputs(10648) <= a xor b;
    outputs(10649) <= b;
    outputs(10650) <= not a or b;
    outputs(10651) <= b;
    outputs(10652) <= a;
    outputs(10653) <= b;
    outputs(10654) <= not a;
    outputs(10655) <= not b or a;
    outputs(10656) <= not a or b;
    outputs(10657) <= a xor b;
    outputs(10658) <= not (a xor b);
    outputs(10659) <= not a;
    outputs(10660) <= not b or a;
    outputs(10661) <= not b;
    outputs(10662) <= not a;
    outputs(10663) <= b and not a;
    outputs(10664) <= not b or a;
    outputs(10665) <= a xor b;
    outputs(10666) <= b;
    outputs(10667) <= a;
    outputs(10668) <= not (a xor b);
    outputs(10669) <= a xor b;
    outputs(10670) <= a;
    outputs(10671) <= a;
    outputs(10672) <= a xor b;
    outputs(10673) <= a or b;
    outputs(10674) <= a xor b;
    outputs(10675) <= not (a and b);
    outputs(10676) <= not a or b;
    outputs(10677) <= not (a and b);
    outputs(10678) <= not a;
    outputs(10679) <= b;
    outputs(10680) <= not (a xor b);
    outputs(10681) <= a xor b;
    outputs(10682) <= not b or a;
    outputs(10683) <= not a or b;
    outputs(10684) <= not (a xor b);
    outputs(10685) <= not b or a;
    outputs(10686) <= a xor b;
    outputs(10687) <= a xor b;
    outputs(10688) <= a xor b;
    outputs(10689) <= not (a xor b);
    outputs(10690) <= not (a xor b);
    outputs(10691) <= not (a xor b);
    outputs(10692) <= not (a or b);
    outputs(10693) <= not b;
    outputs(10694) <= not b;
    outputs(10695) <= a and not b;
    outputs(10696) <= not a or b;
    outputs(10697) <= b;
    outputs(10698) <= b;
    outputs(10699) <= b;
    outputs(10700) <= not b;
    outputs(10701) <= not (a xor b);
    outputs(10702) <= not b;
    outputs(10703) <= a xor b;
    outputs(10704) <= b;
    outputs(10705) <= a;
    outputs(10706) <= not (a and b);
    outputs(10707) <= a and not b;
    outputs(10708) <= not (a or b);
    outputs(10709) <= a;
    outputs(10710) <= a xor b;
    outputs(10711) <= a and b;
    outputs(10712) <= a xor b;
    outputs(10713) <= not a;
    outputs(10714) <= a and not b;
    outputs(10715) <= a and b;
    outputs(10716) <= not a;
    outputs(10717) <= a;
    outputs(10718) <= not b or a;
    outputs(10719) <= not (a xor b);
    outputs(10720) <= a xor b;
    outputs(10721) <= a xor b;
    outputs(10722) <= not a;
    outputs(10723) <= b;
    outputs(10724) <= b;
    outputs(10725) <= a and not b;
    outputs(10726) <= a;
    outputs(10727) <= not (a xor b);
    outputs(10728) <= b and not a;
    outputs(10729) <= a;
    outputs(10730) <= not b;
    outputs(10731) <= a or b;
    outputs(10732) <= b;
    outputs(10733) <= a or b;
    outputs(10734) <= a xor b;
    outputs(10735) <= a xor b;
    outputs(10736) <= not a;
    outputs(10737) <= not b or a;
    outputs(10738) <= a xor b;
    outputs(10739) <= a;
    outputs(10740) <= not b or a;
    outputs(10741) <= not (a xor b);
    outputs(10742) <= not a;
    outputs(10743) <= a xor b;
    outputs(10744) <= not a;
    outputs(10745) <= not a or b;
    outputs(10746) <= not a;
    outputs(10747) <= not (a xor b);
    outputs(10748) <= not b;
    outputs(10749) <= a xor b;
    outputs(10750) <= not b or a;
    outputs(10751) <= not (a xor b);
    outputs(10752) <= a;
    outputs(10753) <= a xor b;
    outputs(10754) <= not a;
    outputs(10755) <= a;
    outputs(10756) <= not (a xor b);
    outputs(10757) <= not b;
    outputs(10758) <= not (a and b);
    outputs(10759) <= not a or b;
    outputs(10760) <= not a;
    outputs(10761) <= b and not a;
    outputs(10762) <= b and not a;
    outputs(10763) <= not b;
    outputs(10764) <= not a;
    outputs(10765) <= not (a xor b);
    outputs(10766) <= a or b;
    outputs(10767) <= a;
    outputs(10768) <= b;
    outputs(10769) <= b and not a;
    outputs(10770) <= not (a xor b);
    outputs(10771) <= not a;
    outputs(10772) <= a or b;
    outputs(10773) <= a xor b;
    outputs(10774) <= not (a xor b);
    outputs(10775) <= not a;
    outputs(10776) <= b;
    outputs(10777) <= a or b;
    outputs(10778) <= not a;
    outputs(10779) <= not (a or b);
    outputs(10780) <= not b;
    outputs(10781) <= a xor b;
    outputs(10782) <= not (a xor b);
    outputs(10783) <= a xor b;
    outputs(10784) <= not a or b;
    outputs(10785) <= not (a xor b);
    outputs(10786) <= a xor b;
    outputs(10787) <= not (a and b);
    outputs(10788) <= a xor b;
    outputs(10789) <= a xor b;
    outputs(10790) <= not a;
    outputs(10791) <= not a;
    outputs(10792) <= not a;
    outputs(10793) <= a xor b;
    outputs(10794) <= a xor b;
    outputs(10795) <= a or b;
    outputs(10796) <= a and b;
    outputs(10797) <= a and not b;
    outputs(10798) <= a or b;
    outputs(10799) <= b;
    outputs(10800) <= a;
    outputs(10801) <= a;
    outputs(10802) <= a and b;
    outputs(10803) <= a;
    outputs(10804) <= b;
    outputs(10805) <= not b;
    outputs(10806) <= b;
    outputs(10807) <= not (a xor b);
    outputs(10808) <= b;
    outputs(10809) <= a xor b;
    outputs(10810) <= not b or a;
    outputs(10811) <= a xor b;
    outputs(10812) <= not b;
    outputs(10813) <= b;
    outputs(10814) <= a and not b;
    outputs(10815) <= not b;
    outputs(10816) <= a xor b;
    outputs(10817) <= not a;
    outputs(10818) <= a xor b;
    outputs(10819) <= a and not b;
    outputs(10820) <= not (a xor b);
    outputs(10821) <= not (a or b);
    outputs(10822) <= not (a xor b);
    outputs(10823) <= not b;
    outputs(10824) <= not a;
    outputs(10825) <= not a or b;
    outputs(10826) <= a and b;
    outputs(10827) <= b and not a;
    outputs(10828) <= a and not b;
    outputs(10829) <= a or b;
    outputs(10830) <= not (a xor b);
    outputs(10831) <= not (a xor b);
    outputs(10832) <= a;
    outputs(10833) <= not a;
    outputs(10834) <= a or b;
    outputs(10835) <= a or b;
    outputs(10836) <= a xor b;
    outputs(10837) <= b and not a;
    outputs(10838) <= b;
    outputs(10839) <= not (a xor b);
    outputs(10840) <= not b or a;
    outputs(10841) <= not a or b;
    outputs(10842) <= not (a xor b);
    outputs(10843) <= not b;
    outputs(10844) <= b;
    outputs(10845) <= a;
    outputs(10846) <= not (a xor b);
    outputs(10847) <= b;
    outputs(10848) <= not b;
    outputs(10849) <= a xor b;
    outputs(10850) <= not b;
    outputs(10851) <= not (a and b);
    outputs(10852) <= a xor b;
    outputs(10853) <= not b;
    outputs(10854) <= b;
    outputs(10855) <= a or b;
    outputs(10856) <= not (a xor b);
    outputs(10857) <= not (a and b);
    outputs(10858) <= not b;
    outputs(10859) <= b and not a;
    outputs(10860) <= not (a xor b);
    outputs(10861) <= a xor b;
    outputs(10862) <= not a;
    outputs(10863) <= not (a xor b);
    outputs(10864) <= b;
    outputs(10865) <= not b;
    outputs(10866) <= a xor b;
    outputs(10867) <= not b;
    outputs(10868) <= b;
    outputs(10869) <= not (a and b);
    outputs(10870) <= a xor b;
    outputs(10871) <= not (a xor b);
    outputs(10872) <= a and not b;
    outputs(10873) <= not (a xor b);
    outputs(10874) <= a and b;
    outputs(10875) <= not (a xor b);
    outputs(10876) <= not (a xor b);
    outputs(10877) <= not a;
    outputs(10878) <= a or b;
    outputs(10879) <= a;
    outputs(10880) <= not (a xor b);
    outputs(10881) <= not (a xor b);
    outputs(10882) <= not b;
    outputs(10883) <= not a or b;
    outputs(10884) <= a xor b;
    outputs(10885) <= not (a xor b);
    outputs(10886) <= a;
    outputs(10887) <= not a;
    outputs(10888) <= not b;
    outputs(10889) <= a and not b;
    outputs(10890) <= b and not a;
    outputs(10891) <= not a;
    outputs(10892) <= not b or a;
    outputs(10893) <= not (a or b);
    outputs(10894) <= a xor b;
    outputs(10895) <= a;
    outputs(10896) <= a and b;
    outputs(10897) <= not b;
    outputs(10898) <= not a or b;
    outputs(10899) <= not (a xor b);
    outputs(10900) <= a or b;
    outputs(10901) <= a;
    outputs(10902) <= b;
    outputs(10903) <= not a or b;
    outputs(10904) <= b;
    outputs(10905) <= b;
    outputs(10906) <= not (a xor b);
    outputs(10907) <= a xor b;
    outputs(10908) <= a xor b;
    outputs(10909) <= not (a xor b);
    outputs(10910) <= not (a or b);
    outputs(10911) <= not (a xor b);
    outputs(10912) <= a and not b;
    outputs(10913) <= a or b;
    outputs(10914) <= not (a xor b);
    outputs(10915) <= not (a xor b);
    outputs(10916) <= not (a xor b);
    outputs(10917) <= not (a xor b);
    outputs(10918) <= a;
    outputs(10919) <= 1'b1;
    outputs(10920) <= a xor b;
    outputs(10921) <= not (a xor b);
    outputs(10922) <= a;
    outputs(10923) <= not a;
    outputs(10924) <= not b;
    outputs(10925) <= not (a xor b);
    outputs(10926) <= a xor b;
    outputs(10927) <= not b;
    outputs(10928) <= a xor b;
    outputs(10929) <= b and not a;
    outputs(10930) <= b;
    outputs(10931) <= b;
    outputs(10932) <= not a;
    outputs(10933) <= not b;
    outputs(10934) <= not b;
    outputs(10935) <= not (a xor b);
    outputs(10936) <= a xor b;
    outputs(10937) <= not b;
    outputs(10938) <= a;
    outputs(10939) <= a xor b;
    outputs(10940) <= not (a xor b);
    outputs(10941) <= b;
    outputs(10942) <= a;
    outputs(10943) <= not (a or b);
    outputs(10944) <= a;
    outputs(10945) <= a xor b;
    outputs(10946) <= b and not a;
    outputs(10947) <= not (a or b);
    outputs(10948) <= a and b;
    outputs(10949) <= not b or a;
    outputs(10950) <= a xor b;
    outputs(10951) <= a xor b;
    outputs(10952) <= not (a xor b);
    outputs(10953) <= b and not a;
    outputs(10954) <= a;
    outputs(10955) <= not (a and b);
    outputs(10956) <= not a;
    outputs(10957) <= not b or a;
    outputs(10958) <= a xor b;
    outputs(10959) <= a xor b;
    outputs(10960) <= b;
    outputs(10961) <= a xor b;
    outputs(10962) <= a xor b;
    outputs(10963) <= not a;
    outputs(10964) <= not (a xor b);
    outputs(10965) <= a xor b;
    outputs(10966) <= not (a xor b);
    outputs(10967) <= a xor b;
    outputs(10968) <= a xor b;
    outputs(10969) <= not (a and b);
    outputs(10970) <= a or b;
    outputs(10971) <= a xor b;
    outputs(10972) <= a xor b;
    outputs(10973) <= a xor b;
    outputs(10974) <= not a or b;
    outputs(10975) <= a and b;
    outputs(10976) <= a;
    outputs(10977) <= a and b;
    outputs(10978) <= not (a xor b);
    outputs(10979) <= not b;
    outputs(10980) <= not (a or b);
    outputs(10981) <= a;
    outputs(10982) <= not (a and b);
    outputs(10983) <= a xor b;
    outputs(10984) <= not (a and b);
    outputs(10985) <= a;
    outputs(10986) <= not a;
    outputs(10987) <= not (a and b);
    outputs(10988) <= b;
    outputs(10989) <= not a;
    outputs(10990) <= not (a xor b);
    outputs(10991) <= a;
    outputs(10992) <= a xor b;
    outputs(10993) <= a or b;
    outputs(10994) <= a;
    outputs(10995) <= a and b;
    outputs(10996) <= a and not b;
    outputs(10997) <= not (a xor b);
    outputs(10998) <= b;
    outputs(10999) <= not a or b;
    outputs(11000) <= a;
    outputs(11001) <= not a;
    outputs(11002) <= not a or b;
    outputs(11003) <= not a;
    outputs(11004) <= a xor b;
    outputs(11005) <= not a or b;
    outputs(11006) <= not b or a;
    outputs(11007) <= b and not a;
    outputs(11008) <= a;
    outputs(11009) <= not b or a;
    outputs(11010) <= a;
    outputs(11011) <= b;
    outputs(11012) <= not b;
    outputs(11013) <= b and not a;
    outputs(11014) <= a xor b;
    outputs(11015) <= not (a xor b);
    outputs(11016) <= not b or a;
    outputs(11017) <= b;
    outputs(11018) <= not b or a;
    outputs(11019) <= not (a and b);
    outputs(11020) <= a and not b;
    outputs(11021) <= not (a xor b);
    outputs(11022) <= not (a xor b);
    outputs(11023) <= not (a xor b);
    outputs(11024) <= a xor b;
    outputs(11025) <= not (a and b);
    outputs(11026) <= not (a xor b);
    outputs(11027) <= not b;
    outputs(11028) <= b;
    outputs(11029) <= a and b;
    outputs(11030) <= not a;
    outputs(11031) <= not b;
    outputs(11032) <= a or b;
    outputs(11033) <= not (a xor b);
    outputs(11034) <= a;
    outputs(11035) <= not (a or b);
    outputs(11036) <= b;
    outputs(11037) <= a or b;
    outputs(11038) <= b;
    outputs(11039) <= not a;
    outputs(11040) <= a xor b;
    outputs(11041) <= b;
    outputs(11042) <= a;
    outputs(11043) <= not (a xor b);
    outputs(11044) <= not (a and b);
    outputs(11045) <= not (a xor b);
    outputs(11046) <= a xor b;
    outputs(11047) <= b and not a;
    outputs(11048) <= not (a or b);
    outputs(11049) <= a xor b;
    outputs(11050) <= not b or a;
    outputs(11051) <= not (a xor b);
    outputs(11052) <= not a;
    outputs(11053) <= not a;
    outputs(11054) <= b;
    outputs(11055) <= not b;
    outputs(11056) <= a or b;
    outputs(11057) <= not (a xor b);
    outputs(11058) <= a xor b;
    outputs(11059) <= b;
    outputs(11060) <= not a;
    outputs(11061) <= a xor b;
    outputs(11062) <= a xor b;
    outputs(11063) <= not a;
    outputs(11064) <= a or b;
    outputs(11065) <= not (a and b);
    outputs(11066) <= not (a xor b);
    outputs(11067) <= a and b;
    outputs(11068) <= a or b;
    outputs(11069) <= a xor b;
    outputs(11070) <= not (a xor b);
    outputs(11071) <= not (a xor b);
    outputs(11072) <= not b;
    outputs(11073) <= not b or a;
    outputs(11074) <= a xor b;
    outputs(11075) <= not (a or b);
    outputs(11076) <= a xor b;
    outputs(11077) <= not (a xor b);
    outputs(11078) <= a xor b;
    outputs(11079) <= not (a xor b);
    outputs(11080) <= not (a xor b);
    outputs(11081) <= not a or b;
    outputs(11082) <= not (a xor b);
    outputs(11083) <= not (a xor b);
    outputs(11084) <= b;
    outputs(11085) <= a;
    outputs(11086) <= not (a and b);
    outputs(11087) <= a and not b;
    outputs(11088) <= not a or b;
    outputs(11089) <= not (a xor b);
    outputs(11090) <= not a;
    outputs(11091) <= a xor b;
    outputs(11092) <= b;
    outputs(11093) <= a xor b;
    outputs(11094) <= a xor b;
    outputs(11095) <= a;
    outputs(11096) <= not a;
    outputs(11097) <= not b;
    outputs(11098) <= not (a xor b);
    outputs(11099) <= b;
    outputs(11100) <= not a;
    outputs(11101) <= not a or b;
    outputs(11102) <= not b;
    outputs(11103) <= not a;
    outputs(11104) <= a xor b;
    outputs(11105) <= a;
    outputs(11106) <= a;
    outputs(11107) <= not (a xor b);
    outputs(11108) <= a xor b;
    outputs(11109) <= not a;
    outputs(11110) <= not (a xor b);
    outputs(11111) <= a xor b;
    outputs(11112) <= a xor b;
    outputs(11113) <= a and not b;
    outputs(11114) <= not a;
    outputs(11115) <= not b;
    outputs(11116) <= a and not b;
    outputs(11117) <= not b;
    outputs(11118) <= a;
    outputs(11119) <= not (a and b);
    outputs(11120) <= a xor b;
    outputs(11121) <= not b;
    outputs(11122) <= not (a xor b);
    outputs(11123) <= a;
    outputs(11124) <= b;
    outputs(11125) <= not (a xor b);
    outputs(11126) <= a or b;
    outputs(11127) <= b;
    outputs(11128) <= a xor b;
    outputs(11129) <= not b;
    outputs(11130) <= not (a xor b);
    outputs(11131) <= a or b;
    outputs(11132) <= a;
    outputs(11133) <= a xor b;
    outputs(11134) <= not (a or b);
    outputs(11135) <= b;
    outputs(11136) <= a xor b;
    outputs(11137) <= not a or b;
    outputs(11138) <= a;
    outputs(11139) <= a and b;
    outputs(11140) <= not (a or b);
    outputs(11141) <= b;
    outputs(11142) <= a xor b;
    outputs(11143) <= not b;
    outputs(11144) <= a;
    outputs(11145) <= b;
    outputs(11146) <= not (a or b);
    outputs(11147) <= a;
    outputs(11148) <= b;
    outputs(11149) <= a;
    outputs(11150) <= a;
    outputs(11151) <= a or b;
    outputs(11152) <= not b;
    outputs(11153) <= b and not a;
    outputs(11154) <= not (a and b);
    outputs(11155) <= not a;
    outputs(11156) <= a;
    outputs(11157) <= a xor b;
    outputs(11158) <= not b;
    outputs(11159) <= a;
    outputs(11160) <= not a or b;
    outputs(11161) <= a xor b;
    outputs(11162) <= not a;
    outputs(11163) <= not b or a;
    outputs(11164) <= not (a xor b);
    outputs(11165) <= not b or a;
    outputs(11166) <= a xor b;
    outputs(11167) <= not a or b;
    outputs(11168) <= not (a or b);
    outputs(11169) <= b;
    outputs(11170) <= not (a xor b);
    outputs(11171) <= a;
    outputs(11172) <= a xor b;
    outputs(11173) <= a;
    outputs(11174) <= not (a xor b);
    outputs(11175) <= not a;
    outputs(11176) <= b;
    outputs(11177) <= a xor b;
    outputs(11178) <= not (a xor b);
    outputs(11179) <= not a;
    outputs(11180) <= a xor b;
    outputs(11181) <= not (a xor b);
    outputs(11182) <= a xor b;
    outputs(11183) <= not a;
    outputs(11184) <= a xor b;
    outputs(11185) <= a and not b;
    outputs(11186) <= not a;
    outputs(11187) <= not (a and b);
    outputs(11188) <= b;
    outputs(11189) <= not a;
    outputs(11190) <= a;
    outputs(11191) <= not a or b;
    outputs(11192) <= not (a xor b);
    outputs(11193) <= not a;
    outputs(11194) <= a xor b;
    outputs(11195) <= a;
    outputs(11196) <= not (a xor b);
    outputs(11197) <= not a;
    outputs(11198) <= b;
    outputs(11199) <= a or b;
    outputs(11200) <= not (a xor b);
    outputs(11201) <= b;
    outputs(11202) <= not (a and b);
    outputs(11203) <= not a;
    outputs(11204) <= a xor b;
    outputs(11205) <= not (a and b);
    outputs(11206) <= not (a xor b);
    outputs(11207) <= 1'b1;
    outputs(11208) <= a or b;
    outputs(11209) <= not a or b;
    outputs(11210) <= b and not a;
    outputs(11211) <= a xor b;
    outputs(11212) <= not a or b;
    outputs(11213) <= not b;
    outputs(11214) <= b;
    outputs(11215) <= not (a and b);
    outputs(11216) <= b;
    outputs(11217) <= not (a xor b);
    outputs(11218) <= not (a xor b);
    outputs(11219) <= not (a xor b);
    outputs(11220) <= not a;
    outputs(11221) <= not a or b;
    outputs(11222) <= not b or a;
    outputs(11223) <= not b;
    outputs(11224) <= b;
    outputs(11225) <= not a;
    outputs(11226) <= b and not a;
    outputs(11227) <= not (a xor b);
    outputs(11228) <= a or b;
    outputs(11229) <= b;
    outputs(11230) <= not (a xor b);
    outputs(11231) <= not (a and b);
    outputs(11232) <= not (a xor b);
    outputs(11233) <= not a or b;
    outputs(11234) <= b;
    outputs(11235) <= not (a or b);
    outputs(11236) <= not (a xor b);
    outputs(11237) <= b;
    outputs(11238) <= a or b;
    outputs(11239) <= a xor b;
    outputs(11240) <= not (a and b);
    outputs(11241) <= a xor b;
    outputs(11242) <= a xor b;
    outputs(11243) <= not (a xor b);
    outputs(11244) <= not b;
    outputs(11245) <= a or b;
    outputs(11246) <= b and not a;
    outputs(11247) <= not b;
    outputs(11248) <= a or b;
    outputs(11249) <= not (a xor b);
    outputs(11250) <= not b;
    outputs(11251) <= not b;
    outputs(11252) <= b;
    outputs(11253) <= not (a xor b);
    outputs(11254) <= not (a xor b);
    outputs(11255) <= a;
    outputs(11256) <= not (a xor b);
    outputs(11257) <= a xor b;
    outputs(11258) <= a and not b;
    outputs(11259) <= not (a xor b);
    outputs(11260) <= not b;
    outputs(11261) <= a xor b;
    outputs(11262) <= not (a xor b);
    outputs(11263) <= a;
    outputs(11264) <= b;
    outputs(11265) <= not b;
    outputs(11266) <= a or b;
    outputs(11267) <= a xor b;
    outputs(11268) <= not (a xor b);
    outputs(11269) <= not a or b;
    outputs(11270) <= a;
    outputs(11271) <= a xor b;
    outputs(11272) <= not (a xor b);
    outputs(11273) <= a and b;
    outputs(11274) <= not (a or b);
    outputs(11275) <= not (a or b);
    outputs(11276) <= b;
    outputs(11277) <= not a;
    outputs(11278) <= not b;
    outputs(11279) <= b and not a;
    outputs(11280) <= not b or a;
    outputs(11281) <= not b;
    outputs(11282) <= not (a xor b);
    outputs(11283) <= not (a xor b);
    outputs(11284) <= not a or b;
    outputs(11285) <= not a;
    outputs(11286) <= not a or b;
    outputs(11287) <= not b;
    outputs(11288) <= a xor b;
    outputs(11289) <= a xor b;
    outputs(11290) <= not a;
    outputs(11291) <= a xor b;
    outputs(11292) <= a xor b;
    outputs(11293) <= a xor b;
    outputs(11294) <= not (a xor b);
    outputs(11295) <= not b;
    outputs(11296) <= not (a xor b);
    outputs(11297) <= b;
    outputs(11298) <= a xor b;
    outputs(11299) <= a xor b;
    outputs(11300) <= a;
    outputs(11301) <= not (a xor b);
    outputs(11302) <= a;
    outputs(11303) <= a and b;
    outputs(11304) <= not (a and b);
    outputs(11305) <= a and not b;
    outputs(11306) <= a;
    outputs(11307) <= a xor b;
    outputs(11308) <= a and b;
    outputs(11309) <= b;
    outputs(11310) <= not a;
    outputs(11311) <= a;
    outputs(11312) <= not (a and b);
    outputs(11313) <= a xor b;
    outputs(11314) <= not a;
    outputs(11315) <= not b;
    outputs(11316) <= a and b;
    outputs(11317) <= not (a xor b);
    outputs(11318) <= not (a and b);
    outputs(11319) <= a;
    outputs(11320) <= not (a xor b);
    outputs(11321) <= a and not b;
    outputs(11322) <= a xor b;
    outputs(11323) <= not a;
    outputs(11324) <= a and not b;
    outputs(11325) <= not (a xor b);
    outputs(11326) <= a xor b;
    outputs(11327) <= not (a or b);
    outputs(11328) <= a xor b;
    outputs(11329) <= not (a xor b);
    outputs(11330) <= a xor b;
    outputs(11331) <= not (a and b);
    outputs(11332) <= not a;
    outputs(11333) <= a or b;
    outputs(11334) <= not a;
    outputs(11335) <= not (a xor b);
    outputs(11336) <= a xor b;
    outputs(11337) <= a xor b;
    outputs(11338) <= b and not a;
    outputs(11339) <= not (a xor b);
    outputs(11340) <= b;
    outputs(11341) <= not b;
    outputs(11342) <= not a;
    outputs(11343) <= a or b;
    outputs(11344) <= b and not a;
    outputs(11345) <= b;
    outputs(11346) <= b and not a;
    outputs(11347) <= a xor b;
    outputs(11348) <= not (a xor b);
    outputs(11349) <= a xor b;
    outputs(11350) <= not (a xor b);
    outputs(11351) <= not (a xor b);
    outputs(11352) <= b;
    outputs(11353) <= not (a xor b);
    outputs(11354) <= not a or b;
    outputs(11355) <= a;
    outputs(11356) <= b;
    outputs(11357) <= a;
    outputs(11358) <= not (a xor b);
    outputs(11359) <= not (a xor b);
    outputs(11360) <= a;
    outputs(11361) <= b;
    outputs(11362) <= b;
    outputs(11363) <= not a;
    outputs(11364) <= a xor b;
    outputs(11365) <= b;
    outputs(11366) <= not (a xor b);
    outputs(11367) <= b;
    outputs(11368) <= not b;
    outputs(11369) <= not b;
    outputs(11370) <= a;
    outputs(11371) <= not (a xor b);
    outputs(11372) <= a;
    outputs(11373) <= a or b;
    outputs(11374) <= a and b;
    outputs(11375) <= not b;
    outputs(11376) <= not (a and b);
    outputs(11377) <= b;
    outputs(11378) <= a;
    outputs(11379) <= a;
    outputs(11380) <= not b;
    outputs(11381) <= not b;
    outputs(11382) <= a xor b;
    outputs(11383) <= not a;
    outputs(11384) <= b;
    outputs(11385) <= a;
    outputs(11386) <= a and b;
    outputs(11387) <= not a;
    outputs(11388) <= not (a and b);
    outputs(11389) <= a;
    outputs(11390) <= b and not a;
    outputs(11391) <= b and not a;
    outputs(11392) <= not b;
    outputs(11393) <= not a;
    outputs(11394) <= a xor b;
    outputs(11395) <= a or b;
    outputs(11396) <= not (a xor b);
    outputs(11397) <= not a or b;
    outputs(11398) <= a and not b;
    outputs(11399) <= a xor b;
    outputs(11400) <= not a or b;
    outputs(11401) <= not (a or b);
    outputs(11402) <= b and not a;
    outputs(11403) <= not (a xor b);
    outputs(11404) <= a or b;
    outputs(11405) <= not b;
    outputs(11406) <= a and not b;
    outputs(11407) <= a xor b;
    outputs(11408) <= a;
    outputs(11409) <= a xor b;
    outputs(11410) <= a xor b;
    outputs(11411) <= not a;
    outputs(11412) <= b and not a;
    outputs(11413) <= not (a xor b);
    outputs(11414) <= not (a or b);
    outputs(11415) <= not b;
    outputs(11416) <= a or b;
    outputs(11417) <= b;
    outputs(11418) <= a xor b;
    outputs(11419) <= a;
    outputs(11420) <= a xor b;
    outputs(11421) <= a xor b;
    outputs(11422) <= a xor b;
    outputs(11423) <= not b;
    outputs(11424) <= not (a xor b);
    outputs(11425) <= not b;
    outputs(11426) <= not (a xor b);
    outputs(11427) <= b and not a;
    outputs(11428) <= not (a and b);
    outputs(11429) <= a;
    outputs(11430) <= a xor b;
    outputs(11431) <= a xor b;
    outputs(11432) <= not (a xor b);
    outputs(11433) <= not b;
    outputs(11434) <= b and not a;
    outputs(11435) <= a or b;
    outputs(11436) <= a xor b;
    outputs(11437) <= not (a xor b);
    outputs(11438) <= not (a xor b);
    outputs(11439) <= a xor b;
    outputs(11440) <= a or b;
    outputs(11441) <= not (a xor b);
    outputs(11442) <= a and b;
    outputs(11443) <= b;
    outputs(11444) <= not a or b;
    outputs(11445) <= not (a xor b);
    outputs(11446) <= not b;
    outputs(11447) <= not (a xor b);
    outputs(11448) <= not (a or b);
    outputs(11449) <= not a;
    outputs(11450) <= not a;
    outputs(11451) <= not (a and b);
    outputs(11452) <= not b;
    outputs(11453) <= a and b;
    outputs(11454) <= b;
    outputs(11455) <= not (a or b);
    outputs(11456) <= b;
    outputs(11457) <= b and not a;
    outputs(11458) <= a or b;
    outputs(11459) <= a xor b;
    outputs(11460) <= a or b;
    outputs(11461) <= a;
    outputs(11462) <= not (a or b);
    outputs(11463) <= a xor b;
    outputs(11464) <= not (a or b);
    outputs(11465) <= a xor b;
    outputs(11466) <= a xor b;
    outputs(11467) <= a;
    outputs(11468) <= not b;
    outputs(11469) <= not (a and b);
    outputs(11470) <= a xor b;
    outputs(11471) <= not a;
    outputs(11472) <= a xor b;
    outputs(11473) <= a xor b;
    outputs(11474) <= b;
    outputs(11475) <= a or b;
    outputs(11476) <= not (a and b);
    outputs(11477) <= not (a xor b);
    outputs(11478) <= not a;
    outputs(11479) <= a xor b;
    outputs(11480) <= not (a and b);
    outputs(11481) <= not a or b;
    outputs(11482) <= a and b;
    outputs(11483) <= a and not b;
    outputs(11484) <= not (a xor b);
    outputs(11485) <= b;
    outputs(11486) <= a;
    outputs(11487) <= not a or b;
    outputs(11488) <= a and not b;
    outputs(11489) <= not a or b;
    outputs(11490) <= a xor b;
    outputs(11491) <= not (a xor b);
    outputs(11492) <= not a;
    outputs(11493) <= b;
    outputs(11494) <= b;
    outputs(11495) <= not (a and b);
    outputs(11496) <= a xor b;
    outputs(11497) <= b;
    outputs(11498) <= not a or b;
    outputs(11499) <= b;
    outputs(11500) <= a xor b;
    outputs(11501) <= a xor b;
    outputs(11502) <= a;
    outputs(11503) <= b;
    outputs(11504) <= a;
    outputs(11505) <= a xor b;
    outputs(11506) <= not b;
    outputs(11507) <= b and not a;
    outputs(11508) <= not (a xor b);
    outputs(11509) <= a xor b;
    outputs(11510) <= not (a xor b);
    outputs(11511) <= b;
    outputs(11512) <= not a or b;
    outputs(11513) <= not b;
    outputs(11514) <= a xor b;
    outputs(11515) <= not (a xor b);
    outputs(11516) <= not (a or b);
    outputs(11517) <= not a;
    outputs(11518) <= not a;
    outputs(11519) <= not a or b;
    outputs(11520) <= not b;
    outputs(11521) <= not a or b;
    outputs(11522) <= not (a xor b);
    outputs(11523) <= a and not b;
    outputs(11524) <= not b;
    outputs(11525) <= not (a xor b);
    outputs(11526) <= b and not a;
    outputs(11527) <= not (a xor b);
    outputs(11528) <= a and b;
    outputs(11529) <= a xor b;
    outputs(11530) <= not (a xor b);
    outputs(11531) <= a and b;
    outputs(11532) <= not (a and b);
    outputs(11533) <= b;
    outputs(11534) <= not b;
    outputs(11535) <= not b;
    outputs(11536) <= not a;
    outputs(11537) <= not b;
    outputs(11538) <= b and not a;
    outputs(11539) <= a and b;
    outputs(11540) <= not (a or b);
    outputs(11541) <= b;
    outputs(11542) <= not a;
    outputs(11543) <= b;
    outputs(11544) <= a xor b;
    outputs(11545) <= not (a xor b);
    outputs(11546) <= b;
    outputs(11547) <= a;
    outputs(11548) <= not b;
    outputs(11549) <= not b or a;
    outputs(11550) <= b;
    outputs(11551) <= a and not b;
    outputs(11552) <= a xor b;
    outputs(11553) <= b;
    outputs(11554) <= not b;
    outputs(11555) <= a;
    outputs(11556) <= not (a xor b);
    outputs(11557) <= b;
    outputs(11558) <= b;
    outputs(11559) <= a;
    outputs(11560) <= not b or a;
    outputs(11561) <= not (a xor b);
    outputs(11562) <= b;
    outputs(11563) <= not (a xor b);
    outputs(11564) <= b;
    outputs(11565) <= not a;
    outputs(11566) <= a and not b;
    outputs(11567) <= b and not a;
    outputs(11568) <= a;
    outputs(11569) <= a or b;
    outputs(11570) <= not b;
    outputs(11571) <= a;
    outputs(11572) <= a xor b;
    outputs(11573) <= a and not b;
    outputs(11574) <= a and not b;
    outputs(11575) <= a and b;
    outputs(11576) <= b and not a;
    outputs(11577) <= not (a or b);
    outputs(11578) <= a and b;
    outputs(11579) <= a xor b;
    outputs(11580) <= not (a xor b);
    outputs(11581) <= not b;
    outputs(11582) <= not a;
    outputs(11583) <= a xor b;
    outputs(11584) <= not (a xor b);
    outputs(11585) <= a;
    outputs(11586) <= a xor b;
    outputs(11587) <= a;
    outputs(11588) <= a xor b;
    outputs(11589) <= a and not b;
    outputs(11590) <= not b;
    outputs(11591) <= a or b;
    outputs(11592) <= not (a xor b);
    outputs(11593) <= not (a xor b);
    outputs(11594) <= not (a xor b);
    outputs(11595) <= not (a xor b);
    outputs(11596) <= b and not a;
    outputs(11597) <= a and b;
    outputs(11598) <= not (a and b);
    outputs(11599) <= not (a and b);
    outputs(11600) <= not b;
    outputs(11601) <= not (a and b);
    outputs(11602) <= a xor b;
    outputs(11603) <= not (a and b);
    outputs(11604) <= a;
    outputs(11605) <= not (a xor b);
    outputs(11606) <= not a or b;
    outputs(11607) <= not b or a;
    outputs(11608) <= not (a xor b);
    outputs(11609) <= a and not b;
    outputs(11610) <= a;
    outputs(11611) <= not (a xor b);
    outputs(11612) <= a or b;
    outputs(11613) <= a;
    outputs(11614) <= a;
    outputs(11615) <= not (a xor b);
    outputs(11616) <= a;
    outputs(11617) <= not (a xor b);
    outputs(11618) <= a xor b;
    outputs(11619) <= not b;
    outputs(11620) <= b;
    outputs(11621) <= not (a xor b);
    outputs(11622) <= not (a xor b);
    outputs(11623) <= a xor b;
    outputs(11624) <= a xor b;
    outputs(11625) <= not (a xor b);
    outputs(11626) <= not b;
    outputs(11627) <= not (a xor b);
    outputs(11628) <= not b;
    outputs(11629) <= b and not a;
    outputs(11630) <= a xor b;
    outputs(11631) <= a and b;
    outputs(11632) <= b and not a;
    outputs(11633) <= b;
    outputs(11634) <= a and b;
    outputs(11635) <= not (a xor b);
    outputs(11636) <= b;
    outputs(11637) <= a and not b;
    outputs(11638) <= not (a xor b);
    outputs(11639) <= a xor b;
    outputs(11640) <= a xor b;
    outputs(11641) <= not (a xor b);
    outputs(11642) <= b;
    outputs(11643) <= a or b;
    outputs(11644) <= not (a or b);
    outputs(11645) <= not a;
    outputs(11646) <= a and not b;
    outputs(11647) <= a;
    outputs(11648) <= a and not b;
    outputs(11649) <= not b;
    outputs(11650) <= not b;
    outputs(11651) <= not b or a;
    outputs(11652) <= a and b;
    outputs(11653) <= b;
    outputs(11654) <= a;
    outputs(11655) <= not a;
    outputs(11656) <= not a or b;
    outputs(11657) <= b and not a;
    outputs(11658) <= a;
    outputs(11659) <= b;
    outputs(11660) <= a and b;
    outputs(11661) <= not (a xor b);
    outputs(11662) <= not (a xor b);
    outputs(11663) <= a xor b;
    outputs(11664) <= not (a xor b);
    outputs(11665) <= not (a and b);
    outputs(11666) <= a xor b;
    outputs(11667) <= not b;
    outputs(11668) <= not b;
    outputs(11669) <= b;
    outputs(11670) <= not (a xor b);
    outputs(11671) <= a;
    outputs(11672) <= not (a xor b);
    outputs(11673) <= not a;
    outputs(11674) <= b;
    outputs(11675) <= a xor b;
    outputs(11676) <= not (a or b);
    outputs(11677) <= a xor b;
    outputs(11678) <= b and not a;
    outputs(11679) <= not (a or b);
    outputs(11680) <= not (a or b);
    outputs(11681) <= not (a or b);
    outputs(11682) <= b;
    outputs(11683) <= not b;
    outputs(11684) <= a;
    outputs(11685) <= not (a and b);
    outputs(11686) <= a and b;
    outputs(11687) <= not (a xor b);
    outputs(11688) <= not (a xor b);
    outputs(11689) <= a xor b;
    outputs(11690) <= a;
    outputs(11691) <= a and not b;
    outputs(11692) <= b;
    outputs(11693) <= b and not a;
    outputs(11694) <= not a;
    outputs(11695) <= not (a xor b);
    outputs(11696) <= not a;
    outputs(11697) <= a and not b;
    outputs(11698) <= not a;
    outputs(11699) <= a xor b;
    outputs(11700) <= a and not b;
    outputs(11701) <= not a;
    outputs(11702) <= not (a xor b);
    outputs(11703) <= not b or a;
    outputs(11704) <= a xor b;
    outputs(11705) <= a xor b;
    outputs(11706) <= not (a xor b);
    outputs(11707) <= not (a xor b);
    outputs(11708) <= not a;
    outputs(11709) <= not b;
    outputs(11710) <= not b;
    outputs(11711) <= not b;
    outputs(11712) <= not a or b;
    outputs(11713) <= not a;
    outputs(11714) <= not b or a;
    outputs(11715) <= not b;
    outputs(11716) <= not b;
    outputs(11717) <= a;
    outputs(11718) <= a and not b;
    outputs(11719) <= not a or b;
    outputs(11720) <= a and b;
    outputs(11721) <= b;
    outputs(11722) <= not a;
    outputs(11723) <= b;
    outputs(11724) <= a or b;
    outputs(11725) <= b;
    outputs(11726) <= not (a xor b);
    outputs(11727) <= not a;
    outputs(11728) <= not (a xor b);
    outputs(11729) <= not a;
    outputs(11730) <= b;
    outputs(11731) <= a xor b;
    outputs(11732) <= a xor b;
    outputs(11733) <= a and b;
    outputs(11734) <= a xor b;
    outputs(11735) <= a xor b;
    outputs(11736) <= a;
    outputs(11737) <= not (a and b);
    outputs(11738) <= b and not a;
    outputs(11739) <= a xor b;
    outputs(11740) <= a xor b;
    outputs(11741) <= not (a xor b);
    outputs(11742) <= a xor b;
    outputs(11743) <= not a;
    outputs(11744) <= not a;
    outputs(11745) <= b;
    outputs(11746) <= a;
    outputs(11747) <= a and b;
    outputs(11748) <= not (a and b);
    outputs(11749) <= a;
    outputs(11750) <= not a;
    outputs(11751) <= a xor b;
    outputs(11752) <= a;
    outputs(11753) <= b;
    outputs(11754) <= not (a xor b);
    outputs(11755) <= 1'b0;
    outputs(11756) <= not (a xor b);
    outputs(11757) <= a xor b;
    outputs(11758) <= a;
    outputs(11759) <= a;
    outputs(11760) <= not a;
    outputs(11761) <= a xor b;
    outputs(11762) <= not a;
    outputs(11763) <= not a;
    outputs(11764) <= a xor b;
    outputs(11765) <= not b;
    outputs(11766) <= not b;
    outputs(11767) <= not a or b;
    outputs(11768) <= b;
    outputs(11769) <= a and not b;
    outputs(11770) <= a;
    outputs(11771) <= b;
    outputs(11772) <= not (a xor b);
    outputs(11773) <= a xor b;
    outputs(11774) <= a xor b;
    outputs(11775) <= not b;
    outputs(11776) <= a xor b;
    outputs(11777) <= not (a xor b);
    outputs(11778) <= b and not a;
    outputs(11779) <= b and not a;
    outputs(11780) <= not a or b;
    outputs(11781) <= not (a xor b);
    outputs(11782) <= a xor b;
    outputs(11783) <= not b;
    outputs(11784) <= a;
    outputs(11785) <= not (a xor b);
    outputs(11786) <= b and not a;
    outputs(11787) <= a or b;
    outputs(11788) <= a xor b;
    outputs(11789) <= not (a xor b);
    outputs(11790) <= a xor b;
    outputs(11791) <= a;
    outputs(11792) <= not b;
    outputs(11793) <= a xor b;
    outputs(11794) <= not (a xor b);
    outputs(11795) <= not (a xor b);
    outputs(11796) <= a xor b;
    outputs(11797) <= not (a or b);
    outputs(11798) <= not a;
    outputs(11799) <= a;
    outputs(11800) <= a xor b;
    outputs(11801) <= b;
    outputs(11802) <= a xor b;
    outputs(11803) <= a or b;
    outputs(11804) <= a xor b;
    outputs(11805) <= not b;
    outputs(11806) <= not (a or b);
    outputs(11807) <= not a;
    outputs(11808) <= b;
    outputs(11809) <= not a;
    outputs(11810) <= not (a or b);
    outputs(11811) <= b and not a;
    outputs(11812) <= a xor b;
    outputs(11813) <= not b;
    outputs(11814) <= not a;
    outputs(11815) <= not b;
    outputs(11816) <= not (a or b);
    outputs(11817) <= not b or a;
    outputs(11818) <= b;
    outputs(11819) <= b;
    outputs(11820) <= not (a xor b);
    outputs(11821) <= not (a xor b);
    outputs(11822) <= a xor b;
    outputs(11823) <= not (a xor b);
    outputs(11824) <= not (a xor b);
    outputs(11825) <= b and not a;
    outputs(11826) <= b and not a;
    outputs(11827) <= not b or a;
    outputs(11828) <= not (a xor b);
    outputs(11829) <= a and b;
    outputs(11830) <= not (a xor b);
    outputs(11831) <= a xor b;
    outputs(11832) <= a and not b;
    outputs(11833) <= a xor b;
    outputs(11834) <= not b;
    outputs(11835) <= not (a xor b);
    outputs(11836) <= not (a xor b);
    outputs(11837) <= not a;
    outputs(11838) <= not b;
    outputs(11839) <= a xor b;
    outputs(11840) <= not b or a;
    outputs(11841) <= not a or b;
    outputs(11842) <= a xor b;
    outputs(11843) <= not a or b;
    outputs(11844) <= a xor b;
    outputs(11845) <= a and b;
    outputs(11846) <= b and not a;
    outputs(11847) <= not (a or b);
    outputs(11848) <= a;
    outputs(11849) <= not a;
    outputs(11850) <= not (a xor b);
    outputs(11851) <= a xor b;
    outputs(11852) <= not b;
    outputs(11853) <= not (a and b);
    outputs(11854) <= a and not b;
    outputs(11855) <= not (a and b);
    outputs(11856) <= a xor b;
    outputs(11857) <= not b;
    outputs(11858) <= not b;
    outputs(11859) <= b;
    outputs(11860) <= a and not b;
    outputs(11861) <= not (a xor b);
    outputs(11862) <= b and not a;
    outputs(11863) <= b and not a;
    outputs(11864) <= not b;
    outputs(11865) <= b and not a;
    outputs(11866) <= not b;
    outputs(11867) <= not b or a;
    outputs(11868) <= not (a or b);
    outputs(11869) <= a or b;
    outputs(11870) <= a;
    outputs(11871) <= not a;
    outputs(11872) <= b;
    outputs(11873) <= b;
    outputs(11874) <= not (a xor b);
    outputs(11875) <= not (a xor b);
    outputs(11876) <= not b or a;
    outputs(11877) <= not (a xor b);
    outputs(11878) <= not (a xor b);
    outputs(11879) <= a and b;
    outputs(11880) <= not b or a;
    outputs(11881) <= not (a xor b);
    outputs(11882) <= a and b;
    outputs(11883) <= not b;
    outputs(11884) <= a xor b;
    outputs(11885) <= a and not b;
    outputs(11886) <= not a;
    outputs(11887) <= a xor b;
    outputs(11888) <= a xor b;
    outputs(11889) <= not (a xor b);
    outputs(11890) <= not (a xor b);
    outputs(11891) <= not a;
    outputs(11892) <= a xor b;
    outputs(11893) <= not b;
    outputs(11894) <= not b;
    outputs(11895) <= not a;
    outputs(11896) <= not (a xor b);
    outputs(11897) <= not (a xor b);
    outputs(11898) <= b;
    outputs(11899) <= not b or a;
    outputs(11900) <= a xor b;
    outputs(11901) <= not a;
    outputs(11902) <= not a or b;
    outputs(11903) <= b;
    outputs(11904) <= a;
    outputs(11905) <= not (a xor b);
    outputs(11906) <= a xor b;
    outputs(11907) <= not (a xor b);
    outputs(11908) <= not b;
    outputs(11909) <= not a;
    outputs(11910) <= a xor b;
    outputs(11911) <= not a;
    outputs(11912) <= a xor b;
    outputs(11913) <= a xor b;
    outputs(11914) <= a and b;
    outputs(11915) <= not a;
    outputs(11916) <= not (a xor b);
    outputs(11917) <= a;
    outputs(11918) <= not a;
    outputs(11919) <= b and not a;
    outputs(11920) <= not (a xor b);
    outputs(11921) <= a and b;
    outputs(11922) <= not b;
    outputs(11923) <= a xor b;
    outputs(11924) <= not (a or b);
    outputs(11925) <= not (a xor b);
    outputs(11926) <= a and b;
    outputs(11927) <= a xor b;
    outputs(11928) <= b;
    outputs(11929) <= a xor b;
    outputs(11930) <= a;
    outputs(11931) <= not (a and b);
    outputs(11932) <= a xor b;
    outputs(11933) <= not (a xor b);
    outputs(11934) <= b and not a;
    outputs(11935) <= not (a xor b);
    outputs(11936) <= b;
    outputs(11937) <= not (a xor b);
    outputs(11938) <= not (a xor b);
    outputs(11939) <= not (a and b);
    outputs(11940) <= not b;
    outputs(11941) <= not (a xor b);
    outputs(11942) <= a;
    outputs(11943) <= not b or a;
    outputs(11944) <= not b or a;
    outputs(11945) <= b;
    outputs(11946) <= a and b;
    outputs(11947) <= a xor b;
    outputs(11948) <= not a;
    outputs(11949) <= not (a xor b);
    outputs(11950) <= not (a xor b);
    outputs(11951) <= b;
    outputs(11952) <= a and b;
    outputs(11953) <= not b or a;
    outputs(11954) <= a xor b;
    outputs(11955) <= a and b;
    outputs(11956) <= b and not a;
    outputs(11957) <= not a;
    outputs(11958) <= a xor b;
    outputs(11959) <= not (a xor b);
    outputs(11960) <= not (a xor b);
    outputs(11961) <= not a;
    outputs(11962) <= a xor b;
    outputs(11963) <= not (a xor b);
    outputs(11964) <= not a or b;
    outputs(11965) <= not (a and b);
    outputs(11966) <= not b or a;
    outputs(11967) <= a xor b;
    outputs(11968) <= a or b;
    outputs(11969) <= not a or b;
    outputs(11970) <= a and not b;
    outputs(11971) <= a xor b;
    outputs(11972) <= not (a xor b);
    outputs(11973) <= not a;
    outputs(11974) <= a xor b;
    outputs(11975) <= not b;
    outputs(11976) <= b and not a;
    outputs(11977) <= not b;
    outputs(11978) <= b and not a;
    outputs(11979) <= not b;
    outputs(11980) <= b;
    outputs(11981) <= a and b;
    outputs(11982) <= b;
    outputs(11983) <= a and not b;
    outputs(11984) <= not (a xor b);
    outputs(11985) <= not a;
    outputs(11986) <= not (a or b);
    outputs(11987) <= a;
    outputs(11988) <= not (a xor b);
    outputs(11989) <= not b;
    outputs(11990) <= a and not b;
    outputs(11991) <= a and b;
    outputs(11992) <= a;
    outputs(11993) <= a and not b;
    outputs(11994) <= a;
    outputs(11995) <= a xor b;
    outputs(11996) <= not (a xor b);
    outputs(11997) <= a and b;
    outputs(11998) <= a and b;
    outputs(11999) <= b;
    outputs(12000) <= b and not a;
    outputs(12001) <= not a;
    outputs(12002) <= b;
    outputs(12003) <= not (a xor b);
    outputs(12004) <= not (a xor b);
    outputs(12005) <= b and not a;
    outputs(12006) <= not b;
    outputs(12007) <= not (a xor b);
    outputs(12008) <= a or b;
    outputs(12009) <= not (a xor b);
    outputs(12010) <= not (a xor b);
    outputs(12011) <= not (a xor b);
    outputs(12012) <= not (a xor b);
    outputs(12013) <= a and b;
    outputs(12014) <= b;
    outputs(12015) <= not (a xor b);
    outputs(12016) <= a;
    outputs(12017) <= a;
    outputs(12018) <= b;
    outputs(12019) <= not (a xor b);
    outputs(12020) <= a;
    outputs(12021) <= not (a xor b);
    outputs(12022) <= a xor b;
    outputs(12023) <= a xor b;
    outputs(12024) <= a;
    outputs(12025) <= a;
    outputs(12026) <= not (a xor b);
    outputs(12027) <= not a;
    outputs(12028) <= not b or a;
    outputs(12029) <= b;
    outputs(12030) <= a xor b;
    outputs(12031) <= a and b;
    outputs(12032) <= a xor b;
    outputs(12033) <= not b;
    outputs(12034) <= a xor b;
    outputs(12035) <= b and not a;
    outputs(12036) <= a;
    outputs(12037) <= not (a xor b);
    outputs(12038) <= b;
    outputs(12039) <= not a;
    outputs(12040) <= a xor b;
    outputs(12041) <= a;
    outputs(12042) <= not (a and b);
    outputs(12043) <= a xor b;
    outputs(12044) <= b;
    outputs(12045) <= not b;
    outputs(12046) <= b;
    outputs(12047) <= not a or b;
    outputs(12048) <= b;
    outputs(12049) <= b and not a;
    outputs(12050) <= a;
    outputs(12051) <= not (a and b);
    outputs(12052) <= not (a xor b);
    outputs(12053) <= not a;
    outputs(12054) <= not (a xor b);
    outputs(12055) <= a xor b;
    outputs(12056) <= a and not b;
    outputs(12057) <= not a;
    outputs(12058) <= a xor b;
    outputs(12059) <= b and not a;
    outputs(12060) <= not (a xor b);
    outputs(12061) <= not (a xor b);
    outputs(12062) <= not a or b;
    outputs(12063) <= a xor b;
    outputs(12064) <= not (a or b);
    outputs(12065) <= not (a xor b);
    outputs(12066) <= a xor b;
    outputs(12067) <= a xor b;
    outputs(12068) <= a;
    outputs(12069) <= not b;
    outputs(12070) <= a xor b;
    outputs(12071) <= a xor b;
    outputs(12072) <= a and b;
    outputs(12073) <= not (a and b);
    outputs(12074) <= not (a xor b);
    outputs(12075) <= not (a xor b);
    outputs(12076) <= b and not a;
    outputs(12077) <= a xor b;
    outputs(12078) <= not (a xor b);
    outputs(12079) <= not a or b;
    outputs(12080) <= not b;
    outputs(12081) <= not a or b;
    outputs(12082) <= a and b;
    outputs(12083) <= not (a xor b);
    outputs(12084) <= a xor b;
    outputs(12085) <= a xor b;
    outputs(12086) <= a;
    outputs(12087) <= not (a xor b);
    outputs(12088) <= not b;
    outputs(12089) <= b;
    outputs(12090) <= not (a xor b);
    outputs(12091) <= not a;
    outputs(12092) <= not (a xor b);
    outputs(12093) <= b and not a;
    outputs(12094) <= a xor b;
    outputs(12095) <= not (a xor b);
    outputs(12096) <= a and not b;
    outputs(12097) <= b;
    outputs(12098) <= b;
    outputs(12099) <= not a;
    outputs(12100) <= not b or a;
    outputs(12101) <= b;
    outputs(12102) <= not a;
    outputs(12103) <= not (a xor b);
    outputs(12104) <= a and b;
    outputs(12105) <= a xor b;
    outputs(12106) <= a and not b;
    outputs(12107) <= not b;
    outputs(12108) <= not (a xor b);
    outputs(12109) <= not (a or b);
    outputs(12110) <= not b;
    outputs(12111) <= a xor b;
    outputs(12112) <= not (a xor b);
    outputs(12113) <= a xor b;
    outputs(12114) <= b;
    outputs(12115) <= not a;
    outputs(12116) <= a and b;
    outputs(12117) <= a;
    outputs(12118) <= not (a or b);
    outputs(12119) <= b;
    outputs(12120) <= not b;
    outputs(12121) <= not b;
    outputs(12122) <= a and not b;
    outputs(12123) <= not (a xor b);
    outputs(12124) <= not (a xor b);
    outputs(12125) <= not b or a;
    outputs(12126) <= b;
    outputs(12127) <= a xor b;
    outputs(12128) <= not b;
    outputs(12129) <= a and b;
    outputs(12130) <= a xor b;
    outputs(12131) <= not b or a;
    outputs(12132) <= not a or b;
    outputs(12133) <= b;
    outputs(12134) <= a and b;
    outputs(12135) <= not (a xor b);
    outputs(12136) <= not (a xor b);
    outputs(12137) <= a or b;
    outputs(12138) <= not a;
    outputs(12139) <= b;
    outputs(12140) <= not (a and b);
    outputs(12141) <= not (a and b);
    outputs(12142) <= not (a or b);
    outputs(12143) <= a and not b;
    outputs(12144) <= b;
    outputs(12145) <= b and not a;
    outputs(12146) <= not (a or b);
    outputs(12147) <= not a;
    outputs(12148) <= a xor b;
    outputs(12149) <= not a;
    outputs(12150) <= not b;
    outputs(12151) <= b;
    outputs(12152) <= not (a xor b);
    outputs(12153) <= not (a or b);
    outputs(12154) <= a xor b;
    outputs(12155) <= not b;
    outputs(12156) <= a;
    outputs(12157) <= b;
    outputs(12158) <= b;
    outputs(12159) <= a;
    outputs(12160) <= a and b;
    outputs(12161) <= not b;
    outputs(12162) <= not b or a;
    outputs(12163) <= b;
    outputs(12164) <= a;
    outputs(12165) <= not (a xor b);
    outputs(12166) <= not a or b;
    outputs(12167) <= not b;
    outputs(12168) <= not b;
    outputs(12169) <= not (a or b);
    outputs(12170) <= not b;
    outputs(12171) <= not a;
    outputs(12172) <= a;
    outputs(12173) <= not (a xor b);
    outputs(12174) <= not (a xor b);
    outputs(12175) <= not (a xor b);
    outputs(12176) <= a and b;
    outputs(12177) <= b;
    outputs(12178) <= a;
    outputs(12179) <= a and not b;
    outputs(12180) <= not (a xor b);
    outputs(12181) <= a and not b;
    outputs(12182) <= a xor b;
    outputs(12183) <= b;
    outputs(12184) <= a xor b;
    outputs(12185) <= a;
    outputs(12186) <= not (a xor b);
    outputs(12187) <= a xor b;
    outputs(12188) <= a;
    outputs(12189) <= a and not b;
    outputs(12190) <= a or b;
    outputs(12191) <= a;
    outputs(12192) <= not b;
    outputs(12193) <= a xor b;
    outputs(12194) <= not (a xor b);
    outputs(12195) <= not b;
    outputs(12196) <= b;
    outputs(12197) <= not (a or b);
    outputs(12198) <= not (a xor b);
    outputs(12199) <= not (a xor b);
    outputs(12200) <= not (a xor b);
    outputs(12201) <= not (a or b);
    outputs(12202) <= a;
    outputs(12203) <= a xor b;
    outputs(12204) <= not (a xor b);
    outputs(12205) <= a xor b;
    outputs(12206) <= a xor b;
    outputs(12207) <= b and not a;
    outputs(12208) <= a xor b;
    outputs(12209) <= b and not a;
    outputs(12210) <= not (a xor b);
    outputs(12211) <= not (a or b);
    outputs(12212) <= not (a or b);
    outputs(12213) <= not (a xor b);
    outputs(12214) <= a xor b;
    outputs(12215) <= not b;
    outputs(12216) <= b and not a;
    outputs(12217) <= not b;
    outputs(12218) <= a xor b;
    outputs(12219) <= not b;
    outputs(12220) <= not a;
    outputs(12221) <= b and not a;
    outputs(12222) <= not (a or b);
    outputs(12223) <= a xor b;
    outputs(12224) <= a and not b;
    outputs(12225) <= a;
    outputs(12226) <= b;
    outputs(12227) <= not b;
    outputs(12228) <= not b;
    outputs(12229) <= a and not b;
    outputs(12230) <= not (a xor b);
    outputs(12231) <= a and b;
    outputs(12232) <= not a;
    outputs(12233) <= not b;
    outputs(12234) <= a xor b;
    outputs(12235) <= a xor b;
    outputs(12236) <= not (a or b);
    outputs(12237) <= not a;
    outputs(12238) <= not b;
    outputs(12239) <= a;
    outputs(12240) <= a and not b;
    outputs(12241) <= a xor b;
    outputs(12242) <= a xor b;
    outputs(12243) <= a xor b;
    outputs(12244) <= not (a or b);
    outputs(12245) <= b;
    outputs(12246) <= b and not a;
    outputs(12247) <= a xor b;
    outputs(12248) <= not (a xor b);
    outputs(12249) <= not (a xor b);
    outputs(12250) <= not a or b;
    outputs(12251) <= a xor b;
    outputs(12252) <= not (a or b);
    outputs(12253) <= b and not a;
    outputs(12254) <= not a or b;
    outputs(12255) <= not (a xor b);
    outputs(12256) <= not (a or b);
    outputs(12257) <= not a or b;
    outputs(12258) <= b and not a;
    outputs(12259) <= a xor b;
    outputs(12260) <= a xor b;
    outputs(12261) <= not (a xor b);
    outputs(12262) <= not a or b;
    outputs(12263) <= a and b;
    outputs(12264) <= b;
    outputs(12265) <= not (a or b);
    outputs(12266) <= not b or a;
    outputs(12267) <= a or b;
    outputs(12268) <= not (a xor b);
    outputs(12269) <= not (a xor b);
    outputs(12270) <= a and not b;
    outputs(12271) <= not a;
    outputs(12272) <= not b;
    outputs(12273) <= b;
    outputs(12274) <= not (a or b);
    outputs(12275) <= a and not b;
    outputs(12276) <= a or b;
    outputs(12277) <= not (a xor b);
    outputs(12278) <= not (a xor b);
    outputs(12279) <= not b;
    outputs(12280) <= not (a or b);
    outputs(12281) <= a xor b;
    outputs(12282) <= b and not a;
    outputs(12283) <= not b;
    outputs(12284) <= not a or b;
    outputs(12285) <= not b;
    outputs(12286) <= b;
    outputs(12287) <= a and b;
    outputs(12288) <= not (a xor b);
    outputs(12289) <= not a;
    outputs(12290) <= not (a xor b);
    outputs(12291) <= a xor b;
    outputs(12292) <= not a;
    outputs(12293) <= a xor b;
    outputs(12294) <= not b;
    outputs(12295) <= b;
    outputs(12296) <= a;
    outputs(12297) <= not a;
    outputs(12298) <= not a;
    outputs(12299) <= a;
    outputs(12300) <= not (a or b);
    outputs(12301) <= a xor b;
    outputs(12302) <= not (a or b);
    outputs(12303) <= a xor b;
    outputs(12304) <= a and not b;
    outputs(12305) <= not b;
    outputs(12306) <= a xor b;
    outputs(12307) <= not (a xor b);
    outputs(12308) <= not (a or b);
    outputs(12309) <= b and not a;
    outputs(12310) <= not b;
    outputs(12311) <= not (a xor b);
    outputs(12312) <= b;
    outputs(12313) <= a and not b;
    outputs(12314) <= not (a xor b);
    outputs(12315) <= a;
    outputs(12316) <= not a;
    outputs(12317) <= a xor b;
    outputs(12318) <= not (a xor b);
    outputs(12319) <= a and not b;
    outputs(12320) <= a;
    outputs(12321) <= not (a xor b);
    outputs(12322) <= a;
    outputs(12323) <= a;
    outputs(12324) <= not (a xor b);
    outputs(12325) <= not b;
    outputs(12326) <= a;
    outputs(12327) <= not b;
    outputs(12328) <= not a;
    outputs(12329) <= a xor b;
    outputs(12330) <= a and not b;
    outputs(12331) <= not b or a;
    outputs(12332) <= b;
    outputs(12333) <= b;
    outputs(12334) <= not a;
    outputs(12335) <= b;
    outputs(12336) <= not (a xor b);
    outputs(12337) <= not (a or b);
    outputs(12338) <= not a;
    outputs(12339) <= not (a and b);
    outputs(12340) <= not (a or b);
    outputs(12341) <= a xor b;
    outputs(12342) <= not (a xor b);
    outputs(12343) <= not (a xor b);
    outputs(12344) <= a xor b;
    outputs(12345) <= a and b;
    outputs(12346) <= not (a or b);
    outputs(12347) <= a;
    outputs(12348) <= not (a xor b);
    outputs(12349) <= not (a xor b);
    outputs(12350) <= not b;
    outputs(12351) <= not (a xor b);
    outputs(12352) <= b and not a;
    outputs(12353) <= b and not a;
    outputs(12354) <= b;
    outputs(12355) <= a;
    outputs(12356) <= a and not b;
    outputs(12357) <= a;
    outputs(12358) <= a xor b;
    outputs(12359) <= not a;
    outputs(12360) <= a xor b;
    outputs(12361) <= not (a xor b);
    outputs(12362) <= a xor b;
    outputs(12363) <= not (a xor b);
    outputs(12364) <= b and not a;
    outputs(12365) <= not (a or b);
    outputs(12366) <= not (a or b);
    outputs(12367) <= b;
    outputs(12368) <= not (a xor b);
    outputs(12369) <= b;
    outputs(12370) <= b and not a;
    outputs(12371) <= not (a xor b);
    outputs(12372) <= not b or a;
    outputs(12373) <= not b or a;
    outputs(12374) <= not (a or b);
    outputs(12375) <= b;
    outputs(12376) <= a xor b;
    outputs(12377) <= not (a xor b);
    outputs(12378) <= not (a xor b);
    outputs(12379) <= a xor b;
    outputs(12380) <= b;
    outputs(12381) <= b and not a;
    outputs(12382) <= a xor b;
    outputs(12383) <= not b or a;
    outputs(12384) <= a xor b;
    outputs(12385) <= a xor b;
    outputs(12386) <= not (a xor b);
    outputs(12387) <= not (a xor b);
    outputs(12388) <= not b;
    outputs(12389) <= a and not b;
    outputs(12390) <= a and b;
    outputs(12391) <= a and b;
    outputs(12392) <= b and not a;
    outputs(12393) <= b;
    outputs(12394) <= not a;
    outputs(12395) <= not a;
    outputs(12396) <= a xor b;
    outputs(12397) <= a and not b;
    outputs(12398) <= a;
    outputs(12399) <= a;
    outputs(12400) <= not b;
    outputs(12401) <= a;
    outputs(12402) <= a xor b;
    outputs(12403) <= a xor b;
    outputs(12404) <= b and not a;
    outputs(12405) <= not (a or b);
    outputs(12406) <= b;
    outputs(12407) <= a xor b;
    outputs(12408) <= a xor b;
    outputs(12409) <= a;
    outputs(12410) <= not (a or b);
    outputs(12411) <= not (a xor b);
    outputs(12412) <= a and not b;
    outputs(12413) <= 1'b0;
    outputs(12414) <= a and b;
    outputs(12415) <= a and b;
    outputs(12416) <= a;
    outputs(12417) <= not (a xor b);
    outputs(12418) <= not b or a;
    outputs(12419) <= not b;
    outputs(12420) <= a xor b;
    outputs(12421) <= a or b;
    outputs(12422) <= not b or a;
    outputs(12423) <= b;
    outputs(12424) <= not (a or b);
    outputs(12425) <= not (a xor b);
    outputs(12426) <= not (a xor b);
    outputs(12427) <= not (a xor b);
    outputs(12428) <= a xor b;
    outputs(12429) <= a xor b;
    outputs(12430) <= b;
    outputs(12431) <= a xor b;
    outputs(12432) <= not (a xor b);
    outputs(12433) <= b and not a;
    outputs(12434) <= not (a xor b);
    outputs(12435) <= a xor b;
    outputs(12436) <= not b;
    outputs(12437) <= a and b;
    outputs(12438) <= not b;
    outputs(12439) <= a xor b;
    outputs(12440) <= not (a xor b);
    outputs(12441) <= not a or b;
    outputs(12442) <= not (a xor b);
    outputs(12443) <= not (a and b);
    outputs(12444) <= not (a or b);
    outputs(12445) <= b;
    outputs(12446) <= not (a xor b);
    outputs(12447) <= a xor b;
    outputs(12448) <= a and b;
    outputs(12449) <= not a;
    outputs(12450) <= b;
    outputs(12451) <= not (a xor b);
    outputs(12452) <= b and not a;
    outputs(12453) <= not (a xor b);
    outputs(12454) <= b;
    outputs(12455) <= b and not a;
    outputs(12456) <= not a or b;
    outputs(12457) <= b;
    outputs(12458) <= b;
    outputs(12459) <= not (a xor b);
    outputs(12460) <= a and b;
    outputs(12461) <= not (a xor b);
    outputs(12462) <= a or b;
    outputs(12463) <= a and b;
    outputs(12464) <= not (a xor b);
    outputs(12465) <= not a;
    outputs(12466) <= a xor b;
    outputs(12467) <= not (a xor b);
    outputs(12468) <= b;
    outputs(12469) <= not b;
    outputs(12470) <= a xor b;
    outputs(12471) <= a xor b;
    outputs(12472) <= not a;
    outputs(12473) <= not (a xor b);
    outputs(12474) <= a xor b;
    outputs(12475) <= a;
    outputs(12476) <= not (a and b);
    outputs(12477) <= a and b;
    outputs(12478) <= a xor b;
    outputs(12479) <= not (a xor b);
    outputs(12480) <= a xor b;
    outputs(12481) <= not a or b;
    outputs(12482) <= b and not a;
    outputs(12483) <= b and not a;
    outputs(12484) <= not b;
    outputs(12485) <= b and not a;
    outputs(12486) <= not (a xor b);
    outputs(12487) <= a or b;
    outputs(12488) <= not (a xor b);
    outputs(12489) <= a;
    outputs(12490) <= a xor b;
    outputs(12491) <= a;
    outputs(12492) <= not (a xor b);
    outputs(12493) <= a;
    outputs(12494) <= b;
    outputs(12495) <= not b;
    outputs(12496) <= b and not a;
    outputs(12497) <= not (a xor b);
    outputs(12498) <= b;
    outputs(12499) <= not a;
    outputs(12500) <= not b;
    outputs(12501) <= b and not a;
    outputs(12502) <= a xor b;
    outputs(12503) <= b and not a;
    outputs(12504) <= not (a xor b);
    outputs(12505) <= a xor b;
    outputs(12506) <= b and not a;
    outputs(12507) <= not b;
    outputs(12508) <= not (a xor b);
    outputs(12509) <= a and b;
    outputs(12510) <= a and b;
    outputs(12511) <= a and b;
    outputs(12512) <= not (a or b);
    outputs(12513) <= a xor b;
    outputs(12514) <= a xor b;
    outputs(12515) <= not (a or b);
    outputs(12516) <= not (a xor b);
    outputs(12517) <= not (a xor b);
    outputs(12518) <= b;
    outputs(12519) <= a xor b;
    outputs(12520) <= b;
    outputs(12521) <= not (a xor b);
    outputs(12522) <= a xor b;
    outputs(12523) <= a xor b;
    outputs(12524) <= a xor b;
    outputs(12525) <= b;
    outputs(12526) <= a and b;
    outputs(12527) <= a;
    outputs(12528) <= a;
    outputs(12529) <= a xor b;
    outputs(12530) <= a xor b;
    outputs(12531) <= b;
    outputs(12532) <= not (a xor b);
    outputs(12533) <= not b;
    outputs(12534) <= not b or a;
    outputs(12535) <= a xor b;
    outputs(12536) <= not a;
    outputs(12537) <= not (a xor b);
    outputs(12538) <= a or b;
    outputs(12539) <= b;
    outputs(12540) <= not (a xor b);
    outputs(12541) <= a;
    outputs(12542) <= a or b;
    outputs(12543) <= a and b;
    outputs(12544) <= a;
    outputs(12545) <= a xor b;
    outputs(12546) <= a xor b;
    outputs(12547) <= not (a xor b);
    outputs(12548) <= a xor b;
    outputs(12549) <= a xor b;
    outputs(12550) <= a;
    outputs(12551) <= a xor b;
    outputs(12552) <= a xor b;
    outputs(12553) <= b;
    outputs(12554) <= not b;
    outputs(12555) <= b;
    outputs(12556) <= b and not a;
    outputs(12557) <= a;
    outputs(12558) <= not (a xor b);
    outputs(12559) <= not a;
    outputs(12560) <= not (a xor b);
    outputs(12561) <= not (a xor b);
    outputs(12562) <= not (a xor b);
    outputs(12563) <= not (a xor b);
    outputs(12564) <= b and not a;
    outputs(12565) <= a and not b;
    outputs(12566) <= a or b;
    outputs(12567) <= a and not b;
    outputs(12568) <= b;
    outputs(12569) <= a xor b;
    outputs(12570) <= not a or b;
    outputs(12571) <= a xor b;
    outputs(12572) <= b;
    outputs(12573) <= a and not b;
    outputs(12574) <= not b or a;
    outputs(12575) <= not (a xor b);
    outputs(12576) <= a and not b;
    outputs(12577) <= not a or b;
    outputs(12578) <= a or b;
    outputs(12579) <= not (a xor b);
    outputs(12580) <= a and not b;
    outputs(12581) <= not (a xor b);
    outputs(12582) <= not (a xor b);
    outputs(12583) <= not a;
    outputs(12584) <= not b;
    outputs(12585) <= not b;
    outputs(12586) <= not (a or b);
    outputs(12587) <= not (a xor b);
    outputs(12588) <= not (a or b);
    outputs(12589) <= a;
    outputs(12590) <= b;
    outputs(12591) <= a and b;
    outputs(12592) <= a or b;
    outputs(12593) <= a;
    outputs(12594) <= a and not b;
    outputs(12595) <= b;
    outputs(12596) <= not (a and b);
    outputs(12597) <= b and not a;
    outputs(12598) <= not a;
    outputs(12599) <= b;
    outputs(12600) <= not (a and b);
    outputs(12601) <= not b;
    outputs(12602) <= not b;
    outputs(12603) <= not b;
    outputs(12604) <= a xor b;
    outputs(12605) <= not b or a;
    outputs(12606) <= not (a xor b);
    outputs(12607) <= a xor b;
    outputs(12608) <= a xor b;
    outputs(12609) <= a and not b;
    outputs(12610) <= not (a xor b);
    outputs(12611) <= a and not b;
    outputs(12612) <= not (a or b);
    outputs(12613) <= not b;
    outputs(12614) <= not a;
    outputs(12615) <= a and not b;
    outputs(12616) <= not (a xor b);
    outputs(12617) <= a or b;
    outputs(12618) <= not (a xor b);
    outputs(12619) <= a;
    outputs(12620) <= not b;
    outputs(12621) <= not a;
    outputs(12622) <= not (a or b);
    outputs(12623) <= not (a and b);
    outputs(12624) <= a xor b;
    outputs(12625) <= a and not b;
    outputs(12626) <= not b or a;
    outputs(12627) <= not (a xor b);
    outputs(12628) <= not (a or b);
    outputs(12629) <= b and not a;
    outputs(12630) <= not a;
    outputs(12631) <= not a;
    outputs(12632) <= b and not a;
    outputs(12633) <= b and not a;
    outputs(12634) <= not (a xor b);
    outputs(12635) <= not b;
    outputs(12636) <= b and not a;
    outputs(12637) <= not (a xor b);
    outputs(12638) <= not b;
    outputs(12639) <= a xor b;
    outputs(12640) <= not a;
    outputs(12641) <= not b;
    outputs(12642) <= a xor b;
    outputs(12643) <= a;
    outputs(12644) <= a;
    outputs(12645) <= not a or b;
    outputs(12646) <= b and not a;
    outputs(12647) <= a and b;
    outputs(12648) <= a;
    outputs(12649) <= not (a xor b);
    outputs(12650) <= not b or a;
    outputs(12651) <= b and not a;
    outputs(12652) <= a and b;
    outputs(12653) <= a;
    outputs(12654) <= not (a xor b);
    outputs(12655) <= a and not b;
    outputs(12656) <= not a or b;
    outputs(12657) <= not a;
    outputs(12658) <= a and b;
    outputs(12659) <= not (a xor b);
    outputs(12660) <= a xor b;
    outputs(12661) <= a or b;
    outputs(12662) <= a;
    outputs(12663) <= a;
    outputs(12664) <= a xor b;
    outputs(12665) <= b;
    outputs(12666) <= a xor b;
    outputs(12667) <= not (a xor b);
    outputs(12668) <= a;
    outputs(12669) <= not (a or b);
    outputs(12670) <= not b;
    outputs(12671) <= not a;
    outputs(12672) <= not (a xor b);
    outputs(12673) <= a and not b;
    outputs(12674) <= not b;
    outputs(12675) <= not b;
    outputs(12676) <= not (a xor b);
    outputs(12677) <= a;
    outputs(12678) <= b;
    outputs(12679) <= b;
    outputs(12680) <= not b;
    outputs(12681) <= not (a and b);
    outputs(12682) <= a xor b;
    outputs(12683) <= a;
    outputs(12684) <= not (a or b);
    outputs(12685) <= b;
    outputs(12686) <= not a;
    outputs(12687) <= not b;
    outputs(12688) <= not b;
    outputs(12689) <= not (a xor b);
    outputs(12690) <= a;
    outputs(12691) <= not a;
    outputs(12692) <= a xor b;
    outputs(12693) <= not (a xor b);
    outputs(12694) <= not (a xor b);
    outputs(12695) <= not a;
    outputs(12696) <= not (a xor b);
    outputs(12697) <= not (a xor b);
    outputs(12698) <= a and b;
    outputs(12699) <= a;
    outputs(12700) <= a xor b;
    outputs(12701) <= not (a xor b);
    outputs(12702) <= a xor b;
    outputs(12703) <= b and not a;
    outputs(12704) <= not a;
    outputs(12705) <= not b;
    outputs(12706) <= a or b;
    outputs(12707) <= not b;
    outputs(12708) <= not (a and b);
    outputs(12709) <= not (a xor b);
    outputs(12710) <= not (a xor b);
    outputs(12711) <= a and not b;
    outputs(12712) <= b;
    outputs(12713) <= not a;
    outputs(12714) <= b and not a;
    outputs(12715) <= not (a xor b);
    outputs(12716) <= not (a or b);
    outputs(12717) <= a and b;
    outputs(12718) <= not a;
    outputs(12719) <= b and not a;
    outputs(12720) <= not a;
    outputs(12721) <= not (a xor b);
    outputs(12722) <= b;
    outputs(12723) <= not (a xor b);
    outputs(12724) <= not (a and b);
    outputs(12725) <= b and not a;
    outputs(12726) <= not a;
    outputs(12727) <= not (a xor b);
    outputs(12728) <= not a;
    outputs(12729) <= not a;
    outputs(12730) <= a;
    outputs(12731) <= a and b;
    outputs(12732) <= b and not a;
    outputs(12733) <= not a;
    outputs(12734) <= not (a xor b);
    outputs(12735) <= not (a and b);
    outputs(12736) <= not (a xor b);
    outputs(12737) <= not (a and b);
    outputs(12738) <= not b;
    outputs(12739) <= a;
    outputs(12740) <= a xor b;
    outputs(12741) <= a;
    outputs(12742) <= not (a xor b);
    outputs(12743) <= b and not a;
    outputs(12744) <= not (a xor b);
    outputs(12745) <= not (a xor b);
    outputs(12746) <= a and b;
    outputs(12747) <= b and not a;
    outputs(12748) <= a xor b;
    outputs(12749) <= not (a xor b);
    outputs(12750) <= not (a xor b);
    outputs(12751) <= a xor b;
    outputs(12752) <= not a or b;
    outputs(12753) <= not (a xor b);
    outputs(12754) <= not (a xor b);
    outputs(12755) <= not (a xor b);
    outputs(12756) <= a or b;
    outputs(12757) <= not (a or b);
    outputs(12758) <= not a;
    outputs(12759) <= a xor b;
    outputs(12760) <= a or b;
    outputs(12761) <= a xor b;
    outputs(12762) <= not a or b;
    outputs(12763) <= not b;
    outputs(12764) <= not b;
    outputs(12765) <= not a;
    outputs(12766) <= not b;
    outputs(12767) <= a xor b;
    outputs(12768) <= a and not b;
    outputs(12769) <= not a;
    outputs(12770) <= not (a or b);
    outputs(12771) <= b and not a;
    outputs(12772) <= b;
    outputs(12773) <= a xor b;
    outputs(12774) <= not a;
    outputs(12775) <= a xor b;
    outputs(12776) <= a;
    outputs(12777) <= not (a xor b);
    outputs(12778) <= not a;
    outputs(12779) <= b and not a;
    outputs(12780) <= not (a xor b);
    outputs(12781) <= not a;
    outputs(12782) <= a;
    outputs(12783) <= not (a xor b);
    outputs(12784) <= b;
    outputs(12785) <= a xor b;
    outputs(12786) <= not (a or b);
    outputs(12787) <= b;
    outputs(12788) <= not (a xor b);
    outputs(12789) <= a xor b;
    outputs(12790) <= a xor b;
    outputs(12791) <= not (a xor b);
    outputs(12792) <= b and not a;
    outputs(12793) <= not b;
    outputs(12794) <= b;
    outputs(12795) <= b;
    outputs(12796) <= not a;
    outputs(12797) <= not (a or b);
    outputs(12798) <= not a;
    outputs(12799) <= b;
end Behavioral;
