library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(2559 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);
    signal layer1_outputs : std_logic_vector(2559 downto 0);
    signal layer2_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not((inputs(224)) or (inputs(73)));
    layer0_outputs(1) <= inputs(166);
    layer0_outputs(2) <= not(inputs(247)) or (inputs(199));
    layer0_outputs(3) <= '0';
    layer0_outputs(4) <= not(inputs(94));
    layer0_outputs(5) <= (inputs(155)) or (inputs(236));
    layer0_outputs(6) <= not((inputs(224)) xor (inputs(193)));
    layer0_outputs(7) <= inputs(198);
    layer0_outputs(8) <= inputs(177);
    layer0_outputs(9) <= inputs(120);
    layer0_outputs(10) <= (inputs(187)) or (inputs(247));
    layer0_outputs(11) <= '0';
    layer0_outputs(12) <= not(inputs(108));
    layer0_outputs(13) <= (inputs(219)) or (inputs(98));
    layer0_outputs(14) <= (inputs(14)) or (inputs(168));
    layer0_outputs(15) <= inputs(194);
    layer0_outputs(16) <= (inputs(109)) and not (inputs(123));
    layer0_outputs(17) <= inputs(50);
    layer0_outputs(18) <= inputs(190);
    layer0_outputs(19) <= (inputs(118)) and not (inputs(91));
    layer0_outputs(20) <= inputs(6);
    layer0_outputs(21) <= (inputs(183)) and not (inputs(1));
    layer0_outputs(22) <= not(inputs(3)) or (inputs(78));
    layer0_outputs(23) <= '0';
    layer0_outputs(24) <= not(inputs(108)) or (inputs(5));
    layer0_outputs(25) <= not((inputs(226)) or (inputs(216)));
    layer0_outputs(26) <= not(inputs(224)) or (inputs(223));
    layer0_outputs(27) <= not(inputs(88));
    layer0_outputs(28) <= inputs(155);
    layer0_outputs(29) <= inputs(68);
    layer0_outputs(30) <= not(inputs(29)) or (inputs(223));
    layer0_outputs(31) <= not(inputs(91));
    layer0_outputs(32) <= (inputs(214)) or (inputs(254));
    layer0_outputs(33) <= not(inputs(102));
    layer0_outputs(34) <= inputs(101);
    layer0_outputs(35) <= inputs(135);
    layer0_outputs(36) <= not(inputs(17)) or (inputs(112));
    layer0_outputs(37) <= (inputs(244)) or (inputs(142));
    layer0_outputs(38) <= not(inputs(118)) or (inputs(170));
    layer0_outputs(39) <= '1';
    layer0_outputs(40) <= not((inputs(201)) or (inputs(234)));
    layer0_outputs(41) <= not(inputs(63)) or (inputs(229));
    layer0_outputs(42) <= not(inputs(123)) or (inputs(133));
    layer0_outputs(43) <= (inputs(225)) or (inputs(129));
    layer0_outputs(44) <= (inputs(46)) or (inputs(112));
    layer0_outputs(45) <= not(inputs(247)) or (inputs(208));
    layer0_outputs(46) <= not((inputs(204)) or (inputs(254)));
    layer0_outputs(47) <= (inputs(238)) and not (inputs(36));
    layer0_outputs(48) <= (inputs(230)) or (inputs(111));
    layer0_outputs(49) <= not((inputs(183)) and (inputs(70)));
    layer0_outputs(50) <= inputs(142);
    layer0_outputs(51) <= inputs(156);
    layer0_outputs(52) <= not(inputs(228)) or (inputs(208));
    layer0_outputs(53) <= '1';
    layer0_outputs(54) <= not(inputs(119));
    layer0_outputs(55) <= (inputs(127)) and not (inputs(53));
    layer0_outputs(56) <= not(inputs(31));
    layer0_outputs(57) <= not(inputs(10)) or (inputs(180));
    layer0_outputs(58) <= not(inputs(69));
    layer0_outputs(59) <= not(inputs(85)) or (inputs(6));
    layer0_outputs(60) <= not(inputs(50));
    layer0_outputs(61) <= (inputs(28)) and not (inputs(27));
    layer0_outputs(62) <= not(inputs(105));
    layer0_outputs(63) <= not(inputs(188)) or (inputs(223));
    layer0_outputs(64) <= inputs(93);
    layer0_outputs(65) <= (inputs(185)) and (inputs(72));
    layer0_outputs(66) <= not(inputs(29));
    layer0_outputs(67) <= not(inputs(73));
    layer0_outputs(68) <= (inputs(88)) or (inputs(144));
    layer0_outputs(69) <= inputs(231);
    layer0_outputs(70) <= not(inputs(69)) or (inputs(21));
    layer0_outputs(71) <= not((inputs(123)) or (inputs(216)));
    layer0_outputs(72) <= '0';
    layer0_outputs(73) <= (inputs(251)) or (inputs(185));
    layer0_outputs(74) <= '1';
    layer0_outputs(75) <= (inputs(158)) or (inputs(190));
    layer0_outputs(76) <= not(inputs(41));
    layer0_outputs(77) <= not(inputs(228)) or (inputs(111));
    layer0_outputs(78) <= inputs(204);
    layer0_outputs(79) <= not(inputs(142));
    layer0_outputs(80) <= not(inputs(124));
    layer0_outputs(81) <= '1';
    layer0_outputs(82) <= not(inputs(47));
    layer0_outputs(83) <= inputs(143);
    layer0_outputs(84) <= not(inputs(22)) or (inputs(127));
    layer0_outputs(85) <= (inputs(179)) or (inputs(127));
    layer0_outputs(86) <= not(inputs(238));
    layer0_outputs(87) <= inputs(231);
    layer0_outputs(88) <= not(inputs(136)) or (inputs(116));
    layer0_outputs(89) <= '0';
    layer0_outputs(90) <= (inputs(59)) or (inputs(53));
    layer0_outputs(91) <= (inputs(126)) and not (inputs(207));
    layer0_outputs(92) <= inputs(195);
    layer0_outputs(93) <= not(inputs(204));
    layer0_outputs(94) <= inputs(119);
    layer0_outputs(95) <= '0';
    layer0_outputs(96) <= (inputs(232)) and not (inputs(67));
    layer0_outputs(97) <= inputs(181);
    layer0_outputs(98) <= not((inputs(66)) xor (inputs(70)));
    layer0_outputs(99) <= not((inputs(199)) or (inputs(179)));
    layer0_outputs(100) <= (inputs(62)) or (inputs(163));
    layer0_outputs(101) <= inputs(151);
    layer0_outputs(102) <= '0';
    layer0_outputs(103) <= '1';
    layer0_outputs(104) <= not(inputs(254)) or (inputs(205));
    layer0_outputs(105) <= (inputs(229)) and not (inputs(59));
    layer0_outputs(106) <= not(inputs(188));
    layer0_outputs(107) <= (inputs(100)) and not (inputs(210));
    layer0_outputs(108) <= not((inputs(69)) or (inputs(135)));
    layer0_outputs(109) <= not((inputs(85)) or (inputs(115)));
    layer0_outputs(110) <= inputs(127);
    layer0_outputs(111) <= '0';
    layer0_outputs(112) <= not(inputs(37)) or (inputs(174));
    layer0_outputs(113) <= (inputs(224)) and (inputs(65));
    layer0_outputs(114) <= (inputs(161)) or (inputs(146));
    layer0_outputs(115) <= '1';
    layer0_outputs(116) <= not(inputs(222)) or (inputs(156));
    layer0_outputs(117) <= not(inputs(69));
    layer0_outputs(118) <= not((inputs(246)) and (inputs(78)));
    layer0_outputs(119) <= not(inputs(248)) or (inputs(77));
    layer0_outputs(120) <= not((inputs(194)) or (inputs(116)));
    layer0_outputs(121) <= (inputs(38)) and (inputs(104));
    layer0_outputs(122) <= inputs(102);
    layer0_outputs(123) <= not(inputs(69)) or (inputs(236));
    layer0_outputs(124) <= not(inputs(187));
    layer0_outputs(125) <= not(inputs(219)) or (inputs(106));
    layer0_outputs(126) <= (inputs(74)) and not (inputs(15));
    layer0_outputs(127) <= (inputs(66)) or (inputs(110));
    layer0_outputs(128) <= not((inputs(45)) or (inputs(68)));
    layer0_outputs(129) <= not((inputs(48)) or (inputs(76)));
    layer0_outputs(130) <= not(inputs(41));
    layer0_outputs(131) <= inputs(86);
    layer0_outputs(132) <= inputs(60);
    layer0_outputs(133) <= (inputs(36)) and not (inputs(180));
    layer0_outputs(134) <= inputs(23);
    layer0_outputs(135) <= inputs(198);
    layer0_outputs(136) <= not((inputs(237)) or (inputs(184)));
    layer0_outputs(137) <= not(inputs(212));
    layer0_outputs(138) <= inputs(188);
    layer0_outputs(139) <= not(inputs(223)) or (inputs(55));
    layer0_outputs(140) <= inputs(119);
    layer0_outputs(141) <= (inputs(189)) or (inputs(89));
    layer0_outputs(142) <= not(inputs(27));
    layer0_outputs(143) <= not((inputs(120)) xor (inputs(45)));
    layer0_outputs(144) <= not(inputs(174)) or (inputs(228));
    layer0_outputs(145) <= (inputs(111)) or (inputs(17));
    layer0_outputs(146) <= not(inputs(43));
    layer0_outputs(147) <= not((inputs(114)) xor (inputs(217)));
    layer0_outputs(148) <= not((inputs(143)) or (inputs(140)));
    layer0_outputs(149) <= inputs(253);
    layer0_outputs(150) <= (inputs(208)) or (inputs(4));
    layer0_outputs(151) <= not((inputs(110)) or (inputs(155)));
    layer0_outputs(152) <= '1';
    layer0_outputs(153) <= (inputs(80)) and not (inputs(235));
    layer0_outputs(154) <= (inputs(29)) and not (inputs(252));
    layer0_outputs(155) <= inputs(117);
    layer0_outputs(156) <= not(inputs(177)) or (inputs(182));
    layer0_outputs(157) <= (inputs(145)) and not (inputs(119));
    layer0_outputs(158) <= not((inputs(33)) and (inputs(114)));
    layer0_outputs(159) <= not((inputs(108)) and (inputs(70)));
    layer0_outputs(160) <= not(inputs(179));
    layer0_outputs(161) <= not((inputs(73)) xor (inputs(13)));
    layer0_outputs(162) <= (inputs(96)) or (inputs(123));
    layer0_outputs(163) <= (inputs(141)) or (inputs(47));
    layer0_outputs(164) <= inputs(39);
    layer0_outputs(165) <= not(inputs(196));
    layer0_outputs(166) <= (inputs(7)) or (inputs(215));
    layer0_outputs(167) <= inputs(69);
    layer0_outputs(168) <= '1';
    layer0_outputs(169) <= (inputs(52)) or (inputs(97));
    layer0_outputs(170) <= (inputs(117)) and not (inputs(172));
    layer0_outputs(171) <= (inputs(122)) or (inputs(131));
    layer0_outputs(172) <= not((inputs(171)) or (inputs(223)));
    layer0_outputs(173) <= not((inputs(172)) or (inputs(203)));
    layer0_outputs(174) <= not(inputs(149));
    layer0_outputs(175) <= not(inputs(19)) or (inputs(156));
    layer0_outputs(176) <= not(inputs(29)) or (inputs(206));
    layer0_outputs(177) <= inputs(146);
    layer0_outputs(178) <= not(inputs(1)) or (inputs(255));
    layer0_outputs(179) <= (inputs(187)) and not (inputs(46));
    layer0_outputs(180) <= (inputs(166)) or (inputs(119));
    layer0_outputs(181) <= not((inputs(201)) or (inputs(35)));
    layer0_outputs(182) <= inputs(123);
    layer0_outputs(183) <= inputs(160);
    layer0_outputs(184) <= not((inputs(57)) and (inputs(44)));
    layer0_outputs(185) <= (inputs(171)) and (inputs(184));
    layer0_outputs(186) <= not(inputs(87));
    layer0_outputs(187) <= not((inputs(91)) or (inputs(10)));
    layer0_outputs(188) <= (inputs(211)) or (inputs(239));
    layer0_outputs(189) <= (inputs(60)) xor (inputs(72));
    layer0_outputs(190) <= inputs(59);
    layer0_outputs(191) <= not(inputs(168));
    layer0_outputs(192) <= not((inputs(82)) or (inputs(248)));
    layer0_outputs(193) <= (inputs(175)) and (inputs(79));
    layer0_outputs(194) <= not(inputs(119));
    layer0_outputs(195) <= not((inputs(159)) or (inputs(66)));
    layer0_outputs(196) <= not((inputs(66)) or (inputs(171)));
    layer0_outputs(197) <= '0';
    layer0_outputs(198) <= (inputs(154)) and not (inputs(63));
    layer0_outputs(199) <= not(inputs(188));
    layer0_outputs(200) <= not(inputs(107));
    layer0_outputs(201) <= (inputs(7)) and not (inputs(217));
    layer0_outputs(202) <= not(inputs(197)) or (inputs(30));
    layer0_outputs(203) <= (inputs(244)) or (inputs(88));
    layer0_outputs(204) <= inputs(203);
    layer0_outputs(205) <= inputs(178);
    layer0_outputs(206) <= inputs(191);
    layer0_outputs(207) <= not(inputs(11));
    layer0_outputs(208) <= (inputs(130)) and not (inputs(192));
    layer0_outputs(209) <= inputs(216);
    layer0_outputs(210) <= not((inputs(13)) and (inputs(31)));
    layer0_outputs(211) <= not((inputs(20)) or (inputs(191)));
    layer0_outputs(212) <= '1';
    layer0_outputs(213) <= not(inputs(235));
    layer0_outputs(214) <= inputs(241);
    layer0_outputs(215) <= inputs(183);
    layer0_outputs(216) <= (inputs(164)) and not (inputs(62));
    layer0_outputs(217) <= not(inputs(44));
    layer0_outputs(218) <= (inputs(131)) or (inputs(116));
    layer0_outputs(219) <= (inputs(162)) and not (inputs(25));
    layer0_outputs(220) <= not(inputs(183)) or (inputs(177));
    layer0_outputs(221) <= not(inputs(255)) or (inputs(13));
    layer0_outputs(222) <= not((inputs(38)) or (inputs(79)));
    layer0_outputs(223) <= inputs(244);
    layer0_outputs(224) <= (inputs(12)) xor (inputs(24));
    layer0_outputs(225) <= (inputs(202)) or (inputs(82));
    layer0_outputs(226) <= inputs(221);
    layer0_outputs(227) <= not(inputs(84));
    layer0_outputs(228) <= not((inputs(96)) and (inputs(8)));
    layer0_outputs(229) <= (inputs(42)) or (inputs(65));
    layer0_outputs(230) <= not(inputs(92));
    layer0_outputs(231) <= (inputs(79)) xor (inputs(20));
    layer0_outputs(232) <= inputs(138);
    layer0_outputs(233) <= (inputs(219)) or (inputs(201));
    layer0_outputs(234) <= not(inputs(68)) or (inputs(61));
    layer0_outputs(235) <= not(inputs(178));
    layer0_outputs(236) <= not(inputs(164));
    layer0_outputs(237) <= not((inputs(57)) or (inputs(176)));
    layer0_outputs(238) <= not(inputs(69));
    layer0_outputs(239) <= (inputs(188)) and not (inputs(147));
    layer0_outputs(240) <= (inputs(52)) or (inputs(67));
    layer0_outputs(241) <= not(inputs(226));
    layer0_outputs(242) <= not(inputs(148)) or (inputs(176));
    layer0_outputs(243) <= not((inputs(156)) and (inputs(70)));
    layer0_outputs(244) <= not((inputs(197)) or (inputs(215)));
    layer0_outputs(245) <= inputs(74);
    layer0_outputs(246) <= not((inputs(134)) or (inputs(192)));
    layer0_outputs(247) <= (inputs(63)) or (inputs(46));
    layer0_outputs(248) <= inputs(168);
    layer0_outputs(249) <= not(inputs(202));
    layer0_outputs(250) <= not(inputs(168)) or (inputs(62));
    layer0_outputs(251) <= not(inputs(223)) or (inputs(107));
    layer0_outputs(252) <= (inputs(147)) and not (inputs(175));
    layer0_outputs(253) <= (inputs(51)) xor (inputs(55));
    layer0_outputs(254) <= (inputs(190)) or (inputs(146));
    layer0_outputs(255) <= inputs(146);
    layer0_outputs(256) <= not(inputs(83));
    layer0_outputs(257) <= '1';
    layer0_outputs(258) <= (inputs(50)) and (inputs(161));
    layer0_outputs(259) <= inputs(201);
    layer0_outputs(260) <= inputs(217);
    layer0_outputs(261) <= not(inputs(123));
    layer0_outputs(262) <= (inputs(173)) and not (inputs(249));
    layer0_outputs(263) <= (inputs(150)) and not (inputs(141));
    layer0_outputs(264) <= (inputs(247)) and not (inputs(0));
    layer0_outputs(265) <= not(inputs(228)) or (inputs(142));
    layer0_outputs(266) <= inputs(247);
    layer0_outputs(267) <= (inputs(188)) and not (inputs(110));
    layer0_outputs(268) <= not((inputs(132)) and (inputs(179)));
    layer0_outputs(269) <= (inputs(163)) and not (inputs(191));
    layer0_outputs(270) <= not((inputs(96)) or (inputs(195)));
    layer0_outputs(271) <= not(inputs(255)) or (inputs(179));
    layer0_outputs(272) <= (inputs(213)) or (inputs(129));
    layer0_outputs(273) <= (inputs(32)) or (inputs(169));
    layer0_outputs(274) <= (inputs(37)) and not (inputs(203));
    layer0_outputs(275) <= not(inputs(128));
    layer0_outputs(276) <= inputs(110);
    layer0_outputs(277) <= '1';
    layer0_outputs(278) <= not((inputs(91)) or (inputs(83)));
    layer0_outputs(279) <= not((inputs(144)) and (inputs(39)));
    layer0_outputs(280) <= '0';
    layer0_outputs(281) <= not(inputs(102));
    layer0_outputs(282) <= not(inputs(27)) or (inputs(150));
    layer0_outputs(283) <= not((inputs(42)) or (inputs(236)));
    layer0_outputs(284) <= not(inputs(247)) or (inputs(151));
    layer0_outputs(285) <= inputs(2);
    layer0_outputs(286) <= inputs(251);
    layer0_outputs(287) <= (inputs(148)) xor (inputs(68));
    layer0_outputs(288) <= (inputs(70)) and not (inputs(105));
    layer0_outputs(289) <= not((inputs(154)) or (inputs(191)));
    layer0_outputs(290) <= not(inputs(115)) or (inputs(32));
    layer0_outputs(291) <= inputs(84);
    layer0_outputs(292) <= (inputs(127)) and not (inputs(175));
    layer0_outputs(293) <= (inputs(233)) or (inputs(240));
    layer0_outputs(294) <= inputs(99);
    layer0_outputs(295) <= not((inputs(232)) xor (inputs(234)));
    layer0_outputs(296) <= not(inputs(115));
    layer0_outputs(297) <= not(inputs(82));
    layer0_outputs(298) <= not(inputs(20)) or (inputs(94));
    layer0_outputs(299) <= (inputs(52)) and not (inputs(205));
    layer0_outputs(300) <= inputs(195);
    layer0_outputs(301) <= (inputs(177)) xor (inputs(209));
    layer0_outputs(302) <= not(inputs(167));
    layer0_outputs(303) <= inputs(160);
    layer0_outputs(304) <= inputs(68);
    layer0_outputs(305) <= not((inputs(104)) xor (inputs(10)));
    layer0_outputs(306) <= not((inputs(185)) or (inputs(144)));
    layer0_outputs(307) <= not(inputs(246));
    layer0_outputs(308) <= (inputs(59)) or (inputs(141));
    layer0_outputs(309) <= not(inputs(114)) or (inputs(240));
    layer0_outputs(310) <= '1';
    layer0_outputs(311) <= not(inputs(10)) or (inputs(238));
    layer0_outputs(312) <= not(inputs(231)) or (inputs(167));
    layer0_outputs(313) <= inputs(141);
    layer0_outputs(314) <= '1';
    layer0_outputs(315) <= not((inputs(141)) or (inputs(138)));
    layer0_outputs(316) <= (inputs(41)) and (inputs(28));
    layer0_outputs(317) <= (inputs(52)) or (inputs(153));
    layer0_outputs(318) <= inputs(1);
    layer0_outputs(319) <= not((inputs(238)) xor (inputs(1)));
    layer0_outputs(320) <= inputs(76);
    layer0_outputs(321) <= inputs(75);
    layer0_outputs(322) <= inputs(83);
    layer0_outputs(323) <= not(inputs(147)) or (inputs(11));
    layer0_outputs(324) <= inputs(94);
    layer0_outputs(325) <= '0';
    layer0_outputs(326) <= not((inputs(74)) and (inputs(195)));
    layer0_outputs(327) <= not(inputs(34)) or (inputs(250));
    layer0_outputs(328) <= not(inputs(178));
    layer0_outputs(329) <= (inputs(231)) and (inputs(182));
    layer0_outputs(330) <= (inputs(230)) or (inputs(80));
    layer0_outputs(331) <= not((inputs(13)) xor (inputs(122)));
    layer0_outputs(332) <= not((inputs(101)) or (inputs(8)));
    layer0_outputs(333) <= not((inputs(143)) or (inputs(159)));
    layer0_outputs(334) <= (inputs(122)) and not (inputs(216));
    layer0_outputs(335) <= not((inputs(170)) or (inputs(108)));
    layer0_outputs(336) <= not((inputs(117)) or (inputs(147)));
    layer0_outputs(337) <= inputs(69);
    layer0_outputs(338) <= not((inputs(105)) or (inputs(153)));
    layer0_outputs(339) <= '1';
    layer0_outputs(340) <= inputs(22);
    layer0_outputs(341) <= inputs(9);
    layer0_outputs(342) <= (inputs(250)) and not (inputs(116));
    layer0_outputs(343) <= not(inputs(158)) or (inputs(28));
    layer0_outputs(344) <= (inputs(142)) and not (inputs(41));
    layer0_outputs(345) <= not(inputs(71)) or (inputs(4));
    layer0_outputs(346) <= not(inputs(115));
    layer0_outputs(347) <= (inputs(51)) and not (inputs(112));
    layer0_outputs(348) <= (inputs(49)) or (inputs(164));
    layer0_outputs(349) <= not((inputs(85)) xor (inputs(88)));
    layer0_outputs(350) <= not(inputs(247));
    layer0_outputs(351) <= inputs(167);
    layer0_outputs(352) <= not(inputs(214)) or (inputs(152));
    layer0_outputs(353) <= (inputs(155)) or (inputs(139));
    layer0_outputs(354) <= not((inputs(52)) or (inputs(162)));
    layer0_outputs(355) <= (inputs(17)) or (inputs(35));
    layer0_outputs(356) <= '0';
    layer0_outputs(357) <= not((inputs(106)) or (inputs(83)));
    layer0_outputs(358) <= not(inputs(247));
    layer0_outputs(359) <= inputs(133);
    layer0_outputs(360) <= (inputs(220)) and not (inputs(233));
    layer0_outputs(361) <= (inputs(108)) and not (inputs(104));
    layer0_outputs(362) <= (inputs(157)) xor (inputs(121));
    layer0_outputs(363) <= not((inputs(59)) or (inputs(58)));
    layer0_outputs(364) <= not((inputs(63)) or (inputs(76)));
    layer0_outputs(365) <= inputs(239);
    layer0_outputs(366) <= (inputs(131)) and (inputs(212));
    layer0_outputs(367) <= inputs(105);
    layer0_outputs(368) <= inputs(66);
    layer0_outputs(369) <= inputs(62);
    layer0_outputs(370) <= (inputs(35)) xor (inputs(207));
    layer0_outputs(371) <= inputs(227);
    layer0_outputs(372) <= inputs(61);
    layer0_outputs(373) <= not((inputs(241)) or (inputs(56)));
    layer0_outputs(374) <= inputs(147);
    layer0_outputs(375) <= '0';
    layer0_outputs(376) <= inputs(127);
    layer0_outputs(377) <= (inputs(208)) or (inputs(99));
    layer0_outputs(378) <= '0';
    layer0_outputs(379) <= not((inputs(162)) xor (inputs(249)));
    layer0_outputs(380) <= not(inputs(29));
    layer0_outputs(381) <= '1';
    layer0_outputs(382) <= not(inputs(137)) or (inputs(205));
    layer0_outputs(383) <= (inputs(213)) and not (inputs(85));
    layer0_outputs(384) <= not(inputs(103));
    layer0_outputs(385) <= not(inputs(211));
    layer0_outputs(386) <= (inputs(105)) and (inputs(205));
    layer0_outputs(387) <= not(inputs(102)) or (inputs(83));
    layer0_outputs(388) <= not(inputs(171));
    layer0_outputs(389) <= not(inputs(9));
    layer0_outputs(390) <= (inputs(90)) and not (inputs(133));
    layer0_outputs(391) <= not(inputs(20)) or (inputs(100));
    layer0_outputs(392) <= (inputs(167)) and not (inputs(4));
    layer0_outputs(393) <= (inputs(196)) or (inputs(237));
    layer0_outputs(394) <= (inputs(197)) or (inputs(97));
    layer0_outputs(395) <= not(inputs(111)) or (inputs(98));
    layer0_outputs(396) <= '0';
    layer0_outputs(397) <= not(inputs(185)) or (inputs(210));
    layer0_outputs(398) <= (inputs(38)) and not (inputs(132));
    layer0_outputs(399) <= (inputs(173)) or (inputs(222));
    layer0_outputs(400) <= not((inputs(79)) and (inputs(200)));
    layer0_outputs(401) <= not(inputs(108));
    layer0_outputs(402) <= (inputs(152)) and not (inputs(217));
    layer0_outputs(403) <= '1';
    layer0_outputs(404) <= not((inputs(131)) xor (inputs(80)));
    layer0_outputs(405) <= inputs(249);
    layer0_outputs(406) <= inputs(23);
    layer0_outputs(407) <= not((inputs(58)) or (inputs(108)));
    layer0_outputs(408) <= not(inputs(163)) or (inputs(161));
    layer0_outputs(409) <= (inputs(120)) xor (inputs(245));
    layer0_outputs(410) <= not(inputs(228));
    layer0_outputs(411) <= (inputs(160)) or (inputs(41));
    layer0_outputs(412) <= (inputs(172)) and not (inputs(139));
    layer0_outputs(413) <= not(inputs(106)) or (inputs(237));
    layer0_outputs(414) <= (inputs(160)) or (inputs(227));
    layer0_outputs(415) <= not((inputs(232)) or (inputs(21)));
    layer0_outputs(416) <= (inputs(221)) xor (inputs(251));
    layer0_outputs(417) <= (inputs(121)) and not (inputs(157));
    layer0_outputs(418) <= not(inputs(59)) or (inputs(13));
    layer0_outputs(419) <= '0';
    layer0_outputs(420) <= not(inputs(192)) or (inputs(47));
    layer0_outputs(421) <= not(inputs(245));
    layer0_outputs(422) <= not(inputs(70)) or (inputs(116));
    layer0_outputs(423) <= (inputs(68)) or (inputs(194));
    layer0_outputs(424) <= inputs(180);
    layer0_outputs(425) <= (inputs(137)) and not (inputs(57));
    layer0_outputs(426) <= not((inputs(147)) or (inputs(147)));
    layer0_outputs(427) <= inputs(104);
    layer0_outputs(428) <= not(inputs(54)) or (inputs(110));
    layer0_outputs(429) <= (inputs(181)) and (inputs(54));
    layer0_outputs(430) <= '1';
    layer0_outputs(431) <= inputs(105);
    layer0_outputs(432) <= not(inputs(229)) or (inputs(166));
    layer0_outputs(433) <= (inputs(189)) or (inputs(187));
    layer0_outputs(434) <= inputs(176);
    layer0_outputs(435) <= inputs(172);
    layer0_outputs(436) <= (inputs(16)) and (inputs(201));
    layer0_outputs(437) <= '0';
    layer0_outputs(438) <= not(inputs(245));
    layer0_outputs(439) <= inputs(152);
    layer0_outputs(440) <= not(inputs(57));
    layer0_outputs(441) <= not((inputs(71)) or (inputs(83)));
    layer0_outputs(442) <= (inputs(211)) and (inputs(30));
    layer0_outputs(443) <= not(inputs(100));
    layer0_outputs(444) <= not(inputs(118));
    layer0_outputs(445) <= not(inputs(155));
    layer0_outputs(446) <= not((inputs(75)) and (inputs(215)));
    layer0_outputs(447) <= not(inputs(158));
    layer0_outputs(448) <= inputs(83);
    layer0_outputs(449) <= not(inputs(119));
    layer0_outputs(450) <= '1';
    layer0_outputs(451) <= (inputs(23)) and not (inputs(77));
    layer0_outputs(452) <= not(inputs(98)) or (inputs(93));
    layer0_outputs(453) <= not(inputs(119)) or (inputs(56));
    layer0_outputs(454) <= (inputs(234)) or (inputs(226));
    layer0_outputs(455) <= not(inputs(246));
    layer0_outputs(456) <= not(inputs(68));
    layer0_outputs(457) <= (inputs(9)) or (inputs(73));
    layer0_outputs(458) <= (inputs(97)) and not (inputs(62));
    layer0_outputs(459) <= inputs(19);
    layer0_outputs(460) <= (inputs(241)) or (inputs(108));
    layer0_outputs(461) <= inputs(119);
    layer0_outputs(462) <= not(inputs(231));
    layer0_outputs(463) <= inputs(27);
    layer0_outputs(464) <= inputs(191);
    layer0_outputs(465) <= (inputs(104)) or (inputs(66));
    layer0_outputs(466) <= not(inputs(89));
    layer0_outputs(467) <= (inputs(30)) xor (inputs(1));
    layer0_outputs(468) <= inputs(151);
    layer0_outputs(469) <= (inputs(184)) and (inputs(43));
    layer0_outputs(470) <= (inputs(24)) or (inputs(62));
    layer0_outputs(471) <= '1';
    layer0_outputs(472) <= not((inputs(252)) xor (inputs(43)));
    layer0_outputs(473) <= not((inputs(32)) and (inputs(149)));
    layer0_outputs(474) <= (inputs(191)) and not (inputs(66));
    layer0_outputs(475) <= not((inputs(169)) or (inputs(83)));
    layer0_outputs(476) <= not((inputs(82)) or (inputs(47)));
    layer0_outputs(477) <= not(inputs(156));
    layer0_outputs(478) <= not(inputs(169));
    layer0_outputs(479) <= inputs(150);
    layer0_outputs(480) <= (inputs(174)) and not (inputs(91));
    layer0_outputs(481) <= not(inputs(72)) or (inputs(88));
    layer0_outputs(482) <= inputs(39);
    layer0_outputs(483) <= not(inputs(118));
    layer0_outputs(484) <= not((inputs(239)) and (inputs(247)));
    layer0_outputs(485) <= (inputs(172)) and not (inputs(122));
    layer0_outputs(486) <= (inputs(85)) and not (inputs(255));
    layer0_outputs(487) <= not(inputs(101));
    layer0_outputs(488) <= inputs(86);
    layer0_outputs(489) <= not(inputs(46));
    layer0_outputs(490) <= not(inputs(122));
    layer0_outputs(491) <= (inputs(173)) or (inputs(181));
    layer0_outputs(492) <= not(inputs(139));
    layer0_outputs(493) <= not(inputs(58)) or (inputs(136));
    layer0_outputs(494) <= not(inputs(42));
    layer0_outputs(495) <= not(inputs(22)) or (inputs(201));
    layer0_outputs(496) <= not(inputs(102));
    layer0_outputs(497) <= not(inputs(6));
    layer0_outputs(498) <= inputs(218);
    layer0_outputs(499) <= not((inputs(188)) and (inputs(44)));
    layer0_outputs(500) <= '1';
    layer0_outputs(501) <= not((inputs(124)) or (inputs(145)));
    layer0_outputs(502) <= not(inputs(165));
    layer0_outputs(503) <= not(inputs(146));
    layer0_outputs(504) <= inputs(77);
    layer0_outputs(505) <= '1';
    layer0_outputs(506) <= not((inputs(3)) or (inputs(14)));
    layer0_outputs(507) <= (inputs(95)) or (inputs(255));
    layer0_outputs(508) <= not(inputs(22));
    layer0_outputs(509) <= inputs(147);
    layer0_outputs(510) <= not(inputs(140));
    layer0_outputs(511) <= not((inputs(240)) or (inputs(160)));
    layer0_outputs(512) <= '1';
    layer0_outputs(513) <= '1';
    layer0_outputs(514) <= not((inputs(58)) and (inputs(218)));
    layer0_outputs(515) <= (inputs(89)) or (inputs(58));
    layer0_outputs(516) <= (inputs(0)) and not (inputs(205));
    layer0_outputs(517) <= not(inputs(143));
    layer0_outputs(518) <= not(inputs(243)) or (inputs(145));
    layer0_outputs(519) <= not((inputs(1)) or (inputs(204)));
    layer0_outputs(520) <= not(inputs(145)) or (inputs(56));
    layer0_outputs(521) <= inputs(195);
    layer0_outputs(522) <= not(inputs(76));
    layer0_outputs(523) <= '0';
    layer0_outputs(524) <= '0';
    layer0_outputs(525) <= (inputs(85)) or (inputs(69));
    layer0_outputs(526) <= not((inputs(22)) or (inputs(32)));
    layer0_outputs(527) <= inputs(64);
    layer0_outputs(528) <= (inputs(49)) or (inputs(243));
    layer0_outputs(529) <= not(inputs(213));
    layer0_outputs(530) <= not((inputs(249)) or (inputs(22)));
    layer0_outputs(531) <= not(inputs(229));
    layer0_outputs(532) <= inputs(131);
    layer0_outputs(533) <= not(inputs(34));
    layer0_outputs(534) <= inputs(165);
    layer0_outputs(535) <= (inputs(36)) and (inputs(34));
    layer0_outputs(536) <= inputs(135);
    layer0_outputs(537) <= not(inputs(118)) or (inputs(115));
    layer0_outputs(538) <= (inputs(183)) and not (inputs(186));
    layer0_outputs(539) <= '0';
    layer0_outputs(540) <= '1';
    layer0_outputs(541) <= (inputs(178)) or (inputs(148));
    layer0_outputs(542) <= inputs(227);
    layer0_outputs(543) <= '1';
    layer0_outputs(544) <= not((inputs(55)) and (inputs(156)));
    layer0_outputs(545) <= inputs(63);
    layer0_outputs(546) <= (inputs(149)) and not (inputs(160));
    layer0_outputs(547) <= not(inputs(175));
    layer0_outputs(548) <= not((inputs(200)) or (inputs(21)));
    layer0_outputs(549) <= not(inputs(85));
    layer0_outputs(550) <= (inputs(211)) and not (inputs(144));
    layer0_outputs(551) <= '0';
    layer0_outputs(552) <= not(inputs(213));
    layer0_outputs(553) <= not((inputs(73)) or (inputs(190)));
    layer0_outputs(554) <= (inputs(202)) and not (inputs(144));
    layer0_outputs(555) <= (inputs(91)) or (inputs(32));
    layer0_outputs(556) <= not(inputs(76)) or (inputs(181));
    layer0_outputs(557) <= not(inputs(180)) or (inputs(31));
    layer0_outputs(558) <= '1';
    layer0_outputs(559) <= (inputs(96)) or (inputs(220));
    layer0_outputs(560) <= inputs(60);
    layer0_outputs(561) <= (inputs(19)) and not (inputs(222));
    layer0_outputs(562) <= (inputs(166)) or (inputs(89));
    layer0_outputs(563) <= (inputs(74)) and not (inputs(2));
    layer0_outputs(564) <= not(inputs(210));
    layer0_outputs(565) <= '1';
    layer0_outputs(566) <= (inputs(255)) or (inputs(91));
    layer0_outputs(567) <= not(inputs(202));
    layer0_outputs(568) <= inputs(24);
    layer0_outputs(569) <= inputs(81);
    layer0_outputs(570) <= not((inputs(136)) or (inputs(253)));
    layer0_outputs(571) <= not((inputs(91)) or (inputs(68)));
    layer0_outputs(572) <= not(inputs(104));
    layer0_outputs(573) <= (inputs(30)) or (inputs(35));
    layer0_outputs(574) <= not(inputs(59));
    layer0_outputs(575) <= not(inputs(238)) or (inputs(65));
    layer0_outputs(576) <= (inputs(159)) or (inputs(174));
    layer0_outputs(577) <= not(inputs(21));
    layer0_outputs(578) <= inputs(127);
    layer0_outputs(579) <= (inputs(82)) or (inputs(101));
    layer0_outputs(580) <= inputs(102);
    layer0_outputs(581) <= not(inputs(217)) or (inputs(237));
    layer0_outputs(582) <= (inputs(31)) or (inputs(211));
    layer0_outputs(583) <= inputs(217);
    layer0_outputs(584) <= inputs(152);
    layer0_outputs(585) <= inputs(177);
    layer0_outputs(586) <= (inputs(169)) and (inputs(219));
    layer0_outputs(587) <= not(inputs(109));
    layer0_outputs(588) <= not(inputs(192)) or (inputs(46));
    layer0_outputs(589) <= inputs(229);
    layer0_outputs(590) <= (inputs(219)) and not (inputs(185));
    layer0_outputs(591) <= not(inputs(35)) or (inputs(207));
    layer0_outputs(592) <= (inputs(118)) and not (inputs(253));
    layer0_outputs(593) <= not((inputs(88)) xor (inputs(113)));
    layer0_outputs(594) <= not(inputs(156)) or (inputs(149));
    layer0_outputs(595) <= not(inputs(223));
    layer0_outputs(596) <= (inputs(80)) and (inputs(69));
    layer0_outputs(597) <= not(inputs(205));
    layer0_outputs(598) <= '1';
    layer0_outputs(599) <= not(inputs(215)) or (inputs(15));
    layer0_outputs(600) <= not((inputs(217)) and (inputs(48)));
    layer0_outputs(601) <= (inputs(168)) and not (inputs(160));
    layer0_outputs(602) <= not(inputs(228)) or (inputs(20));
    layer0_outputs(603) <= not(inputs(149)) or (inputs(14));
    layer0_outputs(604) <= not(inputs(7));
    layer0_outputs(605) <= (inputs(10)) and not (inputs(109));
    layer0_outputs(606) <= inputs(84);
    layer0_outputs(607) <= not(inputs(163));
    layer0_outputs(608) <= (inputs(136)) xor (inputs(81));
    layer0_outputs(609) <= not(inputs(121));
    layer0_outputs(610) <= inputs(198);
    layer0_outputs(611) <= not((inputs(140)) or (inputs(193)));
    layer0_outputs(612) <= inputs(250);
    layer0_outputs(613) <= inputs(166);
    layer0_outputs(614) <= '1';
    layer0_outputs(615) <= (inputs(104)) or (inputs(29));
    layer0_outputs(616) <= not((inputs(148)) or (inputs(98)));
    layer0_outputs(617) <= (inputs(219)) and not (inputs(31));
    layer0_outputs(618) <= '0';
    layer0_outputs(619) <= not(inputs(130)) or (inputs(136));
    layer0_outputs(620) <= (inputs(199)) and not (inputs(158));
    layer0_outputs(621) <= inputs(229);
    layer0_outputs(622) <= '0';
    layer0_outputs(623) <= (inputs(130)) and (inputs(76));
    layer0_outputs(624) <= (inputs(12)) and not (inputs(59));
    layer0_outputs(625) <= (inputs(45)) and not (inputs(81));
    layer0_outputs(626) <= not(inputs(142));
    layer0_outputs(627) <= '0';
    layer0_outputs(628) <= (inputs(134)) and (inputs(242));
    layer0_outputs(629) <= not((inputs(43)) or (inputs(232)));
    layer0_outputs(630) <= inputs(80);
    layer0_outputs(631) <= not((inputs(178)) or (inputs(95)));
    layer0_outputs(632) <= (inputs(161)) or (inputs(239));
    layer0_outputs(633) <= (inputs(69)) or (inputs(209));
    layer0_outputs(634) <= '1';
    layer0_outputs(635) <= not(inputs(236));
    layer0_outputs(636) <= (inputs(62)) and not (inputs(141));
    layer0_outputs(637) <= not(inputs(44)) or (inputs(79));
    layer0_outputs(638) <= not(inputs(70));
    layer0_outputs(639) <= not((inputs(45)) and (inputs(157)));
    layer0_outputs(640) <= not(inputs(167));
    layer0_outputs(641) <= (inputs(185)) or (inputs(237));
    layer0_outputs(642) <= not((inputs(153)) or (inputs(158)));
    layer0_outputs(643) <= not((inputs(18)) or (inputs(163)));
    layer0_outputs(644) <= not((inputs(16)) xor (inputs(81)));
    layer0_outputs(645) <= not((inputs(19)) xor (inputs(130)));
    layer0_outputs(646) <= '1';
    layer0_outputs(647) <= not(inputs(87));
    layer0_outputs(648) <= inputs(122);
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= not(inputs(213)) or (inputs(78));
    layer0_outputs(651) <= not((inputs(246)) or (inputs(173)));
    layer0_outputs(652) <= not(inputs(208)) or (inputs(68));
    layer0_outputs(653) <= inputs(166);
    layer0_outputs(654) <= (inputs(184)) and (inputs(157));
    layer0_outputs(655) <= (inputs(182)) and (inputs(7));
    layer0_outputs(656) <= (inputs(189)) or (inputs(173));
    layer0_outputs(657) <= inputs(4);
    layer0_outputs(658) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(659) <= not(inputs(197)) or (inputs(98));
    layer0_outputs(660) <= inputs(163);
    layer0_outputs(661) <= not(inputs(130));
    layer0_outputs(662) <= not((inputs(168)) or (inputs(66)));
    layer0_outputs(663) <= (inputs(196)) and (inputs(164));
    layer0_outputs(664) <= not(inputs(138)) or (inputs(39));
    layer0_outputs(665) <= (inputs(190)) and not (inputs(239));
    layer0_outputs(666) <= inputs(83);
    layer0_outputs(667) <= '0';
    layer0_outputs(668) <= not(inputs(119));
    layer0_outputs(669) <= inputs(181);
    layer0_outputs(670) <= not(inputs(55));
    layer0_outputs(671) <= not(inputs(6));
    layer0_outputs(672) <= (inputs(34)) or (inputs(196));
    layer0_outputs(673) <= inputs(122);
    layer0_outputs(674) <= not((inputs(250)) or (inputs(152)));
    layer0_outputs(675) <= (inputs(65)) or (inputs(51));
    layer0_outputs(676) <= (inputs(169)) or (inputs(157));
    layer0_outputs(677) <= inputs(109);
    layer0_outputs(678) <= not(inputs(109));
    layer0_outputs(679) <= not((inputs(50)) or (inputs(152)));
    layer0_outputs(680) <= not(inputs(101));
    layer0_outputs(681) <= (inputs(47)) and not (inputs(15));
    layer0_outputs(682) <= not(inputs(92)) or (inputs(223));
    layer0_outputs(683) <= not(inputs(197));
    layer0_outputs(684) <= inputs(215);
    layer0_outputs(685) <= (inputs(165)) and not (inputs(133));
    layer0_outputs(686) <= not((inputs(88)) or (inputs(215)));
    layer0_outputs(687) <= not(inputs(118));
    layer0_outputs(688) <= not(inputs(73)) or (inputs(77));
    layer0_outputs(689) <= '1';
    layer0_outputs(690) <= (inputs(55)) and not (inputs(240));
    layer0_outputs(691) <= (inputs(97)) and not (inputs(254));
    layer0_outputs(692) <= inputs(156);
    layer0_outputs(693) <= not(inputs(37)) or (inputs(152));
    layer0_outputs(694) <= not((inputs(94)) and (inputs(145)));
    layer0_outputs(695) <= not((inputs(6)) and (inputs(57)));
    layer0_outputs(696) <= not(inputs(98)) or (inputs(186));
    layer0_outputs(697) <= (inputs(225)) or (inputs(228));
    layer0_outputs(698) <= (inputs(130)) and not (inputs(87));
    layer0_outputs(699) <= inputs(115);
    layer0_outputs(700) <= inputs(139);
    layer0_outputs(701) <= inputs(139);
    layer0_outputs(702) <= (inputs(71)) or (inputs(98));
    layer0_outputs(703) <= not(inputs(230));
    layer0_outputs(704) <= inputs(21);
    layer0_outputs(705) <= (inputs(234)) and (inputs(79));
    layer0_outputs(706) <= (inputs(85)) and not (inputs(145));
    layer0_outputs(707) <= not((inputs(111)) xor (inputs(254)));
    layer0_outputs(708) <= (inputs(6)) xor (inputs(78));
    layer0_outputs(709) <= not(inputs(254));
    layer0_outputs(710) <= inputs(74);
    layer0_outputs(711) <= '1';
    layer0_outputs(712) <= (inputs(246)) or (inputs(95));
    layer0_outputs(713) <= not(inputs(95));
    layer0_outputs(714) <= not((inputs(196)) or (inputs(134)));
    layer0_outputs(715) <= inputs(116);
    layer0_outputs(716) <= not((inputs(204)) or (inputs(253)));
    layer0_outputs(717) <= not((inputs(161)) or (inputs(244)));
    layer0_outputs(718) <= not(inputs(115));
    layer0_outputs(719) <= '1';
    layer0_outputs(720) <= inputs(151);
    layer0_outputs(721) <= (inputs(221)) or (inputs(228));
    layer0_outputs(722) <= not(inputs(134));
    layer0_outputs(723) <= not(inputs(153));
    layer0_outputs(724) <= (inputs(244)) or (inputs(248));
    layer0_outputs(725) <= not((inputs(148)) or (inputs(131)));
    layer0_outputs(726) <= inputs(95);
    layer0_outputs(727) <= not(inputs(217)) or (inputs(62));
    layer0_outputs(728) <= (inputs(250)) and not (inputs(79));
    layer0_outputs(729) <= inputs(46);
    layer0_outputs(730) <= not((inputs(164)) or (inputs(178)));
    layer0_outputs(731) <= (inputs(163)) and not (inputs(203));
    layer0_outputs(732) <= inputs(176);
    layer0_outputs(733) <= inputs(185);
    layer0_outputs(734) <= not(inputs(116)) or (inputs(71));
    layer0_outputs(735) <= not(inputs(212));
    layer0_outputs(736) <= (inputs(215)) and not (inputs(31));
    layer0_outputs(737) <= (inputs(251)) and not (inputs(152));
    layer0_outputs(738) <= inputs(164);
    layer0_outputs(739) <= '0';
    layer0_outputs(740) <= '0';
    layer0_outputs(741) <= (inputs(148)) and not (inputs(170));
    layer0_outputs(742) <= inputs(60);
    layer0_outputs(743) <= inputs(102);
    layer0_outputs(744) <= not((inputs(39)) or (inputs(214)));
    layer0_outputs(745) <= inputs(130);
    layer0_outputs(746) <= not(inputs(99));
    layer0_outputs(747) <= (inputs(107)) and not (inputs(194));
    layer0_outputs(748) <= not(inputs(157));
    layer0_outputs(749) <= (inputs(217)) or (inputs(165));
    layer0_outputs(750) <= (inputs(46)) or (inputs(52));
    layer0_outputs(751) <= not(inputs(131));
    layer0_outputs(752) <= not(inputs(235));
    layer0_outputs(753) <= not(inputs(23));
    layer0_outputs(754) <= not(inputs(157));
    layer0_outputs(755) <= (inputs(236)) or (inputs(105));
    layer0_outputs(756) <= not(inputs(92));
    layer0_outputs(757) <= inputs(77);
    layer0_outputs(758) <= inputs(180);
    layer0_outputs(759) <= not(inputs(88));
    layer0_outputs(760) <= '0';
    layer0_outputs(761) <= (inputs(25)) or (inputs(240));
    layer0_outputs(762) <= not(inputs(165));
    layer0_outputs(763) <= inputs(23);
    layer0_outputs(764) <= (inputs(100)) and not (inputs(141));
    layer0_outputs(765) <= not(inputs(69)) or (inputs(162));
    layer0_outputs(766) <= not(inputs(120));
    layer0_outputs(767) <= not(inputs(200));
    layer0_outputs(768) <= inputs(131);
    layer0_outputs(769) <= not(inputs(161));
    layer0_outputs(770) <= not(inputs(208));
    layer0_outputs(771) <= not(inputs(197));
    layer0_outputs(772) <= inputs(212);
    layer0_outputs(773) <= not(inputs(16)) or (inputs(65));
    layer0_outputs(774) <= inputs(85);
    layer0_outputs(775) <= not(inputs(65)) or (inputs(91));
    layer0_outputs(776) <= not((inputs(5)) and (inputs(7)));
    layer0_outputs(777) <= not(inputs(201));
    layer0_outputs(778) <= (inputs(153)) and not (inputs(136));
    layer0_outputs(779) <= inputs(237);
    layer0_outputs(780) <= not(inputs(226));
    layer0_outputs(781) <= (inputs(134)) and (inputs(167));
    layer0_outputs(782) <= not((inputs(126)) or (inputs(247)));
    layer0_outputs(783) <= (inputs(84)) and not (inputs(35));
    layer0_outputs(784) <= not((inputs(34)) or (inputs(187)));
    layer0_outputs(785) <= inputs(94);
    layer0_outputs(786) <= inputs(239);
    layer0_outputs(787) <= not((inputs(106)) or (inputs(183)));
    layer0_outputs(788) <= (inputs(203)) or (inputs(219));
    layer0_outputs(789) <= (inputs(125)) and not (inputs(120));
    layer0_outputs(790) <= (inputs(232)) and not (inputs(30));
    layer0_outputs(791) <= inputs(120);
    layer0_outputs(792) <= (inputs(83)) or (inputs(249));
    layer0_outputs(793) <= inputs(177);
    layer0_outputs(794) <= not((inputs(119)) or (inputs(166)));
    layer0_outputs(795) <= inputs(126);
    layer0_outputs(796) <= (inputs(4)) and (inputs(92));
    layer0_outputs(797) <= not(inputs(21));
    layer0_outputs(798) <= not(inputs(194));
    layer0_outputs(799) <= inputs(182);
    layer0_outputs(800) <= (inputs(3)) or (inputs(30));
    layer0_outputs(801) <= inputs(18);
    layer0_outputs(802) <= not((inputs(125)) or (inputs(90)));
    layer0_outputs(803) <= not(inputs(206));
    layer0_outputs(804) <= not(inputs(89));
    layer0_outputs(805) <= inputs(166);
    layer0_outputs(806) <= not(inputs(59));
    layer0_outputs(807) <= '0';
    layer0_outputs(808) <= not(inputs(21)) or (inputs(190));
    layer0_outputs(809) <= inputs(121);
    layer0_outputs(810) <= not(inputs(233));
    layer0_outputs(811) <= inputs(254);
    layer0_outputs(812) <= '0';
    layer0_outputs(813) <= not(inputs(89)) or (inputs(99));
    layer0_outputs(814) <= inputs(32);
    layer0_outputs(815) <= (inputs(208)) or (inputs(222));
    layer0_outputs(816) <= not((inputs(201)) or (inputs(148)));
    layer0_outputs(817) <= '0';
    layer0_outputs(818) <= not(inputs(106));
    layer0_outputs(819) <= not((inputs(116)) or (inputs(206)));
    layer0_outputs(820) <= (inputs(82)) and (inputs(82));
    layer0_outputs(821) <= inputs(201);
    layer0_outputs(822) <= not(inputs(36));
    layer0_outputs(823) <= inputs(246);
    layer0_outputs(824) <= '1';
    layer0_outputs(825) <= not(inputs(182));
    layer0_outputs(826) <= inputs(32);
    layer0_outputs(827) <= not((inputs(87)) or (inputs(203)));
    layer0_outputs(828) <= not(inputs(164));
    layer0_outputs(829) <= inputs(110);
    layer0_outputs(830) <= '0';
    layer0_outputs(831) <= not((inputs(7)) xor (inputs(65)));
    layer0_outputs(832) <= '1';
    layer0_outputs(833) <= (inputs(95)) or (inputs(38));
    layer0_outputs(834) <= not(inputs(197)) or (inputs(175));
    layer0_outputs(835) <= not((inputs(53)) or (inputs(210)));
    layer0_outputs(836) <= not(inputs(230));
    layer0_outputs(837) <= not(inputs(107));
    layer0_outputs(838) <= (inputs(215)) and (inputs(240));
    layer0_outputs(839) <= not(inputs(186)) or (inputs(86));
    layer0_outputs(840) <= (inputs(139)) xor (inputs(149));
    layer0_outputs(841) <= (inputs(76)) and not (inputs(152));
    layer0_outputs(842) <= inputs(171);
    layer0_outputs(843) <= inputs(155);
    layer0_outputs(844) <= not((inputs(206)) xor (inputs(79)));
    layer0_outputs(845) <= not((inputs(7)) or (inputs(193)));
    layer0_outputs(846) <= not(inputs(39));
    layer0_outputs(847) <= inputs(6);
    layer0_outputs(848) <= (inputs(121)) and (inputs(234));
    layer0_outputs(849) <= (inputs(158)) or (inputs(111));
    layer0_outputs(850) <= not(inputs(98));
    layer0_outputs(851) <= not((inputs(168)) or (inputs(238)));
    layer0_outputs(852) <= (inputs(136)) and not (inputs(131));
    layer0_outputs(853) <= not(inputs(109)) or (inputs(129));
    layer0_outputs(854) <= not(inputs(166));
    layer0_outputs(855) <= not((inputs(50)) or (inputs(206)));
    layer0_outputs(856) <= (inputs(162)) or (inputs(253));
    layer0_outputs(857) <= inputs(109);
    layer0_outputs(858) <= not(inputs(149));
    layer0_outputs(859) <= not(inputs(145)) or (inputs(105));
    layer0_outputs(860) <= inputs(77);
    layer0_outputs(861) <= not(inputs(12));
    layer0_outputs(862) <= not(inputs(84));
    layer0_outputs(863) <= inputs(133);
    layer0_outputs(864) <= (inputs(91)) and not (inputs(193));
    layer0_outputs(865) <= not(inputs(93)) or (inputs(238));
    layer0_outputs(866) <= inputs(229);
    layer0_outputs(867) <= not(inputs(200));
    layer0_outputs(868) <= (inputs(221)) and not (inputs(101));
    layer0_outputs(869) <= not((inputs(67)) or (inputs(113)));
    layer0_outputs(870) <= (inputs(172)) xor (inputs(238));
    layer0_outputs(871) <= inputs(178);
    layer0_outputs(872) <= (inputs(52)) and not (inputs(221));
    layer0_outputs(873) <= inputs(199);
    layer0_outputs(874) <= inputs(224);
    layer0_outputs(875) <= not((inputs(175)) xor (inputs(45)));
    layer0_outputs(876) <= not((inputs(38)) and (inputs(220)));
    layer0_outputs(877) <= inputs(243);
    layer0_outputs(878) <= inputs(21);
    layer0_outputs(879) <= '1';
    layer0_outputs(880) <= inputs(107);
    layer0_outputs(881) <= inputs(137);
    layer0_outputs(882) <= inputs(247);
    layer0_outputs(883) <= '1';
    layer0_outputs(884) <= (inputs(38)) and not (inputs(198));
    layer0_outputs(885) <= not((inputs(127)) or (inputs(75)));
    layer0_outputs(886) <= '0';
    layer0_outputs(887) <= inputs(113);
    layer0_outputs(888) <= not((inputs(163)) or (inputs(31)));
    layer0_outputs(889) <= not(inputs(184));
    layer0_outputs(890) <= (inputs(192)) or (inputs(216));
    layer0_outputs(891) <= not(inputs(33)) or (inputs(81));
    layer0_outputs(892) <= not(inputs(120));
    layer0_outputs(893) <= inputs(103);
    layer0_outputs(894) <= (inputs(189)) or (inputs(156));
    layer0_outputs(895) <= not(inputs(67));
    layer0_outputs(896) <= (inputs(167)) and not (inputs(98));
    layer0_outputs(897) <= (inputs(197)) and not (inputs(68));
    layer0_outputs(898) <= not(inputs(151));
    layer0_outputs(899) <= not((inputs(218)) or (inputs(140)));
    layer0_outputs(900) <= (inputs(103)) or (inputs(116));
    layer0_outputs(901) <= (inputs(163)) or (inputs(54));
    layer0_outputs(902) <= inputs(113);
    layer0_outputs(903) <= not((inputs(171)) or (inputs(161)));
    layer0_outputs(904) <= not(inputs(210)) or (inputs(60));
    layer0_outputs(905) <= (inputs(244)) or (inputs(129));
    layer0_outputs(906) <= (inputs(124)) and (inputs(29));
    layer0_outputs(907) <= inputs(97);
    layer0_outputs(908) <= not((inputs(147)) or (inputs(36)));
    layer0_outputs(909) <= (inputs(214)) and not (inputs(98));
    layer0_outputs(910) <= (inputs(192)) or (inputs(185));
    layer0_outputs(911) <= not((inputs(78)) and (inputs(46)));
    layer0_outputs(912) <= inputs(83);
    layer0_outputs(913) <= (inputs(154)) or (inputs(93));
    layer0_outputs(914) <= not((inputs(52)) or (inputs(80)));
    layer0_outputs(915) <= (inputs(120)) or (inputs(151));
    layer0_outputs(916) <= inputs(24);
    layer0_outputs(917) <= (inputs(143)) or (inputs(188));
    layer0_outputs(918) <= not(inputs(179)) or (inputs(239));
    layer0_outputs(919) <= not((inputs(139)) or (inputs(207)));
    layer0_outputs(920) <= inputs(239);
    layer0_outputs(921) <= not(inputs(171)) or (inputs(31));
    layer0_outputs(922) <= not(inputs(117));
    layer0_outputs(923) <= '0';
    layer0_outputs(924) <= '1';
    layer0_outputs(925) <= not(inputs(7));
    layer0_outputs(926) <= (inputs(209)) or (inputs(41));
    layer0_outputs(927) <= not(inputs(66)) or (inputs(55));
    layer0_outputs(928) <= '1';
    layer0_outputs(929) <= inputs(245);
    layer0_outputs(930) <= not(inputs(49)) or (inputs(183));
    layer0_outputs(931) <= not((inputs(115)) xor (inputs(102)));
    layer0_outputs(932) <= inputs(115);
    layer0_outputs(933) <= not(inputs(177));
    layer0_outputs(934) <= inputs(42);
    layer0_outputs(935) <= (inputs(206)) or (inputs(255));
    layer0_outputs(936) <= not((inputs(20)) xor (inputs(253)));
    layer0_outputs(937) <= not((inputs(101)) or (inputs(215)));
    layer0_outputs(938) <= not((inputs(220)) or (inputs(239)));
    layer0_outputs(939) <= not(inputs(181));
    layer0_outputs(940) <= inputs(142);
    layer0_outputs(941) <= (inputs(187)) or (inputs(160));
    layer0_outputs(942) <= not(inputs(4));
    layer0_outputs(943) <= not(inputs(151)) or (inputs(109));
    layer0_outputs(944) <= (inputs(220)) and (inputs(212));
    layer0_outputs(945) <= inputs(175);
    layer0_outputs(946) <= (inputs(230)) or (inputs(106));
    layer0_outputs(947) <= not(inputs(139)) or (inputs(237));
    layer0_outputs(948) <= not(inputs(22)) or (inputs(17));
    layer0_outputs(949) <= (inputs(10)) or (inputs(79));
    layer0_outputs(950) <= inputs(27);
    layer0_outputs(951) <= not((inputs(1)) and (inputs(109)));
    layer0_outputs(952) <= not((inputs(32)) or (inputs(131)));
    layer0_outputs(953) <= not((inputs(169)) xor (inputs(16)));
    layer0_outputs(954) <= not(inputs(104));
    layer0_outputs(955) <= inputs(107);
    layer0_outputs(956) <= not((inputs(111)) or (inputs(118)));
    layer0_outputs(957) <= not(inputs(153));
    layer0_outputs(958) <= '0';
    layer0_outputs(959) <= '1';
    layer0_outputs(960) <= not(inputs(151));
    layer0_outputs(961) <= not((inputs(63)) or (inputs(210)));
    layer0_outputs(962) <= not(inputs(116));
    layer0_outputs(963) <= (inputs(192)) or (inputs(203));
    layer0_outputs(964) <= inputs(179);
    layer0_outputs(965) <= not(inputs(50));
    layer0_outputs(966) <= not(inputs(145));
    layer0_outputs(967) <= (inputs(19)) and (inputs(37));
    layer0_outputs(968) <= inputs(41);
    layer0_outputs(969) <= (inputs(30)) or (inputs(253));
    layer0_outputs(970) <= not(inputs(231));
    layer0_outputs(971) <= '1';
    layer0_outputs(972) <= not(inputs(16));
    layer0_outputs(973) <= not(inputs(26)) or (inputs(127));
    layer0_outputs(974) <= not(inputs(90));
    layer0_outputs(975) <= (inputs(205)) and (inputs(102));
    layer0_outputs(976) <= (inputs(19)) or (inputs(90));
    layer0_outputs(977) <= inputs(74);
    layer0_outputs(978) <= (inputs(176)) xor (inputs(233));
    layer0_outputs(979) <= (inputs(239)) or (inputs(135));
    layer0_outputs(980) <= not(inputs(23));
    layer0_outputs(981) <= not((inputs(255)) or (inputs(193)));
    layer0_outputs(982) <= (inputs(175)) and not (inputs(33));
    layer0_outputs(983) <= not(inputs(215));
    layer0_outputs(984) <= '1';
    layer0_outputs(985) <= not(inputs(77));
    layer0_outputs(986) <= not((inputs(144)) or (inputs(97)));
    layer0_outputs(987) <= '1';
    layer0_outputs(988) <= not((inputs(0)) xor (inputs(112)));
    layer0_outputs(989) <= (inputs(13)) and not (inputs(254));
    layer0_outputs(990) <= not(inputs(34));
    layer0_outputs(991) <= not(inputs(196));
    layer0_outputs(992) <= not(inputs(220)) or (inputs(110));
    layer0_outputs(993) <= (inputs(176)) or (inputs(92));
    layer0_outputs(994) <= not(inputs(24)) or (inputs(18));
    layer0_outputs(995) <= not(inputs(204)) or (inputs(65));
    layer0_outputs(996) <= inputs(189);
    layer0_outputs(997) <= not((inputs(56)) and (inputs(70)));
    layer0_outputs(998) <= not(inputs(233));
    layer0_outputs(999) <= not(inputs(216));
    layer0_outputs(1000) <= (inputs(7)) and not (inputs(248));
    layer0_outputs(1001) <= not(inputs(144)) or (inputs(15));
    layer0_outputs(1002) <= not(inputs(104)) or (inputs(147));
    layer0_outputs(1003) <= '0';
    layer0_outputs(1004) <= inputs(100);
    layer0_outputs(1005) <= (inputs(94)) and not (inputs(123));
    layer0_outputs(1006) <= not(inputs(2));
    layer0_outputs(1007) <= (inputs(59)) and (inputs(0));
    layer0_outputs(1008) <= not(inputs(220));
    layer0_outputs(1009) <= not(inputs(17));
    layer0_outputs(1010) <= (inputs(18)) and not (inputs(129));
    layer0_outputs(1011) <= (inputs(253)) xor (inputs(241));
    layer0_outputs(1012) <= inputs(120);
    layer0_outputs(1013) <= not((inputs(211)) xor (inputs(31)));
    layer0_outputs(1014) <= (inputs(212)) and (inputs(238));
    layer0_outputs(1015) <= not(inputs(27));
    layer0_outputs(1016) <= inputs(245);
    layer0_outputs(1017) <= (inputs(7)) or (inputs(40));
    layer0_outputs(1018) <= (inputs(97)) and not (inputs(237));
    layer0_outputs(1019) <= not(inputs(69));
    layer0_outputs(1020) <= '0';
    layer0_outputs(1021) <= not((inputs(154)) or (inputs(67)));
    layer0_outputs(1022) <= (inputs(238)) or (inputs(181));
    layer0_outputs(1023) <= '1';
    layer0_outputs(1024) <= (inputs(208)) or (inputs(18));
    layer0_outputs(1025) <= (inputs(197)) xor (inputs(194));
    layer0_outputs(1026) <= '0';
    layer0_outputs(1027) <= not((inputs(22)) and (inputs(26)));
    layer0_outputs(1028) <= inputs(181);
    layer0_outputs(1029) <= not(inputs(165)) or (inputs(143));
    layer0_outputs(1030) <= '1';
    layer0_outputs(1031) <= not(inputs(26));
    layer0_outputs(1032) <= not(inputs(203)) or (inputs(29));
    layer0_outputs(1033) <= not(inputs(20));
    layer0_outputs(1034) <= (inputs(105)) and not (inputs(115));
    layer0_outputs(1035) <= '1';
    layer0_outputs(1036) <= inputs(76);
    layer0_outputs(1037) <= not(inputs(25));
    layer0_outputs(1038) <= inputs(161);
    layer0_outputs(1039) <= inputs(163);
    layer0_outputs(1040) <= not((inputs(247)) or (inputs(99)));
    layer0_outputs(1041) <= not((inputs(86)) or (inputs(96)));
    layer0_outputs(1042) <= not(inputs(85));
    layer0_outputs(1043) <= not((inputs(248)) and (inputs(180)));
    layer0_outputs(1044) <= not(inputs(155)) or (inputs(154));
    layer0_outputs(1045) <= not(inputs(84));
    layer0_outputs(1046) <= '1';
    layer0_outputs(1047) <= inputs(52);
    layer0_outputs(1048) <= not(inputs(167));
    layer0_outputs(1049) <= inputs(165);
    layer0_outputs(1050) <= (inputs(188)) or (inputs(54));
    layer0_outputs(1051) <= not(inputs(10)) or (inputs(33));
    layer0_outputs(1052) <= (inputs(159)) or (inputs(96));
    layer0_outputs(1053) <= not(inputs(232)) or (inputs(243));
    layer0_outputs(1054) <= (inputs(172)) and not (inputs(234));
    layer0_outputs(1055) <= '1';
    layer0_outputs(1056) <= not(inputs(196)) or (inputs(241));
    layer0_outputs(1057) <= not(inputs(106));
    layer0_outputs(1058) <= '1';
    layer0_outputs(1059) <= not(inputs(128));
    layer0_outputs(1060) <= (inputs(155)) and not (inputs(110));
    layer0_outputs(1061) <= '0';
    layer0_outputs(1062) <= (inputs(113)) or (inputs(219));
    layer0_outputs(1063) <= (inputs(5)) and not (inputs(119));
    layer0_outputs(1064) <= not((inputs(196)) or (inputs(94)));
    layer0_outputs(1065) <= not(inputs(219));
    layer0_outputs(1066) <= not((inputs(29)) or (inputs(31)));
    layer0_outputs(1067) <= not((inputs(111)) or (inputs(171)));
    layer0_outputs(1068) <= not(inputs(60)) or (inputs(220));
    layer0_outputs(1069) <= not((inputs(140)) and (inputs(137)));
    layer0_outputs(1070) <= not((inputs(162)) or (inputs(121)));
    layer0_outputs(1071) <= (inputs(44)) and (inputs(14));
    layer0_outputs(1072) <= not(inputs(90)) or (inputs(57));
    layer0_outputs(1073) <= not((inputs(239)) and (inputs(65)));
    layer0_outputs(1074) <= (inputs(193)) or (inputs(235));
    layer0_outputs(1075) <= inputs(170);
    layer0_outputs(1076) <= (inputs(16)) and (inputs(218));
    layer0_outputs(1077) <= (inputs(136)) and not (inputs(48));
    layer0_outputs(1078) <= not((inputs(240)) xor (inputs(27)));
    layer0_outputs(1079) <= not(inputs(142));
    layer0_outputs(1080) <= not((inputs(26)) and (inputs(91)));
    layer0_outputs(1081) <= not(inputs(147)) or (inputs(13));
    layer0_outputs(1082) <= (inputs(250)) or (inputs(255));
    layer0_outputs(1083) <= not(inputs(232));
    layer0_outputs(1084) <= (inputs(88)) and not (inputs(219));
    layer0_outputs(1085) <= (inputs(227)) and not (inputs(57));
    layer0_outputs(1086) <= not((inputs(194)) or (inputs(211)));
    layer0_outputs(1087) <= (inputs(20)) and not (inputs(146));
    layer0_outputs(1088) <= '1';
    layer0_outputs(1089) <= not(inputs(66));
    layer0_outputs(1090) <= not(inputs(21));
    layer0_outputs(1091) <= not(inputs(67));
    layer0_outputs(1092) <= inputs(20);
    layer0_outputs(1093) <= (inputs(223)) xor (inputs(139));
    layer0_outputs(1094) <= (inputs(26)) and not (inputs(230));
    layer0_outputs(1095) <= (inputs(212)) and (inputs(200));
    layer0_outputs(1096) <= (inputs(210)) or (inputs(0));
    layer0_outputs(1097) <= not(inputs(187));
    layer0_outputs(1098) <= inputs(126);
    layer0_outputs(1099) <= not((inputs(226)) or (inputs(211)));
    layer0_outputs(1100) <= not(inputs(110));
    layer0_outputs(1101) <= inputs(185);
    layer0_outputs(1102) <= not(inputs(169));
    layer0_outputs(1103) <= not(inputs(141)) or (inputs(138));
    layer0_outputs(1104) <= (inputs(178)) or (inputs(135));
    layer0_outputs(1105) <= '1';
    layer0_outputs(1106) <= not((inputs(78)) or (inputs(24)));
    layer0_outputs(1107) <= not(inputs(191)) or (inputs(112));
    layer0_outputs(1108) <= '1';
    layer0_outputs(1109) <= inputs(171);
    layer0_outputs(1110) <= (inputs(18)) or (inputs(244));
    layer0_outputs(1111) <= (inputs(150)) or (inputs(194));
    layer0_outputs(1112) <= '0';
    layer0_outputs(1113) <= (inputs(53)) or (inputs(9));
    layer0_outputs(1114) <= not(inputs(204)) or (inputs(204));
    layer0_outputs(1115) <= not((inputs(175)) or (inputs(227)));
    layer0_outputs(1116) <= inputs(228);
    layer0_outputs(1117) <= '1';
    layer0_outputs(1118) <= (inputs(4)) xor (inputs(160));
    layer0_outputs(1119) <= not(inputs(173));
    layer0_outputs(1120) <= (inputs(81)) and not (inputs(103));
    layer0_outputs(1121) <= inputs(154);
    layer0_outputs(1122) <= inputs(150);
    layer0_outputs(1123) <= not(inputs(101));
    layer0_outputs(1124) <= inputs(163);
    layer0_outputs(1125) <= (inputs(145)) or (inputs(111));
    layer0_outputs(1126) <= not((inputs(114)) xor (inputs(12)));
    layer0_outputs(1127) <= not((inputs(230)) or (inputs(188)));
    layer0_outputs(1128) <= '0';
    layer0_outputs(1129) <= inputs(166);
    layer0_outputs(1130) <= (inputs(93)) and not (inputs(126));
    layer0_outputs(1131) <= (inputs(85)) or (inputs(207));
    layer0_outputs(1132) <= not((inputs(2)) and (inputs(37)));
    layer0_outputs(1133) <= not(inputs(164));
    layer0_outputs(1134) <= inputs(103);
    layer0_outputs(1135) <= not(inputs(248)) or (inputs(95));
    layer0_outputs(1136) <= '0';
    layer0_outputs(1137) <= inputs(234);
    layer0_outputs(1138) <= (inputs(125)) and not (inputs(39));
    layer0_outputs(1139) <= not(inputs(185)) or (inputs(43));
    layer0_outputs(1140) <= (inputs(145)) and not (inputs(155));
    layer0_outputs(1141) <= '0';
    layer0_outputs(1142) <= not(inputs(51));
    layer0_outputs(1143) <= not(inputs(13)) or (inputs(74));
    layer0_outputs(1144) <= not((inputs(156)) xor (inputs(240)));
    layer0_outputs(1145) <= not((inputs(16)) or (inputs(209)));
    layer0_outputs(1146) <= not((inputs(227)) xor (inputs(142)));
    layer0_outputs(1147) <= not(inputs(194));
    layer0_outputs(1148) <= inputs(152);
    layer0_outputs(1149) <= inputs(80);
    layer0_outputs(1150) <= not(inputs(87));
    layer0_outputs(1151) <= not(inputs(214)) or (inputs(45));
    layer0_outputs(1152) <= not(inputs(172));
    layer0_outputs(1153) <= not(inputs(228));
    layer0_outputs(1154) <= '0';
    layer0_outputs(1155) <= '0';
    layer0_outputs(1156) <= inputs(226);
    layer0_outputs(1157) <= not(inputs(133)) or (inputs(2));
    layer0_outputs(1158) <= not((inputs(221)) or (inputs(211)));
    layer0_outputs(1159) <= inputs(248);
    layer0_outputs(1160) <= not(inputs(77));
    layer0_outputs(1161) <= not(inputs(248));
    layer0_outputs(1162) <= not(inputs(167));
    layer0_outputs(1163) <= inputs(181);
    layer0_outputs(1164) <= not(inputs(38));
    layer0_outputs(1165) <= not((inputs(192)) or (inputs(129)));
    layer0_outputs(1166) <= inputs(196);
    layer0_outputs(1167) <= not(inputs(100));
    layer0_outputs(1168) <= not(inputs(151)) or (inputs(243));
    layer0_outputs(1169) <= (inputs(58)) and not (inputs(150));
    layer0_outputs(1170) <= (inputs(169)) and not (inputs(9));
    layer0_outputs(1171) <= '0';
    layer0_outputs(1172) <= (inputs(212)) or (inputs(186));
    layer0_outputs(1173) <= inputs(178);
    layer0_outputs(1174) <= '1';
    layer0_outputs(1175) <= (inputs(207)) and not (inputs(159));
    layer0_outputs(1176) <= (inputs(218)) or (inputs(206));
    layer0_outputs(1177) <= not((inputs(247)) and (inputs(149)));
    layer0_outputs(1178) <= not(inputs(120)) or (inputs(192));
    layer0_outputs(1179) <= not(inputs(233)) or (inputs(35));
    layer0_outputs(1180) <= (inputs(242)) and not (inputs(56));
    layer0_outputs(1181) <= inputs(83);
    layer0_outputs(1182) <= not(inputs(144));
    layer0_outputs(1183) <= not((inputs(59)) and (inputs(183)));
    layer0_outputs(1184) <= not(inputs(113));
    layer0_outputs(1185) <= not(inputs(112));
    layer0_outputs(1186) <= (inputs(238)) and not (inputs(124));
    layer0_outputs(1187) <= not(inputs(193)) or (inputs(167));
    layer0_outputs(1188) <= inputs(84);
    layer0_outputs(1189) <= '0';
    layer0_outputs(1190) <= inputs(117);
    layer0_outputs(1191) <= (inputs(88)) and not (inputs(160));
    layer0_outputs(1192) <= '1';
    layer0_outputs(1193) <= not(inputs(226));
    layer0_outputs(1194) <= (inputs(250)) and not (inputs(148));
    layer0_outputs(1195) <= not(inputs(197)) or (inputs(1));
    layer0_outputs(1196) <= not(inputs(103));
    layer0_outputs(1197) <= inputs(193);
    layer0_outputs(1198) <= not(inputs(40));
    layer0_outputs(1199) <= not(inputs(93)) or (inputs(106));
    layer0_outputs(1200) <= inputs(111);
    layer0_outputs(1201) <= (inputs(113)) or (inputs(63));
    layer0_outputs(1202) <= (inputs(227)) xor (inputs(181));
    layer0_outputs(1203) <= '1';
    layer0_outputs(1204) <= not((inputs(163)) or (inputs(204)));
    layer0_outputs(1205) <= not(inputs(77));
    layer0_outputs(1206) <= not(inputs(254)) or (inputs(161));
    layer0_outputs(1207) <= not((inputs(125)) or (inputs(134)));
    layer0_outputs(1208) <= inputs(231);
    layer0_outputs(1209) <= (inputs(82)) or (inputs(149));
    layer0_outputs(1210) <= (inputs(22)) and not (inputs(112));
    layer0_outputs(1211) <= (inputs(14)) or (inputs(101));
    layer0_outputs(1212) <= (inputs(51)) or (inputs(251));
    layer0_outputs(1213) <= not(inputs(105));
    layer0_outputs(1214) <= not(inputs(62));
    layer0_outputs(1215) <= inputs(77);
    layer0_outputs(1216) <= (inputs(47)) and not (inputs(128));
    layer0_outputs(1217) <= (inputs(198)) or (inputs(229));
    layer0_outputs(1218) <= (inputs(187)) or (inputs(148));
    layer0_outputs(1219) <= not((inputs(191)) or (inputs(246)));
    layer0_outputs(1220) <= not((inputs(175)) or (inputs(171)));
    layer0_outputs(1221) <= not(inputs(160));
    layer0_outputs(1222) <= not(inputs(99)) or (inputs(15));
    layer0_outputs(1223) <= (inputs(69)) and not (inputs(126));
    layer0_outputs(1224) <= (inputs(9)) xor (inputs(3));
    layer0_outputs(1225) <= not(inputs(164));
    layer0_outputs(1226) <= (inputs(30)) and not (inputs(191));
    layer0_outputs(1227) <= not(inputs(56)) or (inputs(125));
    layer0_outputs(1228) <= not(inputs(24)) or (inputs(163));
    layer0_outputs(1229) <= not(inputs(194));
    layer0_outputs(1230) <= (inputs(35)) or (inputs(32));
    layer0_outputs(1231) <= not((inputs(172)) or (inputs(98)));
    layer0_outputs(1232) <= not(inputs(24)) or (inputs(225));
    layer0_outputs(1233) <= not((inputs(190)) xor (inputs(139)));
    layer0_outputs(1234) <= inputs(164);
    layer0_outputs(1235) <= '1';
    layer0_outputs(1236) <= not(inputs(145)) or (inputs(198));
    layer0_outputs(1237) <= inputs(151);
    layer0_outputs(1238) <= not(inputs(163));
    layer0_outputs(1239) <= '0';
    layer0_outputs(1240) <= (inputs(18)) xor (inputs(113));
    layer0_outputs(1241) <= not((inputs(98)) xor (inputs(202)));
    layer0_outputs(1242) <= not((inputs(173)) or (inputs(215)));
    layer0_outputs(1243) <= (inputs(199)) and (inputs(162));
    layer0_outputs(1244) <= not(inputs(113));
    layer0_outputs(1245) <= (inputs(195)) or (inputs(149));
    layer0_outputs(1246) <= inputs(24);
    layer0_outputs(1247) <= not(inputs(205)) or (inputs(50));
    layer0_outputs(1248) <= inputs(183);
    layer0_outputs(1249) <= (inputs(78)) or (inputs(194));
    layer0_outputs(1250) <= inputs(100);
    layer0_outputs(1251) <= inputs(161);
    layer0_outputs(1252) <= not(inputs(140)) or (inputs(205));
    layer0_outputs(1253) <= inputs(154);
    layer0_outputs(1254) <= not(inputs(75));
    layer0_outputs(1255) <= (inputs(35)) and not (inputs(81));
    layer0_outputs(1256) <= inputs(157);
    layer0_outputs(1257) <= inputs(112);
    layer0_outputs(1258) <= not(inputs(166));
    layer0_outputs(1259) <= '0';
    layer0_outputs(1260) <= not(inputs(187)) or (inputs(146));
    layer0_outputs(1261) <= not(inputs(209));
    layer0_outputs(1262) <= (inputs(128)) or (inputs(189));
    layer0_outputs(1263) <= not((inputs(180)) or (inputs(32)));
    layer0_outputs(1264) <= not(inputs(154));
    layer0_outputs(1265) <= (inputs(1)) and (inputs(243));
    layer0_outputs(1266) <= inputs(84);
    layer0_outputs(1267) <= not(inputs(29));
    layer0_outputs(1268) <= not((inputs(53)) or (inputs(52)));
    layer0_outputs(1269) <= not(inputs(104));
    layer0_outputs(1270) <= inputs(105);
    layer0_outputs(1271) <= not((inputs(235)) xor (inputs(175)));
    layer0_outputs(1272) <= (inputs(77)) or (inputs(8));
    layer0_outputs(1273) <= inputs(44);
    layer0_outputs(1274) <= not((inputs(108)) and (inputs(228)));
    layer0_outputs(1275) <= (inputs(231)) and not (inputs(138));
    layer0_outputs(1276) <= not((inputs(64)) and (inputs(86)));
    layer0_outputs(1277) <= inputs(132);
    layer0_outputs(1278) <= (inputs(213)) or (inputs(233));
    layer0_outputs(1279) <= not((inputs(214)) or (inputs(208)));
    layer0_outputs(1280) <= '1';
    layer0_outputs(1281) <= not((inputs(128)) and (inputs(49)));
    layer0_outputs(1282) <= (inputs(241)) and (inputs(184));
    layer0_outputs(1283) <= not(inputs(170)) or (inputs(124));
    layer0_outputs(1284) <= inputs(76);
    layer0_outputs(1285) <= (inputs(85)) and not (inputs(93));
    layer0_outputs(1286) <= not((inputs(154)) and (inputs(9)));
    layer0_outputs(1287) <= (inputs(228)) and (inputs(114));
    layer0_outputs(1288) <= not((inputs(225)) or (inputs(223)));
    layer0_outputs(1289) <= not(inputs(168));
    layer0_outputs(1290) <= not(inputs(193)) or (inputs(161));
    layer0_outputs(1291) <= inputs(146);
    layer0_outputs(1292) <= (inputs(61)) and not (inputs(11));
    layer0_outputs(1293) <= not(inputs(22));
    layer0_outputs(1294) <= '0';
    layer0_outputs(1295) <= (inputs(153)) and (inputs(144));
    layer0_outputs(1296) <= not(inputs(36));
    layer0_outputs(1297) <= inputs(116);
    layer0_outputs(1298) <= not((inputs(249)) xor (inputs(217)));
    layer0_outputs(1299) <= not(inputs(53));
    layer0_outputs(1300) <= (inputs(242)) or (inputs(132));
    layer0_outputs(1301) <= not((inputs(217)) or (inputs(248)));
    layer0_outputs(1302) <= (inputs(130)) and (inputs(142));
    layer0_outputs(1303) <= '0';
    layer0_outputs(1304) <= not((inputs(3)) and (inputs(24)));
    layer0_outputs(1305) <= not((inputs(129)) or (inputs(22)));
    layer0_outputs(1306) <= '1';
    layer0_outputs(1307) <= inputs(193);
    layer0_outputs(1308) <= inputs(230);
    layer0_outputs(1309) <= not(inputs(141));
    layer0_outputs(1310) <= (inputs(9)) and not (inputs(144));
    layer0_outputs(1311) <= inputs(112);
    layer0_outputs(1312) <= (inputs(62)) and not (inputs(128));
    layer0_outputs(1313) <= inputs(25);
    layer0_outputs(1314) <= inputs(135);
    layer0_outputs(1315) <= inputs(56);
    layer0_outputs(1316) <= (inputs(84)) and not (inputs(210));
    layer0_outputs(1317) <= not((inputs(126)) or (inputs(146)));
    layer0_outputs(1318) <= (inputs(122)) or (inputs(74));
    layer0_outputs(1319) <= not(inputs(28)) or (inputs(184));
    layer0_outputs(1320) <= not(inputs(2));
    layer0_outputs(1321) <= not(inputs(27));
    layer0_outputs(1322) <= (inputs(179)) or (inputs(60));
    layer0_outputs(1323) <= inputs(222);
    layer0_outputs(1324) <= not(inputs(146)) or (inputs(224));
    layer0_outputs(1325) <= not((inputs(154)) and (inputs(166)));
    layer0_outputs(1326) <= not(inputs(238)) or (inputs(45));
    layer0_outputs(1327) <= not(inputs(107));
    layer0_outputs(1328) <= not(inputs(22)) or (inputs(173));
    layer0_outputs(1329) <= (inputs(171)) or (inputs(13));
    layer0_outputs(1330) <= inputs(141);
    layer0_outputs(1331) <= not((inputs(242)) or (inputs(192)));
    layer0_outputs(1332) <= not(inputs(44));
    layer0_outputs(1333) <= (inputs(34)) or (inputs(60));
    layer0_outputs(1334) <= '0';
    layer0_outputs(1335) <= not(inputs(94));
    layer0_outputs(1336) <= not((inputs(123)) or (inputs(89)));
    layer0_outputs(1337) <= not(inputs(132)) or (inputs(254));
    layer0_outputs(1338) <= (inputs(3)) or (inputs(29));
    layer0_outputs(1339) <= (inputs(6)) or (inputs(93));
    layer0_outputs(1340) <= not(inputs(183));
    layer0_outputs(1341) <= not((inputs(6)) or (inputs(72)));
    layer0_outputs(1342) <= not(inputs(107));
    layer0_outputs(1343) <= not(inputs(109)) or (inputs(243));
    layer0_outputs(1344) <= not(inputs(204));
    layer0_outputs(1345) <= (inputs(233)) and not (inputs(54));
    layer0_outputs(1346) <= inputs(68);
    layer0_outputs(1347) <= not(inputs(71)) or (inputs(252));
    layer0_outputs(1348) <= inputs(50);
    layer0_outputs(1349) <= '0';
    layer0_outputs(1350) <= not(inputs(165));
    layer0_outputs(1351) <= (inputs(198)) and not (inputs(209));
    layer0_outputs(1352) <= not(inputs(12)) or (inputs(210));
    layer0_outputs(1353) <= inputs(75);
    layer0_outputs(1354) <= not(inputs(185)) or (inputs(81));
    layer0_outputs(1355) <= '0';
    layer0_outputs(1356) <= not(inputs(230)) or (inputs(165));
    layer0_outputs(1357) <= not(inputs(79)) or (inputs(185));
    layer0_outputs(1358) <= (inputs(121)) and not (inputs(11));
    layer0_outputs(1359) <= not(inputs(131));
    layer0_outputs(1360) <= inputs(103);
    layer0_outputs(1361) <= inputs(104);
    layer0_outputs(1362) <= not((inputs(82)) and (inputs(153)));
    layer0_outputs(1363) <= (inputs(240)) and (inputs(244));
    layer0_outputs(1364) <= not((inputs(99)) xor (inputs(200)));
    layer0_outputs(1365) <= inputs(80);
    layer0_outputs(1366) <= not(inputs(246));
    layer0_outputs(1367) <= '1';
    layer0_outputs(1368) <= not(inputs(235)) or (inputs(97));
    layer0_outputs(1369) <= '0';
    layer0_outputs(1370) <= (inputs(5)) or (inputs(71));
    layer0_outputs(1371) <= not((inputs(130)) or (inputs(216)));
    layer0_outputs(1372) <= '1';
    layer0_outputs(1373) <= not((inputs(236)) or (inputs(196)));
    layer0_outputs(1374) <= (inputs(167)) and not (inputs(31));
    layer0_outputs(1375) <= not(inputs(89));
    layer0_outputs(1376) <= (inputs(240)) or (inputs(153));
    layer0_outputs(1377) <= not(inputs(184)) or (inputs(102));
    layer0_outputs(1378) <= '0';
    layer0_outputs(1379) <= inputs(11);
    layer0_outputs(1380) <= not(inputs(107)) or (inputs(234));
    layer0_outputs(1381) <= (inputs(148)) and not (inputs(242));
    layer0_outputs(1382) <= not(inputs(3));
    layer0_outputs(1383) <= inputs(20);
    layer0_outputs(1384) <= not(inputs(86));
    layer0_outputs(1385) <= not(inputs(79));
    layer0_outputs(1386) <= not(inputs(99));
    layer0_outputs(1387) <= (inputs(104)) and (inputs(49));
    layer0_outputs(1388) <= '1';
    layer0_outputs(1389) <= (inputs(82)) and not (inputs(222));
    layer0_outputs(1390) <= inputs(59);
    layer0_outputs(1391) <= not(inputs(233));
    layer0_outputs(1392) <= not((inputs(42)) and (inputs(39)));
    layer0_outputs(1393) <= (inputs(212)) and not (inputs(48));
    layer0_outputs(1394) <= not((inputs(4)) or (inputs(122)));
    layer0_outputs(1395) <= (inputs(3)) or (inputs(125));
    layer0_outputs(1396) <= (inputs(230)) xor (inputs(177));
    layer0_outputs(1397) <= inputs(136);
    layer0_outputs(1398) <= not(inputs(15)) or (inputs(154));
    layer0_outputs(1399) <= not(inputs(27)) or (inputs(231));
    layer0_outputs(1400) <= (inputs(95)) or (inputs(23));
    layer0_outputs(1401) <= (inputs(96)) and not (inputs(33));
    layer0_outputs(1402) <= not((inputs(195)) or (inputs(3)));
    layer0_outputs(1403) <= not(inputs(134));
    layer0_outputs(1404) <= inputs(211);
    layer0_outputs(1405) <= inputs(53);
    layer0_outputs(1406) <= not(inputs(11)) or (inputs(89));
    layer0_outputs(1407) <= not((inputs(253)) or (inputs(131)));
    layer0_outputs(1408) <= inputs(217);
    layer0_outputs(1409) <= (inputs(192)) or (inputs(24));
    layer0_outputs(1410) <= (inputs(87)) or (inputs(113));
    layer0_outputs(1411) <= (inputs(74)) or (inputs(88));
    layer0_outputs(1412) <= not((inputs(53)) or (inputs(114)));
    layer0_outputs(1413) <= inputs(94);
    layer0_outputs(1414) <= '0';
    layer0_outputs(1415) <= not(inputs(77));
    layer0_outputs(1416) <= not(inputs(150));
    layer0_outputs(1417) <= not(inputs(121));
    layer0_outputs(1418) <= not((inputs(95)) or (inputs(252)));
    layer0_outputs(1419) <= (inputs(99)) and not (inputs(157));
    layer0_outputs(1420) <= (inputs(189)) or (inputs(56));
    layer0_outputs(1421) <= not((inputs(195)) xor (inputs(174)));
    layer0_outputs(1422) <= not((inputs(28)) or (inputs(238)));
    layer0_outputs(1423) <= not(inputs(47));
    layer0_outputs(1424) <= not(inputs(204));
    layer0_outputs(1425) <= not(inputs(43)) or (inputs(137));
    layer0_outputs(1426) <= '0';
    layer0_outputs(1427) <= not(inputs(24));
    layer0_outputs(1428) <= not((inputs(36)) or (inputs(242)));
    layer0_outputs(1429) <= not(inputs(138));
    layer0_outputs(1430) <= not((inputs(247)) and (inputs(120)));
    layer0_outputs(1431) <= inputs(247);
    layer0_outputs(1432) <= not(inputs(141));
    layer0_outputs(1433) <= (inputs(41)) or (inputs(95));
    layer0_outputs(1434) <= not(inputs(172)) or (inputs(93));
    layer0_outputs(1435) <= not(inputs(156)) or (inputs(193));
    layer0_outputs(1436) <= inputs(143);
    layer0_outputs(1437) <= inputs(106);
    layer0_outputs(1438) <= not((inputs(187)) or (inputs(26)));
    layer0_outputs(1439) <= not(inputs(117));
    layer0_outputs(1440) <= (inputs(136)) and not (inputs(222));
    layer0_outputs(1441) <= inputs(129);
    layer0_outputs(1442) <= not(inputs(237));
    layer0_outputs(1443) <= not((inputs(107)) or (inputs(124)));
    layer0_outputs(1444) <= not(inputs(205));
    layer0_outputs(1445) <= inputs(137);
    layer0_outputs(1446) <= not(inputs(16)) or (inputs(38));
    layer0_outputs(1447) <= not((inputs(67)) and (inputs(190)));
    layer0_outputs(1448) <= '0';
    layer0_outputs(1449) <= not(inputs(178));
    layer0_outputs(1450) <= not(inputs(8)) or (inputs(151));
    layer0_outputs(1451) <= '0';
    layer0_outputs(1452) <= (inputs(2)) xor (inputs(72));
    layer0_outputs(1453) <= not(inputs(28)) or (inputs(187));
    layer0_outputs(1454) <= not(inputs(78));
    layer0_outputs(1455) <= not(inputs(133));
    layer0_outputs(1456) <= (inputs(45)) and not (inputs(134));
    layer0_outputs(1457) <= inputs(93);
    layer0_outputs(1458) <= not(inputs(62));
    layer0_outputs(1459) <= '0';
    layer0_outputs(1460) <= (inputs(7)) and (inputs(21));
    layer0_outputs(1461) <= (inputs(101)) and not (inputs(125));
    layer0_outputs(1462) <= not((inputs(157)) or (inputs(202)));
    layer0_outputs(1463) <= not(inputs(122));
    layer0_outputs(1464) <= (inputs(158)) or (inputs(63));
    layer0_outputs(1465) <= not(inputs(65));
    layer0_outputs(1466) <= inputs(230);
    layer0_outputs(1467) <= inputs(226);
    layer0_outputs(1468) <= not(inputs(180)) or (inputs(158));
    layer0_outputs(1469) <= not(inputs(150));
    layer0_outputs(1470) <= (inputs(168)) or (inputs(144));
    layer0_outputs(1471) <= (inputs(1)) or (inputs(207));
    layer0_outputs(1472) <= '1';
    layer0_outputs(1473) <= (inputs(107)) or (inputs(239));
    layer0_outputs(1474) <= not((inputs(138)) or (inputs(115)));
    layer0_outputs(1475) <= (inputs(83)) and not (inputs(78));
    layer0_outputs(1476) <= not((inputs(151)) or (inputs(227)));
    layer0_outputs(1477) <= (inputs(165)) or (inputs(4));
    layer0_outputs(1478) <= (inputs(131)) or (inputs(117));
    layer0_outputs(1479) <= not(inputs(235)) or (inputs(87));
    layer0_outputs(1480) <= (inputs(23)) and not (inputs(167));
    layer0_outputs(1481) <= not(inputs(103));
    layer0_outputs(1482) <= '1';
    layer0_outputs(1483) <= inputs(26);
    layer0_outputs(1484) <= not(inputs(95));
    layer0_outputs(1485) <= inputs(80);
    layer0_outputs(1486) <= (inputs(151)) and not (inputs(137));
    layer0_outputs(1487) <= not(inputs(205));
    layer0_outputs(1488) <= not(inputs(192));
    layer0_outputs(1489) <= (inputs(76)) and not (inputs(173));
    layer0_outputs(1490) <= '1';
    layer0_outputs(1491) <= (inputs(54)) or (inputs(125));
    layer0_outputs(1492) <= (inputs(9)) or (inputs(67));
    layer0_outputs(1493) <= (inputs(159)) xor (inputs(208));
    layer0_outputs(1494) <= not(inputs(37));
    layer0_outputs(1495) <= inputs(230);
    layer0_outputs(1496) <= (inputs(175)) or (inputs(197));
    layer0_outputs(1497) <= (inputs(242)) and not (inputs(153));
    layer0_outputs(1498) <= inputs(124);
    layer0_outputs(1499) <= (inputs(148)) or (inputs(128));
    layer0_outputs(1500) <= not((inputs(240)) or (inputs(248)));
    layer0_outputs(1501) <= '1';
    layer0_outputs(1502) <= '0';
    layer0_outputs(1503) <= '0';
    layer0_outputs(1504) <= '0';
    layer0_outputs(1505) <= not(inputs(22));
    layer0_outputs(1506) <= inputs(67);
    layer0_outputs(1507) <= not(inputs(186));
    layer0_outputs(1508) <= not(inputs(204)) or (inputs(238));
    layer0_outputs(1509) <= not((inputs(208)) or (inputs(23)));
    layer0_outputs(1510) <= '0';
    layer0_outputs(1511) <= not(inputs(255));
    layer0_outputs(1512) <= not((inputs(152)) xor (inputs(121)));
    layer0_outputs(1513) <= not(inputs(45));
    layer0_outputs(1514) <= not(inputs(29));
    layer0_outputs(1515) <= inputs(138);
    layer0_outputs(1516) <= inputs(21);
    layer0_outputs(1517) <= (inputs(132)) and not (inputs(61));
    layer0_outputs(1518) <= (inputs(203)) and not (inputs(61));
    layer0_outputs(1519) <= '1';
    layer0_outputs(1520) <= not((inputs(150)) or (inputs(162)));
    layer0_outputs(1521) <= not(inputs(101));
    layer0_outputs(1522) <= (inputs(57)) or (inputs(196));
    layer0_outputs(1523) <= not((inputs(19)) or (inputs(21)));
    layer0_outputs(1524) <= (inputs(71)) or (inputs(158));
    layer0_outputs(1525) <= not(inputs(210));
    layer0_outputs(1526) <= (inputs(220)) and not (inputs(33));
    layer0_outputs(1527) <= (inputs(157)) and (inputs(117));
    layer0_outputs(1528) <= (inputs(126)) or (inputs(217));
    layer0_outputs(1529) <= '1';
    layer0_outputs(1530) <= inputs(212);
    layer0_outputs(1531) <= (inputs(170)) or (inputs(22));
    layer0_outputs(1532) <= not((inputs(162)) or (inputs(15)));
    layer0_outputs(1533) <= not(inputs(220));
    layer0_outputs(1534) <= not(inputs(71)) or (inputs(12));
    layer0_outputs(1535) <= (inputs(77)) and not (inputs(170));
    layer0_outputs(1536) <= (inputs(132)) and not (inputs(181));
    layer0_outputs(1537) <= (inputs(245)) or (inputs(176));
    layer0_outputs(1538) <= inputs(155);
    layer0_outputs(1539) <= (inputs(120)) or (inputs(207));
    layer0_outputs(1540) <= not(inputs(11));
    layer0_outputs(1541) <= (inputs(64)) and not (inputs(174));
    layer0_outputs(1542) <= not(inputs(234));
    layer0_outputs(1543) <= not(inputs(202));
    layer0_outputs(1544) <= (inputs(192)) or (inputs(194));
    layer0_outputs(1545) <= inputs(98);
    layer0_outputs(1546) <= (inputs(82)) or (inputs(115));
    layer0_outputs(1547) <= (inputs(21)) and not (inputs(43));
    layer0_outputs(1548) <= inputs(30);
    layer0_outputs(1549) <= not(inputs(229));
    layer0_outputs(1550) <= inputs(136);
    layer0_outputs(1551) <= not(inputs(153)) or (inputs(138));
    layer0_outputs(1552) <= (inputs(180)) and not (inputs(0));
    layer0_outputs(1553) <= '0';
    layer0_outputs(1554) <= inputs(149);
    layer0_outputs(1555) <= (inputs(70)) and not (inputs(158));
    layer0_outputs(1556) <= (inputs(177)) or (inputs(123));
    layer0_outputs(1557) <= (inputs(28)) and (inputs(113));
    layer0_outputs(1558) <= not(inputs(195));
    layer0_outputs(1559) <= inputs(90);
    layer0_outputs(1560) <= not((inputs(12)) or (inputs(14)));
    layer0_outputs(1561) <= (inputs(118)) and not (inputs(164));
    layer0_outputs(1562) <= not(inputs(255)) or (inputs(109));
    layer0_outputs(1563) <= not((inputs(35)) or (inputs(108)));
    layer0_outputs(1564) <= not(inputs(23));
    layer0_outputs(1565) <= inputs(27);
    layer0_outputs(1566) <= (inputs(231)) or (inputs(248));
    layer0_outputs(1567) <= not(inputs(37));
    layer0_outputs(1568) <= inputs(230);
    layer0_outputs(1569) <= '1';
    layer0_outputs(1570) <= (inputs(207)) and not (inputs(234));
    layer0_outputs(1571) <= not(inputs(31));
    layer0_outputs(1572) <= not(inputs(233));
    layer0_outputs(1573) <= not(inputs(69)) or (inputs(1));
    layer0_outputs(1574) <= inputs(91);
    layer0_outputs(1575) <= not((inputs(227)) and (inputs(10)));
    layer0_outputs(1576) <= not(inputs(121));
    layer0_outputs(1577) <= not(inputs(222));
    layer0_outputs(1578) <= (inputs(84)) and not (inputs(93));
    layer0_outputs(1579) <= not(inputs(231));
    layer0_outputs(1580) <= not(inputs(138));
    layer0_outputs(1581) <= not(inputs(170)) or (inputs(63));
    layer0_outputs(1582) <= (inputs(171)) or (inputs(154));
    layer0_outputs(1583) <= (inputs(80)) or (inputs(211));
    layer0_outputs(1584) <= inputs(88);
    layer0_outputs(1585) <= (inputs(31)) and (inputs(106));
    layer0_outputs(1586) <= not((inputs(18)) xor (inputs(111)));
    layer0_outputs(1587) <= not((inputs(135)) or (inputs(213)));
    layer0_outputs(1588) <= (inputs(225)) xor (inputs(176));
    layer0_outputs(1589) <= not((inputs(232)) or (inputs(217)));
    layer0_outputs(1590) <= (inputs(52)) or (inputs(130));
    layer0_outputs(1591) <= inputs(89);
    layer0_outputs(1592) <= not(inputs(114));
    layer0_outputs(1593) <= not(inputs(96));
    layer0_outputs(1594) <= not(inputs(243));
    layer0_outputs(1595) <= (inputs(95)) xor (inputs(47));
    layer0_outputs(1596) <= inputs(178);
    layer0_outputs(1597) <= '1';
    layer0_outputs(1598) <= inputs(25);
    layer0_outputs(1599) <= not((inputs(170)) or (inputs(124)));
    layer0_outputs(1600) <= inputs(180);
    layer0_outputs(1601) <= not(inputs(40));
    layer0_outputs(1602) <= '1';
    layer0_outputs(1603) <= (inputs(229)) or (inputs(115));
    layer0_outputs(1604) <= (inputs(201)) xor (inputs(176));
    layer0_outputs(1605) <= (inputs(11)) and (inputs(62));
    layer0_outputs(1606) <= not(inputs(114));
    layer0_outputs(1607) <= (inputs(241)) and not (inputs(183));
    layer0_outputs(1608) <= not(inputs(223));
    layer0_outputs(1609) <= not((inputs(179)) or (inputs(40)));
    layer0_outputs(1610) <= not(inputs(115));
    layer0_outputs(1611) <= inputs(203);
    layer0_outputs(1612) <= '1';
    layer0_outputs(1613) <= not((inputs(18)) or (inputs(94)));
    layer0_outputs(1614) <= not(inputs(198)) or (inputs(97));
    layer0_outputs(1615) <= not(inputs(87));
    layer0_outputs(1616) <= not((inputs(140)) or (inputs(155)));
    layer0_outputs(1617) <= inputs(168);
    layer0_outputs(1618) <= not(inputs(116));
    layer0_outputs(1619) <= inputs(29);
    layer0_outputs(1620) <= not(inputs(139)) or (inputs(193));
    layer0_outputs(1621) <= not(inputs(134)) or (inputs(200));
    layer0_outputs(1622) <= inputs(114);
    layer0_outputs(1623) <= not((inputs(198)) or (inputs(228)));
    layer0_outputs(1624) <= inputs(219);
    layer0_outputs(1625) <= not((inputs(115)) or (inputs(98)));
    layer0_outputs(1626) <= (inputs(186)) or (inputs(248));
    layer0_outputs(1627) <= not(inputs(200));
    layer0_outputs(1628) <= not((inputs(23)) or (inputs(4)));
    layer0_outputs(1629) <= '0';
    layer0_outputs(1630) <= (inputs(67)) and not (inputs(50));
    layer0_outputs(1631) <= not((inputs(152)) or (inputs(186)));
    layer0_outputs(1632) <= '1';
    layer0_outputs(1633) <= (inputs(151)) and not (inputs(108));
    layer0_outputs(1634) <= (inputs(15)) and not (inputs(61));
    layer0_outputs(1635) <= not(inputs(188));
    layer0_outputs(1636) <= not(inputs(240)) or (inputs(92));
    layer0_outputs(1637) <= not(inputs(149));
    layer0_outputs(1638) <= not((inputs(179)) or (inputs(84)));
    layer0_outputs(1639) <= not((inputs(225)) or (inputs(120)));
    layer0_outputs(1640) <= inputs(199);
    layer0_outputs(1641) <= not(inputs(218));
    layer0_outputs(1642) <= (inputs(90)) and (inputs(41));
    layer0_outputs(1643) <= not(inputs(215)) or (inputs(101));
    layer0_outputs(1644) <= inputs(170);
    layer0_outputs(1645) <= not(inputs(70)) or (inputs(22));
    layer0_outputs(1646) <= not(inputs(229)) or (inputs(76));
    layer0_outputs(1647) <= (inputs(179)) or (inputs(199));
    layer0_outputs(1648) <= inputs(173);
    layer0_outputs(1649) <= (inputs(177)) xor (inputs(2));
    layer0_outputs(1650) <= (inputs(182)) and not (inputs(236));
    layer0_outputs(1651) <= '1';
    layer0_outputs(1652) <= inputs(52);
    layer0_outputs(1653) <= (inputs(110)) or (inputs(125));
    layer0_outputs(1654) <= (inputs(74)) and not (inputs(246));
    layer0_outputs(1655) <= not((inputs(189)) or (inputs(122)));
    layer0_outputs(1656) <= not(inputs(130)) or (inputs(17));
    layer0_outputs(1657) <= (inputs(126)) and not (inputs(90));
    layer0_outputs(1658) <= not(inputs(50));
    layer0_outputs(1659) <= (inputs(213)) and not (inputs(47));
    layer0_outputs(1660) <= not(inputs(218));
    layer0_outputs(1661) <= '0';
    layer0_outputs(1662) <= '1';
    layer0_outputs(1663) <= (inputs(58)) and not (inputs(149));
    layer0_outputs(1664) <= inputs(145);
    layer0_outputs(1665) <= not(inputs(75)) or (inputs(102));
    layer0_outputs(1666) <= (inputs(146)) or (inputs(156));
    layer0_outputs(1667) <= not((inputs(251)) and (inputs(184)));
    layer0_outputs(1668) <= (inputs(31)) and not (inputs(57));
    layer0_outputs(1669) <= not(inputs(106));
    layer0_outputs(1670) <= (inputs(18)) and not (inputs(106));
    layer0_outputs(1671) <= (inputs(54)) xor (inputs(201));
    layer0_outputs(1672) <= not((inputs(86)) xor (inputs(45)));
    layer0_outputs(1673) <= not(inputs(160)) or (inputs(253));
    layer0_outputs(1674) <= not(inputs(230)) or (inputs(121));
    layer0_outputs(1675) <= not(inputs(8)) or (inputs(3));
    layer0_outputs(1676) <= (inputs(129)) or (inputs(149));
    layer0_outputs(1677) <= not(inputs(129));
    layer0_outputs(1678) <= (inputs(163)) or (inputs(180));
    layer0_outputs(1679) <= not(inputs(243)) or (inputs(140));
    layer0_outputs(1680) <= inputs(136);
    layer0_outputs(1681) <= not(inputs(148));
    layer0_outputs(1682) <= not(inputs(255));
    layer0_outputs(1683) <= inputs(228);
    layer0_outputs(1684) <= not(inputs(227));
    layer0_outputs(1685) <= '0';
    layer0_outputs(1686) <= not((inputs(210)) or (inputs(132)));
    layer0_outputs(1687) <= not(inputs(165));
    layer0_outputs(1688) <= not((inputs(129)) or (inputs(100)));
    layer0_outputs(1689) <= (inputs(105)) and not (inputs(229));
    layer0_outputs(1690) <= not(inputs(73)) or (inputs(67));
    layer0_outputs(1691) <= (inputs(0)) and not (inputs(165));
    layer0_outputs(1692) <= not((inputs(85)) or (inputs(187)));
    layer0_outputs(1693) <= not(inputs(135));
    layer0_outputs(1694) <= not(inputs(133));
    layer0_outputs(1695) <= not((inputs(132)) or (inputs(68)));
    layer0_outputs(1696) <= '1';
    layer0_outputs(1697) <= not(inputs(116));
    layer0_outputs(1698) <= not(inputs(230));
    layer0_outputs(1699) <= (inputs(104)) and not (inputs(140));
    layer0_outputs(1700) <= '0';
    layer0_outputs(1701) <= inputs(186);
    layer0_outputs(1702) <= inputs(84);
    layer0_outputs(1703) <= (inputs(186)) and (inputs(48));
    layer0_outputs(1704) <= inputs(90);
    layer0_outputs(1705) <= inputs(207);
    layer0_outputs(1706) <= (inputs(28)) and not (inputs(160));
    layer0_outputs(1707) <= not(inputs(128));
    layer0_outputs(1708) <= '0';
    layer0_outputs(1709) <= not(inputs(253));
    layer0_outputs(1710) <= inputs(253);
    layer0_outputs(1711) <= inputs(163);
    layer0_outputs(1712) <= (inputs(227)) or (inputs(225));
    layer0_outputs(1713) <= inputs(123);
    layer0_outputs(1714) <= not((inputs(249)) and (inputs(206)));
    layer0_outputs(1715) <= not((inputs(166)) or (inputs(4)));
    layer0_outputs(1716) <= (inputs(253)) or (inputs(92));
    layer0_outputs(1717) <= not(inputs(47));
    layer0_outputs(1718) <= inputs(180);
    layer0_outputs(1719) <= '1';
    layer0_outputs(1720) <= (inputs(250)) and not (inputs(234));
    layer0_outputs(1721) <= not(inputs(67)) or (inputs(152));
    layer0_outputs(1722) <= (inputs(104)) and not (inputs(145));
    layer0_outputs(1723) <= not((inputs(92)) or (inputs(64)));
    layer0_outputs(1724) <= inputs(43);
    layer0_outputs(1725) <= not(inputs(173));
    layer0_outputs(1726) <= (inputs(23)) or (inputs(19));
    layer0_outputs(1727) <= (inputs(121)) or (inputs(79));
    layer0_outputs(1728) <= (inputs(171)) and not (inputs(52));
    layer0_outputs(1729) <= not(inputs(104)) or (inputs(160));
    layer0_outputs(1730) <= not(inputs(18)) or (inputs(81));
    layer0_outputs(1731) <= '0';
    layer0_outputs(1732) <= not(inputs(137));
    layer0_outputs(1733) <= '0';
    layer0_outputs(1734) <= not(inputs(56)) or (inputs(181));
    layer0_outputs(1735) <= not(inputs(191));
    layer0_outputs(1736) <= (inputs(236)) and not (inputs(128));
    layer0_outputs(1737) <= inputs(116);
    layer0_outputs(1738) <= (inputs(58)) or (inputs(78));
    layer0_outputs(1739) <= not(inputs(192));
    layer0_outputs(1740) <= (inputs(5)) xor (inputs(47));
    layer0_outputs(1741) <= (inputs(117)) or (inputs(166));
    layer0_outputs(1742) <= not((inputs(28)) or (inputs(61)));
    layer0_outputs(1743) <= not(inputs(24));
    layer0_outputs(1744) <= (inputs(169)) and not (inputs(120));
    layer0_outputs(1745) <= (inputs(180)) and not (inputs(249));
    layer0_outputs(1746) <= not(inputs(99));
    layer0_outputs(1747) <= not(inputs(25)) or (inputs(202));
    layer0_outputs(1748) <= (inputs(146)) or (inputs(86));
    layer0_outputs(1749) <= (inputs(235)) and not (inputs(239));
    layer0_outputs(1750) <= (inputs(90)) and not (inputs(126));
    layer0_outputs(1751) <= (inputs(140)) or (inputs(110));
    layer0_outputs(1752) <= not(inputs(68));
    layer0_outputs(1753) <= (inputs(41)) or (inputs(242));
    layer0_outputs(1754) <= not(inputs(107));
    layer0_outputs(1755) <= inputs(221);
    layer0_outputs(1756) <= inputs(212);
    layer0_outputs(1757) <= not(inputs(22)) or (inputs(132));
    layer0_outputs(1758) <= (inputs(9)) or (inputs(188));
    layer0_outputs(1759) <= not((inputs(232)) and (inputs(170)));
    layer0_outputs(1760) <= not(inputs(210));
    layer0_outputs(1761) <= inputs(120);
    layer0_outputs(1762) <= not(inputs(252));
    layer0_outputs(1763) <= (inputs(161)) or (inputs(159));
    layer0_outputs(1764) <= (inputs(65)) and not (inputs(239));
    layer0_outputs(1765) <= not((inputs(170)) or (inputs(249)));
    layer0_outputs(1766) <= (inputs(59)) or (inputs(136));
    layer0_outputs(1767) <= (inputs(34)) and not (inputs(118));
    layer0_outputs(1768) <= not(inputs(49)) or (inputs(59));
    layer0_outputs(1769) <= (inputs(120)) and not (inputs(216));
    layer0_outputs(1770) <= not(inputs(57));
    layer0_outputs(1771) <= (inputs(32)) or (inputs(11));
    layer0_outputs(1772) <= not(inputs(227));
    layer0_outputs(1773) <= (inputs(27)) or (inputs(103));
    layer0_outputs(1774) <= not((inputs(29)) and (inputs(255)));
    layer0_outputs(1775) <= (inputs(169)) or (inputs(63));
    layer0_outputs(1776) <= (inputs(94)) and (inputs(143));
    layer0_outputs(1777) <= (inputs(80)) xor (inputs(19));
    layer0_outputs(1778) <= (inputs(234)) or (inputs(230));
    layer0_outputs(1779) <= '1';
    layer0_outputs(1780) <= inputs(25);
    layer0_outputs(1781) <= not((inputs(178)) or (inputs(182)));
    layer0_outputs(1782) <= (inputs(173)) and not (inputs(43));
    layer0_outputs(1783) <= not(inputs(224)) or (inputs(224));
    layer0_outputs(1784) <= (inputs(6)) and not (inputs(236));
    layer0_outputs(1785) <= not(inputs(128));
    layer0_outputs(1786) <= not((inputs(109)) or (inputs(227)));
    layer0_outputs(1787) <= inputs(204);
    layer0_outputs(1788) <= not(inputs(109));
    layer0_outputs(1789) <= not(inputs(8));
    layer0_outputs(1790) <= '1';
    layer0_outputs(1791) <= (inputs(98)) or (inputs(131));
    layer0_outputs(1792) <= (inputs(103)) and not (inputs(253));
    layer0_outputs(1793) <= (inputs(96)) or (inputs(139));
    layer0_outputs(1794) <= not((inputs(203)) or (inputs(114)));
    layer0_outputs(1795) <= '1';
    layer0_outputs(1796) <= inputs(33);
    layer0_outputs(1797) <= not((inputs(62)) or (inputs(164)));
    layer0_outputs(1798) <= not(inputs(157));
    layer0_outputs(1799) <= (inputs(37)) and not (inputs(200));
    layer0_outputs(1800) <= not(inputs(218));
    layer0_outputs(1801) <= inputs(73);
    layer0_outputs(1802) <= inputs(84);
    layer0_outputs(1803) <= not(inputs(122));
    layer0_outputs(1804) <= (inputs(140)) and not (inputs(180));
    layer0_outputs(1805) <= '0';
    layer0_outputs(1806) <= (inputs(164)) or (inputs(246));
    layer0_outputs(1807) <= not((inputs(76)) or (inputs(161)));
    layer0_outputs(1808) <= not((inputs(172)) xor (inputs(252)));
    layer0_outputs(1809) <= not((inputs(19)) xor (inputs(64)));
    layer0_outputs(1810) <= not(inputs(90));
    layer0_outputs(1811) <= not((inputs(33)) or (inputs(120)));
    layer0_outputs(1812) <= not((inputs(61)) or (inputs(174)));
    layer0_outputs(1813) <= (inputs(186)) or (inputs(141));
    layer0_outputs(1814) <= not(inputs(70));
    layer0_outputs(1815) <= not(inputs(215));
    layer0_outputs(1816) <= not((inputs(10)) or (inputs(39)));
    layer0_outputs(1817) <= not((inputs(189)) or (inputs(73)));
    layer0_outputs(1818) <= inputs(51);
    layer0_outputs(1819) <= inputs(181);
    layer0_outputs(1820) <= (inputs(74)) and not (inputs(186));
    layer0_outputs(1821) <= inputs(91);
    layer0_outputs(1822) <= inputs(77);
    layer0_outputs(1823) <= not((inputs(190)) or (inputs(218)));
    layer0_outputs(1824) <= not(inputs(243)) or (inputs(103));
    layer0_outputs(1825) <= (inputs(172)) or (inputs(223));
    layer0_outputs(1826) <= (inputs(123)) or (inputs(236));
    layer0_outputs(1827) <= not(inputs(46)) or (inputs(165));
    layer0_outputs(1828) <= (inputs(53)) or (inputs(16));
    layer0_outputs(1829) <= not(inputs(27)) or (inputs(228));
    layer0_outputs(1830) <= inputs(31);
    layer0_outputs(1831) <= not((inputs(177)) or (inputs(10)));
    layer0_outputs(1832) <= not(inputs(222));
    layer0_outputs(1833) <= not(inputs(239)) or (inputs(14));
    layer0_outputs(1834) <= (inputs(222)) and (inputs(243));
    layer0_outputs(1835) <= not((inputs(156)) xor (inputs(97)));
    layer0_outputs(1836) <= (inputs(19)) and (inputs(49));
    layer0_outputs(1837) <= not((inputs(100)) or (inputs(15)));
    layer0_outputs(1838) <= not(inputs(103)) or (inputs(145));
    layer0_outputs(1839) <= (inputs(176)) and (inputs(48));
    layer0_outputs(1840) <= not((inputs(57)) xor (inputs(0)));
    layer0_outputs(1841) <= not(inputs(209));
    layer0_outputs(1842) <= inputs(34);
    layer0_outputs(1843) <= inputs(25);
    layer0_outputs(1844) <= inputs(194);
    layer0_outputs(1845) <= '1';
    layer0_outputs(1846) <= not(inputs(199));
    layer0_outputs(1847) <= (inputs(26)) or (inputs(176));
    layer0_outputs(1848) <= not(inputs(180));
    layer0_outputs(1849) <= inputs(105);
    layer0_outputs(1850) <= '0';
    layer0_outputs(1851) <= '1';
    layer0_outputs(1852) <= not(inputs(57));
    layer0_outputs(1853) <= inputs(63);
    layer0_outputs(1854) <= (inputs(114)) and (inputs(178));
    layer0_outputs(1855) <= (inputs(126)) and not (inputs(14));
    layer0_outputs(1856) <= inputs(19);
    layer0_outputs(1857) <= (inputs(194)) and not (inputs(233));
    layer0_outputs(1858) <= not((inputs(206)) or (inputs(237)));
    layer0_outputs(1859) <= inputs(125);
    layer0_outputs(1860) <= inputs(76);
    layer0_outputs(1861) <= (inputs(118)) and (inputs(24));
    layer0_outputs(1862) <= '1';
    layer0_outputs(1863) <= not((inputs(176)) or (inputs(214)));
    layer0_outputs(1864) <= not((inputs(38)) or (inputs(162)));
    layer0_outputs(1865) <= (inputs(76)) or (inputs(6));
    layer0_outputs(1866) <= (inputs(130)) or (inputs(118));
    layer0_outputs(1867) <= not((inputs(87)) or (inputs(38)));
    layer0_outputs(1868) <= not(inputs(232)) or (inputs(242));
    layer0_outputs(1869) <= not((inputs(26)) or (inputs(67)));
    layer0_outputs(1870) <= '1';
    layer0_outputs(1871) <= (inputs(213)) and (inputs(6));
    layer0_outputs(1872) <= not(inputs(138));
    layer0_outputs(1873) <= inputs(93);
    layer0_outputs(1874) <= (inputs(58)) xor (inputs(1));
    layer0_outputs(1875) <= not(inputs(159));
    layer0_outputs(1876) <= (inputs(210)) and not (inputs(75));
    layer0_outputs(1877) <= not((inputs(144)) xor (inputs(181)));
    layer0_outputs(1878) <= not(inputs(148)) or (inputs(139));
    layer0_outputs(1879) <= inputs(99);
    layer0_outputs(1880) <= (inputs(34)) or (inputs(64));
    layer0_outputs(1881) <= (inputs(201)) and not (inputs(216));
    layer0_outputs(1882) <= not(inputs(85)) or (inputs(189));
    layer0_outputs(1883) <= not(inputs(237)) or (inputs(2));
    layer0_outputs(1884) <= inputs(98);
    layer0_outputs(1885) <= inputs(157);
    layer0_outputs(1886) <= not(inputs(40));
    layer0_outputs(1887) <= not(inputs(145)) or (inputs(31));
    layer0_outputs(1888) <= not(inputs(107));
    layer0_outputs(1889) <= not(inputs(172)) or (inputs(89));
    layer0_outputs(1890) <= not((inputs(191)) or (inputs(197)));
    layer0_outputs(1891) <= not((inputs(253)) or (inputs(114)));
    layer0_outputs(1892) <= (inputs(179)) or (inputs(191));
    layer0_outputs(1893) <= not((inputs(195)) or (inputs(202)));
    layer0_outputs(1894) <= not(inputs(155)) or (inputs(241));
    layer0_outputs(1895) <= not((inputs(12)) xor (inputs(73)));
    layer0_outputs(1896) <= not((inputs(38)) and (inputs(9)));
    layer0_outputs(1897) <= not((inputs(72)) or (inputs(126)));
    layer0_outputs(1898) <= not(inputs(226));
    layer0_outputs(1899) <= inputs(138);
    layer0_outputs(1900) <= not(inputs(84));
    layer0_outputs(1901) <= (inputs(226)) and not (inputs(95));
    layer0_outputs(1902) <= not((inputs(252)) and (inputs(45)));
    layer0_outputs(1903) <= (inputs(142)) or (inputs(72));
    layer0_outputs(1904) <= not(inputs(90));
    layer0_outputs(1905) <= not((inputs(198)) or (inputs(17)));
    layer0_outputs(1906) <= not(inputs(105)) or (inputs(17));
    layer0_outputs(1907) <= inputs(178);
    layer0_outputs(1908) <= inputs(100);
    layer0_outputs(1909) <= not(inputs(93)) or (inputs(107));
    layer0_outputs(1910) <= not((inputs(25)) and (inputs(62)));
    layer0_outputs(1911) <= not((inputs(177)) or (inputs(211)));
    layer0_outputs(1912) <= not(inputs(56));
    layer0_outputs(1913) <= not(inputs(94));
    layer0_outputs(1914) <= inputs(153);
    layer0_outputs(1915) <= inputs(35);
    layer0_outputs(1916) <= not(inputs(219));
    layer0_outputs(1917) <= not(inputs(75));
    layer0_outputs(1918) <= inputs(60);
    layer0_outputs(1919) <= not((inputs(178)) or (inputs(234)));
    layer0_outputs(1920) <= not(inputs(192)) or (inputs(14));
    layer0_outputs(1921) <= not(inputs(53)) or (inputs(139));
    layer0_outputs(1922) <= not(inputs(113));
    layer0_outputs(1923) <= (inputs(224)) and not (inputs(146));
    layer0_outputs(1924) <= inputs(102);
    layer0_outputs(1925) <= inputs(97);
    layer0_outputs(1926) <= (inputs(8)) or (inputs(33));
    layer0_outputs(1927) <= not((inputs(222)) or (inputs(106)));
    layer0_outputs(1928) <= '0';
    layer0_outputs(1929) <= not(inputs(40)) or (inputs(153));
    layer0_outputs(1930) <= (inputs(167)) and not (inputs(128));
    layer0_outputs(1931) <= (inputs(61)) or (inputs(124));
    layer0_outputs(1932) <= not(inputs(106));
    layer0_outputs(1933) <= (inputs(70)) and (inputs(229));
    layer0_outputs(1934) <= not((inputs(38)) or (inputs(22)));
    layer0_outputs(1935) <= inputs(116);
    layer0_outputs(1936) <= not(inputs(115));
    layer0_outputs(1937) <= (inputs(54)) and not (inputs(136));
    layer0_outputs(1938) <= '0';
    layer0_outputs(1939) <= (inputs(153)) or (inputs(98));
    layer0_outputs(1940) <= (inputs(62)) and not (inputs(134));
    layer0_outputs(1941) <= not(inputs(69));
    layer0_outputs(1942) <= inputs(203);
    layer0_outputs(1943) <= not(inputs(36)) or (inputs(142));
    layer0_outputs(1944) <= (inputs(0)) and not (inputs(96));
    layer0_outputs(1945) <= inputs(197);
    layer0_outputs(1946) <= (inputs(36)) or (inputs(178));
    layer0_outputs(1947) <= '0';
    layer0_outputs(1948) <= not((inputs(228)) or (inputs(80)));
    layer0_outputs(1949) <= not(inputs(135)) or (inputs(27));
    layer0_outputs(1950) <= inputs(145);
    layer0_outputs(1951) <= not(inputs(49)) or (inputs(152));
    layer0_outputs(1952) <= not(inputs(163));
    layer0_outputs(1953) <= (inputs(110)) or (inputs(56));
    layer0_outputs(1954) <= inputs(92);
    layer0_outputs(1955) <= not((inputs(149)) or (inputs(238)));
    layer0_outputs(1956) <= (inputs(207)) or (inputs(104));
    layer0_outputs(1957) <= (inputs(94)) or (inputs(143));
    layer0_outputs(1958) <= '0';
    layer0_outputs(1959) <= inputs(5);
    layer0_outputs(1960) <= not((inputs(252)) or (inputs(60)));
    layer0_outputs(1961) <= '0';
    layer0_outputs(1962) <= not((inputs(168)) or (inputs(69)));
    layer0_outputs(1963) <= not((inputs(198)) or (inputs(5)));
    layer0_outputs(1964) <= inputs(114);
    layer0_outputs(1965) <= '0';
    layer0_outputs(1966) <= (inputs(169)) xor (inputs(0));
    layer0_outputs(1967) <= (inputs(64)) and not (inputs(206));
    layer0_outputs(1968) <= inputs(130);
    layer0_outputs(1969) <= (inputs(142)) or (inputs(76));
    layer0_outputs(1970) <= (inputs(215)) and not (inputs(195));
    layer0_outputs(1971) <= not((inputs(174)) or (inputs(208)));
    layer0_outputs(1972) <= inputs(199);
    layer0_outputs(1973) <= inputs(213);
    layer0_outputs(1974) <= not(inputs(68));
    layer0_outputs(1975) <= not(inputs(245));
    layer0_outputs(1976) <= inputs(90);
    layer0_outputs(1977) <= not(inputs(149));
    layer0_outputs(1978) <= '0';
    layer0_outputs(1979) <= inputs(2);
    layer0_outputs(1980) <= inputs(99);
    layer0_outputs(1981) <= inputs(196);
    layer0_outputs(1982) <= not(inputs(31));
    layer0_outputs(1983) <= not((inputs(223)) or (inputs(211)));
    layer0_outputs(1984) <= (inputs(126)) or (inputs(52));
    layer0_outputs(1985) <= inputs(150);
    layer0_outputs(1986) <= inputs(246);
    layer0_outputs(1987) <= inputs(92);
    layer0_outputs(1988) <= not(inputs(128));
    layer0_outputs(1989) <= not((inputs(35)) or (inputs(49)));
    layer0_outputs(1990) <= (inputs(17)) and not (inputs(13));
    layer0_outputs(1991) <= inputs(97);
    layer0_outputs(1992) <= inputs(246);
    layer0_outputs(1993) <= '1';
    layer0_outputs(1994) <= not((inputs(152)) or (inputs(152)));
    layer0_outputs(1995) <= not(inputs(72));
    layer0_outputs(1996) <= (inputs(243)) and not (inputs(97));
    layer0_outputs(1997) <= inputs(60);
    layer0_outputs(1998) <= (inputs(43)) and (inputs(221));
    layer0_outputs(1999) <= (inputs(123)) or (inputs(16));
    layer0_outputs(2000) <= '0';
    layer0_outputs(2001) <= (inputs(161)) or (inputs(197));
    layer0_outputs(2002) <= inputs(165);
    layer0_outputs(2003) <= (inputs(124)) and not (inputs(119));
    layer0_outputs(2004) <= not(inputs(248)) or (inputs(11));
    layer0_outputs(2005) <= (inputs(33)) and (inputs(133));
    layer0_outputs(2006) <= inputs(121);
    layer0_outputs(2007) <= (inputs(251)) and (inputs(224));
    layer0_outputs(2008) <= '1';
    layer0_outputs(2009) <= not((inputs(104)) and (inputs(144)));
    layer0_outputs(2010) <= '1';
    layer0_outputs(2011) <= not(inputs(36)) or (inputs(125));
    layer0_outputs(2012) <= '1';
    layer0_outputs(2013) <= '0';
    layer0_outputs(2014) <= not((inputs(218)) or (inputs(201)));
    layer0_outputs(2015) <= not(inputs(152));
    layer0_outputs(2016) <= inputs(153);
    layer0_outputs(2017) <= not(inputs(22));
    layer0_outputs(2018) <= not(inputs(212));
    layer0_outputs(2019) <= (inputs(9)) and (inputs(48));
    layer0_outputs(2020) <= (inputs(43)) and not (inputs(220));
    layer0_outputs(2021) <= inputs(11);
    layer0_outputs(2022) <= not((inputs(142)) or (inputs(63)));
    layer0_outputs(2023) <= not((inputs(234)) or (inputs(72)));
    layer0_outputs(2024) <= not((inputs(246)) or (inputs(190)));
    layer0_outputs(2025) <= not(inputs(133));
    layer0_outputs(2026) <= not(inputs(99));
    layer0_outputs(2027) <= inputs(134);
    layer0_outputs(2028) <= not(inputs(236)) or (inputs(121));
    layer0_outputs(2029) <= not(inputs(172));
    layer0_outputs(2030) <= (inputs(193)) and not (inputs(232));
    layer0_outputs(2031) <= inputs(156);
    layer0_outputs(2032) <= inputs(99);
    layer0_outputs(2033) <= not((inputs(38)) or (inputs(2)));
    layer0_outputs(2034) <= (inputs(208)) and not (inputs(81));
    layer0_outputs(2035) <= (inputs(68)) and not (inputs(0));
    layer0_outputs(2036) <= (inputs(71)) and not (inputs(157));
    layer0_outputs(2037) <= not(inputs(127)) or (inputs(16));
    layer0_outputs(2038) <= inputs(141);
    layer0_outputs(2039) <= not(inputs(210));
    layer0_outputs(2040) <= (inputs(90)) and not (inputs(58));
    layer0_outputs(2041) <= not(inputs(173));
    layer0_outputs(2042) <= inputs(134);
    layer0_outputs(2043) <= not(inputs(121));
    layer0_outputs(2044) <= not((inputs(253)) or (inputs(155)));
    layer0_outputs(2045) <= not(inputs(233)) or (inputs(9));
    layer0_outputs(2046) <= not(inputs(89)) or (inputs(188));
    layer0_outputs(2047) <= not(inputs(216)) or (inputs(0));
    layer0_outputs(2048) <= not((inputs(161)) xor (inputs(52)));
    layer0_outputs(2049) <= inputs(180);
    layer0_outputs(2050) <= '1';
    layer0_outputs(2051) <= not(inputs(34)) or (inputs(17));
    layer0_outputs(2052) <= (inputs(46)) and not (inputs(64));
    layer0_outputs(2053) <= inputs(52);
    layer0_outputs(2054) <= (inputs(91)) or (inputs(88));
    layer0_outputs(2055) <= not(inputs(102)) or (inputs(156));
    layer0_outputs(2056) <= '1';
    layer0_outputs(2057) <= (inputs(251)) or (inputs(176));
    layer0_outputs(2058) <= (inputs(216)) and not (inputs(155));
    layer0_outputs(2059) <= (inputs(188)) and (inputs(249));
    layer0_outputs(2060) <= inputs(99);
    layer0_outputs(2061) <= inputs(173);
    layer0_outputs(2062) <= not(inputs(195));
    layer0_outputs(2063) <= (inputs(215)) or (inputs(233));
    layer0_outputs(2064) <= not((inputs(95)) or (inputs(229)));
    layer0_outputs(2065) <= (inputs(182)) and not (inputs(108));
    layer0_outputs(2066) <= not((inputs(226)) or (inputs(176)));
    layer0_outputs(2067) <= (inputs(121)) and not (inputs(209));
    layer0_outputs(2068) <= inputs(131);
    layer0_outputs(2069) <= (inputs(54)) or (inputs(18));
    layer0_outputs(2070) <= not(inputs(85)) or (inputs(2));
    layer0_outputs(2071) <= not(inputs(136)) or (inputs(1));
    layer0_outputs(2072) <= not(inputs(118)) or (inputs(186));
    layer0_outputs(2073) <= inputs(127);
    layer0_outputs(2074) <= '0';
    layer0_outputs(2075) <= (inputs(227)) xor (inputs(220));
    layer0_outputs(2076) <= '1';
    layer0_outputs(2077) <= (inputs(144)) or (inputs(239));
    layer0_outputs(2078) <= not((inputs(237)) or (inputs(222)));
    layer0_outputs(2079) <= inputs(201);
    layer0_outputs(2080) <= (inputs(139)) or (inputs(66));
    layer0_outputs(2081) <= not((inputs(112)) xor (inputs(55)));
    layer0_outputs(2082) <= not(inputs(230)) or (inputs(237));
    layer0_outputs(2083) <= inputs(157);
    layer0_outputs(2084) <= (inputs(21)) xor (inputs(78));
    layer0_outputs(2085) <= not(inputs(43)) or (inputs(88));
    layer0_outputs(2086) <= (inputs(3)) or (inputs(177));
    layer0_outputs(2087) <= not(inputs(156));
    layer0_outputs(2088) <= (inputs(26)) or (inputs(77));
    layer0_outputs(2089) <= not((inputs(125)) or (inputs(191)));
    layer0_outputs(2090) <= not(inputs(159));
    layer0_outputs(2091) <= not((inputs(41)) or (inputs(110)));
    layer0_outputs(2092) <= not((inputs(54)) or (inputs(144)));
    layer0_outputs(2093) <= not(inputs(108));
    layer0_outputs(2094) <= not(inputs(182));
    layer0_outputs(2095) <= (inputs(131)) or (inputs(218));
    layer0_outputs(2096) <= (inputs(146)) or (inputs(20));
    layer0_outputs(2097) <= not(inputs(159));
    layer0_outputs(2098) <= (inputs(221)) or (inputs(99));
    layer0_outputs(2099) <= (inputs(131)) and not (inputs(7));
    layer0_outputs(2100) <= not((inputs(170)) or (inputs(47)));
    layer0_outputs(2101) <= not(inputs(124)) or (inputs(83));
    layer0_outputs(2102) <= (inputs(114)) or (inputs(96));
    layer0_outputs(2103) <= not(inputs(189));
    layer0_outputs(2104) <= (inputs(177)) or (inputs(189));
    layer0_outputs(2105) <= inputs(3);
    layer0_outputs(2106) <= (inputs(208)) or (inputs(25));
    layer0_outputs(2107) <= inputs(162);
    layer0_outputs(2108) <= not(inputs(170));
    layer0_outputs(2109) <= not(inputs(36)) or (inputs(128));
    layer0_outputs(2110) <= not(inputs(190));
    layer0_outputs(2111) <= (inputs(109)) and not (inputs(34));
    layer0_outputs(2112) <= inputs(169);
    layer0_outputs(2113) <= not((inputs(50)) and (inputs(63)));
    layer0_outputs(2114) <= inputs(196);
    layer0_outputs(2115) <= '0';
    layer0_outputs(2116) <= not(inputs(202));
    layer0_outputs(2117) <= not(inputs(173));
    layer0_outputs(2118) <= not((inputs(34)) or (inputs(3)));
    layer0_outputs(2119) <= (inputs(108)) xor (inputs(51));
    layer0_outputs(2120) <= not(inputs(237));
    layer0_outputs(2121) <= (inputs(103)) or (inputs(208));
    layer0_outputs(2122) <= not((inputs(221)) or (inputs(235)));
    layer0_outputs(2123) <= not(inputs(16));
    layer0_outputs(2124) <= (inputs(230)) and not (inputs(62));
    layer0_outputs(2125) <= (inputs(68)) or (inputs(85));
    layer0_outputs(2126) <= inputs(10);
    layer0_outputs(2127) <= not(inputs(22));
    layer0_outputs(2128) <= not(inputs(39)) or (inputs(253));
    layer0_outputs(2129) <= (inputs(67)) or (inputs(35));
    layer0_outputs(2130) <= inputs(40);
    layer0_outputs(2131) <= not((inputs(25)) or (inputs(49)));
    layer0_outputs(2132) <= not(inputs(219));
    layer0_outputs(2133) <= '1';
    layer0_outputs(2134) <= (inputs(202)) or (inputs(16));
    layer0_outputs(2135) <= inputs(13);
    layer0_outputs(2136) <= (inputs(19)) or (inputs(222));
    layer0_outputs(2137) <= (inputs(79)) or (inputs(206));
    layer0_outputs(2138) <= not(inputs(162));
    layer0_outputs(2139) <= not((inputs(106)) or (inputs(73)));
    layer0_outputs(2140) <= (inputs(254)) or (inputs(225));
    layer0_outputs(2141) <= not(inputs(133)) or (inputs(25));
    layer0_outputs(2142) <= not(inputs(146));
    layer0_outputs(2143) <= inputs(182);
    layer0_outputs(2144) <= inputs(75);
    layer0_outputs(2145) <= not(inputs(45)) or (inputs(244));
    layer0_outputs(2146) <= not(inputs(97));
    layer0_outputs(2147) <= inputs(136);
    layer0_outputs(2148) <= not((inputs(107)) or (inputs(196)));
    layer0_outputs(2149) <= inputs(231);
    layer0_outputs(2150) <= not((inputs(49)) or (inputs(168)));
    layer0_outputs(2151) <= inputs(24);
    layer0_outputs(2152) <= (inputs(253)) or (inputs(184));
    layer0_outputs(2153) <= not(inputs(82));
    layer0_outputs(2154) <= not((inputs(133)) and (inputs(73)));
    layer0_outputs(2155) <= not((inputs(108)) or (inputs(126)));
    layer0_outputs(2156) <= not((inputs(51)) or (inputs(198)));
    layer0_outputs(2157) <= not(inputs(138));
    layer0_outputs(2158) <= not((inputs(189)) xor (inputs(177)));
    layer0_outputs(2159) <= '0';
    layer0_outputs(2160) <= (inputs(115)) or (inputs(164));
    layer0_outputs(2161) <= (inputs(87)) and not (inputs(143));
    layer0_outputs(2162) <= not((inputs(236)) or (inputs(199)));
    layer0_outputs(2163) <= not((inputs(236)) or (inputs(141)));
    layer0_outputs(2164) <= not(inputs(104)) or (inputs(4));
    layer0_outputs(2165) <= (inputs(237)) xor (inputs(157));
    layer0_outputs(2166) <= not((inputs(55)) and (inputs(100)));
    layer0_outputs(2167) <= not(inputs(100));
    layer0_outputs(2168) <= not((inputs(176)) or (inputs(215)));
    layer0_outputs(2169) <= not((inputs(55)) or (inputs(250)));
    layer0_outputs(2170) <= '1';
    layer0_outputs(2171) <= not(inputs(233)) or (inputs(111));
    layer0_outputs(2172) <= (inputs(150)) and not (inputs(209));
    layer0_outputs(2173) <= (inputs(84)) and not (inputs(159));
    layer0_outputs(2174) <= not(inputs(208));
    layer0_outputs(2175) <= not(inputs(44));
    layer0_outputs(2176) <= inputs(183);
    layer0_outputs(2177) <= inputs(82);
    layer0_outputs(2178) <= (inputs(188)) and not (inputs(49));
    layer0_outputs(2179) <= not(inputs(20)) or (inputs(172));
    layer0_outputs(2180) <= not((inputs(137)) or (inputs(254)));
    layer0_outputs(2181) <= not(inputs(187));
    layer0_outputs(2182) <= not(inputs(122));
    layer0_outputs(2183) <= inputs(102);
    layer0_outputs(2184) <= inputs(214);
    layer0_outputs(2185) <= not(inputs(14)) or (inputs(200));
    layer0_outputs(2186) <= (inputs(37)) and not (inputs(1));
    layer0_outputs(2187) <= not((inputs(1)) or (inputs(43)));
    layer0_outputs(2188) <= not((inputs(162)) or (inputs(209)));
    layer0_outputs(2189) <= (inputs(106)) or (inputs(48));
    layer0_outputs(2190) <= (inputs(169)) and not (inputs(29));
    layer0_outputs(2191) <= not(inputs(117));
    layer0_outputs(2192) <= '0';
    layer0_outputs(2193) <= not(inputs(21)) or (inputs(222));
    layer0_outputs(2194) <= not(inputs(10)) or (inputs(209));
    layer0_outputs(2195) <= (inputs(225)) xor (inputs(71));
    layer0_outputs(2196) <= inputs(230);
    layer0_outputs(2197) <= inputs(218);
    layer0_outputs(2198) <= not(inputs(179));
    layer0_outputs(2199) <= '0';
    layer0_outputs(2200) <= inputs(132);
    layer0_outputs(2201) <= not((inputs(4)) or (inputs(45)));
    layer0_outputs(2202) <= inputs(117);
    layer0_outputs(2203) <= (inputs(130)) or (inputs(107));
    layer0_outputs(2204) <= not((inputs(245)) or (inputs(71)));
    layer0_outputs(2205) <= '1';
    layer0_outputs(2206) <= (inputs(21)) and not (inputs(51));
    layer0_outputs(2207) <= not(inputs(99));
    layer0_outputs(2208) <= '1';
    layer0_outputs(2209) <= (inputs(103)) or (inputs(190));
    layer0_outputs(2210) <= (inputs(193)) or (inputs(10));
    layer0_outputs(2211) <= not(inputs(122)) or (inputs(15));
    layer0_outputs(2212) <= not(inputs(211));
    layer0_outputs(2213) <= inputs(213);
    layer0_outputs(2214) <= not((inputs(18)) or (inputs(6)));
    layer0_outputs(2215) <= not((inputs(68)) or (inputs(66)));
    layer0_outputs(2216) <= not(inputs(129)) or (inputs(63));
    layer0_outputs(2217) <= not((inputs(252)) xor (inputs(5)));
    layer0_outputs(2218) <= (inputs(197)) or (inputs(104));
    layer0_outputs(2219) <= not((inputs(221)) or (inputs(0)));
    layer0_outputs(2220) <= not(inputs(95)) or (inputs(135));
    layer0_outputs(2221) <= not(inputs(216));
    layer0_outputs(2222) <= '0';
    layer0_outputs(2223) <= inputs(189);
    layer0_outputs(2224) <= not(inputs(182));
    layer0_outputs(2225) <= not(inputs(92));
    layer0_outputs(2226) <= not((inputs(9)) or (inputs(42)));
    layer0_outputs(2227) <= not((inputs(83)) or (inputs(181)));
    layer0_outputs(2228) <= '0';
    layer0_outputs(2229) <= inputs(182);
    layer0_outputs(2230) <= not((inputs(241)) or (inputs(245)));
    layer0_outputs(2231) <= not((inputs(45)) or (inputs(53)));
    layer0_outputs(2232) <= not(inputs(225));
    layer0_outputs(2233) <= '1';
    layer0_outputs(2234) <= not(inputs(119)) or (inputs(162));
    layer0_outputs(2235) <= (inputs(221)) or (inputs(136));
    layer0_outputs(2236) <= not(inputs(245));
    layer0_outputs(2237) <= not(inputs(146));
    layer0_outputs(2238) <= (inputs(23)) and not (inputs(130));
    layer0_outputs(2239) <= not(inputs(151)) or (inputs(209));
    layer0_outputs(2240) <= inputs(105);
    layer0_outputs(2241) <= inputs(190);
    layer0_outputs(2242) <= not((inputs(178)) or (inputs(189)));
    layer0_outputs(2243) <= (inputs(51)) xor (inputs(2));
    layer0_outputs(2244) <= inputs(180);
    layer0_outputs(2245) <= not((inputs(140)) or (inputs(85)));
    layer0_outputs(2246) <= not(inputs(87));
    layer0_outputs(2247) <= not(inputs(3)) or (inputs(162));
    layer0_outputs(2248) <= not(inputs(210));
    layer0_outputs(2249) <= not((inputs(86)) or (inputs(146)));
    layer0_outputs(2250) <= inputs(72);
    layer0_outputs(2251) <= not(inputs(240)) or (inputs(8));
    layer0_outputs(2252) <= not(inputs(18)) or (inputs(204));
    layer0_outputs(2253) <= not(inputs(6));
    layer0_outputs(2254) <= (inputs(120)) and not (inputs(52));
    layer0_outputs(2255) <= not(inputs(5));
    layer0_outputs(2256) <= not(inputs(86)) or (inputs(20));
    layer0_outputs(2257) <= (inputs(162)) or (inputs(179));
    layer0_outputs(2258) <= '1';
    layer0_outputs(2259) <= inputs(133);
    layer0_outputs(2260) <= inputs(233);
    layer0_outputs(2261) <= '0';
    layer0_outputs(2262) <= inputs(213);
    layer0_outputs(2263) <= not(inputs(203));
    layer0_outputs(2264) <= not((inputs(161)) or (inputs(70)));
    layer0_outputs(2265) <= not(inputs(125)) or (inputs(166));
    layer0_outputs(2266) <= (inputs(113)) or (inputs(211));
    layer0_outputs(2267) <= not(inputs(210));
    layer0_outputs(2268) <= not((inputs(251)) and (inputs(76)));
    layer0_outputs(2269) <= not((inputs(198)) and (inputs(232)));
    layer0_outputs(2270) <= inputs(190);
    layer0_outputs(2271) <= (inputs(127)) and (inputs(36));
    layer0_outputs(2272) <= not(inputs(118));
    layer0_outputs(2273) <= not((inputs(189)) or (inputs(134)));
    layer0_outputs(2274) <= inputs(132);
    layer0_outputs(2275) <= '1';
    layer0_outputs(2276) <= inputs(19);
    layer0_outputs(2277) <= not((inputs(25)) or (inputs(124)));
    layer0_outputs(2278) <= inputs(129);
    layer0_outputs(2279) <= (inputs(101)) and (inputs(123));
    layer0_outputs(2280) <= '0';
    layer0_outputs(2281) <= (inputs(108)) and not (inputs(114));
    layer0_outputs(2282) <= not(inputs(51)) or (inputs(111));
    layer0_outputs(2283) <= not(inputs(233));
    layer0_outputs(2284) <= inputs(177);
    layer0_outputs(2285) <= not((inputs(225)) or (inputs(228)));
    layer0_outputs(2286) <= not((inputs(204)) or (inputs(181)));
    layer0_outputs(2287) <= (inputs(157)) or (inputs(159));
    layer0_outputs(2288) <= inputs(183);
    layer0_outputs(2289) <= (inputs(118)) and not (inputs(72));
    layer0_outputs(2290) <= not((inputs(166)) or (inputs(218)));
    layer0_outputs(2291) <= not(inputs(130));
    layer0_outputs(2292) <= not(inputs(231));
    layer0_outputs(2293) <= not(inputs(99));
    layer0_outputs(2294) <= '0';
    layer0_outputs(2295) <= (inputs(149)) and not (inputs(190));
    layer0_outputs(2296) <= not(inputs(125));
    layer0_outputs(2297) <= inputs(176);
    layer0_outputs(2298) <= (inputs(224)) and (inputs(18));
    layer0_outputs(2299) <= inputs(112);
    layer0_outputs(2300) <= not(inputs(188));
    layer0_outputs(2301) <= not(inputs(117));
    layer0_outputs(2302) <= inputs(102);
    layer0_outputs(2303) <= (inputs(14)) and (inputs(84));
    layer0_outputs(2304) <= '0';
    layer0_outputs(2305) <= not(inputs(219)) or (inputs(48));
    layer0_outputs(2306) <= (inputs(47)) and not (inputs(241));
    layer0_outputs(2307) <= not((inputs(169)) and (inputs(195)));
    layer0_outputs(2308) <= (inputs(47)) or (inputs(74));
    layer0_outputs(2309) <= not((inputs(20)) or (inputs(32)));
    layer0_outputs(2310) <= not(inputs(78));
    layer0_outputs(2311) <= not(inputs(231)) or (inputs(0));
    layer0_outputs(2312) <= not(inputs(52)) or (inputs(155));
    layer0_outputs(2313) <= not(inputs(120)) or (inputs(204));
    layer0_outputs(2314) <= '0';
    layer0_outputs(2315) <= not(inputs(251)) or (inputs(50));
    layer0_outputs(2316) <= '1';
    layer0_outputs(2317) <= inputs(203);
    layer0_outputs(2318) <= (inputs(102)) and not (inputs(149));
    layer0_outputs(2319) <= not(inputs(198));
    layer0_outputs(2320) <= not(inputs(23)) or (inputs(200));
    layer0_outputs(2321) <= not(inputs(213)) or (inputs(179));
    layer0_outputs(2322) <= (inputs(245)) or (inputs(241));
    layer0_outputs(2323) <= inputs(166);
    layer0_outputs(2324) <= not(inputs(112));
    layer0_outputs(2325) <= (inputs(204)) or (inputs(217));
    layer0_outputs(2326) <= not(inputs(101));
    layer0_outputs(2327) <= not((inputs(127)) or (inputs(142)));
    layer0_outputs(2328) <= (inputs(138)) or (inputs(10));
    layer0_outputs(2329) <= (inputs(84)) or (inputs(20));
    layer0_outputs(2330) <= inputs(144);
    layer0_outputs(2331) <= not(inputs(251));
    layer0_outputs(2332) <= not((inputs(146)) or (inputs(102)));
    layer0_outputs(2333) <= not(inputs(116));
    layer0_outputs(2334) <= not((inputs(217)) xor (inputs(140)));
    layer0_outputs(2335) <= inputs(14);
    layer0_outputs(2336) <= (inputs(247)) and not (inputs(8));
    layer0_outputs(2337) <= not((inputs(68)) or (inputs(127)));
    layer0_outputs(2338) <= not(inputs(229)) or (inputs(96));
    layer0_outputs(2339) <= not((inputs(177)) or (inputs(199)));
    layer0_outputs(2340) <= inputs(53);
    layer0_outputs(2341) <= '0';
    layer0_outputs(2342) <= not(inputs(132)) or (inputs(184));
    layer0_outputs(2343) <= inputs(17);
    layer0_outputs(2344) <= not(inputs(140));
    layer0_outputs(2345) <= '1';
    layer0_outputs(2346) <= (inputs(195)) or (inputs(205));
    layer0_outputs(2347) <= not(inputs(82));
    layer0_outputs(2348) <= inputs(75);
    layer0_outputs(2349) <= (inputs(123)) or (inputs(178));
    layer0_outputs(2350) <= not((inputs(13)) xor (inputs(117)));
    layer0_outputs(2351) <= inputs(177);
    layer0_outputs(2352) <= not(inputs(164)) or (inputs(81));
    layer0_outputs(2353) <= (inputs(186)) or (inputs(221));
    layer0_outputs(2354) <= not((inputs(137)) and (inputs(203)));
    layer0_outputs(2355) <= not((inputs(217)) or (inputs(159)));
    layer0_outputs(2356) <= not(inputs(197)) or (inputs(30));
    layer0_outputs(2357) <= not((inputs(179)) or (inputs(8)));
    layer0_outputs(2358) <= not((inputs(115)) and (inputs(133)));
    layer0_outputs(2359) <= (inputs(132)) xor (inputs(34));
    layer0_outputs(2360) <= (inputs(242)) and (inputs(92));
    layer0_outputs(2361) <= not(inputs(182));
    layer0_outputs(2362) <= (inputs(120)) and not (inputs(197));
    layer0_outputs(2363) <= not(inputs(176));
    layer0_outputs(2364) <= inputs(167);
    layer0_outputs(2365) <= not((inputs(203)) or (inputs(6)));
    layer0_outputs(2366) <= (inputs(150)) xor (inputs(135));
    layer0_outputs(2367) <= (inputs(112)) and not (inputs(196));
    layer0_outputs(2368) <= not(inputs(110)) or (inputs(40));
    layer0_outputs(2369) <= (inputs(89)) and not (inputs(239));
    layer0_outputs(2370) <= inputs(117);
    layer0_outputs(2371) <= (inputs(175)) and (inputs(12));
    layer0_outputs(2372) <= not(inputs(25));
    layer0_outputs(2373) <= (inputs(91)) or (inputs(37));
    layer0_outputs(2374) <= not((inputs(149)) xor (inputs(167)));
    layer0_outputs(2375) <= (inputs(7)) and not (inputs(141));
    layer0_outputs(2376) <= (inputs(113)) or (inputs(112));
    layer0_outputs(2377) <= (inputs(65)) or (inputs(236));
    layer0_outputs(2378) <= not(inputs(59)) or (inputs(75));
    layer0_outputs(2379) <= not((inputs(118)) or (inputs(74)));
    layer0_outputs(2380) <= not(inputs(25));
    layer0_outputs(2381) <= inputs(147);
    layer0_outputs(2382) <= (inputs(168)) and (inputs(143));
    layer0_outputs(2383) <= '1';
    layer0_outputs(2384) <= not((inputs(172)) and (inputs(198)));
    layer0_outputs(2385) <= (inputs(23)) and not (inputs(192));
    layer0_outputs(2386) <= not(inputs(92));
    layer0_outputs(2387) <= not((inputs(184)) or (inputs(116)));
    layer0_outputs(2388) <= inputs(91);
    layer0_outputs(2389) <= not((inputs(110)) or (inputs(111)));
    layer0_outputs(2390) <= inputs(93);
    layer0_outputs(2391) <= inputs(147);
    layer0_outputs(2392) <= (inputs(51)) or (inputs(94));
    layer0_outputs(2393) <= inputs(80);
    layer0_outputs(2394) <= inputs(106);
    layer0_outputs(2395) <= (inputs(145)) and (inputs(143));
    layer0_outputs(2396) <= not((inputs(253)) and (inputs(136)));
    layer0_outputs(2397) <= not(inputs(190)) or (inputs(87));
    layer0_outputs(2398) <= '1';
    layer0_outputs(2399) <= inputs(195);
    layer0_outputs(2400) <= '0';
    layer0_outputs(2401) <= (inputs(181)) or (inputs(165));
    layer0_outputs(2402) <= '1';
    layer0_outputs(2403) <= not(inputs(100)) or (inputs(16));
    layer0_outputs(2404) <= not(inputs(247)) or (inputs(15));
    layer0_outputs(2405) <= not(inputs(102)) or (inputs(252));
    layer0_outputs(2406) <= (inputs(168)) and not (inputs(57));
    layer0_outputs(2407) <= not(inputs(238)) or (inputs(252));
    layer0_outputs(2408) <= not(inputs(8)) or (inputs(8));
    layer0_outputs(2409) <= (inputs(124)) and not (inputs(161));
    layer0_outputs(2410) <= not((inputs(35)) xor (inputs(145)));
    layer0_outputs(2411) <= inputs(30);
    layer0_outputs(2412) <= (inputs(255)) and (inputs(129));
    layer0_outputs(2413) <= not(inputs(116)) or (inputs(189));
    layer0_outputs(2414) <= inputs(182);
    layer0_outputs(2415) <= not((inputs(247)) or (inputs(132)));
    layer0_outputs(2416) <= '1';
    layer0_outputs(2417) <= not(inputs(181));
    layer0_outputs(2418) <= not((inputs(24)) or (inputs(207)));
    layer0_outputs(2419) <= not(inputs(101));
    layer0_outputs(2420) <= not(inputs(147));
    layer0_outputs(2421) <= not(inputs(210));
    layer0_outputs(2422) <= inputs(239);
    layer0_outputs(2423) <= not(inputs(168));
    layer0_outputs(2424) <= not(inputs(110));
    layer0_outputs(2425) <= (inputs(79)) and not (inputs(185));
    layer0_outputs(2426) <= not((inputs(60)) or (inputs(209)));
    layer0_outputs(2427) <= inputs(63);
    layer0_outputs(2428) <= '1';
    layer0_outputs(2429) <= inputs(168);
    layer0_outputs(2430) <= inputs(55);
    layer0_outputs(2431) <= not((inputs(19)) or (inputs(122)));
    layer0_outputs(2432) <= not(inputs(40)) or (inputs(140));
    layer0_outputs(2433) <= inputs(23);
    layer0_outputs(2434) <= (inputs(49)) and (inputs(133));
    layer0_outputs(2435) <= (inputs(100)) and not (inputs(211));
    layer0_outputs(2436) <= '1';
    layer0_outputs(2437) <= not(inputs(158));
    layer0_outputs(2438) <= not((inputs(37)) or (inputs(248)));
    layer0_outputs(2439) <= (inputs(97)) or (inputs(179));
    layer0_outputs(2440) <= inputs(212);
    layer0_outputs(2441) <= not(inputs(147));
    layer0_outputs(2442) <= (inputs(188)) and (inputs(140));
    layer0_outputs(2443) <= inputs(25);
    layer0_outputs(2444) <= (inputs(220)) or (inputs(73));
    layer0_outputs(2445) <= not(inputs(150));
    layer0_outputs(2446) <= not((inputs(191)) or (inputs(19)));
    layer0_outputs(2447) <= (inputs(32)) or (inputs(175));
    layer0_outputs(2448) <= '0';
    layer0_outputs(2449) <= (inputs(68)) and not (inputs(4));
    layer0_outputs(2450) <= (inputs(16)) and not (inputs(136));
    layer0_outputs(2451) <= not((inputs(57)) and (inputs(214)));
    layer0_outputs(2452) <= (inputs(46)) and not (inputs(92));
    layer0_outputs(2453) <= not(inputs(202)) or (inputs(114));
    layer0_outputs(2454) <= (inputs(86)) or (inputs(172));
    layer0_outputs(2455) <= inputs(250);
    layer0_outputs(2456) <= inputs(117);
    layer0_outputs(2457) <= not((inputs(45)) and (inputs(148)));
    layer0_outputs(2458) <= (inputs(89)) and (inputs(11));
    layer0_outputs(2459) <= inputs(69);
    layer0_outputs(2460) <= (inputs(46)) and not (inputs(12));
    layer0_outputs(2461) <= not((inputs(191)) or (inputs(153)));
    layer0_outputs(2462) <= not(inputs(42));
    layer0_outputs(2463) <= not(inputs(219));
    layer0_outputs(2464) <= (inputs(168)) and (inputs(109));
    layer0_outputs(2465) <= (inputs(92)) and not (inputs(165));
    layer0_outputs(2466) <= not((inputs(146)) and (inputs(238)));
    layer0_outputs(2467) <= not((inputs(182)) and (inputs(239)));
    layer0_outputs(2468) <= not(inputs(53)) or (inputs(18));
    layer0_outputs(2469) <= not(inputs(119));
    layer0_outputs(2470) <= (inputs(255)) or (inputs(7));
    layer0_outputs(2471) <= (inputs(2)) or (inputs(220));
    layer0_outputs(2472) <= not(inputs(135));
    layer0_outputs(2473) <= (inputs(178)) or (inputs(222));
    layer0_outputs(2474) <= not((inputs(129)) and (inputs(56)));
    layer0_outputs(2475) <= (inputs(194)) or (inputs(170));
    layer0_outputs(2476) <= (inputs(94)) and not (inputs(125));
    layer0_outputs(2477) <= (inputs(153)) or (inputs(119));
    layer0_outputs(2478) <= inputs(92);
    layer0_outputs(2479) <= inputs(77);
    layer0_outputs(2480) <= (inputs(128)) and (inputs(11));
    layer0_outputs(2481) <= not(inputs(94)) or (inputs(37));
    layer0_outputs(2482) <= (inputs(138)) and not (inputs(164));
    layer0_outputs(2483) <= not(inputs(75));
    layer0_outputs(2484) <= inputs(43);
    layer0_outputs(2485) <= not(inputs(106));
    layer0_outputs(2486) <= (inputs(59)) and not (inputs(223));
    layer0_outputs(2487) <= inputs(191);
    layer0_outputs(2488) <= (inputs(164)) or (inputs(100));
    layer0_outputs(2489) <= (inputs(212)) and not (inputs(105));
    layer0_outputs(2490) <= (inputs(175)) and not (inputs(173));
    layer0_outputs(2491) <= (inputs(204)) or (inputs(224));
    layer0_outputs(2492) <= (inputs(139)) xor (inputs(105));
    layer0_outputs(2493) <= inputs(183);
    layer0_outputs(2494) <= (inputs(13)) and not (inputs(29));
    layer0_outputs(2495) <= not((inputs(41)) or (inputs(54)));
    layer0_outputs(2496) <= '0';
    layer0_outputs(2497) <= not(inputs(135));
    layer0_outputs(2498) <= not(inputs(153));
    layer0_outputs(2499) <= not((inputs(104)) or (inputs(14)));
    layer0_outputs(2500) <= (inputs(246)) or (inputs(147));
    layer0_outputs(2501) <= inputs(177);
    layer0_outputs(2502) <= not(inputs(117));
    layer0_outputs(2503) <= not(inputs(234));
    layer0_outputs(2504) <= inputs(85);
    layer0_outputs(2505) <= (inputs(0)) or (inputs(94));
    layer0_outputs(2506) <= not((inputs(218)) xor (inputs(218)));
    layer0_outputs(2507) <= inputs(228);
    layer0_outputs(2508) <= not((inputs(69)) and (inputs(201)));
    layer0_outputs(2509) <= '1';
    layer0_outputs(2510) <= inputs(102);
    layer0_outputs(2511) <= not(inputs(130));
    layer0_outputs(2512) <= inputs(76);
    layer0_outputs(2513) <= (inputs(47)) or (inputs(30));
    layer0_outputs(2514) <= (inputs(76)) and not (inputs(216));
    layer0_outputs(2515) <= not(inputs(73));
    layer0_outputs(2516) <= (inputs(155)) or (inputs(51));
    layer0_outputs(2517) <= inputs(75);
    layer0_outputs(2518) <= not((inputs(80)) xor (inputs(33)));
    layer0_outputs(2519) <= not(inputs(108));
    layer0_outputs(2520) <= (inputs(49)) and not (inputs(2));
    layer0_outputs(2521) <= '1';
    layer0_outputs(2522) <= (inputs(173)) or (inputs(216));
    layer0_outputs(2523) <= '1';
    layer0_outputs(2524) <= inputs(186);
    layer0_outputs(2525) <= (inputs(123)) or (inputs(137));
    layer0_outputs(2526) <= '0';
    layer0_outputs(2527) <= inputs(90);
    layer0_outputs(2528) <= (inputs(58)) xor (inputs(45));
    layer0_outputs(2529) <= (inputs(48)) or (inputs(226));
    layer0_outputs(2530) <= inputs(164);
    layer0_outputs(2531) <= (inputs(40)) xor (inputs(130));
    layer0_outputs(2532) <= (inputs(96)) xor (inputs(24));
    layer0_outputs(2533) <= (inputs(138)) and not (inputs(77));
    layer0_outputs(2534) <= (inputs(213)) or (inputs(87));
    layer0_outputs(2535) <= not(inputs(233)) or (inputs(144));
    layer0_outputs(2536) <= not(inputs(218));
    layer0_outputs(2537) <= (inputs(100)) or (inputs(193));
    layer0_outputs(2538) <= inputs(53);
    layer0_outputs(2539) <= not(inputs(42)) or (inputs(147));
    layer0_outputs(2540) <= (inputs(100)) or (inputs(132));
    layer0_outputs(2541) <= (inputs(160)) or (inputs(133));
    layer0_outputs(2542) <= not(inputs(232)) or (inputs(1));
    layer0_outputs(2543) <= not(inputs(17)) or (inputs(160));
    layer0_outputs(2544) <= not(inputs(93));
    layer0_outputs(2545) <= (inputs(66)) or (inputs(141));
    layer0_outputs(2546) <= not(inputs(231));
    layer0_outputs(2547) <= inputs(122);
    layer0_outputs(2548) <= not(inputs(112));
    layer0_outputs(2549) <= inputs(60);
    layer0_outputs(2550) <= not((inputs(228)) or (inputs(117)));
    layer0_outputs(2551) <= '0';
    layer0_outputs(2552) <= not(inputs(242)) or (inputs(28));
    layer0_outputs(2553) <= '1';
    layer0_outputs(2554) <= not(inputs(212)) or (inputs(1));
    layer0_outputs(2555) <= inputs(154);
    layer0_outputs(2556) <= not(inputs(129)) or (inputs(191));
    layer0_outputs(2557) <= (inputs(28)) and (inputs(191));
    layer0_outputs(2558) <= inputs(124);
    layer0_outputs(2559) <= not(inputs(61));
    layer1_outputs(0) <= (layer0_outputs(2044)) xor (layer0_outputs(1605));
    layer1_outputs(1) <= (layer0_outputs(232)) or (layer0_outputs(455));
    layer1_outputs(2) <= not(layer0_outputs(482));
    layer1_outputs(3) <= layer0_outputs(1724);
    layer1_outputs(4) <= '0';
    layer1_outputs(5) <= not((layer0_outputs(2457)) and (layer0_outputs(1336)));
    layer1_outputs(6) <= not((layer0_outputs(2334)) and (layer0_outputs(2463)));
    layer1_outputs(7) <= '1';
    layer1_outputs(8) <= not(layer0_outputs(216)) or (layer0_outputs(1705));
    layer1_outputs(9) <= not(layer0_outputs(218));
    layer1_outputs(10) <= (layer0_outputs(1788)) and not (layer0_outputs(1390));
    layer1_outputs(11) <= not((layer0_outputs(1927)) and (layer0_outputs(1214)));
    layer1_outputs(12) <= not(layer0_outputs(1656)) or (layer0_outputs(1524));
    layer1_outputs(13) <= not(layer0_outputs(283));
    layer1_outputs(14) <= (layer0_outputs(2440)) and not (layer0_outputs(1374));
    layer1_outputs(15) <= not(layer0_outputs(715));
    layer1_outputs(16) <= (layer0_outputs(1789)) or (layer0_outputs(665));
    layer1_outputs(17) <= not(layer0_outputs(616));
    layer1_outputs(18) <= (layer0_outputs(2548)) and not (layer0_outputs(2098));
    layer1_outputs(19) <= (layer0_outputs(208)) and not (layer0_outputs(177));
    layer1_outputs(20) <= '1';
    layer1_outputs(21) <= layer0_outputs(1096);
    layer1_outputs(22) <= layer0_outputs(2183);
    layer1_outputs(23) <= (layer0_outputs(696)) and not (layer0_outputs(1980));
    layer1_outputs(24) <= layer0_outputs(2332);
    layer1_outputs(25) <= layer0_outputs(37);
    layer1_outputs(26) <= layer0_outputs(2165);
    layer1_outputs(27) <= (layer0_outputs(1279)) and not (layer0_outputs(847));
    layer1_outputs(28) <= not(layer0_outputs(1669));
    layer1_outputs(29) <= (layer0_outputs(1662)) and not (layer0_outputs(706));
    layer1_outputs(30) <= '1';
    layer1_outputs(31) <= '1';
    layer1_outputs(32) <= layer0_outputs(664);
    layer1_outputs(33) <= not(layer0_outputs(1147));
    layer1_outputs(34) <= (layer0_outputs(334)) or (layer0_outputs(2221));
    layer1_outputs(35) <= '0';
    layer1_outputs(36) <= (layer0_outputs(583)) and not (layer0_outputs(282));
    layer1_outputs(37) <= layer0_outputs(2027);
    layer1_outputs(38) <= not(layer0_outputs(593)) or (layer0_outputs(92));
    layer1_outputs(39) <= not(layer0_outputs(1318)) or (layer0_outputs(301));
    layer1_outputs(40) <= not((layer0_outputs(1460)) or (layer0_outputs(596)));
    layer1_outputs(41) <= layer0_outputs(1664);
    layer1_outputs(42) <= layer0_outputs(1487);
    layer1_outputs(43) <= not(layer0_outputs(932));
    layer1_outputs(44) <= '1';
    layer1_outputs(45) <= layer0_outputs(33);
    layer1_outputs(46) <= '1';
    layer1_outputs(47) <= layer0_outputs(2121);
    layer1_outputs(48) <= not(layer0_outputs(537));
    layer1_outputs(49) <= not(layer0_outputs(945));
    layer1_outputs(50) <= (layer0_outputs(2183)) and not (layer0_outputs(1767));
    layer1_outputs(51) <= not(layer0_outputs(269));
    layer1_outputs(52) <= not((layer0_outputs(1984)) or (layer0_outputs(175)));
    layer1_outputs(53) <= not(layer0_outputs(1319));
    layer1_outputs(54) <= not((layer0_outputs(2141)) and (layer0_outputs(769)));
    layer1_outputs(55) <= not((layer0_outputs(754)) and (layer0_outputs(2552)));
    layer1_outputs(56) <= (layer0_outputs(1197)) or (layer0_outputs(1974));
    layer1_outputs(57) <= not((layer0_outputs(1324)) and (layer0_outputs(2403)));
    layer1_outputs(58) <= not(layer0_outputs(1477));
    layer1_outputs(59) <= not((layer0_outputs(1257)) and (layer0_outputs(1419)));
    layer1_outputs(60) <= (layer0_outputs(946)) xor (layer0_outputs(1736));
    layer1_outputs(61) <= '1';
    layer1_outputs(62) <= not(layer0_outputs(1647));
    layer1_outputs(63) <= layer0_outputs(2482);
    layer1_outputs(64) <= layer0_outputs(653);
    layer1_outputs(65) <= not((layer0_outputs(2467)) and (layer0_outputs(1165)));
    layer1_outputs(66) <= layer0_outputs(2262);
    layer1_outputs(67) <= (layer0_outputs(1525)) and (layer0_outputs(2130));
    layer1_outputs(68) <= layer0_outputs(1610);
    layer1_outputs(69) <= not(layer0_outputs(2263)) or (layer0_outputs(18));
    layer1_outputs(70) <= not((layer0_outputs(2278)) or (layer0_outputs(2063)));
    layer1_outputs(71) <= not(layer0_outputs(2205)) or (layer0_outputs(1309));
    layer1_outputs(72) <= layer0_outputs(340);
    layer1_outputs(73) <= (layer0_outputs(623)) or (layer0_outputs(2030));
    layer1_outputs(74) <= not(layer0_outputs(2139));
    layer1_outputs(75) <= (layer0_outputs(1712)) or (layer0_outputs(916));
    layer1_outputs(76) <= not((layer0_outputs(534)) and (layer0_outputs(1114)));
    layer1_outputs(77) <= (layer0_outputs(1377)) and not (layer0_outputs(1127));
    layer1_outputs(78) <= not(layer0_outputs(172)) or (layer0_outputs(1787));
    layer1_outputs(79) <= not((layer0_outputs(1450)) and (layer0_outputs(1274)));
    layer1_outputs(80) <= not((layer0_outputs(2410)) or (layer0_outputs(2481)));
    layer1_outputs(81) <= not(layer0_outputs(548)) or (layer0_outputs(460));
    layer1_outputs(82) <= layer0_outputs(1838);
    layer1_outputs(83) <= layer0_outputs(2212);
    layer1_outputs(84) <= not(layer0_outputs(1514)) or (layer0_outputs(2525));
    layer1_outputs(85) <= not(layer0_outputs(582)) or (layer0_outputs(178));
    layer1_outputs(86) <= not(layer0_outputs(479));
    layer1_outputs(87) <= not((layer0_outputs(953)) or (layer0_outputs(1933)));
    layer1_outputs(88) <= layer0_outputs(699);
    layer1_outputs(89) <= not(layer0_outputs(1678));
    layer1_outputs(90) <= layer0_outputs(2372);
    layer1_outputs(91) <= not((layer0_outputs(542)) xor (layer0_outputs(1427)));
    layer1_outputs(92) <= layer0_outputs(192);
    layer1_outputs(93) <= not((layer0_outputs(917)) or (layer0_outputs(356)));
    layer1_outputs(94) <= not(layer0_outputs(357)) or (layer0_outputs(237));
    layer1_outputs(95) <= not((layer0_outputs(338)) and (layer0_outputs(163)));
    layer1_outputs(96) <= not(layer0_outputs(1416));
    layer1_outputs(97) <= (layer0_outputs(129)) and (layer0_outputs(2254));
    layer1_outputs(98) <= '0';
    layer1_outputs(99) <= (layer0_outputs(301)) and not (layer0_outputs(1318));
    layer1_outputs(100) <= not(layer0_outputs(1981));
    layer1_outputs(101) <= (layer0_outputs(1928)) and not (layer0_outputs(1367));
    layer1_outputs(102) <= (layer0_outputs(1837)) and not (layer0_outputs(681));
    layer1_outputs(103) <= not((layer0_outputs(24)) and (layer0_outputs(1843)));
    layer1_outputs(104) <= (layer0_outputs(459)) xor (layer0_outputs(1653));
    layer1_outputs(105) <= (layer0_outputs(404)) and (layer0_outputs(140));
    layer1_outputs(106) <= not(layer0_outputs(1686));
    layer1_outputs(107) <= (layer0_outputs(2076)) and (layer0_outputs(1485));
    layer1_outputs(108) <= not((layer0_outputs(2310)) and (layer0_outputs(831)));
    layer1_outputs(109) <= not(layer0_outputs(2257));
    layer1_outputs(110) <= '0';
    layer1_outputs(111) <= not(layer0_outputs(1272));
    layer1_outputs(112) <= layer0_outputs(2451);
    layer1_outputs(113) <= (layer0_outputs(802)) and (layer0_outputs(2337));
    layer1_outputs(114) <= '0';
    layer1_outputs(115) <= (layer0_outputs(2454)) and (layer0_outputs(2441));
    layer1_outputs(116) <= not(layer0_outputs(2495)) or (layer0_outputs(371));
    layer1_outputs(117) <= not(layer0_outputs(484)) or (layer0_outputs(119));
    layer1_outputs(118) <= layer0_outputs(2180);
    layer1_outputs(119) <= (layer0_outputs(1954)) and not (layer0_outputs(912));
    layer1_outputs(120) <= (layer0_outputs(2041)) and not (layer0_outputs(1943));
    layer1_outputs(121) <= not(layer0_outputs(1359)) or (layer0_outputs(1382));
    layer1_outputs(122) <= not(layer0_outputs(322));
    layer1_outputs(123) <= not((layer0_outputs(1637)) or (layer0_outputs(747)));
    layer1_outputs(124) <= (layer0_outputs(2357)) and (layer0_outputs(1187));
    layer1_outputs(125) <= not(layer0_outputs(983));
    layer1_outputs(126) <= layer0_outputs(1221);
    layer1_outputs(127) <= not(layer0_outputs(1478));
    layer1_outputs(128) <= '1';
    layer1_outputs(129) <= (layer0_outputs(478)) and not (layer0_outputs(1674));
    layer1_outputs(130) <= not((layer0_outputs(409)) xor (layer0_outputs(1975)));
    layer1_outputs(131) <= not((layer0_outputs(806)) and (layer0_outputs(930)));
    layer1_outputs(132) <= not(layer0_outputs(2370));
    layer1_outputs(133) <= layer0_outputs(179);
    layer1_outputs(134) <= not(layer0_outputs(1861));
    layer1_outputs(135) <= not(layer0_outputs(554));
    layer1_outputs(136) <= not(layer0_outputs(220));
    layer1_outputs(137) <= layer0_outputs(2292);
    layer1_outputs(138) <= not(layer0_outputs(1538));
    layer1_outputs(139) <= not(layer0_outputs(1566)) or (layer0_outputs(292));
    layer1_outputs(140) <= (layer0_outputs(1772)) and not (layer0_outputs(1844));
    layer1_outputs(141) <= '0';
    layer1_outputs(142) <= not((layer0_outputs(1329)) or (layer0_outputs(1379)));
    layer1_outputs(143) <= not(layer0_outputs(336));
    layer1_outputs(144) <= not(layer0_outputs(1707));
    layer1_outputs(145) <= (layer0_outputs(555)) or (layer0_outputs(771));
    layer1_outputs(146) <= layer0_outputs(1299);
    layer1_outputs(147) <= not((layer0_outputs(243)) xor (layer0_outputs(1349)));
    layer1_outputs(148) <= not(layer0_outputs(2185)) or (layer0_outputs(1177));
    layer1_outputs(149) <= layer0_outputs(358);
    layer1_outputs(150) <= '1';
    layer1_outputs(151) <= not(layer0_outputs(1713));
    layer1_outputs(152) <= layer0_outputs(46);
    layer1_outputs(153) <= not(layer0_outputs(1175));
    layer1_outputs(154) <= (layer0_outputs(2109)) and not (layer0_outputs(321));
    layer1_outputs(155) <= not(layer0_outputs(730));
    layer1_outputs(156) <= (layer0_outputs(1418)) and not (layer0_outputs(1));
    layer1_outputs(157) <= layer0_outputs(1619);
    layer1_outputs(158) <= layer0_outputs(1664);
    layer1_outputs(159) <= (layer0_outputs(1875)) and not (layer0_outputs(2149));
    layer1_outputs(160) <= not((layer0_outputs(884)) or (layer0_outputs(757)));
    layer1_outputs(161) <= not(layer0_outputs(1134)) or (layer0_outputs(252));
    layer1_outputs(162) <= not(layer0_outputs(1861)) or (layer0_outputs(1209));
    layer1_outputs(163) <= (layer0_outputs(1495)) and not (layer0_outputs(2517));
    layer1_outputs(164) <= (layer0_outputs(2446)) and not (layer0_outputs(412));
    layer1_outputs(165) <= not(layer0_outputs(568)) or (layer0_outputs(1509));
    layer1_outputs(166) <= not(layer0_outputs(1599)) or (layer0_outputs(509));
    layer1_outputs(167) <= not((layer0_outputs(2443)) xor (layer0_outputs(288)));
    layer1_outputs(168) <= layer0_outputs(794);
    layer1_outputs(169) <= not(layer0_outputs(2432));
    layer1_outputs(170) <= '0';
    layer1_outputs(171) <= (layer0_outputs(2273)) and (layer0_outputs(992));
    layer1_outputs(172) <= not(layer0_outputs(592));
    layer1_outputs(173) <= (layer0_outputs(2090)) and (layer0_outputs(2553));
    layer1_outputs(174) <= not(layer0_outputs(794));
    layer1_outputs(175) <= not((layer0_outputs(1872)) and (layer0_outputs(1533)));
    layer1_outputs(176) <= layer0_outputs(1306);
    layer1_outputs(177) <= not((layer0_outputs(279)) and (layer0_outputs(1826)));
    layer1_outputs(178) <= not(layer0_outputs(184)) or (layer0_outputs(951));
    layer1_outputs(179) <= layer0_outputs(2515);
    layer1_outputs(180) <= (layer0_outputs(137)) and (layer0_outputs(770));
    layer1_outputs(181) <= not(layer0_outputs(711)) or (layer0_outputs(2524));
    layer1_outputs(182) <= (layer0_outputs(1850)) and not (layer0_outputs(997));
    layer1_outputs(183) <= '1';
    layer1_outputs(184) <= not(layer0_outputs(284));
    layer1_outputs(185) <= '1';
    layer1_outputs(186) <= layer0_outputs(2308);
    layer1_outputs(187) <= layer0_outputs(853);
    layer1_outputs(188) <= not(layer0_outputs(1088)) or (layer0_outputs(281));
    layer1_outputs(189) <= not(layer0_outputs(1361)) or (layer0_outputs(50));
    layer1_outputs(190) <= not((layer0_outputs(1825)) or (layer0_outputs(2325)));
    layer1_outputs(191) <= (layer0_outputs(2008)) and not (layer0_outputs(477));
    layer1_outputs(192) <= layer0_outputs(2126);
    layer1_outputs(193) <= (layer0_outputs(587)) and not (layer0_outputs(235));
    layer1_outputs(194) <= layer0_outputs(716);
    layer1_outputs(195) <= (layer0_outputs(1479)) and (layer0_outputs(809));
    layer1_outputs(196) <= not(layer0_outputs(324));
    layer1_outputs(197) <= (layer0_outputs(1506)) and not (layer0_outputs(261));
    layer1_outputs(198) <= not((layer0_outputs(171)) and (layer0_outputs(970)));
    layer1_outputs(199) <= not(layer0_outputs(1432));
    layer1_outputs(200) <= not((layer0_outputs(1046)) and (layer0_outputs(1752)));
    layer1_outputs(201) <= (layer0_outputs(1394)) and not (layer0_outputs(1098));
    layer1_outputs(202) <= (layer0_outputs(1165)) and not (layer0_outputs(591));
    layer1_outputs(203) <= not(layer0_outputs(926));
    layer1_outputs(204) <= not((layer0_outputs(673)) and (layer0_outputs(2361)));
    layer1_outputs(205) <= not(layer0_outputs(117));
    layer1_outputs(206) <= not(layer0_outputs(994));
    layer1_outputs(207) <= layer0_outputs(1142);
    layer1_outputs(208) <= layer0_outputs(1124);
    layer1_outputs(209) <= not(layer0_outputs(181));
    layer1_outputs(210) <= not((layer0_outputs(2541)) and (layer0_outputs(906)));
    layer1_outputs(211) <= '0';
    layer1_outputs(212) <= not(layer0_outputs(2396)) or (layer0_outputs(2071));
    layer1_outputs(213) <= (layer0_outputs(114)) or (layer0_outputs(1799));
    layer1_outputs(214) <= (layer0_outputs(832)) and not (layer0_outputs(2253));
    layer1_outputs(215) <= not(layer0_outputs(1760));
    layer1_outputs(216) <= layer0_outputs(2559);
    layer1_outputs(217) <= not((layer0_outputs(387)) and (layer0_outputs(207)));
    layer1_outputs(218) <= '0';
    layer1_outputs(219) <= layer0_outputs(631);
    layer1_outputs(220) <= (layer0_outputs(1260)) and (layer0_outputs(1747));
    layer1_outputs(221) <= not(layer0_outputs(1512));
    layer1_outputs(222) <= not(layer0_outputs(1126)) or (layer0_outputs(229));
    layer1_outputs(223) <= not(layer0_outputs(2336)) or (layer0_outputs(1549));
    layer1_outputs(224) <= not(layer0_outputs(1129));
    layer1_outputs(225) <= (layer0_outputs(1194)) and (layer0_outputs(75));
    layer1_outputs(226) <= '0';
    layer1_outputs(227) <= layer0_outputs(1956);
    layer1_outputs(228) <= layer0_outputs(299);
    layer1_outputs(229) <= '0';
    layer1_outputs(230) <= not(layer0_outputs(2523));
    layer1_outputs(231) <= layer0_outputs(2037);
    layer1_outputs(232) <= not((layer0_outputs(1577)) and (layer0_outputs(1555)));
    layer1_outputs(233) <= '1';
    layer1_outputs(234) <= not(layer0_outputs(736));
    layer1_outputs(235) <= layer0_outputs(2088);
    layer1_outputs(236) <= (layer0_outputs(483)) or (layer0_outputs(1557));
    layer1_outputs(237) <= not(layer0_outputs(47));
    layer1_outputs(238) <= (layer0_outputs(2152)) and (layer0_outputs(65));
    layer1_outputs(239) <= (layer0_outputs(1786)) xor (layer0_outputs(223));
    layer1_outputs(240) <= not(layer0_outputs(368));
    layer1_outputs(241) <= not(layer0_outputs(602));
    layer1_outputs(242) <= layer0_outputs(518);
    layer1_outputs(243) <= (layer0_outputs(1168)) or (layer0_outputs(2276));
    layer1_outputs(244) <= layer0_outputs(1042);
    layer1_outputs(245) <= (layer0_outputs(2389)) and (layer0_outputs(265));
    layer1_outputs(246) <= not(layer0_outputs(2539));
    layer1_outputs(247) <= (layer0_outputs(1453)) and (layer0_outputs(2085));
    layer1_outputs(248) <= not(layer0_outputs(2524)) or (layer0_outputs(1828));
    layer1_outputs(249) <= '1';
    layer1_outputs(250) <= '0';
    layer1_outputs(251) <= layer0_outputs(1640);
    layer1_outputs(252) <= not(layer0_outputs(740)) or (layer0_outputs(2550));
    layer1_outputs(253) <= not(layer0_outputs(1263));
    layer1_outputs(254) <= not((layer0_outputs(946)) and (layer0_outputs(1066)));
    layer1_outputs(255) <= not(layer0_outputs(885)) or (layer0_outputs(2284));
    layer1_outputs(256) <= (layer0_outputs(525)) or (layer0_outputs(907));
    layer1_outputs(257) <= not(layer0_outputs(1695));
    layer1_outputs(258) <= not((layer0_outputs(2448)) or (layer0_outputs(230)));
    layer1_outputs(259) <= not(layer0_outputs(2131));
    layer1_outputs(260) <= layer0_outputs(757);
    layer1_outputs(261) <= not(layer0_outputs(2498));
    layer1_outputs(262) <= not((layer0_outputs(1793)) and (layer0_outputs(1043)));
    layer1_outputs(263) <= not(layer0_outputs(60)) or (layer0_outputs(1144));
    layer1_outputs(264) <= '0';
    layer1_outputs(265) <= (layer0_outputs(447)) and not (layer0_outputs(2011));
    layer1_outputs(266) <= not((layer0_outputs(1258)) or (layer0_outputs(943)));
    layer1_outputs(267) <= not(layer0_outputs(1904));
    layer1_outputs(268) <= not(layer0_outputs(2103)) or (layer0_outputs(1118));
    layer1_outputs(269) <= not(layer0_outputs(1059));
    layer1_outputs(270) <= (layer0_outputs(347)) and not (layer0_outputs(1782));
    layer1_outputs(271) <= not(layer0_outputs(597));
    layer1_outputs(272) <= layer0_outputs(2224);
    layer1_outputs(273) <= layer0_outputs(2423);
    layer1_outputs(274) <= (layer0_outputs(75)) or (layer0_outputs(456));
    layer1_outputs(275) <= not((layer0_outputs(705)) or (layer0_outputs(858)));
    layer1_outputs(276) <= layer0_outputs(196);
    layer1_outputs(277) <= (layer0_outputs(109)) and not (layer0_outputs(1776));
    layer1_outputs(278) <= (layer0_outputs(1068)) and (layer0_outputs(1966));
    layer1_outputs(279) <= not(layer0_outputs(1816)) or (layer0_outputs(1986));
    layer1_outputs(280) <= not(layer0_outputs(967)) or (layer0_outputs(574));
    layer1_outputs(281) <= (layer0_outputs(1031)) and (layer0_outputs(325));
    layer1_outputs(282) <= not(layer0_outputs(179));
    layer1_outputs(283) <= (layer0_outputs(1099)) and not (layer0_outputs(1111));
    layer1_outputs(284) <= not((layer0_outputs(1280)) xor (layer0_outputs(1001)));
    layer1_outputs(285) <= (layer0_outputs(706)) xor (layer0_outputs(1925));
    layer1_outputs(286) <= '1';
    layer1_outputs(287) <= not(layer0_outputs(82)) or (layer0_outputs(87));
    layer1_outputs(288) <= not(layer0_outputs(1212));
    layer1_outputs(289) <= layer0_outputs(2355);
    layer1_outputs(290) <= not(layer0_outputs(2253));
    layer1_outputs(291) <= not(layer0_outputs(1645));
    layer1_outputs(292) <= layer0_outputs(244);
    layer1_outputs(293) <= not(layer0_outputs(2462));
    layer1_outputs(294) <= layer0_outputs(915);
    layer1_outputs(295) <= (layer0_outputs(376)) or (layer0_outputs(2018));
    layer1_outputs(296) <= '0';
    layer1_outputs(297) <= (layer0_outputs(1473)) and not (layer0_outputs(571));
    layer1_outputs(298) <= not(layer0_outputs(1062));
    layer1_outputs(299) <= layer0_outputs(1614);
    layer1_outputs(300) <= not((layer0_outputs(1169)) or (layer0_outputs(1413)));
    layer1_outputs(301) <= layer0_outputs(550);
    layer1_outputs(302) <= not(layer0_outputs(1396));
    layer1_outputs(303) <= (layer0_outputs(1115)) and not (layer0_outputs(1672));
    layer1_outputs(304) <= (layer0_outputs(1572)) or (layer0_outputs(2286));
    layer1_outputs(305) <= (layer0_outputs(2395)) xor (layer0_outputs(2078));
    layer1_outputs(306) <= layer0_outputs(1754);
    layer1_outputs(307) <= layer0_outputs(1403);
    layer1_outputs(308) <= not(layer0_outputs(98));
    layer1_outputs(309) <= '0';
    layer1_outputs(310) <= not(layer0_outputs(1269)) or (layer0_outputs(1432));
    layer1_outputs(311) <= not(layer0_outputs(1373));
    layer1_outputs(312) <= not(layer0_outputs(39)) or (layer0_outputs(1178));
    layer1_outputs(313) <= not(layer0_outputs(966)) or (layer0_outputs(793));
    layer1_outputs(314) <= '0';
    layer1_outputs(315) <= not((layer0_outputs(1275)) and (layer0_outputs(327)));
    layer1_outputs(316) <= not((layer0_outputs(1358)) and (layer0_outputs(2388)));
    layer1_outputs(317) <= not((layer0_outputs(2064)) xor (layer0_outputs(788)));
    layer1_outputs(318) <= (layer0_outputs(2358)) and not (layer0_outputs(825));
    layer1_outputs(319) <= (layer0_outputs(2091)) and not (layer0_outputs(731));
    layer1_outputs(320) <= not(layer0_outputs(1908)) or (layer0_outputs(2073));
    layer1_outputs(321) <= (layer0_outputs(281)) and not (layer0_outputs(1934));
    layer1_outputs(322) <= layer0_outputs(97);
    layer1_outputs(323) <= '0';
    layer1_outputs(324) <= not((layer0_outputs(1393)) and (layer0_outputs(361)));
    layer1_outputs(325) <= not((layer0_outputs(611)) xor (layer0_outputs(1677)));
    layer1_outputs(326) <= not(layer0_outputs(113)) or (layer0_outputs(1779));
    layer1_outputs(327) <= layer0_outputs(2190);
    layer1_outputs(328) <= layer0_outputs(1653);
    layer1_outputs(329) <= layer0_outputs(2369);
    layer1_outputs(330) <= (layer0_outputs(1168)) or (layer0_outputs(1862));
    layer1_outputs(331) <= not(layer0_outputs(589));
    layer1_outputs(332) <= (layer0_outputs(778)) or (layer0_outputs(219));
    layer1_outputs(333) <= '1';
    layer1_outputs(334) <= (layer0_outputs(783)) and not (layer0_outputs(1839));
    layer1_outputs(335) <= not(layer0_outputs(2519));
    layer1_outputs(336) <= not(layer0_outputs(847));
    layer1_outputs(337) <= layer0_outputs(2342);
    layer1_outputs(338) <= not(layer0_outputs(391));
    layer1_outputs(339) <= layer0_outputs(1135);
    layer1_outputs(340) <= not(layer0_outputs(1477)) or (layer0_outputs(2303));
    layer1_outputs(341) <= not((layer0_outputs(880)) and (layer0_outputs(1123)));
    layer1_outputs(342) <= '0';
    layer1_outputs(343) <= layer0_outputs(1988);
    layer1_outputs(344) <= not(layer0_outputs(701));
    layer1_outputs(345) <= not((layer0_outputs(366)) xor (layer0_outputs(2037)));
    layer1_outputs(346) <= not(layer0_outputs(750));
    layer1_outputs(347) <= not((layer0_outputs(1499)) or (layer0_outputs(1044)));
    layer1_outputs(348) <= layer0_outputs(1635);
    layer1_outputs(349) <= not(layer0_outputs(839));
    layer1_outputs(350) <= (layer0_outputs(2003)) and not (layer0_outputs(1762));
    layer1_outputs(351) <= not((layer0_outputs(568)) and (layer0_outputs(1391)));
    layer1_outputs(352) <= not(layer0_outputs(309));
    layer1_outputs(353) <= not((layer0_outputs(2289)) or (layer0_outputs(316)));
    layer1_outputs(354) <= not((layer0_outputs(84)) and (layer0_outputs(2333)));
    layer1_outputs(355) <= not((layer0_outputs(2150)) and (layer0_outputs(1918)));
    layer1_outputs(356) <= not((layer0_outputs(991)) or (layer0_outputs(828)));
    layer1_outputs(357) <= (layer0_outputs(761)) or (layer0_outputs(1839));
    layer1_outputs(358) <= not(layer0_outputs(2288)) or (layer0_outputs(1774));
    layer1_outputs(359) <= not((layer0_outputs(1794)) and (layer0_outputs(58)));
    layer1_outputs(360) <= (layer0_outputs(496)) or (layer0_outputs(931));
    layer1_outputs(361) <= layer0_outputs(679);
    layer1_outputs(362) <= layer0_outputs(1286);
    layer1_outputs(363) <= (layer0_outputs(748)) and not (layer0_outputs(434));
    layer1_outputs(364) <= not(layer0_outputs(759));
    layer1_outputs(365) <= (layer0_outputs(2192)) or (layer0_outputs(1270));
    layer1_outputs(366) <= not(layer0_outputs(323)) or (layer0_outputs(2475));
    layer1_outputs(367) <= layer0_outputs(242);
    layer1_outputs(368) <= (layer0_outputs(2547)) and not (layer0_outputs(1624));
    layer1_outputs(369) <= not(layer0_outputs(2544));
    layer1_outputs(370) <= (layer0_outputs(1829)) and (layer0_outputs(792));
    layer1_outputs(371) <= not(layer0_outputs(1745));
    layer1_outputs(372) <= (layer0_outputs(2181)) and not (layer0_outputs(1461));
    layer1_outputs(373) <= '1';
    layer1_outputs(374) <= (layer0_outputs(2123)) and not (layer0_outputs(687));
    layer1_outputs(375) <= (layer0_outputs(1387)) xor (layer0_outputs(1543));
    layer1_outputs(376) <= not(layer0_outputs(1401));
    layer1_outputs(377) <= not(layer0_outputs(198));
    layer1_outputs(378) <= (layer0_outputs(309)) and (layer0_outputs(1970));
    layer1_outputs(379) <= not(layer0_outputs(1040));
    layer1_outputs(380) <= layer0_outputs(1600);
    layer1_outputs(381) <= not((layer0_outputs(2191)) xor (layer0_outputs(450)));
    layer1_outputs(382) <= (layer0_outputs(1549)) and (layer0_outputs(883));
    layer1_outputs(383) <= not(layer0_outputs(606));
    layer1_outputs(384) <= (layer0_outputs(1714)) and not (layer0_outputs(1461));
    layer1_outputs(385) <= (layer0_outputs(2285)) and not (layer0_outputs(1631));
    layer1_outputs(386) <= not((layer0_outputs(1277)) or (layer0_outputs(31)));
    layer1_outputs(387) <= (layer0_outputs(1641)) and (layer0_outputs(2503));
    layer1_outputs(388) <= layer0_outputs(19);
    layer1_outputs(389) <= not(layer0_outputs(1208));
    layer1_outputs(390) <= (layer0_outputs(413)) and not (layer0_outputs(285));
    layer1_outputs(391) <= layer0_outputs(1864);
    layer1_outputs(392) <= not((layer0_outputs(2296)) and (layer0_outputs(1263)));
    layer1_outputs(393) <= not(layer0_outputs(791));
    layer1_outputs(394) <= '1';
    layer1_outputs(395) <= layer0_outputs(1573);
    layer1_outputs(396) <= not(layer0_outputs(528));
    layer1_outputs(397) <= not(layer0_outputs(1006)) or (layer0_outputs(656));
    layer1_outputs(398) <= layer0_outputs(846);
    layer1_outputs(399) <= not((layer0_outputs(1964)) or (layer0_outputs(511)));
    layer1_outputs(400) <= (layer0_outputs(718)) and not (layer0_outputs(1257));
    layer1_outputs(401) <= not((layer0_outputs(277)) or (layer0_outputs(1735)));
    layer1_outputs(402) <= layer0_outputs(2419);
    layer1_outputs(403) <= '0';
    layer1_outputs(404) <= not((layer0_outputs(1700)) or (layer0_outputs(405)));
    layer1_outputs(405) <= not(layer0_outputs(495));
    layer1_outputs(406) <= not(layer0_outputs(2159));
    layer1_outputs(407) <= (layer0_outputs(2045)) and not (layer0_outputs(256));
    layer1_outputs(408) <= not((layer0_outputs(487)) or (layer0_outputs(318)));
    layer1_outputs(409) <= (layer0_outputs(236)) and not (layer0_outputs(2266));
    layer1_outputs(410) <= not(layer0_outputs(2293));
    layer1_outputs(411) <= not(layer0_outputs(762));
    layer1_outputs(412) <= not((layer0_outputs(1205)) and (layer0_outputs(319)));
    layer1_outputs(413) <= '1';
    layer1_outputs(414) <= '0';
    layer1_outputs(415) <= not(layer0_outputs(110)) or (layer0_outputs(1337));
    layer1_outputs(416) <= (layer0_outputs(1725)) and not (layer0_outputs(1747));
    layer1_outputs(417) <= not(layer0_outputs(127));
    layer1_outputs(418) <= not(layer0_outputs(1596));
    layer1_outputs(419) <= '0';
    layer1_outputs(420) <= (layer0_outputs(1330)) and not (layer0_outputs(2035));
    layer1_outputs(421) <= '1';
    layer1_outputs(422) <= not(layer0_outputs(975));
    layer1_outputs(423) <= '1';
    layer1_outputs(424) <= not(layer0_outputs(307)) or (layer0_outputs(359));
    layer1_outputs(425) <= not(layer0_outputs(1692)) or (layer0_outputs(630));
    layer1_outputs(426) <= not((layer0_outputs(825)) and (layer0_outputs(939)));
    layer1_outputs(427) <= not(layer0_outputs(1900)) or (layer0_outputs(44));
    layer1_outputs(428) <= not(layer0_outputs(2332));
    layer1_outputs(429) <= '0';
    layer1_outputs(430) <= (layer0_outputs(1343)) and not (layer0_outputs(247));
    layer1_outputs(431) <= (layer0_outputs(2122)) and not (layer0_outputs(1633));
    layer1_outputs(432) <= (layer0_outputs(44)) or (layer0_outputs(1552));
    layer1_outputs(433) <= (layer0_outputs(2396)) and (layer0_outputs(1579));
    layer1_outputs(434) <= not(layer0_outputs(515));
    layer1_outputs(435) <= not((layer0_outputs(811)) and (layer0_outputs(2526)));
    layer1_outputs(436) <= (layer0_outputs(1993)) or (layer0_outputs(2368));
    layer1_outputs(437) <= not(layer0_outputs(1145)) or (layer0_outputs(1300));
    layer1_outputs(438) <= (layer0_outputs(17)) and not (layer0_outputs(16));
    layer1_outputs(439) <= layer0_outputs(1581);
    layer1_outputs(440) <= layer0_outputs(522);
    layer1_outputs(441) <= not(layer0_outputs(1350)) or (layer0_outputs(793));
    layer1_outputs(442) <= layer0_outputs(887);
    layer1_outputs(443) <= not((layer0_outputs(1377)) and (layer0_outputs(854)));
    layer1_outputs(444) <= layer0_outputs(1554);
    layer1_outputs(445) <= not(layer0_outputs(2026));
    layer1_outputs(446) <= not(layer0_outputs(114));
    layer1_outputs(447) <= not((layer0_outputs(1604)) and (layer0_outputs(1868)));
    layer1_outputs(448) <= layer0_outputs(1936);
    layer1_outputs(449) <= layer0_outputs(230);
    layer1_outputs(450) <= not(layer0_outputs(2489)) or (layer0_outputs(795));
    layer1_outputs(451) <= layer0_outputs(1133);
    layer1_outputs(452) <= not(layer0_outputs(2363)) or (layer0_outputs(632));
    layer1_outputs(453) <= layer0_outputs(156);
    layer1_outputs(454) <= (layer0_outputs(342)) and not (layer0_outputs(1966));
    layer1_outputs(455) <= not(layer0_outputs(208));
    layer1_outputs(456) <= not((layer0_outputs(247)) and (layer0_outputs(1484)));
    layer1_outputs(457) <= (layer0_outputs(93)) and not (layer0_outputs(1923));
    layer1_outputs(458) <= layer0_outputs(475);
    layer1_outputs(459) <= '0';
    layer1_outputs(460) <= layer0_outputs(9);
    layer1_outputs(461) <= (layer0_outputs(1397)) and not (layer0_outputs(467));
    layer1_outputs(462) <= '1';
    layer1_outputs(463) <= not((layer0_outputs(2197)) xor (layer0_outputs(34)));
    layer1_outputs(464) <= layer0_outputs(2160);
    layer1_outputs(465) <= not(layer0_outputs(836));
    layer1_outputs(466) <= not(layer0_outputs(2270));
    layer1_outputs(467) <= not((layer0_outputs(867)) or (layer0_outputs(2318)));
    layer1_outputs(468) <= not(layer0_outputs(1416));
    layer1_outputs(469) <= (layer0_outputs(78)) or (layer0_outputs(1526));
    layer1_outputs(470) <= layer0_outputs(738);
    layer1_outputs(471) <= (layer0_outputs(1562)) and not (layer0_outputs(401));
    layer1_outputs(472) <= not(layer0_outputs(2223));
    layer1_outputs(473) <= layer0_outputs(699);
    layer1_outputs(474) <= (layer0_outputs(2042)) and not (layer0_outputs(365));
    layer1_outputs(475) <= not((layer0_outputs(2283)) and (layer0_outputs(2)));
    layer1_outputs(476) <= not(layer0_outputs(1866));
    layer1_outputs(477) <= not(layer0_outputs(1353));
    layer1_outputs(478) <= (layer0_outputs(1335)) and not (layer0_outputs(320));
    layer1_outputs(479) <= not(layer0_outputs(837)) or (layer0_outputs(2077));
    layer1_outputs(480) <= (layer0_outputs(2200)) and not (layer0_outputs(849));
    layer1_outputs(481) <= layer0_outputs(677);
    layer1_outputs(482) <= not(layer0_outputs(566));
    layer1_outputs(483) <= '0';
    layer1_outputs(484) <= '1';
    layer1_outputs(485) <= not(layer0_outputs(536)) or (layer0_outputs(1967));
    layer1_outputs(486) <= '1';
    layer1_outputs(487) <= (layer0_outputs(2481)) and not (layer0_outputs(1191));
    layer1_outputs(488) <= (layer0_outputs(2513)) or (layer0_outputs(2335));
    layer1_outputs(489) <= layer0_outputs(1601);
    layer1_outputs(490) <= '1';
    layer1_outputs(491) <= '1';
    layer1_outputs(492) <= layer0_outputs(751);
    layer1_outputs(493) <= not(layer0_outputs(2391));
    layer1_outputs(494) <= not(layer0_outputs(584));
    layer1_outputs(495) <= layer0_outputs(1884);
    layer1_outputs(496) <= layer0_outputs(2291);
    layer1_outputs(497) <= not((layer0_outputs(2550)) and (layer0_outputs(595)));
    layer1_outputs(498) <= (layer0_outputs(629)) or (layer0_outputs(1743));
    layer1_outputs(499) <= layer0_outputs(693);
    layer1_outputs(500) <= layer0_outputs(556);
    layer1_outputs(501) <= '0';
    layer1_outputs(502) <= not((layer0_outputs(479)) and (layer0_outputs(904)));
    layer1_outputs(503) <= (layer0_outputs(1550)) and not (layer0_outputs(1545));
    layer1_outputs(504) <= (layer0_outputs(1810)) and not (layer0_outputs(2348));
    layer1_outputs(505) <= layer0_outputs(389);
    layer1_outputs(506) <= not((layer0_outputs(633)) or (layer0_outputs(2080)));
    layer1_outputs(507) <= not(layer0_outputs(264)) or (layer0_outputs(2136));
    layer1_outputs(508) <= layer0_outputs(1610);
    layer1_outputs(509) <= layer0_outputs(2542);
    layer1_outputs(510) <= not(layer0_outputs(2444)) or (layer0_outputs(2069));
    layer1_outputs(511) <= not(layer0_outputs(2504));
    layer1_outputs(512) <= layer0_outputs(379);
    layer1_outputs(513) <= not(layer0_outputs(2310));
    layer1_outputs(514) <= layer0_outputs(565);
    layer1_outputs(515) <= layer0_outputs(541);
    layer1_outputs(516) <= (layer0_outputs(786)) and not (layer0_outputs(2142));
    layer1_outputs(517) <= not(layer0_outputs(2173));
    layer1_outputs(518) <= not(layer0_outputs(1955));
    layer1_outputs(519) <= not((layer0_outputs(158)) and (layer0_outputs(933)));
    layer1_outputs(520) <= not((layer0_outputs(1190)) or (layer0_outputs(1931)));
    layer1_outputs(521) <= not(layer0_outputs(319)) or (layer0_outputs(160));
    layer1_outputs(522) <= (layer0_outputs(947)) or (layer0_outputs(1246));
    layer1_outputs(523) <= layer0_outputs(1325);
    layer1_outputs(524) <= not(layer0_outputs(607));
    layer1_outputs(525) <= not(layer0_outputs(870));
    layer1_outputs(526) <= not(layer0_outputs(1097)) or (layer0_outputs(2353));
    layer1_outputs(527) <= not(layer0_outputs(2507));
    layer1_outputs(528) <= not(layer0_outputs(217)) or (layer0_outputs(2542));
    layer1_outputs(529) <= not(layer0_outputs(2544)) or (layer0_outputs(1441));
    layer1_outputs(530) <= not(layer0_outputs(1487)) or (layer0_outputs(1768));
    layer1_outputs(531) <= not(layer0_outputs(290)) or (layer0_outputs(887));
    layer1_outputs(532) <= not((layer0_outputs(1543)) or (layer0_outputs(1924)));
    layer1_outputs(533) <= layer0_outputs(1443);
    layer1_outputs(534) <= not((layer0_outputs(91)) and (layer0_outputs(1667)));
    layer1_outputs(535) <= layer0_outputs(1107);
    layer1_outputs(536) <= '1';
    layer1_outputs(537) <= not((layer0_outputs(1812)) and (layer0_outputs(1978)));
    layer1_outputs(538) <= not(layer0_outputs(2479)) or (layer0_outputs(333));
    layer1_outputs(539) <= (layer0_outputs(708)) and (layer0_outputs(233));
    layer1_outputs(540) <= layer0_outputs(502);
    layer1_outputs(541) <= (layer0_outputs(2393)) xor (layer0_outputs(345));
    layer1_outputs(542) <= '1';
    layer1_outputs(543) <= not(layer0_outputs(2002)) or (layer0_outputs(729));
    layer1_outputs(544) <= (layer0_outputs(2406)) and not (layer0_outputs(1069));
    layer1_outputs(545) <= not(layer0_outputs(2437)) or (layer0_outputs(978));
    layer1_outputs(546) <= (layer0_outputs(1235)) and not (layer0_outputs(2136));
    layer1_outputs(547) <= not(layer0_outputs(861));
    layer1_outputs(548) <= not(layer0_outputs(1476));
    layer1_outputs(549) <= not((layer0_outputs(2232)) and (layer0_outputs(2053)));
    layer1_outputs(550) <= (layer0_outputs(2415)) and not (layer0_outputs(1523));
    layer1_outputs(551) <= (layer0_outputs(1583)) and (layer0_outputs(1352));
    layer1_outputs(552) <= (layer0_outputs(669)) or (layer0_outputs(1897));
    layer1_outputs(553) <= (layer0_outputs(149)) or (layer0_outputs(510));
    layer1_outputs(554) <= '1';
    layer1_outputs(555) <= layer0_outputs(45);
    layer1_outputs(556) <= not(layer0_outputs(1045));
    layer1_outputs(557) <= (layer0_outputs(1282)) or (layer0_outputs(613));
    layer1_outputs(558) <= not(layer0_outputs(2285)) or (layer0_outputs(1502));
    layer1_outputs(559) <= '0';
    layer1_outputs(560) <= layer0_outputs(1751);
    layer1_outputs(561) <= not((layer0_outputs(899)) xor (layer0_outputs(575)));
    layer1_outputs(562) <= not((layer0_outputs(1574)) and (layer0_outputs(151)));
    layer1_outputs(563) <= not((layer0_outputs(28)) xor (layer0_outputs(1395)));
    layer1_outputs(564) <= (layer0_outputs(1241)) and (layer0_outputs(7));
    layer1_outputs(565) <= not(layer0_outputs(1483));
    layer1_outputs(566) <= (layer0_outputs(1317)) and (layer0_outputs(125));
    layer1_outputs(567) <= not((layer0_outputs(88)) and (layer0_outputs(2179)));
    layer1_outputs(568) <= layer0_outputs(1470);
    layer1_outputs(569) <= layer0_outputs(1015);
    layer1_outputs(570) <= not(layer0_outputs(99)) or (layer0_outputs(2252));
    layer1_outputs(571) <= not((layer0_outputs(2453)) and (layer0_outputs(1090)));
    layer1_outputs(572) <= not(layer0_outputs(1789)) or (layer0_outputs(1835));
    layer1_outputs(573) <= not((layer0_outputs(38)) or (layer0_outputs(1567)));
    layer1_outputs(574) <= layer0_outputs(765);
    layer1_outputs(575) <= not(layer0_outputs(1032)) or (layer0_outputs(772));
    layer1_outputs(576) <= layer0_outputs(1791);
    layer1_outputs(577) <= not(layer0_outputs(2020)) or (layer0_outputs(1650));
    layer1_outputs(578) <= not(layer0_outputs(746)) or (layer0_outputs(2456));
    layer1_outputs(579) <= not((layer0_outputs(2232)) and (layer0_outputs(841)));
    layer1_outputs(580) <= not(layer0_outputs(1002)) or (layer0_outputs(344));
    layer1_outputs(581) <= (layer0_outputs(287)) and not (layer0_outputs(277));
    layer1_outputs(582) <= (layer0_outputs(2148)) or (layer0_outputs(386));
    layer1_outputs(583) <= layer0_outputs(2182);
    layer1_outputs(584) <= '1';
    layer1_outputs(585) <= (layer0_outputs(780)) and (layer0_outputs(36));
    layer1_outputs(586) <= (layer0_outputs(961)) and (layer0_outputs(2320));
    layer1_outputs(587) <= not(layer0_outputs(1819)) or (layer0_outputs(1112));
    layer1_outputs(588) <= not(layer0_outputs(1350));
    layer1_outputs(589) <= '1';
    layer1_outputs(590) <= (layer0_outputs(349)) and not (layer0_outputs(929));
    layer1_outputs(591) <= layer0_outputs(669);
    layer1_outputs(592) <= '0';
    layer1_outputs(593) <= not(layer0_outputs(1025));
    layer1_outputs(594) <= (layer0_outputs(1504)) and (layer0_outputs(2023));
    layer1_outputs(595) <= layer0_outputs(808);
    layer1_outputs(596) <= layer0_outputs(2114);
    layer1_outputs(597) <= layer0_outputs(262);
    layer1_outputs(598) <= not(layer0_outputs(741)) or (layer0_outputs(2153));
    layer1_outputs(599) <= not(layer0_outputs(1063));
    layer1_outputs(600) <= not(layer0_outputs(443));
    layer1_outputs(601) <= not(layer0_outputs(1661)) or (layer0_outputs(234));
    layer1_outputs(602) <= (layer0_outputs(53)) or (layer0_outputs(853));
    layer1_outputs(603) <= (layer0_outputs(2317)) and not (layer0_outputs(1863));
    layer1_outputs(604) <= layer0_outputs(1843);
    layer1_outputs(605) <= not((layer0_outputs(1884)) or (layer0_outputs(1991)));
    layer1_outputs(606) <= not((layer0_outputs(66)) and (layer0_outputs(451)));
    layer1_outputs(607) <= layer0_outputs(733);
    layer1_outputs(608) <= '0';
    layer1_outputs(609) <= layer0_outputs(191);
    layer1_outputs(610) <= not((layer0_outputs(2128)) and (layer0_outputs(2248)));
    layer1_outputs(611) <= not(layer0_outputs(1468));
    layer1_outputs(612) <= (layer0_outputs(17)) and (layer0_outputs(1514));
    layer1_outputs(613) <= (layer0_outputs(308)) or (layer0_outputs(1946));
    layer1_outputs(614) <= not(layer0_outputs(15));
    layer1_outputs(615) <= not(layer0_outputs(1449));
    layer1_outputs(616) <= (layer0_outputs(2384)) and not (layer0_outputs(1293));
    layer1_outputs(617) <= '0';
    layer1_outputs(618) <= layer0_outputs(2549);
    layer1_outputs(619) <= (layer0_outputs(888)) and (layer0_outputs(2138));
    layer1_outputs(620) <= not(layer0_outputs(420)) or (layer0_outputs(641));
    layer1_outputs(621) <= not((layer0_outputs(1749)) and (layer0_outputs(505)));
    layer1_outputs(622) <= not((layer0_outputs(1472)) or (layer0_outputs(999)));
    layer1_outputs(623) <= not(layer0_outputs(692));
    layer1_outputs(624) <= (layer0_outputs(2239)) and (layer0_outputs(2141));
    layer1_outputs(625) <= not(layer0_outputs(912));
    layer1_outputs(626) <= not(layer0_outputs(619)) or (layer0_outputs(2222));
    layer1_outputs(627) <= not(layer0_outputs(727));
    layer1_outputs(628) <= not(layer0_outputs(1179));
    layer1_outputs(629) <= not(layer0_outputs(274));
    layer1_outputs(630) <= (layer0_outputs(372)) or (layer0_outputs(2029));
    layer1_outputs(631) <= not(layer0_outputs(2234));
    layer1_outputs(632) <= not(layer0_outputs(715));
    layer1_outputs(633) <= layer0_outputs(774);
    layer1_outputs(634) <= layer0_outputs(980);
    layer1_outputs(635) <= '0';
    layer1_outputs(636) <= (layer0_outputs(1400)) and not (layer0_outputs(416));
    layer1_outputs(637) <= '0';
    layer1_outputs(638) <= not(layer0_outputs(711));
    layer1_outputs(639) <= layer0_outputs(949);
    layer1_outputs(640) <= (layer0_outputs(1148)) and not (layer0_outputs(1965));
    layer1_outputs(641) <= layer0_outputs(235);
    layer1_outputs(642) <= not((layer0_outputs(146)) and (layer0_outputs(1906)));
    layer1_outputs(643) <= not(layer0_outputs(1856));
    layer1_outputs(644) <= not(layer0_outputs(503));
    layer1_outputs(645) <= layer0_outputs(129);
    layer1_outputs(646) <= (layer0_outputs(1728)) or (layer0_outputs(1913));
    layer1_outputs(647) <= not(layer0_outputs(1505));
    layer1_outputs(648) <= not(layer0_outputs(1942));
    layer1_outputs(649) <= (layer0_outputs(2456)) or (layer0_outputs(893));
    layer1_outputs(650) <= (layer0_outputs(1627)) and not (layer0_outputs(712));
    layer1_outputs(651) <= not(layer0_outputs(2000)) or (layer0_outputs(1774));
    layer1_outputs(652) <= (layer0_outputs(1110)) or (layer0_outputs(288));
    layer1_outputs(653) <= not(layer0_outputs(1176)) or (layer0_outputs(527));
    layer1_outputs(654) <= (layer0_outputs(87)) and (layer0_outputs(311));
    layer1_outputs(655) <= not((layer0_outputs(1507)) and (layer0_outputs(567)));
    layer1_outputs(656) <= layer0_outputs(914);
    layer1_outputs(657) <= not((layer0_outputs(1790)) or (layer0_outputs(1030)));
    layer1_outputs(658) <= (layer0_outputs(1920)) and not (layer0_outputs(2172));
    layer1_outputs(659) <= not(layer0_outputs(449)) or (layer0_outputs(2246));
    layer1_outputs(660) <= not(layer0_outputs(1271));
    layer1_outputs(661) <= not((layer0_outputs(1415)) and (layer0_outputs(913)));
    layer1_outputs(662) <= (layer0_outputs(862)) and (layer0_outputs(927));
    layer1_outputs(663) <= (layer0_outputs(1320)) and not (layer0_outputs(190));
    layer1_outputs(664) <= not((layer0_outputs(176)) and (layer0_outputs(2085)));
    layer1_outputs(665) <= (layer0_outputs(1187)) and (layer0_outputs(2474));
    layer1_outputs(666) <= layer0_outputs(726);
    layer1_outputs(667) <= (layer0_outputs(1157)) and not (layer0_outputs(843));
    layer1_outputs(668) <= layer0_outputs(2313);
    layer1_outputs(669) <= not((layer0_outputs(1457)) or (layer0_outputs(849)));
    layer1_outputs(670) <= not(layer0_outputs(2436)) or (layer0_outputs(500));
    layer1_outputs(671) <= not(layer0_outputs(2537));
    layer1_outputs(672) <= layer0_outputs(1660);
    layer1_outputs(673) <= layer0_outputs(2023);
    layer1_outputs(674) <= not((layer0_outputs(2414)) and (layer0_outputs(2146)));
    layer1_outputs(675) <= layer0_outputs(224);
    layer1_outputs(676) <= (layer0_outputs(827)) or (layer0_outputs(58));
    layer1_outputs(677) <= not(layer0_outputs(2145));
    layer1_outputs(678) <= not(layer0_outputs(911)) or (layer0_outputs(1473));
    layer1_outputs(679) <= not(layer0_outputs(2423));
    layer1_outputs(680) <= not(layer0_outputs(459));
    layer1_outputs(681) <= not(layer0_outputs(1068)) or (layer0_outputs(489));
    layer1_outputs(682) <= not((layer0_outputs(1907)) or (layer0_outputs(2226)));
    layer1_outputs(683) <= (layer0_outputs(2479)) or (layer0_outputs(1880));
    layer1_outputs(684) <= layer0_outputs(966);
    layer1_outputs(685) <= layer0_outputs(392);
    layer1_outputs(686) <= (layer0_outputs(1823)) and not (layer0_outputs(51));
    layer1_outputs(687) <= not(layer0_outputs(1236));
    layer1_outputs(688) <= layer0_outputs(931);
    layer1_outputs(689) <= (layer0_outputs(942)) and not (layer0_outputs(826));
    layer1_outputs(690) <= layer0_outputs(2506);
    layer1_outputs(691) <= (layer0_outputs(1082)) and not (layer0_outputs(1444));
    layer1_outputs(692) <= (layer0_outputs(636)) and not (layer0_outputs(891));
    layer1_outputs(693) <= layer0_outputs(25);
    layer1_outputs(694) <= '1';
    layer1_outputs(695) <= not(layer0_outputs(2368));
    layer1_outputs(696) <= not(layer0_outputs(1298));
    layer1_outputs(697) <= not(layer0_outputs(1486));
    layer1_outputs(698) <= (layer0_outputs(2477)) and (layer0_outputs(1679));
    layer1_outputs(699) <= layer0_outputs(185);
    layer1_outputs(700) <= not((layer0_outputs(1809)) xor (layer0_outputs(10)));
    layer1_outputs(701) <= not((layer0_outputs(349)) xor (layer0_outputs(1089)));
    layer1_outputs(702) <= not((layer0_outputs(1962)) and (layer0_outputs(2084)));
    layer1_outputs(703) <= not(layer0_outputs(2151));
    layer1_outputs(704) <= '0';
    layer1_outputs(705) <= layer0_outputs(1877);
    layer1_outputs(706) <= '0';
    layer1_outputs(707) <= not(layer0_outputs(1162));
    layer1_outputs(708) <= not((layer0_outputs(616)) and (layer0_outputs(2431)));
    layer1_outputs(709) <= (layer0_outputs(2458)) xor (layer0_outputs(1608));
    layer1_outputs(710) <= not(layer0_outputs(431)) or (layer0_outputs(606));
    layer1_outputs(711) <= not(layer0_outputs(806));
    layer1_outputs(712) <= not((layer0_outputs(480)) xor (layer0_outputs(278)));
    layer1_outputs(713) <= not(layer0_outputs(432)) or (layer0_outputs(423));
    layer1_outputs(714) <= layer0_outputs(1489);
    layer1_outputs(715) <= (layer0_outputs(1411)) and (layer0_outputs(198));
    layer1_outputs(716) <= '1';
    layer1_outputs(717) <= not((layer0_outputs(74)) or (layer0_outputs(2417)));
    layer1_outputs(718) <= not(layer0_outputs(2518));
    layer1_outputs(719) <= not(layer0_outputs(1103));
    layer1_outputs(720) <= layer0_outputs(2040);
    layer1_outputs(721) <= not((layer0_outputs(661)) or (layer0_outputs(1901)));
    layer1_outputs(722) <= not(layer0_outputs(1360));
    layer1_outputs(723) <= layer0_outputs(1777);
    layer1_outputs(724) <= not(layer0_outputs(724));
    layer1_outputs(725) <= layer0_outputs(1313);
    layer1_outputs(726) <= not((layer0_outputs(1689)) or (layer0_outputs(1302)));
    layer1_outputs(727) <= not((layer0_outputs(1521)) and (layer0_outputs(1955)));
    layer1_outputs(728) <= (layer0_outputs(923)) and not (layer0_outputs(2319));
    layer1_outputs(729) <= layer0_outputs(440);
    layer1_outputs(730) <= (layer0_outputs(1703)) or (layer0_outputs(950));
    layer1_outputs(731) <= not(layer0_outputs(2420));
    layer1_outputs(732) <= (layer0_outputs(644)) and (layer0_outputs(1722));
    layer1_outputs(733) <= not((layer0_outputs(637)) and (layer0_outputs(2410)));
    layer1_outputs(734) <= not((layer0_outputs(964)) or (layer0_outputs(2107)));
    layer1_outputs(735) <= (layer0_outputs(1019)) and not (layer0_outputs(2340));
    layer1_outputs(736) <= (layer0_outputs(373)) and not (layer0_outputs(2195));
    layer1_outputs(737) <= layer0_outputs(1084);
    layer1_outputs(738) <= (layer0_outputs(1673)) and not (layer0_outputs(2245));
    layer1_outputs(739) <= not(layer0_outputs(1024));
    layer1_outputs(740) <= not(layer0_outputs(1953));
    layer1_outputs(741) <= not((layer0_outputs(2405)) and (layer0_outputs(2288)));
    layer1_outputs(742) <= (layer0_outputs(2466)) and not (layer0_outputs(1831));
    layer1_outputs(743) <= not(layer0_outputs(101));
    layer1_outputs(744) <= (layer0_outputs(2016)) and (layer0_outputs(2187));
    layer1_outputs(745) <= not(layer0_outputs(1893)) or (layer0_outputs(1125));
    layer1_outputs(746) <= (layer0_outputs(2272)) and not (layer0_outputs(351));
    layer1_outputs(747) <= layer0_outputs(1658);
    layer1_outputs(748) <= layer0_outputs(2082);
    layer1_outputs(749) <= layer0_outputs(1338);
    layer1_outputs(750) <= not(layer0_outputs(174));
    layer1_outputs(751) <= (layer0_outputs(1032)) and (layer0_outputs(813));
    layer1_outputs(752) <= not(layer0_outputs(2513));
    layer1_outputs(753) <= layer0_outputs(1199);
    layer1_outputs(754) <= not(layer0_outputs(1591));
    layer1_outputs(755) <= '1';
    layer1_outputs(756) <= not(layer0_outputs(1482)) or (layer0_outputs(1440));
    layer1_outputs(757) <= not(layer0_outputs(903));
    layer1_outputs(758) <= layer0_outputs(2032);
    layer1_outputs(759) <= layer0_outputs(990);
    layer1_outputs(760) <= not((layer0_outputs(1720)) or (layer0_outputs(2184)));
    layer1_outputs(761) <= (layer0_outputs(1188)) and not (layer0_outputs(795));
    layer1_outputs(762) <= not(layer0_outputs(1886)) or (layer0_outputs(1753));
    layer1_outputs(763) <= not(layer0_outputs(1115));
    layer1_outputs(764) <= not(layer0_outputs(2216)) or (layer0_outputs(1196));
    layer1_outputs(765) <= layer0_outputs(1386);
    layer1_outputs(766) <= not((layer0_outputs(1087)) or (layer0_outputs(819)));
    layer1_outputs(767) <= not(layer0_outputs(985));
    layer1_outputs(768) <= (layer0_outputs(919)) and not (layer0_outputs(1060));
    layer1_outputs(769) <= (layer0_outputs(2089)) and (layer0_outputs(275));
    layer1_outputs(770) <= layer0_outputs(872);
    layer1_outputs(771) <= layer0_outputs(1443);
    layer1_outputs(772) <= (layer0_outputs(226)) or (layer0_outputs(266));
    layer1_outputs(773) <= not(layer0_outputs(2046));
    layer1_outputs(774) <= not(layer0_outputs(1976)) or (layer0_outputs(2139));
    layer1_outputs(775) <= '1';
    layer1_outputs(776) <= not(layer0_outputs(1848)) or (layer0_outputs(412));
    layer1_outputs(777) <= not(layer0_outputs(1938)) or (layer0_outputs(1781));
    layer1_outputs(778) <= layer0_outputs(851);
    layer1_outputs(779) <= not(layer0_outputs(240));
    layer1_outputs(780) <= (layer0_outputs(350)) and not (layer0_outputs(908));
    layer1_outputs(781) <= '0';
    layer1_outputs(782) <= (layer0_outputs(1431)) and (layer0_outputs(2101));
    layer1_outputs(783) <= (layer0_outputs(1138)) and not (layer0_outputs(1290));
    layer1_outputs(784) <= (layer0_outputs(1093)) and not (layer0_outputs(164));
    layer1_outputs(785) <= (layer0_outputs(1586)) xor (layer0_outputs(2519));
    layer1_outputs(786) <= (layer0_outputs(725)) and not (layer0_outputs(147));
    layer1_outputs(787) <= layer0_outputs(2375);
    layer1_outputs(788) <= not((layer0_outputs(1688)) and (layer0_outputs(39)));
    layer1_outputs(789) <= not(layer0_outputs(1822));
    layer1_outputs(790) <= layer0_outputs(1848);
    layer1_outputs(791) <= layer0_outputs(909);
    layer1_outputs(792) <= not(layer0_outputs(1128)) or (layer0_outputs(2027));
    layer1_outputs(793) <= layer0_outputs(94);
    layer1_outputs(794) <= not(layer0_outputs(707)) or (layer0_outputs(185));
    layer1_outputs(795) <= not((layer0_outputs(1691)) xor (layer0_outputs(1211)));
    layer1_outputs(796) <= not((layer0_outputs(1717)) and (layer0_outputs(2487)));
    layer1_outputs(797) <= (layer0_outputs(1771)) and not (layer0_outputs(2241));
    layer1_outputs(798) <= (layer0_outputs(1206)) and (layer0_outputs(1888));
    layer1_outputs(799) <= (layer0_outputs(1261)) and not (layer0_outputs(576));
    layer1_outputs(800) <= (layer0_outputs(1244)) and (layer0_outputs(2344));
    layer1_outputs(801) <= '0';
    layer1_outputs(802) <= (layer0_outputs(1816)) and (layer0_outputs(1525));
    layer1_outputs(803) <= not(layer0_outputs(2124)) or (layer0_outputs(2546));
    layer1_outputs(804) <= not(layer0_outputs(2385)) or (layer0_outputs(768));
    layer1_outputs(805) <= (layer0_outputs(816)) and not (layer0_outputs(1670));
    layer1_outputs(806) <= not(layer0_outputs(326)) or (layer0_outputs(1792));
    layer1_outputs(807) <= layer0_outputs(188);
    layer1_outputs(808) <= layer0_outputs(2335);
    layer1_outputs(809) <= '0';
    layer1_outputs(810) <= not(layer0_outputs(131));
    layer1_outputs(811) <= '0';
    layer1_outputs(812) <= (layer0_outputs(2215)) and not (layer0_outputs(1745));
    layer1_outputs(813) <= layer0_outputs(2256);
    layer1_outputs(814) <= (layer0_outputs(1231)) and not (layer0_outputs(1436));
    layer1_outputs(815) <= '1';
    layer1_outputs(816) <= (layer0_outputs(1628)) and not (layer0_outputs(1866));
    layer1_outputs(817) <= not(layer0_outputs(438)) or (layer0_outputs(2450));
    layer1_outputs(818) <= (layer0_outputs(1896)) and not (layer0_outputs(2244));
    layer1_outputs(819) <= (layer0_outputs(1856)) or (layer0_outputs(398));
    layer1_outputs(820) <= '1';
    layer1_outputs(821) <= not(layer0_outputs(905)) or (layer0_outputs(1599));
    layer1_outputs(822) <= not(layer0_outputs(499)) or (layer0_outputs(1638));
    layer1_outputs(823) <= not((layer0_outputs(1849)) and (layer0_outputs(1099)));
    layer1_outputs(824) <= not(layer0_outputs(1036));
    layer1_outputs(825) <= (layer0_outputs(1374)) and not (layer0_outputs(573));
    layer1_outputs(826) <= not(layer0_outputs(1092)) or (layer0_outputs(1612));
    layer1_outputs(827) <= '1';
    layer1_outputs(828) <= (layer0_outputs(1859)) or (layer0_outputs(2164));
    layer1_outputs(829) <= layer0_outputs(2433);
    layer1_outputs(830) <= not(layer0_outputs(2118)) or (layer0_outputs(1974));
    layer1_outputs(831) <= '0';
    layer1_outputs(832) <= '1';
    layer1_outputs(833) <= (layer0_outputs(1405)) or (layer0_outputs(527));
    layer1_outputs(834) <= not((layer0_outputs(476)) or (layer0_outputs(807)));
    layer1_outputs(835) <= not((layer0_outputs(1613)) or (layer0_outputs(1243)));
    layer1_outputs(836) <= not(layer0_outputs(1351)) or (layer0_outputs(2159));
    layer1_outputs(837) <= not(layer0_outputs(1100));
    layer1_outputs(838) <= layer0_outputs(860);
    layer1_outputs(839) <= not(layer0_outputs(2447)) or (layer0_outputs(1117));
    layer1_outputs(840) <= not((layer0_outputs(1948)) xor (layer0_outputs(773)));
    layer1_outputs(841) <= layer0_outputs(2348);
    layer1_outputs(842) <= (layer0_outputs(1983)) and not (layer0_outputs(801));
    layer1_outputs(843) <= not(layer0_outputs(2242)) or (layer0_outputs(405));
    layer1_outputs(844) <= '0';
    layer1_outputs(845) <= not((layer0_outputs(2282)) or (layer0_outputs(1657)));
    layer1_outputs(846) <= layer0_outputs(933);
    layer1_outputs(847) <= not(layer0_outputs(2220)) or (layer0_outputs(1123));
    layer1_outputs(848) <= not((layer0_outputs(1873)) and (layer0_outputs(178)));
    layer1_outputs(849) <= not(layer0_outputs(1764)) or (layer0_outputs(204));
    layer1_outputs(850) <= not(layer0_outputs(2477));
    layer1_outputs(851) <= '0';
    layer1_outputs(852) <= not(layer0_outputs(1592)) or (layer0_outputs(658));
    layer1_outputs(853) <= (layer0_outputs(212)) or (layer0_outputs(1593));
    layer1_outputs(854) <= not(layer0_outputs(96));
    layer1_outputs(855) <= not((layer0_outputs(776)) and (layer0_outputs(1968)));
    layer1_outputs(856) <= not(layer0_outputs(162));
    layer1_outputs(857) <= not(layer0_outputs(175)) or (layer0_outputs(2329));
    layer1_outputs(858) <= layer0_outputs(562);
    layer1_outputs(859) <= layer0_outputs(956);
    layer1_outputs(860) <= not((layer0_outputs(2157)) xor (layer0_outputs(1254)));
    layer1_outputs(861) <= (layer0_outputs(2191)) and not (layer0_outputs(1756));
    layer1_outputs(862) <= not((layer0_outputs(1039)) and (layer0_outputs(1910)));
    layer1_outputs(863) <= not(layer0_outputs(1563));
    layer1_outputs(864) <= layer0_outputs(876);
    layer1_outputs(865) <= not(layer0_outputs(334));
    layer1_outputs(866) <= layer0_outputs(1878);
    layer1_outputs(867) <= not(layer0_outputs(1588));
    layer1_outputs(868) <= not(layer0_outputs(2207));
    layer1_outputs(869) <= not((layer0_outputs(2126)) or (layer0_outputs(299)));
    layer1_outputs(870) <= not(layer0_outputs(710));
    layer1_outputs(871) <= layer0_outputs(1578);
    layer1_outputs(872) <= (layer0_outputs(1401)) and not (layer0_outputs(94));
    layer1_outputs(873) <= layer0_outputs(881);
    layer1_outputs(874) <= layer0_outputs(1310);
    layer1_outputs(875) <= not((layer0_outputs(2024)) and (layer0_outputs(1463)));
    layer1_outputs(876) <= not((layer0_outputs(1110)) or (layer0_outputs(357)));
    layer1_outputs(877) <= (layer0_outputs(675)) xor (layer0_outputs(1493));
    layer1_outputs(878) <= (layer0_outputs(999)) and not (layer0_outputs(2179));
    layer1_outputs(879) <= not((layer0_outputs(395)) or (layer0_outputs(1192)));
    layer1_outputs(880) <= (layer0_outputs(29)) and not (layer0_outputs(1904));
    layer1_outputs(881) <= (layer0_outputs(280)) and not (layer0_outputs(704));
    layer1_outputs(882) <= not(layer0_outputs(1172)) or (layer0_outputs(83));
    layer1_outputs(883) <= not(layer0_outputs(1034));
    layer1_outputs(884) <= (layer0_outputs(243)) and not (layer0_outputs(829));
    layer1_outputs(885) <= layer0_outputs(1804);
    layer1_outputs(886) <= not(layer0_outputs(2377));
    layer1_outputs(887) <= layer0_outputs(1913);
    layer1_outputs(888) <= not(layer0_outputs(2106));
    layer1_outputs(889) <= layer0_outputs(1213);
    layer1_outputs(890) <= not(layer0_outputs(367)) or (layer0_outputs(1512));
    layer1_outputs(891) <= not(layer0_outputs(120));
    layer1_outputs(892) <= layer0_outputs(2113);
    layer1_outputs(893) <= '0';
    layer1_outputs(894) <= not(layer0_outputs(2236)) or (layer0_outputs(1208));
    layer1_outputs(895) <= (layer0_outputs(2271)) and not (layer0_outputs(453));
    layer1_outputs(896) <= layer0_outputs(1334);
    layer1_outputs(897) <= (layer0_outputs(1450)) and not (layer0_outputs(470));
    layer1_outputs(898) <= not(layer0_outputs(1786)) or (layer0_outputs(1990));
    layer1_outputs(899) <= not(layer0_outputs(1607));
    layer1_outputs(900) <= (layer0_outputs(2279)) xor (layer0_outputs(2240));
    layer1_outputs(901) <= '0';
    layer1_outputs(902) <= not((layer0_outputs(2282)) xor (layer0_outputs(428)));
    layer1_outputs(903) <= layer0_outputs(2469);
    layer1_outputs(904) <= '1';
    layer1_outputs(905) <= (layer0_outputs(1103)) or (layer0_outputs(146));
    layer1_outputs(906) <= not(layer0_outputs(1737));
    layer1_outputs(907) <= not(layer0_outputs(2049));
    layer1_outputs(908) <= layer0_outputs(1980);
    layer1_outputs(909) <= '0';
    layer1_outputs(910) <= not(layer0_outputs(40));
    layer1_outputs(911) <= (layer0_outputs(448)) and not (layer0_outputs(61));
    layer1_outputs(912) <= not(layer0_outputs(993));
    layer1_outputs(913) <= (layer0_outputs(1154)) and not (layer0_outputs(1874));
    layer1_outputs(914) <= not((layer0_outputs(1151)) or (layer0_outputs(2488)));
    layer1_outputs(915) <= '0';
    layer1_outputs(916) <= not(layer0_outputs(1678));
    layer1_outputs(917) <= not(layer0_outputs(782)) or (layer0_outputs(37));
    layer1_outputs(918) <= (layer0_outputs(1177)) and (layer0_outputs(2293));
    layer1_outputs(919) <= not(layer0_outputs(2226));
    layer1_outputs(920) <= not(layer0_outputs(1191)) or (layer0_outputs(521));
    layer1_outputs(921) <= '0';
    layer1_outputs(922) <= not((layer0_outputs(876)) or (layer0_outputs(1462)));
    layer1_outputs(923) <= not(layer0_outputs(273));
    layer1_outputs(924) <= (layer0_outputs(1812)) and not (layer0_outputs(2349));
    layer1_outputs(925) <= not((layer0_outputs(1733)) or (layer0_outputs(1682)));
    layer1_outputs(926) <= layer0_outputs(410);
    layer1_outputs(927) <= layer0_outputs(138);
    layer1_outputs(928) <= (layer0_outputs(2238)) and not (layer0_outputs(1278));
    layer1_outputs(929) <= (layer0_outputs(1722)) and not (layer0_outputs(2208));
    layer1_outputs(930) <= layer0_outputs(1734);
    layer1_outputs(931) <= layer0_outputs(2052);
    layer1_outputs(932) <= '1';
    layer1_outputs(933) <= not(layer0_outputs(2043));
    layer1_outputs(934) <= (layer0_outputs(1276)) and (layer0_outputs(359));
    layer1_outputs(935) <= layer0_outputs(2204);
    layer1_outputs(936) <= not(layer0_outputs(1051));
    layer1_outputs(937) <= not((layer0_outputs(1185)) and (layer0_outputs(1040)));
    layer1_outputs(938) <= (layer0_outputs(525)) and not (layer0_outputs(149));
    layer1_outputs(939) <= (layer0_outputs(1328)) and not (layer0_outputs(1153));
    layer1_outputs(940) <= (layer0_outputs(1697)) or (layer0_outputs(1395));
    layer1_outputs(941) <= (layer0_outputs(1166)) and (layer0_outputs(1528));
    layer1_outputs(942) <= not(layer0_outputs(1383));
    layer1_outputs(943) <= not(layer0_outputs(2276));
    layer1_outputs(944) <= not(layer0_outputs(69));
    layer1_outputs(945) <= layer0_outputs(1801);
    layer1_outputs(946) <= (layer0_outputs(250)) and (layer0_outputs(1761));
    layer1_outputs(947) <= (layer0_outputs(1055)) and not (layer0_outputs(418));
    layer1_outputs(948) <= not((layer0_outputs(1365)) or (layer0_outputs(2532)));
    layer1_outputs(949) <= (layer0_outputs(713)) or (layer0_outputs(2199));
    layer1_outputs(950) <= '1';
    layer1_outputs(951) <= not(layer0_outputs(2066)) or (layer0_outputs(963));
    layer1_outputs(952) <= not(layer0_outputs(1763));
    layer1_outputs(953) <= not(layer0_outputs(2527));
    layer1_outputs(954) <= not((layer0_outputs(491)) or (layer0_outputs(2435)));
    layer1_outputs(955) <= layer0_outputs(1337);
    layer1_outputs(956) <= '0';
    layer1_outputs(957) <= (layer0_outputs(1726)) and not (layer0_outputs(29));
    layer1_outputs(958) <= not(layer0_outputs(951)) or (layer0_outputs(1038));
    layer1_outputs(959) <= (layer0_outputs(2515)) and (layer0_outputs(1342));
    layer1_outputs(960) <= not((layer0_outputs(516)) or (layer0_outputs(2511)));
    layer1_outputs(961) <= (layer0_outputs(2413)) and not (layer0_outputs(157));
    layer1_outputs(962) <= layer0_outputs(979);
    layer1_outputs(963) <= (layer0_outputs(1953)) or (layer0_outputs(978));
    layer1_outputs(964) <= (layer0_outputs(1102)) and not (layer0_outputs(1819));
    layer1_outputs(965) <= not(layer0_outputs(1392));
    layer1_outputs(966) <= (layer0_outputs(200)) and not (layer0_outputs(737));
    layer1_outputs(967) <= '1';
    layer1_outputs(968) <= '0';
    layer1_outputs(969) <= layer0_outputs(918);
    layer1_outputs(970) <= (layer0_outputs(1993)) or (layer0_outputs(2506));
    layer1_outputs(971) <= not(layer0_outputs(1155));
    layer1_outputs(972) <= not((layer0_outputs(2424)) or (layer0_outputs(514)));
    layer1_outputs(973) <= layer0_outputs(502);
    layer1_outputs(974) <= not(layer0_outputs(856));
    layer1_outputs(975) <= layer0_outputs(1425);
    layer1_outputs(976) <= '1';
    layer1_outputs(977) <= not(layer0_outputs(234)) or (layer0_outputs(1049));
    layer1_outputs(978) <= not(layer0_outputs(2168)) or (layer0_outputs(2439));
    layer1_outputs(979) <= not((layer0_outputs(2077)) or (layer0_outputs(1266)));
    layer1_outputs(980) <= (layer0_outputs(642)) and (layer0_outputs(597));
    layer1_outputs(981) <= (layer0_outputs(1956)) and not (layer0_outputs(2331));
    layer1_outputs(982) <= not(layer0_outputs(934));
    layer1_outputs(983) <= (layer0_outputs(767)) and not (layer0_outputs(1082));
    layer1_outputs(984) <= not(layer0_outputs(1748)) or (layer0_outputs(1917));
    layer1_outputs(985) <= (layer0_outputs(1893)) and (layer0_outputs(2307));
    layer1_outputs(986) <= not(layer0_outputs(2171));
    layer1_outputs(987) <= not((layer0_outputs(1491)) xor (layer0_outputs(19)));
    layer1_outputs(988) <= not((layer0_outputs(612)) xor (layer0_outputs(1218)));
    layer1_outputs(989) <= layer0_outputs(2401);
    layer1_outputs(990) <= not(layer0_outputs(1462)) or (layer0_outputs(251));
    layer1_outputs(991) <= layer0_outputs(896);
    layer1_outputs(992) <= not(layer0_outputs(1313));
    layer1_outputs(993) <= not(layer0_outputs(1270));
    layer1_outputs(994) <= not(layer0_outputs(1683));
    layer1_outputs(995) <= not(layer0_outputs(709));
    layer1_outputs(996) <= (layer0_outputs(1345)) and not (layer0_outputs(1021));
    layer1_outputs(997) <= (layer0_outputs(1881)) or (layer0_outputs(805));
    layer1_outputs(998) <= (layer0_outputs(1811)) and not (layer0_outputs(1011));
    layer1_outputs(999) <= not(layer0_outputs(1198));
    layer1_outputs(1000) <= not(layer0_outputs(173));
    layer1_outputs(1001) <= (layer0_outputs(855)) or (layer0_outputs(1244));
    layer1_outputs(1002) <= (layer0_outputs(141)) and (layer0_outputs(2092));
    layer1_outputs(1003) <= not(layer0_outputs(684));
    layer1_outputs(1004) <= layer0_outputs(353);
    layer1_outputs(1005) <= not((layer0_outputs(2387)) or (layer0_outputs(355)));
    layer1_outputs(1006) <= not(layer0_outputs(1513));
    layer1_outputs(1007) <= (layer0_outputs(2251)) and not (layer0_outputs(2245));
    layer1_outputs(1008) <= layer0_outputs(660);
    layer1_outputs(1009) <= (layer0_outputs(1702)) and not (layer0_outputs(789));
    layer1_outputs(1010) <= not((layer0_outputs(779)) or (layer0_outputs(428)));
    layer1_outputs(1011) <= (layer0_outputs(720)) or (layer0_outputs(2099));
    layer1_outputs(1012) <= not((layer0_outputs(2112)) xor (layer0_outputs(1311)));
    layer1_outputs(1013) <= (layer0_outputs(2140)) and (layer0_outputs(355));
    layer1_outputs(1014) <= not(layer0_outputs(837));
    layer1_outputs(1015) <= not(layer0_outputs(1190)) or (layer0_outputs(201));
    layer1_outputs(1016) <= not(layer0_outputs(328)) or (layer0_outputs(1446));
    layer1_outputs(1017) <= not(layer0_outputs(1289));
    layer1_outputs(1018) <= not(layer0_outputs(635)) or (layer0_outputs(2118));
    layer1_outputs(1019) <= layer0_outputs(444);
    layer1_outputs(1020) <= (layer0_outputs(567)) and not (layer0_outputs(407));
    layer1_outputs(1021) <= not(layer0_outputs(2102));
    layer1_outputs(1022) <= not((layer0_outputs(1703)) or (layer0_outputs(1696)));
    layer1_outputs(1023) <= (layer0_outputs(1558)) and (layer0_outputs(1381));
    layer1_outputs(1024) <= (layer0_outputs(2463)) or (layer0_outputs(159));
    layer1_outputs(1025) <= not(layer0_outputs(2066)) or (layer0_outputs(2358));
    layer1_outputs(1026) <= (layer0_outputs(2474)) and not (layer0_outputs(970));
    layer1_outputs(1027) <= not(layer0_outputs(222));
    layer1_outputs(1028) <= (layer0_outputs(433)) xor (layer0_outputs(1271));
    layer1_outputs(1029) <= (layer0_outputs(844)) and (layer0_outputs(2309));
    layer1_outputs(1030) <= not((layer0_outputs(864)) or (layer0_outputs(920)));
    layer1_outputs(1031) <= not(layer0_outputs(2379));
    layer1_outputs(1032) <= (layer0_outputs(1415)) and not (layer0_outputs(429));
    layer1_outputs(1033) <= not((layer0_outputs(2385)) or (layer0_outputs(2450)));
    layer1_outputs(1034) <= layer0_outputs(1568);
    layer1_outputs(1035) <= not(layer0_outputs(1729));
    layer1_outputs(1036) <= (layer0_outputs(2266)) and (layer0_outputs(6));
    layer1_outputs(1037) <= not(layer0_outputs(618)) or (layer0_outputs(638));
    layer1_outputs(1038) <= layer0_outputs(1799);
    layer1_outputs(1039) <= not(layer0_outputs(1717)) or (layer0_outputs(800));
    layer1_outputs(1040) <= '1';
    layer1_outputs(1041) <= (layer0_outputs(1408)) and not (layer0_outputs(1295));
    layer1_outputs(1042) <= not(layer0_outputs(1232));
    layer1_outputs(1043) <= (layer0_outputs(2407)) and (layer0_outputs(1915));
    layer1_outputs(1044) <= (layer0_outputs(1864)) and not (layer0_outputs(593));
    layer1_outputs(1045) <= (layer0_outputs(2198)) and not (layer0_outputs(1307));
    layer1_outputs(1046) <= not(layer0_outputs(1708)) or (layer0_outputs(2331));
    layer1_outputs(1047) <= not(layer0_outputs(1273)) or (layer0_outputs(580));
    layer1_outputs(1048) <= layer0_outputs(1480);
    layer1_outputs(1049) <= (layer0_outputs(1932)) xor (layer0_outputs(138));
    layer1_outputs(1050) <= not((layer0_outputs(262)) or (layer0_outputs(743)));
    layer1_outputs(1051) <= (layer0_outputs(734)) or (layer0_outputs(296));
    layer1_outputs(1052) <= (layer0_outputs(2169)) and (layer0_outputs(1229));
    layer1_outputs(1053) <= layer0_outputs(1899);
    layer1_outputs(1054) <= (layer0_outputs(1943)) and (layer0_outputs(2131));
    layer1_outputs(1055) <= not(layer0_outputs(2217));
    layer1_outputs(1056) <= (layer0_outputs(1094)) or (layer0_outputs(2147));
    layer1_outputs(1057) <= not(layer0_outputs(1121)) or (layer0_outputs(366));
    layer1_outputs(1058) <= (layer0_outputs(307)) or (layer0_outputs(85));
    layer1_outputs(1059) <= not(layer0_outputs(105));
    layer1_outputs(1060) <= not(layer0_outputs(97));
    layer1_outputs(1061) <= not(layer0_outputs(993));
    layer1_outputs(1062) <= not((layer0_outputs(394)) or (layer0_outputs(77)));
    layer1_outputs(1063) <= not(layer0_outputs(504));
    layer1_outputs(1064) <= '0';
    layer1_outputs(1065) <= (layer0_outputs(550)) or (layer0_outputs(818));
    layer1_outputs(1066) <= not(layer0_outputs(472)) or (layer0_outputs(1813));
    layer1_outputs(1067) <= not(layer0_outputs(170));
    layer1_outputs(1068) <= (layer0_outputs(1125)) or (layer0_outputs(760));
    layer1_outputs(1069) <= not((layer0_outputs(1684)) xor (layer0_outputs(1508)));
    layer1_outputs(1070) <= (layer0_outputs(2320)) and (layer0_outputs(1575));
    layer1_outputs(1071) <= not((layer0_outputs(874)) or (layer0_outputs(2541)));
    layer1_outputs(1072) <= not((layer0_outputs(8)) or (layer0_outputs(209)));
    layer1_outputs(1073) <= '1';
    layer1_outputs(1074) <= layer0_outputs(988);
    layer1_outputs(1075) <= (layer0_outputs(2278)) and not (layer0_outputs(1453));
    layer1_outputs(1076) <= not(layer0_outputs(1496));
    layer1_outputs(1077) <= layer0_outputs(1306);
    layer1_outputs(1078) <= (layer0_outputs(1435)) and not (layer0_outputs(174));
    layer1_outputs(1079) <= not((layer0_outputs(1776)) or (layer0_outputs(1356)));
    layer1_outputs(1080) <= (layer0_outputs(1380)) xor (layer0_outputs(2186));
    layer1_outputs(1081) <= not((layer0_outputs(2235)) and (layer0_outputs(2343)));
    layer1_outputs(1082) <= not(layer0_outputs(1465)) or (layer0_outputs(526));
    layer1_outputs(1083) <= (layer0_outputs(2447)) and not (layer0_outputs(1996));
    layer1_outputs(1084) <= '1';
    layer1_outputs(1085) <= (layer0_outputs(558)) xor (layer0_outputs(2086));
    layer1_outputs(1086) <= not(layer0_outputs(614));
    layer1_outputs(1087) <= not(layer0_outputs(549)) or (layer0_outputs(226));
    layer1_outputs(1088) <= not((layer0_outputs(1101)) or (layer0_outputs(1842)));
    layer1_outputs(1089) <= not(layer0_outputs(312));
    layer1_outputs(1090) <= layer0_outputs(902);
    layer1_outputs(1091) <= (layer0_outputs(452)) and not (layer0_outputs(369));
    layer1_outputs(1092) <= (layer0_outputs(2020)) and not (layer0_outputs(2399));
    layer1_outputs(1093) <= layer0_outputs(1316);
    layer1_outputs(1094) <= (layer0_outputs(71)) and not (layer0_outputs(41));
    layer1_outputs(1095) <= not(layer0_outputs(1469)) or (layer0_outputs(1035));
    layer1_outputs(1096) <= layer0_outputs(1215);
    layer1_outputs(1097) <= (layer0_outputs(835)) and not (layer0_outputs(1120));
    layer1_outputs(1098) <= not(layer0_outputs(495));
    layer1_outputs(1099) <= not(layer0_outputs(2157)) or (layer0_outputs(2065));
    layer1_outputs(1100) <= (layer0_outputs(1322)) xor (layer0_outputs(1958));
    layer1_outputs(1101) <= not((layer0_outputs(1077)) xor (layer0_outputs(2354)));
    layer1_outputs(1102) <= not(layer0_outputs(2502)) or (layer0_outputs(1830));
    layer1_outputs(1103) <= not((layer0_outputs(1542)) xor (layer0_outputs(1075)));
    layer1_outputs(1104) <= not(layer0_outputs(1195)) or (layer0_outputs(2227));
    layer1_outputs(1105) <= not(layer0_outputs(276));
    layer1_outputs(1106) <= not((layer0_outputs(2359)) and (layer0_outputs(298)));
    layer1_outputs(1107) <= (layer0_outputs(558)) and not (layer0_outputs(14));
    layer1_outputs(1108) <= not(layer0_outputs(703));
    layer1_outputs(1109) <= (layer0_outputs(2555)) and not (layer0_outputs(1224));
    layer1_outputs(1110) <= '1';
    layer1_outputs(1111) <= (layer0_outputs(1005)) or (layer0_outputs(1256));
    layer1_outputs(1112) <= not((layer0_outputs(2299)) xor (layer0_outputs(1384)));
    layer1_outputs(1113) <= not(layer0_outputs(2265)) or (layer0_outputs(841));
    layer1_outputs(1114) <= (layer0_outputs(1917)) and (layer0_outputs(89));
    layer1_outputs(1115) <= not(layer0_outputs(1146)) or (layer0_outputs(90));
    layer1_outputs(1116) <= not((layer0_outputs(1217)) or (layer0_outputs(1383)));
    layer1_outputs(1117) <= layer0_outputs(227);
    layer1_outputs(1118) <= '0';
    layer1_outputs(1119) <= (layer0_outputs(2083)) or (layer0_outputs(2038));
    layer1_outputs(1120) <= not((layer0_outputs(1098)) and (layer0_outputs(2182)));
    layer1_outputs(1121) <= '1';
    layer1_outputs(1122) <= (layer0_outputs(562)) or (layer0_outputs(2057));
    layer1_outputs(1123) <= not((layer0_outputs(2054)) or (layer0_outputs(2185)));
    layer1_outputs(1124) <= layer0_outputs(1327);
    layer1_outputs(1125) <= not((layer0_outputs(998)) and (layer0_outputs(1593)));
    layer1_outputs(1126) <= not(layer0_outputs(554));
    layer1_outputs(1127) <= not((layer0_outputs(2321)) and (layer0_outputs(1023)));
    layer1_outputs(1128) <= not((layer0_outputs(1481)) and (layer0_outputs(1520)));
    layer1_outputs(1129) <= not(layer0_outputs(687)) or (layer0_outputs(872));
    layer1_outputs(1130) <= layer0_outputs(2327);
    layer1_outputs(1131) <= '1';
    layer1_outputs(1132) <= not((layer0_outputs(258)) or (layer0_outputs(231)));
    layer1_outputs(1133) <= (layer0_outputs(1846)) or (layer0_outputs(967));
    layer1_outputs(1134) <= not(layer0_outputs(1033));
    layer1_outputs(1135) <= not(layer0_outputs(647)) or (layer0_outputs(1106));
    layer1_outputs(1136) <= '1';
    layer1_outputs(1137) <= not((layer0_outputs(2211)) and (layer0_outputs(773)));
    layer1_outputs(1138) <= (layer0_outputs(289)) and (layer0_outputs(2075));
    layer1_outputs(1139) <= not((layer0_outputs(1874)) and (layer0_outputs(1138)));
    layer1_outputs(1140) <= not((layer0_outputs(2323)) and (layer0_outputs(533)));
    layer1_outputs(1141) <= (layer0_outputs(885)) or (layer0_outputs(2298));
    layer1_outputs(1142) <= not(layer0_outputs(510));
    layer1_outputs(1143) <= not(layer0_outputs(1037));
    layer1_outputs(1144) <= not((layer0_outputs(2192)) or (layer0_outputs(1814)));
    layer1_outputs(1145) <= not(layer0_outputs(2470)) or (layer0_outputs(649));
    layer1_outputs(1146) <= (layer0_outputs(1308)) and not (layer0_outputs(1915));
    layer1_outputs(1147) <= not(layer0_outputs(1147)) or (layer0_outputs(897));
    layer1_outputs(1148) <= layer0_outputs(1386);
    layer1_outputs(1149) <= not(layer0_outputs(286));
    layer1_outputs(1150) <= not(layer0_outputs(1156));
    layer1_outputs(1151) <= not(layer0_outputs(636)) or (layer0_outputs(1510));
    layer1_outputs(1152) <= not(layer0_outputs(2070)) or (layer0_outputs(2330));
    layer1_outputs(1153) <= (layer0_outputs(1238)) and (layer0_outputs(2142));
    layer1_outputs(1154) <= not(layer0_outputs(1400)) or (layer0_outputs(1687));
    layer1_outputs(1155) <= '1';
    layer1_outputs(1156) <= layer0_outputs(674);
    layer1_outputs(1157) <= (layer0_outputs(2061)) and not (layer0_outputs(2536));
    layer1_outputs(1158) <= not(layer0_outputs(1596));
    layer1_outputs(1159) <= layer0_outputs(2429);
    layer1_outputs(1160) <= not((layer0_outputs(1070)) and (layer0_outputs(544)));
    layer1_outputs(1161) <= not(layer0_outputs(659));
    layer1_outputs(1162) <= (layer0_outputs(2006)) or (layer0_outputs(2394));
    layer1_outputs(1163) <= not((layer0_outputs(975)) or (layer0_outputs(1927)));
    layer1_outputs(1164) <= not((layer0_outputs(1732)) and (layer0_outputs(2499)));
    layer1_outputs(1165) <= '0';
    layer1_outputs(1166) <= (layer0_outputs(2384)) and (layer0_outputs(1303));
    layer1_outputs(1167) <= '1';
    layer1_outputs(1168) <= not((layer0_outputs(388)) or (layer0_outputs(1053)));
    layer1_outputs(1169) <= (layer0_outputs(1210)) and not (layer0_outputs(1623));
    layer1_outputs(1170) <= not((layer0_outputs(797)) and (layer0_outputs(798)));
    layer1_outputs(1171) <= not(layer0_outputs(249));
    layer1_outputs(1172) <= layer0_outputs(2301);
    layer1_outputs(1173) <= not((layer0_outputs(1821)) and (layer0_outputs(2217)));
    layer1_outputs(1174) <= '0';
    layer1_outputs(1175) <= not(layer0_outputs(834)) or (layer0_outputs(1718));
    layer1_outputs(1176) <= (layer0_outputs(2407)) and (layer0_outputs(2083));
    layer1_outputs(1177) <= not((layer0_outputs(799)) and (layer0_outputs(454)));
    layer1_outputs(1178) <= not(layer0_outputs(488));
    layer1_outputs(1179) <= not((layer0_outputs(1075)) xor (layer0_outputs(620)));
    layer1_outputs(1180) <= not(layer0_outputs(1261)) or (layer0_outputs(2470));
    layer1_outputs(1181) <= not((layer0_outputs(2120)) and (layer0_outputs(1809)));
    layer1_outputs(1182) <= not((layer0_outputs(1194)) or (layer0_outputs(1116)));
    layer1_outputs(1183) <= '0';
    layer1_outputs(1184) <= not(layer0_outputs(1606));
    layer1_outputs(1185) <= not(layer0_outputs(317));
    layer1_outputs(1186) <= not(layer0_outputs(373));
    layer1_outputs(1187) <= '1';
    layer1_outputs(1188) <= not(layer0_outputs(1069)) or (layer0_outputs(1331));
    layer1_outputs(1189) <= layer0_outputs(1402);
    layer1_outputs(1190) <= not(layer0_outputs(383));
    layer1_outputs(1191) <= layer0_outputs(435);
    layer1_outputs(1192) <= not(layer0_outputs(1100)) or (layer0_outputs(1969));
    layer1_outputs(1193) <= not(layer0_outputs(1757)) or (layer0_outputs(1249));
    layer1_outputs(1194) <= (layer0_outputs(2460)) and not (layer0_outputs(26));
    layer1_outputs(1195) <= (layer0_outputs(2440)) or (layer0_outputs(1017));
    layer1_outputs(1196) <= not(layer0_outputs(1171));
    layer1_outputs(1197) <= not((layer0_outputs(1646)) or (layer0_outputs(977)));
    layer1_outputs(1198) <= not((layer0_outputs(2465)) or (layer0_outputs(1918)));
    layer1_outputs(1199) <= not(layer0_outputs(652)) or (layer0_outputs(1577));
    layer1_outputs(1200) <= not(layer0_outputs(1398)) or (layer0_outputs(1379));
    layer1_outputs(1201) <= (layer0_outputs(828)) or (layer0_outputs(254));
    layer1_outputs(1202) <= not(layer0_outputs(1781));
    layer1_outputs(1203) <= not(layer0_outputs(2302));
    layer1_outputs(1204) <= '1';
    layer1_outputs(1205) <= not((layer0_outputs(1183)) and (layer0_outputs(1048)));
    layer1_outputs(1206) <= not((layer0_outputs(835)) and (layer0_outputs(2467)));
    layer1_outputs(1207) <= not(layer0_outputs(1130)) or (layer0_outputs(2014));
    layer1_outputs(1208) <= not(layer0_outputs(76)) or (layer0_outputs(956));
    layer1_outputs(1209) <= (layer0_outputs(2155)) and not (layer0_outputs(464));
    layer1_outputs(1210) <= '0';
    layer1_outputs(1211) <= not(layer0_outputs(888)) or (layer0_outputs(1743));
    layer1_outputs(1212) <= not(layer0_outputs(35));
    layer1_outputs(1213) <= '1';
    layer1_outputs(1214) <= not((layer0_outputs(1648)) and (layer0_outputs(1636)));
    layer1_outputs(1215) <= not(layer0_outputs(2163)) or (layer0_outputs(910));
    layer1_outputs(1216) <= not(layer0_outputs(1322)) or (layer0_outputs(682));
    layer1_outputs(1217) <= layer0_outputs(1272);
    layer1_outputs(1218) <= not((layer0_outputs(2162)) and (layer0_outputs(833)));
    layer1_outputs(1219) <= layer0_outputs(1792);
    layer1_outputs(1220) <= layer0_outputs(462);
    layer1_outputs(1221) <= not(layer0_outputs(1371));
    layer1_outputs(1222) <= layer0_outputs(1254);
    layer1_outputs(1223) <= (layer0_outputs(1135)) or (layer0_outputs(2376));
    layer1_outputs(1224) <= not(layer0_outputs(271)) or (layer0_outputs(976));
    layer1_outputs(1225) <= not(layer0_outputs(128));
    layer1_outputs(1226) <= (layer0_outputs(696)) and (layer0_outputs(5));
    layer1_outputs(1227) <= layer0_outputs(1644);
    layer1_outputs(1228) <= not(layer0_outputs(332)) or (layer0_outputs(403));
    layer1_outputs(1229) <= not(layer0_outputs(224));
    layer1_outputs(1230) <= (layer0_outputs(169)) or (layer0_outputs(1268));
    layer1_outputs(1231) <= (layer0_outputs(1561)) and not (layer0_outputs(293));
    layer1_outputs(1232) <= not(layer0_outputs(503));
    layer1_outputs(1233) <= (layer0_outputs(1312)) and not (layer0_outputs(1925));
    layer1_outputs(1234) <= (layer0_outputs(332)) and not (layer0_outputs(2004));
    layer1_outputs(1235) <= (layer0_outputs(476)) or (layer0_outputs(1072));
    layer1_outputs(1236) <= not(layer0_outputs(628)) or (layer0_outputs(589));
    layer1_outputs(1237) <= not(layer0_outputs(1005));
    layer1_outputs(1238) <= not(layer0_outputs(1640)) or (layer0_outputs(2053));
    layer1_outputs(1239) <= not((layer0_outputs(1903)) or (layer0_outputs(424)));
    layer1_outputs(1240) <= not(layer0_outputs(260));
    layer1_outputs(1241) <= not(layer0_outputs(1006)) or (layer0_outputs(2031));
    layer1_outputs(1242) <= (layer0_outputs(752)) and (layer0_outputs(2096));
    layer1_outputs(1243) <= '0';
    layer1_outputs(1244) <= not((layer0_outputs(1012)) or (layer0_outputs(2369)));
    layer1_outputs(1245) <= not((layer0_outputs(840)) and (layer0_outputs(516)));
    layer1_outputs(1246) <= '1';
    layer1_outputs(1247) <= (layer0_outputs(1940)) xor (layer0_outputs(1847));
    layer1_outputs(1248) <= layer0_outputs(2060);
    layer1_outputs(1249) <= (layer0_outputs(1375)) or (layer0_outputs(1109));
    layer1_outputs(1250) <= not(layer0_outputs(206)) or (layer0_outputs(1490));
    layer1_outputs(1251) <= (layer0_outputs(2374)) and not (layer0_outputs(169));
    layer1_outputs(1252) <= (layer0_outputs(80)) and not (layer0_outputs(1309));
    layer1_outputs(1253) <= not(layer0_outputs(2367));
    layer1_outputs(1254) <= '1';
    layer1_outputs(1255) <= not(layer0_outputs(384));
    layer1_outputs(1256) <= not(layer0_outputs(2221)) or (layer0_outputs(2073));
    layer1_outputs(1257) <= layer0_outputs(1558);
    layer1_outputs(1258) <= '1';
    layer1_outputs(1259) <= (layer0_outputs(604)) and (layer0_outputs(1143));
    layer1_outputs(1260) <= (layer0_outputs(2393)) and not (layer0_outputs(2322));
    layer1_outputs(1261) <= (layer0_outputs(1972)) or (layer0_outputs(2015));
    layer1_outputs(1262) <= (layer0_outputs(2457)) and not (layer0_outputs(2121));
    layer1_outputs(1263) <= (layer0_outputs(1320)) and not (layer0_outputs(582));
    layer1_outputs(1264) <= not(layer0_outputs(1827)) or (layer0_outputs(2538));
    layer1_outputs(1265) <= not((layer0_outputs(623)) or (layer0_outputs(1480)));
    layer1_outputs(1266) <= '1';
    layer1_outputs(1267) <= '0';
    layer1_outputs(1268) <= not(layer0_outputs(1811));
    layer1_outputs(1269) <= not((layer0_outputs(1538)) and (layer0_outputs(539)));
    layer1_outputs(1270) <= layer0_outputs(1806);
    layer1_outputs(1271) <= not((layer0_outputs(1404)) or (layer0_outputs(1527)));
    layer1_outputs(1272) <= '0';
    layer1_outputs(1273) <= not(layer0_outputs(1969));
    layer1_outputs(1274) <= not(layer0_outputs(1868)) or (layer0_outputs(2302));
    layer1_outputs(1275) <= not(layer0_outputs(2048)) or (layer0_outputs(2516));
    layer1_outputs(1276) <= not(layer0_outputs(588)) or (layer0_outputs(922));
    layer1_outputs(1277) <= (layer0_outputs(1875)) and not (layer0_outputs(1028));
    layer1_outputs(1278) <= not(layer0_outputs(717));
    layer1_outputs(1279) <= not((layer0_outputs(457)) or (layer0_outputs(2322)));
    layer1_outputs(1280) <= '1';
    layer1_outputs(1281) <= layer0_outputs(2025);
    layer1_outputs(1282) <= (layer0_outputs(1407)) and (layer0_outputs(620));
    layer1_outputs(1283) <= (layer0_outputs(187)) and not (layer0_outputs(2134));
    layer1_outputs(1284) <= layer0_outputs(1458);
    layer1_outputs(1285) <= layer0_outputs(1222);
    layer1_outputs(1286) <= (layer0_outputs(652)) and not (layer0_outputs(426));
    layer1_outputs(1287) <= layer0_outputs(1029);
    layer1_outputs(1288) <= (layer0_outputs(1284)) or (layer0_outputs(880));
    layer1_outputs(1289) <= layer0_outputs(707);
    layer1_outputs(1290) <= '0';
    layer1_outputs(1291) <= not(layer0_outputs(1357));
    layer1_outputs(1292) <= not((layer0_outputs(284)) or (layer0_outputs(2422)));
    layer1_outputs(1293) <= not(layer0_outputs(544)) or (layer0_outputs(940));
    layer1_outputs(1294) <= not((layer0_outputs(2426)) or (layer0_outputs(1902)));
    layer1_outputs(1295) <= layer0_outputs(1258);
    layer1_outputs(1296) <= not((layer0_outputs(1014)) or (layer0_outputs(1693)));
    layer1_outputs(1297) <= (layer0_outputs(1001)) and (layer0_outputs(810));
    layer1_outputs(1298) <= not(layer0_outputs(107));
    layer1_outputs(1299) <= layer0_outputs(814);
    layer1_outputs(1300) <= '0';
    layer1_outputs(1301) <= not(layer0_outputs(569));
    layer1_outputs(1302) <= not(layer0_outputs(1594));
    layer1_outputs(1303) <= (layer0_outputs(1921)) and not (layer0_outputs(2520));
    layer1_outputs(1304) <= (layer0_outputs(1569)) and not (layer0_outputs(2272));
    layer1_outputs(1305) <= not(layer0_outputs(2502)) or (layer0_outputs(1476));
    layer1_outputs(1306) <= not(layer0_outputs(1104));
    layer1_outputs(1307) <= not(layer0_outputs(560));
    layer1_outputs(1308) <= (layer0_outputs(1033)) and (layer0_outputs(2468));
    layer1_outputs(1309) <= not(layer0_outputs(293));
    layer1_outputs(1310) <= not(layer0_outputs(446)) or (layer0_outputs(1151));
    layer1_outputs(1311) <= layer0_outputs(1354);
    layer1_outputs(1312) <= not((layer0_outputs(1858)) and (layer0_outputs(603)));
    layer1_outputs(1313) <= not(layer0_outputs(1389));
    layer1_outputs(1314) <= (layer0_outputs(1296)) and (layer0_outputs(2242));
    layer1_outputs(1315) <= layer0_outputs(1022);
    layer1_outputs(1316) <= layer0_outputs(1617);
    layer1_outputs(1317) <= not(layer0_outputs(1618));
    layer1_outputs(1318) <= layer0_outputs(650);
    layer1_outputs(1319) <= '1';
    layer1_outputs(1320) <= '1';
    layer1_outputs(1321) <= (layer0_outputs(2249)) and not (layer0_outputs(2200));
    layer1_outputs(1322) <= not((layer0_outputs(542)) and (layer0_outputs(2198)));
    layer1_outputs(1323) <= not(layer0_outputs(1828));
    layer1_outputs(1324) <= (layer0_outputs(895)) and (layer0_outputs(2153));
    layer1_outputs(1325) <= (layer0_outputs(326)) and not (layer0_outputs(1429));
    layer1_outputs(1326) <= layer0_outputs(290);
    layer1_outputs(1327) <= not(layer0_outputs(2473)) or (layer0_outputs(767));
    layer1_outputs(1328) <= not(layer0_outputs(2451)) or (layer0_outputs(1566));
    layer1_outputs(1329) <= (layer0_outputs(2071)) xor (layer0_outputs(1493));
    layer1_outputs(1330) <= (layer0_outputs(1794)) and not (layer0_outputs(122));
    layer1_outputs(1331) <= layer0_outputs(134);
    layer1_outputs(1332) <= not((layer0_outputs(1114)) and (layer0_outputs(2104)));
    layer1_outputs(1333) <= (layer0_outputs(1330)) and not (layer0_outputs(1064));
    layer1_outputs(1334) <= not(layer0_outputs(92));
    layer1_outputs(1335) <= not(layer0_outputs(1949));
    layer1_outputs(1336) <= layer0_outputs(2318);
    layer1_outputs(1337) <= (layer0_outputs(1530)) or (layer0_outputs(2260));
    layer1_outputs(1338) <= layer0_outputs(1858);
    layer1_outputs(1339) <= not(layer0_outputs(547)) or (layer0_outputs(2111));
    layer1_outputs(1340) <= layer0_outputs(703);
    layer1_outputs(1341) <= not(layer0_outputs(762)) or (layer0_outputs(811));
    layer1_outputs(1342) <= (layer0_outputs(259)) or (layer0_outputs(584));
    layer1_outputs(1343) <= not((layer0_outputs(594)) or (layer0_outputs(1964)));
    layer1_outputs(1344) <= layer0_outputs(2504);
    layer1_outputs(1345) <= '0';
    layer1_outputs(1346) <= layer0_outputs(785);
    layer1_outputs(1347) <= not(layer0_outputs(399)) or (layer0_outputs(530));
    layer1_outputs(1348) <= (layer0_outputs(1367)) and not (layer0_outputs(475));
    layer1_outputs(1349) <= not(layer0_outputs(585));
    layer1_outputs(1350) <= not(layer0_outputs(1785)) or (layer0_outputs(2323));
    layer1_outputs(1351) <= (layer0_outputs(285)) or (layer0_outputs(840));
    layer1_outputs(1352) <= layer0_outputs(160);
    layer1_outputs(1353) <= layer0_outputs(1748);
    layer1_outputs(1354) <= layer0_outputs(676);
    layer1_outputs(1355) <= layer0_outputs(2497);
    layer1_outputs(1356) <= not(layer0_outputs(1428)) or (layer0_outputs(1333));
    layer1_outputs(1357) <= not((layer0_outputs(2304)) or (layer0_outputs(1665)));
    layer1_outputs(1358) <= (layer0_outputs(1889)) xor (layer0_outputs(635));
    layer1_outputs(1359) <= (layer0_outputs(818)) and not (layer0_outputs(2493));
    layer1_outputs(1360) <= not(layer0_outputs(163));
    layer1_outputs(1361) <= '0';
    layer1_outputs(1362) <= not(layer0_outputs(508));
    layer1_outputs(1363) <= layer0_outputs(167);
    layer1_outputs(1364) <= not(layer0_outputs(2230));
    layer1_outputs(1365) <= layer0_outputs(1930);
    layer1_outputs(1366) <= not((layer0_outputs(591)) or (layer0_outputs(1262)));
    layer1_outputs(1367) <= (layer0_outputs(1855)) or (layer0_outputs(2326));
    layer1_outputs(1368) <= layer0_outputs(233);
    layer1_outputs(1369) <= layer0_outputs(820);
    layer1_outputs(1370) <= (layer0_outputs(1481)) and not (layer0_outputs(683));
    layer1_outputs(1371) <= '0';
    layer1_outputs(1372) <= (layer0_outputs(1548)) or (layer0_outputs(2347));
    layer1_outputs(1373) <= (layer0_outputs(56)) or (layer0_outputs(1174));
    layer1_outputs(1374) <= layer0_outputs(1207);
    layer1_outputs(1375) <= not((layer0_outputs(1556)) and (layer0_outputs(2143)));
    layer1_outputs(1376) <= layer0_outputs(1499);
    layer1_outputs(1377) <= not((layer0_outputs(141)) and (layer0_outputs(1160)));
    layer1_outputs(1378) <= '0';
    layer1_outputs(1379) <= layer0_outputs(994);
    layer1_outputs(1380) <= not((layer0_outputs(2237)) and (layer0_outputs(1494)));
    layer1_outputs(1381) <= not(layer0_outputs(297));
    layer1_outputs(1382) <= (layer0_outputs(22)) and not (layer0_outputs(2267));
    layer1_outputs(1383) <= not(layer0_outputs(62));
    layer1_outputs(1384) <= not(layer0_outputs(2488));
    layer1_outputs(1385) <= (layer0_outputs(1362)) and (layer0_outputs(1992));
    layer1_outputs(1386) <= layer0_outputs(1587);
    layer1_outputs(1387) <= '1';
    layer1_outputs(1388) <= not((layer0_outputs(449)) or (layer0_outputs(337)));
    layer1_outputs(1389) <= layer0_outputs(638);
    layer1_outputs(1390) <= not((layer0_outputs(1791)) and (layer0_outputs(308)));
    layer1_outputs(1391) <= not(layer0_outputs(2167)) or (layer0_outputs(2514));
    layer1_outputs(1392) <= (layer0_outputs(2347)) xor (layer0_outputs(2351));
    layer1_outputs(1393) <= (layer0_outputs(93)) and (layer0_outputs(1419));
    layer1_outputs(1394) <= '0';
    layer1_outputs(1395) <= layer0_outputs(2319);
    layer1_outputs(1396) <= (layer0_outputs(501)) xor (layer0_outputs(2485));
    layer1_outputs(1397) <= (layer0_outputs(1642)) xor (layer0_outputs(2390));
    layer1_outputs(1398) <= layer0_outputs(304);
    layer1_outputs(1399) <= layer0_outputs(1167);
    layer1_outputs(1400) <= not(layer0_outputs(1544)) or (layer0_outputs(725));
    layer1_outputs(1401) <= not((layer0_outputs(564)) and (layer0_outputs(1983)));
    layer1_outputs(1402) <= layer0_outputs(2172);
    layer1_outputs(1403) <= (layer0_outputs(1738)) and not (layer0_outputs(1769));
    layer1_outputs(1404) <= (layer0_outputs(1654)) and not (layer0_outputs(984));
    layer1_outputs(1405) <= not(layer0_outputs(577));
    layer1_outputs(1406) <= not((layer0_outputs(70)) and (layer0_outputs(1210)));
    layer1_outputs(1407) <= not(layer0_outputs(2514)) or (layer0_outputs(2151));
    layer1_outputs(1408) <= not((layer0_outputs(1957)) or (layer0_outputs(2218)));
    layer1_outputs(1409) <= layer0_outputs(2111);
    layer1_outputs(1410) <= (layer0_outputs(57)) and not (layer0_outputs(1083));
    layer1_outputs(1411) <= (layer0_outputs(1926)) and not (layer0_outputs(2099));
    layer1_outputs(1412) <= not(layer0_outputs(2435)) or (layer0_outputs(1463));
    layer1_outputs(1413) <= (layer0_outputs(2116)) and not (layer0_outputs(1285));
    layer1_outputs(1414) <= (layer0_outputs(150)) or (layer0_outputs(2134));
    layer1_outputs(1415) <= not(layer0_outputs(1440)) or (layer0_outputs(274));
    layer1_outputs(1416) <= (layer0_outputs(2048)) and (layer0_outputs(1803));
    layer1_outputs(1417) <= not(layer0_outputs(1575)) or (layer0_outputs(735));
    layer1_outputs(1418) <= '0';
    layer1_outputs(1419) <= not(layer0_outputs(534));
    layer1_outputs(1420) <= (layer0_outputs(1368)) and (layer0_outputs(154));
    layer1_outputs(1421) <= '0';
    layer1_outputs(1422) <= '1';
    layer1_outputs(1423) <= (layer0_outputs(2427)) and not (layer0_outputs(1770));
    layer1_outputs(1424) <= layer0_outputs(2196);
    layer1_outputs(1425) <= '1';
    layer1_outputs(1426) <= (layer0_outputs(81)) or (layer0_outputs(445));
    layer1_outputs(1427) <= layer0_outputs(1413);
    layer1_outputs(1428) <= not((layer0_outputs(745)) or (layer0_outputs(766)));
    layer1_outputs(1429) <= not(layer0_outputs(1376));
    layer1_outputs(1430) <= not((layer0_outputs(1622)) or (layer0_outputs(612)));
    layer1_outputs(1431) <= not(layer0_outputs(1057));
    layer1_outputs(1432) <= not(layer0_outputs(690)) or (layer0_outputs(443));
    layer1_outputs(1433) <= not(layer0_outputs(680));
    layer1_outputs(1434) <= not((layer0_outputs(2225)) and (layer0_outputs(2101)));
    layer1_outputs(1435) <= (layer0_outputs(32)) and not (layer0_outputs(2161));
    layer1_outputs(1436) <= layer0_outputs(1037);
    layer1_outputs(1437) <= (layer0_outputs(2491)) and not (layer0_outputs(427));
    layer1_outputs(1438) <= not(layer0_outputs(1683));
    layer1_outputs(1439) <= not((layer0_outputs(2343)) or (layer0_outputs(2059)));
    layer1_outputs(1440) <= not(layer0_outputs(1833));
    layer1_outputs(1441) <= not(layer0_outputs(836));
    layer1_outputs(1442) <= not(layer0_outputs(1891));
    layer1_outputs(1443) <= not(layer0_outputs(2372));
    layer1_outputs(1444) <= (layer0_outputs(1948)) and not (layer0_outputs(540));
    layer1_outputs(1445) <= not(layer0_outputs(603));
    layer1_outputs(1446) <= not(layer0_outputs(186));
    layer1_outputs(1447) <= layer0_outputs(439);
    layer1_outputs(1448) <= layer0_outputs(389);
    layer1_outputs(1449) <= layer0_outputs(745);
    layer1_outputs(1450) <= layer0_outputs(222);
    layer1_outputs(1451) <= not(layer0_outputs(641));
    layer1_outputs(1452) <= (layer0_outputs(1198)) and (layer0_outputs(1668));
    layer1_outputs(1453) <= not(layer0_outputs(650));
    layer1_outputs(1454) <= not(layer0_outputs(1158));
    layer1_outputs(1455) <= layer0_outputs(1779);
    layer1_outputs(1456) <= not(layer0_outputs(1412));
    layer1_outputs(1457) <= (layer0_outputs(1494)) and (layer0_outputs(1540));
    layer1_outputs(1458) <= layer0_outputs(1438);
    layer1_outputs(1459) <= not(layer0_outputs(331)) or (layer0_outputs(2442));
    layer1_outputs(1460) <= not(layer0_outputs(1034));
    layer1_outputs(1461) <= '1';
    layer1_outputs(1462) <= not(layer0_outputs(2088));
    layer1_outputs(1463) <= not(layer0_outputs(2055));
    layer1_outputs(1464) <= not((layer0_outputs(1200)) xor (layer0_outputs(878)));
    layer1_outputs(1465) <= (layer0_outputs(407)) or (layer0_outputs(255));
    layer1_outputs(1466) <= not(layer0_outputs(135));
    layer1_outputs(1467) <= layer0_outputs(2483);
    layer1_outputs(1468) <= (layer0_outputs(100)) and not (layer0_outputs(431));
    layer1_outputs(1469) <= (layer0_outputs(2112)) and not (layer0_outputs(2346));
    layer1_outputs(1470) <= not((layer0_outputs(2003)) xor (layer0_outputs(1343)));
    layer1_outputs(1471) <= (layer0_outputs(2123)) and not (layer0_outputs(660));
    layer1_outputs(1472) <= (layer0_outputs(1977)) and not (layer0_outputs(815));
    layer1_outputs(1473) <= (layer0_outputs(116)) and not (layer0_outputs(2500));
    layer1_outputs(1474) <= not(layer0_outputs(723));
    layer1_outputs(1475) <= (layer0_outputs(106)) and not (layer0_outputs(2165));
    layer1_outputs(1476) <= '1';
    layer1_outputs(1477) <= (layer0_outputs(957)) and not (layer0_outputs(390));
    layer1_outputs(1478) <= layer0_outputs(189);
    layer1_outputs(1479) <= not((layer0_outputs(2311)) or (layer0_outputs(1315)));
    layer1_outputs(1480) <= (layer0_outputs(621)) and (layer0_outputs(1482));
    layer1_outputs(1481) <= layer0_outputs(980);
    layer1_outputs(1482) <= (layer0_outputs(1842)) and not (layer0_outputs(688));
    layer1_outputs(1483) <= not(layer0_outputs(915));
    layer1_outputs(1484) <= (layer0_outputs(1775)) and not (layer0_outputs(1977));
    layer1_outputs(1485) <= (layer0_outputs(1159)) or (layer0_outputs(267));
    layer1_outputs(1486) <= '1';
    layer1_outputs(1487) <= '0';
    layer1_outputs(1488) <= not(layer0_outputs(922)) or (layer0_outputs(1002));
    layer1_outputs(1489) <= (layer0_outputs(1179)) and not (layer0_outputs(860));
    layer1_outputs(1490) <= not(layer0_outputs(944));
    layer1_outputs(1491) <= layer0_outputs(2032);
    layer1_outputs(1492) <= layer0_outputs(352);
    layer1_outputs(1493) <= not(layer0_outputs(1853));
    layer1_outputs(1494) <= layer0_outputs(341);
    layer1_outputs(1495) <= not((layer0_outputs(1924)) and (layer0_outputs(49)));
    layer1_outputs(1496) <= (layer0_outputs(2127)) or (layer0_outputs(768));
    layer1_outputs(1497) <= not((layer0_outputs(615)) and (layer0_outputs(2300)));
    layer1_outputs(1498) <= not(layer0_outputs(1576));
    layer1_outputs(1499) <= not(layer0_outputs(1427));
    layer1_outputs(1500) <= '0';
    layer1_outputs(1501) <= not((layer0_outputs(1681)) or (layer0_outputs(1365)));
    layer1_outputs(1502) <= not(layer0_outputs(2194));
    layer1_outputs(1503) <= layer0_outputs(983);
    layer1_outputs(1504) <= not(layer0_outputs(850));
    layer1_outputs(1505) <= layer0_outputs(2379);
    layer1_outputs(1506) <= (layer0_outputs(329)) and not (layer0_outputs(2452));
    layer1_outputs(1507) <= (layer0_outputs(1104)) or (layer0_outputs(1467));
    layer1_outputs(1508) <= not(layer0_outputs(13));
    layer1_outputs(1509) <= (layer0_outputs(1324)) and (layer0_outputs(2441));
    layer1_outputs(1510) <= (layer0_outputs(928)) and (layer0_outputs(2469));
    layer1_outputs(1511) <= layer0_outputs(1380);
    layer1_outputs(1512) <= '0';
    layer1_outputs(1513) <= not((layer0_outputs(1770)) or (layer0_outputs(263)));
    layer1_outputs(1514) <= not((layer0_outputs(576)) and (layer0_outputs(2100)));
    layer1_outputs(1515) <= layer0_outputs(205);
    layer1_outputs(1516) <= not((layer0_outputs(1611)) or (layer0_outputs(663)));
    layer1_outputs(1517) <= not(layer0_outputs(1572));
    layer1_outputs(1518) <= not(layer0_outputs(2074)) or (layer0_outputs(1942));
    layer1_outputs(1519) <= not(layer0_outputs(2381));
    layer1_outputs(1520) <= (layer0_outputs(1616)) and not (layer0_outputs(157));
    layer1_outputs(1521) <= not(layer0_outputs(83)) or (layer0_outputs(1036));
    layer1_outputs(1522) <= (layer0_outputs(1399)) and not (layer0_outputs(1713));
    layer1_outputs(1523) <= not(layer0_outputs(474));
    layer1_outputs(1524) <= (layer0_outputs(2439)) and not (layer0_outputs(1164));
    layer1_outputs(1525) <= (layer0_outputs(1997)) and (layer0_outputs(1393));
    layer1_outputs(1526) <= '1';
    layer1_outputs(1527) <= (layer0_outputs(2214)) and not (layer0_outputs(2373));
    layer1_outputs(1528) <= (layer0_outputs(563)) and not (layer0_outputs(1677));
    layer1_outputs(1529) <= (layer0_outputs(404)) and not (layer0_outputs(433));
    layer1_outputs(1530) <= not((layer0_outputs(2091)) and (layer0_outputs(2538)));
    layer1_outputs(1531) <= (layer0_outputs(1238)) and not (layer0_outputs(1218));
    layer1_outputs(1532) <= not(layer0_outputs(489)) or (layer0_outputs(2100));
    layer1_outputs(1533) <= layer0_outputs(1004);
    layer1_outputs(1534) <= layer0_outputs(1988);
    layer1_outputs(1535) <= (layer0_outputs(4)) and not (layer0_outputs(1780));
    layer1_outputs(1536) <= not(layer0_outputs(189));
    layer1_outputs(1537) <= layer0_outputs(1960);
    layer1_outputs(1538) <= (layer0_outputs(886)) or (layer0_outputs(2518));
    layer1_outputs(1539) <= (layer0_outputs(962)) and (layer0_outputs(803));
    layer1_outputs(1540) <= not(layer0_outputs(2507));
    layer1_outputs(1541) <= '0';
    layer1_outputs(1542) <= not((layer0_outputs(949)) or (layer0_outputs(294)));
    layer1_outputs(1543) <= '1';
    layer1_outputs(1544) <= (layer0_outputs(95)) xor (layer0_outputs(981));
    layer1_outputs(1545) <= not(layer0_outputs(2490));
    layer1_outputs(1546) <= not(layer0_outputs(106));
    layer1_outputs(1547) <= not(layer0_outputs(2144));
    layer1_outputs(1548) <= (layer0_outputs(1091)) or (layer0_outputs(2202));
    layer1_outputs(1549) <= (layer0_outputs(117)) and not (layer0_outputs(1242));
    layer1_outputs(1550) <= not(layer0_outputs(1087));
    layer1_outputs(1551) <= '0';
    layer1_outputs(1552) <= (layer0_outputs(1586)) and not (layer0_outputs(1935));
    layer1_outputs(1553) <= (layer0_outputs(137)) and not (layer0_outputs(866));
    layer1_outputs(1554) <= not(layer0_outputs(753));
    layer1_outputs(1555) <= not(layer0_outputs(1516));
    layer1_outputs(1556) <= layer0_outputs(1994);
    layer1_outputs(1557) <= not(layer0_outputs(2243)) or (layer0_outputs(666));
    layer1_outputs(1558) <= layer0_outputs(511);
    layer1_outputs(1559) <= (layer0_outputs(1773)) and (layer0_outputs(1802));
    layer1_outputs(1560) <= (layer0_outputs(2315)) and (layer0_outputs(702));
    layer1_outputs(1561) <= (layer0_outputs(918)) and not (layer0_outputs(1857));
    layer1_outputs(1562) <= not(layer0_outputs(648));
    layer1_outputs(1563) <= (layer0_outputs(2072)) and (layer0_outputs(418));
    layer1_outputs(1564) <= not(layer0_outputs(2401));
    layer1_outputs(1565) <= not((layer0_outputs(2132)) or (layer0_outputs(317)));
    layer1_outputs(1566) <= not(layer0_outputs(1663));
    layer1_outputs(1567) <= (layer0_outputs(86)) or (layer0_outputs(272));
    layer1_outputs(1568) <= layer0_outputs(808);
    layer1_outputs(1569) <= (layer0_outputs(396)) and not (layer0_outputs(2056));
    layer1_outputs(1570) <= (layer0_outputs(1200)) or (layer0_outputs(799));
    layer1_outputs(1571) <= layer0_outputs(1137);
    layer1_outputs(1572) <= not(layer0_outputs(1335)) or (layer0_outputs(48));
    layer1_outputs(1573) <= (layer0_outputs(2012)) and (layer0_outputs(2203));
    layer1_outputs(1574) <= not(layer0_outputs(653));
    layer1_outputs(1575) <= (layer0_outputs(2062)) and (layer0_outputs(1800));
    layer1_outputs(1576) <= not((layer0_outputs(2195)) and (layer0_outputs(195)));
    layer1_outputs(1577) <= not(layer0_outputs(1992));
    layer1_outputs(1578) <= not(layer0_outputs(2291));
    layer1_outputs(1579) <= not((layer0_outputs(856)) or (layer0_outputs(2095)));
    layer1_outputs(1580) <= not((layer0_outputs(11)) or (layer0_outputs(1028)));
    layer1_outputs(1581) <= layer0_outputs(601);
    layer1_outputs(1582) <= not((layer0_outputs(340)) and (layer0_outputs(2188)));
    layer1_outputs(1583) <= not(layer0_outputs(1952)) or (layer0_outputs(625));
    layer1_outputs(1584) <= layer0_outputs(559);
    layer1_outputs(1585) <= not(layer0_outputs(803)) or (layer0_outputs(870));
    layer1_outputs(1586) <= (layer0_outputs(1814)) and not (layer0_outputs(1031));
    layer1_outputs(1587) <= not((layer0_outputs(1961)) or (layer0_outputs(1204)));
    layer1_outputs(1588) <= layer0_outputs(1688);
    layer1_outputs(1589) <= not((layer0_outputs(416)) and (layer0_outputs(1500)));
    layer1_outputs(1590) <= not((layer0_outputs(1564)) or (layer0_outputs(632)));
    layer1_outputs(1591) <= layer0_outputs(1559);
    layer1_outputs(1592) <= (layer0_outputs(756)) and (layer0_outputs(608));
    layer1_outputs(1593) <= layer0_outputs(1402);
    layer1_outputs(1594) <= not(layer0_outputs(1158));
    layer1_outputs(1595) <= not(layer0_outputs(2260)) or (layer0_outputs(1090));
    layer1_outputs(1596) <= not(layer0_outputs(12)) or (layer0_outputs(1716));
    layer1_outputs(1597) <= not(layer0_outputs(457));
    layer1_outputs(1598) <= (layer0_outputs(381)) and (layer0_outputs(165));
    layer1_outputs(1599) <= (layer0_outputs(2300)) xor (layer0_outputs(809));
    layer1_outputs(1600) <= not(layer0_outputs(822)) or (layer0_outputs(2274));
    layer1_outputs(1601) <= not(layer0_outputs(294));
    layer1_outputs(1602) <= (layer0_outputs(677)) or (layer0_outputs(1718));
    layer1_outputs(1603) <= '0';
    layer1_outputs(1604) <= not(layer0_outputs(1609));
    layer1_outputs(1605) <= (layer0_outputs(1798)) and (layer0_outputs(289));
    layer1_outputs(1606) <= not(layer0_outputs(1628));
    layer1_outputs(1607) <= not((layer0_outputs(2068)) and (layer0_outputs(422)));
    layer1_outputs(1608) <= not(layer0_outputs(1676)) or (layer0_outputs(2486));
    layer1_outputs(1609) <= layer0_outputs(955);
    layer1_outputs(1610) <= (layer0_outputs(1999)) or (layer0_outputs(2164));
    layer1_outputs(1611) <= layer0_outputs(2309);
    layer1_outputs(1612) <= not(layer0_outputs(2156));
    layer1_outputs(1613) <= (layer0_outputs(2363)) xor (layer0_outputs(1441));
    layer1_outputs(1614) <= (layer0_outputs(133)) and (layer0_outputs(2548));
    layer1_outputs(1615) <= (layer0_outputs(1714)) and (layer0_outputs(998));
    layer1_outputs(1616) <= not((layer0_outputs(947)) or (layer0_outputs(444)));
    layer1_outputs(1617) <= layer0_outputs(531);
    layer1_outputs(1618) <= not(layer0_outputs(1278)) or (layer0_outputs(16));
    layer1_outputs(1619) <= (layer0_outputs(645)) and not (layer0_outputs(877));
    layer1_outputs(1620) <= layer0_outputs(1478);
    layer1_outputs(1621) <= not(layer0_outputs(436)) or (layer0_outputs(2233));
    layer1_outputs(1622) <= not(layer0_outputs(1226));
    layer1_outputs(1623) <= '1';
    layer1_outputs(1624) <= not(layer0_outputs(1439)) or (layer0_outputs(2001));
    layer1_outputs(1625) <= not(layer0_outputs(2267));
    layer1_outputs(1626) <= not(layer0_outputs(453)) or (layer0_outputs(353));
    layer1_outputs(1627) <= layer0_outputs(1164);
    layer1_outputs(1628) <= (layer0_outputs(1485)) and (layer0_outputs(2386));
    layer1_outputs(1629) <= not(layer0_outputs(2475)) or (layer0_outputs(2042));
    layer1_outputs(1630) <= not(layer0_outputs(1788)) or (layer0_outputs(2051));
    layer1_outputs(1631) <= (layer0_outputs(602)) and not (layer0_outputs(458));
    layer1_outputs(1632) <= (layer0_outputs(682)) and not (layer0_outputs(173));
    layer1_outputs(1633) <= (layer0_outputs(2097)) and not (layer0_outputs(866));
    layer1_outputs(1634) <= not(layer0_outputs(1067));
    layer1_outputs(1635) <= not((layer0_outputs(59)) or (layer0_outputs(232)));
    layer1_outputs(1636) <= layer0_outputs(2236);
    layer1_outputs(1637) <= not(layer0_outputs(150));
    layer1_outputs(1638) <= layer0_outputs(1092);
    layer1_outputs(1639) <= layer0_outputs(136);
    layer1_outputs(1640) <= layer0_outputs(968);
    layer1_outputs(1641) <= not(layer0_outputs(609));
    layer1_outputs(1642) <= (layer0_outputs(22)) and not (layer0_outputs(1196));
    layer1_outputs(1643) <= layer0_outputs(694);
    layer1_outputs(1644) <= not((layer0_outputs(759)) and (layer0_outputs(2094)));
    layer1_outputs(1645) <= not((layer0_outputs(1209)) and (layer0_outputs(2487)));
    layer1_outputs(1646) <= (layer0_outputs(1081)) and not (layer0_outputs(1406));
    layer1_outputs(1647) <= (layer0_outputs(1470)) and not (layer0_outputs(118));
    layer1_outputs(1648) <= (layer0_outputs(1366)) and not (layer0_outputs(2314));
    layer1_outputs(1649) <= (layer0_outputs(2483)) and not (layer0_outputs(186));
    layer1_outputs(1650) <= layer0_outputs(354);
    layer1_outputs(1651) <= not(layer0_outputs(165)) or (layer0_outputs(1711));
    layer1_outputs(1652) <= (layer0_outputs(80)) and not (layer0_outputs(64));
    layer1_outputs(1653) <= not((layer0_outputs(2230)) and (layer0_outputs(2051)));
    layer1_outputs(1654) <= not(layer0_outputs(1757));
    layer1_outputs(1655) <= not(layer0_outputs(590)) or (layer0_outputs(2459));
    layer1_outputs(1656) <= (layer0_outputs(894)) and not (layer0_outputs(778));
    layer1_outputs(1657) <= not((layer0_outputs(2352)) xor (layer0_outputs(54)));
    layer1_outputs(1658) <= not(layer0_outputs(2427)) or (layer0_outputs(791));
    layer1_outputs(1659) <= layer0_outputs(246);
    layer1_outputs(1660) <= not(layer0_outputs(2106)) or (layer0_outputs(1723));
    layer1_outputs(1661) <= (layer0_outputs(823)) and (layer0_outputs(297));
    layer1_outputs(1662) <= not(layer0_outputs(2536));
    layer1_outputs(1663) <= (layer0_outputs(63)) and not (layer0_outputs(303));
    layer1_outputs(1664) <= (layer0_outputs(1580)) and (layer0_outputs(855));
    layer1_outputs(1665) <= layer0_outputs(1113);
    layer1_outputs(1666) <= not(layer0_outputs(2177)) or (layer0_outputs(1522));
    layer1_outputs(1667) <= not(layer0_outputs(854));
    layer1_outputs(1668) <= (layer0_outputs(586)) and not (layer0_outputs(2012));
    layer1_outputs(1669) <= not(layer0_outputs(2062));
    layer1_outputs(1670) <= not(layer0_outputs(488));
    layer1_outputs(1671) <= (layer0_outputs(1697)) and not (layer0_outputs(2080));
    layer1_outputs(1672) <= not((layer0_outputs(1540)) or (layer0_outputs(797)));
    layer1_outputs(1673) <= layer0_outputs(2326);
    layer1_outputs(1674) <= layer0_outputs(859);
    layer1_outputs(1675) <= (layer0_outputs(691)) or (layer0_outputs(2356));
    layer1_outputs(1676) <= layer0_outputs(2517);
    layer1_outputs(1677) <= not(layer0_outputs(1578)) or (layer0_outputs(1173));
    layer1_outputs(1678) <= layer0_outputs(535);
    layer1_outputs(1679) <= layer0_outputs(100);
    layer1_outputs(1680) <= layer0_outputs(1796);
    layer1_outputs(1681) <= not(layer0_outputs(6));
    layer1_outputs(1682) <= not((layer0_outputs(42)) and (layer0_outputs(1311)));
    layer1_outputs(1683) <= not((layer0_outputs(1639)) and (layer0_outputs(954)));
    layer1_outputs(1684) <= layer0_outputs(974);
    layer1_outputs(1685) <= not(layer0_outputs(1667)) or (layer0_outputs(1049));
    layer1_outputs(1686) <= '1';
    layer1_outputs(1687) <= not((layer0_outputs(1883)) or (layer0_outputs(193)));
    layer1_outputs(1688) <= layer0_outputs(1666);
    layer1_outputs(1689) <= layer0_outputs(1314);
    layer1_outputs(1690) <= not(layer0_outputs(421)) or (layer0_outputs(2262));
    layer1_outputs(1691) <= (layer0_outputs(1972)) or (layer0_outputs(1267));
    layer1_outputs(1692) <= not((layer0_outputs(2360)) and (layer0_outputs(2261)));
    layer1_outputs(1693) <= not(layer0_outputs(2445)) or (layer0_outputs(170));
    layer1_outputs(1694) <= (layer0_outputs(1852)) and not (layer0_outputs(1568));
    layer1_outputs(1695) <= layer0_outputs(1285);
    layer1_outputs(1696) <= not(layer0_outputs(184)) or (layer0_outputs(2084));
    layer1_outputs(1697) <= (layer0_outputs(506)) and not (layer0_outputs(1346));
    layer1_outputs(1698) <= '0';
    layer1_outputs(1699) <= not(layer0_outputs(492)) or (layer0_outputs(386));
    layer1_outputs(1700) <= '0';
    layer1_outputs(1701) <= layer0_outputs(948);
    layer1_outputs(1702) <= layer0_outputs(1506);
    layer1_outputs(1703) <= layer0_outputs(1157);
    layer1_outputs(1704) <= not(layer0_outputs(902));
    layer1_outputs(1705) <= not(layer0_outputs(203)) or (layer0_outputs(2119));
    layer1_outputs(1706) <= (layer0_outputs(2269)) and not (layer0_outputs(2223));
    layer1_outputs(1707) <= not((layer0_outputs(147)) or (layer0_outputs(2011)));
    layer1_outputs(1708) <= layer0_outputs(1289);
    layer1_outputs(1709) <= not(layer0_outputs(982));
    layer1_outputs(1710) <= layer0_outputs(1170);
    layer1_outputs(1711) <= not((layer0_outputs(1048)) or (layer0_outputs(1018)));
    layer1_outputs(1712) <= not(layer0_outputs(330));
    layer1_outputs(1713) <= (layer0_outputs(1012)) and not (layer0_outputs(1600));
    layer1_outputs(1714) <= layer0_outputs(1353);
    layer1_outputs(1715) <= (layer0_outputs(2175)) and not (layer0_outputs(65));
    layer1_outputs(1716) <= not(layer0_outputs(1994));
    layer1_outputs(1717) <= layer0_outputs(2558);
    layer1_outputs(1718) <= not(layer0_outputs(629));
    layer1_outputs(1719) <= not(layer0_outputs(1877));
    layer1_outputs(1720) <= layer0_outputs(240);
    layer1_outputs(1721) <= not(layer0_outputs(1091)) or (layer0_outputs(43));
    layer1_outputs(1722) <= not(layer0_outputs(547));
    layer1_outputs(1723) <= '0';
    layer1_outputs(1724) <= (layer0_outputs(826)) and not (layer0_outputs(691));
    layer1_outputs(1725) <= not(layer0_outputs(26)) or (layer0_outputs(570));
    layer1_outputs(1726) <= layer0_outputs(1865);
    layer1_outputs(1727) <= (layer0_outputs(2497)) or (layer0_outputs(2244));
    layer1_outputs(1728) <= '1';
    layer1_outputs(1729) <= layer0_outputs(1622);
    layer1_outputs(1730) <= not(layer0_outputs(1645)) or (layer0_outputs(1356));
    layer1_outputs(1731) <= not(layer0_outputs(132)) or (layer0_outputs(1979));
    layer1_outputs(1732) <= (layer0_outputs(2228)) or (layer0_outputs(730));
    layer1_outputs(1733) <= '1';
    layer1_outputs(1734) <= '1';
    layer1_outputs(1735) <= not((layer0_outputs(1944)) or (layer0_outputs(1916)));
    layer1_outputs(1736) <= (layer0_outputs(12)) and (layer0_outputs(851));
    layer1_outputs(1737) <= (layer0_outputs(283)) or (layer0_outputs(2521));
    layer1_outputs(1738) <= (layer0_outputs(577)) or (layer0_outputs(868));
    layer1_outputs(1739) <= '1';
    layer1_outputs(1740) <= not(layer0_outputs(1686));
    layer1_outputs(1741) <= not(layer0_outputs(33));
    layer1_outputs(1742) <= not(layer0_outputs(882));
    layer1_outputs(1743) <= (layer0_outputs(1995)) and not (layer0_outputs(2292));
    layer1_outputs(1744) <= layer0_outputs(2130);
    layer1_outputs(1745) <= (layer0_outputs(549)) and not (layer0_outputs(1693));
    layer1_outputs(1746) <= '1';
    layer1_outputs(1747) <= layer0_outputs(1908);
    layer1_outputs(1748) <= layer0_outputs(254);
    layer1_outputs(1749) <= not(layer0_outputs(1466)) or (layer0_outputs(417));
    layer1_outputs(1750) <= layer0_outputs(506);
    layer1_outputs(1751) <= not(layer0_outputs(961));
    layer1_outputs(1752) <= layer0_outputs(748);
    layer1_outputs(1753) <= not(layer0_outputs(2411));
    layer1_outputs(1754) <= (layer0_outputs(819)) and not (layer0_outputs(1611));
    layer1_outputs(1755) <= not(layer0_outputs(672));
    layer1_outputs(1756) <= not((layer0_outputs(2460)) or (layer0_outputs(1056)));
    layer1_outputs(1757) <= '0';
    layer1_outputs(1758) <= not(layer0_outputs(1630)) or (layer0_outputs(1867));
    layer1_outputs(1759) <= not((layer0_outputs(2442)) or (layer0_outputs(2468)));
    layer1_outputs(1760) <= not((layer0_outputs(987)) or (layer0_outputs(1888)));
    layer1_outputs(1761) <= layer0_outputs(218);
    layer1_outputs(1762) <= not(layer0_outputs(743));
    layer1_outputs(1763) <= layer0_outputs(1488);
    layer1_outputs(1764) <= layer0_outputs(1095);
    layer1_outputs(1765) <= not((layer0_outputs(1797)) or (layer0_outputs(401)));
    layer1_outputs(1766) <= layer0_outputs(1746);
    layer1_outputs(1767) <= not(layer0_outputs(1251));
    layer1_outputs(1768) <= '1';
    layer1_outputs(1769) <= layer0_outputs(898);
    layer1_outputs(1770) <= not(layer0_outputs(1648));
    layer1_outputs(1771) <= not((layer0_outputs(1464)) and (layer0_outputs(668)));
    layer1_outputs(1772) <= not(layer0_outputs(1709));
    layer1_outputs(1773) <= (layer0_outputs(498)) or (layer0_outputs(1511));
    layer1_outputs(1774) <= not(layer0_outputs(2259));
    layer1_outputs(1775) <= not(layer0_outputs(328));
    layer1_outputs(1776) <= (layer0_outputs(215)) and (layer0_outputs(1684));
    layer1_outputs(1777) <= layer0_outputs(1434);
    layer1_outputs(1778) <= not(layer0_outputs(1240));
    layer1_outputs(1779) <= not(layer0_outputs(833));
    layer1_outputs(1780) <= (layer0_outputs(1603)) xor (layer0_outputs(1614));
    layer1_outputs(1781) <= not(layer0_outputs(955));
    layer1_outputs(1782) <= (layer0_outputs(1423)) and not (layer0_outputs(1579));
    layer1_outputs(1783) <= not(layer0_outputs(2432));
    layer1_outputs(1784) <= layer0_outputs(2109);
    layer1_outputs(1785) <= (layer0_outputs(242)) and (layer0_outputs(183));
    layer1_outputs(1786) <= (layer0_outputs(1454)) and not (layer0_outputs(1326));
    layer1_outputs(1787) <= not(layer0_outputs(2045));
    layer1_outputs(1788) <= not(layer0_outputs(2160));
    layer1_outputs(1789) <= not(layer0_outputs(755)) or (layer0_outputs(1838));
    layer1_outputs(1790) <= not(layer0_outputs(1139));
    layer1_outputs(1791) <= layer0_outputs(619);
    layer1_outputs(1792) <= not(layer0_outputs(1521));
    layer1_outputs(1793) <= layer0_outputs(202);
    layer1_outputs(1794) <= not(layer0_outputs(1841));
    layer1_outputs(1795) <= not(layer0_outputs(2150));
    layer1_outputs(1796) <= not(layer0_outputs(338));
    layer1_outputs(1797) <= layer0_outputs(2152);
    layer1_outputs(1798) <= layer0_outputs(788);
    layer1_outputs(1799) <= not(layer0_outputs(109));
    layer1_outputs(1800) <= '0';
    layer1_outputs(1801) <= not(layer0_outputs(1815));
    layer1_outputs(1802) <= layer0_outputs(2034);
    layer1_outputs(1803) <= layer0_outputs(801);
    layer1_outputs(1804) <= (layer0_outputs(1570)) or (layer0_outputs(2529));
    layer1_outputs(1805) <= (layer0_outputs(86)) and not (layer0_outputs(2110));
    layer1_outputs(1806) <= layer0_outputs(199);
    layer1_outputs(1807) <= (layer0_outputs(31)) xor (layer0_outputs(539));
    layer1_outputs(1808) <= '1';
    layer1_outputs(1809) <= not((layer0_outputs(1475)) or (layer0_outputs(315)));
    layer1_outputs(1810) <= not((layer0_outputs(382)) xor (layer0_outputs(779)));
    layer1_outputs(1811) <= (layer0_outputs(119)) and not (layer0_outputs(1202));
    layer1_outputs(1812) <= not(layer0_outputs(2203));
    layer1_outputs(1813) <= (layer0_outputs(2249)) and not (layer0_outputs(1561));
    layer1_outputs(1814) <= not(layer0_outputs(1920)) or (layer0_outputs(2486));
    layer1_outputs(1815) <= (layer0_outputs(614)) and not (layer0_outputs(1728));
    layer1_outputs(1816) <= not(layer0_outputs(869)) or (layer0_outputs(889));
    layer1_outputs(1817) <= not((layer0_outputs(1255)) or (layer0_outputs(248)));
    layer1_outputs(1818) <= not(layer0_outputs(515));
    layer1_outputs(1819) <= not(layer0_outputs(501));
    layer1_outputs(1820) <= not((layer0_outputs(1699)) and (layer0_outputs(1119)));
    layer1_outputs(1821) <= not((layer0_outputs(1)) or (layer0_outputs(2411)));
    layer1_outputs(1822) <= not(layer0_outputs(1434)) or (layer0_outputs(1912));
    layer1_outputs(1823) <= not((layer0_outputs(316)) and (layer0_outputs(2125)));
    layer1_outputs(1824) <= not(layer0_outputs(125));
    layer1_outputs(1825) <= not(layer0_outputs(2079));
    layer1_outputs(1826) <= (layer0_outputs(2125)) and (layer0_outputs(775));
    layer1_outputs(1827) <= (layer0_outputs(427)) and not (layer0_outputs(276));
    layer1_outputs(1828) <= layer0_outputs(2072);
    layer1_outputs(1829) <= (layer0_outputs(1140)) and not (layer0_outputs(1253));
    layer1_outputs(1830) <= layer0_outputs(1203);
    layer1_outputs(1831) <= (layer0_outputs(1029)) or (layer0_outputs(698));
    layer1_outputs(1832) <= not(layer0_outputs(1674)) or (layer0_outputs(761));
    layer1_outputs(1833) <= (layer0_outputs(99)) and not (layer0_outputs(644));
    layer1_outputs(1834) <= not(layer0_outputs(1381));
    layer1_outputs(1835) <= not(layer0_outputs(335));
    layer1_outputs(1836) <= not(layer0_outputs(816));
    layer1_outputs(1837) <= not(layer0_outputs(1184));
    layer1_outputs(1838) <= not((layer0_outputs(1871)) or (layer0_outputs(700)));
    layer1_outputs(1839) <= not(layer0_outputs(1618));
    layer1_outputs(1840) <= not((layer0_outputs(1665)) and (layer0_outputs(988)));
    layer1_outputs(1841) <= not(layer0_outputs(566)) or (layer0_outputs(982));
    layer1_outputs(1842) <= not((layer0_outputs(2426)) and (layer0_outputs(908)));
    layer1_outputs(1843) <= layer0_outputs(1508);
    layer1_outputs(1844) <= not(layer0_outputs(1268));
    layer1_outputs(1845) <= '1';
    layer1_outputs(1846) <= (layer0_outputs(8)) or (layer0_outputs(2339));
    layer1_outputs(1847) <= not(layer0_outputs(153));
    layer1_outputs(1848) <= layer0_outputs(2459);
    layer1_outputs(1849) <= not(layer0_outputs(1520)) or (layer0_outputs(2405));
    layer1_outputs(1850) <= (layer0_outputs(346)) and (layer0_outputs(424));
    layer1_outputs(1851) <= not((layer0_outputs(2516)) or (layer0_outputs(300)));
    layer1_outputs(1852) <= not(layer0_outputs(626)) or (layer0_outputs(264));
    layer1_outputs(1853) <= layer0_outputs(300);
    layer1_outputs(1854) <= (layer0_outputs(1778)) and not (layer0_outputs(456));
    layer1_outputs(1855) <= (layer0_outputs(2024)) and not (layer0_outputs(2030));
    layer1_outputs(1856) <= not(layer0_outputs(1065));
    layer1_outputs(1857) <= not(layer0_outputs(484)) or (layer0_outputs(216));
    layer1_outputs(1858) <= (layer0_outputs(221)) and not (layer0_outputs(148));
    layer1_outputs(1859) <= layer0_outputs(659);
    layer1_outputs(1860) <= not(layer0_outputs(1359)) or (layer0_outputs(2299));
    layer1_outputs(1861) <= (layer0_outputs(304)) and not (layer0_outputs(965));
    layer1_outputs(1862) <= not(layer0_outputs(425)) or (layer0_outputs(1555));
    layer1_outputs(1863) <= not(layer0_outputs(461));
    layer1_outputs(1864) <= (layer0_outputs(464)) or (layer0_outputs(2250));
    layer1_outputs(1865) <= not(layer0_outputs(685));
    layer1_outputs(1866) <= (layer0_outputs(2543)) and (layer0_outputs(1690));
    layer1_outputs(1867) <= layer0_outputs(986);
    layer1_outputs(1868) <= layer0_outputs(2530);
    layer1_outputs(1869) <= not(layer0_outputs(1730)) or (layer0_outputs(38));
    layer1_outputs(1870) <= (layer0_outputs(132)) or (layer0_outputs(182));
    layer1_outputs(1871) <= not(layer0_outputs(938)) or (layer0_outputs(613));
    layer1_outputs(1872) <= (layer0_outputs(1952)) and not (layer0_outputs(2060));
    layer1_outputs(1873) <= layer0_outputs(545);
    layer1_outputs(1874) <= '1';
    layer1_outputs(1875) <= not(layer0_outputs(858));
    layer1_outputs(1876) <= not(layer0_outputs(213)) or (layer0_outputs(2018));
    layer1_outputs(1877) <= '0';
    layer1_outputs(1878) <= layer0_outputs(1184);
    layer1_outputs(1879) <= layer0_outputs(1183);
    layer1_outputs(1880) <= not((layer0_outputs(1109)) or (layer0_outputs(2273)));
    layer1_outputs(1881) <= (layer0_outputs(2493)) and not (layer0_outputs(2009));
    layer1_outputs(1882) <= not((layer0_outputs(1589)) and (layer0_outputs(1243)));
    layer1_outputs(1883) <= (layer0_outputs(2472)) or (layer0_outputs(1834));
    layer1_outputs(1884) <= '0';
    layer1_outputs(1885) <= not((layer0_outputs(469)) or (layer0_outputs(2338)));
    layer1_outputs(1886) <= (layer0_outputs(1916)) and not (layer0_outputs(1570));
    layer1_outputs(1887) <= layer0_outputs(1876);
    layer1_outputs(1888) <= not(layer0_outputs(1351));
    layer1_outputs(1889) <= layer0_outputs(2546);
    layer1_outputs(1890) <= (layer0_outputs(1247)) and not (layer0_outputs(2376));
    layer1_outputs(1891) <= layer0_outputs(248);
    layer1_outputs(1892) <= (layer0_outputs(590)) or (layer0_outputs(1245));
    layer1_outputs(1893) <= not(layer0_outputs(143));
    layer1_outputs(1894) <= (layer0_outputs(679)) and not (layer0_outputs(1192));
    layer1_outputs(1895) <= not((layer0_outputs(2408)) and (layer0_outputs(907)));
    layer1_outputs(1896) <= layer0_outputs(1574);
    layer1_outputs(1897) <= (layer0_outputs(59)) and not (layer0_outputs(1176));
    layer1_outputs(1898) <= not(layer0_outputs(905));
    layer1_outputs(1899) <= not(layer0_outputs(1750));
    layer1_outputs(1900) <= not((layer0_outputs(852)) and (layer0_outputs(1041)));
    layer1_outputs(1901) <= layer0_outputs(245);
    layer1_outputs(1902) <= '0';
    layer1_outputs(1903) <= layer0_outputs(658);
    layer1_outputs(1904) <= layer0_outputs(741);
    layer1_outputs(1905) <= (layer0_outputs(749)) or (layer0_outputs(971));
    layer1_outputs(1906) <= not(layer0_outputs(2193));
    layer1_outputs(1907) <= not(layer0_outputs(2377)) or (layer0_outputs(1354));
    layer1_outputs(1908) <= (layer0_outputs(596)) or (layer0_outputs(2527));
    layer1_outputs(1909) <= (layer0_outputs(1007)) or (layer0_outputs(815));
    layer1_outputs(1910) <= layer0_outputs(1498);
    layer1_outputs(1911) <= not((layer0_outputs(1410)) and (layer0_outputs(1505)));
    layer1_outputs(1912) <= layer0_outputs(1250);
    layer1_outputs(1913) <= layer0_outputs(2251);
    layer1_outputs(1914) <= (layer0_outputs(2556)) and not (layer0_outputs(245));
    layer1_outputs(1915) <= not((layer0_outputs(378)) and (layer0_outputs(807)));
    layer1_outputs(1916) <= (layer0_outputs(1283)) and not (layer0_outputs(203));
    layer1_outputs(1917) <= not((layer0_outputs(1849)) or (layer0_outputs(1390)));
    layer1_outputs(1918) <= not(layer0_outputs(1010));
    layer1_outputs(1919) <= not(layer0_outputs(1772)) or (layer0_outputs(1700));
    layer1_outputs(1920) <= layer0_outputs(1898);
    layer1_outputs(1921) <= not((layer0_outputs(2471)) or (layer0_outputs(751)));
    layer1_outputs(1922) <= not((layer0_outputs(2270)) or (layer0_outputs(932)));
    layer1_outputs(1923) <= (layer0_outputs(1744)) or (layer0_outputs(193));
    layer1_outputs(1924) <= layer0_outputs(1981);
    layer1_outputs(1925) <= layer0_outputs(891);
    layer1_outputs(1926) <= layer0_outputs(2225);
    layer1_outputs(1927) <= not(layer0_outputs(1345));
    layer1_outputs(1928) <= not((layer0_outputs(2268)) and (layer0_outputs(672)));
    layer1_outputs(1929) <= (layer0_outputs(1057)) and not (layer0_outputs(1460));
    layer1_outputs(1930) <= not((layer0_outputs(318)) or (layer0_outputs(1666)));
    layer1_outputs(1931) <= layer0_outputs(889);
    layer1_outputs(1932) <= layer0_outputs(1449);
    layer1_outputs(1933) <= not(layer0_outputs(531));
    layer1_outputs(1934) <= layer0_outputs(238);
    layer1_outputs(1935) <= (layer0_outputs(2231)) and not (layer0_outputs(1657));
    layer1_outputs(1936) <= not(layer0_outputs(2534));
    layer1_outputs(1937) <= layer0_outputs(107);
    layer1_outputs(1938) <= '0';
    layer1_outputs(1939) <= not(layer0_outputs(1193));
    layer1_outputs(1940) <= (layer0_outputs(199)) and (layer0_outputs(439));
    layer1_outputs(1941) <= not(layer0_outputs(255));
    layer1_outputs(1942) <= (layer0_outputs(2038)) and not (layer0_outputs(1617));
    layer1_outputs(1943) <= not(layer0_outputs(508));
    layer1_outputs(1944) <= layer0_outputs(120);
    layer1_outputs(1945) <= (layer0_outputs(535)) or (layer0_outputs(2394));
    layer1_outputs(1946) <= not(layer0_outputs(2554));
    layer1_outputs(1947) <= not(layer0_outputs(217)) or (layer0_outputs(1911));
    layer1_outputs(1948) <= not((layer0_outputs(1652)) or (layer0_outputs(2306)));
    layer1_outputs(1949) <= (layer0_outputs(780)) and not (layer0_outputs(842));
    layer1_outputs(1950) <= not((layer0_outputs(1997)) and (layer0_outputs(2420)));
    layer1_outputs(1951) <= not((layer0_outputs(787)) and (layer0_outputs(1947)));
    layer1_outputs(1952) <= not((layer0_outputs(1331)) xor (layer0_outputs(1149)));
    layer1_outputs(1953) <= (layer0_outputs(1355)) and (layer0_outputs(2438));
    layer1_outputs(1954) <= not((layer0_outputs(2)) or (layer0_outputs(532)));
    layer1_outputs(1955) <= not(layer0_outputs(438));
    layer1_outputs(1956) <= (layer0_outputs(692)) and not (layer0_outputs(1264));
    layer1_outputs(1957) <= not(layer0_outputs(478)) or (layer0_outputs(1541));
    layer1_outputs(1958) <= layer0_outputs(917);
    layer1_outputs(1959) <= (layer0_outputs(2498)) or (layer0_outputs(214));
    layer1_outputs(1960) <= not(layer0_outputs(561));
    layer1_outputs(1961) <= layer0_outputs(490);
    layer1_outputs(1962) <= not(layer0_outputs(1407));
    layer1_outputs(1963) <= layer0_outputs(1433);
    layer1_outputs(1964) <= layer0_outputs(1301);
    layer1_outputs(1965) <= not(layer0_outputs(2466)) or (layer0_outputs(763));
    layer1_outputs(1966) <= not(layer0_outputs(490));
    layer1_outputs(1967) <= layer0_outputs(2238);
    layer1_outputs(1968) <= not(layer0_outputs(1065));
    layer1_outputs(1969) <= not(layer0_outputs(2403));
    layer1_outputs(1970) <= layer0_outputs(214);
    layer1_outputs(1971) <= not(layer0_outputs(1737));
    layer1_outputs(1972) <= not(layer0_outputs(1909)) or (layer0_outputs(1248));
    layer1_outputs(1973) <= not(layer0_outputs(2311));
    layer1_outputs(1974) <= not((layer0_outputs(2353)) or (layer0_outputs(5)));
    layer1_outputs(1975) <= layer0_outputs(1765);
    layer1_outputs(1976) <= '0';
    layer1_outputs(1977) <= (layer0_outputs(2227)) and not (layer0_outputs(2035));
    layer1_outputs(1978) <= not(layer0_outputs(2532));
    layer1_outputs(1979) <= not((layer0_outputs(2255)) and (layer0_outputs(335)));
    layer1_outputs(1980) <= (layer0_outputs(509)) and (layer0_outputs(1155));
    layer1_outputs(1981) <= layer0_outputs(1780);
    layer1_outputs(1982) <= (layer0_outputs(500)) and (layer0_outputs(2303));
    layer1_outputs(1983) <= not(layer0_outputs(1532)) or (layer0_outputs(252));
    layer1_outputs(1984) <= (layer0_outputs(952)) and not (layer0_outputs(628));
    layer1_outputs(1985) <= (layer0_outputs(1991)) or (layer0_outputs(377));
    layer1_outputs(1986) <= not((layer0_outputs(51)) and (layer0_outputs(1929)));
    layer1_outputs(1987) <= (layer0_outputs(965)) and not (layer0_outputs(1429));
    layer1_outputs(1988) <= (layer0_outputs(1804)) xor (layer0_outputs(1305));
    layer1_outputs(1989) <= layer0_outputs(2511);
    layer1_outputs(1990) <= '1';
    layer1_outputs(1991) <= not((layer0_outputs(314)) and (layer0_outputs(197)));
    layer1_outputs(1992) <= not(layer0_outputs(2114)) or (layer0_outputs(1820));
    layer1_outputs(1993) <= layer0_outputs(1711);
    layer1_outputs(1994) <= not(layer0_outputs(52)) or (layer0_outputs(1837));
    layer1_outputs(1995) <= (layer0_outputs(1317)) and (layer0_outputs(1655));
    layer1_outputs(1996) <= layer0_outputs(1222);
    layer1_outputs(1997) <= layer0_outputs(320);
    layer1_outputs(1998) <= layer0_outputs(1906);
    layer1_outputs(1999) <= (layer0_outputs(1421)) xor (layer0_outputs(1901));
    layer1_outputs(2000) <= layer0_outputs(2433);
    layer1_outputs(2001) <= not(layer0_outputs(2417));
    layer1_outputs(2002) <= layer0_outputs(329);
    layer1_outputs(2003) <= not(layer0_outputs(2189));
    layer1_outputs(2004) <= (layer0_outputs(2352)) and not (layer0_outputs(1954));
    layer1_outputs(2005) <= not(layer0_outputs(2362));
    layer1_outputs(2006) <= '0';
    layer1_outputs(2007) <= not(layer0_outputs(1403));
    layer1_outputs(2008) <= (layer0_outputs(1560)) and (layer0_outputs(30));
    layer1_outputs(2009) <= not(layer0_outputs(498));
    layer1_outputs(2010) <= not((layer0_outputs(2452)) or (layer0_outputs(1232)));
    layer1_outputs(2011) <= (layer0_outputs(461)) and (layer0_outputs(2312));
    layer1_outputs(2012) <= not(layer0_outputs(1000)) or (layer0_outputs(824));
    layer1_outputs(2013) <= not((layer0_outputs(2001)) and (layer0_outputs(116)));
    layer1_outputs(2014) <= layer0_outputs(2346);
    layer1_outputs(2015) <= not(layer0_outputs(2067)) or (layer0_outputs(738));
    layer1_outputs(2016) <= not(layer0_outputs(1534));
    layer1_outputs(2017) <= (layer0_outputs(896)) or (layer0_outputs(1471));
    layer1_outputs(2018) <= not(layer0_outputs(462)) or (layer0_outputs(73));
    layer1_outputs(2019) <= not((layer0_outputs(941)) and (layer0_outputs(1286)));
    layer1_outputs(2020) <= layer0_outputs(1552);
    layer1_outputs(2021) <= not(layer0_outputs(1680));
    layer1_outputs(2022) <= layer0_outputs(1370);
    layer1_outputs(2023) <= (layer0_outputs(1430)) and not (layer0_outputs(1410));
    layer1_outputs(2024) <= layer0_outputs(1759);
    layer1_outputs(2025) <= not(layer0_outputs(1339));
    layer1_outputs(2026) <= layer0_outputs(2090);
    layer1_outputs(2027) <= '0';
    layer1_outputs(2028) <= not(layer0_outputs(1659));
    layer1_outputs(2029) <= not((layer0_outputs(1820)) xor (layer0_outputs(95)));
    layer1_outputs(2030) <= not((layer0_outputs(1030)) xor (layer0_outputs(736)));
    layer1_outputs(2031) <= not(layer0_outputs(2095));
    layer1_outputs(2032) <= not(layer0_outputs(1554));
    layer1_outputs(2033) <= layer0_outputs(2482);
    layer1_outputs(2034) <= layer0_outputs(2404);
    layer1_outputs(2035) <= not(layer0_outputs(1394));
    layer1_outputs(2036) <= '0';
    layer1_outputs(2037) <= layer0_outputs(1211);
    layer1_outputs(2038) <= (layer0_outputs(709)) xor (layer0_outputs(2117));
    layer1_outputs(2039) <= layer0_outputs(579);
    layer1_outputs(2040) <= not((layer0_outputs(272)) and (layer0_outputs(639)));
    layer1_outputs(2041) <= not((layer0_outputs(2476)) or (layer0_outputs(2484)));
    layer1_outputs(2042) <= (layer0_outputs(296)) and not (layer0_outputs(448));
    layer1_outputs(2043) <= (layer0_outputs(1860)) or (layer0_outputs(2269));
    layer1_outputs(2044) <= layer0_outputs(237);
    layer1_outputs(2045) <= not(layer0_outputs(749));
    layer1_outputs(2046) <= layer0_outputs(180);
    layer1_outputs(2047) <= not(layer0_outputs(1635));
    layer1_outputs(2048) <= '1';
    layer1_outputs(2049) <= (layer0_outputs(2148)) and not (layer0_outputs(737));
    layer1_outputs(2050) <= layer0_outputs(592);
    layer1_outputs(2051) <= not(layer0_outputs(2049));
    layer1_outputs(2052) <= layer0_outputs(1725);
    layer1_outputs(2053) <= (layer0_outputs(1616)) and not (layer0_outputs(1844));
    layer1_outputs(2054) <= layer0_outputs(2455);
    layer1_outputs(2055) <= not(layer0_outputs(557));
    layer1_outputs(2056) <= not(layer0_outputs(1847)) or (layer0_outputs(857));
    layer1_outputs(2057) <= (layer0_outputs(2022)) and not (layer0_outputs(1899));
    layer1_outputs(2058) <= '0';
    layer1_outputs(2059) <= not(layer0_outputs(2028)) or (layer0_outputs(1234));
    layer1_outputs(2060) <= not(layer0_outputs(2097)) or (layer0_outputs(583));
    layer1_outputs(2061) <= layer0_outputs(2338);
    layer1_outputs(2062) <= not(layer0_outputs(2279)) or (layer0_outputs(2531));
    layer1_outputs(2063) <= layer0_outputs(1004);
    layer1_outputs(2064) <= not((layer0_outputs(466)) xor (layer0_outputs(1716)));
    layer1_outputs(2065) <= not(layer0_outputs(2337));
    layer1_outputs(2066) <= not((layer0_outputs(727)) and (layer0_outputs(1696)));
    layer1_outputs(2067) <= (layer0_outputs(194)) and not (layer0_outputs(1122));
    layer1_outputs(2068) <= not((layer0_outputs(387)) or (layer0_outputs(2025)));
    layer1_outputs(2069) <= layer0_outputs(1437);
    layer1_outputs(2070) <= not((layer0_outputs(2366)) or (layer0_outputs(1078)));
    layer1_outputs(2071) <= (layer0_outputs(1273)) and (layer0_outputs(2004));
    layer1_outputs(2072) <= not(layer0_outputs(1971)) or (layer0_outputs(411));
    layer1_outputs(2073) <= (layer0_outputs(529)) and not (layer0_outputs(823));
    layer1_outputs(2074) <= (layer0_outputs(360)) and (layer0_outputs(2252));
    layer1_outputs(2075) <= not(layer0_outputs(1361));
    layer1_outputs(2076) <= not(layer0_outputs(1148)) or (layer0_outputs(2325));
    layer1_outputs(2077) <= (layer0_outputs(700)) and not (layer0_outputs(201));
    layer1_outputs(2078) <= (layer0_outputs(526)) and (layer0_outputs(151));
    layer1_outputs(2079) <= '0';
    layer1_outputs(2080) <= layer0_outputs(354);
    layer1_outputs(2081) <= (layer0_outputs(1646)) and not (layer0_outputs(916));
    layer1_outputs(2082) <= (layer0_outputs(324)) or (layer0_outputs(406));
    layer1_outputs(2083) <= not(layer0_outputs(688)) or (layer0_outputs(1689));
    layer1_outputs(2084) <= not(layer0_outputs(1841));
    layer1_outputs(2085) <= not((layer0_outputs(1986)) and (layer0_outputs(990)));
    layer1_outputs(2086) <= not(layer0_outputs(1675));
    layer1_outputs(2087) <= not((layer0_outputs(85)) or (layer0_outputs(571)));
    layer1_outputs(2088) <= not(layer0_outputs(722));
    layer1_outputs(2089) <= not(layer0_outputs(1457));
    layer1_outputs(2090) <= (layer0_outputs(134)) and not (layer0_outputs(2529));
    layer1_outputs(2091) <= layer0_outputs(1829);
    layer1_outputs(2092) <= layer0_outputs(84);
    layer1_outputs(2093) <= (layer0_outputs(2237)) and (layer0_outputs(2354));
    layer1_outputs(2094) <= not((layer0_outputs(732)) or (layer0_outputs(166)));
    layer1_outputs(2095) <= (layer0_outputs(385)) and (layer0_outputs(1502));
    layer1_outputs(2096) <= not((layer0_outputs(964)) or (layer0_outputs(2234)));
    layer1_outputs(2097) <= not(layer0_outputs(1368));
    layer1_outputs(2098) <= not(layer0_outputs(2173)) or (layer0_outputs(2086));
    layer1_outputs(2099) <= not((layer0_outputs(1724)) xor (layer0_outputs(1307)));
    layer1_outputs(2100) <= not(layer0_outputs(2501));
    layer1_outputs(2101) <= layer0_outputs(2039);
    layer1_outputs(2102) <= (layer0_outputs(1907)) and not (layer0_outputs(1530));
    layer1_outputs(2103) <= not(layer0_outputs(537));
    layer1_outputs(2104) <= not(layer0_outputs(1690)) or (layer0_outputs(766));
    layer1_outputs(2105) <= (layer0_outputs(2461)) or (layer0_outputs(1939));
    layer1_outputs(2106) <= layer0_outputs(1807);
    layer1_outputs(2107) <= (layer0_outputs(1835)) and not (layer0_outputs(1251));
    layer1_outputs(2108) <= not((layer0_outputs(2137)) or (layer0_outputs(1052)));
    layer1_outputs(2109) <= layer0_outputs(610);
    layer1_outputs(2110) <= (layer0_outputs(695)) and not (layer0_outputs(2250));
    layer1_outputs(2111) <= not((layer0_outputs(397)) or (layer0_outputs(228)));
    layer1_outputs(2112) <= not(layer0_outputs(2492));
    layer1_outputs(2113) <= not(layer0_outputs(560));
    layer1_outputs(2114) <= not(layer0_outputs(2494));
    layer1_outputs(2115) <= not(layer0_outputs(1911));
    layer1_outputs(2116) <= layer0_outputs(820);
    layer1_outputs(2117) <= layer0_outputs(2505);
    layer1_outputs(2118) <= layer0_outputs(1637);
    layer1_outputs(2119) <= (layer0_outputs(2075)) and not (layer0_outputs(937));
    layer1_outputs(2120) <= layer0_outputs(455);
    layer1_outputs(2121) <= (layer0_outputs(1467)) and (layer0_outputs(2525));
    layer1_outputs(2122) <= not(layer0_outputs(997));
    layer1_outputs(2123) <= not(layer0_outputs(1638));
    layer1_outputs(2124) <= (layer0_outputs(2082)) or (layer0_outputs(2367));
    layer1_outputs(2125) <= layer0_outputs(1900);
    layer1_outputs(2126) <= layer0_outputs(1559);
    layer1_outputs(2127) <= not(layer0_outputs(130));
    layer1_outputs(2128) <= '0';
    layer1_outputs(2129) <= not((layer0_outputs(598)) and (layer0_outputs(1095)));
    layer1_outputs(2130) <= layer0_outputs(729);
    layer1_outputs(2131) <= (layer0_outputs(1963)) and not (layer0_outputs(2180));
    layer1_outputs(2132) <= (layer0_outputs(450)) and (layer0_outputs(2387));
    layer1_outputs(2133) <= '1';
    layer1_outputs(2134) <= not(layer0_outputs(2175));
    layer1_outputs(2135) <= not(layer0_outputs(491));
    layer1_outputs(2136) <= layer0_outputs(1292);
    layer1_outputs(2137) <= (layer0_outputs(1584)) or (layer0_outputs(1615));
    layer1_outputs(2138) <= (layer0_outputs(1808)) and (layer0_outputs(1230));
    layer1_outputs(2139) <= not(layer0_outputs(1321)) or (layer0_outputs(1959));
    layer1_outputs(2140) <= layer0_outputs(441);
    layer1_outputs(2141) <= not(layer0_outputs(2510));
    layer1_outputs(2142) <= '0';
    layer1_outputs(2143) <= not(layer0_outputs(1009)) or (layer0_outputs(1892));
    layer1_outputs(2144) <= (layer0_outputs(1357)) and not (layer0_outputs(2549));
    layer1_outputs(2145) <= (layer0_outputs(551)) and not (layer0_outputs(1503));
    layer1_outputs(2146) <= layer0_outputs(291);
    layer1_outputs(2147) <= not(layer0_outputs(2135));
    layer1_outputs(2148) <= not(layer0_outputs(2341)) or (layer0_outputs(1366));
    layer1_outputs(2149) <= layer0_outputs(2043);
    layer1_outputs(2150) <= not(layer0_outputs(607));
    layer1_outputs(2151) <= not((layer0_outputs(1431)) or (layer0_outputs(1156)));
    layer1_outputs(2152) <= (layer0_outputs(686)) or (layer0_outputs(742));
    layer1_outputs(2153) <= not(layer0_outputs(239));
    layer1_outputs(2154) <= not(layer0_outputs(1879));
    layer1_outputs(2155) <= not((layer0_outputs(1488)) xor (layer0_outputs(645)));
    layer1_outputs(2156) <= not(layer0_outputs(697)) or (layer0_outputs(1754));
    layer1_outputs(2157) <= not(layer0_outputs(1537)) or (layer0_outputs(2429));
    layer1_outputs(2158) <= not(layer0_outputs(1852));
    layer1_outputs(2159) <= (layer0_outputs(2149)) and not (layer0_outputs(1445));
    layer1_outputs(2160) <= not(layer0_outputs(867)) or (layer0_outputs(1894));
    layer1_outputs(2161) <= layer0_outputs(790);
    layer1_outputs(2162) <= not((layer0_outputs(1152)) xor (layer0_outputs(1749)));
    layer1_outputs(2163) <= not((layer0_outputs(1649)) or (layer0_outputs(989)));
    layer1_outputs(2164) <= not(layer0_outputs(2308));
    layer1_outputs(2165) <= layer0_outputs(892);
    layer1_outputs(2166) <= layer0_outputs(460);
    layer1_outputs(2167) <= not(layer0_outputs(2364));
    layer1_outputs(2168) <= not(layer0_outputs(194));
    layer1_outputs(2169) <= layer0_outputs(1887);
    layer1_outputs(2170) <= (layer0_outputs(1880)) and (layer0_outputs(595));
    layer1_outputs(2171) <= not(layer0_outputs(1584)) or (layer0_outputs(573));
    layer1_outputs(2172) <= not(layer0_outputs(2138));
    layer1_outputs(2173) <= not((layer0_outputs(1710)) or (layer0_outputs(960)));
    layer1_outputs(2174) <= not((layer0_outputs(372)) or (layer0_outputs(2240)));
    layer1_outputs(2175) <= not((layer0_outputs(2283)) or (layer0_outputs(913)));
    layer1_outputs(2176) <= layer0_outputs(27);
    layer1_outputs(2177) <= (layer0_outputs(336)) or (layer0_outputs(585));
    layer1_outputs(2178) <= layer0_outputs(63);
    layer1_outputs(2179) <= not(layer0_outputs(1340));
    layer1_outputs(2180) <= not(layer0_outputs(477)) or (layer0_outputs(758));
    layer1_outputs(2181) <= layer0_outputs(1945);
    layer1_outputs(2182) <= not(layer0_outputs(1740)) or (layer0_outputs(977));
    layer1_outputs(2183) <= not(layer0_outputs(1544)) or (layer0_outputs(1471));
    layer1_outputs(2184) <= not(layer0_outputs(2105)) or (layer0_outputs(1602));
    layer1_outputs(2185) <= not(layer0_outputs(1409));
    layer1_outputs(2186) <= (layer0_outputs(123)) and not (layer0_outputs(2176));
    layer1_outputs(2187) <= (layer0_outputs(518)) and not (layer0_outputs(206));
    layer1_outputs(2188) <= (layer0_outputs(1985)) and not (layer0_outputs(1937));
    layer1_outputs(2189) <= layer0_outputs(2196);
    layer1_outputs(2190) <= (layer0_outputs(1241)) and (layer0_outputs(2132));
    layer1_outputs(2191) <= layer0_outputs(2500);
    layer1_outputs(2192) <= not(layer0_outputs(1921)) or (layer0_outputs(2171));
    layer1_outputs(2193) <= (layer0_outputs(1598)) and not (layer0_outputs(1468));
    layer1_outputs(2194) <= not(layer0_outputs(1435)) or (layer0_outputs(1373));
    layer1_outputs(2195) <= not(layer0_outputs(2438));
    layer1_outputs(2196) <= not(layer0_outputs(1237)) or (layer0_outputs(1323));
    layer1_outputs(2197) <= not((layer0_outputs(572)) and (layer0_outputs(1308)));
    layer1_outputs(2198) <= not((layer0_outputs(1140)) or (layer0_outputs(2485)));
    layer1_outputs(2199) <= (layer0_outputs(1047)) and not (layer0_outputs(18));
    layer1_outputs(2200) <= '1';
    layer1_outputs(2201) <= not(layer0_outputs(985));
    layer1_outputs(2202) <= not(layer0_outputs(1732));
    layer1_outputs(2203) <= layer0_outputs(110);
    layer1_outputs(2204) <= (layer0_outputs(1221)) xor (layer0_outputs(432));
    layer1_outputs(2205) <= not((layer0_outputs(1504)) and (layer0_outputs(1076)));
    layer1_outputs(2206) <= not(layer0_outputs(579)) or (layer0_outputs(1142));
    layer1_outputs(2207) <= (layer0_outputs(11)) or (layer0_outputs(69));
    layer1_outputs(2208) <= not(layer0_outputs(400)) or (layer0_outputs(986));
    layer1_outputs(2209) <= not(layer0_outputs(1511)) or (layer0_outputs(2328));
    layer1_outputs(2210) <= '0';
    layer1_outputs(2211) <= layer0_outputs(20);
    layer1_outputs(2212) <= not((layer0_outputs(899)) and (layer0_outputs(2033)));
    layer1_outputs(2213) <= not(layer0_outputs(1333));
    layer1_outputs(2214) <= not((layer0_outputs(1670)) or (layer0_outputs(1045)));
    layer1_outputs(2215) <= '1';
    layer1_outputs(2216) <= not(layer0_outputs(1299));
    layer1_outputs(2217) <= not(layer0_outputs(714));
    layer1_outputs(2218) <= not(layer0_outputs(468));
    layer1_outputs(2219) <= (layer0_outputs(1466)) and not (layer0_outputs(402));
    layer1_outputs(2220) <= not(layer0_outputs(1734)) or (layer0_outputs(1885));
    layer1_outputs(2221) <= not(layer0_outputs(1130));
    layer1_outputs(2222) <= not((layer0_outputs(952)) and (layer0_outputs(1079)));
    layer1_outputs(2223) <= (layer0_outputs(2478)) and not (layer0_outputs(1742));
    layer1_outputs(2224) <= (layer0_outputs(211)) and (layer0_outputs(2219));
    layer1_outputs(2225) <= not(layer0_outputs(2344));
    layer1_outputs(2226) <= not((layer0_outputs(704)) or (layer0_outputs(894)));
    layer1_outputs(2227) <= layer0_outputs(919);
    layer1_outputs(2228) <= not((layer0_outputs(1723)) or (layer0_outputs(2019)));
    layer1_outputs(2229) <= layer0_outputs(1669);
    layer1_outputs(2230) <= (layer0_outputs(599)) and not (layer0_outputs(871));
    layer1_outputs(2231) <= not(layer0_outputs(108));
    layer1_outputs(2232) <= (layer0_outputs(694)) and (layer0_outputs(1126));
    layer1_outputs(2233) <= not((layer0_outputs(1332)) xor (layer0_outputs(211)));
    layer1_outputs(2234) <= not(layer0_outputs(2039));
    layer1_outputs(2235) <= not(layer0_outputs(298)) or (layer0_outputs(1201));
    layer1_outputs(2236) <= not((layer0_outputs(599)) and (layer0_outputs(2017)));
    layer1_outputs(2237) <= (layer0_outputs(1013)) and (layer0_outputs(1019));
    layer1_outputs(2238) <= not(layer0_outputs(1987));
    layer1_outputs(2239) <= layer0_outputs(900);
    layer1_outputs(2240) <= not(layer0_outputs(2047)) or (layer0_outputs(482));
    layer1_outputs(2241) <= not(layer0_outputs(1673)) or (layer0_outputs(1341));
    layer1_outputs(2242) <= not(layer0_outputs(877));
    layer1_outputs(2243) <= layer0_outputs(1941);
    layer1_outputs(2244) <= (layer0_outputs(1643)) or (layer0_outputs(219));
    layer1_outputs(2245) <= (layer0_outputs(2271)) or (layer0_outputs(1715));
    layer1_outputs(2246) <= (layer0_outputs(1150)) and not (layer0_outputs(790));
    layer1_outputs(2247) <= not(layer0_outputs(1181));
    layer1_outputs(2248) <= (layer0_outputs(1869)) and (layer0_outputs(1658));
    layer1_outputs(2249) <= not(layer0_outputs(1433));
    layer1_outputs(2250) <= not(layer0_outputs(1483)) or (layer0_outputs(142));
    layer1_outputs(2251) <= not(layer0_outputs(1496));
    layer1_outputs(2252) <= (layer0_outputs(1250)) and not (layer0_outputs(2418));
    layer1_outputs(2253) <= layer0_outputs(1939);
    layer1_outputs(2254) <= not(layer0_outputs(1039));
    layer1_outputs(2255) <= layer0_outputs(605);
    layer1_outputs(2256) <= '0';
    layer1_outputs(2257) <= not((layer0_outputs(507)) xor (layer0_outputs(563)));
    layer1_outputs(2258) <= layer0_outputs(792);
    layer1_outputs(2259) <= not(layer0_outputs(1516)) or (layer0_outputs(1316));
    layer1_outputs(2260) <= not((layer0_outputs(376)) and (layer0_outputs(2496)));
    layer1_outputs(2261) <= (layer0_outputs(2412)) and not (layer0_outputs(928));
    layer1_outputs(2262) <= not((layer0_outputs(2127)) and (layer0_outputs(270)));
    layer1_outputs(2263) <= not((layer0_outputs(1905)) and (layer0_outputs(468)));
    layer1_outputs(2264) <= layer0_outputs(1205);
    layer1_outputs(2265) <= not(layer0_outputs(1985));
    layer1_outputs(2266) <= not(layer0_outputs(1588));
    layer1_outputs(2267) <= (layer0_outputs(20)) and (layer0_outputs(463));
    layer1_outputs(2268) <= layer0_outputs(1710);
    layer1_outputs(2269) <= not(layer0_outputs(371));
    layer1_outputs(2270) <= layer0_outputs(155);
    layer1_outputs(2271) <= not((layer0_outputs(895)) or (layer0_outputs(1172)));
    layer1_outputs(2272) <= '1';
    layer1_outputs(2273) <= (layer0_outputs(1699)) and (layer0_outputs(643));
    layer1_outputs(2274) <= not(layer0_outputs(1059)) or (layer0_outputs(2530));
    layer1_outputs(2275) <= not(layer0_outputs(1412));
    layer1_outputs(2276) <= (layer0_outputs(1763)) xor (layer0_outputs(1826));
    layer1_outputs(2277) <= not(layer0_outputs(241)) or (layer0_outputs(1246));
    layer1_outputs(2278) <= not(layer0_outputs(305));
    layer1_outputs(2279) <= layer0_outputs(1228);
    layer1_outputs(2280) <= (layer0_outputs(310)) and not (layer0_outputs(24));
    layer1_outputs(2281) <= '1';
    layer1_outputs(2282) <= layer0_outputs(732);
    layer1_outputs(2283) <= (layer0_outputs(2339)) and not (layer0_outputs(2557));
    layer1_outputs(2284) <= not((layer0_outputs(1671)) or (layer0_outputs(88)));
    layer1_outputs(2285) <= not((layer0_outputs(575)) xor (layer0_outputs(844)));
    layer1_outputs(2286) <= not((layer0_outputs(640)) or (layer0_outputs(2464)));
    layer1_outputs(2287) <= not(layer0_outputs(1266)) or (layer0_outputs(690));
    layer1_outputs(2288) <= (layer0_outputs(586)) or (layer0_outputs(697));
    layer1_outputs(2289) <= layer0_outputs(848);
    layer1_outputs(2290) <= (layer0_outputs(1175)) or (layer0_outputs(2351));
    layer1_outputs(2291) <= not((layer0_outputs(1016)) or (layer0_outputs(411)));
    layer1_outputs(2292) <= layer0_outputs(2528);
    layer1_outputs(2293) <= not(layer0_outputs(1923));
    layer1_outputs(2294) <= not((layer0_outputs(678)) or (layer0_outputs(1613)));
    layer1_outputs(2295) <= layer0_outputs(486);
    layer1_outputs(2296) <= layer0_outputs(1773);
    layer1_outputs(2297) <= layer0_outputs(2103);
    layer1_outputs(2298) <= (layer0_outputs(2050)) xor (layer0_outputs(754));
    layer1_outputs(2299) <= not((layer0_outputs(2107)) or (layer0_outputs(2297)));
    layer1_outputs(2300) <= (layer0_outputs(2239)) xor (layer0_outputs(271));
    layer1_outputs(2301) <= layer0_outputs(765);
    layer1_outputs(2302) <= layer0_outputs(2218);
    layer1_outputs(2303) <= not(layer0_outputs(546)) or (layer0_outputs(360));
    layer1_outputs(2304) <= not(layer0_outputs(1656));
    layer1_outputs(2305) <= (layer0_outputs(1762)) and not (layer0_outputs(2313));
    layer1_outputs(2306) <= not(layer0_outputs(827));
    layer1_outputs(2307) <= (layer0_outputs(2264)) and (layer0_outputs(166));
    layer1_outputs(2308) <= not(layer0_outputs(21)) or (layer0_outputs(73));
    layer1_outputs(2309) <= not((layer0_outputs(1738)) and (layer0_outputs(64)));
    layer1_outputs(2310) <= not((layer0_outputs(2274)) and (layer0_outputs(102)));
    layer1_outputs(2311) <= not(layer0_outputs(831));
    layer1_outputs(2312) <= layer0_outputs(1704);
    layer1_outputs(2313) <= (layer0_outputs(578)) or (layer0_outputs(1388));
    layer1_outputs(2314) <= not(layer0_outputs(1136)) or (layer0_outputs(1346));
    layer1_outputs(2315) <= not(layer0_outputs(1188));
    layer1_outputs(2316) <= layer0_outputs(805);
    layer1_outputs(2317) <= (layer0_outputs(2454)) and not (layer0_outputs(2365));
    layer1_outputs(2318) <= not((layer0_outputs(2357)) or (layer0_outputs(177)));
    layer1_outputs(2319) <= not((layer0_outputs(726)) and (layer0_outputs(1706)));
    layer1_outputs(2320) <= '0';
    layer1_outputs(2321) <= layer0_outputs(2491);
    layer1_outputs(2322) <= (layer0_outputs(1960)) and not (layer0_outputs(162));
    layer1_outputs(2323) <= not(layer0_outputs(2214));
    layer1_outputs(2324) <= layer0_outputs(1127);
    layer1_outputs(2325) <= not((layer0_outputs(657)) or (layer0_outputs(1755)));
    layer1_outputs(2326) <= (layer0_outputs(1571)) and (layer0_outputs(1707));
    layer1_outputs(2327) <= (layer0_outputs(1709)) and (layer0_outputs(721));
    layer1_outputs(2328) <= not(layer0_outputs(973)) or (layer0_outputs(1730));
    layer1_outputs(2329) <= (layer0_outputs(587)) and not (layer0_outputs(145));
    layer1_outputs(2330) <= layer0_outputs(938);
    layer1_outputs(2331) <= (layer0_outputs(1465)) and not (layer0_outputs(1458));
    layer1_outputs(2332) <= (layer0_outputs(2419)) and not (layer0_outputs(1582));
    layer1_outputs(2333) <= not(layer0_outputs(124)) or (layer0_outputs(1973));
    layer1_outputs(2334) <= '1';
    layer1_outputs(2335) <= not(layer0_outputs(758));
    layer1_outputs(2336) <= not(layer0_outputs(942)) or (layer0_outputs(1515));
    layer1_outputs(2337) <= not(layer0_outputs(973));
    layer1_outputs(2338) <= layer0_outputs(852);
    layer1_outputs(2339) <= not(layer0_outputs(1654)) or (layer0_outputs(901));
    layer1_outputs(2340) <= not(layer0_outputs(2257));
    layer1_outputs(2341) <= layer0_outputs(578);
    layer1_outputs(2342) <= not(layer0_outputs(1332)) or (layer0_outputs(1118));
    layer1_outputs(2343) <= layer0_outputs(111);
    layer1_outputs(2344) <= layer0_outputs(2105);
    layer1_outputs(2345) <= layer0_outputs(782);
    layer1_outputs(2346) <= layer0_outputs(1072);
    layer1_outputs(2347) <= not((layer0_outputs(2034)) or (layer0_outputs(2124)));
    layer1_outputs(2348) <= layer0_outputs(2064);
    layer1_outputs(2349) <= layer0_outputs(1086);
    layer1_outputs(2350) <= layer0_outputs(976);
    layer1_outputs(2351) <= (layer0_outputs(1228)) and (layer0_outputs(41));
    layer1_outputs(2352) <= (layer0_outputs(1247)) and not (layer0_outputs(1758));
    layer1_outputs(2353) <= not(layer0_outputs(1269));
    layer1_outputs(2354) <= not((layer0_outputs(1951)) and (layer0_outputs(2202)));
    layer1_outputs(2355) <= not(layer0_outputs(303)) or (layer0_outputs(1891));
    layer1_outputs(2356) <= not(layer0_outputs(1550)) or (layer0_outputs(1701));
    layer1_outputs(2357) <= not(layer0_outputs(346)) or (layer0_outputs(884));
    layer1_outputs(2358) <= (layer0_outputs(268)) and (layer0_outputs(662));
    layer1_outputs(2359) <= (layer0_outputs(1430)) xor (layer0_outputs(1112));
    layer1_outputs(2360) <= not(layer0_outputs(1385)) or (layer0_outputs(1227));
    layer1_outputs(2361) <= not(layer0_outputs(123));
    layer1_outputs(2362) <= layer0_outputs(1930);
    layer1_outputs(2363) <= (layer0_outputs(2209)) and not (layer0_outputs(553));
    layer1_outputs(2364) <= not(layer0_outputs(393));
    layer1_outputs(2365) <= not(layer0_outputs(1878));
    layer1_outputs(2366) <= not(layer0_outputs(863));
    layer1_outputs(2367) <= not(layer0_outputs(2535));
    layer1_outputs(2368) <= not(layer0_outputs(268)) or (layer0_outputs(380));
    layer1_outputs(2369) <= (layer0_outputs(2219)) and (layer0_outputs(1097));
    layer1_outputs(2370) <= layer0_outputs(363);
    layer1_outputs(2371) <= not((layer0_outputs(228)) and (layer0_outputs(259)));
    layer1_outputs(2372) <= not((layer0_outputs(1803)) or (layer0_outputs(2284)));
    layer1_outputs(2373) <= not(layer0_outputs(333)) or (layer0_outputs(1089));
    layer1_outputs(2374) <= not(layer0_outputs(249));
    layer1_outputs(2375) <= (layer0_outputs(1159)) and not (layer0_outputs(90));
    layer1_outputs(2376) <= (layer0_outputs(2449)) or (layer0_outputs(1784));
    layer1_outputs(2377) <= '0';
    layer1_outputs(2378) <= layer0_outputs(1528);
    layer1_outputs(2379) <= (layer0_outputs(325)) xor (layer0_outputs(467));
    layer1_outputs(2380) <= not(layer0_outputs(868));
    layer1_outputs(2381) <= '1';
    layer1_outputs(2382) <= layer0_outputs(1150);
    layer1_outputs(2383) <= not(layer0_outputs(188));
    layer1_outputs(2384) <= not((layer0_outputs(850)) or (layer0_outputs(671)));
    layer1_outputs(2385) <= not(layer0_outputs(2418));
    layer1_outputs(2386) <= '0';
    layer1_outputs(2387) <= not((layer0_outputs(630)) and (layer0_outputs(1708)));
    layer1_outputs(2388) <= '1';
    layer1_outputs(2389) <= (layer0_outputs(1950)) or (layer0_outputs(68));
    layer1_outputs(2390) <= not(layer0_outputs(56)) or (layer0_outputs(1043));
    layer1_outputs(2391) <= (layer0_outputs(719)) or (layer0_outputs(250));
    layer1_outputs(2392) <= (layer0_outputs(2455)) and (layer0_outputs(1302));
    layer1_outputs(2393) <= not(layer0_outputs(746)) or (layer0_outputs(2330));
    layer1_outputs(2394) <= '1';
    layer1_outputs(2395) <= not(layer0_outputs(559));
    layer1_outputs(2396) <= not(layer0_outputs(154));
    layer1_outputs(2397) <= not(layer0_outputs(1865));
    layer1_outputs(2398) <= not(layer0_outputs(1936)) or (layer0_outputs(1027));
    layer1_outputs(2399) <= not((layer0_outputs(524)) or (layer0_outputs(253)));
    layer1_outputs(2400) <= not((layer0_outputs(445)) and (layer0_outputs(648)));
    layer1_outputs(2401) <= layer0_outputs(656);
    layer1_outputs(2402) <= layer0_outputs(974);
    layer1_outputs(2403) <= not(layer0_outputs(1539));
    layer1_outputs(2404) <= not((layer0_outputs(1230)) or (layer0_outputs(1778)));
    layer1_outputs(2405) <= not((layer0_outputs(2294)) or (layer0_outputs(1695)));
    layer1_outputs(2406) <= (layer0_outputs(865)) and (layer0_outputs(695));
    layer1_outputs(2407) <= '0';
    layer1_outputs(2408) <= '1';
    layer1_outputs(2409) <= (layer0_outputs(1053)) xor (layer0_outputs(2430));
    layer1_outputs(2410) <= (layer0_outputs(1625)) and not (layer0_outputs(1389));
    layer1_outputs(2411) <= not(layer0_outputs(1524)) or (layer0_outputs(2364));
    layer1_outputs(2412) <= (layer0_outputs(1162)) and not (layer0_outputs(1836));
    layer1_outputs(2413) <= not(layer0_outputs(1264));
    layer1_outputs(2414) <= layer0_outputs(929);
    layer1_outputs(2415) <= not((layer0_outputs(1262)) or (layer0_outputs(963)));
    layer1_outputs(2416) <= layer0_outputs(764);
    layer1_outputs(2417) <= (layer0_outputs(1818)) xor (layer0_outputs(1959));
    layer1_outputs(2418) <= not(layer0_outputs(1882)) or (layer0_outputs(2545));
    layer1_outputs(2419) <= not(layer0_outputs(2287));
    layer1_outputs(2420) <= (layer0_outputs(1237)) or (layer0_outputs(1281));
    layer1_outputs(2421) <= (layer0_outputs(395)) and (layer0_outputs(2087));
    layer1_outputs(2422) <= not((layer0_outputs(2145)) or (layer0_outputs(469)));
    layer1_outputs(2423) <= layer0_outputs(1219);
    layer1_outputs(2424) <= (layer0_outputs(2324)) xor (layer0_outputs(1545));
    layer1_outputs(2425) <= (layer0_outputs(2098)) and not (layer0_outputs(1795));
    layer1_outputs(2426) <= layer0_outputs(610);
    layer1_outputs(2427) <= (layer0_outputs(1785)) and not (layer0_outputs(1989));
    layer1_outputs(2428) <= not(layer0_outputs(538)) or (layer0_outputs(1604));
    layer1_outputs(2429) <= (layer0_outputs(519)) and (layer0_outputs(903));
    layer1_outputs(2430) <= (layer0_outputs(45)) or (layer0_outputs(945));
    layer1_outputs(2431) <= (layer0_outputs(2033)) or (layer0_outputs(483));
    layer1_outputs(2432) <= not(layer0_outputs(1987));
    layer1_outputs(2433) <= not(layer0_outputs(1170)) or (layer0_outputs(2007));
    layer1_outputs(2434) <= not(layer0_outputs(136));
    layer1_outputs(2435) <= layer0_outputs(802);
    layer1_outputs(2436) <= (layer0_outputs(728)) and not (layer0_outputs(1995));
    layer1_outputs(2437) <= layer0_outputs(2528);
    layer1_outputs(2438) <= layer0_outputs(1971);
    layer1_outputs(2439) <= (layer0_outputs(1753)) and not (layer0_outputs(1295));
    layer1_outputs(2440) <= (layer0_outputs(1850)) and (layer0_outputs(670));
    layer1_outputs(2441) <= layer0_outputs(769);
    layer1_outputs(2442) <= layer0_outputs(1624);
    layer1_outputs(2443) <= layer0_outputs(1202);
    layer1_outputs(2444) <= not(layer0_outputs(1290));
    layer1_outputs(2445) <= '1';
    layer1_outputs(2446) <= not((layer0_outputs(2208)) and (layer0_outputs(348)));
    layer1_outputs(2447) <= layer0_outputs(322);
    layer1_outputs(2448) <= (layer0_outputs(419)) and not (layer0_outputs(1719));
    layer1_outputs(2449) <= (layer0_outputs(783)) or (layer0_outputs(485));
    layer1_outputs(2450) <= not(layer0_outputs(1687));
    layer1_outputs(2451) <= not((layer0_outputs(1608)) or (layer0_outputs(574)));
    layer1_outputs(2452) <= not((layer0_outputs(1479)) and (layer0_outputs(1735)));
    layer1_outputs(2453) <= (layer0_outputs(54)) and not (layer0_outputs(1698));
    layer1_outputs(2454) <= layer0_outputs(1680);
    layer1_outputs(2455) <= not((layer0_outputs(2373)) and (layer0_outputs(995)));
    layer1_outputs(2456) <= not(layer0_outputs(1342)) or (layer0_outputs(507));
    layer1_outputs(2457) <= not((layer0_outputs(1565)) or (layer0_outputs(1050)));
    layer1_outputs(2458) <= not(layer0_outputs(1120)) or (layer0_outputs(1853));
    layer1_outputs(2459) <= layer0_outputs(1456);
    layer1_outputs(2460) <= not(layer0_outputs(126));
    layer1_outputs(2461) <= (layer0_outputs(1131)) and not (layer0_outputs(399));
    layer1_outputs(2462) <= layer0_outputs(2380);
    layer1_outputs(2463) <= layer0_outputs(379);
    layer1_outputs(2464) <= not(layer0_outputs(292));
    layer1_outputs(2465) <= (layer0_outputs(2117)) and not (layer0_outputs(1806));
    layer1_outputs(2466) <= not((layer0_outputs(1589)) xor (layer0_outputs(1364)));
    layer1_outputs(2467) <= not((layer0_outputs(47)) or (layer0_outputs(2295)));
    layer1_outputs(2468) <= not(layer0_outputs(1404)) or (layer0_outputs(712));
    layer1_outputs(2469) <= layer0_outputs(1694);
    layer1_outputs(2470) <= not(layer0_outputs(666));
    layer1_outputs(2471) <= not((layer0_outputs(968)) or (layer0_outputs(722)));
    layer1_outputs(2472) <= not((layer0_outputs(1963)) xor (layer0_outputs(881)));
    layer1_outputs(2473) <= (layer0_outputs(1621)) and not (layer0_outputs(992));
    layer1_outputs(2474) <= not((layer0_outputs(651)) and (layer0_outputs(763)));
    layer1_outputs(2475) <= (layer0_outputs(227)) and not (layer0_outputs(615));
    layer1_outputs(2476) <= '0';
    layer1_outputs(2477) <= not(layer0_outputs(1919));
    layer1_outputs(2478) <= not((layer0_outputs(1769)) and (layer0_outputs(183)));
    layer1_outputs(2479) <= (layer0_outputs(1931)) and (layer0_outputs(1876));
    layer1_outputs(2480) <= not(layer0_outputs(480));
    layer1_outputs(2481) <= layer0_outputs(2067);
    layer1_outputs(2482) <= not(layer0_outputs(1926));
    layer1_outputs(2483) <= (layer0_outputs(2265)) and not (layer0_outputs(1590));
    layer1_outputs(2484) <= (layer0_outputs(1044)) and (layer0_outputs(996));
    layer1_outputs(2485) <= not(layer0_outputs(2421));
    layer1_outputs(2486) <= (layer0_outputs(153)) and (layer0_outputs(1531));
    layer1_outputs(2487) <= layer0_outputs(1531);
    layer1_outputs(2488) <= layer0_outputs(1546);
    layer1_outputs(2489) <= not(layer0_outputs(532)) or (layer0_outputs(2115));
    layer1_outputs(2490) <= (layer0_outputs(1999)) xor (layer0_outputs(2317));
    layer1_outputs(2491) <= layer0_outputs(1131);
    layer1_outputs(2492) <= layer0_outputs(2421);
    layer1_outputs(2493) <= not((layer0_outputs(674)) and (layer0_outputs(2397)));
    layer1_outputs(2494) <= (layer0_outputs(2533)) and not (layer0_outputs(2063));
    layer1_outputs(2495) <= not(layer0_outputs(2178));
    layer1_outputs(2496) <= layer0_outputs(2446);
    layer1_outputs(2497) <= not((layer0_outputs(2392)) or (layer0_outputs(124)));
    layer1_outputs(2498) <= '0';
    layer1_outputs(2499) <= not(layer0_outputs(420)) or (layer0_outputs(1768));
    layer1_outputs(2500) <= not(layer0_outputs(570));
    layer1_outputs(2501) <= (layer0_outputs(2093)) and not (layer0_outputs(2026));
    layer1_outputs(2502) <= layer0_outputs(382);
    layer1_outputs(2503) <= not(layer0_outputs(1094));
    layer1_outputs(2504) <= (layer0_outputs(1288)) and not (layer0_outputs(724));
    layer1_outputs(2505) <= (layer0_outputs(1079)) and not (layer0_outputs(1411));
    layer1_outputs(2506) <= not(layer0_outputs(364));
    layer1_outputs(2507) <= not((layer0_outputs(890)) and (layer0_outputs(1129)));
    layer1_outputs(2508) <= layer0_outputs(96);
    layer1_outputs(2509) <= '0';
    layer1_outputs(2510) <= not(layer0_outputs(1857));
    layer1_outputs(2511) <= layer0_outputs(552);
    layer1_outputs(2512) <= not((layer0_outputs(904)) and (layer0_outputs(1195)));
    layer1_outputs(2513) <= '0';
    layer1_outputs(2514) <= layer0_outputs(1895);
    layer1_outputs(2515) <= not((layer0_outputs(1145)) and (layer0_outputs(1739)));
    layer1_outputs(2516) <= not(layer0_outputs(1474));
    layer1_outputs(2517) <= not(layer0_outputs(1219));
    layer1_outputs(2518) <= (layer0_outputs(654)) or (layer0_outputs(925));
    layer1_outputs(2519) <= (layer0_outputs(112)) or (layer0_outputs(734));
    layer1_outputs(2520) <= not(layer0_outputs(1712));
    layer1_outputs(2521) <= (layer0_outputs(935)) or (layer0_outputs(423));
    layer1_outputs(2522) <= (layer0_outputs(1619)) and not (layer0_outputs(1213));
    layer1_outputs(2523) <= not(layer0_outputs(2395));
    layer1_outputs(2524) <= not((layer0_outputs(1287)) and (layer0_outputs(2078)));
    layer1_outputs(2525) <= not((layer0_outputs(267)) and (layer0_outputs(1497)));
    layer1_outputs(2526) <= (layer0_outputs(1153)) and not (layer0_outputs(2155));
    layer1_outputs(2527) <= not(layer0_outputs(1417)) or (layer0_outputs(651));
    layer1_outputs(2528) <= not((layer0_outputs(2362)) or (layer0_outputs(1668)));
    layer1_outputs(2529) <= not(layer0_outputs(1694)) or (layer0_outputs(1291));
    layer1_outputs(2530) <= not(layer0_outputs(1420));
    layer1_outputs(2531) <= (layer0_outputs(1922)) and not (layer0_outputs(643));
    layer1_outputs(2532) <= not(layer0_outputs(1752));
    layer1_outputs(2533) <= not(layer0_outputs(2391));
    layer1_outputs(2534) <= not(layer0_outputs(121));
    layer1_outputs(2535) <= layer0_outputs(878);
    layer1_outputs(2536) <= (layer0_outputs(473)) and not (layer0_outputs(713));
    layer1_outputs(2537) <= not(layer0_outputs(205));
    layer1_outputs(2538) <= not((layer0_outputs(40)) or (layer0_outputs(1193)));
    layer1_outputs(2539) <= (layer0_outputs(2140)) or (layer0_outputs(200));
    layer1_outputs(2540) <= layer0_outputs(609);
    layer1_outputs(2541) <= not(layer0_outputs(79));
    layer1_outputs(2542) <= layer0_outputs(2104);
    layer1_outputs(2543) <= layer0_outputs(2522);
    layer1_outputs(2544) <= not((layer0_outputs(2390)) or (layer0_outputs(1894)));
    layer1_outputs(2545) <= (layer0_outputs(1484)) and (layer0_outputs(77));
    layer1_outputs(2546) <= not(layer0_outputs(46)) or (layer0_outputs(413));
    layer1_outputs(2547) <= (layer0_outputs(1647)) or (layer0_outputs(374));
    layer1_outputs(2548) <= (layer0_outputs(1832)) and not (layer0_outputs(2161));
    layer1_outputs(2549) <= '0';
    layer1_outputs(2550) <= layer0_outputs(545);
    layer1_outputs(2551) <= layer0_outputs(1163);
    layer1_outputs(2552) <= not(layer0_outputs(1325)) or (layer0_outputs(1676));
    layer1_outputs(2553) <= layer0_outputs(2247);
    layer1_outputs(2554) <= not(layer0_outputs(723));
    layer1_outputs(2555) <= not(layer0_outputs(786)) or (layer0_outputs(873));
    layer1_outputs(2556) <= not((layer0_outputs(2558)) or (layer0_outputs(1083)));
    layer1_outputs(2557) <= layer0_outputs(1626);
    layer1_outputs(2558) <= not(layer0_outputs(50));
    layer1_outputs(2559) <= '0';
    layer2_outputs(0) <= not(layer1_outputs(2385));
    layer2_outputs(1) <= layer1_outputs(2481);
    layer2_outputs(2) <= (layer1_outputs(969)) and (layer1_outputs(1482));
    layer2_outputs(3) <= not(layer1_outputs(2473));
    layer2_outputs(4) <= layer1_outputs(1574);
    layer2_outputs(5) <= not(layer1_outputs(1325));
    layer2_outputs(6) <= not(layer1_outputs(1015));
    layer2_outputs(7) <= (layer1_outputs(1767)) and (layer1_outputs(183));
    layer2_outputs(8) <= (layer1_outputs(2395)) and not (layer1_outputs(1264));
    layer2_outputs(9) <= not((layer1_outputs(467)) and (layer1_outputs(1302)));
    layer2_outputs(10) <= (layer1_outputs(329)) and (layer1_outputs(705));
    layer2_outputs(11) <= not(layer1_outputs(2153));
    layer2_outputs(12) <= not(layer1_outputs(1500)) or (layer1_outputs(617));
    layer2_outputs(13) <= not(layer1_outputs(587));
    layer2_outputs(14) <= layer1_outputs(1390);
    layer2_outputs(15) <= (layer1_outputs(1387)) and not (layer1_outputs(790));
    layer2_outputs(16) <= not((layer1_outputs(269)) or (layer1_outputs(1027)));
    layer2_outputs(17) <= not(layer1_outputs(914)) or (layer1_outputs(200));
    layer2_outputs(18) <= (layer1_outputs(1025)) and not (layer1_outputs(2044));
    layer2_outputs(19) <= not((layer1_outputs(1089)) and (layer1_outputs(62)));
    layer2_outputs(20) <= '1';
    layer2_outputs(21) <= not(layer1_outputs(2528));
    layer2_outputs(22) <= layer1_outputs(1492);
    layer2_outputs(23) <= not(layer1_outputs(1281));
    layer2_outputs(24) <= layer1_outputs(1443);
    layer2_outputs(25) <= (layer1_outputs(947)) and not (layer1_outputs(1902));
    layer2_outputs(26) <= not(layer1_outputs(288));
    layer2_outputs(27) <= not(layer1_outputs(1313));
    layer2_outputs(28) <= (layer1_outputs(530)) and (layer1_outputs(273));
    layer2_outputs(29) <= layer1_outputs(105);
    layer2_outputs(30) <= layer1_outputs(2010);
    layer2_outputs(31) <= not(layer1_outputs(445));
    layer2_outputs(32) <= (layer1_outputs(296)) xor (layer1_outputs(700));
    layer2_outputs(33) <= (layer1_outputs(606)) and (layer1_outputs(1375));
    layer2_outputs(34) <= not(layer1_outputs(618)) or (layer1_outputs(1090));
    layer2_outputs(35) <= not((layer1_outputs(2323)) and (layer1_outputs(1459)));
    layer2_outputs(36) <= '0';
    layer2_outputs(37) <= (layer1_outputs(317)) and (layer1_outputs(1490));
    layer2_outputs(38) <= not(layer1_outputs(1888));
    layer2_outputs(39) <= not(layer1_outputs(1057));
    layer2_outputs(40) <= (layer1_outputs(1609)) or (layer1_outputs(2337));
    layer2_outputs(41) <= not(layer1_outputs(1947));
    layer2_outputs(42) <= (layer1_outputs(2106)) and not (layer1_outputs(858));
    layer2_outputs(43) <= not(layer1_outputs(888));
    layer2_outputs(44) <= (layer1_outputs(2095)) or (layer1_outputs(1866));
    layer2_outputs(45) <= (layer1_outputs(1566)) and not (layer1_outputs(131));
    layer2_outputs(46) <= layer1_outputs(2059);
    layer2_outputs(47) <= not(layer1_outputs(1219));
    layer2_outputs(48) <= (layer1_outputs(2320)) and not (layer1_outputs(2150));
    layer2_outputs(49) <= (layer1_outputs(857)) and (layer1_outputs(796));
    layer2_outputs(50) <= '0';
    layer2_outputs(51) <= (layer1_outputs(205)) xor (layer1_outputs(717));
    layer2_outputs(52) <= (layer1_outputs(2300)) and (layer1_outputs(1789));
    layer2_outputs(53) <= not(layer1_outputs(18)) or (layer1_outputs(2508));
    layer2_outputs(54) <= layer1_outputs(392);
    layer2_outputs(55) <= (layer1_outputs(49)) and (layer1_outputs(1326));
    layer2_outputs(56) <= not(layer1_outputs(2275));
    layer2_outputs(57) <= not(layer1_outputs(611)) or (layer1_outputs(2047));
    layer2_outputs(58) <= not(layer1_outputs(39)) or (layer1_outputs(1094));
    layer2_outputs(59) <= not((layer1_outputs(1979)) or (layer1_outputs(757)));
    layer2_outputs(60) <= (layer1_outputs(49)) and (layer1_outputs(1944));
    layer2_outputs(61) <= not((layer1_outputs(444)) and (layer1_outputs(1862)));
    layer2_outputs(62) <= layer1_outputs(1960);
    layer2_outputs(63) <= (layer1_outputs(661)) and not (layer1_outputs(551));
    layer2_outputs(64) <= layer1_outputs(1390);
    layer2_outputs(65) <= (layer1_outputs(1407)) and not (layer1_outputs(1575));
    layer2_outputs(66) <= layer1_outputs(1943);
    layer2_outputs(67) <= not(layer1_outputs(1799));
    layer2_outputs(68) <= (layer1_outputs(1468)) or (layer1_outputs(2448));
    layer2_outputs(69) <= (layer1_outputs(739)) and not (layer1_outputs(2417));
    layer2_outputs(70) <= not((layer1_outputs(422)) or (layer1_outputs(1046)));
    layer2_outputs(71) <= not((layer1_outputs(2490)) xor (layer1_outputs(1022)));
    layer2_outputs(72) <= layer1_outputs(765);
    layer2_outputs(73) <= '0';
    layer2_outputs(74) <= '1';
    layer2_outputs(75) <= (layer1_outputs(230)) and not (layer1_outputs(2426));
    layer2_outputs(76) <= '1';
    layer2_outputs(77) <= (layer1_outputs(1637)) and not (layer1_outputs(2525));
    layer2_outputs(78) <= not(layer1_outputs(266));
    layer2_outputs(79) <= not(layer1_outputs(866));
    layer2_outputs(80) <= not(layer1_outputs(1453));
    layer2_outputs(81) <= not(layer1_outputs(1495)) or (layer1_outputs(720));
    layer2_outputs(82) <= not(layer1_outputs(802));
    layer2_outputs(83) <= layer1_outputs(2090);
    layer2_outputs(84) <= (layer1_outputs(374)) and (layer1_outputs(1488));
    layer2_outputs(85) <= not(layer1_outputs(2011));
    layer2_outputs(86) <= not(layer1_outputs(366));
    layer2_outputs(87) <= (layer1_outputs(1041)) and (layer1_outputs(2435));
    layer2_outputs(88) <= not(layer1_outputs(1503));
    layer2_outputs(89) <= not(layer1_outputs(2139));
    layer2_outputs(90) <= not(layer1_outputs(1438));
    layer2_outputs(91) <= layer1_outputs(1991);
    layer2_outputs(92) <= not(layer1_outputs(891));
    layer2_outputs(93) <= layer1_outputs(1226);
    layer2_outputs(94) <= not(layer1_outputs(656));
    layer2_outputs(95) <= (layer1_outputs(1151)) and not (layer1_outputs(1955));
    layer2_outputs(96) <= not(layer1_outputs(353));
    layer2_outputs(97) <= (layer1_outputs(736)) and (layer1_outputs(1965));
    layer2_outputs(98) <= (layer1_outputs(2414)) and not (layer1_outputs(1420));
    layer2_outputs(99) <= not(layer1_outputs(1181));
    layer2_outputs(100) <= (layer1_outputs(1716)) or (layer1_outputs(344));
    layer2_outputs(101) <= layer1_outputs(680);
    layer2_outputs(102) <= not(layer1_outputs(2324));
    layer2_outputs(103) <= layer1_outputs(1314);
    layer2_outputs(104) <= not(layer1_outputs(12));
    layer2_outputs(105) <= not((layer1_outputs(1235)) or (layer1_outputs(967)));
    layer2_outputs(106) <= not(layer1_outputs(382));
    layer2_outputs(107) <= layer1_outputs(1828);
    layer2_outputs(108) <= not(layer1_outputs(1163));
    layer2_outputs(109) <= layer1_outputs(404);
    layer2_outputs(110) <= not(layer1_outputs(523)) or (layer1_outputs(425));
    layer2_outputs(111) <= layer1_outputs(1481);
    layer2_outputs(112) <= not((layer1_outputs(2003)) and (layer1_outputs(727)));
    layer2_outputs(113) <= layer1_outputs(1485);
    layer2_outputs(114) <= not(layer1_outputs(1465));
    layer2_outputs(115) <= not((layer1_outputs(211)) xor (layer1_outputs(2335)));
    layer2_outputs(116) <= not(layer1_outputs(1307));
    layer2_outputs(117) <= not(layer1_outputs(2020));
    layer2_outputs(118) <= not(layer1_outputs(1497));
    layer2_outputs(119) <= layer1_outputs(2224);
    layer2_outputs(120) <= layer1_outputs(987);
    layer2_outputs(121) <= '0';
    layer2_outputs(122) <= layer1_outputs(2455);
    layer2_outputs(123) <= not(layer1_outputs(941));
    layer2_outputs(124) <= not(layer1_outputs(2468)) or (layer1_outputs(1950));
    layer2_outputs(125) <= (layer1_outputs(1594)) and not (layer1_outputs(229));
    layer2_outputs(126) <= layer1_outputs(1843);
    layer2_outputs(127) <= not(layer1_outputs(1602)) or (layer1_outputs(2274));
    layer2_outputs(128) <= (layer1_outputs(619)) and (layer1_outputs(522));
    layer2_outputs(129) <= (layer1_outputs(241)) or (layer1_outputs(519));
    layer2_outputs(130) <= (layer1_outputs(2404)) and (layer1_outputs(1283));
    layer2_outputs(131) <= not(layer1_outputs(1650));
    layer2_outputs(132) <= layer1_outputs(2446);
    layer2_outputs(133) <= (layer1_outputs(1926)) xor (layer1_outputs(657));
    layer2_outputs(134) <= layer1_outputs(656);
    layer2_outputs(135) <= (layer1_outputs(523)) and (layer1_outputs(372));
    layer2_outputs(136) <= (layer1_outputs(163)) xor (layer1_outputs(901));
    layer2_outputs(137) <= not(layer1_outputs(644));
    layer2_outputs(138) <= not(layer1_outputs(1922)) or (layer1_outputs(2506));
    layer2_outputs(139) <= layer1_outputs(1067);
    layer2_outputs(140) <= (layer1_outputs(1668)) xor (layer1_outputs(1756));
    layer2_outputs(141) <= layer1_outputs(318);
    layer2_outputs(142) <= layer1_outputs(1817);
    layer2_outputs(143) <= layer1_outputs(641);
    layer2_outputs(144) <= layer1_outputs(1000);
    layer2_outputs(145) <= layer1_outputs(2385);
    layer2_outputs(146) <= not(layer1_outputs(28));
    layer2_outputs(147) <= layer1_outputs(378);
    layer2_outputs(148) <= not(layer1_outputs(2296));
    layer2_outputs(149) <= (layer1_outputs(621)) and (layer1_outputs(510));
    layer2_outputs(150) <= (layer1_outputs(1605)) and (layer1_outputs(1137));
    layer2_outputs(151) <= not((layer1_outputs(1556)) or (layer1_outputs(2170)));
    layer2_outputs(152) <= (layer1_outputs(1060)) and (layer1_outputs(1973));
    layer2_outputs(153) <= (layer1_outputs(979)) and not (layer1_outputs(1442));
    layer2_outputs(154) <= (layer1_outputs(460)) and not (layer1_outputs(1640));
    layer2_outputs(155) <= not(layer1_outputs(1125));
    layer2_outputs(156) <= not(layer1_outputs(204));
    layer2_outputs(157) <= not(layer1_outputs(2100));
    layer2_outputs(158) <= (layer1_outputs(1504)) or (layer1_outputs(2427));
    layer2_outputs(159) <= not(layer1_outputs(1193));
    layer2_outputs(160) <= layer1_outputs(1638);
    layer2_outputs(161) <= not(layer1_outputs(545));
    layer2_outputs(162) <= not((layer1_outputs(1593)) or (layer1_outputs(1031)));
    layer2_outputs(163) <= not((layer1_outputs(950)) and (layer1_outputs(1263)));
    layer2_outputs(164) <= not(layer1_outputs(2214));
    layer2_outputs(165) <= layer1_outputs(1392);
    layer2_outputs(166) <= not(layer1_outputs(1761));
    layer2_outputs(167) <= (layer1_outputs(616)) and not (layer1_outputs(1921));
    layer2_outputs(168) <= layer1_outputs(318);
    layer2_outputs(169) <= layer1_outputs(165);
    layer2_outputs(170) <= layer1_outputs(42);
    layer2_outputs(171) <= not(layer1_outputs(102));
    layer2_outputs(172) <= layer1_outputs(1956);
    layer2_outputs(173) <= not(layer1_outputs(1276)) or (layer1_outputs(896));
    layer2_outputs(174) <= not(layer1_outputs(892)) or (layer1_outputs(1351));
    layer2_outputs(175) <= not(layer1_outputs(2285)) or (layer1_outputs(1026));
    layer2_outputs(176) <= layer1_outputs(2091);
    layer2_outputs(177) <= not(layer1_outputs(240)) or (layer1_outputs(944));
    layer2_outputs(178) <= not(layer1_outputs(1582));
    layer2_outputs(179) <= '0';
    layer2_outputs(180) <= not((layer1_outputs(462)) or (layer1_outputs(1567)));
    layer2_outputs(181) <= (layer1_outputs(149)) and (layer1_outputs(2081));
    layer2_outputs(182) <= (layer1_outputs(898)) and not (layer1_outputs(1702));
    layer2_outputs(183) <= (layer1_outputs(2002)) and (layer1_outputs(1467));
    layer2_outputs(184) <= (layer1_outputs(1977)) xor (layer1_outputs(2026));
    layer2_outputs(185) <= not(layer1_outputs(202));
    layer2_outputs(186) <= not((layer1_outputs(1181)) or (layer1_outputs(529)));
    layer2_outputs(187) <= (layer1_outputs(791)) xor (layer1_outputs(1512));
    layer2_outputs(188) <= not(layer1_outputs(1076)) or (layer1_outputs(1057));
    layer2_outputs(189) <= not(layer1_outputs(1276));
    layer2_outputs(190) <= not(layer1_outputs(1411));
    layer2_outputs(191) <= not(layer1_outputs(1896));
    layer2_outputs(192) <= layer1_outputs(2264);
    layer2_outputs(193) <= (layer1_outputs(1860)) or (layer1_outputs(1304));
    layer2_outputs(194) <= not((layer1_outputs(1209)) and (layer1_outputs(1144)));
    layer2_outputs(195) <= (layer1_outputs(104)) or (layer1_outputs(13));
    layer2_outputs(196) <= (layer1_outputs(876)) and (layer1_outputs(5));
    layer2_outputs(197) <= layer1_outputs(714);
    layer2_outputs(198) <= not((layer1_outputs(572)) and (layer1_outputs(738)));
    layer2_outputs(199) <= not(layer1_outputs(2470));
    layer2_outputs(200) <= (layer1_outputs(45)) xor (layer1_outputs(2215));
    layer2_outputs(201) <= not(layer1_outputs(1034));
    layer2_outputs(202) <= (layer1_outputs(454)) and not (layer1_outputs(1156));
    layer2_outputs(203) <= layer1_outputs(2234);
    layer2_outputs(204) <= (layer1_outputs(475)) and not (layer1_outputs(1513));
    layer2_outputs(205) <= not(layer1_outputs(1056));
    layer2_outputs(206) <= '1';
    layer2_outputs(207) <= layer1_outputs(573);
    layer2_outputs(208) <= (layer1_outputs(499)) and not (layer1_outputs(270));
    layer2_outputs(209) <= not((layer1_outputs(1665)) or (layer1_outputs(1721)));
    layer2_outputs(210) <= not(layer1_outputs(488));
    layer2_outputs(211) <= not(layer1_outputs(1034));
    layer2_outputs(212) <= not((layer1_outputs(2349)) and (layer1_outputs(2499)));
    layer2_outputs(213) <= not(layer1_outputs(1871)) or (layer1_outputs(1433));
    layer2_outputs(214) <= (layer1_outputs(1560)) and not (layer1_outputs(1299));
    layer2_outputs(215) <= (layer1_outputs(722)) and (layer1_outputs(1434));
    layer2_outputs(216) <= not(layer1_outputs(1007));
    layer2_outputs(217) <= not(layer1_outputs(2520));
    layer2_outputs(218) <= not(layer1_outputs(1207)) or (layer1_outputs(2411));
    layer2_outputs(219) <= (layer1_outputs(1006)) and not (layer1_outputs(1440));
    layer2_outputs(220) <= (layer1_outputs(1689)) or (layer1_outputs(2454));
    layer2_outputs(221) <= (layer1_outputs(1699)) and not (layer1_outputs(14));
    layer2_outputs(222) <= layer1_outputs(2188);
    layer2_outputs(223) <= (layer1_outputs(109)) and not (layer1_outputs(364));
    layer2_outputs(224) <= (layer1_outputs(1132)) and not (layer1_outputs(1292));
    layer2_outputs(225) <= not(layer1_outputs(2401));
    layer2_outputs(226) <= layer1_outputs(1809);
    layer2_outputs(227) <= (layer1_outputs(1366)) or (layer1_outputs(2295));
    layer2_outputs(228) <= not(layer1_outputs(201)) or (layer1_outputs(880));
    layer2_outputs(229) <= layer1_outputs(474);
    layer2_outputs(230) <= layer1_outputs(843);
    layer2_outputs(231) <= not(layer1_outputs(1591));
    layer2_outputs(232) <= (layer1_outputs(1713)) and not (layer1_outputs(1570));
    layer2_outputs(233) <= (layer1_outputs(1740)) or (layer1_outputs(1507));
    layer2_outputs(234) <= not(layer1_outputs(77)) or (layer1_outputs(461));
    layer2_outputs(235) <= not((layer1_outputs(758)) or (layer1_outputs(1839)));
    layer2_outputs(236) <= layer1_outputs(2029);
    layer2_outputs(237) <= layer1_outputs(1729);
    layer2_outputs(238) <= (layer1_outputs(2081)) xor (layer1_outputs(2407));
    layer2_outputs(239) <= layer1_outputs(724);
    layer2_outputs(240) <= (layer1_outputs(347)) and not (layer1_outputs(783));
    layer2_outputs(241) <= layer1_outputs(1120);
    layer2_outputs(242) <= layer1_outputs(1692);
    layer2_outputs(243) <= (layer1_outputs(562)) and not (layer1_outputs(665));
    layer2_outputs(244) <= (layer1_outputs(1653)) and not (layer1_outputs(1435));
    layer2_outputs(245) <= (layer1_outputs(310)) and not (layer1_outputs(2063));
    layer2_outputs(246) <= not(layer1_outputs(1501));
    layer2_outputs(247) <= (layer1_outputs(880)) or (layer1_outputs(997));
    layer2_outputs(248) <= (layer1_outputs(188)) or (layer1_outputs(438));
    layer2_outputs(249) <= not((layer1_outputs(1961)) xor (layer1_outputs(2558)));
    layer2_outputs(250) <= not((layer1_outputs(383)) and (layer1_outputs(2358)));
    layer2_outputs(251) <= not((layer1_outputs(1731)) and (layer1_outputs(2465)));
    layer2_outputs(252) <= layer1_outputs(2379);
    layer2_outputs(253) <= not(layer1_outputs(624));
    layer2_outputs(254) <= not(layer1_outputs(1353)) or (layer1_outputs(780));
    layer2_outputs(255) <= '0';
    layer2_outputs(256) <= not(layer1_outputs(2049)) or (layer1_outputs(1735));
    layer2_outputs(257) <= not((layer1_outputs(392)) and (layer1_outputs(2375)));
    layer2_outputs(258) <= not(layer1_outputs(2542));
    layer2_outputs(259) <= not(layer1_outputs(2037));
    layer2_outputs(260) <= not((layer1_outputs(686)) and (layer1_outputs(905)));
    layer2_outputs(261) <= layer1_outputs(1396);
    layer2_outputs(262) <= not(layer1_outputs(1409));
    layer2_outputs(263) <= (layer1_outputs(799)) and not (layer1_outputs(1598));
    layer2_outputs(264) <= not(layer1_outputs(2338)) or (layer1_outputs(498));
    layer2_outputs(265) <= (layer1_outputs(785)) or (layer1_outputs(258));
    layer2_outputs(266) <= (layer1_outputs(923)) and (layer1_outputs(2327));
    layer2_outputs(267) <= not((layer1_outputs(1544)) and (layer1_outputs(917)));
    layer2_outputs(268) <= layer1_outputs(1779);
    layer2_outputs(269) <= layer1_outputs(147);
    layer2_outputs(270) <= not(layer1_outputs(1027));
    layer2_outputs(271) <= (layer1_outputs(1116)) and not (layer1_outputs(141));
    layer2_outputs(272) <= layer1_outputs(2007);
    layer2_outputs(273) <= '1';
    layer2_outputs(274) <= (layer1_outputs(41)) or (layer1_outputs(1848));
    layer2_outputs(275) <= not((layer1_outputs(1468)) or (layer1_outputs(1073)));
    layer2_outputs(276) <= (layer1_outputs(316)) and not (layer1_outputs(2152));
    layer2_outputs(277) <= not(layer1_outputs(2435)) or (layer1_outputs(2276));
    layer2_outputs(278) <= not(layer1_outputs(1811));
    layer2_outputs(279) <= layer1_outputs(2225);
    layer2_outputs(280) <= '1';
    layer2_outputs(281) <= layer1_outputs(663);
    layer2_outputs(282) <= not(layer1_outputs(2410));
    layer2_outputs(283) <= not(layer1_outputs(2027));
    layer2_outputs(284) <= (layer1_outputs(719)) xor (layer1_outputs(399));
    layer2_outputs(285) <= layer1_outputs(621);
    layer2_outputs(286) <= not(layer1_outputs(187));
    layer2_outputs(287) <= not(layer1_outputs(1755));
    layer2_outputs(288) <= layer1_outputs(1164);
    layer2_outputs(289) <= (layer1_outputs(1564)) and (layer1_outputs(1702));
    layer2_outputs(290) <= layer1_outputs(1678);
    layer2_outputs(291) <= (layer1_outputs(1912)) or (layer1_outputs(1382));
    layer2_outputs(292) <= not(layer1_outputs(1355));
    layer2_outputs(293) <= layer1_outputs(482);
    layer2_outputs(294) <= (layer1_outputs(820)) xor (layer1_outputs(761));
    layer2_outputs(295) <= layer1_outputs(1549);
    layer2_outputs(296) <= not(layer1_outputs(2482));
    layer2_outputs(297) <= not(layer1_outputs(1170));
    layer2_outputs(298) <= layer1_outputs(1215);
    layer2_outputs(299) <= layer1_outputs(1550);
    layer2_outputs(300) <= (layer1_outputs(1393)) or (layer1_outputs(1559));
    layer2_outputs(301) <= not(layer1_outputs(1074)) or (layer1_outputs(1600));
    layer2_outputs(302) <= layer1_outputs(1933);
    layer2_outputs(303) <= layer1_outputs(2040);
    layer2_outputs(304) <= (layer1_outputs(1729)) or (layer1_outputs(2532));
    layer2_outputs(305) <= not((layer1_outputs(1200)) and (layer1_outputs(1895)));
    layer2_outputs(306) <= not(layer1_outputs(1249)) or (layer1_outputs(2392));
    layer2_outputs(307) <= (layer1_outputs(2193)) and not (layer1_outputs(1212));
    layer2_outputs(308) <= layer1_outputs(1338);
    layer2_outputs(309) <= (layer1_outputs(1811)) and not (layer1_outputs(1123));
    layer2_outputs(310) <= layer1_outputs(2252);
    layer2_outputs(311) <= (layer1_outputs(673)) and (layer1_outputs(2171));
    layer2_outputs(312) <= not((layer1_outputs(625)) or (layer1_outputs(2437)));
    layer2_outputs(313) <= not(layer1_outputs(1657)) or (layer1_outputs(2306));
    layer2_outputs(314) <= not(layer1_outputs(244)) or (layer1_outputs(2252));
    layer2_outputs(315) <= layer1_outputs(2307);
    layer2_outputs(316) <= not(layer1_outputs(255));
    layer2_outputs(317) <= (layer1_outputs(1760)) and not (layer1_outputs(1951));
    layer2_outputs(318) <= not(layer1_outputs(1843));
    layer2_outputs(319) <= (layer1_outputs(2496)) or (layer1_outputs(2133));
    layer2_outputs(320) <= layer1_outputs(340);
    layer2_outputs(321) <= not((layer1_outputs(1324)) and (layer1_outputs(1218)));
    layer2_outputs(322) <= not(layer1_outputs(365));
    layer2_outputs(323) <= '1';
    layer2_outputs(324) <= not(layer1_outputs(2271)) or (layer1_outputs(1444));
    layer2_outputs(325) <= layer1_outputs(1604);
    layer2_outputs(326) <= not(layer1_outputs(2514)) or (layer1_outputs(482));
    layer2_outputs(327) <= not(layer1_outputs(1231));
    layer2_outputs(328) <= layer1_outputs(1070);
    layer2_outputs(329) <= not((layer1_outputs(2556)) or (layer1_outputs(1062)));
    layer2_outputs(330) <= not(layer1_outputs(1424));
    layer2_outputs(331) <= layer1_outputs(579);
    layer2_outputs(332) <= layer1_outputs(1505);
    layer2_outputs(333) <= (layer1_outputs(15)) and (layer1_outputs(2017));
    layer2_outputs(334) <= not(layer1_outputs(938)) or (layer1_outputs(1241));
    layer2_outputs(335) <= '0';
    layer2_outputs(336) <= layer1_outputs(387);
    layer2_outputs(337) <= not(layer1_outputs(914)) or (layer1_outputs(2106));
    layer2_outputs(338) <= not((layer1_outputs(576)) or (layer1_outputs(977)));
    layer2_outputs(339) <= layer1_outputs(50);
    layer2_outputs(340) <= not(layer1_outputs(2267)) or (layer1_outputs(1426));
    layer2_outputs(341) <= layer1_outputs(506);
    layer2_outputs(342) <= (layer1_outputs(1708)) and not (layer1_outputs(125));
    layer2_outputs(343) <= not(layer1_outputs(32));
    layer2_outputs(344) <= (layer1_outputs(1606)) and not (layer1_outputs(1075));
    layer2_outputs(345) <= not(layer1_outputs(1327));
    layer2_outputs(346) <= not(layer1_outputs(355)) or (layer1_outputs(809));
    layer2_outputs(347) <= not((layer1_outputs(149)) or (layer1_outputs(872)));
    layer2_outputs(348) <= (layer1_outputs(377)) or (layer1_outputs(1707));
    layer2_outputs(349) <= (layer1_outputs(2107)) and (layer1_outputs(1430));
    layer2_outputs(350) <= layer1_outputs(1763);
    layer2_outputs(351) <= not(layer1_outputs(126)) or (layer1_outputs(776));
    layer2_outputs(352) <= (layer1_outputs(2190)) and (layer1_outputs(1897));
    layer2_outputs(353) <= not(layer1_outputs(1654));
    layer2_outputs(354) <= not(layer1_outputs(1462)) or (layer1_outputs(429));
    layer2_outputs(355) <= not(layer1_outputs(2332));
    layer2_outputs(356) <= not((layer1_outputs(1055)) or (layer1_outputs(1599)));
    layer2_outputs(357) <= not(layer1_outputs(1806)) or (layer1_outputs(757));
    layer2_outputs(358) <= layer1_outputs(531);
    layer2_outputs(359) <= (layer1_outputs(1377)) and not (layer1_outputs(981));
    layer2_outputs(360) <= not(layer1_outputs(2013));
    layer2_outputs(361) <= layer1_outputs(2507);
    layer2_outputs(362) <= not((layer1_outputs(2205)) and (layer1_outputs(302)));
    layer2_outputs(363) <= (layer1_outputs(1742)) and not (layer1_outputs(2365));
    layer2_outputs(364) <= not(layer1_outputs(1220));
    layer2_outputs(365) <= layer1_outputs(1407);
    layer2_outputs(366) <= not(layer1_outputs(2340)) or (layer1_outputs(687));
    layer2_outputs(367) <= not(layer1_outputs(1683));
    layer2_outputs(368) <= not(layer1_outputs(1571));
    layer2_outputs(369) <= not(layer1_outputs(1461)) or (layer1_outputs(351));
    layer2_outputs(370) <= (layer1_outputs(1820)) or (layer1_outputs(1533));
    layer2_outputs(371) <= not(layer1_outputs(81));
    layer2_outputs(372) <= layer1_outputs(442);
    layer2_outputs(373) <= not(layer1_outputs(1175));
    layer2_outputs(374) <= (layer1_outputs(1936)) and not (layer1_outputs(1156));
    layer2_outputs(375) <= (layer1_outputs(1130)) and (layer1_outputs(251));
    layer2_outputs(376) <= not(layer1_outputs(1506)) or (layer1_outputs(1386));
    layer2_outputs(377) <= not(layer1_outputs(1064));
    layer2_outputs(378) <= (layer1_outputs(338)) and not (layer1_outputs(2384));
    layer2_outputs(379) <= layer1_outputs(884);
    layer2_outputs(380) <= not(layer1_outputs(382));
    layer2_outputs(381) <= not((layer1_outputs(1083)) or (layer1_outputs(2308)));
    layer2_outputs(382) <= layer1_outputs(910);
    layer2_outputs(383) <= not(layer1_outputs(2033));
    layer2_outputs(384) <= not(layer1_outputs(659));
    layer2_outputs(385) <= not((layer1_outputs(24)) and (layer1_outputs(1986)));
    layer2_outputs(386) <= not(layer1_outputs(2539));
    layer2_outputs(387) <= not(layer1_outputs(2438)) or (layer1_outputs(11));
    layer2_outputs(388) <= (layer1_outputs(1297)) and (layer1_outputs(34));
    layer2_outputs(389) <= not(layer1_outputs(2185));
    layer2_outputs(390) <= (layer1_outputs(1442)) or (layer1_outputs(836));
    layer2_outputs(391) <= not((layer1_outputs(769)) xor (layer1_outputs(1187)));
    layer2_outputs(392) <= layer1_outputs(17);
    layer2_outputs(393) <= '1';
    layer2_outputs(394) <= (layer1_outputs(1944)) and not (layer1_outputs(1054));
    layer2_outputs(395) <= layer1_outputs(1791);
    layer2_outputs(396) <= not(layer1_outputs(2517));
    layer2_outputs(397) <= not(layer1_outputs(314)) or (layer1_outputs(554));
    layer2_outputs(398) <= not(layer1_outputs(2279));
    layer2_outputs(399) <= not(layer1_outputs(37));
    layer2_outputs(400) <= (layer1_outputs(1469)) or (layer1_outputs(780));
    layer2_outputs(401) <= layer1_outputs(1719);
    layer2_outputs(402) <= layer1_outputs(810);
    layer2_outputs(403) <= not(layer1_outputs(976)) or (layer1_outputs(726));
    layer2_outputs(404) <= (layer1_outputs(2476)) and (layer1_outputs(801));
    layer2_outputs(405) <= not(layer1_outputs(1737)) or (layer1_outputs(2268));
    layer2_outputs(406) <= layer1_outputs(611);
    layer2_outputs(407) <= (layer1_outputs(972)) xor (layer1_outputs(716));
    layer2_outputs(408) <= not(layer1_outputs(2198));
    layer2_outputs(409) <= (layer1_outputs(771)) and not (layer1_outputs(588));
    layer2_outputs(410) <= layer1_outputs(729);
    layer2_outputs(411) <= (layer1_outputs(357)) or (layer1_outputs(1873));
    layer2_outputs(412) <= not(layer1_outputs(238)) or (layer1_outputs(118));
    layer2_outputs(413) <= not((layer1_outputs(2108)) or (layer1_outputs(859)));
    layer2_outputs(414) <= layer1_outputs(939);
    layer2_outputs(415) <= layer1_outputs(1270);
    layer2_outputs(416) <= (layer1_outputs(2116)) and not (layer1_outputs(606));
    layer2_outputs(417) <= layer1_outputs(1840);
    layer2_outputs(418) <= not(layer1_outputs(2123));
    layer2_outputs(419) <= not(layer1_outputs(6)) or (layer1_outputs(1646));
    layer2_outputs(420) <= layer1_outputs(847);
    layer2_outputs(421) <= (layer1_outputs(1872)) and not (layer1_outputs(1075));
    layer2_outputs(422) <= not(layer1_outputs(2512));
    layer2_outputs(423) <= layer1_outputs(1704);
    layer2_outputs(424) <= (layer1_outputs(1259)) and not (layer1_outputs(139));
    layer2_outputs(425) <= not((layer1_outputs(504)) or (layer1_outputs(798)));
    layer2_outputs(426) <= not(layer1_outputs(1379));
    layer2_outputs(427) <= layer1_outputs(908);
    layer2_outputs(428) <= (layer1_outputs(1257)) and not (layer1_outputs(2288));
    layer2_outputs(429) <= (layer1_outputs(1214)) and not (layer1_outputs(2399));
    layer2_outputs(430) <= not((layer1_outputs(99)) or (layer1_outputs(540)));
    layer2_outputs(431) <= layer1_outputs(2085);
    layer2_outputs(432) <= (layer1_outputs(1879)) and not (layer1_outputs(1721));
    layer2_outputs(433) <= not((layer1_outputs(1474)) and (layer1_outputs(1996)));
    layer2_outputs(434) <= not(layer1_outputs(2087));
    layer2_outputs(435) <= layer1_outputs(1441);
    layer2_outputs(436) <= (layer1_outputs(145)) and not (layer1_outputs(146));
    layer2_outputs(437) <= (layer1_outputs(1758)) xor (layer1_outputs(1586));
    layer2_outputs(438) <= not(layer1_outputs(2137)) or (layer1_outputs(519));
    layer2_outputs(439) <= not(layer1_outputs(1117));
    layer2_outputs(440) <= layer1_outputs(540);
    layer2_outputs(441) <= not(layer1_outputs(1774));
    layer2_outputs(442) <= not(layer1_outputs(591));
    layer2_outputs(443) <= not((layer1_outputs(1972)) or (layer1_outputs(1504)));
    layer2_outputs(444) <= not(layer1_outputs(1047));
    layer2_outputs(445) <= not(layer1_outputs(1323));
    layer2_outputs(446) <= not(layer1_outputs(2390)) or (layer1_outputs(167));
    layer2_outputs(447) <= layer1_outputs(83);
    layer2_outputs(448) <= not((layer1_outputs(738)) or (layer1_outputs(1683)));
    layer2_outputs(449) <= not(layer1_outputs(1578));
    layer2_outputs(450) <= layer1_outputs(1863);
    layer2_outputs(451) <= not(layer1_outputs(1803));
    layer2_outputs(452) <= layer1_outputs(390);
    layer2_outputs(453) <= (layer1_outputs(1600)) and not (layer1_outputs(324));
    layer2_outputs(454) <= not(layer1_outputs(627));
    layer2_outputs(455) <= not(layer1_outputs(1318)) or (layer1_outputs(411));
    layer2_outputs(456) <= not(layer1_outputs(1091));
    layer2_outputs(457) <= (layer1_outputs(521)) and not (layer1_outputs(2304));
    layer2_outputs(458) <= '0';
    layer2_outputs(459) <= (layer1_outputs(1256)) or (layer1_outputs(1049));
    layer2_outputs(460) <= not(layer1_outputs(1062));
    layer2_outputs(461) <= not(layer1_outputs(1974)) or (layer1_outputs(875));
    layer2_outputs(462) <= (layer1_outputs(563)) and (layer1_outputs(259));
    layer2_outputs(463) <= layer1_outputs(175);
    layer2_outputs(464) <= layer1_outputs(1762);
    layer2_outputs(465) <= not((layer1_outputs(1874)) and (layer1_outputs(48)));
    layer2_outputs(466) <= (layer1_outputs(1021)) xor (layer1_outputs(439));
    layer2_outputs(467) <= layer1_outputs(2161);
    layer2_outputs(468) <= not(layer1_outputs(1825)) or (layer1_outputs(1013));
    layer2_outputs(469) <= not((layer1_outputs(2487)) xor (layer1_outputs(659)));
    layer2_outputs(470) <= layer1_outputs(893);
    layer2_outputs(471) <= not(layer1_outputs(999));
    layer2_outputs(472) <= not(layer1_outputs(2437));
    layer2_outputs(473) <= not(layer1_outputs(1288));
    layer2_outputs(474) <= layer1_outputs(1648);
    layer2_outputs(475) <= layer1_outputs(515);
    layer2_outputs(476) <= layer1_outputs(696);
    layer2_outputs(477) <= not((layer1_outputs(2269)) and (layer1_outputs(2352)));
    layer2_outputs(478) <= layer1_outputs(1366);
    layer2_outputs(479) <= layer1_outputs(2049);
    layer2_outputs(480) <= layer1_outputs(2021);
    layer2_outputs(481) <= not(layer1_outputs(773));
    layer2_outputs(482) <= (layer1_outputs(395)) xor (layer1_outputs(466));
    layer2_outputs(483) <= not(layer1_outputs(1039)) or (layer1_outputs(1921));
    layer2_outputs(484) <= not(layer1_outputs(77));
    layer2_outputs(485) <= '1';
    layer2_outputs(486) <= layer1_outputs(259);
    layer2_outputs(487) <= not(layer1_outputs(1456));
    layer2_outputs(488) <= (layer1_outputs(503)) and not (layer1_outputs(250));
    layer2_outputs(489) <= (layer1_outputs(1608)) and (layer1_outputs(1321));
    layer2_outputs(490) <= layer1_outputs(2292);
    layer2_outputs(491) <= not(layer1_outputs(410));
    layer2_outputs(492) <= layer1_outputs(1791);
    layer2_outputs(493) <= (layer1_outputs(1360)) and not (layer1_outputs(485));
    layer2_outputs(494) <= not(layer1_outputs(979));
    layer2_outputs(495) <= layer1_outputs(235);
    layer2_outputs(496) <= (layer1_outputs(1932)) and not (layer1_outputs(958));
    layer2_outputs(497) <= not(layer1_outputs(2025)) or (layer1_outputs(660));
    layer2_outputs(498) <= not((layer1_outputs(695)) or (layer1_outputs(120)));
    layer2_outputs(499) <= not(layer1_outputs(130)) or (layer1_outputs(1481));
    layer2_outputs(500) <= not((layer1_outputs(326)) or (layer1_outputs(538)));
    layer2_outputs(501) <= not(layer1_outputs(1800)) or (layer1_outputs(2356));
    layer2_outputs(502) <= layer1_outputs(2482);
    layer2_outputs(503) <= not(layer1_outputs(2028)) or (layer1_outputs(742));
    layer2_outputs(504) <= not(layer1_outputs(2270)) or (layer1_outputs(885));
    layer2_outputs(505) <= (layer1_outputs(1864)) and not (layer1_outputs(630));
    layer2_outputs(506) <= not((layer1_outputs(1118)) or (layer1_outputs(2547)));
    layer2_outputs(507) <= not(layer1_outputs(754));
    layer2_outputs(508) <= layer1_outputs(1849);
    layer2_outputs(509) <= (layer1_outputs(643)) and not (layer1_outputs(2022));
    layer2_outputs(510) <= layer1_outputs(501);
    layer2_outputs(511) <= not((layer1_outputs(610)) and (layer1_outputs(2449)));
    layer2_outputs(512) <= layer1_outputs(1920);
    layer2_outputs(513) <= (layer1_outputs(1)) and not (layer1_outputs(878));
    layer2_outputs(514) <= not((layer1_outputs(1174)) xor (layer1_outputs(2360)));
    layer2_outputs(515) <= layer1_outputs(2546);
    layer2_outputs(516) <= not(layer1_outputs(1771));
    layer2_outputs(517) <= not(layer1_outputs(1043));
    layer2_outputs(518) <= layer1_outputs(1554);
    layer2_outputs(519) <= (layer1_outputs(2515)) or (layer1_outputs(2336));
    layer2_outputs(520) <= '0';
    layer2_outputs(521) <= '1';
    layer2_outputs(522) <= layer1_outputs(1696);
    layer2_outputs(523) <= not(layer1_outputs(2144)) or (layer1_outputs(2192));
    layer2_outputs(524) <= not(layer1_outputs(1143));
    layer2_outputs(525) <= layer1_outputs(2432);
    layer2_outputs(526) <= (layer1_outputs(847)) and (layer1_outputs(918));
    layer2_outputs(527) <= not((layer1_outputs(1475)) or (layer1_outputs(1421)));
    layer2_outputs(528) <= (layer1_outputs(2555)) or (layer1_outputs(1104));
    layer2_outputs(529) <= not((layer1_outputs(1756)) and (layer1_outputs(2397)));
    layer2_outputs(530) <= not(layer1_outputs(493));
    layer2_outputs(531) <= (layer1_outputs(155)) or (layer1_outputs(467));
    layer2_outputs(532) <= layer1_outputs(965);
    layer2_outputs(533) <= not(layer1_outputs(1968));
    layer2_outputs(534) <= (layer1_outputs(1465)) and not (layer1_outputs(1901));
    layer2_outputs(535) <= layer1_outputs(2348);
    layer2_outputs(536) <= layer1_outputs(504);
    layer2_outputs(537) <= (layer1_outputs(518)) and not (layer1_outputs(758));
    layer2_outputs(538) <= layer1_outputs(1344);
    layer2_outputs(539) <= not(layer1_outputs(224)) or (layer1_outputs(1759));
    layer2_outputs(540) <= '1';
    layer2_outputs(541) <= layer1_outputs(2073);
    layer2_outputs(542) <= (layer1_outputs(1401)) and not (layer1_outputs(878));
    layer2_outputs(543) <= layer1_outputs(1940);
    layer2_outputs(544) <= not(layer1_outputs(446));
    layer2_outputs(545) <= layer1_outputs(2398);
    layer2_outputs(546) <= not(layer1_outputs(1766));
    layer2_outputs(547) <= not((layer1_outputs(1014)) and (layer1_outputs(810)));
    layer2_outputs(548) <= layer1_outputs(1854);
    layer2_outputs(549) <= not(layer1_outputs(1615));
    layer2_outputs(550) <= not((layer1_outputs(1191)) or (layer1_outputs(2374)));
    layer2_outputs(551) <= layer1_outputs(289);
    layer2_outputs(552) <= '0';
    layer2_outputs(553) <= (layer1_outputs(2248)) and (layer1_outputs(1568));
    layer2_outputs(554) <= layer1_outputs(2347);
    layer2_outputs(555) <= not(layer1_outputs(698));
    layer2_outputs(556) <= not((layer1_outputs(8)) and (layer1_outputs(192)));
    layer2_outputs(557) <= layer1_outputs(2508);
    layer2_outputs(558) <= layer1_outputs(2312);
    layer2_outputs(559) <= not(layer1_outputs(2363));
    layer2_outputs(560) <= layer1_outputs(851);
    layer2_outputs(561) <= not(layer1_outputs(1585));
    layer2_outputs(562) <= not(layer1_outputs(743));
    layer2_outputs(563) <= '1';
    layer2_outputs(564) <= not(layer1_outputs(2174)) or (layer1_outputs(1446));
    layer2_outputs(565) <= not(layer1_outputs(268));
    layer2_outputs(566) <= not(layer1_outputs(1710));
    layer2_outputs(567) <= (layer1_outputs(1139)) and not (layer1_outputs(1008));
    layer2_outputs(568) <= (layer1_outputs(990)) and not (layer1_outputs(1048));
    layer2_outputs(569) <= not(layer1_outputs(207));
    layer2_outputs(570) <= layer1_outputs(2109);
    layer2_outputs(571) <= not((layer1_outputs(2499)) and (layer1_outputs(118)));
    layer2_outputs(572) <= (layer1_outputs(1113)) xor (layer1_outputs(589));
    layer2_outputs(573) <= not(layer1_outputs(189));
    layer2_outputs(574) <= '1';
    layer2_outputs(575) <= not((layer1_outputs(775)) xor (layer1_outputs(1689)));
    layer2_outputs(576) <= not(layer1_outputs(393));
    layer2_outputs(577) <= layer1_outputs(2164);
    layer2_outputs(578) <= (layer1_outputs(662)) and (layer1_outputs(2155));
    layer2_outputs(579) <= not(layer1_outputs(2302)) or (layer1_outputs(1311));
    layer2_outputs(580) <= layer1_outputs(222);
    layer2_outputs(581) <= layer1_outputs(745);
    layer2_outputs(582) <= layer1_outputs(1271);
    layer2_outputs(583) <= layer1_outputs(195);
    layer2_outputs(584) <= (layer1_outputs(441)) and not (layer1_outputs(524));
    layer2_outputs(585) <= not(layer1_outputs(204));
    layer2_outputs(586) <= not(layer1_outputs(583));
    layer2_outputs(587) <= layer1_outputs(1429);
    layer2_outputs(588) <= layer1_outputs(2418);
    layer2_outputs(589) <= not(layer1_outputs(741));
    layer2_outputs(590) <= not((layer1_outputs(1886)) and (layer1_outputs(348)));
    layer2_outputs(591) <= not(layer1_outputs(528));
    layer2_outputs(592) <= layer1_outputs(247);
    layer2_outputs(593) <= (layer1_outputs(974)) and (layer1_outputs(919));
    layer2_outputs(594) <= not(layer1_outputs(66));
    layer2_outputs(595) <= not(layer1_outputs(1912)) or (layer1_outputs(184));
    layer2_outputs(596) <= (layer1_outputs(469)) xor (layer1_outputs(2160));
    layer2_outputs(597) <= (layer1_outputs(1148)) and (layer1_outputs(2140));
    layer2_outputs(598) <= layer1_outputs(1070);
    layer2_outputs(599) <= not((layer1_outputs(67)) and (layer1_outputs(246)));
    layer2_outputs(600) <= layer1_outputs(1581);
    layer2_outputs(601) <= layer1_outputs(2416);
    layer2_outputs(602) <= not((layer1_outputs(168)) and (layer1_outputs(1808)));
    layer2_outputs(603) <= (layer1_outputs(1280)) and (layer1_outputs(1803));
    layer2_outputs(604) <= not(layer1_outputs(1639));
    layer2_outputs(605) <= not((layer1_outputs(1805)) xor (layer1_outputs(2421)));
    layer2_outputs(606) <= not(layer1_outputs(1483));
    layer2_outputs(607) <= (layer1_outputs(2340)) and not (layer1_outputs(612));
    layer2_outputs(608) <= not(layer1_outputs(203));
    layer2_outputs(609) <= not((layer1_outputs(827)) and (layer1_outputs(1732)));
    layer2_outputs(610) <= not(layer1_outputs(221));
    layer2_outputs(611) <= not(layer1_outputs(1875));
    layer2_outputs(612) <= not(layer1_outputs(871));
    layer2_outputs(613) <= not(layer1_outputs(441));
    layer2_outputs(614) <= not(layer1_outputs(279));
    layer2_outputs(615) <= not(layer1_outputs(113));
    layer2_outputs(616) <= not(layer1_outputs(1021));
    layer2_outputs(617) <= layer1_outputs(2055);
    layer2_outputs(618) <= (layer1_outputs(2103)) or (layer1_outputs(195));
    layer2_outputs(619) <= not(layer1_outputs(2430)) or (layer1_outputs(241));
    layer2_outputs(620) <= not((layer1_outputs(924)) or (layer1_outputs(300)));
    layer2_outputs(621) <= not(layer1_outputs(1821));
    layer2_outputs(622) <= not(layer1_outputs(1778));
    layer2_outputs(623) <= (layer1_outputs(1065)) and (layer1_outputs(2189));
    layer2_outputs(624) <= layer1_outputs(1053);
    layer2_outputs(625) <= not(layer1_outputs(137));
    layer2_outputs(626) <= layer1_outputs(1076);
    layer2_outputs(627) <= not(layer1_outputs(2553));
    layer2_outputs(628) <= not((layer1_outputs(2441)) and (layer1_outputs(1519)));
    layer2_outputs(629) <= layer1_outputs(385);
    layer2_outputs(630) <= not(layer1_outputs(1039));
    layer2_outputs(631) <= not((layer1_outputs(2484)) or (layer1_outputs(172)));
    layer2_outputs(632) <= (layer1_outputs(1579)) and (layer1_outputs(1588));
    layer2_outputs(633) <= not((layer1_outputs(1529)) or (layer1_outputs(2054)));
    layer2_outputs(634) <= (layer1_outputs(337)) or (layer1_outputs(1893));
    layer2_outputs(635) <= (layer1_outputs(43)) and not (layer1_outputs(1786));
    layer2_outputs(636) <= not((layer1_outputs(2136)) xor (layer1_outputs(1306)));
    layer2_outputs(637) <= layer1_outputs(2014);
    layer2_outputs(638) <= layer1_outputs(1477);
    layer2_outputs(639) <= not(layer1_outputs(2041));
    layer2_outputs(640) <= not(layer1_outputs(2309));
    layer2_outputs(641) <= not(layer1_outputs(1643)) or (layer1_outputs(1824));
    layer2_outputs(642) <= not(layer1_outputs(2494)) or (layer1_outputs(1589));
    layer2_outputs(643) <= (layer1_outputs(1104)) and not (layer1_outputs(1900));
    layer2_outputs(644) <= (layer1_outputs(2355)) and (layer1_outputs(1795));
    layer2_outputs(645) <= not(layer1_outputs(2176));
    layer2_outputs(646) <= layer1_outputs(2166);
    layer2_outputs(647) <= not(layer1_outputs(748));
    layer2_outputs(648) <= (layer1_outputs(1085)) xor (layer1_outputs(2391));
    layer2_outputs(649) <= not(layer1_outputs(1868));
    layer2_outputs(650) <= not(layer1_outputs(2300)) or (layer1_outputs(209));
    layer2_outputs(651) <= not(layer1_outputs(1827));
    layer2_outputs(652) <= not((layer1_outputs(581)) and (layer1_outputs(1914)));
    layer2_outputs(653) <= (layer1_outputs(189)) or (layer1_outputs(224));
    layer2_outputs(654) <= (layer1_outputs(794)) or (layer1_outputs(191));
    layer2_outputs(655) <= '0';
    layer2_outputs(656) <= not((layer1_outputs(2419)) and (layer1_outputs(2556)));
    layer2_outputs(657) <= not((layer1_outputs(547)) xor (layer1_outputs(1866)));
    layer2_outputs(658) <= not(layer1_outputs(2468)) or (layer1_outputs(557));
    layer2_outputs(659) <= layer1_outputs(1631);
    layer2_outputs(660) <= '1';
    layer2_outputs(661) <= layer1_outputs(1618);
    layer2_outputs(662) <= layer1_outputs(1558);
    layer2_outputs(663) <= not(layer1_outputs(1274));
    layer2_outputs(664) <= not((layer1_outputs(2452)) and (layer1_outputs(1452)));
    layer2_outputs(665) <= layer1_outputs(645);
    layer2_outputs(666) <= layer1_outputs(1028);
    layer2_outputs(667) <= not(layer1_outputs(1473)) or (layer1_outputs(1802));
    layer2_outputs(668) <= not(layer1_outputs(1180)) or (layer1_outputs(334));
    layer2_outputs(669) <= '0';
    layer2_outputs(670) <= not(layer1_outputs(2292));
    layer2_outputs(671) <= not(layer1_outputs(299));
    layer2_outputs(672) <= layer1_outputs(1649);
    layer2_outputs(673) <= not(layer1_outputs(356));
    layer2_outputs(674) <= not(layer1_outputs(124));
    layer2_outputs(675) <= not(layer1_outputs(174));
    layer2_outputs(676) <= (layer1_outputs(173)) xor (layer1_outputs(2256));
    layer2_outputs(677) <= not((layer1_outputs(492)) and (layer1_outputs(737)));
    layer2_outputs(678) <= layer1_outputs(2415);
    layer2_outputs(679) <= not(layer1_outputs(2275));
    layer2_outputs(680) <= '1';
    layer2_outputs(681) <= layer1_outputs(1761);
    layer2_outputs(682) <= (layer1_outputs(1607)) and (layer1_outputs(2434));
    layer2_outputs(683) <= layer1_outputs(301);
    layer2_outputs(684) <= layer1_outputs(629);
    layer2_outputs(685) <= layer1_outputs(1997);
    layer2_outputs(686) <= not(layer1_outputs(2383));
    layer2_outputs(687) <= not(layer1_outputs(1241));
    layer2_outputs(688) <= not((layer1_outputs(728)) and (layer1_outputs(1086)));
    layer2_outputs(689) <= '1';
    layer2_outputs(690) <= not(layer1_outputs(1102));
    layer2_outputs(691) <= not(layer1_outputs(2030));
    layer2_outputs(692) <= not(layer1_outputs(1093));
    layer2_outputs(693) <= (layer1_outputs(1517)) xor (layer1_outputs(2550));
    layer2_outputs(694) <= not((layer1_outputs(1464)) and (layer1_outputs(535)));
    layer2_outputs(695) <= layer1_outputs(1401);
    layer2_outputs(696) <= layer1_outputs(2512);
    layer2_outputs(697) <= not(layer1_outputs(1042)) or (layer1_outputs(1047));
    layer2_outputs(698) <= layer1_outputs(2165);
    layer2_outputs(699) <= not(layer1_outputs(874)) or (layer1_outputs(1805));
    layer2_outputs(700) <= not((layer1_outputs(198)) and (layer1_outputs(894)));
    layer2_outputs(701) <= layer1_outputs(2485);
    layer2_outputs(702) <= not(layer1_outputs(1195)) or (layer1_outputs(352));
    layer2_outputs(703) <= not((layer1_outputs(2041)) and (layer1_outputs(154)));
    layer2_outputs(704) <= layer1_outputs(89);
    layer2_outputs(705) <= (layer1_outputs(1865)) and (layer1_outputs(1705));
    layer2_outputs(706) <= '0';
    layer2_outputs(707) <= not(layer1_outputs(2321));
    layer2_outputs(708) <= (layer1_outputs(59)) or (layer1_outputs(1358));
    layer2_outputs(709) <= (layer1_outputs(320)) and not (layer1_outputs(925));
    layer2_outputs(710) <= not(layer1_outputs(264)) or (layer1_outputs(1972));
    layer2_outputs(711) <= not(layer1_outputs(153)) or (layer1_outputs(2005));
    layer2_outputs(712) <= (layer1_outputs(1158)) and not (layer1_outputs(911));
    layer2_outputs(713) <= not(layer1_outputs(2419));
    layer2_outputs(714) <= layer1_outputs(2389);
    layer2_outputs(715) <= (layer1_outputs(254)) and (layer1_outputs(2257));
    layer2_outputs(716) <= not(layer1_outputs(479));
    layer2_outputs(717) <= not((layer1_outputs(101)) or (layer1_outputs(1644)));
    layer2_outputs(718) <= (layer1_outputs(502)) and not (layer1_outputs(2169));
    layer2_outputs(719) <= not(layer1_outputs(453)) or (layer1_outputs(1754));
    layer2_outputs(720) <= not(layer1_outputs(2335)) or (layer1_outputs(1790));
    layer2_outputs(721) <= layer1_outputs(1004);
    layer2_outputs(722) <= layer1_outputs(2204);
    layer2_outputs(723) <= not((layer1_outputs(712)) or (layer1_outputs(1275)));
    layer2_outputs(724) <= layer1_outputs(794);
    layer2_outputs(725) <= not(layer1_outputs(615));
    layer2_outputs(726) <= not((layer1_outputs(1154)) and (layer1_outputs(1475)));
    layer2_outputs(727) <= layer1_outputs(2500);
    layer2_outputs(728) <= not(layer1_outputs(1223)) or (layer1_outputs(1658));
    layer2_outputs(729) <= layer1_outputs(1247);
    layer2_outputs(730) <= layer1_outputs(160);
    layer2_outputs(731) <= '0';
    layer2_outputs(732) <= not(layer1_outputs(1511));
    layer2_outputs(733) <= not(layer1_outputs(369));
    layer2_outputs(734) <= not(layer1_outputs(580)) or (layer1_outputs(425));
    layer2_outputs(735) <= (layer1_outputs(1878)) and not (layer1_outputs(2083));
    layer2_outputs(736) <= not(layer1_outputs(466));
    layer2_outputs(737) <= not((layer1_outputs(372)) or (layer1_outputs(1017)));
    layer2_outputs(738) <= not(layer1_outputs(123));
    layer2_outputs(739) <= layer1_outputs(1715);
    layer2_outputs(740) <= not((layer1_outputs(2471)) and (layer1_outputs(904)));
    layer2_outputs(741) <= not((layer1_outputs(1527)) and (layer1_outputs(417)));
    layer2_outputs(742) <= not((layer1_outputs(2061)) and (layer1_outputs(81)));
    layer2_outputs(743) <= layer1_outputs(856);
    layer2_outputs(744) <= not(layer1_outputs(630));
    layer2_outputs(745) <= layer1_outputs(779);
    layer2_outputs(746) <= not(layer1_outputs(74));
    layer2_outputs(747) <= not(layer1_outputs(902));
    layer2_outputs(748) <= not(layer1_outputs(1694));
    layer2_outputs(749) <= (layer1_outputs(1410)) xor (layer1_outputs(1522));
    layer2_outputs(750) <= not((layer1_outputs(2122)) or (layer1_outputs(1359)));
    layer2_outputs(751) <= '0';
    layer2_outputs(752) <= layer1_outputs(591);
    layer2_outputs(753) <= layer1_outputs(1726);
    layer2_outputs(754) <= (layer1_outputs(1541)) xor (layer1_outputs(2209));
    layer2_outputs(755) <= not(layer1_outputs(1203));
    layer2_outputs(756) <= not(layer1_outputs(1981)) or (layer1_outputs(264));
    layer2_outputs(757) <= not((layer1_outputs(2317)) and (layer1_outputs(1324)));
    layer2_outputs(758) <= (layer1_outputs(2544)) and not (layer1_outputs(935));
    layer2_outputs(759) <= layer1_outputs(202);
    layer2_outputs(760) <= not((layer1_outputs(168)) or (layer1_outputs(1381)));
    layer2_outputs(761) <= not((layer1_outputs(672)) or (layer1_outputs(1398)));
    layer2_outputs(762) <= layer1_outputs(194);
    layer2_outputs(763) <= not(layer1_outputs(845));
    layer2_outputs(764) <= not(layer1_outputs(1162));
    layer2_outputs(765) <= not((layer1_outputs(1414)) or (layer1_outputs(104)));
    layer2_outputs(766) <= (layer1_outputs(1980)) or (layer1_outputs(1596));
    layer2_outputs(767) <= not(layer1_outputs(864));
    layer2_outputs(768) <= layer1_outputs(673);
    layer2_outputs(769) <= (layer1_outputs(857)) or (layer1_outputs(1573));
    layer2_outputs(770) <= not(layer1_outputs(1408)) or (layer1_outputs(1470));
    layer2_outputs(771) <= not(layer1_outputs(327));
    layer2_outputs(772) <= (layer1_outputs(2237)) and (layer1_outputs(1308));
    layer2_outputs(773) <= not((layer1_outputs(1770)) and (layer1_outputs(2184)));
    layer2_outputs(774) <= (layer1_outputs(1230)) and (layer1_outputs(862));
    layer2_outputs(775) <= not((layer1_outputs(1961)) and (layer1_outputs(993)));
    layer2_outputs(776) <= (layer1_outputs(975)) and not (layer1_outputs(41));
    layer2_outputs(777) <= not(layer1_outputs(1637));
    layer2_outputs(778) <= layer1_outputs(1113);
    layer2_outputs(779) <= not(layer1_outputs(2450));
    layer2_outputs(780) <= not(layer1_outputs(1116));
    layer2_outputs(781) <= (layer1_outputs(1965)) or (layer1_outputs(2260));
    layer2_outputs(782) <= not(layer1_outputs(2341));
    layer2_outputs(783) <= (layer1_outputs(1520)) and (layer1_outputs(1529));
    layer2_outputs(784) <= '0';
    layer2_outputs(785) <= layer1_outputs(605);
    layer2_outputs(786) <= not(layer1_outputs(561)) or (layer1_outputs(1802));
    layer2_outputs(787) <= not((layer1_outputs(1682)) or (layer1_outputs(949)));
    layer2_outputs(788) <= (layer1_outputs(156)) and not (layer1_outputs(275));
    layer2_outputs(789) <= (layer1_outputs(676)) and (layer1_outputs(1876));
    layer2_outputs(790) <= not(layer1_outputs(575));
    layer2_outputs(791) <= (layer1_outputs(1978)) and not (layer1_outputs(2304));
    layer2_outputs(792) <= (layer1_outputs(1762)) and (layer1_outputs(409));
    layer2_outputs(793) <= layer1_outputs(208);
    layer2_outputs(794) <= layer1_outputs(2120);
    layer2_outputs(795) <= not(layer1_outputs(336)) or (layer1_outputs(1804));
    layer2_outputs(796) <= not(layer1_outputs(2333));
    layer2_outputs(797) <= (layer1_outputs(552)) and not (layer1_outputs(681));
    layer2_outputs(798) <= not(layer1_outputs(894)) or (layer1_outputs(1267));
    layer2_outputs(799) <= (layer1_outputs(39)) or (layer1_outputs(21));
    layer2_outputs(800) <= '1';
    layer2_outputs(801) <= not(layer1_outputs(936));
    layer2_outputs(802) <= not(layer1_outputs(2173));
    layer2_outputs(803) <= (layer1_outputs(1652)) and not (layer1_outputs(408));
    layer2_outputs(804) <= layer1_outputs(2146);
    layer2_outputs(805) <= not(layer1_outputs(2353));
    layer2_outputs(806) <= (layer1_outputs(437)) or (layer1_outputs(691));
    layer2_outputs(807) <= not((layer1_outputs(1717)) or (layer1_outputs(1289)));
    layer2_outputs(808) <= (layer1_outputs(1673)) and not (layer1_outputs(1491));
    layer2_outputs(809) <= layer1_outputs(604);
    layer2_outputs(810) <= (layer1_outputs(869)) or (layer1_outputs(1211));
    layer2_outputs(811) <= layer1_outputs(2065);
    layer2_outputs(812) <= not((layer1_outputs(1284)) and (layer1_outputs(1778)));
    layer2_outputs(813) <= layer1_outputs(1651);
    layer2_outputs(814) <= not((layer1_outputs(1173)) or (layer1_outputs(703)));
    layer2_outputs(815) <= layer1_outputs(1626);
    layer2_outputs(816) <= not(layer1_outputs(1568)) or (layer1_outputs(1413));
    layer2_outputs(817) <= not(layer1_outputs(2219));
    layer2_outputs(818) <= (layer1_outputs(505)) and (layer1_outputs(1686));
    layer2_outputs(819) <= not(layer1_outputs(1480));
    layer2_outputs(820) <= (layer1_outputs(1055)) and not (layer1_outputs(1751));
    layer2_outputs(821) <= (layer1_outputs(1019)) and not (layer1_outputs(1578));
    layer2_outputs(822) <= not(layer1_outputs(728)) or (layer1_outputs(2012));
    layer2_outputs(823) <= not(layer1_outputs(1941));
    layer2_outputs(824) <= not(layer1_outputs(1781)) or (layer1_outputs(2235));
    layer2_outputs(825) <= not(layer1_outputs(2096));
    layer2_outputs(826) <= (layer1_outputs(1236)) and (layer1_outputs(2217));
    layer2_outputs(827) <= (layer1_outputs(1445)) and (layer1_outputs(643));
    layer2_outputs(828) <= not(layer1_outputs(1580)) or (layer1_outputs(1612));
    layer2_outputs(829) <= not(layer1_outputs(770)) or (layer1_outputs(2389));
    layer2_outputs(830) <= not(layer1_outputs(1314));
    layer2_outputs(831) <= layer1_outputs(1934);
    layer2_outputs(832) <= (layer1_outputs(1855)) and not (layer1_outputs(2536));
    layer2_outputs(833) <= not((layer1_outputs(2036)) and (layer1_outputs(666)));
    layer2_outputs(834) <= (layer1_outputs(1867)) and not (layer1_outputs(2267));
    layer2_outputs(835) <= (layer1_outputs(1404)) and (layer1_outputs(1341));
    layer2_outputs(836) <= not(layer1_outputs(1601));
    layer2_outputs(837) <= (layer1_outputs(1374)) and (layer1_outputs(1535));
    layer2_outputs(838) <= (layer1_outputs(1177)) and not (layer1_outputs(2129));
    layer2_outputs(839) <= not(layer1_outputs(689)) or (layer1_outputs(1238));
    layer2_outputs(840) <= layer1_outputs(2134);
    layer2_outputs(841) <= not(layer1_outputs(2453));
    layer2_outputs(842) <= not(layer1_outputs(1695));
    layer2_outputs(843) <= layer1_outputs(1406);
    layer2_outputs(844) <= layer1_outputs(1587);
    layer2_outputs(845) <= not(layer1_outputs(511));
    layer2_outputs(846) <= '0';
    layer2_outputs(847) <= layer1_outputs(234);
    layer2_outputs(848) <= layer1_outputs(94);
    layer2_outputs(849) <= layer1_outputs(776);
    layer2_outputs(850) <= layer1_outputs(2529);
    layer2_outputs(851) <= (layer1_outputs(521)) and (layer1_outputs(450));
    layer2_outputs(852) <= not(layer1_outputs(632));
    layer2_outputs(853) <= not(layer1_outputs(1147));
    layer2_outputs(854) <= (layer1_outputs(387)) and (layer1_outputs(2469));
    layer2_outputs(855) <= (layer1_outputs(2121)) or (layer1_outputs(1836));
    layer2_outputs(856) <= not(layer1_outputs(1369)) or (layer1_outputs(2260));
    layer2_outputs(857) <= not((layer1_outputs(1176)) and (layer1_outputs(2089)));
    layer2_outputs(858) <= '0';
    layer2_outputs(859) <= (layer1_outputs(752)) and not (layer1_outputs(2370));
    layer2_outputs(860) <= not(layer1_outputs(2051)) or (layer1_outputs(107));
    layer2_outputs(861) <= not(layer1_outputs(1943)) or (layer1_outputs(1111));
    layer2_outputs(862) <= layer1_outputs(2046);
    layer2_outputs(863) <= '0';
    layer2_outputs(864) <= layer1_outputs(236);
    layer2_outputs(865) <= (layer1_outputs(1627)) and (layer1_outputs(1626));
    layer2_outputs(866) <= layer1_outputs(1859);
    layer2_outputs(867) <= not(layer1_outputs(1119));
    layer2_outputs(868) <= (layer1_outputs(2105)) and (layer1_outputs(2537));
    layer2_outputs(869) <= (layer1_outputs(2416)) and (layer1_outputs(1417));
    layer2_outputs(870) <= layer1_outputs(1559);
    layer2_outputs(871) <= layer1_outputs(1107);
    layer2_outputs(872) <= not(layer1_outputs(650));
    layer2_outputs(873) <= layer1_outputs(2124);
    layer2_outputs(874) <= (layer1_outputs(2284)) and not (layer1_outputs(55));
    layer2_outputs(875) <= layer1_outputs(1690);
    layer2_outputs(876) <= not(layer1_outputs(1598));
    layer2_outputs(877) <= (layer1_outputs(1029)) and (layer1_outputs(2380));
    layer2_outputs(878) <= (layer1_outputs(835)) xor (layer1_outputs(73));
    layer2_outputs(879) <= (layer1_outputs(1647)) or (layer1_outputs(2291));
    layer2_outputs(880) <= layer1_outputs(254);
    layer2_outputs(881) <= not(layer1_outputs(295));
    layer2_outputs(882) <= (layer1_outputs(110)) or (layer1_outputs(1666));
    layer2_outputs(883) <= layer1_outputs(653);
    layer2_outputs(884) <= (layer1_outputs(870)) and not (layer1_outputs(1054));
    layer2_outputs(885) <= not(layer1_outputs(54)) or (layer1_outputs(2278));
    layer2_outputs(886) <= not(layer1_outputs(2005));
    layer2_outputs(887) <= (layer1_outputs(985)) and (layer1_outputs(1208));
    layer2_outputs(888) <= '0';
    layer2_outputs(889) <= not(layer1_outputs(1594)) or (layer1_outputs(1850));
    layer2_outputs(890) <= layer1_outputs(883);
    layer2_outputs(891) <= (layer1_outputs(1417)) or (layer1_outputs(718));
    layer2_outputs(892) <= not((layer1_outputs(1430)) and (layer1_outputs(2433)));
    layer2_outputs(893) <= not(layer1_outputs(1552)) or (layer1_outputs(613));
    layer2_outputs(894) <= not(layer1_outputs(861));
    layer2_outputs(895) <= not(layer1_outputs(740));
    layer2_outputs(896) <= not(layer1_outputs(1061));
    layer2_outputs(897) <= (layer1_outputs(406)) and not (layer1_outputs(994));
    layer2_outputs(898) <= layer1_outputs(740);
    layer2_outputs(899) <= layer1_outputs(2488);
    layer2_outputs(900) <= (layer1_outputs(1845)) and (layer1_outputs(397));
    layer2_outputs(901) <= not(layer1_outputs(1622)) or (layer1_outputs(1651));
    layer2_outputs(902) <= (layer1_outputs(122)) and not (layer1_outputs(1202));
    layer2_outputs(903) <= layer1_outputs(331);
    layer2_outputs(904) <= not(layer1_outputs(1793));
    layer2_outputs(905) <= not(layer1_outputs(1112)) or (layer1_outputs(1910));
    layer2_outputs(906) <= not(layer1_outputs(1788));
    layer2_outputs(907) <= layer1_outputs(2168);
    layer2_outputs(908) <= (layer1_outputs(1771)) and (layer1_outputs(912));
    layer2_outputs(909) <= (layer1_outputs(196)) and not (layer1_outputs(208));
    layer2_outputs(910) <= (layer1_outputs(452)) xor (layer1_outputs(1435));
    layer2_outputs(911) <= not(layer1_outputs(2194));
    layer2_outputs(912) <= not(layer1_outputs(1245));
    layer2_outputs(913) <= (layer1_outputs(829)) or (layer1_outputs(1484));
    layer2_outputs(914) <= layer1_outputs(1336);
    layer2_outputs(915) <= '0';
    layer2_outputs(916) <= layer1_outputs(2017);
    layer2_outputs(917) <= not(layer1_outputs(304));
    layer2_outputs(918) <= layer1_outputs(756);
    layer2_outputs(919) <= not(layer1_outputs(1111));
    layer2_outputs(920) <= not((layer1_outputs(353)) and (layer1_outputs(1613)));
    layer2_outputs(921) <= (layer1_outputs(1458)) and (layer1_outputs(1050));
    layer2_outputs(922) <= (layer1_outputs(368)) and (layer1_outputs(1250));
    layer2_outputs(923) <= not(layer1_outputs(555)) or (layer1_outputs(1003));
    layer2_outputs(924) <= '1';
    layer2_outputs(925) <= layer1_outputs(1296);
    layer2_outputs(926) <= not(layer1_outputs(2101));
    layer2_outputs(927) <= (layer1_outputs(640)) or (layer1_outputs(1498));
    layer2_outputs(928) <= (layer1_outputs(927)) or (layer1_outputs(2097));
    layer2_outputs(929) <= (layer1_outputs(887)) and not (layer1_outputs(597));
    layer2_outputs(930) <= not((layer1_outputs(1524)) or (layer1_outputs(664)));
    layer2_outputs(931) <= not((layer1_outputs(124)) and (layer1_outputs(1135)));
    layer2_outputs(932) <= (layer1_outputs(1106)) or (layer1_outputs(1966));
    layer2_outputs(933) <= layer1_outputs(1175);
    layer2_outputs(934) <= layer1_outputs(2505);
    layer2_outputs(935) <= not((layer1_outputs(2079)) or (layer1_outputs(1604)));
    layer2_outputs(936) <= (layer1_outputs(1010)) and not (layer1_outputs(513));
    layer2_outputs(937) <= (layer1_outputs(416)) or (layer1_outputs(2071));
    layer2_outputs(938) <= (layer1_outputs(121)) and not (layer1_outputs(1203));
    layer2_outputs(939) <= not((layer1_outputs(822)) xor (layer1_outputs(233)));
    layer2_outputs(940) <= not(layer1_outputs(717)) or (layer1_outputs(601));
    layer2_outputs(941) <= not((layer1_outputs(2382)) and (layer1_outputs(1659)));
    layer2_outputs(942) <= not((layer1_outputs(2337)) and (layer1_outputs(796)));
    layer2_outputs(943) <= layer1_outputs(1948);
    layer2_outputs(944) <= not(layer1_outputs(2151)) or (layer1_outputs(1479));
    layer2_outputs(945) <= not(layer1_outputs(1751));
    layer2_outputs(946) <= layer1_outputs(2096);
    layer2_outputs(947) <= (layer1_outputs(1619)) and not (layer1_outputs(1719));
    layer2_outputs(948) <= not(layer1_outputs(1164));
    layer2_outputs(949) <= not((layer1_outputs(721)) or (layer1_outputs(283)));
    layer2_outputs(950) <= layer1_outputs(628);
    layer2_outputs(951) <= not((layer1_outputs(38)) xor (layer1_outputs(1194)));
    layer2_outputs(952) <= layer1_outputs(578);
    layer2_outputs(953) <= layer1_outputs(68);
    layer2_outputs(954) <= not(layer1_outputs(1584));
    layer2_outputs(955) <= layer1_outputs(1783);
    layer2_outputs(956) <= (layer1_outputs(1511)) and not (layer1_outputs(1434));
    layer2_outputs(957) <= not(layer1_outputs(1230)) or (layer1_outputs(1962));
    layer2_outputs(958) <= not(layer1_outputs(1124));
    layer2_outputs(959) <= not(layer1_outputs(1745));
    layer2_outputs(960) <= not(layer1_outputs(2062)) or (layer1_outputs(708));
    layer2_outputs(961) <= layer1_outputs(561);
    layer2_outputs(962) <= (layer1_outputs(1130)) and not (layer1_outputs(2083));
    layer2_outputs(963) <= layer1_outputs(251);
    layer2_outputs(964) <= not((layer1_outputs(2391)) and (layer1_outputs(588)));
    layer2_outputs(965) <= not(layer1_outputs(1930)) or (layer1_outputs(1574));
    layer2_outputs(966) <= layer1_outputs(1754);
    layer2_outputs(967) <= (layer1_outputs(961)) and not (layer1_outputs(563));
    layer2_outputs(968) <= layer1_outputs(855);
    layer2_outputs(969) <= not((layer1_outputs(333)) and (layer1_outputs(562)));
    layer2_outputs(970) <= not(layer1_outputs(1583));
    layer2_outputs(971) <= not((layer1_outputs(1957)) or (layer1_outputs(2001)));
    layer2_outputs(972) <= layer1_outputs(2305);
    layer2_outputs(973) <= '1';
    layer2_outputs(974) <= layer1_outputs(1454);
    layer2_outputs(975) <= not(layer1_outputs(2469));
    layer2_outputs(976) <= '0';
    layer2_outputs(977) <= layer1_outputs(464);
    layer2_outputs(978) <= not(layer1_outputs(450));
    layer2_outputs(979) <= not(layer1_outputs(1225)) or (layer1_outputs(2452));
    layer2_outputs(980) <= not(layer1_outputs(1588));
    layer2_outputs(981) <= not(layer1_outputs(1797));
    layer2_outputs(982) <= layer1_outputs(247);
    layer2_outputs(983) <= not(layer1_outputs(1890));
    layer2_outputs(984) <= (layer1_outputs(2161)) or (layer1_outputs(432));
    layer2_outputs(985) <= layer1_outputs(639);
    layer2_outputs(986) <= not(layer1_outputs(2206)) or (layer1_outputs(1456));
    layer2_outputs(987) <= (layer1_outputs(1050)) or (layer1_outputs(877));
    layer2_outputs(988) <= not((layer1_outputs(458)) and (layer1_outputs(2510)));
    layer2_outputs(989) <= layer1_outputs(960);
    layer2_outputs(990) <= not(layer1_outputs(2244));
    layer2_outputs(991) <= not(layer1_outputs(1543));
    layer2_outputs(992) <= not(layer1_outputs(2504)) or (layer1_outputs(1319));
    layer2_outputs(993) <= (layer1_outputs(1139)) and not (layer1_outputs(82));
    layer2_outputs(994) <= not(layer1_outputs(747)) or (layer1_outputs(835));
    layer2_outputs(995) <= layer1_outputs(720);
    layer2_outputs(996) <= (layer1_outputs(891)) or (layer1_outputs(1244));
    layer2_outputs(997) <= not(layer1_outputs(427));
    layer2_outputs(998) <= not(layer1_outputs(449)) or (layer1_outputs(120));
    layer2_outputs(999) <= not(layer1_outputs(2162)) or (layer1_outputs(2344));
    layer2_outputs(1000) <= (layer1_outputs(734)) and not (layer1_outputs(2479));
    layer2_outputs(1001) <= not(layer1_outputs(1853));
    layer2_outputs(1002) <= not(layer1_outputs(897));
    layer2_outputs(1003) <= not(layer1_outputs(1128));
    layer2_outputs(1004) <= not(layer1_outputs(1808));
    layer2_outputs(1005) <= layer1_outputs(502);
    layer2_outputs(1006) <= layer1_outputs(2534);
    layer2_outputs(1007) <= (layer1_outputs(1709)) xor (layer1_outputs(1157));
    layer2_outputs(1008) <= layer1_outputs(1069);
    layer2_outputs(1009) <= not(layer1_outputs(1532));
    layer2_outputs(1010) <= not(layer1_outputs(551));
    layer2_outputs(1011) <= layer1_outputs(558);
    layer2_outputs(1012) <= not(layer1_outputs(900));
    layer2_outputs(1013) <= not(layer1_outputs(1334));
    layer2_outputs(1014) <= not((layer1_outputs(2130)) or (layer1_outputs(420)));
    layer2_outputs(1015) <= (layer1_outputs(356)) and (layer1_outputs(1880));
    layer2_outputs(1016) <= layer1_outputs(354);
    layer2_outputs(1017) <= not((layer1_outputs(1281)) and (layer1_outputs(890)));
    layer2_outputs(1018) <= (layer1_outputs(1285)) or (layer1_outputs(127));
    layer2_outputs(1019) <= (layer1_outputs(226)) and not (layer1_outputs(17));
    layer2_outputs(1020) <= not(layer1_outputs(2327)) or (layer1_outputs(1402));
    layer2_outputs(1021) <= not(layer1_outputs(1935));
    layer2_outputs(1022) <= (layer1_outputs(2222)) xor (layer1_outputs(1484));
    layer2_outputs(1023) <= layer1_outputs(1191);
    layer2_outputs(1024) <= not(layer1_outputs(2032)) or (layer1_outputs(2413));
    layer2_outputs(1025) <= layer1_outputs(100);
    layer2_outputs(1026) <= not(layer1_outputs(2339)) or (layer1_outputs(1438));
    layer2_outputs(1027) <= layer1_outputs(8);
    layer2_outputs(1028) <= layer1_outputs(404);
    layer2_outputs(1029) <= not(layer1_outputs(1451));
    layer2_outputs(1030) <= not(layer1_outputs(2345));
    layer2_outputs(1031) <= not(layer1_outputs(315));
    layer2_outputs(1032) <= layer1_outputs(1270);
    layer2_outputs(1033) <= not((layer1_outputs(221)) or (layer1_outputs(2035)));
    layer2_outputs(1034) <= not(layer1_outputs(1018)) or (layer1_outputs(2448));
    layer2_outputs(1035) <= (layer1_outputs(1372)) and (layer1_outputs(863));
    layer2_outputs(1036) <= not((layer1_outputs(981)) or (layer1_outputs(1033)));
    layer2_outputs(1037) <= (layer1_outputs(2)) and not (layer1_outputs(1499));
    layer2_outputs(1038) <= layer1_outputs(2318);
    layer2_outputs(1039) <= not(layer1_outputs(1610));
    layer2_outputs(1040) <= not((layer1_outputs(69)) or (layer1_outputs(731)));
    layer2_outputs(1041) <= not(layer1_outputs(336));
    layer2_outputs(1042) <= layer1_outputs(2250);
    layer2_outputs(1043) <= not(layer1_outputs(1346)) or (layer1_outputs(1603));
    layer2_outputs(1044) <= not(layer1_outputs(1753)) or (layer1_outputs(1033));
    layer2_outputs(1045) <= '1';
    layer2_outputs(1046) <= not((layer1_outputs(320)) or (layer1_outputs(1717)));
    layer2_outputs(1047) <= not(layer1_outputs(2251));
    layer2_outputs(1048) <= (layer1_outputs(2024)) and (layer1_outputs(1605));
    layer2_outputs(1049) <= layer1_outputs(2290);
    layer2_outputs(1050) <= (layer1_outputs(2511)) and not (layer1_outputs(596));
    layer2_outputs(1051) <= layer1_outputs(998);
    layer2_outputs(1052) <= layer1_outputs(1553);
    layer2_outputs(1053) <= not(layer1_outputs(638));
    layer2_outputs(1054) <= not(layer1_outputs(1249));
    layer2_outputs(1055) <= (layer1_outputs(462)) or (layer1_outputs(874));
    layer2_outputs(1056) <= not((layer1_outputs(929)) or (layer1_outputs(2157)));
    layer2_outputs(1057) <= layer1_outputs(1880);
    layer2_outputs(1058) <= not(layer1_outputs(1155)) or (layer1_outputs(1645));
    layer2_outputs(1059) <= layer1_outputs(442);
    layer2_outputs(1060) <= layer1_outputs(1342);
    layer2_outputs(1061) <= not(layer1_outputs(742));
    layer2_outputs(1062) <= layer1_outputs(1923);
    layer2_outputs(1063) <= layer1_outputs(94);
    layer2_outputs(1064) <= not((layer1_outputs(1240)) and (layer1_outputs(1339)));
    layer2_outputs(1065) <= (layer1_outputs(2228)) and not (layer1_outputs(2352));
    layer2_outputs(1066) <= not(layer1_outputs(576));
    layer2_outputs(1067) <= not(layer1_outputs(2007)) or (layer1_outputs(1210));
    layer2_outputs(1068) <= (layer1_outputs(246)) and not (layer1_outputs(1623));
    layer2_outputs(1069) <= not(layer1_outputs(352));
    layer2_outputs(1070) <= layer1_outputs(565);
    layer2_outputs(1071) <= not(layer1_outputs(1672)) or (layer1_outputs(570));
    layer2_outputs(1072) <= layer1_outputs(2558);
    layer2_outputs(1073) <= not((layer1_outputs(1204)) or (layer1_outputs(1216)));
    layer2_outputs(1074) <= '1';
    layer2_outputs(1075) <= not((layer1_outputs(955)) and (layer1_outputs(671)));
    layer2_outputs(1076) <= layer1_outputs(942);
    layer2_outputs(1077) <= layer1_outputs(1788);
    layer2_outputs(1078) <= not((layer1_outputs(1305)) or (layer1_outputs(193)));
    layer2_outputs(1079) <= layer1_outputs(2116);
    layer2_outputs(1080) <= layer1_outputs(67);
    layer2_outputs(1081) <= not(layer1_outputs(186));
    layer2_outputs(1082) <= (layer1_outputs(92)) and (layer1_outputs(72));
    layer2_outputs(1083) <= layer1_outputs(2277);
    layer2_outputs(1084) <= not((layer1_outputs(895)) xor (layer1_outputs(2501)));
    layer2_outputs(1085) <= (layer1_outputs(2238)) or (layer1_outputs(170));
    layer2_outputs(1086) <= not((layer1_outputs(1618)) or (layer1_outputs(3)));
    layer2_outputs(1087) <= (layer1_outputs(1007)) or (layer1_outputs(1952));
    layer2_outputs(1088) <= not(layer1_outputs(1351));
    layer2_outputs(1089) <= layer1_outputs(1340);
    layer2_outputs(1090) <= not((layer1_outputs(916)) and (layer1_outputs(1433)));
    layer2_outputs(1091) <= not(layer1_outputs(1502));
    layer2_outputs(1092) <= not(layer1_outputs(1089));
    layer2_outputs(1093) <= not(layer1_outputs(1224));
    layer2_outputs(1094) <= layer1_outputs(50);
    layer2_outputs(1095) <= '1';
    layer2_outputs(1096) <= not(layer1_outputs(2462));
    layer2_outputs(1097) <= not((layer1_outputs(1812)) or (layer1_outputs(2262)));
    layer2_outputs(1098) <= layer1_outputs(46);
    layer2_outputs(1099) <= layer1_outputs(267);
    layer2_outputs(1100) <= (layer1_outputs(285)) or (layer1_outputs(1826));
    layer2_outputs(1101) <= (layer1_outputs(1831)) and (layer1_outputs(2089));
    layer2_outputs(1102) <= layer1_outputs(1144);
    layer2_outputs(1103) <= layer1_outputs(1920);
    layer2_outputs(1104) <= (layer1_outputs(1352)) and not (layer1_outputs(1376));
    layer2_outputs(1105) <= layer1_outputs(1792);
    layer2_outputs(1106) <= not(layer1_outputs(1017));
    layer2_outputs(1107) <= (layer1_outputs(376)) and (layer1_outputs(402));
    layer2_outputs(1108) <= not(layer1_outputs(782)) or (layer1_outputs(2027));
    layer2_outputs(1109) <= not(layer1_outputs(1711));
    layer2_outputs(1110) <= (layer1_outputs(52)) or (layer1_outputs(2515));
    layer2_outputs(1111) <= not((layer1_outputs(420)) or (layer1_outputs(549)));
    layer2_outputs(1112) <= (layer1_outputs(1985)) xor (layer1_outputs(1046));
    layer2_outputs(1113) <= not(layer1_outputs(1506));
    layer2_outputs(1114) <= not(layer1_outputs(1292)) or (layer1_outputs(111));
    layer2_outputs(1115) <= not(layer1_outputs(1322));
    layer2_outputs(1116) <= not(layer1_outputs(347));
    layer2_outputs(1117) <= not(layer1_outputs(703));
    layer2_outputs(1118) <= layer1_outputs(274);
    layer2_outputs(1119) <= (layer1_outputs(2519)) and not (layer1_outputs(159));
    layer2_outputs(1120) <= '0';
    layer2_outputs(1121) <= not((layer1_outputs(1546)) and (layer1_outputs(609)));
    layer2_outputs(1122) <= not(layer1_outputs(2076));
    layer2_outputs(1123) <= (layer1_outputs(101)) and not (layer1_outputs(2061));
    layer2_outputs(1124) <= not(layer1_outputs(2529)) or (layer1_outputs(1987));
    layer2_outputs(1125) <= not(layer1_outputs(2028));
    layer2_outputs(1126) <= layer1_outputs(2042);
    layer2_outputs(1127) <= not(layer1_outputs(2422));
    layer2_outputs(1128) <= not(layer1_outputs(593));
    layer2_outputs(1129) <= layer1_outputs(525);
    layer2_outputs(1130) <= not(layer1_outputs(2176));
    layer2_outputs(1131) <= layer1_outputs(1160);
    layer2_outputs(1132) <= not(layer1_outputs(1494));
    layer2_outputs(1133) <= not(layer1_outputs(2478)) or (layer1_outputs(138));
    layer2_outputs(1134) <= '0';
    layer2_outputs(1135) <= not(layer1_outputs(1221));
    layer2_outputs(1136) <= not(layer1_outputs(1932));
    layer2_outputs(1137) <= not(layer1_outputs(2033));
    layer2_outputs(1138) <= (layer1_outputs(1833)) xor (layer1_outputs(2338));
    layer2_outputs(1139) <= not((layer1_outputs(163)) and (layer1_outputs(216)));
    layer2_outputs(1140) <= layer1_outputs(343);
    layer2_outputs(1141) <= layer1_outputs(223);
    layer2_outputs(1142) <= not(layer1_outputs(910)) or (layer1_outputs(1597));
    layer2_outputs(1143) <= '0';
    layer2_outputs(1144) <= layer1_outputs(1583);
    layer2_outputs(1145) <= not(layer1_outputs(1189));
    layer2_outputs(1146) <= layer1_outputs(2088);
    layer2_outputs(1147) <= (layer1_outputs(2093)) and not (layer1_outputs(1987));
    layer2_outputs(1148) <= layer1_outputs(1071);
    layer2_outputs(1149) <= (layer1_outputs(1247)) and not (layer1_outputs(2193));
    layer2_outputs(1150) <= not((layer1_outputs(463)) and (layer1_outputs(1032)));
    layer2_outputs(1151) <= layer1_outputs(256);
    layer2_outputs(1152) <= layer1_outputs(1315);
    layer2_outputs(1153) <= not(layer1_outputs(1572));
    layer2_outputs(1154) <= not(layer1_outputs(1307));
    layer2_outputs(1155) <= not(layer1_outputs(828));
    layer2_outputs(1156) <= (layer1_outputs(157)) or (layer1_outputs(1842));
    layer2_outputs(1157) <= layer1_outputs(308);
    layer2_outputs(1158) <= layer1_outputs(718);
    layer2_outputs(1159) <= not(layer1_outputs(2075)) or (layer1_outputs(465));
    layer2_outputs(1160) <= not((layer1_outputs(2143)) or (layer1_outputs(1939)));
    layer2_outputs(1161) <= layer1_outputs(1609);
    layer2_outputs(1162) <= (layer1_outputs(44)) and not (layer1_outputs(1516));
    layer2_outputs(1163) <= not(layer1_outputs(2408));
    layer2_outputs(1164) <= not(layer1_outputs(2325));
    layer2_outputs(1165) <= not((layer1_outputs(2281)) and (layer1_outputs(2055)));
    layer2_outputs(1166) <= (layer1_outputs(1303)) and not (layer1_outputs(1331));
    layer2_outputs(1167) <= (layer1_outputs(558)) and not (layer1_outputs(1387));
    layer2_outputs(1168) <= layer1_outputs(498);
    layer2_outputs(1169) <= not((layer1_outputs(2086)) xor (layer1_outputs(1037)));
    layer2_outputs(1170) <= not((layer1_outputs(1099)) or (layer1_outputs(219)));
    layer2_outputs(1171) <= not(layer1_outputs(789));
    layer2_outputs(1172) <= layer1_outputs(1964);
    layer2_outputs(1173) <= layer1_outputs(587);
    layer2_outputs(1174) <= not((layer1_outputs(1832)) and (layer1_outputs(2368)));
    layer2_outputs(1175) <= not(layer1_outputs(457)) or (layer1_outputs(2125));
    layer2_outputs(1176) <= (layer1_outputs(71)) and not (layer1_outputs(1507));
    layer2_outputs(1177) <= not(layer1_outputs(206));
    layer2_outputs(1178) <= not((layer1_outputs(791)) or (layer1_outputs(768)));
    layer2_outputs(1179) <= layer1_outputs(819);
    layer2_outputs(1180) <= layer1_outputs(2255);
    layer2_outputs(1181) <= not((layer1_outputs(1200)) or (layer1_outputs(292)));
    layer2_outputs(1182) <= not(layer1_outputs(638));
    layer2_outputs(1183) <= layer1_outputs(1198);
    layer2_outputs(1184) <= not(layer1_outputs(1332));
    layer2_outputs(1185) <= layer1_outputs(1973);
    layer2_outputs(1186) <= not(layer1_outputs(227));
    layer2_outputs(1187) <= layer1_outputs(842);
    layer2_outputs(1188) <= not(layer1_outputs(2205));
    layer2_outputs(1189) <= layer1_outputs(609);
    layer2_outputs(1190) <= not(layer1_outputs(1287));
    layer2_outputs(1191) <= not(layer1_outputs(1852));
    layer2_outputs(1192) <= layer1_outputs(786);
    layer2_outputs(1193) <= layer1_outputs(1826);
    layer2_outputs(1194) <= not((layer1_outputs(1706)) and (layer1_outputs(966)));
    layer2_outputs(1195) <= layer1_outputs(719);
    layer2_outputs(1196) <= '1';
    layer2_outputs(1197) <= layer1_outputs(1379);
    layer2_outputs(1198) <= not(layer1_outputs(553)) or (layer1_outputs(2203));
    layer2_outputs(1199) <= layer1_outputs(1841);
    layer2_outputs(1200) <= not(layer1_outputs(1577));
    layer2_outputs(1201) <= (layer1_outputs(1776)) and (layer1_outputs(2242));
    layer2_outputs(1202) <= not((layer1_outputs(679)) or (layer1_outputs(350)));
    layer2_outputs(1203) <= layer1_outputs(36);
    layer2_outputs(1204) <= layer1_outputs(160);
    layer2_outputs(1205) <= not(layer1_outputs(2234));
    layer2_outputs(1206) <= not(layer1_outputs(983));
    layer2_outputs(1207) <= layer1_outputs(1045);
    layer2_outputs(1208) <= (layer1_outputs(1981)) xor (layer1_outputs(303));
    layer2_outputs(1209) <= not(layer1_outputs(930));
    layer2_outputs(1210) <= (layer1_outputs(1187)) and (layer1_outputs(937));
    layer2_outputs(1211) <= (layer1_outputs(1460)) or (layer1_outputs(2440));
    layer2_outputs(1212) <= (layer1_outputs(300)) and not (layer1_outputs(1236));
    layer2_outputs(1213) <= (layer1_outputs(1327)) and not (layer1_outputs(132));
    layer2_outputs(1214) <= (layer1_outputs(31)) and (layer1_outputs(1428));
    layer2_outputs(1215) <= (layer1_outputs(1830)) or (layer1_outputs(517));
    layer2_outputs(1216) <= layer1_outputs(1765);
    layer2_outputs(1217) <= not(layer1_outputs(1224));
    layer2_outputs(1218) <= not((layer1_outputs(2178)) or (layer1_outputs(2289)));
    layer2_outputs(1219) <= not((layer1_outputs(1092)) and (layer1_outputs(598)));
    layer2_outputs(1220) <= not((layer1_outputs(559)) xor (layer1_outputs(1035)));
    layer2_outputs(1221) <= (layer1_outputs(316)) and (layer1_outputs(1725));
    layer2_outputs(1222) <= not(layer1_outputs(346)) or (layer1_outputs(1275));
    layer2_outputs(1223) <= not(layer1_outputs(1001)) or (layer1_outputs(2153));
    layer2_outputs(1224) <= layer1_outputs(1440);
    layer2_outputs(1225) <= not((layer1_outputs(2004)) and (layer1_outputs(755)));
    layer2_outputs(1226) <= not(layer1_outputs(2415)) or (layer1_outputs(2360));
    layer2_outputs(1227) <= layer1_outputs(1641);
    layer2_outputs(1228) <= not(layer1_outputs(833));
    layer2_outputs(1229) <= layer1_outputs(785);
    layer2_outputs(1230) <= not(layer1_outputs(1093));
    layer2_outputs(1231) <= not(layer1_outputs(778));
    layer2_outputs(1232) <= not(layer1_outputs(2413));
    layer2_outputs(1233) <= layer1_outputs(682);
    layer2_outputs(1234) <= not(layer1_outputs(773));
    layer2_outputs(1235) <= layer1_outputs(2465);
    layer2_outputs(1236) <= not(layer1_outputs(1664)) or (layer1_outputs(349));
    layer2_outputs(1237) <= layer1_outputs(212);
    layer2_outputs(1238) <= (layer1_outputs(2261)) or (layer1_outputs(2031));
    layer2_outputs(1239) <= layer1_outputs(605);
    layer2_outputs(1240) <= '1';
    layer2_outputs(1241) <= not(layer1_outputs(66));
    layer2_outputs(1242) <= (layer1_outputs(815)) and not (layer1_outputs(1814));
    layer2_outputs(1243) <= not(layer1_outputs(1960)) or (layer1_outputs(1408));
    layer2_outputs(1244) <= not(layer1_outputs(688));
    layer2_outputs(1245) <= not(layer1_outputs(29));
    layer2_outputs(1246) <= not(layer1_outputs(585));
    layer2_outputs(1247) <= not((layer1_outputs(1949)) and (layer1_outputs(2516)));
    layer2_outputs(1248) <= not((layer1_outputs(1082)) xor (layer1_outputs(190)));
    layer2_outputs(1249) <= layer1_outputs(2259);
    layer2_outputs(1250) <= (layer1_outputs(1316)) or (layer1_outputs(434));
    layer2_outputs(1251) <= layer1_outputs(1206);
    layer2_outputs(1252) <= layer1_outputs(1242);
    layer2_outputs(1253) <= not((layer1_outputs(1171)) or (layer1_outputs(2367)));
    layer2_outputs(1254) <= layer1_outputs(448);
    layer2_outputs(1255) <= layer1_outputs(1854);
    layer2_outputs(1256) <= (layer1_outputs(1878)) xor (layer1_outputs(1424));
    layer2_outputs(1257) <= not(layer1_outputs(268)) or (layer1_outputs(1160));
    layer2_outputs(1258) <= layer1_outputs(1377);
    layer2_outputs(1259) <= not(layer1_outputs(1268));
    layer2_outputs(1260) <= not(layer1_outputs(959)) or (layer1_outputs(1928));
    layer2_outputs(1261) <= not(layer1_outputs(911));
    layer2_outputs(1262) <= not(layer1_outputs(1201));
    layer2_outputs(1263) <= not(layer1_outputs(1922));
    layer2_outputs(1264) <= layer1_outputs(1348);
    layer2_outputs(1265) <= layer1_outputs(155);
    layer2_outputs(1266) <= layer1_outputs(2067);
    layer2_outputs(1267) <= not((layer1_outputs(1124)) or (layer1_outputs(1157)));
    layer2_outputs(1268) <= layer1_outputs(751);
    layer2_outputs(1269) <= not((layer1_outputs(1233)) or (layer1_outputs(13)));
    layer2_outputs(1270) <= (layer1_outputs(1192)) or (layer1_outputs(365));
    layer2_outputs(1271) <= layer1_outputs(526);
    layer2_outputs(1272) <= layer1_outputs(1038);
    layer2_outputs(1273) <= layer1_outputs(973);
    layer2_outputs(1274) <= '1';
    layer2_outputs(1275) <= '0';
    layer2_outputs(1276) <= not(layer1_outputs(1392)) or (layer1_outputs(1244));
    layer2_outputs(1277) <= (layer1_outputs(992)) and not (layer1_outputs(1141));
    layer2_outputs(1278) <= '1';
    layer2_outputs(1279) <= layer1_outputs(1328);
    layer2_outputs(1280) <= not(layer1_outputs(379));
    layer2_outputs(1281) <= layer1_outputs(760);
    layer2_outputs(1282) <= not(layer1_outputs(1298)) or (layer1_outputs(2461));
    layer2_outputs(1283) <= (layer1_outputs(398)) and not (layer1_outputs(2473));
    layer2_outputs(1284) <= not(layer1_outputs(1502));
    layer2_outputs(1285) <= (layer1_outputs(2519)) and (layer1_outputs(1892));
    layer2_outputs(1286) <= layer1_outputs(1950);
    layer2_outputs(1287) <= not((layer1_outputs(206)) and (layer1_outputs(1869)));
    layer2_outputs(1288) <= layer1_outputs(1533);
    layer2_outputs(1289) <= (layer1_outputs(1419)) and not (layer1_outputs(2540));
    layer2_outputs(1290) <= layer1_outputs(683);
    layer2_outputs(1291) <= (layer1_outputs(2545)) and not (layer1_outputs(2204));
    layer2_outputs(1292) <= layer1_outputs(102);
    layer2_outputs(1293) <= not(layer1_outputs(603));
    layer2_outputs(1294) <= (layer1_outputs(938)) or (layer1_outputs(1436));
    layer2_outputs(1295) <= not(layer1_outputs(211));
    layer2_outputs(1296) <= not(layer1_outputs(2557));
    layer2_outputs(1297) <= not(layer1_outputs(969));
    layer2_outputs(1298) <= not(layer1_outputs(1295));
    layer2_outputs(1299) <= not((layer1_outputs(415)) xor (layer1_outputs(1982)));
    layer2_outputs(1300) <= layer1_outputs(1367);
    layer2_outputs(1301) <= layer1_outputs(824);
    layer2_outputs(1302) <= not((layer1_outputs(1838)) xor (layer1_outputs(1635)));
    layer2_outputs(1303) <= (layer1_outputs(1063)) or (layer1_outputs(1982));
    layer2_outputs(1304) <= (layer1_outputs(405)) and not (layer1_outputs(1405));
    layer2_outputs(1305) <= not(layer1_outputs(1));
    layer2_outputs(1306) <= not(layer1_outputs(48));
    layer2_outputs(1307) <= layer1_outputs(275);
    layer2_outputs(1308) <= (layer1_outputs(1174)) xor (layer1_outputs(1087));
    layer2_outputs(1309) <= not(layer1_outputs(1128));
    layer2_outputs(1310) <= (layer1_outputs(22)) and (layer1_outputs(1586));
    layer2_outputs(1311) <= not(layer1_outputs(1822));
    layer2_outputs(1312) <= not((layer1_outputs(1925)) and (layer1_outputs(242)));
    layer2_outputs(1313) <= not(layer1_outputs(2411));
    layer2_outputs(1314) <= not(layer1_outputs(1420));
    layer2_outputs(1315) <= not(layer1_outputs(2485));
    layer2_outputs(1316) <= not(layer1_outputs(964));
    layer2_outputs(1317) <= not(layer1_outputs(52));
    layer2_outputs(1318) <= not(layer1_outputs(2101));
    layer2_outputs(1319) <= layer1_outputs(86);
    layer2_outputs(1320) <= (layer1_outputs(494)) or (layer1_outputs(332));
    layer2_outputs(1321) <= not(layer1_outputs(1799));
    layer2_outputs(1322) <= not(layer1_outputs(2424));
    layer2_outputs(1323) <= not((layer1_outputs(2150)) or (layer1_outputs(410)));
    layer2_outputs(1324) <= not(layer1_outputs(750));
    layer2_outputs(1325) <= not(layer1_outputs(640)) or (layer1_outputs(886));
    layer2_outputs(1326) <= (layer1_outputs(584)) xor (layer1_outputs(952));
    layer2_outputs(1327) <= layer1_outputs(297);
    layer2_outputs(1328) <= not(layer1_outputs(2390)) or (layer1_outputs(311));
    layer2_outputs(1329) <= not(layer1_outputs(623));
    layer2_outputs(1330) <= not((layer1_outputs(626)) or (layer1_outputs(12)));
    layer2_outputs(1331) <= layer1_outputs(674);
    layer2_outputs(1332) <= not(layer1_outputs(2396));
    layer2_outputs(1333) <= (layer1_outputs(245)) or (layer1_outputs(1975));
    layer2_outputs(1334) <= not((layer1_outputs(2065)) or (layer1_outputs(1899)));
    layer2_outputs(1335) <= (layer1_outputs(1225)) and not (layer1_outputs(1723));
    layer2_outputs(1336) <= not((layer1_outputs(1190)) and (layer1_outputs(653)));
    layer2_outputs(1337) <= not(layer1_outputs(2506));
    layer2_outputs(1338) <= layer1_outputs(25);
    layer2_outputs(1339) <= (layer1_outputs(1557)) and not (layer1_outputs(2127));
    layer2_outputs(1340) <= '0';
    layer2_outputs(1341) <= not((layer1_outputs(1168)) or (layer1_outputs(1822)));
    layer2_outputs(1342) <= not(layer1_outputs(1556));
    layer2_outputs(1343) <= not(layer1_outputs(2192));
    layer2_outputs(1344) <= layer1_outputs(1775);
    layer2_outputs(1345) <= layer1_outputs(1472);
    layer2_outputs(1346) <= (layer1_outputs(1091)) and (layer1_outputs(1384));
    layer2_outputs(1347) <= (layer1_outputs(633)) and not (layer1_outputs(2498));
    layer2_outputs(1348) <= (layer1_outputs(2476)) and (layer1_outputs(736));
    layer2_outputs(1349) <= not(layer1_outputs(2497));
    layer2_outputs(1350) <= not(layer1_outputs(1929));
    layer2_outputs(1351) <= (layer1_outputs(678)) and not (layer1_outputs(169));
    layer2_outputs(1352) <= not(layer1_outputs(1736));
    layer2_outputs(1353) <= (layer1_outputs(1204)) and not (layer1_outputs(546));
    layer2_outputs(1354) <= (layer1_outputs(1491)) or (layer1_outputs(882));
    layer2_outputs(1355) <= not(layer1_outputs(1542));
    layer2_outputs(1356) <= (layer1_outputs(1539)) and not (layer1_outputs(2289));
    layer2_outputs(1357) <= (layer1_outputs(797)) and not (layer1_outputs(1958));
    layer2_outputs(1358) <= not((layer1_outputs(2259)) and (layer1_outputs(2197)));
    layer2_outputs(1359) <= not((layer1_outputs(1024)) and (layer1_outputs(1659)));
    layer2_outputs(1360) <= not(layer1_outputs(1688));
    layer2_outputs(1361) <= '1';
    layer2_outputs(1362) <= not((layer1_outputs(545)) or (layer1_outputs(143)));
    layer2_outputs(1363) <= layer1_outputs(257);
    layer2_outputs(1364) <= not(layer1_outputs(1870));
    layer2_outputs(1365) <= not((layer1_outputs(1763)) and (layer1_outputs(550)));
    layer2_outputs(1366) <= layer1_outputs(634);
    layer2_outputs(1367) <= not(layer1_outputs(873));
    layer2_outputs(1368) <= not((layer1_outputs(553)) xor (layer1_outputs(1299)));
    layer2_outputs(1369) <= not(layer1_outputs(166));
    layer2_outputs(1370) <= (layer1_outputs(1178)) and not (layer1_outputs(578));
    layer2_outputs(1371) <= (layer1_outputs(1874)) and (layer1_outputs(946));
    layer2_outputs(1372) <= layer1_outputs(2119);
    layer2_outputs(1373) <= (layer1_outputs(982)) and (layer1_outputs(1837));
    layer2_outputs(1374) <= layer1_outputs(205);
    layer2_outputs(1375) <= not((layer1_outputs(1674)) and (layer1_outputs(806)));
    layer2_outputs(1376) <= (layer1_outputs(2364)) and not (layer1_outputs(1087));
    layer2_outputs(1377) <= '1';
    layer2_outputs(1378) <= not(layer1_outputs(1849)) or (layer1_outputs(2379));
    layer2_outputs(1379) <= not(layer1_outputs(772));
    layer2_outputs(1380) <= not((layer1_outputs(1532)) or (layer1_outputs(838)));
    layer2_outputs(1381) <= not(layer1_outputs(631)) or (layer1_outputs(1668));
    layer2_outputs(1382) <= not(layer1_outputs(2429));
    layer2_outputs(1383) <= not(layer1_outputs(117)) or (layer1_outputs(2450));
    layer2_outputs(1384) <= (layer1_outputs(1389)) or (layer1_outputs(628));
    layer2_outputs(1385) <= (layer1_outputs(1282)) and (layer1_outputs(1429));
    layer2_outputs(1386) <= not(layer1_outputs(1813));
    layer2_outputs(1387) <= not(layer1_outputs(472));
    layer2_outputs(1388) <= (layer1_outputs(1304)) and (layer1_outputs(904));
    layer2_outputs(1389) <= not(layer1_outputs(171));
    layer2_outputs(1390) <= layer1_outputs(963);
    layer2_outputs(1391) <= '0';
    layer2_outputs(1392) <= not(layer1_outputs(1002));
    layer2_outputs(1393) <= layer1_outputs(1749);
    layer2_outputs(1394) <= layer1_outputs(626);
    layer2_outputs(1395) <= layer1_outputs(1146);
    layer2_outputs(1396) <= not(layer1_outputs(2265));
    layer2_outputs(1397) <= not(layer1_outputs(2058));
    layer2_outputs(1398) <= layer1_outputs(2133);
    layer2_outputs(1399) <= not(layer1_outputs(2229)) or (layer1_outputs(1881));
    layer2_outputs(1400) <= layer1_outputs(658);
    layer2_outputs(1401) <= layer1_outputs(2359);
    layer2_outputs(1402) <= (layer1_outputs(1219)) and (layer1_outputs(957));
    layer2_outputs(1403) <= not((layer1_outputs(271)) xor (layer1_outputs(400)));
    layer2_outputs(1404) <= not(layer1_outputs(2493)) or (layer1_outputs(1452));
    layer2_outputs(1405) <= not(layer1_outputs(1362));
    layer2_outputs(1406) <= (layer1_outputs(849)) and not (layer1_outputs(58));
    layer2_outputs(1407) <= (layer1_outputs(2393)) and not (layer1_outputs(2373));
    layer2_outputs(1408) <= layer1_outputs(84);
    layer2_outputs(1409) <= layer1_outputs(228);
    layer2_outputs(1410) <= not(layer1_outputs(1253));
    layer2_outputs(1411) <= (layer1_outputs(2113)) and not (layer1_outputs(1488));
    layer2_outputs(1412) <= (layer1_outputs(584)) and not (layer1_outputs(2322));
    layer2_outputs(1413) <= not(layer1_outputs(1461)) or (layer1_outputs(1555));
    layer2_outputs(1414) <= not(layer1_outputs(577));
    layer2_outputs(1415) <= not(layer1_outputs(715));
    layer2_outputs(1416) <= (layer1_outputs(330)) xor (layer1_outputs(178));
    layer2_outputs(1417) <= not(layer1_outputs(1125));
    layer2_outputs(1418) <= not(layer1_outputs(0)) or (layer1_outputs(1380));
    layer2_outputs(1419) <= (layer1_outputs(129)) and not (layer1_outputs(2316));
    layer2_outputs(1420) <= not((layer1_outputs(106)) or (layer1_outputs(65)));
    layer2_outputs(1421) <= not(layer1_outputs(961));
    layer2_outputs(1422) <= not(layer1_outputs(1096));
    layer2_outputs(1423) <= layer1_outputs(444);
    layer2_outputs(1424) <= not(layer1_outputs(569)) or (layer1_outputs(637));
    layer2_outputs(1425) <= (layer1_outputs(2530)) and (layer1_outputs(1636));
    layer2_outputs(1426) <= layer1_outputs(1852);
    layer2_outputs(1427) <= (layer1_outputs(1534)) and (layer1_outputs(2122));
    layer2_outputs(1428) <= not(layer1_outputs(2006)) or (layer1_outputs(1368));
    layer2_outputs(1429) <= '1';
    layer2_outputs(1430) <= not(layer1_outputs(947));
    layer2_outputs(1431) <= layer1_outputs(889);
    layer2_outputs(1432) <= not((layer1_outputs(2026)) xor (layer1_outputs(335)));
    layer2_outputs(1433) <= not(layer1_outputs(47));
    layer2_outputs(1434) <= layer1_outputs(2172);
    layer2_outputs(1435) <= not(layer1_outputs(1131));
    layer2_outputs(1436) <= layer1_outputs(1527);
    layer2_outputs(1437) <= not(layer1_outputs(2020));
    layer2_outputs(1438) <= (layer1_outputs(1513)) and not (layer1_outputs(1931));
    layer2_outputs(1439) <= not(layer1_outputs(1819));
    layer2_outputs(1440) <= (layer1_outputs(2313)) or (layer1_outputs(956));
    layer2_outputs(1441) <= (layer1_outputs(2457)) or (layer1_outputs(1535));
    layer2_outputs(1442) <= (layer1_outputs(469)) and not (layer1_outputs(1759));
    layer2_outputs(1443) <= not(layer1_outputs(590));
    layer2_outputs(1444) <= not(layer1_outputs(830));
    layer2_outputs(1445) <= (layer1_outputs(2303)) and (layer1_outputs(566));
    layer2_outputs(1446) <= '0';
    layer2_outputs(1447) <= not(layer1_outputs(2526));
    layer2_outputs(1448) <= not(layer1_outputs(620)) or (layer1_outputs(751));
    layer2_outputs(1449) <= '1';
    layer2_outputs(1450) <= not(layer1_outputs(940));
    layer2_outputs(1451) <= (layer1_outputs(596)) or (layer1_outputs(1427));
    layer2_outputs(1452) <= layer1_outputs(418);
    layer2_outputs(1453) <= not(layer1_outputs(2474));
    layer2_outputs(1454) <= not(layer1_outputs(481));
    layer2_outputs(1455) <= not(layer1_outputs(730));
    layer2_outputs(1456) <= layer1_outputs(846);
    layer2_outputs(1457) <= not(layer1_outputs(1140)) or (layer1_outputs(1998));
    layer2_outputs(1458) <= not(layer1_outputs(97));
    layer2_outputs(1459) <= (layer1_outputs(748)) and not (layer1_outputs(1718));
    layer2_outputs(1460) <= not((layer1_outputs(433)) and (layer1_outputs(1531)));
    layer2_outputs(1461) <= not(layer1_outputs(1009));
    layer2_outputs(1462) <= not(layer1_outputs(1450));
    layer2_outputs(1463) <= not(layer1_outputs(1831)) or (layer1_outputs(1904));
    layer2_outputs(1464) <= not(layer1_outputs(177));
    layer2_outputs(1465) <= (layer1_outputs(2397)) and not (layer1_outputs(539));
    layer2_outputs(1466) <= (layer1_outputs(571)) and (layer1_outputs(2428));
    layer2_outputs(1467) <= not(layer1_outputs(2233));
    layer2_outputs(1468) <= not(layer1_outputs(1575));
    layer2_outputs(1469) <= (layer1_outputs(2367)) or (layer1_outputs(2255));
    layer2_outputs(1470) <= not(layer1_outputs(384));
    layer2_outputs(1471) <= (layer1_outputs(2329)) and not (layer1_outputs(900));
    layer2_outputs(1472) <= not(layer1_outputs(980));
    layer2_outputs(1473) <= (layer1_outputs(169)) or (layer1_outputs(1967));
    layer2_outputs(1474) <= not(layer1_outputs(1173));
    layer2_outputs(1475) <= not(layer1_outputs(1509)) or (layer1_outputs(474));
    layer2_outputs(1476) <= not(layer1_outputs(1454));
    layer2_outputs(1477) <= (layer1_outputs(1679)) or (layer1_outputs(529));
    layer2_outputs(1478) <= not(layer1_outputs(850)) or (layer1_outputs(928));
    layer2_outputs(1479) <= not((layer1_outputs(135)) and (layer1_outputs(384)));
    layer2_outputs(1480) <= not(layer1_outputs(534));
    layer2_outputs(1481) <= layer1_outputs(1730);
    layer2_outputs(1482) <= not(layer1_outputs(762));
    layer2_outputs(1483) <= not((layer1_outputs(735)) or (layer1_outputs(1524)));
    layer2_outputs(1484) <= layer1_outputs(2270);
    layer2_outputs(1485) <= layer1_outputs(322);
    layer2_outputs(1486) <= not(layer1_outputs(18)) or (layer1_outputs(1634));
    layer2_outputs(1487) <= layer1_outputs(2180);
    layer2_outputs(1488) <= not(layer1_outputs(152)) or (layer1_outputs(957));
    layer2_outputs(1489) <= layer1_outputs(1350);
    layer2_outputs(1490) <= (layer1_outputs(1658)) xor (layer1_outputs(42));
    layer2_outputs(1491) <= not(layer1_outputs(1008));
    layer2_outputs(1492) <= not(layer1_outputs(83));
    layer2_outputs(1493) <= not((layer1_outputs(614)) and (layer1_outputs(739)));
    layer2_outputs(1494) <= not(layer1_outputs(2412));
    layer2_outputs(1495) <= not((layer1_outputs(2477)) and (layer1_outputs(1510)));
    layer2_outputs(1496) <= not(layer1_outputs(265));
    layer2_outputs(1497) <= (layer1_outputs(476)) and not (layer1_outputs(1402));
    layer2_outputs(1498) <= not(layer1_outputs(782));
    layer2_outputs(1499) <= not(layer1_outputs(1817));
    layer2_outputs(1500) <= (layer1_outputs(1554)) and not (layer1_outputs(1669));
    layer2_outputs(1501) <= layer1_outputs(1673);
    layer2_outputs(1502) <= (layer1_outputs(483)) or (layer1_outputs(2077));
    layer2_outputs(1503) <= not(layer1_outputs(1891));
    layer2_outputs(1504) <= layer1_outputs(321);
    layer2_outputs(1505) <= not(layer1_outputs(2346));
    layer2_outputs(1506) <= not(layer1_outputs(624)) or (layer1_outputs(161));
    layer2_outputs(1507) <= not(layer1_outputs(1872));
    layer2_outputs(1508) <= not(layer1_outputs(1993));
    layer2_outputs(1509) <= (layer1_outputs(1992)) and not (layer1_outputs(2092));
    layer2_outputs(1510) <= not(layer1_outputs(574));
    layer2_outputs(1511) <= not(layer1_outputs(29));
    layer2_outputs(1512) <= layer1_outputs(507);
    layer2_outputs(1513) <= (layer1_outputs(1697)) and not (layer1_outputs(1875));
    layer2_outputs(1514) <= layer1_outputs(2531);
    layer2_outputs(1515) <= layer1_outputs(539);
    layer2_outputs(1516) <= layer1_outputs(186);
    layer2_outputs(1517) <= (layer1_outputs(328)) and (layer1_outputs(119));
    layer2_outputs(1518) <= not(layer1_outputs(2057)) or (layer1_outputs(2162));
    layer2_outputs(1519) <= layer1_outputs(642);
    layer2_outputs(1520) <= layer1_outputs(1419);
    layer2_outputs(1521) <= not((layer1_outputs(428)) xor (layer1_outputs(689)));
    layer2_outputs(1522) <= (layer1_outputs(2241)) and not (layer1_outputs(1101));
    layer2_outputs(1523) <= layer1_outputs(726);
    layer2_outputs(1524) <= (layer1_outputs(1131)) or (layer1_outputs(971));
    layer2_outputs(1525) <= not(layer1_outputs(763));
    layer2_outputs(1526) <= layer1_outputs(427);
    layer2_outputs(1527) <= not(layer1_outputs(1496));
    layer2_outputs(1528) <= layer1_outputs(115);
    layer2_outputs(1529) <= not((layer1_outputs(63)) or (layer1_outputs(105)));
    layer2_outputs(1530) <= layer1_outputs(174);
    layer2_outputs(1531) <= layer1_outputs(1069);
    layer2_outputs(1532) <= not(layer1_outputs(2148));
    layer2_outputs(1533) <= (layer1_outputs(2274)) and (layer1_outputs(1676));
    layer2_outputs(1534) <= not(layer1_outputs(1660)) or (layer1_outputs(1705));
    layer2_outputs(1535) <= layer1_outputs(440);
    layer2_outputs(1536) <= (layer1_outputs(2522)) or (layer1_outputs(2527));
    layer2_outputs(1537) <= not(layer1_outputs(788));
    layer2_outputs(1538) <= not(layer1_outputs(649));
    layer2_outputs(1539) <= (layer1_outputs(377)) and (layer1_outputs(1789));
    layer2_outputs(1540) <= layer1_outputs(1619);
    layer2_outputs(1541) <= layer1_outputs(492);
    layer2_outputs(1542) <= not(layer1_outputs(1150));
    layer2_outputs(1543) <= (layer1_outputs(2449)) and (layer1_outputs(370));
    layer2_outputs(1544) <= layer1_outputs(1884);
    layer2_outputs(1545) <= not(layer1_outputs(1364));
    layer2_outputs(1546) <= not(layer1_outputs(117));
    layer2_outputs(1547) <= layer1_outputs(1029);
    layer2_outputs(1548) <= '0';
    layer2_outputs(1549) <= not(layer1_outputs(903));
    layer2_outputs(1550) <= not((layer1_outputs(1557)) or (layer1_outputs(599)));
    layer2_outputs(1551) <= not(layer1_outputs(2441)) or (layer1_outputs(2119));
    layer2_outputs(1552) <= not(layer1_outputs(1485));
    layer2_outputs(1553) <= not(layer1_outputs(723));
    layer2_outputs(1554) <= not(layer1_outputs(79));
    layer2_outputs(1555) <= not(layer1_outputs(46)) or (layer1_outputs(2353));
    layer2_outputs(1556) <= layer1_outputs(2318);
    layer2_outputs(1557) <= not(layer1_outputs(1494));
    layer2_outputs(1558) <= (layer1_outputs(1942)) or (layer1_outputs(25));
    layer2_outputs(1559) <= not(layer1_outputs(290));
    layer2_outputs(1560) <= (layer1_outputs(1913)) and (layer1_outputs(1555));
    layer2_outputs(1561) <= (layer1_outputs(668)) or (layer1_outputs(2377));
    layer2_outputs(1562) <= (layer1_outputs(2396)) and not (layer1_outputs(1315));
    layer2_outputs(1563) <= not(layer1_outputs(2112));
    layer2_outputs(1564) <= not(layer1_outputs(485));
    layer2_outputs(1565) <= (layer1_outputs(2381)) and not (layer1_outputs(1740));
    layer2_outputs(1566) <= not(layer1_outputs(385)) or (layer1_outputs(2443));
    layer2_outputs(1567) <= not(layer1_outputs(1195));
    layer2_outputs(1568) <= not((layer1_outputs(2040)) or (layer1_outputs(460)));
    layer2_outputs(1569) <= not(layer1_outputs(2418)) or (layer1_outputs(767));
    layer2_outputs(1570) <= (layer1_outputs(1538)) and (layer1_outputs(1112));
    layer2_outputs(1571) <= not(layer1_outputs(2158));
    layer2_outputs(1572) <= not(layer1_outputs(1325)) or (layer1_outputs(1752));
    layer2_outputs(1573) <= layer1_outputs(1694);
    layer2_outputs(1574) <= not(layer1_outputs(2103)) or (layer1_outputs(2225));
    layer2_outputs(1575) <= not((layer1_outputs(1427)) or (layer1_outputs(2090)));
    layer2_outputs(1576) <= not(layer1_outputs(986));
    layer2_outputs(1577) <= (layer1_outputs(1882)) and not (layer1_outputs(2171));
    layer2_outputs(1578) <= (layer1_outputs(411)) and (layer1_outputs(1260));
    layer2_outputs(1579) <= not(layer1_outputs(1792)) or (layer1_outputs(16));
    layer2_outputs(1580) <= layer1_outputs(2044);
    layer2_outputs(1581) <= (layer1_outputs(1114)) and not (layer1_outputs(1868));
    layer2_outputs(1582) <= layer1_outputs(424);
    layer2_outputs(1583) <= not(layer1_outputs(475));
    layer2_outputs(1584) <= not((layer1_outputs(759)) and (layer1_outputs(2254)));
    layer2_outputs(1585) <= (layer1_outputs(1025)) and not (layer1_outputs(2073));
    layer2_outputs(1586) <= layer1_outputs(1564);
    layer2_outputs(1587) <= not(layer1_outputs(2366)) or (layer1_outputs(445));
    layer2_outputs(1588) <= layer1_outputs(1749);
    layer2_outputs(1589) <= not(layer1_outputs(635)) or (layer1_outputs(1548));
    layer2_outputs(1590) <= (layer1_outputs(2266)) and (layer1_outputs(873));
    layer2_outputs(1591) <= not(layer1_outputs(394)) or (layer1_outputs(2042));
    layer2_outputs(1592) <= layer1_outputs(1436);
    layer2_outputs(1593) <= (layer1_outputs(461)) and not (layer1_outputs(1846));
    layer2_outputs(1594) <= not(layer1_outputs(47));
    layer2_outputs(1595) <= (layer1_outputs(1561)) and (layer1_outputs(1579));
    layer2_outputs(1596) <= (layer1_outputs(2299)) xor (layer1_outputs(57));
    layer2_outputs(1597) <= (layer1_outputs(53)) or (layer1_outputs(1310));
    layer2_outputs(1598) <= not((layer1_outputs(26)) and (layer1_outputs(1562)));
    layer2_outputs(1599) <= layer1_outputs(1590);
    layer2_outputs(1600) <= not(layer1_outputs(2336));
    layer2_outputs(1601) <= not(layer1_outputs(1226));
    layer2_outputs(1602) <= not(layer1_outputs(1587));
    layer2_outputs(1603) <= layer1_outputs(1693);
    layer2_outputs(1604) <= (layer1_outputs(1154)) and not (layer1_outputs(2343));
    layer2_outputs(1605) <= not(layer1_outputs(2463)) or (layer1_outputs(1152));
    layer2_outputs(1606) <= not(layer1_outputs(1416)) or (layer1_outputs(2535));
    layer2_outputs(1607) <= not(layer1_outputs(816));
    layer2_outputs(1608) <= not((layer1_outputs(2072)) or (layer1_outputs(808)));
    layer2_outputs(1609) <= not(layer1_outputs(199)) or (layer1_outputs(23));
    layer2_outputs(1610) <= (layer1_outputs(100)) and not (layer1_outputs(2543));
    layer2_outputs(1611) <= not(layer1_outputs(548));
    layer2_outputs(1612) <= layer1_outputs(330);
    layer2_outputs(1613) <= (layer1_outputs(2511)) and not (layer1_outputs(2316));
    layer2_outputs(1614) <= not(layer1_outputs(1898));
    layer2_outputs(1615) <= (layer1_outputs(700)) and not (layer1_outputs(2550));
    layer2_outputs(1616) <= (layer1_outputs(2226)) or (layer1_outputs(487));
    layer2_outputs(1617) <= '0';
    layer2_outputs(1618) <= layer1_outputs(2459);
    layer2_outputs(1619) <= (layer1_outputs(1261)) and not (layer1_outputs(1365));
    layer2_outputs(1620) <= not(layer1_outputs(1780));
    layer2_outputs(1621) <= (layer1_outputs(16)) and not (layer1_outputs(1842));
    layer2_outputs(1622) <= (layer1_outputs(1339)) xor (layer1_outputs(142));
    layer2_outputs(1623) <= '0';
    layer2_outputs(1624) <= layer1_outputs(1206);
    layer2_outputs(1625) <= layer1_outputs(889);
    layer2_outputs(1626) <= layer1_outputs(1383);
    layer2_outputs(1627) <= not((layer1_outputs(552)) or (layer1_outputs(2131)));
    layer2_outputs(1628) <= '1';
    layer2_outputs(1629) <= not(layer1_outputs(1335));
    layer2_outputs(1630) <= layer1_outputs(232);
    layer2_outputs(1631) <= (layer1_outputs(1633)) and not (layer1_outputs(1252));
    layer2_outputs(1632) <= not(layer1_outputs(215));
    layer2_outputs(1633) <= not(layer1_outputs(512));
    layer2_outputs(1634) <= (layer1_outputs(951)) and not (layer1_outputs(2199));
    layer2_outputs(1635) <= layer1_outputs(93);
    layer2_outputs(1636) <= layer1_outputs(1787);
    layer2_outputs(1637) <= not(layer1_outputs(473));
    layer2_outputs(1638) <= not(layer1_outputs(2114)) or (layer1_outputs(27));
    layer2_outputs(1639) <= not(layer1_outputs(1775));
    layer2_outputs(1640) <= layer1_outputs(2131);
    layer2_outputs(1641) <= not(layer1_outputs(1931)) or (layer1_outputs(583));
    layer2_outputs(1642) <= (layer1_outputs(2410)) and (layer1_outputs(1526));
    layer2_outputs(1643) <= (layer1_outputs(1642)) or (layer1_outputs(1194));
    layer2_outputs(1644) <= (layer1_outputs(1355)) and (layer1_outputs(143));
    layer2_outputs(1645) <= layer1_outputs(2156);
    layer2_outputs(1646) <= not(layer1_outputs(1080)) or (layer1_outputs(1363));
    layer2_outputs(1647) <= not((layer1_outputs(2034)) and (layer1_outputs(2481)));
    layer2_outputs(1648) <= (layer1_outputs(641)) and not (layer1_outputs(1457));
    layer2_outputs(1649) <= not(layer1_outputs(2284));
    layer2_outputs(1650) <= not(layer1_outputs(1257)) or (layer1_outputs(1919));
    layer2_outputs(1651) <= (layer1_outputs(1712)) and not (layer1_outputs(691));
    layer2_outputs(1652) <= layer1_outputs(1519);
    layer2_outputs(1653) <= (layer1_outputs(1133)) and not (layer1_outputs(1464));
    layer2_outputs(1654) <= not((layer1_outputs(1103)) or (layer1_outputs(2038)));
    layer2_outputs(1655) <= not(layer1_outputs(2037)) or (layer1_outputs(1723));
    layer2_outputs(1656) <= not(layer1_outputs(282));
    layer2_outputs(1657) <= not(layer1_outputs(1476));
    layer2_outputs(1658) <= (layer1_outputs(2281)) and not (layer1_outputs(96));
    layer2_outputs(1659) <= not(layer1_outputs(725));
    layer2_outputs(1660) <= layer1_outputs(1962);
    layer2_outputs(1661) <= not(layer1_outputs(1916));
    layer2_outputs(1662) <= not(layer1_outputs(2403)) or (layer1_outputs(749));
    layer2_outputs(1663) <= not(layer1_outputs(1261));
    layer2_outputs(1664) <= (layer1_outputs(76)) and not (layer1_outputs(69));
    layer2_outputs(1665) <= layer1_outputs(1837);
    layer2_outputs(1666) <= (layer1_outputs(764)) and not (layer1_outputs(2498));
    layer2_outputs(1667) <= (layer1_outputs(1298)) and (layer1_outputs(2524));
    layer2_outputs(1668) <= not(layer1_outputs(1784)) or (layer1_outputs(213));
    layer2_outputs(1669) <= not((layer1_outputs(1432)) xor (layer1_outputs(2188)));
    layer2_outputs(1670) <= not((layer1_outputs(761)) or (layer1_outputs(229)));
    layer2_outputs(1671) <= not((layer1_outputs(2423)) or (layer1_outputs(581)));
    layer2_outputs(1672) <= layer1_outputs(166);
    layer2_outputs(1673) <= not(layer1_outputs(580));
    layer2_outputs(1674) <= (layer1_outputs(263)) and (layer1_outputs(93));
    layer2_outputs(1675) <= not(layer1_outputs(954)) or (layer1_outputs(1894));
    layer2_outputs(1676) <= not(layer1_outputs(2214));
    layer2_outputs(1677) <= not(layer1_outputs(2053)) or (layer1_outputs(2262));
    layer2_outputs(1678) <= layer1_outputs(1023);
    layer2_outputs(1679) <= not(layer1_outputs(2147));
    layer2_outputs(1680) <= layer1_outputs(1463);
    layer2_outputs(1681) <= not((layer1_outputs(2400)) and (layer1_outputs(1929)));
    layer2_outputs(1682) <= not(layer1_outputs(2183));
    layer2_outputs(1683) <= not(layer1_outputs(433)) or (layer1_outputs(1184));
    layer2_outputs(1684) <= not((layer1_outputs(2324)) and (layer1_outputs(934)));
    layer2_outputs(1685) <= not(layer1_outputs(937)) or (layer1_outputs(2216));
    layer2_outputs(1686) <= not(layer1_outputs(764)) or (layer1_outputs(508));
    layer2_outputs(1687) <= not(layer1_outputs(2185));
    layer2_outputs(1688) <= layer1_outputs(84);
    layer2_outputs(1689) <= (layer1_outputs(2151)) or (layer1_outputs(841));
    layer2_outputs(1690) <= layer1_outputs(480);
    layer2_outputs(1691) <= not(layer1_outputs(655));
    layer2_outputs(1692) <= not((layer1_outputs(70)) or (layer1_outputs(2117)));
    layer2_outputs(1693) <= layer1_outputs(60);
    layer2_outputs(1694) <= '1';
    layer2_outputs(1695) <= not(layer1_outputs(1222));
    layer2_outputs(1696) <= not((layer1_outputs(2287)) and (layer1_outputs(9)));
    layer2_outputs(1697) <= (layer1_outputs(207)) and (layer1_outputs(2051));
    layer2_outputs(1698) <= layer1_outputs(814);
    layer2_outputs(1699) <= not((layer1_outputs(2294)) xor (layer1_outputs(1473)));
    layer2_outputs(1700) <= not(layer1_outputs(693));
    layer2_outputs(1701) <= (layer1_outputs(235)) and (layer1_outputs(2230));
    layer2_outputs(1702) <= not(layer1_outputs(1099));
    layer2_outputs(1703) <= (layer1_outputs(1081)) and (layer1_outputs(288));
    layer2_outputs(1704) <= not(layer1_outputs(36));
    layer2_outputs(1705) <= not(layer1_outputs(220));
    layer2_outputs(1706) <= not(layer1_outputs(1825));
    layer2_outputs(1707) <= layer1_outputs(391);
    layer2_outputs(1708) <= not((layer1_outputs(279)) and (layer1_outputs(1005)));
    layer2_outputs(1709) <= '1';
    layer2_outputs(1710) <= not(layer1_outputs(2406)) or (layer1_outputs(1889));
    layer2_outputs(1711) <= layer1_outputs(481);
    layer2_outputs(1712) <= not(layer1_outputs(802));
    layer2_outputs(1713) <= (layer1_outputs(88)) or (layer1_outputs(713));
    layer2_outputs(1714) <= not(layer1_outputs(1061)) or (layer1_outputs(1406));
    layer2_outputs(1715) <= (layer1_outputs(2111)) and not (layer1_outputs(815));
    layer2_outputs(1716) <= not(layer1_outputs(346));
    layer2_outputs(1717) <= not(layer1_outputs(1255));
    layer2_outputs(1718) <= not(layer1_outputs(1652));
    layer2_outputs(1719) <= not(layer1_outputs(1432));
    layer2_outputs(1720) <= not(layer1_outputs(2527));
    layer2_outputs(1721) <= not(layer1_outputs(1641)) or (layer1_outputs(78));
    layer2_outputs(1722) <= '0';
    layer2_outputs(1723) <= not(layer1_outputs(1796));
    layer2_outputs(1724) <= layer1_outputs(2347);
    layer2_outputs(1725) <= not((layer1_outputs(2412)) or (layer1_outputs(1272)));
    layer2_outputs(1726) <= not(layer1_outputs(1553));
    layer2_outputs(1727) <= (layer1_outputs(150)) or (layer1_outputs(614));
    layer2_outputs(1728) <= not((layer1_outputs(607)) or (layer1_outputs(2066)));
    layer2_outputs(1729) <= not((layer1_outputs(1565)) xor (layer1_outputs(1531)));
    layer2_outputs(1730) <= layer1_outputs(702);
    layer2_outputs(1731) <= '0';
    layer2_outputs(1732) <= layer1_outputs(1003);
    layer2_outputs(1733) <= not(layer1_outputs(721));
    layer2_outputs(1734) <= (layer1_outputs(574)) xor (layer1_outputs(2271));
    layer2_outputs(1735) <= layer1_outputs(494);
    layer2_outputs(1736) <= not(layer1_outputs(1720));
    layer2_outputs(1737) <= layer1_outputs(380);
    layer2_outputs(1738) <= (layer1_outputs(1115)) or (layer1_outputs(1356));
    layer2_outputs(1739) <= layer1_outputs(636);
    layer2_outputs(1740) <= not((layer1_outputs(1907)) and (layer1_outputs(2286)));
    layer2_outputs(1741) <= layer1_outputs(2064);
    layer2_outputs(1742) <= not((layer1_outputs(473)) or (layer1_outputs(2329)));
    layer2_outputs(1743) <= (layer1_outputs(1512)) xor (layer1_outputs(379));
    layer2_outputs(1744) <= (layer1_outputs(129)) and not (layer1_outputs(826));
    layer2_outputs(1745) <= (layer1_outputs(2492)) and not (layer1_outputs(401));
    layer2_outputs(1746) <= not(layer1_outputs(1044));
    layer2_outputs(1747) <= (layer1_outputs(2552)) xor (layer1_outputs(2434));
    layer2_outputs(1748) <= not((layer1_outputs(1352)) xor (layer1_outputs(2408)));
    layer2_outputs(1749) <= (layer1_outputs(2467)) and (layer1_outputs(1067));
    layer2_outputs(1750) <= '1';
    layer2_outputs(1751) <= not((layer1_outputs(1994)) and (layer1_outputs(1329)));
    layer2_outputs(1752) <= (layer1_outputs(2523)) xor (layer1_outputs(1425));
    layer2_outputs(1753) <= (layer1_outputs(1926)) and not (layer1_outputs(1101));
    layer2_outputs(1754) <= not(layer1_outputs(2222));
    layer2_outputs(1755) <= not(layer1_outputs(1834));
    layer2_outputs(1756) <= layer1_outputs(1399);
    layer2_outputs(1757) <= layer1_outputs(1704);
    layer2_outputs(1758) <= layer1_outputs(162);
    layer2_outputs(1759) <= layer1_outputs(698);
    layer2_outputs(1760) <= layer1_outputs(351);
    layer2_outputs(1761) <= (layer1_outputs(2236)) and not (layer1_outputs(744));
    layer2_outputs(1762) <= not((layer1_outputs(1301)) and (layer1_outputs(875)));
    layer2_outputs(1763) <= layer1_outputs(2459);
    layer2_outputs(1764) <= (layer1_outputs(1466)) and not (layer1_outputs(1286));
    layer2_outputs(1765) <= layer1_outputs(90);
    layer2_outputs(1766) <= not(layer1_outputs(824));
    layer2_outputs(1767) <= not(layer1_outputs(74));
    layer2_outputs(1768) <= layer1_outputs(1068);
    layer2_outputs(1769) <= not(layer1_outputs(554)) or (layer1_outputs(2043));
    layer2_outputs(1770) <= not(layer1_outputs(1856));
    layer2_outputs(1771) <= layer1_outputs(616);
    layer2_outputs(1772) <= layer1_outputs(1748);
    layer2_outputs(1773) <= not((layer1_outputs(962)) xor (layer1_outputs(1425)));
    layer2_outputs(1774) <= layer1_outputs(443);
    layer2_outputs(1775) <= not((layer1_outputs(1471)) xor (layer1_outputs(1280)));
    layer2_outputs(1776) <= (layer1_outputs(898)) and (layer1_outputs(814));
    layer2_outputs(1777) <= layer1_outputs(671);
    layer2_outputs(1778) <= layer1_outputs(684);
    layer2_outputs(1779) <= not((layer1_outputs(1367)) or (layer1_outputs(537)));
    layer2_outputs(1780) <= (layer1_outputs(808)) and not (layer1_outputs(495));
    layer2_outputs(1781) <= (layer1_outputs(1037)) xor (layer1_outputs(1103));
    layer2_outputs(1782) <= not(layer1_outputs(311));
    layer2_outputs(1783) <= not(layer1_outputs(945));
    layer2_outputs(1784) <= not(layer1_outputs(992));
    layer2_outputs(1785) <= layer1_outputs(994);
    layer2_outputs(1786) <= (layer1_outputs(134)) and not (layer1_outputs(1954));
    layer2_outputs(1787) <= (layer1_outputs(1259)) and not (layer1_outputs(55));
    layer2_outputs(1788) <= layer1_outputs(865);
    layer2_outputs(1789) <= not(layer1_outputs(511)) or (layer1_outputs(2146));
    layer2_outputs(1790) <= layer1_outputs(2249);
    layer2_outputs(1791) <= layer1_outputs(2223);
    layer2_outputs(1792) <= not(layer1_outputs(14));
    layer2_outputs(1793) <= not(layer1_outputs(2328)) or (layer1_outputs(2077));
    layer2_outputs(1794) <= not(layer1_outputs(868));
    layer2_outputs(1795) <= (layer1_outputs(2325)) xor (layer1_outputs(313));
    layer2_outputs(1796) <= not(layer1_outputs(2025));
    layer2_outputs(1797) <= layer1_outputs(2009);
    layer2_outputs(1798) <= not(layer1_outputs(1338)) or (layer1_outputs(215));
    layer2_outputs(1799) <= not(layer1_outputs(1098));
    layer2_outputs(1800) <= not(layer1_outputs(968)) or (layer1_outputs(569));
    layer2_outputs(1801) <= layer1_outputs(1893);
    layer2_outputs(1802) <= not(layer1_outputs(582)) or (layer1_outputs(1766));
    layer2_outputs(1803) <= not(layer1_outputs(2056));
    layer2_outputs(1804) <= layer1_outputs(56);
    layer2_outputs(1805) <= layer1_outputs(434);
    layer2_outputs(1806) <= (layer1_outputs(1064)) and not (layer1_outputs(341));
    layer2_outputs(1807) <= (layer1_outputs(732)) and (layer1_outputs(566));
    layer2_outputs(1808) <= layer1_outputs(1328);
    layer2_outputs(1809) <= not(layer1_outputs(192));
    layer2_outputs(1810) <= not(layer1_outputs(1832)) or (layer1_outputs(1528));
    layer2_outputs(1811) <= (layer1_outputs(40)) and (layer1_outputs(842));
    layer2_outputs(1812) <= not((layer1_outputs(436)) and (layer1_outputs(723)));
    layer2_outputs(1813) <= not(layer1_outputs(1051)) or (layer1_outputs(180));
    layer2_outputs(1814) <= (layer1_outputs(453)) and not (layer1_outputs(1119));
    layer2_outputs(1815) <= not(layer1_outputs(2342));
    layer2_outputs(1816) <= (layer1_outputs(2311)) and not (layer1_outputs(269));
    layer2_outputs(1817) <= layer1_outputs(861);
    layer2_outputs(1818) <= (layer1_outputs(1596)) or (layer1_outputs(1971));
    layer2_outputs(1819) <= not(layer1_outputs(2242)) or (layer1_outputs(1624));
    layer2_outputs(1820) <= not(layer1_outputs(677));
    layer2_outputs(1821) <= '0';
    layer2_outputs(1822) <= not(layer1_outputs(1449));
    layer2_outputs(1823) <= (layer1_outputs(807)) and not (layer1_outputs(2522));
    layer2_outputs(1824) <= layer1_outputs(2315);
    layer2_outputs(1825) <= not(layer1_outputs(666)) or (layer1_outputs(1378));
    layer2_outputs(1826) <= not((layer1_outputs(497)) xor (layer1_outputs(1845)));
    layer2_outputs(1827) <= not((layer1_outputs(1242)) or (layer1_outputs(34)));
    layer2_outputs(1828) <= layer1_outputs(1510);
    layer2_outputs(1829) <= layer1_outputs(2202);
    layer2_outputs(1830) <= (layer1_outputs(1722)) and not (layer1_outputs(837));
    layer2_outputs(1831) <= (layer1_outputs(1675)) and not (layer1_outputs(954));
    layer2_outputs(1832) <= not(layer1_outputs(2045)) or (layer1_outputs(1462));
    layer2_outputs(1833) <= not((layer1_outputs(1741)) and (layer1_outputs(472)));
    layer2_outputs(1834) <= layer1_outputs(1020);
    layer2_outputs(1835) <= not(layer1_outputs(405));
    layer2_outputs(1836) <= not(layer1_outputs(2163)) or (layer1_outputs(2159));
    layer2_outputs(1837) <= (layer1_outputs(1945)) and (layer1_outputs(686));
    layer2_outputs(1838) <= layer1_outputs(480);
    layer2_outputs(1839) <= not(layer1_outputs(2121));
    layer2_outputs(1840) <= not(layer1_outputs(1661)) or (layer1_outputs(989));
    layer2_outputs(1841) <= not((layer1_outputs(2094)) or (layer1_outputs(1090)));
    layer2_outputs(1842) <= (layer1_outputs(711)) and not (layer1_outputs(1627));
    layer2_outputs(1843) <= layer1_outputs(1844);
    layer2_outputs(1844) <= layer1_outputs(1441);
    layer2_outputs(1845) <= layer1_outputs(1370);
    layer2_outputs(1846) <= not(layer1_outputs(390));
    layer2_outputs(1847) <= not(layer1_outputs(2079)) or (layer1_outputs(2296));
    layer2_outputs(1848) <= layer1_outputs(338);
    layer2_outputs(1849) <= layer1_outputs(1687);
    layer2_outputs(1850) <= '0';
    layer2_outputs(1851) <= not(layer1_outputs(2393));
    layer2_outputs(1852) <= not(layer1_outputs(568)) or (layer1_outputs(358));
    layer2_outputs(1853) <= '0';
    layer2_outputs(1854) <= not(layer1_outputs(1669));
    layer2_outputs(1855) <= (layer1_outputs(2494)) and not (layer1_outputs(1989));
    layer2_outputs(1856) <= layer1_outputs(825);
    layer2_outputs(1857) <= layer1_outputs(1712);
    layer2_outputs(1858) <= (layer1_outputs(582)) xor (layer1_outputs(817));
    layer2_outputs(1859) <= not((layer1_outputs(989)) or (layer1_outputs(1617)));
    layer2_outputs(1860) <= not(layer1_outputs(2350));
    layer2_outputs(1861) <= not(layer1_outputs(2076));
    layer2_outputs(1862) <= not(layer1_outputs(1561)) or (layer1_outputs(1376));
    layer2_outputs(1863) <= not((layer1_outputs(998)) and (layer1_outputs(2540)));
    layer2_outputs(1864) <= (layer1_outputs(30)) and not (layer1_outputs(1632));
    layer2_outputs(1865) <= not(layer1_outputs(821)) or (layer1_outputs(10));
    layer2_outputs(1866) <= not(layer1_outputs(1243));
    layer2_outputs(1867) <= not(layer1_outputs(292));
    layer2_outputs(1868) <= (layer1_outputs(177)) and not (layer1_outputs(87));
    layer2_outputs(1869) <= (layer1_outputs(2155)) and not (layer1_outputs(571));
    layer2_outputs(1870) <= (layer1_outputs(2167)) or (layer1_outputs(1860));
    layer2_outputs(1871) <= not(layer1_outputs(2429));
    layer2_outputs(1872) <= layer1_outputs(2422);
    layer2_outputs(1873) <= layer1_outputs(821);
    layer2_outputs(1874) <= not(layer1_outputs(1153));
    layer2_outputs(1875) <= (layer1_outputs(1297)) and not (layer1_outputs(239));
    layer2_outputs(1876) <= not(layer1_outputs(2169));
    layer2_outputs(1877) <= not((layer1_outputs(595)) and (layer1_outputs(586)));
    layer2_outputs(1878) <= (layer1_outputs(1118)) xor (layer1_outputs(412));
    layer2_outputs(1879) <= layer1_outputs(953);
    layer2_outputs(1880) <= not(layer1_outputs(2078));
    layer2_outputs(1881) <= layer1_outputs(2231);
    layer2_outputs(1882) <= layer1_outputs(95);
    layer2_outputs(1883) <= layer1_outputs(2330);
    layer2_outputs(1884) <= (layer1_outputs(734)) and not (layer1_outputs(568));
    layer2_outputs(1885) <= layer1_outputs(2118);
    layer2_outputs(1886) <= not(layer1_outputs(1563)) or (layer1_outputs(1732));
    layer2_outputs(1887) <= not(layer1_outputs(2362)) or (layer1_outputs(532));
    layer2_outputs(1888) <= not((layer1_outputs(608)) and (layer1_outputs(35)));
    layer2_outputs(1889) <= layer1_outputs(1566);
    layer2_outputs(1890) <= (layer1_outputs(274)) and (layer1_outputs(296));
    layer2_outputs(1891) <= not(layer1_outputs(6)) or (layer1_outputs(733));
    layer2_outputs(1892) <= (layer1_outputs(2107)) and not (layer1_outputs(1066));
    layer2_outputs(1893) <= not(layer1_outputs(1361)) or (layer1_outputs(567));
    layer2_outputs(1894) <= layer1_outputs(1126);
    layer2_outputs(1895) <= (layer1_outputs(1956)) or (layer1_outputs(1903));
    layer2_outputs(1896) <= (layer1_outputs(1149)) and not (layer1_outputs(1266));
    layer2_outputs(1897) <= (layer1_outputs(2226)) and not (layer1_outputs(2357));
    layer2_outputs(1898) <= layer1_outputs(1690);
    layer2_outputs(1899) <= (layer1_outputs(456)) and (layer1_outputs(804));
    layer2_outputs(1900) <= not((layer1_outputs(2241)) and (layer1_outputs(527)));
    layer2_outputs(1901) <= not(layer1_outputs(818));
    layer2_outputs(1902) <= not((layer1_outputs(706)) xor (layer1_outputs(790)));
    layer2_outputs(1903) <= (layer1_outputs(1521)) or (layer1_outputs(1990));
    layer2_outputs(1904) <= (layer1_outputs(2019)) and (layer1_outputs(522));
    layer2_outputs(1905) <= '1';
    layer2_outputs(1906) <= not((layer1_outputs(1471)) or (layer1_outputs(2223)));
    layer2_outputs(1907) <= not((layer1_outputs(95)) and (layer1_outputs(577)));
    layer2_outputs(1908) <= (layer1_outputs(2263)) and not (layer1_outputs(1624));
    layer2_outputs(1909) <= layer1_outputs(1317);
    layer2_outputs(1910) <= not(layer1_outputs(1153)) or (layer1_outputs(1068));
    layer2_outputs(1911) <= layer1_outputs(2149);
    layer2_outputs(1912) <= layer1_outputs(2212);
    layer2_outputs(1913) <= layer1_outputs(335);
    layer2_outputs(1914) <= layer1_outputs(2460);
    layer2_outputs(1915) <= (layer1_outputs(1349)) and not (layer1_outputs(2491));
    layer2_outputs(1916) <= not(layer1_outputs(2126));
    layer2_outputs(1917) <= not(layer1_outputs(409));
    layer2_outputs(1918) <= (layer1_outputs(2518)) and not (layer1_outputs(1233));
    layer2_outputs(1919) <= not((layer1_outputs(895)) or (layer1_outputs(2177)));
    layer2_outputs(1920) <= layer1_outputs(984);
    layer2_outputs(1921) <= not((layer1_outputs(3)) and (layer1_outputs(2303)));
    layer2_outputs(1922) <= layer1_outputs(1516);
    layer2_outputs(1923) <= not(layer1_outputs(933));
    layer2_outputs(1924) <= not((layer1_outputs(1663)) and (layer1_outputs(1331)));
    layer2_outputs(1925) <= layer1_outputs(1288);
    layer2_outputs(1926) <= (layer1_outputs(2297)) and not (layer1_outputs(2154));
    layer2_outputs(1927) <= (layer1_outputs(1514)) and (layer1_outputs(863));
    layer2_outputs(1928) <= (layer1_outputs(280)) and (layer1_outputs(2503));
    layer2_outputs(1929) <= layer1_outputs(2369);
    layer2_outputs(1930) <= not(layer1_outputs(139));
    layer2_outputs(1931) <= layer1_outputs(1212);
    layer2_outputs(1932) <= (layer1_outputs(733)) and not (layer1_outputs(1640));
    layer2_outputs(1933) <= not(layer1_outputs(647));
    layer2_outputs(1934) <= '0';
    layer2_outputs(1935) <= (layer1_outputs(2142)) xor (layer1_outputs(1667));
    layer2_outputs(1936) <= layer1_outputs(2542);
    layer2_outputs(1937) <= (layer1_outputs(1819)) and not (layer1_outputs(564));
    layer2_outputs(1938) <= layer1_outputs(396);
    layer2_outputs(1939) <= layer1_outputs(2232);
    layer2_outputs(1940) <= not((layer1_outputs(197)) and (layer1_outputs(2243)));
    layer2_outputs(1941) <= (layer1_outputs(793)) or (layer1_outputs(2179));
    layer2_outputs(1942) <= layer1_outputs(917);
    layer2_outputs(1943) <= (layer1_outputs(1365)) or (layer1_outputs(1100));
    layer2_outputs(1944) <= (layer1_outputs(1409)) or (layer1_outputs(295));
    layer2_outputs(1945) <= (layer1_outputs(1540)) or (layer1_outputs(2551));
    layer2_outputs(1946) <= not((layer1_outputs(2066)) and (layer1_outputs(162)));
    layer2_outputs(1947) <= layer1_outputs(1030);
    layer2_outputs(1948) <= not(layer1_outputs(1120));
    layer2_outputs(1949) <= not(layer1_outputs(1656)) or (layer1_outputs(2406));
    layer2_outputs(1950) <= layer1_outputs(1023);
    layer2_outputs(1951) <= not(layer1_outputs(1058));
    layer2_outputs(1952) <= (layer1_outputs(1798)) and not (layer1_outputs(1176));
    layer2_outputs(1953) <= not(layer1_outputs(1105));
    layer2_outputs(1954) <= (layer1_outputs(901)) or (layer1_outputs(343));
    layer2_outputs(1955) <= layer1_outputs(2456);
    layer2_outputs(1956) <= (layer1_outputs(1924)) or (layer1_outputs(397));
    layer2_outputs(1957) <= layer1_outputs(1818);
    layer2_outputs(1958) <= (layer1_outputs(1105)) and not (layer1_outputs(1168));
    layer2_outputs(1959) <= layer1_outputs(369);
    layer2_outputs(1960) <= '1';
    layer2_outputs(1961) <= not(layer1_outputs(1074)) or (layer1_outputs(2330));
    layer2_outputs(1962) <= (layer1_outputs(943)) and not (layer1_outputs(1551));
    layer2_outputs(1963) <= (layer1_outputs(2186)) and not (layer1_outputs(944));
    layer2_outputs(1964) <= (layer1_outputs(1550)) xor (layer1_outputs(2228));
    layer2_outputs(1965) <= not(layer1_outputs(2211));
    layer2_outputs(1966) <= layer1_outputs(2546);
    layer2_outputs(1967) <= (layer1_outputs(88)) or (layer1_outputs(2305));
    layer2_outputs(1968) <= (layer1_outputs(866)) and not (layer1_outputs(557));
    layer2_outputs(1969) <= layer1_outputs(1169);
    layer2_outputs(1970) <= not(layer1_outputs(325));
    layer2_outputs(1971) <= not(layer1_outputs(1405));
    layer2_outputs(1972) <= layer1_outputs(1838);
    layer2_outputs(1973) <= not((layer1_outputs(2032)) and (layer1_outputs(389)));
    layer2_outputs(1974) <= (layer1_outputs(2382)) and (layer1_outputs(1727));
    layer2_outputs(1975) <= (layer1_outputs(753)) and (layer1_outputs(684));
    layer2_outputs(1976) <= not(layer1_outputs(1680));
    layer2_outputs(1977) <= (layer1_outputs(1663)) and (layer1_outputs(2012));
    layer2_outputs(1978) <= layer1_outputs(868);
    layer2_outputs(1979) <= layer1_outputs(476);
    layer2_outputs(1980) <= layer1_outputs(2070);
    layer2_outputs(1981) <= not((layer1_outputs(2080)) and (layer1_outputs(428)));
    layer2_outputs(1982) <= not(layer1_outputs(978));
    layer2_outputs(1983) <= not(layer1_outputs(2372));
    layer2_outputs(1984) <= not((layer1_outputs(834)) or (layer1_outputs(2167)));
    layer2_outputs(1985) <= not(layer1_outputs(1829));
    layer2_outputs(1986) <= not((layer1_outputs(164)) and (layer1_outputs(1750)));
    layer2_outputs(1987) <= not(layer1_outputs(1386));
    layer2_outputs(1988) <= layer1_outputs(1060);
    layer2_outputs(1989) <= not((layer1_outputs(239)) or (layer1_outputs(1748)));
    layer2_outputs(1990) <= layer1_outputs(753);
    layer2_outputs(1991) <= not((layer1_outputs(1238)) xor (layer1_outputs(2219)));
    layer2_outputs(1992) <= (layer1_outputs(400)) and not (layer1_outputs(997));
    layer2_outputs(1993) <= layer1_outputs(2034);
    layer2_outputs(1994) <= not(layer1_outputs(5));
    layer2_outputs(1995) <= layer1_outputs(1216);
    layer2_outputs(1996) <= (layer1_outputs(1316)) and not (layer1_outputs(1764));
    layer2_outputs(1997) <= not((layer1_outputs(1864)) or (layer1_outputs(75)));
    layer2_outputs(1998) <= (layer1_outputs(1138)) and not (layer1_outputs(1786));
    layer2_outputs(1999) <= not(layer1_outputs(1820)) or (layer1_outputs(416));
    layer2_outputs(2000) <= not((layer1_outputs(826)) xor (layer1_outputs(512)));
    layer2_outputs(2001) <= not((layer1_outputs(1332)) xor (layer1_outputs(828)));
    layer2_outputs(2002) <= layer1_outputs(767);
    layer2_outputs(2003) <= not(layer1_outputs(1268));
    layer2_outputs(2004) <= (layer1_outputs(11)) and not (layer1_outputs(1963));
    layer2_outputs(2005) <= not((layer1_outputs(518)) or (layer1_outputs(1333)));
    layer2_outputs(2006) <= not((layer1_outputs(1935)) or (layer1_outputs(386)));
    layer2_outputs(2007) <= not(layer1_outputs(1970));
    layer2_outputs(2008) <= layer1_outputs(1794);
    layer2_outputs(2009) <= layer1_outputs(2010);
    layer2_outputs(2010) <= not(layer1_outputs(355));
    layer2_outputs(2011) <= not(layer1_outputs(960)) or (layer1_outputs(1613));
    layer2_outputs(2012) <= not(layer1_outputs(2140));
    layer2_outputs(2013) <= layer1_outputs(2069);
    layer2_outputs(2014) <= not(layer1_outputs(677));
    layer2_outputs(2015) <= not((layer1_outputs(89)) and (layer1_outputs(1508)));
    layer2_outputs(2016) <= (layer1_outputs(28)) or (layer1_outputs(942));
    layer2_outputs(2017) <= layer1_outputs(1857);
    layer2_outputs(2018) <= layer1_outputs(257);
    layer2_outputs(2019) <= (layer1_outputs(1032)) and not (layer1_outputs(2014));
    layer2_outputs(2020) <= layer1_outputs(2236);
    layer2_outputs(2021) <= not(layer1_outputs(1777)) or (layer1_outputs(2321));
    layer2_outputs(2022) <= not(layer1_outputs(1072));
    layer2_outputs(2023) <= not(layer1_outputs(2207));
    layer2_outputs(2024) <= layer1_outputs(1983);
    layer2_outputs(2025) <= layer1_outputs(1346);
    layer2_outputs(2026) <= not(layer1_outputs(1859));
    layer2_outputs(2027) <= (layer1_outputs(1558)) and not (layer1_outputs(1639));
    layer2_outputs(2028) <= layer1_outputs(1998);
    layer2_outputs(2029) <= layer1_outputs(1248);
    layer2_outputs(2030) <= not((layer1_outputs(932)) and (layer1_outputs(1065)));
    layer2_outputs(2031) <= not(layer1_outputs(707));
    layer2_outputs(2032) <= not(layer1_outputs(455));
    layer2_outputs(2033) <= (layer1_outputs(931)) and (layer1_outputs(313));
    layer2_outputs(2034) <= layer1_outputs(1544);
    layer2_outputs(2035) <= (layer1_outputs(2197)) or (layer1_outputs(63));
    layer2_outputs(2036) <= not(layer1_outputs(1431)) or (layer1_outputs(1186));
    layer2_outputs(2037) <= (layer1_outputs(294)) and not (layer1_outputs(858));
    layer2_outputs(2038) <= '1';
    layer2_outputs(2039) <= (layer1_outputs(697)) or (layer1_outputs(1227));
    layer2_outputs(2040) <= (layer1_outputs(1736)) and not (layer1_outputs(1782));
    layer2_outputs(2041) <= layer1_outputs(1159);
    layer2_outputs(2042) <= (layer1_outputs(2378)) and (layer1_outputs(618));
    layer2_outputs(2043) <= layer1_outputs(1927);
    layer2_outputs(2044) <= (layer1_outputs(1913)) xor (layer1_outputs(1271));
    layer2_outputs(2045) <= layer1_outputs(1807);
    layer2_outputs(2046) <= layer1_outputs(2098);
    layer2_outputs(2047) <= layer1_outputs(123);
    layer2_outputs(2048) <= layer1_outputs(1711);
    layer2_outputs(2049) <= (layer1_outputs(478)) or (layer1_outputs(250));
    layer2_outputs(2050) <= not(layer1_outputs(647));
    layer2_outputs(2051) <= (layer1_outputs(1590)) and not (layer1_outputs(1764));
    layer2_outputs(2052) <= not(layer1_outputs(2269)) or (layer1_outputs(1681));
    layer2_outputs(2053) <= '1';
    layer2_outputs(2054) <= (layer1_outputs(1520)) xor (layer1_outputs(422));
    layer2_outputs(2055) <= (layer1_outputs(1946)) and (layer1_outputs(2346));
    layer2_outputs(2056) <= not((layer1_outputs(1294)) or (layer1_outputs(137)));
    layer2_outputs(2057) <= not(layer1_outputs(1399));
    layer2_outputs(2058) <= not(layer1_outputs(193));
    layer2_outputs(2059) <= not(layer1_outputs(489)) or (layer1_outputs(963));
    layer2_outputs(2060) <= (layer1_outputs(1873)) or (layer1_outputs(2312));
    layer2_outputs(2061) <= (layer1_outputs(786)) and not (layer1_outputs(2030));
    layer2_outputs(2062) <= not((layer1_outputs(2474)) and (layer1_outputs(775)));
    layer2_outputs(2063) <= layer1_outputs(2490);
    layer2_outputs(2064) <= not((layer1_outputs(2159)) or (layer1_outputs(1691)));
    layer2_outputs(2065) <= layer1_outputs(852);
    layer2_outputs(2066) <= not((layer1_outputs(1368)) and (layer1_outputs(430)));
    layer2_outputs(2067) <= (layer1_outputs(1018)) and not (layer1_outputs(1952));
    layer2_outputs(2068) <= not(layer1_outputs(388));
    layer2_outputs(2069) <= not(layer1_outputs(2530)) or (layer1_outputs(1724));
    layer2_outputs(2070) <= not(layer1_outputs(1274)) or (layer1_outputs(784));
    layer2_outputs(2071) <= layer1_outputs(2021);
    layer2_outputs(2072) <= not((layer1_outputs(795)) and (layer1_outputs(1585)));
    layer2_outputs(2073) <= (layer1_outputs(589)) and (layer1_outputs(132));
    layer2_outputs(2074) <= not(layer1_outputs(1337));
    layer2_outputs(2075) <= not((layer1_outputs(2483)) or (layer1_outputs(1078)));
    layer2_outputs(2076) <= (layer1_outputs(993)) or (layer1_outputs(1963));
    layer2_outputs(2077) <= not(layer1_outputs(449)) or (layer1_outputs(888));
    layer2_outputs(2078) <= not(layer1_outputs(260));
    layer2_outputs(2079) <= not(layer1_outputs(906)) or (layer1_outputs(2218));
    layer2_outputs(2080) <= not(layer1_outputs(2207));
    layer2_outputs(2081) <= layer1_outputs(946);
    layer2_outputs(2082) <= not((layer1_outputs(2486)) xor (layer1_outputs(2387)));
    layer2_outputs(2083) <= (layer1_outputs(231)) and not (layer1_outputs(479));
    layer2_outputs(2084) <= not((layer1_outputs(237)) xor (layer1_outputs(15)));
    layer2_outputs(2085) <= not(layer1_outputs(1263));
    layer2_outputs(2086) <= '0';
    layer2_outputs(2087) <= '0';
    layer2_outputs(2088) <= (layer1_outputs(1996)) and not (layer1_outputs(108));
    layer2_outputs(2089) <= not(layer1_outputs(2518)) or (layer1_outputs(2127));
    layer2_outputs(2090) <= layer1_outputs(2279);
    layer2_outputs(2091) <= not(layer1_outputs(136));
    layer2_outputs(2092) <= '0';
    layer2_outputs(2093) <= (layer1_outputs(1305)) and (layer1_outputs(22));
    layer2_outputs(2094) <= not(layer1_outputs(2333)) or (layer1_outputs(2417));
    layer2_outputs(2095) <= not(layer1_outputs(899));
    layer2_outputs(2096) <= (layer1_outputs(2366)) and (layer1_outputs(1890));
    layer2_outputs(2097) <= (layer1_outputs(570)) and not (layer1_outputs(724));
    layer2_outputs(2098) <= not(layer1_outputs(374));
    layer2_outputs(2099) <= layer1_outputs(2456);
    layer2_outputs(2100) <= not((layer1_outputs(1501)) or (layer1_outputs(1005)));
    layer2_outputs(2101) <= layer1_outputs(1197);
    layer2_outputs(2102) <= not(layer1_outputs(191));
    layer2_outputs(2103) <= not(layer1_outputs(272)) or (layer1_outputs(2074));
    layer2_outputs(2104) <= not(layer1_outputs(1908));
    layer2_outputs(2105) <= layer1_outputs(2112);
    layer2_outputs(2106) <= not(layer1_outputs(919));
    layer2_outputs(2107) <= not(layer1_outputs(1655));
    layer2_outputs(2108) <= not((layer1_outputs(2283)) and (layer1_outputs(414)));
    layer2_outputs(2109) <= not((layer1_outputs(238)) or (layer1_outputs(1041)));
    layer2_outputs(2110) <= (layer1_outputs(1217)) and (layer1_outputs(76));
    layer2_outputs(2111) <= (layer1_outputs(1266)) xor (layer1_outputs(725));
    layer2_outputs(2112) <= not((layer1_outputs(727)) and (layer1_outputs(1918)));
    layer2_outputs(2113) <= not((layer1_outputs(2462)) and (layer1_outputs(2221)));
    layer2_outputs(2114) <= not((layer1_outputs(2213)) or (layer1_outputs(1445)));
    layer2_outputs(2115) <= (layer1_outputs(451)) and not (layer1_outputs(2553));
    layer2_outputs(2116) <= not(layer1_outputs(669));
    layer2_outputs(2117) <= not(layer1_outputs(1974)) or (layer1_outputs(731));
    layer2_outputs(2118) <= not(layer1_outputs(1394));
    layer2_outputs(2119) <= not(layer1_outputs(439));
    layer2_outputs(2120) <= not(layer1_outputs(812));
    layer2_outputs(2121) <= not(layer1_outputs(443));
    layer2_outputs(2122) <= not(layer1_outputs(276)) or (layer1_outputs(1083));
    layer2_outputs(2123) <= layer1_outputs(2199);
    layer2_outputs(2124) <= layer1_outputs(2104);
    layer2_outputs(2125) <= not(layer1_outputs(2464));
    layer2_outputs(2126) <= layer1_outputs(531);
    layer2_outputs(2127) <= (layer1_outputs(533)) or (layer1_outputs(1451));
    layer2_outputs(2128) <= layer1_outputs(803);
    layer2_outputs(2129) <= (layer1_outputs(9)) and (layer1_outputs(130));
    layer2_outputs(2130) <= layer1_outputs(2404);
    layer2_outputs(2131) <= '0';
    layer2_outputs(2132) <= layer1_outputs(2504);
    layer2_outputs(2133) <= not(layer1_outputs(256)) or (layer1_outputs(2074));
    layer2_outputs(2134) <= not(layer1_outputs(768)) or (layer1_outputs(1797));
    layer2_outputs(2135) <= (layer1_outputs(515)) or (layer1_outputs(2253));
    layer2_outputs(2136) <= not(layer1_outputs(1940));
    layer2_outputs(2137) <= not(layer1_outputs(381)) or (layer1_outputs(1079));
    layer2_outputs(2138) <= not((layer1_outputs(285)) and (layer1_outputs(819)));
    layer2_outputs(2139) <= layer1_outputs(907);
    layer2_outputs(2140) <= not(layer1_outputs(871));
    layer2_outputs(2141) <= layer1_outputs(1152);
    layer2_outputs(2142) <= (layer1_outputs(1975)) xor (layer1_outputs(333));
    layer2_outputs(2143) <= layer1_outputs(2002);
    layer2_outputs(2144) <= (layer1_outputs(1800)) and not (layer1_outputs(2394));
    layer2_outputs(2145) <= layer1_outputs(2239);
    layer2_outputs(2146) <= not(layer1_outputs(1812));
    layer2_outputs(2147) <= not((layer1_outputs(1703)) xor (layer1_outputs(827)));
    layer2_outputs(2148) <= not(layer1_outputs(1813));
    layer2_outputs(2149) <= layer1_outputs(1336);
    layer2_outputs(2150) <= not(layer1_outputs(2374)) or (layer1_outputs(2048));
    layer2_outputs(2151) <= not(layer1_outputs(157));
    layer2_outputs(2152) <= (layer1_outputs(1480)) xor (layer1_outputs(1213));
    layer2_outputs(2153) <= not(layer1_outputs(1337));
    layer2_outputs(2154) <= not(layer1_outputs(654)) or (layer1_outputs(2182));
    layer2_outputs(2155) <= not(layer1_outputs(432));
    layer2_outputs(2156) <= (layer1_outputs(1592)) and (layer1_outputs(402));
    layer2_outputs(2157) <= not((layer1_outputs(2043)) and (layer1_outputs(693)));
    layer2_outputs(2158) <= not(layer1_outputs(1388));
    layer2_outputs(2159) <= not(layer1_outputs(2477));
    layer2_outputs(2160) <= layer1_outputs(497);
    layer2_outputs(2161) <= not(layer1_outputs(364)) or (layer1_outputs(885));
    layer2_outputs(2162) <= (layer1_outputs(948)) and (layer1_outputs(2466));
    layer2_outputs(2163) <= layer1_outputs(667);
    layer2_outputs(2164) <= not(layer1_outputs(2535));
    layer2_outputs(2165) <= layer1_outputs(678);
    layer2_outputs(2166) <= not(layer1_outputs(2402));
    layer2_outputs(2167) <= not(layer1_outputs(2513)) or (layer1_outputs(849));
    layer2_outputs(2168) <= not((layer1_outputs(1538)) and (layer1_outputs(1428)));
    layer2_outputs(2169) <= (layer1_outputs(573)) or (layer1_outputs(649));
    layer2_outputs(2170) <= not(layer1_outputs(600));
    layer2_outputs(2171) <= (layer1_outputs(1995)) and (layer1_outputs(769));
    layer2_outputs(2172) <= layer1_outputs(2139);
    layer2_outputs(2173) <= not(layer1_outputs(1221));
    layer2_outputs(2174) <= not(layer1_outputs(315)) or (layer1_outputs(2467));
    layer2_outputs(2175) <= layer1_outputs(1696);
    layer2_outputs(2176) <= not(layer1_outputs(1134));
    layer2_outputs(2177) <= not(layer1_outputs(1883));
    layer2_outputs(2178) <= '0';
    layer2_outputs(2179) <= layer1_outputs(2432);
    layer2_outputs(2180) <= not(layer1_outputs(586));
    layer2_outputs(2181) <= not(layer1_outputs(2082));
    layer2_outputs(2182) <= not(layer1_outputs(1150)) or (layer1_outputs(1885));
    layer2_outputs(2183) <= not(layer1_outputs(1714));
    layer2_outputs(2184) <= (layer1_outputs(33)) or (layer1_outputs(1211));
    layer2_outputs(2185) <= not(layer1_outputs(133));
    layer2_outputs(2186) <= layer1_outputs(1738);
    layer2_outputs(2187) <= (layer1_outputs(1478)) and (layer1_outputs(430));
    layer2_outputs(2188) <= layer1_outputs(1497);
    layer2_outputs(2189) <= not((layer1_outputs(839)) or (layer1_outputs(1692)));
    layer2_outputs(2190) <= not(layer1_outputs(2247));
    layer2_outputs(2191) <= '1';
    layer2_outputs(2192) <= (layer1_outputs(1977)) and not (layer1_outputs(2320));
    layer2_outputs(2193) <= '1';
    layer2_outputs(2194) <= not(layer1_outputs(674)) or (layer1_outputs(1602));
    layer2_outputs(2195) <= not(layer1_outputs(1447));
    layer2_outputs(2196) <= (layer1_outputs(1648)) or (layer1_outputs(985));
    layer2_outputs(2197) <= layer1_outputs(1147);
    layer2_outputs(2198) <= not(layer1_outputs(1985));
    layer2_outputs(2199) <= '1';
    layer2_outputs(2200) <= (layer1_outputs(348)) and not (layer1_outputs(941));
    layer2_outputs(2201) <= not(layer1_outputs(198));
    layer2_outputs(2202) <= '0';
    layer2_outputs(2203) <= (layer1_outputs(407)) xor (layer1_outputs(770));
    layer2_outputs(2204) <= (layer1_outputs(2235)) and not (layer1_outputs(2458));
    layer2_outputs(2205) <= (layer1_outputs(746)) and not (layer1_outputs(2050));
    layer2_outputs(2206) <= not(layer1_outputs(2057)) or (layer1_outputs(1193));
    layer2_outputs(2207) <= not(layer1_outputs(986));
    layer2_outputs(2208) <= (layer1_outputs(2221)) and not (layer1_outputs(1968));
    layer2_outputs(2209) <= (layer1_outputs(1710)) or (layer1_outputs(506));
    layer2_outputs(2210) <= not(layer1_outputs(1028)) or (layer1_outputs(146));
    layer2_outputs(2211) <= layer1_outputs(412);
    layer2_outputs(2212) <= not(layer1_outputs(2533));
    layer2_outputs(2213) <= '1';
    layer2_outputs(2214) <= layer1_outputs(1412);
    layer2_outputs(2215) <= layer1_outputs(1923);
    layer2_outputs(2216) <= layer1_outputs(2370);
    layer2_outputs(2217) <= not((layer1_outputs(2447)) and (layer1_outputs(319)));
    layer2_outputs(2218) <= layer1_outputs(1278);
    layer2_outputs(2219) <= layer1_outputs(1011);
    layer2_outputs(2220) <= (layer1_outputs(423)) or (layer1_outputs(620));
    layer2_outputs(2221) <= not((layer1_outputs(1149)) and (layer1_outputs(1827)));
    layer2_outputs(2222) <= not((layer1_outputs(64)) or (layer1_outputs(2317)));
    layer2_outputs(2223) <= not(layer1_outputs(91));
    layer2_outputs(2224) <= layer1_outputs(625);
    layer2_outputs(2225) <= not((layer1_outputs(1747)) or (layer1_outputs(73)));
    layer2_outputs(2226) <= '1';
    layer2_outputs(2227) <= not(layer1_outputs(1286));
    layer2_outputs(2228) <= layer1_outputs(145);
    layer2_outputs(2229) <= not(layer1_outputs(359));
    layer2_outputs(2230) <= (layer1_outputs(2492)) and (layer1_outputs(1190));
    layer2_outputs(2231) <= '0';
    layer2_outputs(2232) <= (layer1_outputs(2263)) and not (layer1_outputs(2442));
    layer2_outputs(2233) <= layer1_outputs(363);
    layer2_outputs(2234) <= not(layer1_outputs(1273));
    layer2_outputs(2235) <= not((layer1_outputs(2084)) xor (layer1_outputs(339)));
    layer2_outputs(2236) <= (layer1_outputs(632)) and not (layer1_outputs(2308));
    layer2_outputs(2237) <= not((layer1_outputs(1437)) and (layer1_outputs(1031)));
    layer2_outputs(2238) <= not(layer1_outputs(699)) or (layer1_outputs(1291));
    layer2_outputs(2239) <= (layer1_outputs(1467)) or (layer1_outputs(2286));
    layer2_outputs(2240) <= not(layer1_outputs(765)) or (layer1_outputs(1772));
    layer2_outputs(2241) <= (layer1_outputs(1358)) or (layer1_outputs(1161));
    layer2_outputs(2242) <= '0';
    layer2_outputs(2243) <= not(layer1_outputs(1220));
    layer2_outputs(2244) <= not(layer1_outputs(2351)) or (layer1_outputs(1394));
    layer2_outputs(2245) <= not((layer1_outputs(331)) and (layer1_outputs(499)));
    layer2_outputs(2246) <= not(layer1_outputs(2245)) or (layer1_outputs(933));
    layer2_outputs(2247) <= not((layer1_outputs(1904)) or (layer1_outputs(45)));
    layer2_outputs(2248) <= not(layer1_outputs(258)) or (layer1_outputs(1781));
    layer2_outputs(2249) <= layer1_outputs(2168);
    layer2_outputs(2250) <= layer1_outputs(2216);
    layer2_outputs(2251) <= '1';
    layer2_outputs(2252) <= not(layer1_outputs(478));
    layer2_outputs(2253) <= not(layer1_outputs(2470));
    layer2_outputs(2254) <= layer1_outputs(277);
    layer2_outputs(2255) <= layer1_outputs(982);
    layer2_outputs(2256) <= not(layer1_outputs(623)) or (layer1_outputs(1411));
    layer2_outputs(2257) <= (layer1_outputs(883)) and (layer1_outputs(1151));
    layer2_outputs(2258) <= layer1_outputs(713);
    layer2_outputs(2259) <= layer1_outputs(227);
    layer2_outputs(2260) <= not(layer1_outputs(389));
    layer2_outputs(2261) <= (layer1_outputs(2238)) and not (layer1_outputs(1056));
    layer2_outputs(2262) <= layer1_outputs(181);
    layer2_outputs(2263) <= layer1_outputs(262);
    layer2_outputs(2264) <= not(layer1_outputs(1701));
    layer2_outputs(2265) <= (layer1_outputs(2035)) and not (layer1_outputs(1547));
    layer2_outputs(2266) <= (layer1_outputs(804)) or (layer1_outputs(2541));
    layer2_outputs(2267) <= not(layer1_outputs(302));
    layer2_outputs(2268) <= layer1_outputs(1326);
    layer2_outputs(2269) <= (layer1_outputs(743)) or (layer1_outputs(190));
    layer2_outputs(2270) <= layer1_outputs(965);
    layer2_outputs(2271) <= not(layer1_outputs(1058));
    layer2_outputs(2272) <= layer1_outputs(1202);
    layer2_outputs(2273) <= not((layer1_outputs(2521)) and (layer1_outputs(555)));
    layer2_outputs(2274) <= (layer1_outputs(1020)) and (layer1_outputs(1347));
    layer2_outputs(2275) <= not(layer1_outputs(1229));
    layer2_outputs(2276) <= (layer1_outputs(1933)) xor (layer1_outputs(1284));
    layer2_outputs(2277) <= not(layer1_outputs(1293));
    layer2_outputs(2278) <= not(layer1_outputs(2187));
    layer2_outputs(2279) <= not(layer1_outputs(2141)) or (layer1_outputs(2538));
    layer2_outputs(2280) <= layer1_outputs(1374);
    layer2_outputs(2281) <= (layer1_outputs(1490)) and not (layer1_outputs(737));
    layer2_outputs(2282) <= (layer1_outputs(833)) or (layer1_outputs(1979));
    layer2_outputs(2283) <= not(layer1_outputs(627));
    layer2_outputs(2284) <= layer1_outputs(1703);
    layer2_outputs(2285) <= not(layer1_outputs(1262)) or (layer1_outputs(806));
    layer2_outputs(2286) <= not(layer1_outputs(884));
    layer2_outputs(2287) <= layer1_outputs(1072);
    layer2_outputs(2288) <= not((layer1_outputs(1169)) or (layer1_outputs(2029)));
    layer2_outputs(2289) <= not((layer1_outputs(2502)) and (layer1_outputs(1801)));
    layer2_outputs(2290) <= not(layer1_outputs(26));
    layer2_outputs(2291) <= (layer1_outputs(212)) or (layer1_outputs(1889));
    layer2_outputs(2292) <= not(layer1_outputs(1685)) or (layer1_outputs(892));
    layer2_outputs(2293) <= not(layer1_outputs(2000));
    layer2_outputs(2294) <= not((layer1_outputs(2381)) and (layer1_outputs(2524)));
    layer2_outputs(2295) <= not(layer1_outputs(2356));
    layer2_outputs(2296) <= layer1_outputs(1560);
    layer2_outputs(2297) <= layer1_outputs(1850);
    layer2_outputs(2298) <= layer1_outputs(2047);
    layer2_outputs(2299) <= not(layer1_outputs(2248));
    layer2_outputs(2300) <= not(layer1_outputs(955)) or (layer1_outputs(2520));
    layer2_outputs(2301) <= '1';
    layer2_outputs(2302) <= (layer1_outputs(854)) and not (layer1_outputs(54));
    layer2_outputs(2303) <= (layer1_outputs(1989)) and not (layer1_outputs(2552));
    layer2_outputs(2304) <= not(layer1_outputs(1915));
    layer2_outputs(2305) <= not(layer1_outputs(2178));
    layer2_outputs(2306) <= layer1_outputs(664);
    layer2_outputs(2307) <= not(layer1_outputs(1523));
    layer2_outputs(2308) <= not(layer1_outputs(2008));
    layer2_outputs(2309) <= (layer1_outputs(867)) and not (layer1_outputs(2288));
    layer2_outputs(2310) <= '0';
    layer2_outputs(2311) <= not((layer1_outputs(956)) and (layer1_outputs(1698)));
    layer2_outputs(2312) <= layer1_outputs(106);
    layer2_outputs(2313) <= not(layer1_outputs(1163));
    layer2_outputs(2314) <= (layer1_outputs(273)) and not (layer1_outputs(1078));
    layer2_outputs(2315) <= not(layer1_outputs(1714));
    layer2_outputs(2316) <= not(layer1_outputs(714)) or (layer1_outputs(924));
    layer2_outputs(2317) <= not(layer1_outputs(1088)) or (layer1_outputs(1397));
    layer2_outputs(2318) <= layer1_outputs(854);
    layer2_outputs(2319) <= layer1_outputs(2299);
    layer2_outputs(2320) <= (layer1_outputs(862)) and not (layer1_outputs(707));
    layer2_outputs(2321) <= not((layer1_outputs(2152)) and (layer1_outputs(2093)));
    layer2_outputs(2322) <= not(layer1_outputs(1615));
    layer2_outputs(2323) <= layer1_outputs(1770);
    layer2_outputs(2324) <= layer1_outputs(708);
    layer2_outputs(2325) <= not(layer1_outputs(2102));
    layer2_outputs(2326) <= not(layer1_outputs(2124));
    layer2_outputs(2327) <= not(layer1_outputs(175)) or (layer1_outputs(996));
    layer2_outputs(2328) <= (layer1_outputs(1795)) or (layer1_outputs(361));
    layer2_outputs(2329) <= not((layer1_outputs(1389)) or (layer1_outputs(1341)));
    layer2_outputs(2330) <= not(layer1_outputs(1616));
    layer2_outputs(2331) <= layer1_outputs(1353);
    layer2_outputs(2332) <= (layer1_outputs(1886)) and not (layer1_outputs(1835));
    layer2_outputs(2333) <= not(layer1_outputs(1318));
    layer2_outputs(2334) <= layer1_outputs(1649);
    layer2_outputs(2335) <= not(layer1_outputs(2069));
    layer2_outputs(2336) <= layer1_outputs(72);
    layer2_outputs(2337) <= not((layer1_outputs(1309)) xor (layer1_outputs(702)));
    layer2_outputs(2338) <= (layer1_outputs(2068)) or (layer1_outputs(1515));
    layer2_outputs(2339) <= not((layer1_outputs(1393)) or (layer1_outputs(877)));
    layer2_outputs(2340) <= not(layer1_outputs(565));
    layer2_outputs(2341) <= layer1_outputs(1865);
    layer2_outputs(2342) <= not((layer1_outputs(1911)) and (layer1_outputs(2125)));
    layer2_outputs(2343) <= (layer1_outputs(1403)) and not (layer1_outputs(1036));
    layer2_outputs(2344) <= layer1_outputs(2031);
    layer2_outputs(2345) <= (layer1_outputs(395)) and not (layer1_outputs(2102));
    layer2_outputs(2346) <= not(layer1_outputs(1999));
    layer2_outputs(2347) <= layer1_outputs(2194);
    layer2_outputs(2348) <= not((layer1_outputs(813)) and (layer1_outputs(1941)));
    layer2_outputs(2349) <= not(layer1_outputs(1597)) or (layer1_outputs(2211));
    layer2_outputs(2350) <= not(layer1_outputs(278));
    layer2_outputs(2351) <= not(layer1_outputs(701));
    layer2_outputs(2352) <= layer1_outputs(637);
    layer2_outputs(2353) <= layer1_outputs(1002);
    layer2_outputs(2354) <= not(layer1_outputs(2149));
    layer2_outputs(2355) <= layer1_outputs(948);
    layer2_outputs(2356) <= (layer1_outputs(423)) or (layer1_outputs(1422));
    layer2_outputs(2357) <= (layer1_outputs(1718)) and not (layer1_outputs(2039));
    layer2_outputs(2358) <= not(layer1_outputs(1631));
    layer2_outputs(2359) <= not(layer1_outputs(1256));
    layer2_outputs(2360) <= (layer1_outputs(1350)) or (layer1_outputs(564));
    layer2_outputs(2361) <= layer1_outputs(322);
    layer2_outputs(2362) <= not((layer1_outputs(2509)) and (layer1_outputs(2016)));
    layer2_outputs(2363) <= not(layer1_outputs(1569));
    layer2_outputs(2364) <= '0';
    layer2_outputs(2365) <= not(layer1_outputs(1810));
    layer2_outputs(2366) <= layer1_outputs(2453);
    layer2_outputs(2367) <= layer1_outputs(496);
    layer2_outputs(2368) <= not(layer1_outputs(543));
    layer2_outputs(2369) <= not(layer1_outputs(388));
    layer2_outputs(2370) <= not(layer1_outputs(2254)) or (layer1_outputs(140));
    layer2_outputs(2371) <= layer1_outputs(2354);
    layer2_outputs(2372) <= (layer1_outputs(59)) and not (layer1_outputs(68));
    layer2_outputs(2373) <= not(layer1_outputs(1642));
    layer2_outputs(2374) <= not(layer1_outputs(1182));
    layer2_outputs(2375) <= not((layer1_outputs(2086)) or (layer1_outputs(2426)));
    layer2_outputs(2376) <= (layer1_outputs(1505)) or (layer1_outputs(1919));
    layer2_outputs(2377) <= layer1_outputs(180);
    layer2_outputs(2378) <= not((layer1_outputs(1772)) xor (layer1_outputs(4)));
    layer2_outputs(2379) <= layer1_outputs(1391);
    layer2_outputs(2380) <= not(layer1_outputs(2489)) or (layer1_outputs(1312));
    layer2_outputs(2381) <= not((layer1_outputs(597)) and (layer1_outputs(2488)));
    layer2_outputs(2382) <= (layer1_outputs(1457)) xor (layer1_outputs(1439));
    layer2_outputs(2383) <= (layer1_outputs(381)) and not (layer1_outputs(2442));
    layer2_outputs(2384) <= not(layer1_outputs(926));
    layer2_outputs(2385) <= not(layer1_outputs(811));
    layer2_outputs(2386) <= layer1_outputs(51);
    layer2_outputs(2387) <= layer1_outputs(1115);
    layer2_outputs(2388) <= (layer1_outputs(359)) or (layer1_outputs(1363));
    layer2_outputs(2389) <= layer1_outputs(2078);
    layer2_outputs(2390) <= layer1_outputs(1646);
    layer2_outputs(2391) <= (layer1_outputs(2227)) and (layer1_outputs(2208));
    layer2_outputs(2392) <= '1';
    layer2_outputs(2393) <= not((layer1_outputs(1861)) or (layer1_outputs(749)));
    layer2_outputs(2394) <= (layer1_outputs(648)) and not (layer1_outputs(401));
    layer2_outputs(2395) <= not(layer1_outputs(2543));
    layer2_outputs(2396) <= (layer1_outputs(1081)) and (layer1_outputs(1883));
    layer2_outputs(2397) <= not(layer1_outputs(1246)) or (layer1_outputs(923));
    layer2_outputs(2398) <= not(layer1_outputs(541)) or (layer1_outputs(1881));
    layer2_outputs(2399) <= layer1_outputs(1909);
    layer2_outputs(2400) <= not((layer1_outputs(1785)) xor (layer1_outputs(1321)));
    layer2_outputs(2401) <= not((layer1_outputs(701)) and (layer1_outputs(532)));
    layer2_outputs(2402) <= not((layer1_outputs(2070)) and (layer1_outputs(135)));
    layer2_outputs(2403) <= (layer1_outputs(156)) and not (layer1_outputs(520));
    layer2_outputs(2404) <= (layer1_outputs(1746)) and not (layer1_outputs(2514));
    layer2_outputs(2405) <= (layer1_outputs(1523)) and (layer1_outputs(1697));
    layer2_outputs(2406) <= not(layer1_outputs(864)) or (layer1_outputs(2174));
    layer2_outputs(2407) <= layer1_outputs(575);
    layer2_outputs(2408) <= layer1_outputs(2265);
    layer2_outputs(2409) <= layer1_outputs(1448);
    layer2_outputs(2410) <= layer1_outputs(2018);
    layer2_outputs(2411) <= layer1_outputs(1106);
    layer2_outputs(2412) <= not((layer1_outputs(2293)) and (layer1_outputs(1769)));
    layer2_outputs(2413) <= not(layer1_outputs(2183));
    layer2_outputs(2414) <= not((layer1_outputs(602)) xor (layer1_outputs(798)));
    layer2_outputs(2415) <= not(layer1_outputs(2372));
    layer2_outputs(2416) <= (layer1_outputs(881)) and (layer1_outputs(2046));
    layer2_outputs(2417) <= not(layer1_outputs(615));
    layer2_outputs(2418) <= layer1_outputs(2250);
    layer2_outputs(2419) <= layer1_outputs(685);
    layer2_outputs(2420) <= not((layer1_outputs(831)) or (layer1_outputs(2466)));
    layer2_outputs(2421) <= layer1_outputs(1777);
    layer2_outputs(2422) <= layer1_outputs(2258);
    layer2_outputs(2423) <= not((layer1_outputs(1672)) or (layer1_outputs(662)));
    layer2_outputs(2424) <= '1';
    layer2_outputs(2425) <= not((layer1_outputs(399)) or (layer1_outputs(1580)));
    layer2_outputs(2426) <= not(layer1_outputs(2472));
    layer2_outputs(2427) <= not(layer1_outputs(1666));
    layer2_outputs(2428) <= not((layer1_outputs(1906)) and (layer1_outputs(1514)));
    layer2_outputs(2429) <= not(layer1_outputs(784));
    layer2_outputs(2430) <= layer1_outputs(1899);
    layer2_outputs(2431) <= not(layer1_outputs(746));
    layer2_outputs(2432) <= layer1_outputs(2541);
    layer2_outputs(2433) <= not(layer1_outputs(440)) or (layer1_outputs(1309));
    layer2_outputs(2434) <= not((layer1_outputs(823)) or (layer1_outputs(1680)));
    layer2_outputs(2435) <= '0';
    layer2_outputs(2436) <= layer1_outputs(1572);
    layer2_outputs(2437) <= not(layer1_outputs(595));
    layer2_outputs(2438) <= (layer1_outputs(1172)) and (layer1_outputs(391));
    layer2_outputs(2439) <= layer1_outputs(1343);
    layer2_outputs(2440) <= not(layer1_outputs(2036)) or (layer1_outputs(970));
    layer2_outputs(2441) <= layer1_outputs(1614);
    layer2_outputs(2442) <= not(layer1_outputs(505)) or (layer1_outputs(652));
    layer2_outputs(2443) <= not(layer1_outputs(881));
    layer2_outputs(2444) <= not(layer1_outputs(658));
    layer2_outputs(2445) <= '0';
    layer2_outputs(2446) <= (layer1_outputs(1914)) xor (layer1_outputs(2392));
    layer2_outputs(2447) <= (layer1_outputs(1713)) and not (layer1_outputs(524));
    layer2_outputs(2448) <= not(layer1_outputs(546));
    layer2_outputs(2449) <= not(layer1_outputs(1969));
    layer2_outputs(2450) <= not((layer1_outputs(2420)) or (layer1_outputs(90)));
    layer2_outputs(2451) <= not(layer1_outputs(1655)) or (layer1_outputs(1385));
    layer2_outputs(2452) <= not((layer1_outputs(848)) and (layer1_outputs(1549)));
    layer2_outputs(2453) <= layer1_outputs(312);
    layer2_outputs(2454) <= layer1_outputs(103);
    layer2_outputs(2455) <= not(layer1_outputs(2246));
    layer2_outputs(2456) <= not(layer1_outputs(323));
    layer2_outputs(2457) <= layer1_outputs(57);
    layer2_outputs(2458) <= not((layer1_outputs(639)) or (layer1_outputs(2439)));
    layer2_outputs(2459) <= (layer1_outputs(2018)) and (layer1_outputs(1576));
    layer2_outputs(2460) <= not((layer1_outputs(451)) xor (layer1_outputs(1301)));
    layer2_outputs(2461) <= not((layer1_outputs(1235)) and (layer1_outputs(2548)));
    layer2_outputs(2462) <= layer1_outputs(2023);
    layer2_outputs(2463) <= not(layer1_outputs(1911)) or (layer1_outputs(1562));
    layer2_outputs(2464) <= (layer1_outputs(2243)) and not (layer1_outputs(695));
    layer2_outputs(2465) <= not(layer1_outputs(1607));
    layer2_outputs(2466) <= layer1_outputs(468);
    layer2_outputs(2467) <= not(layer1_outputs(991));
    layer2_outputs(2468) <= (layer1_outputs(284)) and not (layer1_outputs(2464));
    layer2_outputs(2469) <= not(layer1_outputs(1537)) or (layer1_outputs(837));
    layer2_outputs(2470) <= not((layer1_outputs(2398)) or (layer1_outputs(1463)));
    layer2_outputs(2471) <= not(layer1_outputs(2268));
    layer2_outputs(2472) <= (layer1_outputs(140)) and not (layer1_outputs(816));
    layer2_outputs(2473) <= (layer1_outputs(940)) and (layer1_outputs(2277));
    layer2_outputs(2474) <= not(layer1_outputs(2212));
    layer2_outputs(2475) <= not(layer1_outputs(1172)) or (layer1_outputs(2361));
    layer2_outputs(2476) <= not(layer1_outputs(663));
    layer2_outputs(2477) <= layer1_outputs(1601);
    layer2_outputs(2478) <= not(layer1_outputs(1828));
    layer2_outputs(2479) <= not(layer1_outputs(1969));
    layer2_outputs(2480) <= layer1_outputs(680);
    layer2_outputs(2481) <= (layer1_outputs(823)) and (layer1_outputs(709));
    layer2_outputs(2482) <= not((layer1_outputs(1412)) and (layer1_outputs(636)));
    layer2_outputs(2483) <= (layer1_outputs(1052)) and not (layer1_outputs(744));
    layer2_outputs(2484) <= not((layer1_outputs(112)) and (layer1_outputs(509)));
    layer2_outputs(2485) <= layer1_outputs(829);
    layer2_outputs(2486) <= not(layer1_outputs(1071));
    layer2_outputs(2487) <= (layer1_outputs(1496)) and not (layer1_outputs(1210));
    layer2_outputs(2488) <= layer1_outputs(1108);
    layer2_outputs(2489) <= (layer1_outputs(1413)) and (layer1_outputs(306));
    layer2_outputs(2490) <= not(layer1_outputs(1223));
    layer2_outputs(2491) <= not(layer1_outputs(1525)) or (layer1_outputs(2447));
    layer2_outputs(2492) <= (layer1_outputs(1214)) and not (layer1_outputs(560));
    layer2_outputs(2493) <= (layer1_outputs(1487)) and not (layer1_outputs(1654));
    layer2_outputs(2494) <= (layer1_outputs(1798)) and not (layer1_outputs(2126));
    layer2_outputs(2495) <= not(layer1_outputs(287)) or (layer1_outputs(644));
    layer2_outputs(2496) <= not((layer1_outputs(648)) or (layer1_outputs(1768)));
    layer2_outputs(2497) <= not(layer1_outputs(2196));
    layer2_outputs(2498) <= '1';
    layer2_outputs(2499) <= (layer1_outputs(2023)) and not (layer1_outputs(33));
    layer2_outputs(2500) <= not(layer1_outputs(277));
    layer2_outputs(2501) <= layer1_outputs(1097);
    layer2_outputs(2502) <= layer1_outputs(1397);
    layer2_outputs(2503) <= (layer1_outputs(1684)) and (layer1_outputs(1662));
    layer2_outputs(2504) <= layer1_outputs(1727);
    layer2_outputs(2505) <= (layer1_outputs(380)) or (layer1_outputs(1927));
    layer2_outputs(2506) <= (layer1_outputs(421)) and not (layer1_outputs(527));
    layer2_outputs(2507) <= not(layer1_outputs(1946));
    layer2_outputs(2508) <= not(layer1_outputs(310)) or (layer1_outputs(1372));
    layer2_outputs(2509) <= layer1_outputs(426);
    layer2_outputs(2510) <= not(layer1_outputs(2537));
    layer2_outputs(2511) <= layer1_outputs(2229);
    layer2_outputs(2512) <= (layer1_outputs(2364)) xor (layer1_outputs(716));
    layer2_outputs(2513) <= (layer1_outputs(1552)) and not (layer1_outputs(70));
    layer2_outputs(2514) <= layer1_outputs(1818);
    layer2_outputs(2515) <= not((layer1_outputs(236)) or (layer1_outputs(1022)));
    layer2_outputs(2516) <= not(layer1_outputs(23)) or (layer1_outputs(2380));
    layer2_outputs(2517) <= (layer1_outputs(1674)) and not (layer1_outputs(2491));
    layer2_outputs(2518) <= not(layer1_outputs(1179));
    layer2_outputs(2519) <= not(layer1_outputs(2191)) or (layer1_outputs(283));
    layer2_outputs(2520) <= (layer1_outputs(60)) and not (layer1_outputs(1282));
    layer2_outputs(2521) <= not(layer1_outputs(603));
    layer2_outputs(2522) <= layer1_outputs(1716);
    layer2_outputs(2523) <= '1';
    layer2_outputs(2524) <= not(layer1_outputs(1804));
    layer2_outputs(2525) <= layer1_outputs(897);
    layer2_outputs(2526) <= not((layer1_outputs(1986)) and (layer1_outputs(2357)));
    layer2_outputs(2527) <= (layer1_outputs(378)) and not (layer1_outputs(248));
    layer2_outputs(2528) <= (layer1_outputs(2302)) and not (layer1_outputs(2118));
    layer2_outputs(2529) <= not((layer1_outputs(1536)) or (layer1_outputs(2532)));
    layer2_outputs(2530) <= (layer1_outputs(261)) and not (layer1_outputs(138));
    layer2_outputs(2531) <= layer1_outputs(818);
    layer2_outputs(2532) <= layer1_outputs(2075);
    layer2_outputs(2533) <= layer1_outputs(509);
    layer2_outputs(2534) <= not(layer1_outputs(92));
    layer2_outputs(2535) <= not(layer1_outputs(517));
    layer2_outputs(2536) <= not(layer1_outputs(2135));
    layer2_outputs(2537) <= (layer1_outputs(2326)) and not (layer1_outputs(490));
    layer2_outputs(2538) <= not(layer1_outputs(1026));
    layer2_outputs(2539) <= not(layer1_outputs(1385));
    layer2_outputs(2540) <= layer1_outputs(984);
    layer2_outputs(2541) <= layer1_outputs(332);
    layer2_outputs(2542) <= not(layer1_outputs(1570));
    layer2_outputs(2543) <= not(layer1_outputs(805));
    layer2_outputs(2544) <= not(layer1_outputs(1356));
    layer2_outputs(2545) <= (layer1_outputs(2184)) and not (layer1_outputs(56));
    layer2_outputs(2546) <= layer1_outputs(1870);
    layer2_outputs(2547) <= not(layer1_outputs(1671));
    layer2_outputs(2548) <= not(layer1_outputs(1370));
    layer2_outputs(2549) <= layer1_outputs(1934);
    layer2_outputs(2550) <= (layer1_outputs(1239)) or (layer1_outputs(503));
    layer2_outputs(2551) <= layer1_outputs(920);
    layer2_outputs(2552) <= not(layer1_outputs(1251));
    layer2_outputs(2553) <= (layer1_outputs(2503)) and (layer1_outputs(121));
    layer2_outputs(2554) <= not((layer1_outputs(534)) or (layer1_outputs(2237)));
    layer2_outputs(2555) <= not((layer1_outputs(2210)) xor (layer1_outputs(1500)));
    layer2_outputs(2556) <= layer1_outputs(787);
    layer2_outputs(2557) <= layer1_outputs(1495);
    layer2_outputs(2558) <= (layer1_outputs(1182)) or (layer1_outputs(2085));
    layer2_outputs(2559) <= layer1_outputs(1992);
    outputs(0) <= (layer2_outputs(1868)) and not (layer2_outputs(192));
    outputs(1) <= not(layer2_outputs(624));
    outputs(2) <= not((layer2_outputs(1092)) or (layer2_outputs(1505)));
    outputs(3) <= layer2_outputs(587);
    outputs(4) <= layer2_outputs(1477);
    outputs(5) <= (layer2_outputs(1840)) and (layer2_outputs(83));
    outputs(6) <= layer2_outputs(2510);
    outputs(7) <= layer2_outputs(793);
    outputs(8) <= layer2_outputs(414);
    outputs(9) <= not(layer2_outputs(1153));
    outputs(10) <= not((layer2_outputs(1025)) or (layer2_outputs(1070)));
    outputs(11) <= layer2_outputs(480);
    outputs(12) <= not((layer2_outputs(1086)) or (layer2_outputs(1135)));
    outputs(13) <= not(layer2_outputs(862));
    outputs(14) <= (layer2_outputs(940)) and not (layer2_outputs(1975));
    outputs(15) <= not(layer2_outputs(1452));
    outputs(16) <= layer2_outputs(2365);
    outputs(17) <= not(layer2_outputs(1554));
    outputs(18) <= not((layer2_outputs(1140)) and (layer2_outputs(1941)));
    outputs(19) <= not(layer2_outputs(1958));
    outputs(20) <= layer2_outputs(620);
    outputs(21) <= not(layer2_outputs(1939));
    outputs(22) <= (layer2_outputs(698)) and not (layer2_outputs(603));
    outputs(23) <= not(layer2_outputs(1174)) or (layer2_outputs(1434));
    outputs(24) <= layer2_outputs(278);
    outputs(25) <= layer2_outputs(1702);
    outputs(26) <= layer2_outputs(2554);
    outputs(27) <= not(layer2_outputs(2412));
    outputs(28) <= not(layer2_outputs(1536));
    outputs(29) <= layer2_outputs(2272);
    outputs(30) <= not(layer2_outputs(1822));
    outputs(31) <= layer2_outputs(544);
    outputs(32) <= (layer2_outputs(2146)) and not (layer2_outputs(1242));
    outputs(33) <= layer2_outputs(1023);
    outputs(34) <= layer2_outputs(2029);
    outputs(35) <= (layer2_outputs(2463)) and not (layer2_outputs(606));
    outputs(36) <= not((layer2_outputs(292)) or (layer2_outputs(2082)));
    outputs(37) <= not(layer2_outputs(64));
    outputs(38) <= not(layer2_outputs(1654));
    outputs(39) <= not(layer2_outputs(832));
    outputs(40) <= not(layer2_outputs(2550));
    outputs(41) <= not(layer2_outputs(288));
    outputs(42) <= layer2_outputs(359);
    outputs(43) <= not(layer2_outputs(727));
    outputs(44) <= (layer2_outputs(647)) and not (layer2_outputs(1269));
    outputs(45) <= not(layer2_outputs(927));
    outputs(46) <= (layer2_outputs(1137)) and (layer2_outputs(2031));
    outputs(47) <= not(layer2_outputs(2249));
    outputs(48) <= (layer2_outputs(1150)) and (layer2_outputs(1382));
    outputs(49) <= layer2_outputs(203);
    outputs(50) <= (layer2_outputs(310)) or (layer2_outputs(1209));
    outputs(51) <= not(layer2_outputs(1829));
    outputs(52) <= not(layer2_outputs(571));
    outputs(53) <= not((layer2_outputs(1083)) xor (layer2_outputs(465)));
    outputs(54) <= layer2_outputs(2375);
    outputs(55) <= not((layer2_outputs(2440)) and (layer2_outputs(220)));
    outputs(56) <= layer2_outputs(2484);
    outputs(57) <= not(layer2_outputs(1449)) or (layer2_outputs(282));
    outputs(58) <= not(layer2_outputs(1565));
    outputs(59) <= layer2_outputs(948);
    outputs(60) <= (layer2_outputs(1627)) or (layer2_outputs(1644));
    outputs(61) <= (layer2_outputs(703)) xor (layer2_outputs(2441));
    outputs(62) <= not(layer2_outputs(733));
    outputs(63) <= layer2_outputs(205);
    outputs(64) <= not(layer2_outputs(644));
    outputs(65) <= not((layer2_outputs(867)) or (layer2_outputs(1)));
    outputs(66) <= (layer2_outputs(2044)) and (layer2_outputs(285));
    outputs(67) <= not(layer2_outputs(2431));
    outputs(68) <= not(layer2_outputs(932));
    outputs(69) <= layer2_outputs(654);
    outputs(70) <= not(layer2_outputs(2035));
    outputs(71) <= layer2_outputs(1910);
    outputs(72) <= (layer2_outputs(805)) and not (layer2_outputs(2466));
    outputs(73) <= (layer2_outputs(1451)) and (layer2_outputs(2089));
    outputs(74) <= not(layer2_outputs(2347)) or (layer2_outputs(944));
    outputs(75) <= layer2_outputs(1198);
    outputs(76) <= layer2_outputs(1218);
    outputs(77) <= not(layer2_outputs(1000));
    outputs(78) <= not(layer2_outputs(1478));
    outputs(79) <= (layer2_outputs(1693)) and not (layer2_outputs(935));
    outputs(80) <= not(layer2_outputs(930));
    outputs(81) <= layer2_outputs(1056);
    outputs(82) <= not(layer2_outputs(1456)) or (layer2_outputs(732));
    outputs(83) <= layer2_outputs(433);
    outputs(84) <= not(layer2_outputs(1904));
    outputs(85) <= layer2_outputs(1860);
    outputs(86) <= layer2_outputs(2071);
    outputs(87) <= (layer2_outputs(1074)) and not (layer2_outputs(1026));
    outputs(88) <= not(layer2_outputs(1298));
    outputs(89) <= (layer2_outputs(2025)) or (layer2_outputs(1305));
    outputs(90) <= layer2_outputs(358);
    outputs(91) <= (layer2_outputs(1367)) and not (layer2_outputs(2492));
    outputs(92) <= layer2_outputs(1421);
    outputs(93) <= not(layer2_outputs(1814));
    outputs(94) <= layer2_outputs(1195);
    outputs(95) <= (layer2_outputs(861)) and (layer2_outputs(1739));
    outputs(96) <= layer2_outputs(620);
    outputs(97) <= layer2_outputs(778);
    outputs(98) <= not((layer2_outputs(521)) and (layer2_outputs(2134)));
    outputs(99) <= layer2_outputs(2349);
    outputs(100) <= layer2_outputs(2484);
    outputs(101) <= not(layer2_outputs(1882));
    outputs(102) <= not((layer2_outputs(787)) xor (layer2_outputs(1652)));
    outputs(103) <= not((layer2_outputs(380)) xor (layer2_outputs(1045)));
    outputs(104) <= not(layer2_outputs(407)) or (layer2_outputs(718));
    outputs(105) <= (layer2_outputs(1265)) and not (layer2_outputs(211));
    outputs(106) <= layer2_outputs(5);
    outputs(107) <= not(layer2_outputs(1227));
    outputs(108) <= not(layer2_outputs(2417));
    outputs(109) <= not(layer2_outputs(2539));
    outputs(110) <= not(layer2_outputs(1773));
    outputs(111) <= layer2_outputs(214);
    outputs(112) <= (layer2_outputs(1225)) and not (layer2_outputs(1362));
    outputs(113) <= not(layer2_outputs(1142)) or (layer2_outputs(2025));
    outputs(114) <= not(layer2_outputs(999)) or (layer2_outputs(1533));
    outputs(115) <= layer2_outputs(1718);
    outputs(116) <= not(layer2_outputs(916));
    outputs(117) <= not(layer2_outputs(511));
    outputs(118) <= layer2_outputs(1266);
    outputs(119) <= not((layer2_outputs(1464)) or (layer2_outputs(1663)));
    outputs(120) <= (layer2_outputs(1625)) and not (layer2_outputs(1360));
    outputs(121) <= not(layer2_outputs(2246));
    outputs(122) <= layer2_outputs(2055);
    outputs(123) <= (layer2_outputs(1836)) and not (layer2_outputs(1406));
    outputs(124) <= not((layer2_outputs(488)) or (layer2_outputs(993)));
    outputs(125) <= layer2_outputs(2397);
    outputs(126) <= layer2_outputs(2205);
    outputs(127) <= not(layer2_outputs(789));
    outputs(128) <= not(layer2_outputs(2491)) or (layer2_outputs(1543));
    outputs(129) <= layer2_outputs(1876);
    outputs(130) <= layer2_outputs(813);
    outputs(131) <= layer2_outputs(950);
    outputs(132) <= (layer2_outputs(1852)) xor (layer2_outputs(1631));
    outputs(133) <= not(layer2_outputs(775));
    outputs(134) <= (layer2_outputs(1331)) xor (layer2_outputs(1623));
    outputs(135) <= layer2_outputs(1419);
    outputs(136) <= not((layer2_outputs(682)) or (layer2_outputs(2233)));
    outputs(137) <= layer2_outputs(538);
    outputs(138) <= layer2_outputs(1313);
    outputs(139) <= not(layer2_outputs(891)) or (layer2_outputs(360));
    outputs(140) <= layer2_outputs(436);
    outputs(141) <= not(layer2_outputs(1072));
    outputs(142) <= not(layer2_outputs(16));
    outputs(143) <= layer2_outputs(1189);
    outputs(144) <= not(layer2_outputs(1995));
    outputs(145) <= not(layer2_outputs(1920)) or (layer2_outputs(616));
    outputs(146) <= not((layer2_outputs(1615)) xor (layer2_outputs(1095)));
    outputs(147) <= not((layer2_outputs(535)) or (layer2_outputs(1402)));
    outputs(148) <= layer2_outputs(453);
    outputs(149) <= not(layer2_outputs(782));
    outputs(150) <= not(layer2_outputs(457));
    outputs(151) <= not(layer2_outputs(776));
    outputs(152) <= (layer2_outputs(299)) and (layer2_outputs(17));
    outputs(153) <= layer2_outputs(1210);
    outputs(154) <= not((layer2_outputs(953)) and (layer2_outputs(421)));
    outputs(155) <= not(layer2_outputs(1603));
    outputs(156) <= not(layer2_outputs(379));
    outputs(157) <= not(layer2_outputs(1454));
    outputs(158) <= (layer2_outputs(2471)) and (layer2_outputs(628));
    outputs(159) <= (layer2_outputs(1966)) and not (layer2_outputs(1289));
    outputs(160) <= layer2_outputs(18);
    outputs(161) <= not(layer2_outputs(7));
    outputs(162) <= not((layer2_outputs(1275)) xor (layer2_outputs(1588)));
    outputs(163) <= not(layer2_outputs(1541));
    outputs(164) <= not(layer2_outputs(1303));
    outputs(165) <= (layer2_outputs(1198)) or (layer2_outputs(2002));
    outputs(166) <= not(layer2_outputs(2431));
    outputs(167) <= not(layer2_outputs(1001));
    outputs(168) <= (layer2_outputs(1714)) and not (layer2_outputs(1774));
    outputs(169) <= not(layer2_outputs(1066));
    outputs(170) <= not(layer2_outputs(29));
    outputs(171) <= layer2_outputs(1911);
    outputs(172) <= not(layer2_outputs(573));
    outputs(173) <= layer2_outputs(1521);
    outputs(174) <= not(layer2_outputs(1334));
    outputs(175) <= layer2_outputs(1326);
    outputs(176) <= layer2_outputs(895);
    outputs(177) <= layer2_outputs(980);
    outputs(178) <= (layer2_outputs(2059)) and not (layer2_outputs(576));
    outputs(179) <= not((layer2_outputs(600)) or (layer2_outputs(796)));
    outputs(180) <= not(layer2_outputs(841));
    outputs(181) <= (layer2_outputs(1706)) or (layer2_outputs(2204));
    outputs(182) <= layer2_outputs(142);
    outputs(183) <= not((layer2_outputs(1085)) and (layer2_outputs(1337)));
    outputs(184) <= layer2_outputs(1719);
    outputs(185) <= layer2_outputs(157);
    outputs(186) <= not(layer2_outputs(1287));
    outputs(187) <= layer2_outputs(1170);
    outputs(188) <= (layer2_outputs(2366)) xor (layer2_outputs(2352));
    outputs(189) <= layer2_outputs(2286);
    outputs(190) <= not(layer2_outputs(750));
    outputs(191) <= layer2_outputs(1033);
    outputs(192) <= (layer2_outputs(301)) and (layer2_outputs(2245));
    outputs(193) <= not(layer2_outputs(2106));
    outputs(194) <= not(layer2_outputs(2109));
    outputs(195) <= (layer2_outputs(503)) and not (layer2_outputs(1353));
    outputs(196) <= layer2_outputs(1953);
    outputs(197) <= not(layer2_outputs(1580));
    outputs(198) <= (layer2_outputs(2326)) and not (layer2_outputs(2477));
    outputs(199) <= (layer2_outputs(1600)) and not (layer2_outputs(1884));
    outputs(200) <= (layer2_outputs(1093)) and not (layer2_outputs(1089));
    outputs(201) <= not((layer2_outputs(1429)) xor (layer2_outputs(346)));
    outputs(202) <= not(layer2_outputs(908));
    outputs(203) <= layer2_outputs(1030);
    outputs(204) <= not(layer2_outputs(790));
    outputs(205) <= layer2_outputs(1171);
    outputs(206) <= (layer2_outputs(2184)) and not (layer2_outputs(156));
    outputs(207) <= not(layer2_outputs(2239));
    outputs(208) <= not(layer2_outputs(14));
    outputs(209) <= layer2_outputs(1911);
    outputs(210) <= layer2_outputs(1558);
    outputs(211) <= not(layer2_outputs(565));
    outputs(212) <= not(layer2_outputs(1425));
    outputs(213) <= (layer2_outputs(605)) and not (layer2_outputs(759));
    outputs(214) <= layer2_outputs(2314);
    outputs(215) <= not(layer2_outputs(1639));
    outputs(216) <= not(layer2_outputs(1010));
    outputs(217) <= not(layer2_outputs(1183));
    outputs(218) <= layer2_outputs(2010);
    outputs(219) <= layer2_outputs(2432);
    outputs(220) <= (layer2_outputs(2075)) and not (layer2_outputs(229));
    outputs(221) <= layer2_outputs(435);
    outputs(222) <= layer2_outputs(1723);
    outputs(223) <= layer2_outputs(2481);
    outputs(224) <= layer2_outputs(896);
    outputs(225) <= not(layer2_outputs(1191));
    outputs(226) <= not(layer2_outputs(316));
    outputs(227) <= not(layer2_outputs(174));
    outputs(228) <= not(layer2_outputs(1990));
    outputs(229) <= layer2_outputs(1723);
    outputs(230) <= not(layer2_outputs(1662));
    outputs(231) <= layer2_outputs(2500);
    outputs(232) <= not(layer2_outputs(662)) or (layer2_outputs(415));
    outputs(233) <= not(layer2_outputs(2522));
    outputs(234) <= layer2_outputs(1614);
    outputs(235) <= layer2_outputs(1344);
    outputs(236) <= layer2_outputs(1768);
    outputs(237) <= layer2_outputs(2195);
    outputs(238) <= layer2_outputs(2141);
    outputs(239) <= (layer2_outputs(2341)) and not (layer2_outputs(1642));
    outputs(240) <= (layer2_outputs(2391)) xor (layer2_outputs(2102));
    outputs(241) <= not(layer2_outputs(562));
    outputs(242) <= not(layer2_outputs(1598));
    outputs(243) <= not(layer2_outputs(898));
    outputs(244) <= (layer2_outputs(1394)) and not (layer2_outputs(537));
    outputs(245) <= not(layer2_outputs(601));
    outputs(246) <= (layer2_outputs(1529)) and (layer2_outputs(302));
    outputs(247) <= layer2_outputs(588);
    outputs(248) <= (layer2_outputs(2329)) or (layer2_outputs(2294));
    outputs(249) <= not(layer2_outputs(2359));
    outputs(250) <= not(layer2_outputs(241));
    outputs(251) <= (layer2_outputs(366)) and not (layer2_outputs(388));
    outputs(252) <= layer2_outputs(638);
    outputs(253) <= not((layer2_outputs(2277)) or (layer2_outputs(2081)));
    outputs(254) <= not(layer2_outputs(947));
    outputs(255) <= not(layer2_outputs(2419));
    outputs(256) <= not((layer2_outputs(1065)) or (layer2_outputs(2206)));
    outputs(257) <= not((layer2_outputs(786)) or (layer2_outputs(913)));
    outputs(258) <= (layer2_outputs(1524)) xor (layer2_outputs(793));
    outputs(259) <= (layer2_outputs(1817)) and not (layer2_outputs(2305));
    outputs(260) <= not((layer2_outputs(681)) or (layer2_outputs(934)));
    outputs(261) <= (layer2_outputs(63)) and not (layer2_outputs(2234));
    outputs(262) <= (layer2_outputs(2185)) and not (layer2_outputs(221));
    outputs(263) <= layer2_outputs(1984);
    outputs(264) <= (layer2_outputs(851)) and (layer2_outputs(336));
    outputs(265) <= layer2_outputs(1856);
    outputs(266) <= not(layer2_outputs(1468)) or (layer2_outputs(706));
    outputs(267) <= layer2_outputs(341);
    outputs(268) <= not((layer2_outputs(2079)) or (layer2_outputs(2175)));
    outputs(269) <= not(layer2_outputs(1649));
    outputs(270) <= not(layer2_outputs(2282));
    outputs(271) <= not((layer2_outputs(1932)) or (layer2_outputs(43)));
    outputs(272) <= layer2_outputs(2529);
    outputs(273) <= not(layer2_outputs(24));
    outputs(274) <= not(layer2_outputs(812));
    outputs(275) <= not(layer2_outputs(1831));
    outputs(276) <= not((layer2_outputs(1412)) or (layer2_outputs(411)));
    outputs(277) <= not(layer2_outputs(734));
    outputs(278) <= (layer2_outputs(306)) and (layer2_outputs(524));
    outputs(279) <= (layer2_outputs(2164)) and not (layer2_outputs(2453));
    outputs(280) <= not(layer2_outputs(1251));
    outputs(281) <= not((layer2_outputs(1049)) or (layer2_outputs(824)));
    outputs(282) <= (layer2_outputs(2388)) xor (layer2_outputs(76));
    outputs(283) <= not((layer2_outputs(227)) or (layer2_outputs(900)));
    outputs(284) <= not(layer2_outputs(301));
    outputs(285) <= not((layer2_outputs(2015)) or (layer2_outputs(1082)));
    outputs(286) <= (layer2_outputs(1147)) and not (layer2_outputs(48));
    outputs(287) <= not((layer2_outputs(94)) or (layer2_outputs(160)));
    outputs(288) <= layer2_outputs(791);
    outputs(289) <= layer2_outputs(1595);
    outputs(290) <= layer2_outputs(120);
    outputs(291) <= not(layer2_outputs(1534));
    outputs(292) <= (layer2_outputs(1562)) and (layer2_outputs(281));
    outputs(293) <= layer2_outputs(1807);
    outputs(294) <= not(layer2_outputs(1472));
    outputs(295) <= (layer2_outputs(929)) and (layer2_outputs(103));
    outputs(296) <= not(layer2_outputs(741));
    outputs(297) <= not(layer2_outputs(274));
    outputs(298) <= layer2_outputs(792);
    outputs(299) <= layer2_outputs(1441);
    outputs(300) <= layer2_outputs(2474);
    outputs(301) <= layer2_outputs(874);
    outputs(302) <= layer2_outputs(1078);
    outputs(303) <= layer2_outputs(921);
    outputs(304) <= not((layer2_outputs(580)) and (layer2_outputs(390)));
    outputs(305) <= not(layer2_outputs(1746));
    outputs(306) <= not(layer2_outputs(78));
    outputs(307) <= not((layer2_outputs(997)) xor (layer2_outputs(118)));
    outputs(308) <= not((layer2_outputs(1677)) xor (layer2_outputs(1731)));
    outputs(309) <= layer2_outputs(2236);
    outputs(310) <= not(layer2_outputs(1194));
    outputs(311) <= not(layer2_outputs(2258));
    outputs(312) <= not(layer2_outputs(2091));
    outputs(313) <= (layer2_outputs(2355)) and (layer2_outputs(1754));
    outputs(314) <= not((layer2_outputs(265)) or (layer2_outputs(1629)));
    outputs(315) <= layer2_outputs(1411);
    outputs(316) <= not(layer2_outputs(1688));
    outputs(317) <= layer2_outputs(489);
    outputs(318) <= not((layer2_outputs(385)) or (layer2_outputs(814)));
    outputs(319) <= layer2_outputs(963);
    outputs(320) <= (layer2_outputs(1991)) and not (layer2_outputs(1477));
    outputs(321) <= not(layer2_outputs(1486));
    outputs(322) <= not((layer2_outputs(1906)) xor (layer2_outputs(486)));
    outputs(323) <= layer2_outputs(1214);
    outputs(324) <= not((layer2_outputs(2028)) or (layer2_outputs(753)));
    outputs(325) <= (layer2_outputs(1253)) and not (layer2_outputs(648));
    outputs(326) <= (layer2_outputs(716)) and not (layer2_outputs(852));
    outputs(327) <= not(layer2_outputs(461));
    outputs(328) <= (layer2_outputs(573)) and (layer2_outputs(2011));
    outputs(329) <= not(layer2_outputs(1738));
    outputs(330) <= not(layer2_outputs(906)) or (layer2_outputs(1212));
    outputs(331) <= (layer2_outputs(2088)) and not (layer2_outputs(39));
    outputs(332) <= layer2_outputs(276);
    outputs(333) <= not(layer2_outputs(960));
    outputs(334) <= not((layer2_outputs(32)) or (layer2_outputs(2459)));
    outputs(335) <= not(layer2_outputs(1518));
    outputs(336) <= (layer2_outputs(1379)) and (layer2_outputs(209));
    outputs(337) <= not((layer2_outputs(1681)) or (layer2_outputs(1145)));
    outputs(338) <= not((layer2_outputs(344)) and (layer2_outputs(387)));
    outputs(339) <= not((layer2_outputs(325)) or (layer2_outputs(2342)));
    outputs(340) <= not((layer2_outputs(1513)) xor (layer2_outputs(1903)));
    outputs(341) <= not(layer2_outputs(1644));
    outputs(342) <= not((layer2_outputs(158)) or (layer2_outputs(355)));
    outputs(343) <= (layer2_outputs(2208)) and not (layer2_outputs(1798));
    outputs(344) <= (layer2_outputs(2162)) and (layer2_outputs(1807));
    outputs(345) <= (layer2_outputs(479)) and (layer2_outputs(2330));
    outputs(346) <= (layer2_outputs(1384)) and (layer2_outputs(2501));
    outputs(347) <= (layer2_outputs(885)) xor (layer2_outputs(2340));
    outputs(348) <= (layer2_outputs(1964)) and not (layer2_outputs(296));
    outputs(349) <= not((layer2_outputs(1907)) or (layer2_outputs(633)));
    outputs(350) <= not((layer2_outputs(113)) or (layer2_outputs(1319)));
    outputs(351) <= not((layer2_outputs(1250)) xor (layer2_outputs(241)));
    outputs(352) <= (layer2_outputs(352)) and not (layer2_outputs(475));
    outputs(353) <= (layer2_outputs(1422)) and (layer2_outputs(632));
    outputs(354) <= layer2_outputs(147);
    outputs(355) <= (layer2_outputs(1553)) and not (layer2_outputs(1458));
    outputs(356) <= layer2_outputs(578);
    outputs(357) <= not((layer2_outputs(1320)) or (layer2_outputs(1302)));
    outputs(358) <= not((layer2_outputs(260)) or (layer2_outputs(1925)));
    outputs(359) <= not((layer2_outputs(1022)) or (layer2_outputs(376)));
    outputs(360) <= not((layer2_outputs(1771)) or (layer2_outputs(1862)));
    outputs(361) <= (layer2_outputs(297)) and (layer2_outputs(763));
    outputs(362) <= not((layer2_outputs(2413)) or (layer2_outputs(2324)));
    outputs(363) <= layer2_outputs(550);
    outputs(364) <= not(layer2_outputs(1024));
    outputs(365) <= not((layer2_outputs(26)) or (layer2_outputs(1264)));
    outputs(366) <= not(layer2_outputs(1713));
    outputs(367) <= (layer2_outputs(1857)) and not (layer2_outputs(2024));
    outputs(368) <= not(layer2_outputs(2221));
    outputs(369) <= (layer2_outputs(783)) and not (layer2_outputs(2338));
    outputs(370) <= not(layer2_outputs(131));
    outputs(371) <= (layer2_outputs(1239)) and not (layer2_outputs(2006));
    outputs(372) <= layer2_outputs(514);
    outputs(373) <= layer2_outputs(1042);
    outputs(374) <= layer2_outputs(297);
    outputs(375) <= not(layer2_outputs(274));
    outputs(376) <= (layer2_outputs(2078)) and (layer2_outputs(1577));
    outputs(377) <= (layer2_outputs(135)) and not (layer2_outputs(1624));
    outputs(378) <= not(layer2_outputs(1233));
    outputs(379) <= not((layer2_outputs(131)) or (layer2_outputs(466)));
    outputs(380) <= layer2_outputs(907);
    outputs(381) <= (layer2_outputs(1337)) and not (layer2_outputs(681));
    outputs(382) <= (layer2_outputs(993)) and not (layer2_outputs(26));
    outputs(383) <= (layer2_outputs(348)) and not (layer2_outputs(1222));
    outputs(384) <= (layer2_outputs(35)) and not (layer2_outputs(988));
    outputs(385) <= not((layer2_outputs(1683)) xor (layer2_outputs(1385)));
    outputs(386) <= (layer2_outputs(233)) and (layer2_outputs(1283));
    outputs(387) <= not(layer2_outputs(811));
    outputs(388) <= (layer2_outputs(600)) and not (layer2_outputs(2195));
    outputs(389) <= layer2_outputs(1369);
    outputs(390) <= not(layer2_outputs(277));
    outputs(391) <= layer2_outputs(375);
    outputs(392) <= layer2_outputs(745);
    outputs(393) <= layer2_outputs(130);
    outputs(394) <= layer2_outputs(2353);
    outputs(395) <= not(layer2_outputs(1607));
    outputs(396) <= not((layer2_outputs(1355)) or (layer2_outputs(2299)));
    outputs(397) <= not(layer2_outputs(1377)) or (layer2_outputs(8));
    outputs(398) <= (layer2_outputs(2268)) and not (layer2_outputs(1887));
    outputs(399) <= (layer2_outputs(2517)) and not (layer2_outputs(2211));
    outputs(400) <= layer2_outputs(2389);
    outputs(401) <= (layer2_outputs(562)) and not (layer2_outputs(959));
    outputs(402) <= (layer2_outputs(1499)) and not (layer2_outputs(96));
    outputs(403) <= not(layer2_outputs(2117));
    outputs(404) <= layer2_outputs(2489);
    outputs(405) <= (layer2_outputs(1826)) xor (layer2_outputs(2424));
    outputs(406) <= not(layer2_outputs(1848));
    outputs(407) <= layer2_outputs(2187);
    outputs(408) <= layer2_outputs(765);
    outputs(409) <= not(layer2_outputs(1150));
    outputs(410) <= not((layer2_outputs(569)) or (layer2_outputs(1051)));
    outputs(411) <= (layer2_outputs(2156)) and not (layer2_outputs(2161));
    outputs(412) <= not(layer2_outputs(1561));
    outputs(413) <= layer2_outputs(1228);
    outputs(414) <= layer2_outputs(2419);
    outputs(415) <= (layer2_outputs(111)) and not (layer2_outputs(2135));
    outputs(416) <= not(layer2_outputs(463));
    outputs(417) <= layer2_outputs(723);
    outputs(418) <= (layer2_outputs(643)) and not (layer2_outputs(1550));
    outputs(419) <= (layer2_outputs(258)) and (layer2_outputs(119));
    outputs(420) <= not(layer2_outputs(1156));
    outputs(421) <= (layer2_outputs(2501)) and not (layer2_outputs(2547));
    outputs(422) <= (layer2_outputs(1747)) and not (layer2_outputs(1263));
    outputs(423) <= not(layer2_outputs(2380));
    outputs(424) <= not((layer2_outputs(1665)) or (layer2_outputs(1458)));
    outputs(425) <= not(layer2_outputs(1016));
    outputs(426) <= (layer2_outputs(1201)) and not (layer2_outputs(25));
    outputs(427) <= not(layer2_outputs(931));
    outputs(428) <= not((layer2_outputs(694)) or (layer2_outputs(2420)));
    outputs(429) <= layer2_outputs(1341);
    outputs(430) <= not((layer2_outputs(1116)) xor (layer2_outputs(684)));
    outputs(431) <= not((layer2_outputs(1843)) or (layer2_outputs(469)));
    outputs(432) <= not(layer2_outputs(2420));
    outputs(433) <= layer2_outputs(2129);
    outputs(434) <= not((layer2_outputs(1403)) or (layer2_outputs(1901)));
    outputs(435) <= not(layer2_outputs(1511));
    outputs(436) <= (layer2_outputs(1811)) and (layer2_outputs(31));
    outputs(437) <= not(layer2_outputs(893));
    outputs(438) <= (layer2_outputs(2067)) and not (layer2_outputs(901));
    outputs(439) <= (layer2_outputs(1199)) and not (layer2_outputs(2543));
    outputs(440) <= not(layer2_outputs(2122));
    outputs(441) <= (layer2_outputs(2445)) xor (layer2_outputs(2334));
    outputs(442) <= not(layer2_outputs(1418));
    outputs(443) <= layer2_outputs(1627);
    outputs(444) <= not((layer2_outputs(1668)) or (layer2_outputs(1507)));
    outputs(445) <= not(layer2_outputs(193));
    outputs(446) <= layer2_outputs(166);
    outputs(447) <= (layer2_outputs(918)) and not (layer2_outputs(705));
    outputs(448) <= not((layer2_outputs(1272)) xor (layer2_outputs(1740)));
    outputs(449) <= not((layer2_outputs(677)) or (layer2_outputs(804)));
    outputs(450) <= (layer2_outputs(71)) and not (layer2_outputs(650));
    outputs(451) <= layer2_outputs(1040);
    outputs(452) <= layer2_outputs(428);
    outputs(453) <= not((layer2_outputs(450)) or (layer2_outputs(2298)));
    outputs(454) <= (layer2_outputs(2531)) and (layer2_outputs(1754));
    outputs(455) <= (layer2_outputs(877)) and (layer2_outputs(1535));
    outputs(456) <= not((layer2_outputs(81)) or (layer2_outputs(960)));
    outputs(457) <= (layer2_outputs(572)) and not (layer2_outputs(1713));
    outputs(458) <= not((layer2_outputs(716)) xor (layer2_outputs(132)));
    outputs(459) <= layer2_outputs(1370);
    outputs(460) <= layer2_outputs(925);
    outputs(461) <= (layer2_outputs(1240)) xor (layer2_outputs(2396));
    outputs(462) <= (layer2_outputs(59)) and not (layer2_outputs(2403));
    outputs(463) <= (layer2_outputs(697)) and (layer2_outputs(854));
    outputs(464) <= layer2_outputs(1287);
    outputs(465) <= not(layer2_outputs(1234));
    outputs(466) <= layer2_outputs(1856);
    outputs(467) <= (layer2_outputs(216)) and (layer2_outputs(2319));
    outputs(468) <= (layer2_outputs(992)) xor (layer2_outputs(1566));
    outputs(469) <= not(layer2_outputs(370));
    outputs(470) <= (layer2_outputs(493)) and not (layer2_outputs(1584));
    outputs(471) <= (layer2_outputs(2480)) and not (layer2_outputs(2047));
    outputs(472) <= not((layer2_outputs(357)) or (layer2_outputs(1355)));
    outputs(473) <= layer2_outputs(672);
    outputs(474) <= not(layer2_outputs(2258));
    outputs(475) <= (layer2_outputs(561)) and not (layer2_outputs(804));
    outputs(476) <= not(layer2_outputs(996));
    outputs(477) <= layer2_outputs(154);
    outputs(478) <= not((layer2_outputs(199)) or (layer2_outputs(1877)));
    outputs(479) <= layer2_outputs(2019);
    outputs(480) <= layer2_outputs(1048);
    outputs(481) <= (layer2_outputs(383)) and not (layer2_outputs(769));
    outputs(482) <= (layer2_outputs(2183)) and (layer2_outputs(271));
    outputs(483) <= not((layer2_outputs(2031)) xor (layer2_outputs(470)));
    outputs(484) <= (layer2_outputs(526)) and not (layer2_outputs(1329));
    outputs(485) <= not(layer2_outputs(138));
    outputs(486) <= (layer2_outputs(2319)) and not (layer2_outputs(581));
    outputs(487) <= (layer2_outputs(1655)) and (layer2_outputs(218));
    outputs(488) <= layer2_outputs(2438);
    outputs(489) <= (layer2_outputs(706)) xor (layer2_outputs(645));
    outputs(490) <= not(layer2_outputs(2188));
    outputs(491) <= (layer2_outputs(479)) and not (layer2_outputs(1738));
    outputs(492) <= (layer2_outputs(1346)) and not (layer2_outputs(1410));
    outputs(493) <= (layer2_outputs(1962)) and (layer2_outputs(2171));
    outputs(494) <= not(layer2_outputs(519));
    outputs(495) <= not((layer2_outputs(51)) or (layer2_outputs(228)));
    outputs(496) <= not(layer2_outputs(1726));
    outputs(497) <= layer2_outputs(1591);
    outputs(498) <= (layer2_outputs(816)) and (layer2_outputs(224));
    outputs(499) <= (layer2_outputs(1293)) and (layer2_outputs(1457));
    outputs(500) <= layer2_outputs(818);
    outputs(501) <= (layer2_outputs(966)) and not (layer2_outputs(1308));
    outputs(502) <= (layer2_outputs(421)) and (layer2_outputs(1593));
    outputs(503) <= (layer2_outputs(89)) and not (layer2_outputs(1226));
    outputs(504) <= layer2_outputs(1869);
    outputs(505) <= layer2_outputs(803);
    outputs(506) <= not(layer2_outputs(965));
    outputs(507) <= layer2_outputs(2332);
    outputs(508) <= not(layer2_outputs(1487));
    outputs(509) <= layer2_outputs(1892);
    outputs(510) <= (layer2_outputs(1026)) and not (layer2_outputs(1570));
    outputs(511) <= layer2_outputs(29);
    outputs(512) <= not((layer2_outputs(1752)) xor (layer2_outputs(196)));
    outputs(513) <= layer2_outputs(210);
    outputs(514) <= layer2_outputs(375);
    outputs(515) <= not(layer2_outputs(2467));
    outputs(516) <= not(layer2_outputs(790));
    outputs(517) <= (layer2_outputs(1461)) and not (layer2_outputs(1484));
    outputs(518) <= layer2_outputs(1952);
    outputs(519) <= not(layer2_outputs(213));
    outputs(520) <= layer2_outputs(1280);
    outputs(521) <= not(layer2_outputs(616));
    outputs(522) <= layer2_outputs(1049);
    outputs(523) <= not(layer2_outputs(1587)) or (layer2_outputs(1459));
    outputs(524) <= not(layer2_outputs(2331));
    outputs(525) <= layer2_outputs(570);
    outputs(526) <= (layer2_outputs(362)) and (layer2_outputs(1676));
    outputs(527) <= (layer2_outputs(1364)) xor (layer2_outputs(1051));
    outputs(528) <= layer2_outputs(187);
    outputs(529) <= not((layer2_outputs(2455)) or (layer2_outputs(2559)));
    outputs(530) <= (layer2_outputs(419)) xor (layer2_outputs(1028));
    outputs(531) <= layer2_outputs(2262);
    outputs(532) <= not(layer2_outputs(1249));
    outputs(533) <= not((layer2_outputs(2153)) or (layer2_outputs(871)));
    outputs(534) <= layer2_outputs(1801);
    outputs(535) <= (layer2_outputs(2218)) or (layer2_outputs(873));
    outputs(536) <= not((layer2_outputs(2016)) and (layer2_outputs(2351)));
    outputs(537) <= (layer2_outputs(254)) and not (layer2_outputs(2030));
    outputs(538) <= not(layer2_outputs(2273));
    outputs(539) <= layer2_outputs(1124);
    outputs(540) <= not((layer2_outputs(1617)) xor (layer2_outputs(1870)));
    outputs(541) <= not(layer2_outputs(2072));
    outputs(542) <= (layer2_outputs(212)) xor (layer2_outputs(1896));
    outputs(543) <= layer2_outputs(916);
    outputs(544) <= not((layer2_outputs(306)) or (layer2_outputs(2260)));
    outputs(545) <= (layer2_outputs(1702)) xor (layer2_outputs(1133));
    outputs(546) <= (layer2_outputs(1819)) and (layer2_outputs(1804));
    outputs(547) <= layer2_outputs(1979);
    outputs(548) <= not(layer2_outputs(1808));
    outputs(549) <= (layer2_outputs(47)) or (layer2_outputs(1855));
    outputs(550) <= not((layer2_outputs(1868)) or (layer2_outputs(2040)));
    outputs(551) <= not((layer2_outputs(2033)) xor (layer2_outputs(1540)));
    outputs(552) <= not(layer2_outputs(1546));
    outputs(553) <= layer2_outputs(2412);
    outputs(554) <= layer2_outputs(527);
    outputs(555) <= not((layer2_outputs(219)) xor (layer2_outputs(2432)));
    outputs(556) <= not((layer2_outputs(1985)) xor (layer2_outputs(1983)));
    outputs(557) <= layer2_outputs(2317);
    outputs(558) <= not((layer2_outputs(2019)) or (layer2_outputs(1638)));
    outputs(559) <= not(layer2_outputs(1632));
    outputs(560) <= layer2_outputs(855);
    outputs(561) <= (layer2_outputs(1954)) and (layer2_outputs(1060));
    outputs(562) <= (layer2_outputs(2402)) and (layer2_outputs(682));
    outputs(563) <= layer2_outputs(2215);
    outputs(564) <= (layer2_outputs(1300)) and not (layer2_outputs(28));
    outputs(565) <= layer2_outputs(1667);
    outputs(566) <= layer2_outputs(1534);
    outputs(567) <= (layer2_outputs(2194)) and not (layer2_outputs(1968));
    outputs(568) <= layer2_outputs(589);
    outputs(569) <= layer2_outputs(235);
    outputs(570) <= layer2_outputs(1251);
    outputs(571) <= not(layer2_outputs(1770)) or (layer2_outputs(382));
    outputs(572) <= not(layer2_outputs(1210));
    outputs(573) <= not(layer2_outputs(165));
    outputs(574) <= not(layer2_outputs(1386));
    outputs(575) <= (layer2_outputs(1084)) and not (layer2_outputs(2290));
    outputs(576) <= layer2_outputs(1721);
    outputs(577) <= layer2_outputs(2272);
    outputs(578) <= not(layer2_outputs(2238));
    outputs(579) <= layer2_outputs(1871);
    outputs(580) <= layer2_outputs(686);
    outputs(581) <= (layer2_outputs(1684)) and not (layer2_outputs(2314));
    outputs(582) <= (layer2_outputs(785)) and (layer2_outputs(230));
    outputs(583) <= (layer2_outputs(491)) and not (layer2_outputs(1640));
    outputs(584) <= (layer2_outputs(449)) and (layer2_outputs(1206));
    outputs(585) <= layer2_outputs(1504);
    outputs(586) <= not(layer2_outputs(1785));
    outputs(587) <= not(layer2_outputs(551));
    outputs(588) <= layer2_outputs(1537);
    outputs(589) <= (layer2_outputs(1152)) or (layer2_outputs(663));
    outputs(590) <= (layer2_outputs(1236)) and not (layer2_outputs(1978));
    outputs(591) <= not((layer2_outputs(1165)) and (layer2_outputs(2007)));
    outputs(592) <= not(layer2_outputs(1448));
    outputs(593) <= layer2_outputs(46);
    outputs(594) <= layer2_outputs(468);
    outputs(595) <= not(layer2_outputs(498));
    outputs(596) <= layer2_outputs(406);
    outputs(597) <= not(layer2_outputs(69));
    outputs(598) <= not(layer2_outputs(1273));
    outputs(599) <= not(layer2_outputs(1745));
    outputs(600) <= layer2_outputs(2267);
    outputs(601) <= (layer2_outputs(1310)) xor (layer2_outputs(1609));
    outputs(602) <= layer2_outputs(821);
    outputs(603) <= not(layer2_outputs(2520));
    outputs(604) <= (layer2_outputs(1589)) and not (layer2_outputs(877));
    outputs(605) <= not((layer2_outputs(1441)) xor (layer2_outputs(2127)));
    outputs(606) <= (layer2_outputs(2459)) and (layer2_outputs(1072));
    outputs(607) <= layer2_outputs(1673);
    outputs(608) <= not(layer2_outputs(668));
    outputs(609) <= layer2_outputs(1958);
    outputs(610) <= (layer2_outputs(47)) and (layer2_outputs(1254));
    outputs(611) <= not(layer2_outputs(384));
    outputs(612) <= layer2_outputs(1584);
    outputs(613) <= not(layer2_outputs(631));
    outputs(614) <= not((layer2_outputs(1332)) or (layer2_outputs(1212)));
    outputs(615) <= not(layer2_outputs(33));
    outputs(616) <= layer2_outputs(366);
    outputs(617) <= layer2_outputs(2297);
    outputs(618) <= not(layer2_outputs(1919));
    outputs(619) <= layer2_outputs(1164);
    outputs(620) <= layer2_outputs(904);
    outputs(621) <= (layer2_outputs(137)) xor (layer2_outputs(2208));
    outputs(622) <= (layer2_outputs(1622)) or (layer2_outputs(2541));
    outputs(623) <= (layer2_outputs(109)) and not (layer2_outputs(2350));
    outputs(624) <= layer2_outputs(531);
    outputs(625) <= (layer2_outputs(1514)) and not (layer2_outputs(1193));
    outputs(626) <= (layer2_outputs(1314)) and (layer2_outputs(254));
    outputs(627) <= not(layer2_outputs(1728));
    outputs(628) <= layer2_outputs(1460);
    outputs(629) <= layer2_outputs(2241);
    outputs(630) <= not(layer2_outputs(1811));
    outputs(631) <= layer2_outputs(1939);
    outputs(632) <= layer2_outputs(13);
    outputs(633) <= layer2_outputs(1529);
    outputs(634) <= not(layer2_outputs(213));
    outputs(635) <= not(layer2_outputs(142));
    outputs(636) <= not(layer2_outputs(171));
    outputs(637) <= (layer2_outputs(844)) and not (layer2_outputs(506));
    outputs(638) <= not(layer2_outputs(1586));
    outputs(639) <= not(layer2_outputs(971));
    outputs(640) <= (layer2_outputs(658)) and not (layer2_outputs(1869));
    outputs(641) <= (layer2_outputs(979)) and (layer2_outputs(455));
    outputs(642) <= layer2_outputs(65);
    outputs(643) <= layer2_outputs(604);
    outputs(644) <= not(layer2_outputs(2535));
    outputs(645) <= layer2_outputs(1737);
    outputs(646) <= not(layer2_outputs(2148));
    outputs(647) <= not(layer2_outputs(173));
    outputs(648) <= layer2_outputs(2449);
    outputs(649) <= layer2_outputs(515);
    outputs(650) <= not(layer2_outputs(361));
    outputs(651) <= not(layer2_outputs(2534));
    outputs(652) <= layer2_outputs(259);
    outputs(653) <= not(layer2_outputs(548));
    outputs(654) <= layer2_outputs(911);
    outputs(655) <= not((layer2_outputs(1701)) or (layer2_outputs(2372)));
    outputs(656) <= layer2_outputs(648);
    outputs(657) <= not(layer2_outputs(1938));
    outputs(658) <= not(layer2_outputs(1691));
    outputs(659) <= layer2_outputs(1641);
    outputs(660) <= layer2_outputs(1246);
    outputs(661) <= not(layer2_outputs(685));
    outputs(662) <= (layer2_outputs(2410)) and (layer2_outputs(1756));
    outputs(663) <= not(layer2_outputs(2400));
    outputs(664) <= (layer2_outputs(492)) and not (layer2_outputs(1474));
    outputs(665) <= not((layer2_outputs(1696)) or (layer2_outputs(237)));
    outputs(666) <= layer2_outputs(203);
    outputs(667) <= layer2_outputs(1312);
    outputs(668) <= not(layer2_outputs(1881));
    outputs(669) <= not(layer2_outputs(2029));
    outputs(670) <= not(layer2_outputs(2524)) or (layer2_outputs(1550));
    outputs(671) <= layer2_outputs(933);
    outputs(672) <= not((layer2_outputs(2237)) and (layer2_outputs(2079)));
    outputs(673) <= (layer2_outputs(2479)) and not (layer2_outputs(342));
    outputs(674) <= (layer2_outputs(1981)) and (layer2_outputs(1851));
    outputs(675) <= not(layer2_outputs(1883));
    outputs(676) <= not(layer2_outputs(613));
    outputs(677) <= layer2_outputs(2291);
    outputs(678) <= (layer2_outputs(1673)) and not (layer2_outputs(456));
    outputs(679) <= layer2_outputs(679);
    outputs(680) <= layer2_outputs(904);
    outputs(681) <= layer2_outputs(1110);
    outputs(682) <= layer2_outputs(1969);
    outputs(683) <= layer2_outputs(2366);
    outputs(684) <= not(layer2_outputs(308));
    outputs(685) <= not(layer2_outputs(1363));
    outputs(686) <= layer2_outputs(1190);
    outputs(687) <= not(layer2_outputs(1343)) or (layer2_outputs(2556));
    outputs(688) <= not(layer2_outputs(850));
    outputs(689) <= (layer2_outputs(234)) and not (layer2_outputs(972));
    outputs(690) <= not(layer2_outputs(538));
    outputs(691) <= layer2_outputs(1499);
    outputs(692) <= layer2_outputs(711);
    outputs(693) <= (layer2_outputs(497)) and (layer2_outputs(1121));
    outputs(694) <= layer2_outputs(683);
    outputs(695) <= not(layer2_outputs(1000));
    outputs(696) <= not((layer2_outputs(765)) or (layer2_outputs(1595)));
    outputs(697) <= not(layer2_outputs(361));
    outputs(698) <= not(layer2_outputs(1160));
    outputs(699) <= (layer2_outputs(2164)) xor (layer2_outputs(1750));
    outputs(700) <= not(layer2_outputs(2341));
    outputs(701) <= not(layer2_outputs(704));
    outputs(702) <= layer2_outputs(2284);
    outputs(703) <= (layer2_outputs(1149)) xor (layer2_outputs(195));
    outputs(704) <= layer2_outputs(2361);
    outputs(705) <= not(layer2_outputs(1333));
    outputs(706) <= layer2_outputs(671);
    outputs(707) <= layer2_outputs(2297);
    outputs(708) <= layer2_outputs(1542);
    outputs(709) <= not(layer2_outputs(758));
    outputs(710) <= layer2_outputs(928);
    outputs(711) <= (layer2_outputs(744)) xor (layer2_outputs(2011));
    outputs(712) <= (layer2_outputs(1447)) and (layer2_outputs(1082));
    outputs(713) <= layer2_outputs(2371);
    outputs(714) <= (layer2_outputs(825)) and not (layer2_outputs(737));
    outputs(715) <= not((layer2_outputs(945)) or (layer2_outputs(899)));
    outputs(716) <= not(layer2_outputs(666));
    outputs(717) <= (layer2_outputs(1488)) and not (layer2_outputs(27));
    outputs(718) <= not(layer2_outputs(1701));
    outputs(719) <= layer2_outputs(85);
    outputs(720) <= layer2_outputs(1556);
    outputs(721) <= not(layer2_outputs(303)) or (layer2_outputs(602));
    outputs(722) <= layer2_outputs(1318);
    outputs(723) <= (layer2_outputs(849)) and (layer2_outputs(1512));
    outputs(724) <= not(layer2_outputs(512));
    outputs(725) <= (layer2_outputs(2098)) and not (layer2_outputs(1100));
    outputs(726) <= not(layer2_outputs(69));
    outputs(727) <= not(layer2_outputs(1017));
    outputs(728) <= (layer2_outputs(1126)) and not (layer2_outputs(371));
    outputs(729) <= not(layer2_outputs(1553));
    outputs(730) <= not(layer2_outputs(1883));
    outputs(731) <= layer2_outputs(694);
    outputs(732) <= (layer2_outputs(2399)) and not (layer2_outputs(1073));
    outputs(733) <= layer2_outputs(168);
    outputs(734) <= not((layer2_outputs(639)) xor (layer2_outputs(1373)));
    outputs(735) <= not(layer2_outputs(2379));
    outputs(736) <= (layer2_outputs(2046)) and not (layer2_outputs(2531));
    outputs(737) <= (layer2_outputs(1002)) and not (layer2_outputs(1059));
    outputs(738) <= not(layer2_outputs(1105));
    outputs(739) <= not(layer2_outputs(99));
    outputs(740) <= layer2_outputs(1382);
    outputs(741) <= not(layer2_outputs(771));
    outputs(742) <= layer2_outputs(1917);
    outputs(743) <= not((layer2_outputs(2521)) and (layer2_outputs(923)));
    outputs(744) <= (layer2_outputs(823)) xor (layer2_outputs(2430));
    outputs(745) <= layer2_outputs(1756);
    outputs(746) <= not(layer2_outputs(2480));
    outputs(747) <= (layer2_outputs(155)) or (layer2_outputs(261));
    outputs(748) <= (layer2_outputs(2144)) xor (layer2_outputs(808));
    outputs(749) <= (layer2_outputs(2263)) and (layer2_outputs(1557));
    outputs(750) <= layer2_outputs(1845);
    outputs(751) <= layer2_outputs(1038);
    outputs(752) <= not(layer2_outputs(1967));
    outputs(753) <= not(layer2_outputs(2300));
    outputs(754) <= layer2_outputs(1497);
    outputs(755) <= (layer2_outputs(1537)) xor (layer2_outputs(1744));
    outputs(756) <= not(layer2_outputs(80));
    outputs(757) <= not(layer2_outputs(1354));
    outputs(758) <= not(layer2_outputs(1050));
    outputs(759) <= not((layer2_outputs(813)) xor (layer2_outputs(248)));
    outputs(760) <= layer2_outputs(1776);
    outputs(761) <= (layer2_outputs(1493)) and not (layer2_outputs(938));
    outputs(762) <= not(layer2_outputs(1781));
    outputs(763) <= (layer2_outputs(1906)) or (layer2_outputs(1231));
    outputs(764) <= (layer2_outputs(1758)) and (layer2_outputs(803));
    outputs(765) <= not(layer2_outputs(866));
    outputs(766) <= (layer2_outputs(2103)) and (layer2_outputs(420));
    outputs(767) <= (layer2_outputs(1140)) and not (layer2_outputs(199));
    outputs(768) <= not((layer2_outputs(1824)) xor (layer2_outputs(76)));
    outputs(769) <= layer2_outputs(2052);
    outputs(770) <= (layer2_outputs(760)) and not (layer2_outputs(752));
    outputs(771) <= not(layer2_outputs(1774));
    outputs(772) <= (layer2_outputs(432)) and (layer2_outputs(1408));
    outputs(773) <= not(layer2_outputs(177));
    outputs(774) <= layer2_outputs(2192);
    outputs(775) <= layer2_outputs(56);
    outputs(776) <= layer2_outputs(1466);
    outputs(777) <= not((layer2_outputs(1918)) or (layer2_outputs(1392)));
    outputs(778) <= not(layer2_outputs(183));
    outputs(779) <= (layer2_outputs(1824)) and not (layer2_outputs(2190));
    outputs(780) <= layer2_outputs(2439);
    outputs(781) <= layer2_outputs(1350);
    outputs(782) <= not(layer2_outputs(1223));
    outputs(783) <= not(layer2_outputs(140));
    outputs(784) <= (layer2_outputs(1106)) and not (layer2_outputs(1725));
    outputs(785) <= not(layer2_outputs(661));
    outputs(786) <= not(layer2_outputs(1020));
    outputs(787) <= layer2_outputs(1350);
    outputs(788) <= not((layer2_outputs(2115)) xor (layer2_outputs(2401)));
    outputs(789) <= layer2_outputs(160);
    outputs(790) <= not(layer2_outputs(2524)) or (layer2_outputs(2182));
    outputs(791) <= not(layer2_outputs(1465));
    outputs(792) <= (layer2_outputs(1992)) and not (layer2_outputs(38));
    outputs(793) <= layer2_outputs(2411);
    outputs(794) <= (layer2_outputs(1343)) or (layer2_outputs(2435));
    outputs(795) <= not((layer2_outputs(1348)) xor (layer2_outputs(248)));
    outputs(796) <= not(layer2_outputs(44));
    outputs(797) <= layer2_outputs(907);
    outputs(798) <= not(layer2_outputs(906));
    outputs(799) <= not(layer2_outputs(764));
    outputs(800) <= not(layer2_outputs(1787));
    outputs(801) <= not((layer2_outputs(15)) or (layer2_outputs(1510)));
    outputs(802) <= (layer2_outputs(357)) and (layer2_outputs(487));
    outputs(803) <= not(layer2_outputs(598));
    outputs(804) <= not(layer2_outputs(2552));
    outputs(805) <= not(layer2_outputs(1250));
    outputs(806) <= not(layer2_outputs(1211));
    outputs(807) <= layer2_outputs(1963);
    outputs(808) <= not(layer2_outputs(336));
    outputs(809) <= (layer2_outputs(689)) xor (layer2_outputs(1758));
    outputs(810) <= (layer2_outputs(1257)) and (layer2_outputs(1705));
    outputs(811) <= (layer2_outputs(2334)) or (layer2_outputs(643));
    outputs(812) <= not(layer2_outputs(817));
    outputs(813) <= not((layer2_outputs(1129)) or (layer2_outputs(1394)));
    outputs(814) <= (layer2_outputs(418)) and not (layer2_outputs(961));
    outputs(815) <= (layer2_outputs(2353)) and not (layer2_outputs(2207));
    outputs(816) <= (layer2_outputs(2471)) and (layer2_outputs(971));
    outputs(817) <= (layer2_outputs(939)) and (layer2_outputs(1069));
    outputs(818) <= (layer2_outputs(1859)) and not (layer2_outputs(1984));
    outputs(819) <= not((layer2_outputs(2495)) or (layer2_outputs(2018)));
    outputs(820) <= layer2_outputs(709);
    outputs(821) <= layer2_outputs(167);
    outputs(822) <= (layer2_outputs(1564)) and not (layer2_outputs(2444));
    outputs(823) <= layer2_outputs(2345);
    outputs(824) <= not(layer2_outputs(757)) or (layer2_outputs(797));
    outputs(825) <= (layer2_outputs(1662)) and not (layer2_outputs(1142));
    outputs(826) <= not((layer2_outputs(936)) or (layer2_outputs(1725)));
    outputs(827) <= not(layer2_outputs(2511));
    outputs(828) <= not(layer2_outputs(1425));
    outputs(829) <= layer2_outputs(777);
    outputs(830) <= (layer2_outputs(4)) and not (layer2_outputs(823));
    outputs(831) <= not(layer2_outputs(559));
    outputs(832) <= layer2_outputs(1323);
    outputs(833) <= not(layer2_outputs(933));
    outputs(834) <= not(layer2_outputs(2551));
    outputs(835) <= layer2_outputs(2081);
    outputs(836) <= (layer2_outputs(1880)) and not (layer2_outputs(698));
    outputs(837) <= (layer2_outputs(2219)) xor (layer2_outputs(2378));
    outputs(838) <= layer2_outputs(2198);
    outputs(839) <= not((layer2_outputs(295)) xor (layer2_outputs(1087)));
    outputs(840) <= not(layer2_outputs(1129)) or (layer2_outputs(967));
    outputs(841) <= not(layer2_outputs(46));
    outputs(842) <= not(layer2_outputs(1276));
    outputs(843) <= not((layer2_outputs(1494)) or (layer2_outputs(307)));
    outputs(844) <= layer2_outputs(11);
    outputs(845) <= not((layer2_outputs(1244)) xor (layer2_outputs(1164)));
    outputs(846) <= (layer2_outputs(1047)) xor (layer2_outputs(106));
    outputs(847) <= layer2_outputs(90);
    outputs(848) <= layer2_outputs(2549);
    outputs(849) <= (layer2_outputs(1642)) and not (layer2_outputs(2219));
    outputs(850) <= not(layer2_outputs(168));
    outputs(851) <= not(layer2_outputs(1563));
    outputs(852) <= layer2_outputs(761);
    outputs(853) <= not(layer2_outputs(100));
    outputs(854) <= not(layer2_outputs(1974));
    outputs(855) <= not((layer2_outputs(2176)) or (layer2_outputs(702)));
    outputs(856) <= not(layer2_outputs(2017));
    outputs(857) <= layer2_outputs(1131);
    outputs(858) <= layer2_outputs(134);
    outputs(859) <= (layer2_outputs(1378)) and not (layer2_outputs(1861));
    outputs(860) <= (layer2_outputs(964)) and not (layer2_outputs(124));
    outputs(861) <= not(layer2_outputs(1696));
    outputs(862) <= not(layer2_outputs(2342));
    outputs(863) <= not(layer2_outputs(1186));
    outputs(864) <= not(layer2_outputs(225));
    outputs(865) <= not(layer2_outputs(437));
    outputs(866) <= not((layer2_outputs(1516)) xor (layer2_outputs(822)));
    outputs(867) <= layer2_outputs(722);
    outputs(868) <= layer2_outputs(809);
    outputs(869) <= (layer2_outputs(2548)) and not (layer2_outputs(1033));
    outputs(870) <= layer2_outputs(639);
    outputs(871) <= layer2_outputs(1503);
    outputs(872) <= (layer2_outputs(738)) and not (layer2_outputs(1755));
    outputs(873) <= (layer2_outputs(1334)) and not (layer2_outputs(2201));
    outputs(874) <= not(layer2_outputs(2370));
    outputs(875) <= not(layer2_outputs(952));
    outputs(876) <= layer2_outputs(2259);
    outputs(877) <= not(layer2_outputs(2003));
    outputs(878) <= not(layer2_outputs(1592)) or (layer2_outputs(672));
    outputs(879) <= layer2_outputs(2110);
    outputs(880) <= not(layer2_outputs(1730));
    outputs(881) <= layer2_outputs(1697);
    outputs(882) <= not((layer2_outputs(263)) or (layer2_outputs(1375)));
    outputs(883) <= layer2_outputs(347);
    outputs(884) <= (layer2_outputs(251)) and not (layer2_outputs(2509));
    outputs(885) <= layer2_outputs(30);
    outputs(886) <= layer2_outputs(1515);
    outputs(887) <= not(layer2_outputs(2370));
    outputs(888) <= not(layer2_outputs(250));
    outputs(889) <= (layer2_outputs(1520)) xor (layer2_outputs(2024));
    outputs(890) <= layer2_outputs(2305);
    outputs(891) <= (layer2_outputs(692)) and not (layer2_outputs(1341));
    outputs(892) <= not((layer2_outputs(1850)) or (layer2_outputs(1401)));
    outputs(893) <= (layer2_outputs(1431)) xor (layer2_outputs(74));
    outputs(894) <= layer2_outputs(557);
    outputs(895) <= layer2_outputs(1951);
    outputs(896) <= not(layer2_outputs(828));
    outputs(897) <= (layer2_outputs(2178)) or (layer2_outputs(443));
    outputs(898) <= not(layer2_outputs(1151));
    outputs(899) <= layer2_outputs(2021);
    outputs(900) <= layer2_outputs(2326);
    outputs(901) <= not(layer2_outputs(617));
    outputs(902) <= not(layer2_outputs(1616));
    outputs(903) <= not((layer2_outputs(609)) or (layer2_outputs(2158)));
    outputs(904) <= not((layer2_outputs(439)) or (layer2_outputs(1294)));
    outputs(905) <= (layer2_outputs(2035)) and (layer2_outputs(1816));
    outputs(906) <= not(layer2_outputs(798));
    outputs(907) <= not(layer2_outputs(2120));
    outputs(908) <= not(layer2_outputs(1840));
    outputs(909) <= not(layer2_outputs(2323));
    outputs(910) <= not((layer2_outputs(312)) or (layer2_outputs(247)));
    outputs(911) <= layer2_outputs(506);
    outputs(912) <= not(layer2_outputs(1902));
    outputs(913) <= not(layer2_outputs(1916));
    outputs(914) <= not(layer2_outputs(1929));
    outputs(915) <= layer2_outputs(2479);
    outputs(916) <= not(layer2_outputs(2360));
    outputs(917) <= layer2_outputs(2166);
    outputs(918) <= (layer2_outputs(1023)) and not (layer2_outputs(1264));
    outputs(919) <= not(layer2_outputs(867));
    outputs(920) <= layer2_outputs(93);
    outputs(921) <= not((layer2_outputs(1962)) and (layer2_outputs(22)));
    outputs(922) <= not((layer2_outputs(253)) or (layer2_outputs(2361)));
    outputs(923) <= (layer2_outputs(1634)) and not (layer2_outputs(1910));
    outputs(924) <= (layer2_outputs(928)) or (layer2_outputs(279));
    outputs(925) <= layer2_outputs(946);
    outputs(926) <= (layer2_outputs(748)) and not (layer2_outputs(1342));
    outputs(927) <= not((layer2_outputs(1704)) xor (layer2_outputs(2307)));
    outputs(928) <= layer2_outputs(315);
    outputs(929) <= not(layer2_outputs(1133));
    outputs(930) <= not(layer2_outputs(2466));
    outputs(931) <= layer2_outputs(232);
    outputs(932) <= (layer2_outputs(1699)) or (layer2_outputs(1878));
    outputs(933) <= not(layer2_outputs(2318));
    outputs(934) <= (layer2_outputs(1989)) or (layer2_outputs(138));
    outputs(935) <= not(layer2_outputs(2358));
    outputs(936) <= not(layer2_outputs(19));
    outputs(937) <= not(layer2_outputs(460)) or (layer2_outputs(1830));
    outputs(938) <= not(layer2_outputs(1961));
    outputs(939) <= not((layer2_outputs(2504)) and (layer2_outputs(1114)));
    outputs(940) <= not((layer2_outputs(1447)) xor (layer2_outputs(853)));
    outputs(941) <= not((layer2_outputs(148)) or (layer2_outputs(1296)));
    outputs(942) <= (layer2_outputs(1370)) or (layer2_outputs(507));
    outputs(943) <= not(layer2_outputs(1298));
    outputs(944) <= layer2_outputs(1106);
    outputs(945) <= layer2_outputs(902);
    outputs(946) <= not(layer2_outputs(1964));
    outputs(947) <= (layer2_outputs(2013)) and (layer2_outputs(1461));
    outputs(948) <= layer2_outputs(2451);
    outputs(949) <= (layer2_outputs(1402)) and (layer2_outputs(1069));
    outputs(950) <= layer2_outputs(1963);
    outputs(951) <= not(layer2_outputs(2006));
    outputs(952) <= layer2_outputs(1518);
    outputs(953) <= not(layer2_outputs(702));
    outputs(954) <= not((layer2_outputs(1560)) or (layer2_outputs(311)));
    outputs(955) <= layer2_outputs(2107);
    outputs(956) <= layer2_outputs(10);
    outputs(957) <= not(layer2_outputs(439));
    outputs(958) <= not(layer2_outputs(707));
    outputs(959) <= not(layer2_outputs(2505));
    outputs(960) <= layer2_outputs(871);
    outputs(961) <= (layer2_outputs(4)) and (layer2_outputs(504));
    outputs(962) <= layer2_outputs(2534);
    outputs(963) <= not(layer2_outputs(1783));
    outputs(964) <= layer2_outputs(1500);
    outputs(965) <= not((layer2_outputs(1589)) and (layer2_outputs(568)));
    outputs(966) <= layer2_outputs(2246);
    outputs(967) <= (layer2_outputs(1599)) and not (layer2_outputs(430));
    outputs(968) <= (layer2_outputs(1739)) and not (layer2_outputs(539));
    outputs(969) <= not((layer2_outputs(381)) or (layer2_outputs(696)));
    outputs(970) <= not((layer2_outputs(1429)) xor (layer2_outputs(2354)));
    outputs(971) <= (layer2_outputs(2464)) xor (layer2_outputs(1015));
    outputs(972) <= (layer2_outputs(704)) and not (layer2_outputs(2257));
    outputs(973) <= not((layer2_outputs(438)) or (layer2_outputs(1111)));
    outputs(974) <= (layer2_outputs(1969)) and (layer2_outputs(376));
    outputs(975) <= layer2_outputs(2546);
    outputs(976) <= not(layer2_outputs(2239));
    outputs(977) <= layer2_outputs(318);
    outputs(978) <= (layer2_outputs(1652)) and (layer2_outputs(498));
    outputs(979) <= layer2_outputs(2320);
    outputs(980) <= not(layer2_outputs(651));
    outputs(981) <= not((layer2_outputs(1762)) or (layer2_outputs(1157)));
    outputs(982) <= (layer2_outputs(2112)) and not (layer2_outputs(2304));
    outputs(983) <= not(layer2_outputs(986));
    outputs(984) <= not(layer2_outputs(169));
    outputs(985) <= (layer2_outputs(2210)) and not (layer2_outputs(1660));
    outputs(986) <= not(layer2_outputs(304));
    outputs(987) <= not(layer2_outputs(1433));
    outputs(988) <= layer2_outputs(2014);
    outputs(989) <= (layer2_outputs(1757)) and not (layer2_outputs(1583));
    outputs(990) <= layer2_outputs(1321);
    outputs(991) <= not(layer2_outputs(1889)) or (layer2_outputs(2490));
    outputs(992) <= layer2_outputs(2256);
    outputs(993) <= layer2_outputs(1884);
    outputs(994) <= layer2_outputs(611);
    outputs(995) <= not((layer2_outputs(1532)) xor (layer2_outputs(85)));
    outputs(996) <= (layer2_outputs(2488)) and not (layer2_outputs(921));
    outputs(997) <= not((layer2_outputs(530)) or (layer2_outputs(429)));
    outputs(998) <= layer2_outputs(788);
    outputs(999) <= not(layer2_outputs(1396));
    outputs(1000) <= (layer2_outputs(2357)) and (layer2_outputs(251));
    outputs(1001) <= (layer2_outputs(1697)) and not (layer2_outputs(2348));
    outputs(1002) <= not(layer2_outputs(1867)) or (layer2_outputs(2165));
    outputs(1003) <= layer2_outputs(1323);
    outputs(1004) <= layer2_outputs(1687);
    outputs(1005) <= (layer2_outputs(1005)) and not (layer2_outputs(764));
    outputs(1006) <= (layer2_outputs(1416)) xor (layer2_outputs(145));
    outputs(1007) <= not(layer2_outputs(1809));
    outputs(1008) <= not((layer2_outputs(1522)) or (layer2_outputs(2048)));
    outputs(1009) <= (layer2_outputs(2500)) xor (layer2_outputs(1976));
    outputs(1010) <= not(layer2_outputs(2158)) or (layer2_outputs(736));
    outputs(1011) <= (layer2_outputs(1942)) and not (layer2_outputs(1316));
    outputs(1012) <= not(layer2_outputs(1510));
    outputs(1013) <= layer2_outputs(338);
    outputs(1014) <= (layer2_outputs(266)) and (layer2_outputs(585));
    outputs(1015) <= (layer2_outputs(1942)) and (layer2_outputs(1509));
    outputs(1016) <= not(layer2_outputs(988));
    outputs(1017) <= not(layer2_outputs(1481));
    outputs(1018) <= not(layer2_outputs(1506));
    outputs(1019) <= not(layer2_outputs(1641));
    outputs(1020) <= (layer2_outputs(2169)) and not (layer2_outputs(670));
    outputs(1021) <= (layer2_outputs(31)) and not (layer2_outputs(1379));
    outputs(1022) <= not(layer2_outputs(1100));
    outputs(1023) <= layer2_outputs(1389);
    outputs(1024) <= (layer2_outputs(2507)) and not (layer2_outputs(674));
    outputs(1025) <= (layer2_outputs(668)) and not (layer2_outputs(2365));
    outputs(1026) <= (layer2_outputs(1545)) and not (layer2_outputs(2229));
    outputs(1027) <= layer2_outputs(1366);
    outputs(1028) <= not(layer2_outputs(670));
    outputs(1029) <= layer2_outputs(2201);
    outputs(1030) <= layer2_outputs(143);
    outputs(1031) <= not((layer2_outputs(43)) or (layer2_outputs(625)));
    outputs(1032) <= (layer2_outputs(571)) and not (layer2_outputs(637));
    outputs(1033) <= layer2_outputs(1741);
    outputs(1034) <= not(layer2_outputs(182));
    outputs(1035) <= not(layer2_outputs(1749));
    outputs(1036) <= (layer2_outputs(2292)) and (layer2_outputs(1223));
    outputs(1037) <= not(layer2_outputs(92));
    outputs(1038) <= layer2_outputs(1695);
    outputs(1039) <= not((layer2_outputs(2278)) or (layer2_outputs(2390)));
    outputs(1040) <= (layer2_outputs(1751)) and not (layer2_outputs(2414));
    outputs(1041) <= (layer2_outputs(2144)) xor (layer2_outputs(1789));
    outputs(1042) <= layer2_outputs(2457);
    outputs(1043) <= layer2_outputs(1567);
    outputs(1044) <= not(layer2_outputs(1466));
    outputs(1045) <= not(layer2_outputs(5));
    outputs(1046) <= layer2_outputs(253);
    outputs(1047) <= not(layer2_outputs(1975));
    outputs(1048) <= not((layer2_outputs(48)) or (layer2_outputs(146)));
    outputs(1049) <= not(layer2_outputs(1700));
    outputs(1050) <= not(layer2_outputs(774)) or (layer2_outputs(958));
    outputs(1051) <= not(layer2_outputs(146));
    outputs(1052) <= layer2_outputs(6);
    outputs(1053) <= layer2_outputs(1178);
    outputs(1054) <= layer2_outputs(1997);
    outputs(1055) <= layer2_outputs(2128);
    outputs(1056) <= (layer2_outputs(767)) xor (layer2_outputs(1564));
    outputs(1057) <= not(layer2_outputs(389));
    outputs(1058) <= (layer2_outputs(1476)) xor (layer2_outputs(2496));
    outputs(1059) <= (layer2_outputs(2427)) or (layer2_outputs(2057));
    outputs(1060) <= not((layer2_outputs(278)) and (layer2_outputs(642)));
    outputs(1061) <= not(layer2_outputs(2473));
    outputs(1062) <= layer2_outputs(2487);
    outputs(1063) <= layer2_outputs(1091);
    outputs(1064) <= layer2_outputs(1020);
    outputs(1065) <= not(layer2_outputs(1221));
    outputs(1066) <= layer2_outputs(977);
    outputs(1067) <= not((layer2_outputs(1753)) or (layer2_outputs(2367)));
    outputs(1068) <= layer2_outputs(1351);
    outputs(1069) <= (layer2_outputs(2274)) or (layer2_outputs(2119));
    outputs(1070) <= (layer2_outputs(624)) or (layer2_outputs(1890));
    outputs(1071) <= not(layer2_outputs(326)) or (layer2_outputs(1838));
    outputs(1072) <= not(layer2_outputs(1415)) or (layer2_outputs(1161));
    outputs(1073) <= layer2_outputs(832);
    outputs(1074) <= not(layer2_outputs(2429));
    outputs(1075) <= layer2_outputs(873);
    outputs(1076) <= not((layer2_outputs(1013)) or (layer2_outputs(2436)));
    outputs(1077) <= not(layer2_outputs(477));
    outputs(1078) <= not(layer2_outputs(542));
    outputs(1079) <= not((layer2_outputs(2406)) or (layer2_outputs(2536)));
    outputs(1080) <= not(layer2_outputs(1712));
    outputs(1081) <= (layer2_outputs(818)) and not (layer2_outputs(1798));
    outputs(1082) <= layer2_outputs(400);
    outputs(1083) <= not(layer2_outputs(897));
    outputs(1084) <= not(layer2_outputs(1311));
    outputs(1085) <= not((layer2_outputs(1232)) or (layer2_outputs(990)));
    outputs(1086) <= layer2_outputs(1037);
    outputs(1087) <= layer2_outputs(568);
    outputs(1088) <= not(layer2_outputs(1426));
    outputs(1089) <= not(layer2_outputs(1247));
    outputs(1090) <= (layer2_outputs(1547)) and (layer2_outputs(533));
    outputs(1091) <= layer2_outputs(614);
    outputs(1092) <= layer2_outputs(39);
    outputs(1093) <= layer2_outputs(899);
    outputs(1094) <= not((layer2_outputs(1381)) xor (layer2_outputs(1617)));
    outputs(1095) <= (layer2_outputs(1854)) and not (layer2_outputs(578));
    outputs(1096) <= layer2_outputs(154);
    outputs(1097) <= layer2_outputs(1525);
    outputs(1098) <= not((layer2_outputs(2523)) and (layer2_outputs(1655)));
    outputs(1099) <= layer2_outputs(1857);
    outputs(1100) <= layer2_outputs(181);
    outputs(1101) <= layer2_outputs(1909);
    outputs(1102) <= not(layer2_outputs(491));
    outputs(1103) <= not(layer2_outputs(2504));
    outputs(1104) <= (layer2_outputs(2181)) and (layer2_outputs(2324));
    outputs(1105) <= not(layer2_outputs(1940)) or (layer2_outputs(2200));
    outputs(1106) <= layer2_outputs(1831);
    outputs(1107) <= (layer2_outputs(843)) and not (layer2_outputs(1994));
    outputs(1108) <= not(layer2_outputs(555));
    outputs(1109) <= (layer2_outputs(21)) and not (layer2_outputs(489));
    outputs(1110) <= (layer2_outputs(1672)) and not (layer2_outputs(623));
    outputs(1111) <= layer2_outputs(1396);
    outputs(1112) <= layer2_outputs(1786);
    outputs(1113) <= not(layer2_outputs(175));
    outputs(1114) <= not(layer2_outputs(635));
    outputs(1115) <= (layer2_outputs(1933)) and not (layer2_outputs(1497));
    outputs(1116) <= not(layer2_outputs(1761));
    outputs(1117) <= not(layer2_outputs(603));
    outputs(1118) <= (layer2_outputs(337)) and not (layer2_outputs(1753));
    outputs(1119) <= (layer2_outputs(2146)) xor (layer2_outputs(1391));
    outputs(1120) <= layer2_outputs(1283);
    outputs(1121) <= layer2_outputs(2377);
    outputs(1122) <= (layer2_outputs(1571)) and (layer2_outputs(1592));
    outputs(1123) <= layer2_outputs(374);
    outputs(1124) <= layer2_outputs(852);
    outputs(1125) <= (layer2_outputs(2255)) and not (layer2_outputs(1136));
    outputs(1126) <= (layer2_outputs(283)) and not (layer2_outputs(1232));
    outputs(1127) <= not(layer2_outputs(1445));
    outputs(1128) <= layer2_outputs(1909);
    outputs(1129) <= layer2_outputs(267);
    outputs(1130) <= not(layer2_outputs(1110));
    outputs(1131) <= layer2_outputs(1052);
    outputs(1132) <= not(layer2_outputs(296));
    outputs(1133) <= layer2_outputs(588);
    outputs(1134) <= not(layer2_outputs(1670));
    outputs(1135) <= layer2_outputs(1573);
    outputs(1136) <= not(layer2_outputs(2429));
    outputs(1137) <= (layer2_outputs(1418)) and (layer2_outputs(898));
    outputs(1138) <= not(layer2_outputs(1569));
    outputs(1139) <= not(layer2_outputs(2436));
    outputs(1140) <= layer2_outputs(222);
    outputs(1141) <= layer2_outputs(1790);
    outputs(1142) <= not(layer2_outputs(1290));
    outputs(1143) <= (layer2_outputs(817)) and (layer2_outputs(721));
    outputs(1144) <= not((layer2_outputs(188)) or (layer2_outputs(315)));
    outputs(1145) <= (layer2_outputs(460)) and (layer2_outputs(1813));
    outputs(1146) <= layer2_outputs(0);
    outputs(1147) <= not((layer2_outputs(1152)) or (layer2_outputs(1345)));
    outputs(1148) <= (layer2_outputs(2293)) and not (layer2_outputs(955));
    outputs(1149) <= layer2_outputs(2169);
    outputs(1150) <= layer2_outputs(1547);
    outputs(1151) <= layer2_outputs(1482);
    outputs(1152) <= layer2_outputs(1895);
    outputs(1153) <= not(layer2_outputs(2214));
    outputs(1154) <= not(layer2_outputs(780));
    outputs(1155) <= layer2_outputs(2032);
    outputs(1156) <= layer2_outputs(2475);
    outputs(1157) <= not((layer2_outputs(563)) and (layer2_outputs(1788)));
    outputs(1158) <= (layer2_outputs(662)) xor (layer2_outputs(2235));
    outputs(1159) <= not(layer2_outputs(2020));
    outputs(1160) <= layer2_outputs(1932);
    outputs(1161) <= layer2_outputs(952);
    outputs(1162) <= layer2_outputs(1926);
    outputs(1163) <= not(layer2_outputs(2557)) or (layer2_outputs(2520));
    outputs(1164) <= not(layer2_outputs(549));
    outputs(1165) <= layer2_outputs(27);
    outputs(1166) <= not((layer2_outputs(520)) xor (layer2_outputs(860)));
    outputs(1167) <= layer2_outputs(1895);
    outputs(1168) <= layer2_outputs(2465);
    outputs(1169) <= layer2_outputs(1573);
    outputs(1170) <= layer2_outputs(1552);
    outputs(1171) <= (layer2_outputs(559)) and not (layer2_outputs(1112));
    outputs(1172) <= not(layer2_outputs(882)) or (layer2_outputs(1399));
    outputs(1173) <= layer2_outputs(386);
    outputs(1174) <= not(layer2_outputs(608));
    outputs(1175) <= (layer2_outputs(1665)) xor (layer2_outputs(1123));
    outputs(1176) <= not(layer2_outputs(1851));
    outputs(1177) <= not(layer2_outputs(2442));
    outputs(1178) <= layer2_outputs(471);
    outputs(1179) <= not(layer2_outputs(2102)) or (layer2_outputs(300));
    outputs(1180) <= (layer2_outputs(1789)) and not (layer2_outputs(1328));
    outputs(1181) <= layer2_outputs(594);
    outputs(1182) <= (layer2_outputs(2174)) xor (layer2_outputs(2251));
    outputs(1183) <= not(layer2_outputs(740));
    outputs(1184) <= not(layer2_outputs(2136));
    outputs(1185) <= (layer2_outputs(475)) and not (layer2_outputs(2510));
    outputs(1186) <= (layer2_outputs(1071)) xor (layer2_outputs(1279));
    outputs(1187) <= not(layer2_outputs(2245));
    outputs(1188) <= not(layer2_outputs(477));
    outputs(1189) <= (layer2_outputs(1494)) or (layer2_outputs(1768));
    outputs(1190) <= (layer2_outputs(396)) and (layer2_outputs(530));
    outputs(1191) <= layer2_outputs(1997);
    outputs(1192) <= layer2_outputs(1747);
    outputs(1193) <= not(layer2_outputs(1794));
    outputs(1194) <= layer2_outputs(474);
    outputs(1195) <= layer2_outputs(422);
    outputs(1196) <= not(layer2_outputs(1647));
    outputs(1197) <= (layer2_outputs(2059)) xor (layer2_outputs(1045));
    outputs(1198) <= layer2_outputs(343);
    outputs(1199) <= not(layer2_outputs(1784));
    outputs(1200) <= (layer2_outputs(1691)) and not (layer2_outputs(359));
    outputs(1201) <= not(layer2_outputs(2374));
    outputs(1202) <= not(layer2_outputs(325));
    outputs(1203) <= layer2_outputs(1291);
    outputs(1204) <= not(layer2_outputs(2268));
    outputs(1205) <= layer2_outputs(2525);
    outputs(1206) <= layer2_outputs(975);
    outputs(1207) <= not(layer2_outputs(1336));
    outputs(1208) <= not(layer2_outputs(1469));
    outputs(1209) <= (layer2_outputs(1359)) xor (layer2_outputs(2008));
    outputs(1210) <= layer2_outputs(1103);
    outputs(1211) <= not(layer2_outputs(246));
    outputs(1212) <= layer2_outputs(1277);
    outputs(1213) <= not(layer2_outputs(2089));
    outputs(1214) <= layer2_outputs(1315);
    outputs(1215) <= layer2_outputs(1293);
    outputs(1216) <= not(layer2_outputs(217));
    outputs(1217) <= not(layer2_outputs(1667)) or (layer2_outputs(1678));
    outputs(1218) <= not(layer2_outputs(452));
    outputs(1219) <= (layer2_outputs(170)) and not (layer2_outputs(1490));
    outputs(1220) <= (layer2_outputs(629)) and not (layer2_outputs(83));
    outputs(1221) <= layer2_outputs(1269);
    outputs(1222) <= layer2_outputs(2160);
    outputs(1223) <= layer2_outputs(2004);
    outputs(1224) <= not(layer2_outputs(2267));
    outputs(1225) <= not(layer2_outputs(2227));
    outputs(1226) <= (layer2_outputs(2491)) and not (layer2_outputs(82));
    outputs(1227) <= layer2_outputs(239);
    outputs(1228) <= not(layer2_outputs(1230));
    outputs(1229) <= layer2_outputs(2423);
    outputs(1230) <= layer2_outputs(1178);
    outputs(1231) <= not(layer2_outputs(566));
    outputs(1232) <= not(layer2_outputs(1493));
    outputs(1233) <= (layer2_outputs(845)) and not (layer2_outputs(1823));
    outputs(1234) <= layer2_outputs(2240);
    outputs(1235) <= (layer2_outputs(1945)) and not (layer2_outputs(2446));
    outputs(1236) <= not(layer2_outputs(1468));
    outputs(1237) <= not(layer2_outputs(1096));
    outputs(1238) <= not(layer2_outputs(1900));
    outputs(1239) <= layer2_outputs(1810);
    outputs(1240) <= not(layer2_outputs(1179));
    outputs(1241) <= (layer2_outputs(2379)) and not (layer2_outputs(2244));
    outputs(1242) <= not(layer2_outputs(809));
    outputs(1243) <= layer2_outputs(661);
    outputs(1244) <= not(layer2_outputs(175));
    outputs(1245) <= (layer2_outputs(1559)) and (layer2_outputs(1545));
    outputs(1246) <= (layer2_outputs(1554)) and (layer2_outputs(1978));
    outputs(1247) <= layer2_outputs(879);
    outputs(1248) <= not(layer2_outputs(953));
    outputs(1249) <= not(layer2_outputs(2336));
    outputs(1250) <= not(layer2_outputs(532));
    outputs(1251) <= not(layer2_outputs(695));
    outputs(1252) <= not(layer2_outputs(136));
    outputs(1253) <= layer2_outputs(1765);
    outputs(1254) <= not(layer2_outputs(476));
    outputs(1255) <= layer2_outputs(1061);
    outputs(1256) <= not(layer2_outputs(66));
    outputs(1257) <= layer2_outputs(238);
    outputs(1258) <= not((layer2_outputs(1980)) or (layer2_outputs(452)));
    outputs(1259) <= (layer2_outputs(2067)) and (layer2_outputs(1797));
    outputs(1260) <= not(layer2_outputs(1637));
    outputs(1261) <= layer2_outputs(2458);
    outputs(1262) <= (layer2_outputs(848)) and not (layer2_outputs(1687));
    outputs(1263) <= layer2_outputs(2553);
    outputs(1264) <= not(layer2_outputs(1735));
    outputs(1265) <= not((layer2_outputs(1127)) and (layer2_outputs(735)));
    outputs(1266) <= (layer2_outputs(2058)) and (layer2_outputs(1659));
    outputs(1267) <= not((layer2_outputs(778)) xor (layer2_outputs(2386)));
    outputs(1268) <= (layer2_outputs(268)) and not (layer2_outputs(245));
    outputs(1269) <= (layer2_outputs(355)) and not (layer2_outputs(235));
    outputs(1270) <= layer2_outputs(1222);
    outputs(1271) <= not(layer2_outputs(1841));
    outputs(1272) <= layer2_outputs(2065);
    outputs(1273) <= (layer2_outputs(1472)) and not (layer2_outputs(2163));
    outputs(1274) <= layer2_outputs(2375);
    outputs(1275) <= not((layer2_outputs(653)) xor (layer2_outputs(2462)));
    outputs(1276) <= not(layer2_outputs(566));
    outputs(1277) <= layer2_outputs(2545);
    outputs(1278) <= layer2_outputs(2312);
    outputs(1279) <= not(layer2_outputs(1629));
    outputs(1280) <= (layer2_outputs(2514)) xor (layer2_outputs(1184));
    outputs(1281) <= layer2_outputs(962);
    outputs(1282) <= not((layer2_outputs(1207)) and (layer2_outputs(1239)));
    outputs(1283) <= (layer2_outputs(967)) xor (layer2_outputs(910));
    outputs(1284) <= not(layer2_outputs(2165));
    outputs(1285) <= layer2_outputs(2037);
    outputs(1286) <= not((layer2_outputs(1007)) xor (layer2_outputs(409)));
    outputs(1287) <= layer2_outputs(2137);
    outputs(1288) <= layer2_outputs(1263);
    outputs(1289) <= not((layer2_outputs(97)) xor (layer2_outputs(739)));
    outputs(1290) <= not(layer2_outputs(1734));
    outputs(1291) <= layer2_outputs(909);
    outputs(1292) <= (layer2_outputs(791)) xor (layer2_outputs(159));
    outputs(1293) <= (layer2_outputs(1308)) or (layer2_outputs(1926));
    outputs(1294) <= not(layer2_outputs(2013)) or (layer2_outputs(2115));
    outputs(1295) <= layer2_outputs(1679);
    outputs(1296) <= not(layer2_outputs(1131));
    outputs(1297) <= (layer2_outputs(331)) and (layer2_outputs(1991));
    outputs(1298) <= (layer2_outputs(1923)) and not (layer2_outputs(1406));
    outputs(1299) <= (layer2_outputs(522)) xor (layer2_outputs(73));
    outputs(1300) <= not(layer2_outputs(2276));
    outputs(1301) <= layer2_outputs(2012);
    outputs(1302) <= layer2_outputs(2101);
    outputs(1303) <= layer2_outputs(1115);
    outputs(1304) <= layer2_outputs(980);
    outputs(1305) <= not(layer2_outputs(2469));
    outputs(1306) <= not(layer2_outputs(1944));
    outputs(1307) <= layer2_outputs(755);
    outputs(1308) <= not(layer2_outputs(508));
    outputs(1309) <= layer2_outputs(1174);
    outputs(1310) <= (layer2_outputs(2175)) and not (layer2_outputs(226));
    outputs(1311) <= not(layer2_outputs(1225));
    outputs(1312) <= layer2_outputs(749);
    outputs(1313) <= not(layer2_outputs(636));
    outputs(1314) <= not(layer2_outputs(151));
    outputs(1315) <= (layer2_outputs(2271)) and not (layer2_outputs(1485));
    outputs(1316) <= not((layer2_outputs(2368)) or (layer2_outputs(1171)));
    outputs(1317) <= not(layer2_outputs(54));
    outputs(1318) <= not(layer2_outputs(842));
    outputs(1319) <= (layer2_outputs(926)) and not (layer2_outputs(1796));
    outputs(1320) <= not(layer2_outputs(1538));
    outputs(1321) <= (layer2_outputs(2269)) and (layer2_outputs(1530));
    outputs(1322) <= layer2_outputs(1093);
    outputs(1323) <= layer2_outputs(601);
    outputs(1324) <= not(layer2_outputs(2063));
    outputs(1325) <= not(layer2_outputs(323)) or (layer2_outputs(1653));
    outputs(1326) <= layer2_outputs(42);
    outputs(1327) <= layer2_outputs(1005);
    outputs(1328) <= (layer2_outputs(875)) xor (layer2_outputs(1435));
    outputs(1329) <= not((layer2_outputs(2042)) or (layer2_outputs(2027)));
    outputs(1330) <= (layer2_outputs(456)) xor (layer2_outputs(2033));
    outputs(1331) <= (layer2_outputs(1203)) or (layer2_outputs(1600));
    outputs(1332) <= (layer2_outputs(1970)) xor (layer2_outputs(1009));
    outputs(1333) <= layer2_outputs(1775);
    outputs(1334) <= not((layer2_outputs(2209)) or (layer2_outputs(685)));
    outputs(1335) <= layer2_outputs(2180);
    outputs(1336) <= not((layer2_outputs(2050)) xor (layer2_outputs(2043)));
    outputs(1337) <= (layer2_outputs(2009)) xor (layer2_outputs(1864));
    outputs(1338) <= (layer2_outputs(1102)) and not (layer2_outputs(592));
    outputs(1339) <= not(layer2_outputs(1464));
    outputs(1340) <= (layer2_outputs(625)) and not (layer2_outputs(896));
    outputs(1341) <= not(layer2_outputs(1565));
    outputs(1342) <= layer2_outputs(217);
    outputs(1343) <= not(layer2_outputs(1432));
    outputs(1344) <= not((layer2_outputs(324)) xor (layer2_outputs(1643)));
    outputs(1345) <= layer2_outputs(403);
    outputs(1346) <= layer2_outputs(999);
    outputs(1347) <= not((layer2_outputs(517)) and (layer2_outputs(260)));
    outputs(1348) <= not(layer2_outputs(849));
    outputs(1349) <= (layer2_outputs(402)) xor (layer2_outputs(1708));
    outputs(1350) <= not((layer2_outputs(356)) or (layer2_outputs(2265)));
    outputs(1351) <= not(layer2_outputs(753));
    outputs(1352) <= layer2_outputs(2105);
    outputs(1353) <= (layer2_outputs(826)) xor (layer2_outputs(145));
    outputs(1354) <= layer2_outputs(1826);
    outputs(1355) <= not(layer2_outputs(1693));
    outputs(1356) <= (layer2_outputs(282)) or (layer2_outputs(1597));
    outputs(1357) <= layer2_outputs(2542);
    outputs(1358) <= not(layer2_outputs(1300));
    outputs(1359) <= layer2_outputs(304);
    outputs(1360) <= not(layer2_outputs(2151)) or (layer2_outputs(70));
    outputs(1361) <= not((layer2_outputs(194)) and (layer2_outputs(2454)));
    outputs(1362) <= layer2_outputs(442);
    outputs(1363) <= layer2_outputs(1288);
    outputs(1364) <= layer2_outputs(1470);
    outputs(1365) <= not(layer2_outputs(1772));
    outputs(1366) <= not(layer2_outputs(265));
    outputs(1367) <= (layer2_outputs(1960)) xor (layer2_outputs(531));
    outputs(1368) <= layer2_outputs(1202);
    outputs(1369) <= layer2_outputs(547);
    outputs(1370) <= layer2_outputs(1508);
    outputs(1371) <= layer2_outputs(1217);
    outputs(1372) <= layer2_outputs(1471);
    outputs(1373) <= not(layer2_outputs(349));
    outputs(1374) <= not(layer2_outputs(726));
    outputs(1375) <= not(layer2_outputs(1945));
    outputs(1376) <= layer2_outputs(2149);
    outputs(1377) <= (layer2_outputs(956)) and (layer2_outputs(1282));
    outputs(1378) <= layer2_outputs(1721);
    outputs(1379) <= layer2_outputs(472);
    outputs(1380) <= layer2_outputs(673);
    outputs(1381) <= not((layer2_outputs(1882)) xor (layer2_outputs(1914)));
    outputs(1382) <= layer2_outputs(2329);
    outputs(1383) <= not(layer2_outputs(859));
    outputs(1384) <= layer2_outputs(482);
    outputs(1385) <= (layer2_outputs(771)) and not (layer2_outputs(141));
    outputs(1386) <= layer2_outputs(1101);
    outputs(1387) <= not(layer2_outputs(1818));
    outputs(1388) <= not(layer2_outputs(228)) or (layer2_outputs(1183));
    outputs(1389) <= not(layer2_outputs(333));
    outputs(1390) <= not((layer2_outputs(2398)) xor (layer2_outputs(474)));
    outputs(1391) <= layer2_outputs(2104);
    outputs(1392) <= not(layer2_outputs(1569));
    outputs(1393) <= not((layer2_outputs(165)) and (layer2_outputs(1506)));
    outputs(1394) <= (layer2_outputs(1520)) and not (layer2_outputs(879));
    outputs(1395) <= not((layer2_outputs(79)) xor (layer2_outputs(2499)));
    outputs(1396) <= not(layer2_outputs(1042));
    outputs(1397) <= not((layer2_outputs(1265)) or (layer2_outputs(1107)));
    outputs(1398) <= not(layer2_outputs(1327));
    outputs(1399) <= not((layer2_outputs(112)) or (layer2_outputs(1488)));
    outputs(1400) <= (layer2_outputs(2148)) and (layer2_outputs(2083));
    outputs(1401) <= not((layer2_outputs(1256)) or (layer2_outputs(2041)));
    outputs(1402) <= layer2_outputs(884);
    outputs(1403) <= layer2_outputs(300);
    outputs(1404) <= not(layer2_outputs(185));
    outputs(1405) <= layer2_outputs(2303);
    outputs(1406) <= layer2_outputs(1968);
    outputs(1407) <= (layer2_outputs(162)) xor (layer2_outputs(890));
    outputs(1408) <= layer2_outputs(472);
    outputs(1409) <= not(layer2_outputs(1766));
    outputs(1410) <= (layer2_outputs(1526)) or (layer2_outputs(1543));
    outputs(1411) <= not(layer2_outputs(528)) or (layer2_outputs(1522));
    outputs(1412) <= layer2_outputs(981);
    outputs(1413) <= layer2_outputs(920);
    outputs(1414) <= (layer2_outputs(1433)) xor (layer2_outputs(965));
    outputs(1415) <= not(layer2_outputs(2068));
    outputs(1416) <= (layer2_outputs(133)) and not (layer2_outputs(1959));
    outputs(1417) <= layer2_outputs(929);
    outputs(1418) <= (layer2_outputs(346)) xor (layer2_outputs(2052));
    outputs(1419) <= (layer2_outputs(607)) and not (layer2_outputs(690));
    outputs(1420) <= not(layer2_outputs(1793)) or (layer2_outputs(2123));
    outputs(1421) <= (layer2_outputs(1575)) and not (layer2_outputs(32));
    outputs(1422) <= layer2_outputs(1149);
    outputs(1423) <= not((layer2_outputs(2063)) or (layer2_outputs(497)));
    outputs(1424) <= layer2_outputs(2044);
    outputs(1425) <= layer2_outputs(184);
    outputs(1426) <= layer2_outputs(1439);
    outputs(1427) <= not(layer2_outputs(770)) or (layer2_outputs(1528));
    outputs(1428) <= not(layer2_outputs(2275));
    outputs(1429) <= layer2_outputs(1288);
    outputs(1430) <= not(layer2_outputs(1759));
    outputs(1431) <= layer2_outputs(1012);
    outputs(1432) <= layer2_outputs(42);
    outputs(1433) <= not(layer2_outputs(2187));
    outputs(1434) <= not((layer2_outputs(612)) and (layer2_outputs(708)));
    outputs(1435) <= not(layer2_outputs(2077));
    outputs(1436) <= layer2_outputs(1115);
    outputs(1437) <= (layer2_outputs(649)) and (layer2_outputs(1825));
    outputs(1438) <= not(layer2_outputs(1555));
    outputs(1439) <= not(layer2_outputs(334));
    outputs(1440) <= (layer2_outputs(152)) and not (layer2_outputs(1996));
    outputs(1441) <= not(layer2_outputs(865));
    outputs(1442) <= not((layer2_outputs(972)) xor (layer2_outputs(68)));
    outputs(1443) <= (layer2_outputs(1803)) and not (layer2_outputs(2116));
    outputs(1444) <= not((layer2_outputs(1229)) or (layer2_outputs(597)));
    outputs(1445) <= not(layer2_outputs(461));
    outputs(1446) <= not(layer2_outputs(775));
    outputs(1447) <= not(layer2_outputs(2371));
    outputs(1448) <= layer2_outputs(2126);
    outputs(1449) <= layer2_outputs(96);
    outputs(1450) <= (layer2_outputs(2253)) and (layer2_outputs(1043));
    outputs(1451) <= not((layer2_outputs(2256)) or (layer2_outputs(1948)));
    outputs(1452) <= layer2_outputs(2296);
    outputs(1453) <= (layer2_outputs(1450)) and (layer2_outputs(653));
    outputs(1454) <= not(layer2_outputs(2194));
    outputs(1455) <= not(layer2_outputs(507));
    outputs(1456) <= not((layer2_outputs(894)) xor (layer2_outputs(781)));
    outputs(1457) <= not(layer2_outputs(1943));
    outputs(1458) <= not((layer2_outputs(164)) or (layer2_outputs(646)));
    outputs(1459) <= not(layer2_outputs(1128));
    outputs(1460) <= (layer2_outputs(1602)) and not (layer2_outputs(752));
    outputs(1461) <= not((layer2_outputs(1456)) xor (layer2_outputs(427)));
    outputs(1462) <= layer2_outputs(880);
    outputs(1463) <= not((layer2_outputs(1401)) xor (layer2_outputs(1360)));
    outputs(1464) <= not(layer2_outputs(754));
    outputs(1465) <= (layer2_outputs(525)) xor (layer2_outputs(73));
    outputs(1466) <= layer2_outputs(1951);
    outputs(1467) <= (layer2_outputs(1467)) xor (layer2_outputs(41));
    outputs(1468) <= layer2_outputs(2313);
    outputs(1469) <= not(layer2_outputs(827));
    outputs(1470) <= layer2_outputs(799);
    outputs(1471) <= (layer2_outputs(1276)) xor (layer2_outputs(1618));
    outputs(1472) <= not((layer2_outputs(2023)) and (layer2_outputs(1060)));
    outputs(1473) <= (layer2_outputs(579)) and (layer2_outputs(1109));
    outputs(1474) <= (layer2_outputs(316)) and not (layer2_outputs(1837));
    outputs(1475) <= not(layer2_outputs(834));
    outputs(1476) <= (layer2_outputs(2145)) or (layer2_outputs(2261));
    outputs(1477) <= not((layer2_outputs(822)) xor (layer2_outputs(1712)));
    outputs(1478) <= not(layer2_outputs(38));
    outputs(1479) <= layer2_outputs(136);
    outputs(1480) <= not((layer2_outputs(267)) xor (layer2_outputs(1929)));
    outputs(1481) <= not((layer2_outputs(1489)) xor (layer2_outputs(50)));
    outputs(1482) <= (layer2_outputs(130)) or (layer2_outputs(884));
    outputs(1483) <= layer2_outputs(1762);
    outputs(1484) <= not(layer2_outputs(2143));
    outputs(1485) <= not((layer2_outputs(221)) or (layer2_outputs(630)));
    outputs(1486) <= not(layer2_outputs(1676));
    outputs(1487) <= not(layer2_outputs(750));
    outputs(1488) <= layer2_outputs(934);
    outputs(1489) <= not(layer2_outputs(115));
    outputs(1490) <= layer2_outputs(1491);
    outputs(1491) <= not(layer2_outputs(1257)) or (layer2_outputs(223));
    outputs(1492) <= not((layer2_outputs(1128)) xor (layer2_outputs(1742)));
    outputs(1493) <= layer2_outputs(836);
    outputs(1494) <= not(layer2_outputs(115)) or (layer2_outputs(416));
    outputs(1495) <= layer2_outputs(722);
    outputs(1496) <= not(layer2_outputs(72));
    outputs(1497) <= (layer2_outputs(1238)) xor (layer2_outputs(1207));
    outputs(1498) <= layer2_outputs(1213);
    outputs(1499) <= not((layer2_outputs(2197)) xor (layer2_outputs(1821)));
    outputs(1500) <= not(layer2_outputs(1899));
    outputs(1501) <= (layer2_outputs(2343)) xor (layer2_outputs(1527));
    outputs(1502) <= not(layer2_outputs(2369));
    outputs(1503) <= layer2_outputs(788);
    outputs(1504) <= not(layer2_outputs(1194));
    outputs(1505) <= layer2_outputs(740);
    outputs(1506) <= layer2_outputs(227);
    outputs(1507) <= not(layer2_outputs(215));
    outputs(1508) <= not((layer2_outputs(2295)) or (layer2_outputs(1375)));
    outputs(1509) <= not(layer2_outputs(889));
    outputs(1510) <= layer2_outputs(1248);
    outputs(1511) <= not((layer2_outputs(2087)) xor (layer2_outputs(210)));
    outputs(1512) <= layer2_outputs(1690);
    outputs(1513) <= not((layer2_outputs(1590)) or (layer2_outputs(745)));
    outputs(1514) <= not(layer2_outputs(2133));
    outputs(1515) <= not(layer2_outputs(678)) or (layer2_outputs(289));
    outputs(1516) <= layer2_outputs(1102);
    outputs(1517) <= (layer2_outputs(1268)) and not (layer2_outputs(1352));
    outputs(1518) <= layer2_outputs(1318);
    outputs(1519) <= layer2_outputs(2346);
    outputs(1520) <= layer2_outputs(914);
    outputs(1521) <= not(layer2_outputs(1084));
    outputs(1522) <= (layer2_outputs(2325)) xor (layer2_outputs(2211));
    outputs(1523) <= not(layer2_outputs(261));
    outputs(1524) <= (layer2_outputs(1192)) and not (layer2_outputs(935));
    outputs(1525) <= not((layer2_outputs(1802)) and (layer2_outputs(1630)));
    outputs(1526) <= not(layer2_outputs(2254));
    outputs(1527) <= layer2_outputs(838);
    outputs(1528) <= (layer2_outputs(238)) xor (layer2_outputs(2490));
    outputs(1529) <= layer2_outputs(231);
    outputs(1530) <= not(layer2_outputs(2166));
    outputs(1531) <= not(layer2_outputs(1187)) or (layer2_outputs(2056));
    outputs(1532) <= (layer2_outputs(1430)) and not (layer2_outputs(943));
    outputs(1533) <= (layer2_outputs(1598)) and not (layer2_outputs(1014));
    outputs(1534) <= layer2_outputs(2005);
    outputs(1535) <= not((layer2_outputs(2234)) xor (layer2_outputs(1459)));
    outputs(1536) <= not(layer2_outputs(368));
    outputs(1537) <= layer2_outputs(844);
    outputs(1538) <= not(layer2_outputs(1708));
    outputs(1539) <= layer2_outputs(1465);
    outputs(1540) <= not(layer2_outputs(1710));
    outputs(1541) <= layer2_outputs(1956);
    outputs(1542) <= layer2_outputs(183);
    outputs(1543) <= (layer2_outputs(1919)) and (layer2_outputs(2512));
    outputs(1544) <= not(layer2_outputs(1863));
    outputs(1545) <= not(layer2_outputs(348));
    outputs(1546) <= not(layer2_outputs(833)) or (layer2_outputs(364));
    outputs(1547) <= layer2_outputs(2514);
    outputs(1548) <= layer2_outputs(2407);
    outputs(1549) <= not(layer2_outputs(2253));
    outputs(1550) <= not((layer2_outputs(1446)) or (layer2_outputs(1235)));
    outputs(1551) <= not(layer2_outputs(2113));
    outputs(1552) <= not(layer2_outputs(1260));
    outputs(1553) <= layer2_outputs(98);
    outputs(1554) <= not(layer2_outputs(2521));
    outputs(1555) <= (layer2_outputs(1297)) and not (layer2_outputs(2502));
    outputs(1556) <= (layer2_outputs(176)) and not (layer2_outputs(394));
    outputs(1557) <= (layer2_outputs(825)) and not (layer2_outputs(1216));
    outputs(1558) <= not((layer2_outputs(1229)) or (layer2_outputs(1946)));
    outputs(1559) <= not(layer2_outputs(396));
    outputs(1560) <= not((layer2_outputs(1959)) or (layer2_outputs(2060)));
    outputs(1561) <= not(layer2_outputs(490));
    outputs(1562) <= not(layer2_outputs(615));
    outputs(1563) <= not(layer2_outputs(847));
    outputs(1564) <= layer2_outputs(2179);
    outputs(1565) <= not(layer2_outputs(1139));
    outputs(1566) <= (layer2_outputs(2544)) and not (layer2_outputs(425));
    outputs(1567) <= not((layer2_outputs(1872)) or (layer2_outputs(1816)));
    outputs(1568) <= layer2_outputs(536);
    outputs(1569) <= not(layer2_outputs(1955));
    outputs(1570) <= layer2_outputs(1185);
    outputs(1571) <= (layer2_outputs(2117)) and not (layer2_outputs(1937));
    outputs(1572) <= not((layer2_outputs(1141)) xor (layer2_outputs(105)));
    outputs(1573) <= not(layer2_outputs(1801));
    outputs(1574) <= not(layer2_outputs(2519));
    outputs(1575) <= not(layer2_outputs(1495));
    outputs(1576) <= not(layer2_outputs(1377)) or (layer2_outputs(45));
    outputs(1577) <= not(layer2_outputs(741));
    outputs(1578) <= not((layer2_outputs(1035)) or (layer2_outputs(878)));
    outputs(1579) <= (layer2_outputs(1889)) and (layer2_outputs(1422));
    outputs(1580) <= not(layer2_outputs(1154));
    outputs(1581) <= not(layer2_outputs(1208));
    outputs(1582) <= not((layer2_outputs(1764)) or (layer2_outputs(1369)));
    outputs(1583) <= layer2_outputs(1339);
    outputs(1584) <= (layer2_outputs(2151)) and not (layer2_outputs(1155));
    outputs(1585) <= not(layer2_outputs(757));
    outputs(1586) <= layer2_outputs(1204);
    outputs(1587) <= not(layer2_outputs(1191));
    outputs(1588) <= layer2_outputs(392);
    outputs(1589) <= not(layer2_outputs(1552));
    outputs(1590) <= layer2_outputs(1930);
    outputs(1591) <= not(layer2_outputs(394));
    outputs(1592) <= layer2_outputs(2331);
    outputs(1593) <= layer2_outputs(293);
    outputs(1594) <= (layer2_outputs(180)) xor (layer2_outputs(281));
    outputs(1595) <= (layer2_outputs(665)) and not (layer2_outputs(2040));
    outputs(1596) <= layer2_outputs(110);
    outputs(1597) <= (layer2_outputs(577)) and not (layer2_outputs(795));
    outputs(1598) <= not(layer2_outputs(779));
    outputs(1599) <= not(layer2_outputs(1886));
    outputs(1600) <= not(layer2_outputs(1751));
    outputs(1601) <= (layer2_outputs(2396)) and (layer2_outputs(432));
    outputs(1602) <= not(layer2_outputs(1597));
    outputs(1603) <= not(layer2_outputs(181));
    outputs(1604) <= (layer2_outputs(2216)) and not (layer2_outputs(1875));
    outputs(1605) <= layer2_outputs(446);
    outputs(1606) <= not(layer2_outputs(2538));
    outputs(1607) <= layer2_outputs(2181);
    outputs(1608) <= not((layer2_outputs(2533)) or (layer2_outputs(1054)));
    outputs(1609) <= not((layer2_outputs(1500)) or (layer2_outputs(1277)));
    outputs(1610) <= not(layer2_outputs(1527));
    outputs(1611) <= layer2_outputs(204);
    outputs(1612) <= layer2_outputs(746);
    outputs(1613) <= layer2_outputs(98);
    outputs(1614) <= not((layer2_outputs(798)) or (layer2_outputs(1453)));
    outputs(1615) <= not(layer2_outputs(309));
    outputs(1616) <= not(layer2_outputs(2356)) or (layer2_outputs(761));
    outputs(1617) <= not(layer2_outputs(2121));
    outputs(1618) <= layer2_outputs(1181);
    outputs(1619) <= not(layer2_outputs(2094)) or (layer2_outputs(1492));
    outputs(1620) <= layer2_outputs(1395);
    outputs(1621) <= layer2_outputs(1151);
    outputs(1622) <= not(layer2_outputs(526));
    outputs(1623) <= not((layer2_outputs(1972)) xor (layer2_outputs(164)));
    outputs(1624) <= not(layer2_outputs(1445));
    outputs(1625) <= layer2_outputs(408);
    outputs(1626) <= not((layer2_outputs(240)) or (layer2_outputs(1695)));
    outputs(1627) <= layer2_outputs(720);
    outputs(1628) <= not(layer2_outputs(1113));
    outputs(1629) <= layer2_outputs(978);
    outputs(1630) <= layer2_outputs(1971);
    outputs(1631) <= not(layer2_outputs(2548));
    outputs(1632) <= not(layer2_outputs(1335));
    outputs(1633) <= not(layer2_outputs(857));
    outputs(1634) <= layer2_outputs(744);
    outputs(1635) <= not(layer2_outputs(523));
    outputs(1636) <= layer2_outputs(2553);
    outputs(1637) <= (layer2_outputs(1820)) and (layer2_outputs(2056));
    outputs(1638) <= not(layer2_outputs(462));
    outputs(1639) <= not((layer2_outputs(581)) xor (layer2_outputs(1628)));
    outputs(1640) <= not(layer2_outputs(354));
    outputs(1641) <= not(layer2_outputs(1027));
    outputs(1642) <= not((layer2_outputs(286)) or (layer2_outputs(880)));
    outputs(1643) <= not((layer2_outputs(1068)) xor (layer2_outputs(998)));
    outputs(1644) <= (layer2_outputs(51)) xor (layer2_outputs(709));
    outputs(1645) <= (layer2_outputs(2049)) and (layer2_outputs(2335));
    outputs(1646) <= not(layer2_outputs(2285));
    outputs(1647) <= layer2_outputs(577);
    outputs(1648) <= layer2_outputs(473);
    outputs(1649) <= layer2_outputs(1047);
    outputs(1650) <= layer2_outputs(730);
    outputs(1651) <= layer2_outputs(2065);
    outputs(1652) <= layer2_outputs(15);
    outputs(1653) <= (layer2_outputs(1297)) and (layer2_outputs(1234));
    outputs(1654) <= (layer2_outputs(19)) and not (layer2_outputs(966));
    outputs(1655) <= (layer2_outputs(445)) xor (layer2_outputs(1126));
    outputs(1656) <= not(layer2_outputs(2228));
    outputs(1657) <= not(layer2_outputs(1664));
    outputs(1658) <= layer2_outputs(1475);
    outputs(1659) <= not(layer2_outputs(840));
    outputs(1660) <= layer2_outputs(1032);
    outputs(1661) <= not(layer2_outputs(2318));
    outputs(1662) <= not((layer2_outputs(335)) xor (layer2_outputs(277)));
    outputs(1663) <= (layer2_outputs(881)) and not (layer2_outputs(286));
    outputs(1664) <= layer2_outputs(1081);
    outputs(1665) <= layer2_outputs(455);
    outputs(1666) <= (layer2_outputs(2105)) xor (layer2_outputs(1368));
    outputs(1667) <= layer2_outputs(1037);
    outputs(1668) <= not(layer2_outputs(1922));
    outputs(1669) <= layer2_outputs(534);
    outputs(1670) <= (layer2_outputs(121)) or (layer2_outputs(1024));
    outputs(1671) <= not((layer2_outputs(1267)) or (layer2_outputs(2074)));
    outputs(1672) <= (layer2_outputs(2007)) and (layer2_outputs(1805));
    outputs(1673) <= (layer2_outputs(249)) and not (layer2_outputs(1907));
    outputs(1674) <= not(layer2_outputs(1290));
    outputs(1675) <= layer2_outputs(1767);
    outputs(1676) <= layer2_outputs(481);
    outputs(1677) <= layer2_outputs(208);
    outputs(1678) <= (layer2_outputs(1615)) and (layer2_outputs(414));
    outputs(1679) <= (layer2_outputs(2488)) and not (layer2_outputs(883));
    outputs(1680) <= not(layer2_outputs(114)) or (layer2_outputs(2111));
    outputs(1681) <= (layer2_outputs(1271)) and not (layer2_outputs(1776));
    outputs(1682) <= not(layer2_outputs(2476));
    outputs(1683) <= not(layer2_outputs(1139));
    outputs(1684) <= not(layer2_outputs(1769)) or (layer2_outputs(915));
    outputs(1685) <= layer2_outputs(1314);
    outputs(1686) <= layer2_outputs(982);
    outputs(1687) <= not(layer2_outputs(104));
    outputs(1688) <= (layer2_outputs(122)) and not (layer2_outputs(1631));
    outputs(1689) <= not((layer2_outputs(272)) xor (layer2_outputs(1404)));
    outputs(1690) <= not(layer2_outputs(1113));
    outputs(1691) <= not(layer2_outputs(725));
    outputs(1692) <= layer2_outputs(876);
    outputs(1693) <= layer2_outputs(1471);
    outputs(1694) <= (layer2_outputs(780)) and (layer2_outputs(1220));
    outputs(1695) <= layer2_outputs(2184);
    outputs(1696) <= not((layer2_outputs(994)) and (layer2_outputs(1746)));
    outputs(1697) <= not((layer2_outputs(1785)) or (layer2_outputs(1796)));
    outputs(1698) <= (layer2_outputs(1933)) and not (layer2_outputs(1241));
    outputs(1699) <= (layer2_outputs(2078)) and not (layer2_outputs(2485));
    outputs(1700) <= layer2_outputs(1860);
    outputs(1701) <= not(layer2_outputs(2460));
    outputs(1702) <= layer2_outputs(1364);
    outputs(1703) <= (layer2_outputs(1426)) and (layer2_outputs(2536));
    outputs(1704) <= layer2_outputs(385);
    outputs(1705) <= layer2_outputs(723);
    outputs(1706) <= not(layer2_outputs(1096));
    outputs(1707) <= not(layer2_outputs(518));
    outputs(1708) <= (layer2_outputs(1125)) and not (layer2_outputs(470));
    outputs(1709) <= not(layer2_outputs(1021));
    outputs(1710) <= not(layer2_outputs(118));
    outputs(1711) <= not(layer2_outputs(703));
    outputs(1712) <= not(layer2_outputs(2173));
    outputs(1713) <= layer2_outputs(172);
    outputs(1714) <= (layer2_outputs(996)) and not (layer2_outputs(80));
    outputs(1715) <= layer2_outputs(696);
    outputs(1716) <= (layer2_outputs(2104)) xor (layer2_outputs(1416));
    outputs(1717) <= not(layer2_outputs(2485));
    outputs(1718) <= not(layer2_outputs(1208));
    outputs(1719) <= (layer2_outputs(1081)) and not (layer2_outputs(1158));
    outputs(1720) <= layer2_outputs(2041);
    outputs(1721) <= not(layer2_outputs(1324)) or (layer2_outputs(2012));
    outputs(1722) <= not((layer2_outputs(2468)) or (layer2_outputs(1108)));
    outputs(1723) <= (layer2_outputs(106)) and not (layer2_outputs(2110));
    outputs(1724) <= not(layer2_outputs(529));
    outputs(1725) <= not(layer2_outputs(1586));
    outputs(1726) <= (layer2_outputs(397)) xor (layer2_outputs(1635));
    outputs(1727) <= not((layer2_outputs(1748)) or (layer2_outputs(207)));
    outputs(1728) <= layer2_outputs(502);
    outputs(1729) <= not((layer2_outputs(2139)) or (layer2_outputs(1583)));
    outputs(1730) <= layer2_outputs(1568);
    outputs(1731) <= not((layer2_outputs(2023)) or (layer2_outputs(1716)));
    outputs(1732) <= not((layer2_outputs(831)) xor (layer2_outputs(23)));
    outputs(1733) <= layer2_outputs(1431);
    outputs(1734) <= (layer2_outputs(1874)) and not (layer2_outputs(1653));
    outputs(1735) <= layer2_outputs(1062);
    outputs(1736) <= (layer2_outputs(805)) and not (layer2_outputs(783));
    outputs(1737) <= layer2_outputs(1560);
    outputs(1738) <= (layer2_outputs(1380)) or (layer2_outputs(448));
    outputs(1739) <= (layer2_outputs(2039)) and not (layer2_outputs(824));
    outputs(1740) <= not(layer2_outputs(886));
    outputs(1741) <= layer2_outputs(1086);
    outputs(1742) <= not(layer2_outputs(1782));
    outputs(1743) <= (layer2_outputs(1546)) and not (layer2_outputs(657));
    outputs(1744) <= (layer2_outputs(2527)) xor (layer2_outputs(2358));
    outputs(1745) <= not(layer2_outputs(2084)) or (layer2_outputs(1486));
    outputs(1746) <= layer2_outputs(979);
    outputs(1747) <= not(layer2_outputs(700));
    outputs(1748) <= layer2_outputs(392);
    outputs(1749) <= not((layer2_outputs(413)) or (layer2_outputs(1270)));
    outputs(1750) <= (layer2_outputs(89)) and not (layer2_outputs(2163));
    outputs(1751) <= not(layer2_outputs(1817));
    outputs(1752) <= (layer2_outputs(250)) and (layer2_outputs(434));
    outputs(1753) <= (layer2_outputs(2142)) and not (layer2_outputs(2259));
    outputs(1754) <= layer2_outputs(424);
    outputs(1755) <= not(layer2_outputs(905));
    outputs(1756) <= layer2_outputs(591);
    outputs(1757) <= not((layer2_outputs(1498)) or (layer2_outputs(1834)));
    outputs(1758) <= not((layer2_outputs(673)) or (layer2_outputs(2030)));
    outputs(1759) <= not((layer2_outputs(398)) or (layer2_outputs(219)));
    outputs(1760) <= not(layer2_outputs(2058)) or (layer2_outputs(448));
    outputs(1761) <= (layer2_outputs(2339)) and not (layer2_outputs(2060));
    outputs(1762) <= not((layer2_outputs(710)) xor (layer2_outputs(1720)));
    outputs(1763) <= not((layer2_outputs(646)) or (layer2_outputs(1606)));
    outputs(1764) <= (layer2_outputs(2351)) and (layer2_outputs(892));
    outputs(1765) <= not(layer2_outputs(1891));
    outputs(1766) <= not(layer2_outputs(1572)) or (layer2_outputs(2425));
    outputs(1767) <= layer2_outputs(2494);
    outputs(1768) <= not((layer2_outputs(1519)) or (layer2_outputs(1549)));
    outputs(1769) <= not((layer2_outputs(807)) or (layer2_outputs(1724)));
    outputs(1770) <= not(layer2_outputs(841));
    outputs(1771) <= (layer2_outputs(1923)) and not (layer2_outputs(105));
    outputs(1772) <= layer2_outputs(360);
    outputs(1773) <= layer2_outputs(295);
    outputs(1774) <= not(layer2_outputs(126));
    outputs(1775) <= not((layer2_outputs(2082)) or (layer2_outputs(1351)));
    outputs(1776) <= layer2_outputs(2338);
    outputs(1777) <= layer2_outputs(1819);
    outputs(1778) <= not(layer2_outputs(1576));
    outputs(1779) <= not(layer2_outputs(1141));
    outputs(1780) <= (layer2_outputs(917)) or (layer2_outputs(917));
    outputs(1781) <= layer2_outputs(1743);
    outputs(1782) <= (layer2_outputs(2356)) xor (layer2_outputs(1349));
    outputs(1783) <= layer2_outputs(1656);
    outputs(1784) <= not(layer2_outputs(1904)) or (layer2_outputs(87));
    outputs(1785) <= layer2_outputs(1987);
    outputs(1786) <= not(layer2_outputs(937));
    outputs(1787) <= not(layer2_outputs(2320));
    outputs(1788) <= not(layer2_outputs(2196));
    outputs(1789) <= not(layer2_outputs(2096));
    outputs(1790) <= not((layer2_outputs(2525)) xor (layer2_outputs(2362)));
    outputs(1791) <= not(layer2_outputs(78));
    outputs(1792) <= not((layer2_outputs(482)) or (layer2_outputs(1157)));
    outputs(1793) <= layer2_outputs(1356);
    outputs(1794) <= not(layer2_outputs(2186));
    outputs(1795) <= layer2_outputs(116);
    outputs(1796) <= (layer2_outputs(2539)) and (layer2_outputs(1908));
    outputs(1797) <= (layer2_outputs(1674)) and not (layer2_outputs(272));
    outputs(1798) <= (layer2_outputs(1118)) or (layer2_outputs(1480));
    outputs(1799) <= (layer2_outputs(395)) and (layer2_outputs(2132));
    outputs(1800) <= not((layer2_outputs(2145)) or (layer2_outputs(553)));
    outputs(1801) <= layer2_outputs(215);
    outputs(1802) <= not(layer2_outputs(451));
    outputs(1803) <= not(layer2_outputs(1706));
    outputs(1804) <= not(layer2_outputs(1365));
    outputs(1805) <= layer2_outputs(1763);
    outputs(1806) <= layer2_outputs(1040);
    outputs(1807) <= layer2_outputs(678);
    outputs(1808) <= not(layer2_outputs(270));
    outputs(1809) <= (layer2_outputs(1437)) and (layer2_outputs(440));
    outputs(1810) <= layer2_outputs(1688);
    outputs(1811) <= not((layer2_outputs(2150)) xor (layer2_outputs(554)));
    outputs(1812) <= (layer2_outputs(635)) and not (layer2_outputs(2407));
    outputs(1813) <= (layer2_outputs(1432)) and not (layer2_outputs(2444));
    outputs(1814) <= layer2_outputs(1837);
    outputs(1815) <= layer2_outputs(2200);
    outputs(1816) <= not(layer2_outputs(1017));
    outputs(1817) <= not(layer2_outputs(1389));
    outputs(1818) <= (layer2_outputs(1077)) and (layer2_outputs(2373));
    outputs(1819) <= not(layer2_outputs(773));
    outputs(1820) <= not(layer2_outputs(930));
    outputs(1821) <= not(layer2_outputs(185));
    outputs(1822) <= not(layer2_outputs(2321));
    outputs(1823) <= (layer2_outputs(1632)) and not (layer2_outputs(101));
    outputs(1824) <= not(layer2_outputs(1413));
    outputs(1825) <= (layer2_outputs(580)) and not (layer2_outputs(1436));
    outputs(1826) <= not((layer2_outputs(2380)) or (layer2_outputs(2374)));
    outputs(1827) <= not(layer2_outputs(2188));
    outputs(1828) <= not(layer2_outputs(1076));
    outputs(1829) <= not(layer2_outputs(1773));
    outputs(1830) <= layer2_outputs(1179);
    outputs(1831) <= layer2_outputs(92);
    outputs(1832) <= (layer2_outputs(201)) and not (layer2_outputs(2177));
    outputs(1833) <= layer2_outputs(126);
    outputs(1834) <= layer2_outputs(2051);
    outputs(1835) <= layer2_outputs(951);
    outputs(1836) <= not(layer2_outputs(1436));
    outputs(1837) <= layer2_outputs(1848);
    outputs(1838) <= not(layer2_outputs(1620));
    outputs(1839) <= (layer2_outputs(2147)) and not (layer2_outputs(1815));
    outputs(1840) <= not((layer2_outputs(957)) or (layer2_outputs(2346)));
    outputs(1841) <= (layer2_outputs(2092)) xor (layer2_outputs(55));
    outputs(1842) <= not((layer2_outputs(351)) or (layer2_outputs(737)));
    outputs(1843) <= not(layer2_outputs(1917));
    outputs(1844) <= not((layer2_outputs(404)) or (layer2_outputs(2461)));
    outputs(1845) <= not((layer2_outputs(1650)) or (layer2_outputs(1245)));
    outputs(1846) <= not((layer2_outputs(1866)) xor (layer2_outputs(2502)));
    outputs(1847) <= layer2_outputs(58);
    outputs(1848) <= not(layer2_outputs(233));
    outputs(1849) <= (layer2_outputs(350)) and not (layer2_outputs(53));
    outputs(1850) <= not(layer2_outputs(2015));
    outputs(1851) <= (layer2_outputs(2309)) and not (layer2_outputs(881));
    outputs(1852) <= (layer2_outputs(1345)) and not (layer2_outputs(826));
    outputs(1853) <= not(layer2_outputs(1455));
    outputs(1854) <= not((layer2_outputs(2099)) xor (layer2_outputs(1043)));
    outputs(1855) <= (layer2_outputs(114)) and (layer2_outputs(561));
    outputs(1856) <= layer2_outputs(155);
    outputs(1857) <= not(layer2_outputs(1091)) or (layer2_outputs(94));
    outputs(1858) <= layer2_outputs(2308);
    outputs(1859) <= (layer2_outputs(1108)) and not (layer2_outputs(2106));
    outputs(1860) <= layer2_outputs(1491);
    outputs(1861) <= not((layer2_outputs(623)) or (layer2_outputs(2141)));
    outputs(1862) <= not(layer2_outputs(547));
    outputs(1863) <= not((layer2_outputs(1387)) or (layer2_outputs(409)));
    outputs(1864) <= not(layer2_outputs(1899));
    outputs(1865) <= not(layer2_outputs(313));
    outputs(1866) <= (layer2_outputs(9)) and not (layer2_outputs(2266));
    outputs(1867) <= (layer2_outputs(1854)) and not (layer2_outputs(1587));
    outputs(1868) <= layer2_outputs(1296);
    outputs(1869) <= layer2_outputs(532);
    outputs(1870) <= (layer2_outputs(188)) xor (layer2_outputs(403));
    outputs(1871) <= layer2_outputs(1148);
    outputs(1872) <= not((layer2_outputs(369)) or (layer2_outputs(345)));
    outputs(1873) <= (layer2_outputs(2558)) and not (layer2_outputs(1892));
    outputs(1874) <= layer2_outputs(1393);
    outputs(1875) <= (layer2_outputs(541)) and (layer2_outputs(1055));
    outputs(1876) <= layer2_outputs(1309);
    outputs(1877) <= not(layer2_outputs(1865));
    outputs(1878) <= (layer2_outputs(1281)) and (layer2_outputs(7));
    outputs(1879) <= not(layer2_outputs(1555));
    outputs(1880) <= not(layer2_outputs(437));
    outputs(1881) <= layer2_outputs(49);
    outputs(1882) <= layer2_outputs(258);
    outputs(1883) <= (layer2_outputs(1982)) xor (layer2_outputs(2095));
    outputs(1884) <= not(layer2_outputs(2515));
    outputs(1885) <= layer2_outputs(1003);
    outputs(1886) <= not((layer2_outputs(886)) or (layer2_outputs(0)));
    outputs(1887) <= not(layer2_outputs(125));
    outputs(1888) <= layer2_outputs(1982);
    outputs(1889) <= layer2_outputs(1034);
    outputs(1890) <= layer2_outputs(352);
    outputs(1891) <= layer2_outputs(417);
    outputs(1892) <= (layer2_outputs(1107)) and (layer2_outputs(311));
    outputs(1893) <= not(layer2_outputs(1219));
    outputs(1894) <= not(layer2_outputs(941));
    outputs(1895) <= (layer2_outputs(2468)) or (layer2_outputs(1885));
    outputs(1896) <= not(layer2_outputs(364));
    outputs(1897) <= layer2_outputs(2001);
    outputs(1898) <= layer2_outputs(1717);
    outputs(1899) <= not(layer2_outputs(1328));
    outputs(1900) <= layer2_outputs(367);
    outputs(1901) <= (layer2_outputs(2284)) and not (layer2_outputs(1928));
    outputs(1902) <= not((layer2_outputs(314)) or (layer2_outputs(1030)));
    outputs(1903) <= (layer2_outputs(1777)) and not (layer2_outputs(339));
    outputs(1904) <= (layer2_outputs(484)) and not (layer2_outputs(827));
    outputs(1905) <= (layer2_outputs(1498)) and (layer2_outputs(839));
    outputs(1906) <= not(layer2_outputs(542));
    outputs(1907) <= not(layer2_outputs(982));
    outputs(1908) <= not((layer2_outputs(1772)) or (layer2_outputs(383)));
    outputs(1909) <= not((layer2_outputs(1440)) xor (layer2_outputs(729)));
    outputs(1910) <= layer2_outputs(774);
    outputs(1911) <= not(layer2_outputs(2176));
    outputs(1912) <= (layer2_outputs(1393)) and (layer2_outputs(816));
    outputs(1913) <= not((layer2_outputs(1582)) or (layer2_outputs(1660)));
    outputs(1914) <= not(layer2_outputs(291));
    outputs(1915) <= layer2_outputs(2357);
    outputs(1916) <= not(layer2_outputs(941));
    outputs(1917) <= (layer2_outputs(1980)) and (layer2_outputs(74));
    outputs(1918) <= (layer2_outputs(1648)) and (layer2_outputs(1741));
    outputs(1919) <= not(layer2_outputs(2017));
    outputs(1920) <= (layer2_outputs(1376)) and not (layer2_outputs(758));
    outputs(1921) <= not(layer2_outputs(1031));
    outputs(1922) <= layer2_outputs(1842);
    outputs(1923) <= not(layer2_outputs(1159));
    outputs(1924) <= not(layer2_outputs(1094));
    outputs(1925) <= layer2_outputs(63);
    outputs(1926) <= (layer2_outputs(149)) and not (layer2_outputs(1570));
    outputs(1927) <= (layer2_outputs(2072)) and not (layer2_outputs(108));
    outputs(1928) <= not(layer2_outputs(1966));
    outputs(1929) <= (layer2_outputs(1689)) and not (layer2_outputs(2090));
    outputs(1930) <= not((layer2_outputs(1286)) or (layer2_outputs(10)));
    outputs(1931) <= not(layer2_outputs(2097));
    outputs(1932) <= layer2_outputs(1358);
    outputs(1933) <= (layer2_outputs(766)) and not (layer2_outputs(151));
    outputs(1934) <= (layer2_outputs(714)) xor (layer2_outputs(1324));
    outputs(1935) <= not((layer2_outputs(60)) xor (layer2_outputs(2251)));
    outputs(1936) <= not((layer2_outputs(950)) or (layer2_outputs(144)));
    outputs(1937) <= not(layer2_outputs(133));
    outputs(1938) <= layer2_outputs(1846);
    outputs(1939) <= (layer2_outputs(1258)) and not (layer2_outputs(1755));
    outputs(1940) <= layer2_outputs(1462);
    outputs(1941) <= layer2_outputs(246);
    outputs(1942) <= layer2_outputs(428);
    outputs(1943) <= not(layer2_outputs(2316)) or (layer2_outputs(1414));
    outputs(1944) <= (layer2_outputs(378)) or (layer2_outputs(290));
    outputs(1945) <= (layer2_outputs(2087)) xor (layer2_outputs(819));
    outputs(1946) <= (layer2_outputs(354)) and not (layer2_outputs(1193));
    outputs(1947) <= not(layer2_outputs(476));
    outputs(1948) <= layer2_outputs(178);
    outputs(1949) <= layer2_outputs(1716);
    outputs(1950) <= layer2_outputs(60);
    outputs(1951) <= layer2_outputs(2462);
    outputs(1952) <= (layer2_outputs(2244)) and (layer2_outputs(762));
    outputs(1953) <= not((layer2_outputs(236)) or (layer2_outputs(1120)));
    outputs(1954) <= layer2_outputs(1035);
    outputs(1955) <= not(layer2_outputs(353));
    outputs(1956) <= not(layer2_outputs(2183));
    outputs(1957) <= (layer2_outputs(1080)) and not (layer2_outputs(2261));
    outputs(1958) <= layer2_outputs(2395);
    outputs(1959) <= layer2_outputs(1915);
    outputs(1960) <= not(layer2_outputs(415));
    outputs(1961) <= layer2_outputs(2100);
    outputs(1962) <= layer2_outputs(554);
    outputs(1963) <= not(layer2_outputs(697));
    outputs(1964) <= layer2_outputs(1908);
    outputs(1965) <= not((layer2_outputs(305)) or (layer2_outputs(187)));
    outputs(1966) <= not((layer2_outputs(1420)) xor (layer2_outputs(1628)));
    outputs(1967) <= (layer2_outputs(137)) and (layer2_outputs(2252));
    outputs(1968) <= (layer2_outputs(1668)) and not (layer2_outputs(1184));
    outputs(1969) <= layer2_outputs(2344);
    outputs(1970) <= not(layer2_outputs(1137));
    outputs(1971) <= (layer2_outputs(954)) and not (layer2_outputs(291));
    outputs(1972) <= (layer2_outputs(839)) and not (layer2_outputs(1185));
    outputs(1973) <= (layer2_outputs(478)) or (layer2_outputs(2476));
    outputs(1974) <= not(layer2_outputs(1808));
    outputs(1975) <= layer2_outputs(2383);
    outputs(1976) <= not(layer2_outputs(2393));
    outputs(1977) <= (layer2_outputs(2519)) and (layer2_outputs(40));
    outputs(1978) <= (layer2_outputs(550)) and not (layer2_outputs(1166));
    outputs(1979) <= not(layer2_outputs(1692));
    outputs(1980) <= not(layer2_outputs(2423));
    outputs(1981) <= not(layer2_outputs(2055));
    outputs(1982) <= not((layer2_outputs(1990)) and (layer2_outputs(2422)));
    outputs(1983) <= not(layer2_outputs(176));
    outputs(1984) <= layer2_outputs(1357);
    outputs(1985) <= not(layer2_outputs(1881));
    outputs(1986) <= (layer2_outputs(2227)) and not (layer2_outputs(1383));
    outputs(1987) <= (layer2_outputs(329)) and not (layer2_outputs(6));
    outputs(1988) <= not(layer2_outputs(545));
    outputs(1989) <= (layer2_outputs(659)) and not (layer2_outputs(2428));
    outputs(1990) <= layer2_outputs(444);
    outputs(1991) <= not(layer2_outputs(129));
    outputs(1992) <= layer2_outputs(2198);
    outputs(1993) <= not(layer2_outputs(684));
    outputs(1994) <= (layer2_outputs(1648)) and not (layer2_outputs(200));
    outputs(1995) <= (layer2_outputs(1594)) and (layer2_outputs(218));
    outputs(1996) <= layer2_outputs(1591);
    outputs(1997) <= (layer2_outputs(567)) and (layer2_outputs(1516));
    outputs(1998) <= not(layer2_outputs(1029));
    outputs(1999) <= not(layer2_outputs(62));
    outputs(2000) <= layer2_outputs(349);
    outputs(2001) <= layer2_outputs(2470);
    outputs(2002) <= layer2_outputs(1504);
    outputs(2003) <= (layer2_outputs(1538)) and not (layer2_outputs(915));
    outputs(2004) <= not(layer2_outputs(1823));
    outputs(2005) <= layer2_outputs(759);
    outputs(2006) <= not((layer2_outputs(232)) or (layer2_outputs(1130)));
    outputs(2007) <= not((layer2_outputs(493)) or (layer2_outputs(862)));
    outputs(2008) <= (layer2_outputs(551)) and (layer2_outputs(1066));
    outputs(2009) <= not(layer2_outputs(2285));
    outputs(2010) <= (layer2_outputs(2269)) and not (layer2_outputs(546));
    outputs(2011) <= (layer2_outputs(627)) and not (layer2_outputs(1136));
    outputs(2012) <= layer2_outputs(104);
    outputs(2013) <= not(layer2_outputs(1729));
    outputs(2014) <= not(layer2_outputs(592));
    outputs(2015) <= layer2_outputs(1611);
    outputs(2016) <= layer2_outputs(2084);
    outputs(2017) <= not(layer2_outputs(617)) or (layer2_outputs(2064));
    outputs(2018) <= (layer2_outputs(1090)) and not (layer2_outputs(193));
    outputs(2019) <= layer2_outputs(2437);
    outputs(2020) <= (layer2_outputs(2215)) and not (layer2_outputs(2180));
    outputs(2021) <= (layer2_outputs(610)) and (layer2_outputs(197));
    outputs(2022) <= not(layer2_outputs(2298));
    outputs(2023) <= layer2_outputs(2114);
    outputs(2024) <= not(layer2_outputs(1087));
    outputs(2025) <= not(layer2_outputs(843));
    outputs(2026) <= not(layer2_outputs(2454)) or (layer2_outputs(322));
    outputs(2027) <= (layer2_outputs(1764)) and not (layer2_outputs(1338));
    outputs(2028) <= (layer2_outputs(419)) and not (layer2_outputs(1827));
    outputs(2029) <= (layer2_outputs(2051)) and (layer2_outputs(762));
    outputs(2030) <= (layer2_outputs(2289)) and (layer2_outputs(1709));
    outputs(2031) <= not((layer2_outputs(206)) and (layer2_outputs(667)));
    outputs(2032) <= not(layer2_outputs(236));
    outputs(2033) <= (layer2_outputs(1148)) and not (layer2_outputs(2296));
    outputs(2034) <= layer2_outputs(2225);
    outputs(2035) <= (layer2_outputs(1989)) or (layer2_outputs(820));
    outputs(2036) <= not(layer2_outputs(1973));
    outputs(2037) <= (layer2_outputs(1036)) and (layer2_outputs(444));
    outputs(2038) <= layer2_outputs(1381);
    outputs(2039) <= (layer2_outputs(2499)) and (layer2_outputs(153));
    outputs(2040) <= (layer2_outputs(1346)) or (layer2_outputs(1735));
    outputs(2041) <= not(layer2_outputs(1605));
    outputs(2042) <= not(layer2_outputs(1812));
    outputs(2043) <= (layer2_outputs(2237)) and (layer2_outputs(887));
    outputs(2044) <= not(layer2_outputs(2418));
    outputs(2045) <= not(layer2_outputs(2014));
    outputs(2046) <= not(layer2_outputs(2279));
    outputs(2047) <= (layer2_outputs(67)) and not (layer2_outputs(1971));
    outputs(2048) <= not(layer2_outputs(1437));
    outputs(2049) <= layer2_outputs(1032);
    outputs(2050) <= not(layer2_outputs(2003));
    outputs(2051) <= not(layer2_outputs(738));
    outputs(2052) <= (layer2_outputs(1709)) and not (layer2_outputs(481));
    outputs(2053) <= not(layer2_outputs(1319));
    outputs(2054) <= layer2_outputs(1681);
    outputs(2055) <= layer2_outputs(1117);
    outputs(2056) <= not((layer2_outputs(2433)) xor (layer2_outputs(1682)));
    outputs(2057) <= not(layer2_outputs(649));
    outputs(2058) <= (layer2_outputs(299)) xor (layer2_outputs(1006));
    outputs(2059) <= layer2_outputs(230);
    outputs(2060) <= layer2_outputs(747);
    outputs(2061) <= not(layer2_outputs(2494));
    outputs(2062) <= not(layer2_outputs(794));
    outputs(2063) <= not(layer2_outputs(1619));
    outputs(2064) <= not(layer2_outputs(721));
    outputs(2065) <= not(layer2_outputs(340)) or (layer2_outputs(1813));
    outputs(2066) <= (layer2_outputs(2213)) xor (layer2_outputs(198));
    outputs(2067) <= layer2_outputs(197);
    outputs(2068) <= not((layer2_outputs(418)) and (layer2_outputs(710)));
    outputs(2069) <= layer2_outputs(687);
    outputs(2070) <= not(layer2_outputs(590)) or (layer2_outputs(2322));
    outputs(2071) <= not(layer2_outputs(1321)) or (layer2_outputs(543));
    outputs(2072) <= not(layer2_outputs(484));
    outputs(2073) <= (layer2_outputs(642)) and (layer2_outputs(1423));
    outputs(2074) <= layer2_outputs(184);
    outputs(2075) <= not(layer2_outputs(237));
    outputs(2076) <= not(layer2_outputs(399));
    outputs(2077) <= not(layer2_outputs(2458));
    outputs(2078) <= not(layer2_outputs(1931));
    outputs(2079) <= not(layer2_outputs(2408));
    outputs(2080) <= layer2_outputs(602);
    outputs(2081) <= layer2_outputs(2228);
    outputs(2082) <= (layer2_outputs(426)) xor (layer2_outputs(500));
    outputs(2083) <= not(layer2_outputs(373));
    outputs(2084) <= layer2_outputs(2327);
    outputs(2085) <= not((layer2_outputs(1793)) xor (layer2_outputs(552)));
    outputs(2086) <= not((layer2_outputs(1651)) and (layer2_outputs(691)));
    outputs(2087) <= (layer2_outputs(1054)) or (layer2_outputs(1349));
    outputs(2088) <= not(layer2_outputs(1531));
    outputs(2089) <= (layer2_outputs(1601)) and (layer2_outputs(2120));
    outputs(2090) <= not(layer2_outputs(334));
    outputs(2091) <= layer2_outputs(307);
    outputs(2092) <= not(layer2_outputs(139)) or (layer2_outputs(1));
    outputs(2093) <= not(layer2_outputs(513));
    outputs(2094) <= layer2_outputs(897);
    outputs(2095) <= (layer2_outputs(2402)) xor (layer2_outputs(683));
    outputs(2096) <= not(layer2_outputs(1186));
    outputs(2097) <= (layer2_outputs(845)) and (layer2_outputs(1098));
    outputs(2098) <= not(layer2_outputs(772));
    outputs(2099) <= not((layer2_outputs(2074)) or (layer2_outputs(190)));
    outputs(2100) <= not(layer2_outputs(1220));
    outputs(2101) <= not((layer2_outputs(1442)) and (layer2_outputs(555)));
    outputs(2102) <= not((layer2_outputs(372)) or (layer2_outputs(1405)));
    outputs(2103) <= layer2_outputs(488);
    outputs(2104) <= layer2_outputs(58);
    outputs(2105) <= not(layer2_outputs(2124));
    outputs(2106) <= layer2_outputs(1646);
    outputs(2107) <= not(layer2_outputs(1404));
    outputs(2108) <= not(layer2_outputs(1619));
    outputs(2109) <= (layer2_outputs(1357)) or (layer2_outputs(189));
    outputs(2110) <= not((layer2_outputs(2410)) xor (layer2_outputs(1103)));
    outputs(2111) <= not((layer2_outputs(2291)) and (layer2_outputs(2186)));
    outputs(2112) <= not(layer2_outputs(2152));
    outputs(2113) <= not(layer2_outputs(2325));
    outputs(2114) <= layer2_outputs(944);
    outputs(2115) <= layer2_outputs(1661);
    outputs(2116) <= (layer2_outputs(435)) and not (layer2_outputs(802));
    outputs(2117) <= not(layer2_outputs(1658));
    outputs(2118) <= layer2_outputs(1409);
    outputs(2119) <= not(layer2_outputs(367));
    outputs(2120) <= not(layer2_outputs(864));
    outputs(2121) <= (layer2_outputs(1240)) xor (layer2_outputs(1496));
    outputs(2122) <= not(layer2_outputs(2140));
    outputs(2123) <= (layer2_outputs(644)) xor (layer2_outputs(2287));
    outputs(2124) <= not(layer2_outputs(499));
    outputs(2125) <= not(layer2_outputs(2533)) or (layer2_outputs(695));
    outputs(2126) <= layer2_outputs(2340);
    outputs(2127) <= not((layer2_outputs(1666)) xor (layer2_outputs(787)));
    outputs(2128) <= not(layer2_outputs(663));
    outputs(2129) <= not(layer2_outputs(328));
    outputs(2130) <= layer2_outputs(1244);
    outputs(2131) <= layer2_outputs(2113);
    outputs(2132) <= (layer2_outputs(1292)) xor (layer2_outputs(1630));
    outputs(2133) <= layer2_outputs(1138);
    outputs(2134) <= (layer2_outputs(652)) xor (layer2_outputs(1067));
    outputs(2135) <= (layer2_outputs(2362)) xor (layer2_outputs(633));
    outputs(2136) <= not(layer2_outputs(2028));
    outputs(2137) <= not(layer2_outputs(1306));
    outputs(2138) <= layer2_outputs(2425);
    outputs(2139) <= not(layer2_outputs(1101));
    outputs(2140) <= (layer2_outputs(2457)) xor (layer2_outputs(2387));
    outputs(2141) <= (layer2_outputs(1928)) and not (layer2_outputs(1173));
    outputs(2142) <= not(layer2_outputs(57));
    outputs(2143) <= layer2_outputs(2097);
    outputs(2144) <= layer2_outputs(1469);
    outputs(2145) <= layer2_outputs(2290);
    outputs(2146) <= layer2_outputs(1180);
    outputs(2147) <= layer2_outputs(1146);
    outputs(2148) <= layer2_outputs(925);
    outputs(2149) <= (layer2_outputs(1935)) and not (layer2_outputs(2070));
    outputs(2150) <= layer2_outputs(2177);
    outputs(2151) <= not(layer2_outputs(1259));
    outputs(2152) <= layer2_outputs(2250);
    outputs(2153) <= layer2_outputs(1169);
    outputs(2154) <= not(layer2_outputs(56)) or (layer2_outputs(1829));
    outputs(2155) <= not((layer2_outputs(1670)) or (layer2_outputs(513)));
    outputs(2156) <= (layer2_outputs(1602)) xor (layer2_outputs(2066));
    outputs(2157) <= not(layer2_outputs(2541));
    outputs(2158) <= layer2_outputs(1420);
    outputs(2159) <= not(layer2_outputs(1828));
    outputs(2160) <= not((layer2_outputs(1621)) xor (layer2_outputs(450)));
    outputs(2161) <= not(layer2_outputs(124));
    outputs(2162) <= (layer2_outputs(977)) and not (layer2_outputs(169));
    outputs(2163) <= layer2_outputs(1729);
    outputs(2164) <= not(layer2_outputs(216));
    outputs(2165) <= not(layer2_outputs(1604)) or (layer2_outputs(576));
    outputs(2166) <= (layer2_outputs(1484)) or (layer2_outputs(1846));
    outputs(2167) <= not(layer2_outputs(2124));
    outputs(2168) <= not(layer2_outputs(2403));
    outputs(2169) <= not((layer2_outputs(11)) xor (layer2_outputs(369)));
    outputs(2170) <= not((layer2_outputs(945)) and (layer2_outputs(2328)));
    outputs(2171) <= not((layer2_outputs(1197)) or (layer2_outputs(1097)));
    outputs(2172) <= not(layer2_outputs(1574));
    outputs(2173) <= not(layer2_outputs(1400)) or (layer2_outputs(1262));
    outputs(2174) <= not(layer2_outputs(464));
    outputs(2175) <= not((layer2_outputs(1025)) or (layer2_outputs(2266)));
    outputs(2176) <= layer2_outputs(2515);
    outputs(2177) <= layer2_outputs(548);
    outputs(2178) <= layer2_outputs(229);
    outputs(2179) <= not(layer2_outputs(1804));
    outputs(2180) <= not(layer2_outputs(363));
    outputs(2181) <= layer2_outputs(1967);
    outputs(2182) <= not(layer2_outputs(905));
    outputs(2183) <= not(layer2_outputs(2532));
    outputs(2184) <= not(layer2_outputs(1273));
    outputs(2185) <= not(layer2_outputs(779));
    outputs(2186) <= layer2_outputs(449);
    outputs(2187) <= (layer2_outputs(1999)) and not (layer2_outputs(1059));
    outputs(2188) <= layer2_outputs(2203);
    outputs(2189) <= layer2_outputs(2478);
    outputs(2190) <= not(layer2_outputs(664)) or (layer2_outputs(1098));
    outputs(2191) <= not(layer2_outputs(1920));
    outputs(2192) <= layer2_outputs(1144);
    outputs(2193) <= not(layer2_outputs(1885));
    outputs(2194) <= (layer2_outputs(486)) xor (layer2_outputs(767));
    outputs(2195) <= layer2_outputs(609);
    outputs(2196) <= (layer2_outputs(2277)) and not (layer2_outputs(504));
    outputs(2197) <= layer2_outputs(2327);
    outputs(2198) <= layer2_outputs(1372);
    outputs(2199) <= (layer2_outputs(564)) and not (layer2_outputs(712));
    outputs(2200) <= not(layer2_outputs(2345));
    outputs(2201) <= not(layer2_outputs(502));
    outputs(2202) <= not(layer2_outputs(159));
    outputs(2203) <= not(layer2_outputs(1320));
    outputs(2204) <= layer2_outputs(2535);
    outputs(2205) <= not(layer2_outputs(1748));
    outputs(2206) <= (layer2_outputs(2283)) xor (layer2_outputs(725));
    outputs(2207) <= (layer2_outputs(619)) and not (layer2_outputs(641));
    outputs(2208) <= not((layer2_outputs(2482)) xor (layer2_outputs(2)));
    outputs(2209) <= (layer2_outputs(28)) xor (layer2_outputs(2506));
    outputs(2210) <= layer2_outputs(1654);
    outputs(2211) <= layer2_outputs(462);
    outputs(2212) <= not(layer2_outputs(1124));
    outputs(2213) <= (layer2_outputs(397)) xor (layer2_outputs(821));
    outputs(2214) <= not(layer2_outputs(1740));
    outputs(2215) <= (layer2_outputs(840)) xor (layer2_outputs(2470));
    outputs(2216) <= not(layer2_outputs(990));
    outputs(2217) <= layer2_outputs(25);
    outputs(2218) <= (layer2_outputs(2552)) or (layer2_outputs(244));
    outputs(2219) <= (layer2_outputs(1010)) xor (layer2_outputs(954));
    outputs(2220) <= not(layer2_outputs(2386));
    outputs(2221) <= layer2_outputs(430);
    outputs(2222) <= layer2_outputs(1200);
    outputs(2223) <= (layer2_outputs(1858)) and (layer2_outputs(391));
    outputs(2224) <= not(layer2_outputs(329));
    outputs(2225) <= (layer2_outputs(735)) or (layer2_outputs(467));
    outputs(2226) <= (layer2_outputs(872)) xor (layer2_outputs(629));
    outputs(2227) <= layer2_outputs(1643);
    outputs(2228) <= not(layer2_outputs(675));
    outputs(2229) <= not(layer2_outputs(1833));
    outputs(2230) <= not(layer2_outputs(2138));
    outputs(2231) <= layer2_outputs(37);
    outputs(2232) <= (layer2_outputs(1078)) xor (layer2_outputs(490));
    outputs(2233) <= (layer2_outputs(984)) and not (layer2_outputs(713));
    outputs(2234) <= not(layer2_outputs(612)) or (layer2_outputs(1864));
    outputs(2235) <= (layer2_outputs(2281)) or (layer2_outputs(1167));
    outputs(2236) <= (layer2_outputs(2394)) xor (layer2_outputs(1938));
    outputs(2237) <= (layer2_outputs(1674)) and not (layer2_outputs(93));
    outputs(2238) <= (layer2_outputs(1873)) and not (layer2_outputs(736));
    outputs(2239) <= layer2_outputs(1930);
    outputs(2240) <= (layer2_outputs(1231)) and (layer2_outputs(2160));
    outputs(2241) <= layer2_outputs(1057);
    outputs(2242) <= layer2_outputs(1549);
    outputs(2243) <= layer2_outputs(1190);
    outputs(2244) <= (layer2_outputs(412)) xor (layer2_outputs(1266));
    outputs(2245) <= not((layer2_outputs(2010)) xor (layer2_outputs(1678)));
    outputs(2246) <= (layer2_outputs(225)) and (layer2_outputs(110));
    outputs(2247) <= not(layer2_outputs(2315));
    outputs(2248) <= layer2_outputs(2336);
    outputs(2249) <= layer2_outputs(1698);
    outputs(2250) <= not(layer2_outputs(607));
    outputs(2251) <= layer2_outputs(918);
    outputs(2252) <= layer2_outputs(102);
    outputs(2253) <= not(layer2_outputs(1405));
    outputs(2254) <= not(layer2_outputs(420));
    outputs(2255) <= (layer2_outputs(1039)) or (layer2_outputs(1138));
    outputs(2256) <= layer2_outputs(631);
    outputs(2257) <= (layer2_outputs(1818)) and (layer2_outputs(1439));
    outputs(2258) <= (layer2_outputs(591)) or (layer2_outputs(830));
    outputs(2259) <= not(layer2_outputs(2098));
    outputs(2260) <= not(layer2_outputs(746));
    outputs(2261) <= layer2_outputs(1180);
    outputs(2262) <= (layer2_outputs(919)) and not (layer2_outputs(2232));
    outputs(2263) <= layer2_outputs(1117);
    outputs(2264) <= layer2_outputs(1002);
    outputs(2265) <= layer2_outputs(81);
    outputs(2266) <= (layer2_outputs(2497)) and (layer2_outputs(973));
    outputs(2267) <= not(layer2_outputs(2073));
    outputs(2268) <= layer2_outputs(1424);
    outputs(2269) <= not(layer2_outputs(1719));
    outputs(2270) <= layer2_outputs(1680);
    outputs(2271) <= layer2_outputs(1347);
    outputs(2272) <= layer2_outputs(1633);
    outputs(2273) <= not((layer2_outputs(552)) xor (layer2_outputs(2511)));
    outputs(2274) <= not(layer2_outputs(842));
    outputs(2275) <= not(layer2_outputs(1579)) or (layer2_outputs(1998));
    outputs(2276) <= layer2_outputs(2252);
    outputs(2277) <= (layer2_outputs(441)) and (layer2_outputs(321));
    outputs(2278) <= layer2_outputs(1372);
    outputs(2279) <= (layer2_outputs(1041)) or (layer2_outputs(998));
    outputs(2280) <= (layer2_outputs(2247)) or (layer2_outputs(173));
    outputs(2281) <= not(layer2_outputs(190));
    outputs(2282) <= layer2_outputs(1473);
    outputs(2283) <= not(layer2_outputs(117));
    outputs(2284) <= not((layer2_outputs(1540)) xor (layer2_outputs(2270)));
    outputs(2285) <= not(layer2_outputs(399));
    outputs(2286) <= layer2_outputs(1601);
    outputs(2287) <= (layer2_outputs(2263)) and (layer2_outputs(1609));
    outputs(2288) <= layer2_outputs(1728);
    outputs(2289) <= (layer2_outputs(2020)) and not (layer2_outputs(1336));
    outputs(2290) <= layer2_outputs(44);
    outputs(2291) <= layer2_outputs(1463);
    outputs(2292) <= layer2_outputs(344);
    outputs(2293) <= layer2_outputs(391);
    outputs(2294) <= layer2_outputs(1505);
    outputs(2295) <= not(layer2_outputs(2337)) or (layer2_outputs(969));
    outputs(2296) <= not(layer2_outputs(2070));
    outputs(2297) <= layer2_outputs(2528);
    outputs(2298) <= layer2_outputs(2391);
    outputs(2299) <= not(layer2_outputs(2205));
    outputs(2300) <= not(layer2_outputs(545)) or (layer2_outputs(2513));
    outputs(2301) <= not(layer2_outputs(128)) or (layer2_outputs(875));
    outputs(2302) <= not((layer2_outputs(1767)) or (layer2_outputs(656)));
    outputs(2303) <= not(layer2_outputs(1211));
    outputs(2304) <= (layer2_outputs(1014)) and (layer2_outputs(1664));
    outputs(2305) <= not(layer2_outputs(1760));
    outputs(2306) <= not(layer2_outputs(1044));
    outputs(2307) <= not((layer2_outputs(632)) or (layer2_outputs(1056)));
    outputs(2308) <= (layer2_outputs(2369)) and not (layer2_outputs(1387));
    outputs(2309) <= (layer2_outputs(1863)) and not (layer2_outputs(861));
    outputs(2310) <= not(layer2_outputs(108));
    outputs(2311) <= not((layer2_outputs(2293)) or (layer2_outputs(1726)));
    outputs(2312) <= layer2_outputs(1511);
    outputs(2313) <= not((layer2_outputs(2540)) or (layer2_outputs(243)));
    outputs(2314) <= not(layer2_outputs(1492));
    outputs(2315) <= (layer2_outputs(121)) xor (layer2_outputs(1509));
    outputs(2316) <= (layer2_outputs(1073)) xor (layer2_outputs(30));
    outputs(2317) <= not((layer2_outputs(926)) and (layer2_outputs(1215)));
    outputs(2318) <= not(layer2_outputs(1794));
    outputs(2319) <= layer2_outputs(201);
    outputs(2320) <= not(layer2_outputs(1865));
    outputs(2321) <= not(layer2_outputs(1430));
    outputs(2322) <= layer2_outputs(1021);
    outputs(2323) <= layer2_outputs(1444);
    outputs(2324) <= not(layer2_outputs(658));
    outputs(2325) <= layer2_outputs(211);
    outputs(2326) <= not(layer2_outputs(637));
    outputs(2327) <= not(layer2_outputs(1012));
    outputs(2328) <= layer2_outputs(1281);
    outputs(2329) <= not(layer2_outputs(287));
    outputs(2330) <= layer2_outputs(583);
    outputs(2331) <= (layer2_outputs(1452)) and not (layer2_outputs(2414));
    outputs(2332) <= not(layer2_outputs(2418));
    outputs(2333) <= not(layer2_outputs(1228));
    outputs(2334) <= layer2_outputs(2230);
    outputs(2335) <= not((layer2_outputs(2050)) and (layer2_outputs(1006)));
    outputs(2336) <= not(layer2_outputs(1118));
    outputs(2337) <= (layer2_outputs(529)) and not (layer2_outputs(1585));
    outputs(2338) <= (layer2_outputs(1007)) and not (layer2_outputs(2508));
    outputs(2339) <= not(layer2_outputs(856)) or (layer2_outputs(1412));
    outputs(2340) <= layer2_outputs(947);
    outputs(2341) <= layer2_outputs(86);
    outputs(2342) <= layer2_outputs(1233);
    outputs(2343) <= (layer2_outputs(586)) and (layer2_outputs(1792));
    outputs(2344) <= not(layer2_outputs(287));
    outputs(2345) <= not(layer2_outputs(1832));
    outputs(2346) <= (layer2_outputs(1525)) and not (layer2_outputs(191));
    outputs(2347) <= layer2_outputs(1861);
    outputs(2348) <= (layer2_outputs(2302)) and (layer2_outputs(2475));
    outputs(2349) <= (layer2_outputs(95)) and not (layer2_outputs(1679));
    outputs(2350) <= not(layer2_outputs(1542));
    outputs(2351) <= not((layer2_outputs(1783)) and (layer2_outputs(166)));
    outputs(2352) <= not(layer2_outputs(1175)) or (layer2_outputs(1079));
    outputs(2353) <= layer2_outputs(970);
    outputs(2354) <= not(layer2_outputs(2217));
    outputs(2355) <= layer2_outputs(2009);
    outputs(2356) <= (layer2_outputs(558)) and not (layer2_outputs(2045));
    outputs(2357) <= not((layer2_outputs(1358)) or (layer2_outputs(2355)));
    outputs(2358) <= layer2_outputs(1481);
    outputs(2359) <= layer2_outputs(496);
    outputs(2360) <= layer2_outputs(1111);
    outputs(2361) <= layer2_outputs(1205);
    outputs(2362) <= layer2_outputs(2556);
    outputs(2363) <= not(layer2_outputs(208));
    outputs(2364) <= not(layer2_outputs(974));
    outputs(2365) <= layer2_outputs(1608);
    outputs(2366) <= (layer2_outputs(2062)) and not (layer2_outputs(1119));
    outputs(2367) <= layer2_outputs(1330);
    outputs(2368) <= layer2_outputs(440);
    outputs(2369) <= (layer2_outputs(308)) xor (layer2_outputs(994));
    outputs(2370) <= not(layer2_outputs(2333));
    outputs(2371) <= layer2_outputs(2080);
    outputs(2372) <= (layer2_outputs(1027)) and (layer2_outputs(1050));
    outputs(2373) <= not((layer2_outputs(132)) xor (layer2_outputs(2492)));
    outputs(2374) <= not(layer2_outputs(699));
    outputs(2375) <= not((layer2_outputs(688)) xor (layer2_outputs(2372)));
    outputs(2376) <= layer2_outputs(463);
    outputs(2377) <= not(layer2_outputs(1898));
    outputs(2378) <= not(layer2_outputs(1879));
    outputs(2379) <= not(layer2_outputs(1457));
    outputs(2380) <= not((layer2_outputs(2001)) or (layer2_outputs(537)));
    outputs(2381) <= not(layer2_outputs(1199));
    outputs(2382) <= not((layer2_outputs(2528)) or (layer2_outputs(2489)));
    outputs(2383) <= layer2_outputs(2152);
    outputs(2384) <= layer2_outputs(1160);
    outputs(2385) <= not(layer2_outputs(2335));
    outputs(2386) <= not(layer2_outputs(2210)) or (layer2_outputs(1610));
    outputs(2387) <= not(layer2_outputs(763));
    outputs(2388) <= (layer2_outputs(533)) and not (layer2_outputs(2409));
    outputs(2389) <= layer2_outputs(2121);
    outputs(2390) <= not((layer2_outputs(2551)) or (layer2_outputs(240)));
    outputs(2391) <= (layer2_outputs(1675)) and (layer2_outputs(769));
    outputs(2392) <= (layer2_outputs(1038)) and (layer2_outputs(613));
    outputs(2393) <= (layer2_outputs(1001)) and not (layer2_outputs(13));
    outputs(2394) <= layer2_outputs(1588);
    outputs(2395) <= not(layer2_outputs(2321));
    outputs(2396) <= layer2_outputs(2472);
    outputs(2397) <= layer2_outputs(178);
    outputs(2398) <= not(layer2_outputs(1501));
    outputs(2399) <= layer2_outputs(1176);
    outputs(2400) <= not(layer2_outputs(2315));
    outputs(2401) <= layer2_outputs(1187);
    outputs(2402) <= (layer2_outputs(1612)) xor (layer2_outputs(2243));
    outputs(2403) <= layer2_outputs(1176);
    outputs(2404) <= layer2_outputs(1267);
    outputs(2405) <= (layer2_outputs(2222)) and not (layer2_outputs(1669));
    outputs(2406) <= not(layer2_outputs(2224));
    outputs(2407) <= not((layer2_outputs(2216)) and (layer2_outputs(1684)));
    outputs(2408) <= (layer2_outputs(1083)) and (layer2_outputs(811));
    outputs(2409) <= layer2_outputs(986);
    outputs(2410) <= layer2_outputs(870);
    outputs(2411) <= not((layer2_outputs(2209)) or (layer2_outputs(1874)));
    outputs(2412) <= not((layer2_outputs(1579)) and (layer2_outputs(1018)));
    outputs(2413) <= not(layer2_outputs(2107)) or (layer2_outputs(2486));
    outputs(2414) <= (layer2_outputs(454)) and not (layer2_outputs(549));
    outputs(2415) <= layer2_outputs(1639);
    outputs(2416) <= layer2_outputs(1450);
    outputs(2417) <= not(layer2_outputs(2225));
    outputs(2418) <= (layer2_outputs(1834)) and not (layer2_outputs(79));
    outputs(2419) <= not((layer2_outputs(1200)) or (layer2_outputs(2322)));
    outputs(2420) <= not(layer2_outputs(1924));
    outputs(2421) <= layer2_outputs(1599);
    outputs(2422) <= layer2_outputs(97);
    outputs(2423) <= (layer2_outputs(1795)) and not (layer2_outputs(1252));
    outputs(2424) <= not((layer2_outputs(1252)) or (layer2_outputs(527)));
    outputs(2425) <= (layer2_outputs(593)) and not (layer2_outputs(318));
    outputs(2426) <= not(layer2_outputs(595));
    outputs(2427) <= layer2_outputs(794);
    outputs(2428) <= not((layer2_outputs(1322)) xor (layer2_outputs(939)));
    outputs(2429) <= layer2_outputs(1052);
    outputs(2430) <= not((layer2_outputs(777)) or (layer2_outputs(556)));
    outputs(2431) <= (layer2_outputs(868)) and not (layer2_outputs(2241));
    outputs(2432) <= not(layer2_outputs(198));
    outputs(2433) <= not(layer2_outputs(2108)) or (layer2_outputs(271));
    outputs(2434) <= layer2_outputs(2447);
    outputs(2435) <= (layer2_outputs(806)) xor (layer2_outputs(1325));
    outputs(2436) <= not(layer2_outputs(2316));
    outputs(2437) <= not(layer2_outputs(1799));
    outputs(2438) <= layer2_outputs(1214);
    outputs(2439) <= not(layer2_outputs(2376));
    outputs(2440) <= (layer2_outputs(558)) and not (layer2_outputs(1285));
    outputs(2441) <= layer2_outputs(189);
    outputs(2442) <= not((layer2_outputs(1487)) or (layer2_outputs(2197)));
    outputs(2443) <= layer2_outputs(309);
    outputs(2444) <= not(layer2_outputs(2157));
    outputs(2445) <= (layer2_outputs(985)) and not (layer2_outputs(1558));
    outputs(2446) <= (layer2_outputs(512)) and (layer2_outputs(2126));
    outputs(2447) <= not(layer2_outputs(1390));
    outputs(2448) <= layer2_outputs(1710);
    outputs(2449) <= not(layer2_outputs(1085));
    outputs(2450) <= not(layer2_outputs(942));
    outputs(2451) <= not(layer2_outputs(719));
    outputs(2452) <= layer2_outputs(1409);
    outputs(2453) <= not((layer2_outputs(872)) or (layer2_outputs(2415)));
    outputs(2454) <= not(layer2_outputs(1177));
    outputs(2455) <= layer2_outputs(2309);
    outputs(2456) <= (layer2_outputs(621)) xor (layer2_outputs(407));
    outputs(2457) <= not(layer2_outputs(1924));
    outputs(2458) <= not((layer2_outputs(1284)) or (layer2_outputs(1170)));
    outputs(2459) <= (layer2_outputs(1165)) and not (layer2_outputs(1636));
    outputs(2460) <= not(layer2_outputs(2430));
    outputs(2461) <= not((layer2_outputs(1890)) xor (layer2_outputs(1836)));
    outputs(2462) <= layer2_outputs(1417);
    outputs(2463) <= (layer2_outputs(1769)) and not (layer2_outputs(799));
    outputs(2464) <= (layer2_outputs(2018)) and not (layer2_outputs(2532));
    outputs(2465) <= layer2_outputs(870);
    outputs(2466) <= not(layer2_outputs(2260));
    outputs(2467) <= layer2_outputs(732);
    outputs(2468) <= not((layer2_outputs(895)) or (layer2_outputs(1671)));
    outputs(2469) <= not(layer2_outputs(1682));
    outputs(2470) <= layer2_outputs(1453);
    outputs(2471) <= not(layer2_outputs(122));
    outputs(2472) <= not(layer2_outputs(378));
    outputs(2473) <= not(layer2_outputs(1844));
    outputs(2474) <= not((layer2_outputs(2142)) or (layer2_outputs(1313)));
    outputs(2475) <= not(layer2_outputs(2217)) or (layer2_outputs(196));
    outputs(2476) <= not(layer2_outputs(1986));
    outputs(2477) <= layer2_outputs(161);
    outputs(2478) <= not(layer2_outputs(1243));
    outputs(2479) <= not((layer2_outputs(837)) or (layer2_outputs(2047)));
    outputs(2480) <= layer2_outputs(1771);
    outputs(2481) <= not((layer2_outputs(1361)) and (layer2_outputs(515)));
    outputs(2482) <= not((layer2_outputs(689)) xor (layer2_outputs(1172)));
    outputs(2483) <= not(layer2_outputs(1523));
    outputs(2484) <= layer2_outputs(119);
    outputs(2485) <= (layer2_outputs(2452)) and not (layer2_outputs(1736));
    outputs(2486) <= layer2_outputs(128);
    outputs(2487) <= not(layer2_outputs(1760));
    outputs(2488) <= (layer2_outputs(1065)) or (layer2_outputs(310));
    outputs(2489) <= not(layer2_outputs(1844));
    outputs(2490) <= (layer2_outputs(2377)) and (layer2_outputs(117));
    outputs(2491) <= not(layer2_outputs(2549)) or (layer2_outputs(2123));
    outputs(2492) <= not(layer2_outputs(679));
    outputs(2493) <= layer2_outputs(2128);
    outputs(2494) <= (layer2_outputs(1988)) and not (layer2_outputs(756));
    outputs(2495) <= (layer2_outputs(1950)) or (layer2_outputs(1483));
    outputs(2496) <= layer2_outputs(567);
    outputs(2497) <= layer2_outputs(1766);
    outputs(2498) <= (layer2_outputs(692)) xor (layer2_outputs(1733));
    outputs(2499) <= not((layer2_outputs(942)) xor (layer2_outputs(2092)));
    outputs(2500) <= not(layer2_outputs(1947));
    outputs(2501) <= (layer2_outputs(2323)) and not (layer2_outputs(1383));
    outputs(2502) <= (layer2_outputs(1282)) and (layer2_outputs(1686));
    outputs(2503) <= not((layer2_outputs(1902)) or (layer2_outputs(2223)));
    outputs(2504) <= not((layer2_outputs(1983)) or (layer2_outputs(2530)));
    outputs(2505) <= layer2_outputs(2080);
    outputs(2506) <= (layer2_outputs(52)) xor (layer2_outputs(908));
    outputs(2507) <= (layer2_outputs(330)) and (layer2_outputs(321));
    outputs(2508) <= not(layer2_outputs(1070));
    outputs(2509) <= (layer2_outputs(2103)) and (layer2_outputs(116));
    outputs(2510) <= not(layer2_outputs(163));
    outputs(2511) <= (layer2_outputs(853)) and not (layer2_outputs(949));
    outputs(2512) <= not(layer2_outputs(1090));
    outputs(2513) <= not(layer2_outputs(2085));
    outputs(2514) <= not(layer2_outputs(327));
    outputs(2515) <= not(layer2_outputs(810));
    outputs(2516) <= (layer2_outputs(2503)) xor (layer2_outputs(1912));
    outputs(2517) <= not(layer2_outputs(1867));
    outputs(2518) <= (layer2_outputs(317)) xor (layer2_outputs(2434));
    outputs(2519) <= (layer2_outputs(2289)) and not (layer2_outputs(1261));
    outputs(2520) <= layer2_outputs(869);
    outputs(2521) <= not(layer2_outputs(1132));
    outputs(2522) <= not((layer2_outputs(293)) or (layer2_outputs(2254)));
    outputs(2523) <= not(layer2_outputs(1279));
    outputs(2524) <= not(layer2_outputs(2168));
    outputs(2525) <= not(layer2_outputs(1734));
    outputs(2526) <= (layer2_outputs(2139)) and not (layer2_outputs(438));
    outputs(2527) <= not(layer2_outputs(1809));
    outputs(2528) <= (layer2_outputs(2022)) xor (layer2_outputs(1524));
    outputs(2529) <= (layer2_outputs(868)) and not (layer2_outputs(2156));
    outputs(2530) <= not(layer2_outputs(322));
    outputs(2531) <= not(layer2_outputs(327));
    outputs(2532) <= layer2_outputs(1169);
    outputs(2533) <= (layer2_outputs(127)) and not (layer2_outputs(1585));
    outputs(2534) <= not(layer2_outputs(2046));
    outputs(2535) <= not((layer2_outputs(1460)) or (layer2_outputs(341)));
    outputs(2536) <= (layer2_outputs(903)) and not (layer2_outputs(1480));
    outputs(2537) <= not(layer2_outputs(693));
    outputs(2538) <= (layer2_outputs(1143)) xor (layer2_outputs(2000));
    outputs(2539) <= layer2_outputs(754);
    outputs(2540) <= layer2_outputs(1925);
    outputs(2541) <= not(layer2_outputs(1018));
    outputs(2542) <= layer2_outputs(626);
    outputs(2543) <= layer2_outputs(958);
    outputs(2544) <= not((layer2_outputs(2384)) or (layer2_outputs(801)));
    outputs(2545) <= not((layer2_outputs(2310)) xor (layer2_outputs(1557)));
    outputs(2546) <= not(layer2_outputs(18));
    outputs(2547) <= not(layer2_outputs(628));
    outputs(2548) <= (layer2_outputs(1791)) or (layer2_outputs(167));
    outputs(2549) <= not((layer2_outputs(2170)) or (layer2_outputs(544)));
    outputs(2550) <= (layer2_outputs(2382)) and not (layer2_outputs(67));
    outputs(2551) <= (layer2_outputs(728)) xor (layer2_outputs(1633));
    outputs(2552) <= layer2_outputs(495);
    outputs(2553) <= layer2_outputs(509);
    outputs(2554) <= layer2_outputs(1474);
    outputs(2555) <= not((layer2_outputs(1344)) or (layer2_outputs(1262)));
    outputs(2556) <= layer2_outputs(1310);
    outputs(2557) <= (layer2_outputs(2312)) xor (layer2_outputs(192));
    outputs(2558) <= (layer2_outputs(61)) and not (layer2_outputs(52));
    outputs(2559) <= layer2_outputs(1153);

end Behavioral;
